

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450;

  OAI22_X1 U7273 ( .A1(n13419), .A2(n13418), .B1(n13714), .B2(n8356), .ZN(
        n13407) );
  XNOR2_X1 U7274 ( .A(n11773), .B(n11771), .ZN(n12642) );
  NAND2_X1 U7275 ( .A1(n8199), .A2(n8198), .ZN(n13643) );
  INV_X1 U7276 ( .A(n12909), .ZN(n12883) );
  XNOR2_X1 U7277 ( .A(n15064), .B(n9876), .ZN(n11994) );
  AND4_X1 U7278 ( .A1(n9191), .A2(n9194), .A3(n9192), .A4(n9193), .ZN(n9252)
         );
  INV_X1 U7279 ( .A(n8899), .ZN(n8132) );
  INV_X1 U7280 ( .A(n7832), .ZN(n8133) );
  CLKBUF_X1 U7281 ( .A(n11974), .Z(n6533) );
  CLKBUF_X2 U7282 ( .A(n11974), .Z(n6531) );
  INV_X1 U7283 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  INV_X2 U7284 ( .A(n7645), .ZN(n6893) );
  NAND3_X1 U7285 ( .A1(n8440), .A2(n7205), .A3(n8400), .ZN(n8486) );
  OR2_X2 U7286 ( .A1(n8812), .A2(n14364), .ZN(n11583) );
  BUF_X2 U7287 ( .A(n12222), .Z(n6525) );
  NOR2_X1 U7288 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7705) );
  INV_X1 U7289 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8086) );
  NOR2_X1 U7290 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7704) );
  NAND2_X2 U7291 ( .A1(n9255), .A2(n9254), .ZN(n11789) );
  INV_X1 U7292 ( .A(n12525), .ZN(n12553) );
  INV_X1 U7293 ( .A(n11789), .ZN(n9489) );
  INV_X2 U7294 ( .A(n9489), .ZN(n11786) );
  OR2_X1 U7295 ( .A1(n11943), .A2(n11941), .ZN(n12833) );
  INV_X1 U7296 ( .A(n12854), .ZN(n12882) );
  INV_X1 U7297 ( .A(n11936), .ZN(n11955) );
  NAND2_X1 U7298 ( .A1(n9051), .A2(n11302), .ZN(n6534) );
  OR2_X1 U7299 ( .A1(n6537), .A2(n8445), .ZN(n7833) );
  BUF_X1 U7300 ( .A(n9574), .Z(n13542) );
  OAI211_X1 U7301 ( .C1(n8899), .C2(n8909), .A(n7878), .B(n7877), .ZN(n14936)
         );
  AND2_X1 U7302 ( .A1(n8306), .A2(n9718), .ZN(n12302) );
  AND4_X1 U7303 ( .A1(n7711), .A2(n8281), .A3(n8265), .A4(n7710), .ZN(n7712)
         );
  AND2_X1 U7304 ( .A1(n11581), .A2(n11580), .ZN(n14055) );
  INV_X1 U7305 ( .A(n14055), .ZN(n14284) );
  AND2_X1 U7306 ( .A1(n7134), .A2(n7133), .ZN(n6538) );
  OR2_X1 U7307 ( .A1(n8714), .A2(n8713), .ZN(n7702) );
  NAND2_X1 U7310 ( .A1(n8035), .A2(n8034), .ZN(n12139) );
  NAND2_X1 U7311 ( .A1(n7968), .A2(n7967), .ZN(n13601) );
  INV_X1 U7312 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7891) );
  INV_X2 U7313 ( .A(n14635), .ZN(n11352) );
  NAND2_X1 U7314 ( .A1(n8298), .A2(n8299), .ZN(n9718) );
  XNOR2_X1 U7315 ( .A(n7198), .B(n7197), .ZN(n11635) );
  INV_X1 U7316 ( .A(n12686), .ZN(P3_U3897) );
  NAND2_X2 U7317 ( .A1(n7638), .A2(n7636), .ZN(n13840) );
  AND4_X2 U7318 ( .A1(n9492), .A2(n9490), .A3(n9493), .A4(n9491), .ZN(n15047)
         );
  INV_X2 U7319 ( .A(n9019), .ZN(n12542) );
  NAND3_X2 U7320 ( .A1(n9718), .A2(n8302), .A3(n8301), .ZN(n7130) );
  AOI21_X2 U7321 ( .B1(n7831), .B2(n7830), .A(n7732), .ZN(n7848) );
  NAND4_X4 U7322 ( .A1(n8842), .A2(n8841), .A3(n8840), .A4(n8839), .ZN(n13955)
         );
  NAND2_X1 U7323 ( .A1(n12373), .A2(n7718), .ZN(n12222) );
  AOI21_X2 U7324 ( .B1(n10980), .B2(n10979), .A(n10978), .ZN(n10981) );
  INV_X1 U7326 ( .A(n11608), .ZN(n11489) );
  CLKBUF_X1 U7327 ( .A(n14708), .Z(n6526) );
  XNOR2_X1 U7328 ( .A(n6811), .B(n8612), .ZN(n14708) );
  XNOR2_X1 U7329 ( .A(n8131), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8306) );
  OAI21_X2 U7330 ( .B1(n8397), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8396) );
  INV_X2 U7331 ( .A(n11130), .ZN(n8812) );
  NAND4_X2 U7332 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(
        n12855) );
  OAI21_X2 U7333 ( .B1(n12834), .B2(n11943), .A(n11948), .ZN(n12820) );
  XNOR2_X2 U7334 ( .A(n8811), .B(n8810), .ZN(n14364) );
  NOR2_X2 U7335 ( .A1(n13172), .A2(n6571), .ZN(n9855) );
  OAI22_X2 U7336 ( .A1(n10303), .A2(n8321), .B1(n9863), .B2(n12091), .ZN(
        n10405) );
  NOR2_X4 U7337 ( .A1(n8486), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8543) );
  NOR2_X2 U7338 ( .A1(n11816), .A2(n11815), .ZN(n12907) );
  AND2_X2 U7340 ( .A1(n6956), .A2(n6955), .ZN(n11113) );
  NAND2_X2 U7341 ( .A1(n6794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7818) );
  AND2_X1 U7342 ( .A1(n14122), .A2(n11715), .ZN(n14109) );
  NAND2_X1 U7343 ( .A1(n13189), .A2(n13190), .ZN(n13161) );
  XNOR2_X1 U7344 ( .A(n12347), .B(n6698), .ZN(n6988) );
  OAI21_X1 U7345 ( .B1(n13479), .B2(n8351), .A(n8352), .ZN(n13461) );
  NAND2_X1 U7346 ( .A1(n13216), .A2(n12344), .ZN(n12347) );
  NAND2_X1 U7347 ( .A1(n8350), .A2(n8349), .ZN(n13479) );
  NAND2_X2 U7348 ( .A1(n11934), .A2(n11938), .ZN(n12868) );
  NAND2_X1 U7349 ( .A1(n11202), .A2(n11201), .ZN(n13079) );
  OAI21_X1 U7350 ( .B1(n6719), .B2(n14248), .A(n6717), .ZN(n14242) );
  OAI22_X1 U7351 ( .A1(n10803), .A2(n8030), .B1(n10897), .B2(n10567), .ZN(
        n10883) );
  XNOR2_X1 U7352 ( .A(n13672), .B(n6529), .ZN(n13206) );
  NAND2_X1 U7353 ( .A1(n6708), .A2(n6707), .ZN(n14999) );
  NAND2_X1 U7354 ( .A1(n10735), .A2(n10734), .ZN(n14258) );
  NAND2_X1 U7355 ( .A1(n8054), .A2(n8053), .ZN(n13696) );
  AND2_X1 U7356 ( .A1(n9516), .A2(n6805), .ZN(n9787) );
  INV_X1 U7357 ( .A(n11994), .ZN(n15044) );
  INV_X4 U7358 ( .A(n12542), .ZN(n12554) );
  INV_X1 U7359 ( .A(n14936), .ZN(n10182) );
  INV_X1 U7360 ( .A(n13267), .ZN(n7442) );
  INV_X1 U7361 ( .A(n13952), .ZN(n9781) );
  NOR2_X2 U7362 ( .A1(n9564), .A2(n15063), .ZN(n15061) );
  INV_X1 U7363 ( .A(n13269), .ZN(n6940) );
  INV_X1 U7364 ( .A(n11372), .ZN(n11374) );
  BUF_X1 U7365 ( .A(n9565), .Z(n14901) );
  INV_X2 U7366 ( .A(n11348), .ZN(n11373) );
  AND2_X1 U7367 ( .A1(n8825), .A2(n9746), .ZN(n9019) );
  NAND4_X1 U7368 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n13957)
         );
  CLKBUF_X2 U7369 ( .A(n11626), .Z(n6963) );
  INV_X1 U7370 ( .A(n9432), .ZN(n9564) );
  AND2_X2 U7371 ( .A1(n12302), .A2(n10418), .ZN(n14943) );
  CLKBUF_X2 U7372 ( .A(n11564), .Z(n11582) );
  CLKBUF_X1 U7373 ( .A(n11623), .Z(n6987) );
  NAND2_X1 U7374 ( .A1(n11633), .A2(n11635), .ZN(n11365) );
  CLKBUF_X2 U7376 ( .A(n11974), .Z(n6532) );
  INV_X2 U7377 ( .A(n11516), .ZN(n11455) );
  NAND2_X1 U7378 ( .A1(n14374), .A2(n14635), .ZN(n11307) );
  NAND2_X2 U7379 ( .A1(n9051), .A2(n11302), .ZN(n10868) );
  OAI21_X1 U7380 ( .B1(n9159), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6939), .ZN(
        n7731) );
  INV_X2 U7381 ( .A(n9159), .ZN(n9161) );
  CLKBUF_X3 U7382 ( .A(n6538), .Z(n6536) );
  AND2_X1 U7383 ( .A1(n7134), .A2(n7133), .ZN(n9159) );
  NOR2_X2 U7384 ( .A1(n7377), .A2(n8429), .ZN(n7199) );
  AND4_X1 U7385 ( .A1(n8380), .A2(n8379), .A3(n8378), .A4(n8377), .ZN(n9278)
         );
  CLKBUF_X2 U7386 ( .A(n8440), .Z(n9065) );
  AND3_X2 U7387 ( .A1(n8090), .A2(n8086), .A3(n7485), .ZN(n6651) );
  INV_X2 U7388 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7389 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8392) );
  NOR2_X1 U7390 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8377) );
  NOR2_X1 U7391 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8378) );
  NOR2_X1 U7392 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8379) );
  AND2_X1 U7393 ( .A1(n6898), .A2(n6897), .ZN(n14287) );
  AND2_X1 U7394 ( .A1(n6985), .A2(n14286), .ZN(n6984) );
  AOI21_X1 U7395 ( .B1(n13407), .B2(n12297), .A(n7288), .ZN(n8262) );
  OAI22_X1 U7396 ( .A1(n11605), .A2(n6759), .B1(n6758), .B2(n11604), .ZN(
        n11616) );
  OAI21_X1 U7397 ( .B1(n7361), .B2(n7360), .A(n7266), .ZN(n7265) );
  AND2_X1 U7398 ( .A1(n7145), .A2(n7144), .ZN(n13618) );
  AOI21_X1 U7399 ( .B1(n7235), .B2(n7237), .A(n7234), .ZN(n7233) );
  AOI21_X1 U7400 ( .B1(n14073), .B2(n14494), .A(n14072), .ZN(n14282) );
  XNOR2_X1 U7401 ( .A(n14067), .B(n14075), .ZN(n14073) );
  NAND2_X1 U7402 ( .A1(n12808), .A2(n12812), .ZN(n12807) );
  OAI21_X1 U7403 ( .B1(n7666), .B2(n12193), .A(n7216), .ZN(n6919) );
  NAND2_X1 U7404 ( .A1(n13161), .A2(n12351), .ZN(n6696) );
  AOI21_X1 U7405 ( .B1(n7411), .B2(n7414), .A(n6631), .ZN(n7409) );
  NAND2_X1 U7406 ( .A1(n6575), .A2(n7667), .ZN(n7666) );
  NOR2_X1 U7407 ( .A1(n6727), .A2(n6726), .ZN(n14067) );
  NAND2_X1 U7408 ( .A1(n14309), .A2(n7333), .ZN(n14122) );
  AND2_X1 U7409 ( .A1(n7412), .A2(n6645), .ZN(n7411) );
  NAND2_X1 U7410 ( .A1(n13134), .A2(n12348), .ZN(n13189) );
  AOI21_X1 U7411 ( .B1(n7415), .B2(n7413), .A(n6639), .ZN(n7412) );
  NAND2_X1 U7412 ( .A1(n13493), .A2(n8182), .ZN(n13477) );
  NAND2_X1 U7413 ( .A1(n11330), .A2(n11329), .ZN(n14032) );
  AND2_X1 U7414 ( .A1(n14081), .A2(n6584), .ZN(n14279) );
  NOR3_X1 U7415 ( .A1(n14080), .A2(n14039), .A3(n6821), .ZN(n14035) );
  NAND2_X1 U7416 ( .A1(n6988), .A2(n6676), .ZN(n13134) );
  AND2_X1 U7417 ( .A1(n7418), .A2(n7416), .ZN(n7415) );
  OAI21_X1 U7418 ( .B1(n11286), .B2(n6879), .A(n6877), .ZN(n6885) );
  NAND2_X1 U7419 ( .A1(n7419), .A2(n7420), .ZN(n7418) );
  NAND2_X1 U7420 ( .A1(n12233), .A2(n12232), .ZN(n13396) );
  NAND2_X1 U7421 ( .A1(n14103), .A2(n14102), .ZN(n14101) );
  AOI21_X1 U7422 ( .B1(n6880), .B2(n6878), .A(n6644), .ZN(n6877) );
  INV_X1 U7423 ( .A(n6880), .ZN(n6879) );
  INV_X1 U7424 ( .A(n12294), .ZN(n13432) );
  AND2_X1 U7425 ( .A1(n13409), .A2(n13241), .ZN(n7288) );
  XNOR2_X1 U7426 ( .A(n11129), .B(n11128), .ZN(n12231) );
  CLKBUF_X1 U7427 ( .A(n13790), .Z(n13896) );
  NAND2_X1 U7428 ( .A1(n8239), .A2(n8238), .ZN(n13409) );
  NOR2_X1 U7429 ( .A1(n14118), .A2(n11714), .ZN(n14117) );
  NOR2_X1 U7430 ( .A1(n13457), .A2(n8355), .ZN(n7439) );
  NAND2_X1 U7431 ( .A1(n8254), .A2(n8253), .ZN(n13616) );
  NAND2_X1 U7432 ( .A1(n7111), .A2(n7110), .ZN(n13216) );
  OR2_X1 U7433 ( .A1(n12197), .A2(n7217), .ZN(n7216) );
  OAI211_X1 U7434 ( .C1(n7820), .C2(n7139), .A(n7136), .B(n7135), .ZN(n12294)
         );
  OAI21_X1 U7435 ( .B1(n11269), .B2(n11146), .A(n11147), .ZN(n11273) );
  AOI21_X1 U7436 ( .B1(n7294), .B2(n8193), .A(n6598), .ZN(n7293) );
  NAND2_X1 U7437 ( .A1(n8226), .A2(n8225), .ZN(n13424) );
  AND2_X1 U7438 ( .A1(n11946), .A2(n11942), .ZN(n12850) );
  NAND2_X1 U7439 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  CLKBUF_X1 U7440 ( .A(n13555), .Z(n6967) );
  NAND2_X1 U7441 ( .A1(n11125), .A2(n11124), .ZN(n11321) );
  XNOR2_X1 U7442 ( .A(n11125), .B(n11124), .ZN(n12371) );
  XNOR2_X1 U7443 ( .A(n8250), .B(n8249), .ZN(n13756) );
  OAI22_X1 U7444 ( .A1(n12176), .A2(n6804), .B1(n12175), .B2(n12174), .ZN(
        n7674) );
  NAND2_X1 U7445 ( .A1(n8209), .A2(n8208), .ZN(n13638) );
  NAND2_X1 U7446 ( .A1(n11561), .A2(n11560), .ZN(n14293) );
  AND2_X1 U7447 ( .A1(n7814), .A2(n8223), .ZN(n13763) );
  XNOR2_X1 U7448 ( .A(n8234), .B(n8224), .ZN(n13760) );
  NOR2_X2 U7449 ( .A1(n14201), .A2(n11699), .ZN(n14182) );
  AND2_X1 U7450 ( .A1(n8342), .A2(n8341), .ZN(n13537) );
  NAND2_X1 U7451 ( .A1(n11539), .A2(n11538), .ZN(n14301) );
  AOI21_X1 U7452 ( .B1(n6542), .B2(n7193), .A(n7188), .ZN(n7187) );
  INV_X1 U7453 ( .A(n12879), .ZN(n12886) );
  NAND2_X1 U7454 ( .A1(n11235), .A2(n11234), .ZN(n13008) );
  NAND2_X1 U7455 ( .A1(n7093), .A2(n10798), .ZN(n11142) );
  NAND2_X1 U7456 ( .A1(n8223), .A2(n8222), .ZN(n8234) );
  NAND2_X1 U7457 ( .A1(n7149), .A2(n7148), .ZN(n8223) );
  XNOR2_X1 U7458 ( .A(n8207), .B(n8206), .ZN(n11559) );
  XNOR2_X1 U7459 ( .A(n13012), .B(n12872), .ZN(n12879) );
  OAI21_X1 U7460 ( .B1(n11098), .B2(n7445), .A(n7443), .ZN(n13549) );
  AND2_X1 U7461 ( .A1(n8197), .A2(n8196), .ZN(n11537) );
  AOI21_X1 U7462 ( .B1(n7479), .B2(n6610), .A(n7126), .ZN(n7125) );
  NAND2_X1 U7463 ( .A1(n8197), .A2(n7809), .ZN(n8207) );
  NAND2_X1 U7464 ( .A1(n8197), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U7465 ( .A1(n8185), .A2(n8184), .ZN(n13648) );
  OR2_X1 U7466 ( .A1(n8195), .A2(n8194), .ZN(n8197) );
  AOI21_X1 U7467 ( .B1(n6906), .B2(n12331), .A(n6623), .ZN(n7479) );
  AND2_X1 U7468 ( .A1(n7809), .A2(n7151), .ZN(n7150) );
  OR2_X1 U7469 ( .A1(n10992), .A2(n8333), .ZN(n8335) );
  NAND2_X1 U7470 ( .A1(n7807), .A2(SI_24_), .ZN(n7809) );
  OR2_X1 U7471 ( .A1(n7807), .A2(SI_24_), .ZN(n7808) );
  AND2_X1 U7472 ( .A1(n13229), .A2(n12326), .ZN(n7481) );
  OAI21_X1 U7473 ( .B1(n8170), .B2(n7170), .A(n7166), .ZN(n7807) );
  INV_X1 U7474 ( .A(n7167), .ZN(n7166) );
  OAI21_X1 U7475 ( .B1(n14567), .B2(n11895), .A(n11893), .ZN(n11017) );
  OR2_X1 U7476 ( .A1(n14812), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U7477 ( .A1(n11340), .A2(n11339), .ZN(n14337) );
  NAND2_X1 U7478 ( .A1(n8115), .A2(n8114), .ZN(n13735) );
  NAND2_X1 U7479 ( .A1(n10818), .A2(n6548), .ZN(n13571) );
  NAND2_X1 U7480 ( .A1(n11354), .A2(n11353), .ZN(n14332) );
  AOI21_X1 U7481 ( .B1(n7386), .B2(n10736), .A(n7385), .ZN(n7384) );
  XNOR2_X1 U7482 ( .A(n9833), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9831) );
  OR2_X1 U7483 ( .A1(n11338), .A2(n8171), .ZN(n8115) );
  NAND2_X1 U7484 ( .A1(n10676), .A2(n8325), .ZN(n10771) );
  OR2_X1 U7485 ( .A1(n10572), .A2(n10571), .ZN(n6957) );
  NOR2_X1 U7486 ( .A1(n13696), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U7487 ( .A1(n14573), .A2(n11887), .ZN(n12980) );
  NOR2_X2 U7488 ( .A1(n14623), .A2(n14645), .ZN(n14622) );
  NAND2_X1 U7489 ( .A1(n7498), .A2(n7497), .ZN(n14623) );
  NAND2_X1 U7490 ( .A1(n14999), .A2(n6603), .ZN(n14573) );
  NAND2_X1 U7491 ( .A1(n8158), .A2(n7801), .ZN(n7802) );
  AND2_X2 U7492 ( .A1(n11430), .A2(n11431), .ZN(n14260) );
  OR2_X1 U7493 ( .A1(n14258), .A2(n13882), .ZN(n11430) );
  NOR2_X1 U7494 ( .A1(n12139), .A2(n14819), .ZN(n7369) );
  OAI21_X1 U7495 ( .B1(n10916), .B2(n10915), .A(n12679), .ZN(n10918) );
  NAND2_X1 U7496 ( .A1(n8094), .A2(n8093), .ZN(n13739) );
  AOI21_X1 U7497 ( .B1(n7407), .B2(n10235), .A(n7406), .ZN(n7405) );
  AND2_X1 U7498 ( .A1(n10596), .A2(n10595), .ZN(n14506) );
  NOR2_X1 U7499 ( .A1(n11656), .A2(n7400), .ZN(n7407) );
  XNOR2_X1 U7500 ( .A(n8046), .B(n8045), .ZN(n10732) );
  OR2_X1 U7501 ( .A1(n7131), .A2(n11187), .ZN(n7798) );
  XNOR2_X1 U7502 ( .A(n6981), .B(n8048), .ZN(n10737) );
  AOI21_X1 U7503 ( .B1(n8083), .B2(n7788), .A(n6633), .ZN(n7131) );
  NAND2_X1 U7504 ( .A1(n10601), .A2(n10600), .ZN(n14666) );
  NAND2_X1 U7505 ( .A1(n6825), .A2(n6824), .ZN(n10360) );
  INV_X1 U7506 ( .A(n6713), .ZN(n6981) );
  OAI21_X1 U7507 ( .B1(n8031), .B2(n6716), .A(n6712), .ZN(n8046) );
  NAND2_X1 U7508 ( .A1(n10423), .A2(n11862), .ZN(n10904) );
  NAND2_X1 U7509 ( .A1(n10348), .A2(n10347), .ZN(n14672) );
  INV_X1 U7510 ( .A(n10223), .ZN(n6825) );
  NAND2_X1 U7511 ( .A1(n10051), .A2(n14784), .ZN(n10223) );
  OR2_X1 U7512 ( .A1(n11261), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11263) );
  XNOR2_X1 U7513 ( .A(n7982), .B(n7981), .ZN(n10345) );
  NAND2_X1 U7514 ( .A1(n10027), .A2(n10026), .ZN(n11413) );
  AND2_X1 U7515 ( .A1(n7978), .A2(n7977), .ZN(n7982) );
  OAI21_X1 U7516 ( .B1(n7978), .B2(n7157), .A(n7155), .ZN(n8016) );
  NAND2_X1 U7517 ( .A1(n7951), .A2(n7950), .ZN(n12103) );
  NAND2_X1 U7518 ( .A1(n7961), .A2(n7758), .ZN(n7978) );
  NAND2_X1 U7519 ( .A1(n7945), .A2(n7756), .ZN(n7961) );
  NAND2_X1 U7520 ( .A1(n7920), .A2(n7919), .ZN(n12091) );
  NAND2_X1 U7521 ( .A1(n6722), .A2(n7755), .ZN(n7945) );
  OR2_X1 U7522 ( .A1(n11984), .A2(n6705), .ZN(n6704) );
  NOR2_X2 U7523 ( .A1(n13915), .A2(n14631), .ZN(n8890) );
  OR2_X1 U7524 ( .A1(n12074), .A2(n12073), .ZN(n6786) );
  INV_X2 U7525 ( .A(n14797), .ZN(n6528) );
  AND2_X1 U7526 ( .A1(n6997), .A2(n6996), .ZN(n8903) );
  NAND2_X1 U7527 ( .A1(n7898), .A2(n7746), .ZN(n7915) );
  NAND2_X1 U7528 ( .A1(n9744), .A2(n9743), .ZN(n14758) );
  NAND2_X1 U7529 ( .A1(n7745), .A2(n7744), .ZN(n7898) );
  AND4_X1 U7530 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n11386)
         );
  INV_X1 U7531 ( .A(n14752), .ZN(n7537) );
  NAND2_X1 U7532 ( .A1(n6576), .A2(n7841), .ZN(n13267) );
  NAND4_X1 U7533 ( .A1(n9157), .A2(n9155), .A3(n9158), .A4(n9156), .ZN(n15063)
         );
  NAND4_X1 U7534 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n15064)
         );
  INV_X4 U7535 ( .A(n12356), .ZN(n6529) );
  AND2_X1 U7536 ( .A1(n8879), .A2(n6819), .ZN(n14752) );
  AND2_X1 U7537 ( .A1(n6815), .A2(n9349), .ZN(n14737) );
  INV_X2 U7538 ( .A(n12213), .ZN(n12070) );
  NAND2_X1 U7539 ( .A1(n9224), .A2(n9223), .ZN(n14494) );
  AND2_X1 U7540 ( .A1(n7007), .A2(n7006), .ZN(n8985) );
  OR2_X2 U7541 ( .A1(n11331), .A2(n11633), .ZN(n14674) );
  NAND2_X1 U7542 ( .A1(n8825), .A2(n11365), .ZN(n12543) );
  AND2_X1 U7543 ( .A1(n8419), .A2(n6589), .ZN(n10581) );
  NAND2_X2 U7544 ( .A1(n8812), .A2(n8814), .ZN(n11608) );
  NAND2_X2 U7545 ( .A1(n8812), .A2(n14364), .ZN(n11630) );
  BUF_X2 U7546 ( .A(n9678), .Z(n11216) );
  OR3_X2 U7547 ( .A1(n11799), .A2(n14368), .A3(n11063), .ZN(n8825) );
  INV_X1 U7548 ( .A(n13118), .ZN(n8715) );
  AND2_X1 U7549 ( .A1(n11130), .A2(n14364), .ZN(n11564) );
  XNOR2_X1 U7550 ( .A(n8389), .B(n8388), .ZN(n11799) );
  NAND2_X1 U7551 ( .A1(n7722), .A2(n12375), .ZN(n7857) );
  NAND2_X1 U7552 ( .A1(n8803), .A2(n6730), .ZN(n14635) );
  NAND2_X1 U7553 ( .A1(n8712), .A2(n13111), .ZN(n13118) );
  NAND2_X1 U7554 ( .A1(n8803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7198) );
  NAND3_X1 U7555 ( .A1(n7307), .A2(n7306), .A3(n7308), .ZN(n11130) );
  OAI21_X1 U7556 ( .B1(n8387), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8389) );
  XNOR2_X1 U7557 ( .A(n8304), .B(n8303), .ZN(n10418) );
  NAND2_X1 U7558 ( .A1(n7483), .A2(n7482), .ZN(n8298) );
  MUX2_X1 U7559 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8300), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8301) );
  XNOR2_X1 U7560 ( .A(n8601), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14374) );
  XNOR2_X1 U7561 ( .A(n7716), .B(n7715), .ZN(n12373) );
  NAND2_X1 U7562 ( .A1(n8614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U7563 ( .A1(n8800), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8802) );
  AND4_X1 U7564 ( .A1(n7530), .A2(n7215), .A3(n8543), .A4(n6664), .ZN(n8714)
         );
  AND2_X1 U7565 ( .A1(n8412), .A2(n7257), .ZN(n7215) );
  AND2_X1 U7566 ( .A1(n8407), .A2(n7531), .ZN(n7530) );
  AND3_X1 U7567 ( .A1(n7694), .A2(n7693), .A3(n8408), .ZN(n7531) );
  NOR2_X1 U7568 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  AND2_X1 U7569 ( .A1(n8414), .A2(n8411), .ZN(n8412) );
  AND2_X2 U7570 ( .A1(n9278), .A2(n6563), .ZN(n8611) );
  NAND4_X1 U7571 ( .A1(n14523), .A2(n15357), .A3(P1_ADDR_REG_19__SCAN_IN), 
        .A4(P2_ADDR_REG_19__SCAN_IN), .ZN(n7133) );
  NAND4_X1 U7572 ( .A1(n15392), .A2(n7728), .A3(n15356), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7134) );
  AND3_X1 U7573 ( .A1(n9054), .A2(n9178), .A3(n9053), .ZN(n7694) );
  AND3_X1 U7574 ( .A1(n8417), .A2(n8410), .A3(n6908), .ZN(n8414) );
  INV_X4 U7575 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7576 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8265) );
  NOR2_X1 U7577 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7708) );
  INV_X1 U7578 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8400) );
  NOR2_X2 U7579 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7205) );
  INV_X1 U7580 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8417) );
  INV_X1 U7581 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8516) );
  INV_X1 U7582 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8544) );
  INV_X1 U7583 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9053) );
  INV_X1 U7584 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9054) );
  INV_X1 U7585 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8583) );
  NOR2_X1 U7586 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8401) );
  NOR2_X1 U7587 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8402) );
  INV_X1 U7588 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8537) );
  INV_X4 U7589 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7590 ( .A1(n12820), .A2(n12826), .ZN(n12810) );
  NOR2_X2 U7591 ( .A1(n13420), .A2(n13409), .ZN(n7374) );
  AOI21_X2 U7592 ( .B1(n12810), .B2(n11954), .A(n11953), .ZN(n12020) );
  AND4_X2 U7593 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n11847)
         );
  XNOR2_X1 U7594 ( .A(n10287), .B(n12679), .ZN(n10286) );
  BUF_X8 U7595 ( .A(n10084), .Z(n6530) );
  AND2_X1 U7596 ( .A1(n12569), .A2(n13118), .ZN(n11974) );
  NOR2_X2 U7597 ( .A1(n11263), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10313) );
  NOR2_X2 U7598 ( .A1(n13527), .A2(n13512), .ZN(n7371) );
  NAND2_X4 U7599 ( .A1(n14943), .A2(n12301), .ZN(n12213) );
  NOR4_X2 U7600 ( .A1(n12021), .A2(n12018), .A3(n12011), .A4(n12010), .ZN(
        n12012) );
  OAI222_X1 U7602 ( .A1(n13764), .A2(n8445), .B1(n13766), .B2(n8875), .C1(
        P2_U3088), .C2(n13271), .ZN(P2_U3326) );
  OAI222_X1 U7603 ( .A1(n14372), .A2(n8876), .B1(n14370), .B2(n8875), .C1(
        P1_U3086), .C2(n6931), .ZN(P1_U3354) );
  XNOR2_X1 U7604 ( .A(n7831), .B(n7830), .ZN(n8875) );
  NAND2_X1 U7605 ( .A1(n8899), .A2(n6536), .ZN(n8171) );
  NAND2_X1 U7606 ( .A1(n8899), .A2(n9161), .ZN(n6537) );
  INV_X2 U7607 ( .A(n12053), .ZN(n9451) );
  XNOR2_X1 U7608 ( .A(n12356), .B(n12053), .ZN(n9376) );
  INV_X1 U7609 ( .A(n12143), .ZN(n7660) );
  INV_X1 U7610 ( .A(n12142), .ZN(n7661) );
  INV_X1 U7611 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n6908) );
  INV_X1 U7612 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8403) );
  INV_X1 U7613 ( .A(n14627), .ZN(n7382) );
  OAI21_X1 U7614 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14404), .A(n14403), .ZN(
        n14465) );
  NAND2_X1 U7615 ( .A1(n6837), .A2(n11031), .ZN(n11279) );
  NAND2_X1 U7616 ( .A1(n9035), .A2(n9034), .ZN(n9037) );
  NOR2_X1 U7617 ( .A1(n7416), .A2(n7336), .ZN(n7335) );
  INV_X1 U7618 ( .A(n7339), .ZN(n7336) );
  NAND2_X1 U7619 ( .A1(n7105), .A2(n6754), .ZN(n7462) );
  INV_X1 U7620 ( .A(n12075), .ZN(n6788) );
  NAND2_X1 U7621 ( .A1(n12074), .A2(n12073), .ZN(n6787) );
  NAND2_X1 U7622 ( .A1(n7548), .A2(n11424), .ZN(n7547) );
  NAND2_X1 U7623 ( .A1(n7659), .A2(n7662), .ZN(n7654) );
  INV_X1 U7624 ( .A(n12120), .ZN(n7662) );
  AOI21_X1 U7625 ( .B1(n6972), .B2(n6605), .A(n6742), .ZN(n11503) );
  NOR2_X1 U7626 ( .A1(n11485), .A2(n11486), .ZN(n6742) );
  INV_X1 U7627 ( .A(n12183), .ZN(n6774) );
  INV_X1 U7628 ( .A(n12187), .ZN(n6936) );
  NOR2_X1 U7629 ( .A1(n8047), .A2(n7779), .ZN(n7780) );
  NAND2_X1 U7630 ( .A1(n12227), .A2(n7232), .ZN(n7231) );
  NOR2_X1 U7631 ( .A1(n6570), .A2(n7241), .ZN(n7240) );
  NAND2_X1 U7632 ( .A1(n14289), .A2(n13828), .ZN(n7420) );
  NAND2_X1 U7633 ( .A1(n7775), .A2(n8694), .ZN(n7781) );
  INV_X1 U7634 ( .A(n12855), .ZN(n11784) );
  INV_X1 U7635 ( .A(n15000), .ZN(n11882) );
  NOR2_X1 U7636 ( .A1(n9111), .A2(n6583), .ZN(n9089) );
  AOI21_X1 U7637 ( .B1(n12784), .B2(n12783), .A(n6691), .ZN(n12787) );
  NAND2_X1 U7638 ( .A1(n6865), .A2(n6864), .ZN(n6870) );
  AND2_X1 U7639 ( .A1(n6646), .A2(n11814), .ZN(n6864) );
  AND3_X1 U7640 ( .A1(n9990), .A2(n9989), .A3(n9988), .ZN(n10110) );
  NAND2_X1 U7641 ( .A1(n11286), .A2(n6883), .ZN(n6882) );
  NOR2_X1 U7642 ( .A1(n14568), .A2(n7201), .ZN(n7200) );
  INV_X1 U7643 ( .A(n10931), .ZN(n7201) );
  NAND2_X1 U7644 ( .A1(n7203), .A2(n7202), .ZN(n12974) );
  NAND2_X1 U7645 ( .A1(n6543), .A2(n6568), .ZN(n7202) );
  NAND2_X1 U7646 ( .A1(n7250), .A2(n7252), .ZN(n14997) );
  AND2_X1 U7647 ( .A1(n10906), .A2(n7253), .ZN(n7252) );
  NAND2_X1 U7648 ( .A1(n8626), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U7649 ( .A1(n8598), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U7650 ( .A1(n15259), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U7651 ( .A1(n8555), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8461) );
  INV_X1 U7652 ( .A(n7438), .ZN(n7436) );
  NAND2_X1 U7653 ( .A1(n13243), .A2(n7138), .ZN(n7135) );
  NOR2_X1 U7654 ( .A1(n13243), .A2(n7138), .ZN(n7137) );
  AND2_X1 U7655 ( .A1(n7282), .A2(n6647), .ZN(n7280) );
  NAND2_X1 U7656 ( .A1(n8337), .A2(n7446), .ZN(n7445) );
  NAND2_X1 U7657 ( .A1(n12283), .A2(n8336), .ZN(n7446) );
  NAND2_X1 U7658 ( .A1(n6940), .A2(n12053), .ZN(n8311) );
  INV_X1 U7659 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7815) );
  AND2_X2 U7660 ( .A1(n8049), .A2(n7708), .ZN(n7676) );
  INV_X1 U7661 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7710) );
  OR2_X1 U7662 ( .A1(n8302), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8280) );
  INV_X1 U7663 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6791) );
  INV_X1 U7664 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6790) );
  INV_X1 U7665 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6789) );
  OAI21_X1 U7666 ( .B1(n7183), .B2(n7181), .A(n6682), .ZN(n7180) );
  INV_X1 U7667 ( .A(n13879), .ZN(n7181) );
  INV_X1 U7668 ( .A(n12543), .ZN(n7196) );
  NOR2_X1 U7669 ( .A1(n11707), .A2(n11663), .ZN(n7342) );
  NAND2_X1 U7670 ( .A1(n10739), .A2(n6720), .ZN(n11693) );
  AND2_X1 U7671 ( .A1(n13942), .A2(n10738), .ZN(n6720) );
  NAND2_X1 U7672 ( .A1(n11516), .A2(n6536), .ZN(n11623) );
  NAND2_X1 U7673 ( .A1(n8252), .A2(n8251), .ZN(n11125) );
  INV_X1 U7674 ( .A(n7600), .ZN(n7599) );
  AOI21_X1 U7675 ( .B1(n7602), .B2(n7600), .A(n7598), .ZN(n7597) );
  AND2_X1 U7676 ( .A1(n8082), .A2(n7789), .ZN(n7788) );
  OR2_X1 U7677 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  AND2_X1 U7678 ( .A1(n7770), .A2(n7769), .ZN(n7996) );
  XNOR2_X1 U7679 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n6753) );
  NAND2_X1 U7680 ( .A1(n9496), .A2(n9497), .ZN(n7018) );
  AOI21_X1 U7681 ( .B1(n7039), .B2(n7036), .A(n6630), .ZN(n7035) );
  INV_X1 U7682 ( .A(n11752), .ZN(n7036) );
  AND2_X1 U7683 ( .A1(n11882), .A2(n10708), .ZN(n7534) );
  OR2_X1 U7684 ( .A1(n10689), .A2(n6659), .ZN(n7028) );
  INV_X1 U7685 ( .A(n12019), .ZN(n7360) );
  NOR2_X1 U7686 ( .A1(n12018), .A2(n12017), .ZN(n7266) );
  BUF_X1 U7687 ( .A(n9678), .Z(n6944) );
  AND4_X1 U7688 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n12656) );
  NAND2_X1 U7689 ( .A1(n10868), .A2(n6536), .ZN(n9484) );
  OR2_X1 U7690 ( .A1(n13073), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U7691 ( .A1(n12944), .A2(n11822), .ZN(n7261) );
  NAND2_X1 U7692 ( .A1(n6838), .A2(n11030), .ZN(n11039) );
  INV_X1 U7693 ( .A(n11198), .ZN(n11971) );
  AND2_X1 U7694 ( .A1(n9884), .A2(n11955), .ZN(n15062) );
  INV_X1 U7695 ( .A(n9051), .ZN(n12710) );
  INV_X1 U7696 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8411) );
  AND2_X1 U7697 ( .A1(n15368), .A2(n8409), .ZN(n7693) );
  XNOR2_X1 U7698 ( .A(n9181), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12771) );
  NOR2_X1 U7699 ( .A1(n9214), .A2(n7079), .ZN(n7078) );
  INV_X1 U7700 ( .A(n9212), .ZN(n7079) );
  OAI21_X1 U7701 ( .B1(n8690), .B2(n8689), .A(n8691), .ZN(n8864) );
  NAND2_X1 U7702 ( .A1(n8553), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8458) );
  AND2_X1 U7703 ( .A1(n13266), .A2(n9574), .ZN(n9567) );
  NAND2_X1 U7704 ( .A1(n10378), .A2(n11807), .ZN(n11813) );
  INV_X1 U7705 ( .A(n12299), .ZN(n7147) );
  INV_X1 U7706 ( .A(n12297), .ZN(n13406) );
  NAND2_X1 U7707 ( .A1(n13461), .A2(n13464), .ZN(n8354) );
  INV_X1 U7708 ( .A(n7452), .ZN(n7451) );
  OAI22_X1 U7709 ( .A1(n6565), .A2(n7453), .B1(n13512), .B2(n8347), .ZN(n7452)
         );
  NAND2_X1 U7710 ( .A1(n6640), .A2(n8346), .ZN(n7453) );
  OR2_X1 U7711 ( .A1(n10405), .A2(n8322), .ZN(n7458) );
  NAND2_X1 U7712 ( .A1(n13753), .A2(n12230), .ZN(n7583) );
  OR3_X1 U7713 ( .A1(n13767), .A2(n10954), .A3(n11061), .ZN(n9329) );
  OR2_X1 U7714 ( .A1(n7675), .A2(n7486), .ZN(n7714) );
  INV_X1 U7715 ( .A(n13862), .ZN(n7625) );
  AOI21_X1 U7716 ( .B1(n13862), .B2(n7624), .A(n7623), .ZN(n7622) );
  INV_X1 U7717 ( .A(n13834), .ZN(n7623) );
  NAND2_X1 U7718 ( .A1(n7609), .A2(n7607), .ZN(n10839) );
  NAND2_X1 U7719 ( .A1(n7612), .A2(n7608), .ZN(n7607) );
  NAND2_X1 U7720 ( .A1(n11626), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8842) );
  INV_X1 U7721 ( .A(n14364), .ZN(n8814) );
  NAND2_X1 U7722 ( .A1(n7338), .A2(n6591), .ZN(n14074) );
  NAND2_X1 U7723 ( .A1(n14192), .A2(n7331), .ZN(n14174) );
  NOR2_X1 U7724 ( .A1(n7398), .A2(n7332), .ZN(n7331) );
  INV_X1 U7725 ( .A(n11709), .ZN(n7332) );
  NAND2_X1 U7726 ( .A1(n14209), .A2(n14325), .ZN(n14188) );
  INV_X1 U7727 ( .A(n6718), .ZN(n6717) );
  OAI21_X1 U7728 ( .B1(n6719), .B2(n7386), .A(n11696), .ZN(n6718) );
  NAND2_X1 U7729 ( .A1(n14622), .A2(n14240), .ZN(n14235) );
  INV_X1 U7730 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7380) );
  INV_X1 U7731 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7379) );
  INV_X1 U7732 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U7733 ( .A1(n8802), .A2(n8801), .ZN(n8803) );
  AND2_X1 U7734 ( .A1(n6752), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14433) );
  INV_X1 U7735 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6752) );
  INV_X1 U7736 ( .A(n6744), .ZN(n14445) );
  OAI21_X1 U7737 ( .B1(n15438), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6616), .ZN(
        n6744) );
  INV_X1 U7738 ( .A(n14698), .ZN(n6754) );
  NAND2_X2 U7739 ( .A1(n8307), .A2(n14916), .ZN(n13595) );
  NAND2_X1 U7740 ( .A1(n14287), .A2(n6984), .ZN(n14352) );
  OAI21_X1 U7741 ( .B1(n14696), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6572), .ZN(
        n7105) );
  NAND2_X1 U7742 ( .A1(n12042), .A2(n12213), .ZN(n12048) );
  AOI21_X1 U7743 ( .B1(n6769), .B2(n12056), .A(n12054), .ZN(n12055) );
  NOR2_X1 U7744 ( .A1(n6769), .A2(n12056), .ZN(n12057) );
  INV_X1 U7745 ( .A(n12057), .ZN(n7221) );
  NAND2_X1 U7746 ( .A1(n11397), .A2(n6728), .ZN(n11400) );
  OR2_X1 U7747 ( .A1(n7571), .A2(n11401), .ZN(n7570) );
  INV_X1 U7748 ( .A(n11399), .ZN(n7571) );
  NOR2_X1 U7749 ( .A1(n11402), .A2(n11399), .ZN(n7572) );
  NAND2_X1 U7750 ( .A1(n6785), .A2(n6786), .ZN(n12080) );
  NOR2_X1 U7751 ( .A1(n12088), .A2(n12087), .ZN(n7690) );
  INV_X1 U7752 ( .A(n12079), .ZN(n6784) );
  OAI21_X1 U7753 ( .B1(n11412), .B2(n7566), .A(n6921), .ZN(n11416) );
  OAI21_X1 U7754 ( .B1(n6734), .B2(n6733), .A(n11414), .ZN(n11417) );
  AND2_X1 U7755 ( .A1(n7564), .A2(n7563), .ZN(n6921) );
  NAND2_X1 U7756 ( .A1(n12100), .A2(n6657), .ZN(n7227) );
  AND2_X1 U7757 ( .A1(n11434), .A2(n11429), .ZN(n7551) );
  NAND2_X1 U7758 ( .A1(n7549), .A2(n7547), .ZN(n7546) );
  AND2_X1 U7759 ( .A1(n11425), .A2(n7550), .ZN(n7549) );
  INV_X1 U7760 ( .A(n11424), .ZN(n7550) );
  NOR2_X1 U7761 ( .A1(n6741), .A2(n6740), .ZN(n6739) );
  INV_X1 U7762 ( .A(n11418), .ZN(n6740) );
  NOR2_X1 U7763 ( .A1(n6741), .A2(n11421), .ZN(n6738) );
  NOR2_X1 U7764 ( .A1(n12137), .A2(n12148), .ZN(n12145) );
  NAND2_X1 U7765 ( .A1(n6780), .A2(n6777), .ZN(n12122) );
  NAND2_X1 U7766 ( .A1(n6779), .A2(n6778), .ZN(n6777) );
  NAND2_X1 U7767 ( .A1(n6782), .A2(n6781), .ZN(n6780) );
  INV_X1 U7768 ( .A(n12117), .ZN(n6778) );
  NAND2_X1 U7769 ( .A1(n11451), .A2(n6974), .ZN(n6973) );
  INV_X1 U7770 ( .A(n11452), .ZN(n6974) );
  INV_X1 U7771 ( .A(n12165), .ZN(n7653) );
  INV_X1 U7772 ( .A(n12175), .ZN(n6891) );
  NAND2_X1 U7773 ( .A1(n11503), .A2(n11502), .ZN(n11501) );
  OR2_X1 U7774 ( .A1(n11503), .A2(n11502), .ZN(n11504) );
  NAND2_X1 U7775 ( .A1(n7580), .A2(n11518), .ZN(n7579) );
  INV_X1 U7776 ( .A(n12180), .ZN(n6934) );
  OR2_X1 U7777 ( .A1(n10923), .A2(n10922), .ZN(n10929) );
  NAND2_X1 U7778 ( .A1(n12970), .A2(n10927), .ZN(n10930) );
  OR2_X1 U7779 ( .A1(n7576), .A2(n11589), .ZN(n7574) );
  NAND2_X1 U7780 ( .A1(n7576), .A2(n11589), .ZN(n7575) );
  INV_X1 U7781 ( .A(n11604), .ZN(n6969) );
  NAND2_X1 U7782 ( .A1(n7169), .A2(n7806), .ZN(n7168) );
  INV_X1 U7783 ( .A(n7805), .ZN(n7169) );
  AOI22_X1 U7784 ( .A1(n7787), .A2(n7786), .B1(n7785), .B2(n8110), .ZN(n7792)
         );
  INV_X1 U7785 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U7786 ( .A1(n7682), .A2(n7683), .ZN(n7681) );
  INV_X1 U7787 ( .A(n11700), .ZN(n7389) );
  AND2_X1 U7788 ( .A1(n8106), .A2(n7792), .ZN(n7789) );
  OAI21_X1 U7789 ( .B1(n6535), .B2(n8456), .A(n6926), .ZN(n7739) );
  OR2_X1 U7790 ( .A1(n9161), .A2(n8553), .ZN(n6926) );
  INV_X1 U7791 ( .A(n9673), .ZN(n7525) );
  OR2_X1 U7792 ( .A1(n12628), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U7793 ( .A1(n9144), .A2(n9100), .ZN(n9295) );
  NAND2_X1 U7794 ( .A1(n9440), .A2(n9441), .ZN(n9611) );
  NAND2_X1 U7795 ( .A1(n10963), .A2(n10964), .ZN(n12692) );
  INV_X1 U7796 ( .A(n6870), .ZN(n6871) );
  NAND2_X1 U7797 ( .A1(n10541), .A2(n6613), .ZN(n10907) );
  AND2_X1 U7798 ( .A1(n11867), .A2(n11868), .ZN(n11988) );
  INV_X1 U7799 ( .A(n11841), .ZN(n6705) );
  NAND2_X1 U7800 ( .A1(n15042), .A2(n11994), .ZN(n9889) );
  INV_X1 U7801 ( .A(n12010), .ZN(n7208) );
  AND2_X1 U7802 ( .A1(n12667), .A2(n12855), .ZN(n11943) );
  NOR2_X1 U7803 ( .A1(n12850), .A2(n6881), .ZN(n6880) );
  INV_X1 U7804 ( .A(n11288), .ZN(n6881) );
  INV_X1 U7805 ( .A(n12915), .ZN(n6873) );
  INV_X1 U7806 ( .A(n6847), .ZN(n6846) );
  AND2_X1 U7807 ( .A1(n6845), .A2(n12949), .ZN(n6844) );
  NAND2_X1 U7808 ( .A1(n6847), .A2(n6850), .ZN(n6845) );
  NAND2_X1 U7809 ( .A1(n11901), .A2(n11899), .ZN(n6701) );
  OR2_X1 U7810 ( .A1(n14568), .A2(n10976), .ZN(n11893) );
  AND2_X1 U7811 ( .A1(n14568), .A2(n10976), .ZN(n11895) );
  NAND2_X1 U7812 ( .A1(n15045), .A2(n15044), .ZN(n15043) );
  OR2_X1 U7813 ( .A1(n11198), .A2(n9248), .ZN(n9249) );
  NOR2_X1 U7814 ( .A1(n9056), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U7815 ( .A1(n10585), .A2(n10584), .ZN(n10586) );
  INV_X1 U7816 ( .A(n7076), .ZN(n7075) );
  AND2_X1 U7817 ( .A1(n9834), .A2(n7363), .ZN(n7362) );
  INV_X1 U7818 ( .A(n9837), .ZN(n7363) );
  NAND2_X1 U7819 ( .A1(n9689), .A2(n9688), .ZN(n9833) );
  INV_X1 U7820 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8408) );
  AND2_X1 U7821 ( .A1(n8529), .A2(n8528), .ZN(n8584) );
  INV_X1 U7822 ( .A(n8503), .ZN(n7086) );
  NOR2_X2 U7823 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8440) );
  AND2_X1 U7824 ( .A1(n7701), .A2(n6615), .ZN(n7589) );
  INV_X1 U7825 ( .A(n12257), .ZN(n7236) );
  AND2_X1 U7826 ( .A1(n7231), .A2(n6592), .ZN(n7237) );
  NOR2_X1 U7827 ( .A1(n7238), .A2(n12257), .ZN(n7235) );
  AND2_X1 U7828 ( .A1(n12227), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U7829 ( .A1(n12375), .A2(n12373), .ZN(n7645) );
  INV_X1 U7830 ( .A(n12373), .ZN(n7722) );
  NAND2_X1 U7831 ( .A1(n13424), .A2(n8356), .ZN(n7440) );
  INV_X1 U7832 ( .A(n13525), .ZN(n7454) );
  NAND2_X1 U7833 ( .A1(n13537), .A2(n13536), .ZN(n13535) );
  INV_X1 U7834 ( .A(n10804), .ZN(n7450) );
  INV_X1 U7835 ( .A(n7976), .ZN(n7269) );
  INV_X1 U7836 ( .A(n7896), .ZN(n7273) );
  NAND2_X1 U7837 ( .A1(n7442), .A2(n7852), .ZN(n8313) );
  OAI21_X1 U7838 ( .B1(n7442), .B2(n7852), .A(n8313), .ZN(n8312) );
  INV_X1 U7839 ( .A(n7275), .ZN(n7274) );
  AND2_X1 U7840 ( .A1(n10418), .A2(n9915), .ZN(n9323) );
  OR2_X1 U7841 ( .A1(n7902), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7932) );
  NOR2_X1 U7842 ( .A1(n11639), .A2(n7561), .ZN(n7558) );
  INV_X1 U7843 ( .A(n11583), .ZN(n11626) );
  INV_X1 U7844 ( .A(n6581), .ZN(n7413) );
  NOR2_X1 U7845 ( .A1(n7329), .A2(n14485), .ZN(n7326) );
  INV_X1 U7846 ( .A(n10597), .ZN(n7328) );
  INV_X1 U7847 ( .A(n11656), .ZN(n7304) );
  INV_X1 U7848 ( .A(n10237), .ZN(n7305) );
  INV_X1 U7849 ( .A(n7321), .ZN(n7320) );
  AND2_X1 U7850 ( .A1(n11650), .A2(n7318), .ZN(n7317) );
  NAND2_X1 U7851 ( .A1(n7319), .A2(n7321), .ZN(n7318) );
  INV_X1 U7852 ( .A(n7322), .ZN(n7319) );
  NOR2_X1 U7853 ( .A1(n9389), .A2(n6564), .ZN(n7422) );
  INV_X1 U7854 ( .A(n9525), .ZN(n7425) );
  XNOR2_X1 U7855 ( .A(n7537), .B(n13955), .ZN(n11644) );
  INV_X1 U7856 ( .A(n14374), .ZN(n11305) );
  INV_X1 U7857 ( .A(n8206), .ZN(n7151) );
  NAND2_X1 U7858 ( .A1(n7802), .A2(SI_22_), .ZN(n7805) );
  AOI21_X1 U7859 ( .B1(n7593), .B2(n7595), .A(n7591), .ZN(n7590) );
  INV_X1 U7860 ( .A(n7781), .ZN(n7591) );
  NOR2_X1 U7861 ( .A1(n8045), .A2(SI_14_), .ZN(n6715) );
  NAND2_X1 U7862 ( .A1(n8045), .A2(SI_14_), .ZN(n6714) );
  INV_X1 U7863 ( .A(n7778), .ZN(n8045) );
  NAND2_X1 U7864 ( .A1(n8018), .A2(n7774), .ZN(n8031) );
  NOR2_X1 U7865 ( .A1(n7766), .A2(n7159), .ZN(n7158) );
  INV_X1 U7866 ( .A(n7996), .ZN(n7159) );
  NAND3_X1 U7867 ( .A1(n7376), .A2(n7490), .A3(n7375), .ZN(n8429) );
  INV_X1 U7868 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7375) );
  INV_X1 U7869 ( .A(n6930), .ZN(n14384) );
  INV_X1 U7870 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14385) );
  XNOR2_X1 U7871 ( .A(n14384), .B(n14385), .ZN(n14442) );
  OAI22_X1 U7872 ( .A1(n14446), .A2(n14389), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14388), .ZN(n14390) );
  INV_X1 U7873 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14388) );
  AOI21_X1 U7874 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14395), .A(n14394), .ZN(
        n14454) );
  NOR2_X1 U7875 ( .A1(n14427), .A2(n14426), .ZN(n14394) );
  INV_X1 U7876 ( .A(n11789), .ZN(n11770) );
  INV_X1 U7877 ( .A(n11780), .ZN(n7045) );
  INV_X1 U7878 ( .A(n11782), .ZN(n7521) );
  AOI21_X1 U7879 ( .B1(n12571), .B2(n7519), .A(n7522), .ZN(n7518) );
  AND2_X1 U7880 ( .A1(n11787), .A2(n11788), .ZN(n7522) );
  AND2_X1 U7881 ( .A1(n12610), .A2(n7040), .ZN(n7039) );
  NAND2_X1 U7882 ( .A1(n11753), .A2(n11752), .ZN(n7040) );
  INV_X1 U7883 ( .A(n7018), .ZN(n7527) );
  INV_X1 U7884 ( .A(n7039), .ZN(n7037) );
  OR2_X1 U7885 ( .A1(n9666), .A2(n15047), .ZN(n7526) );
  OR2_X1 U7886 ( .A1(n11882), .A2(n10708), .ZN(n7535) );
  INV_X1 U7887 ( .A(n7534), .ZN(n7532) );
  NAND2_X1 U7888 ( .A1(n9066), .A2(n7053), .ZN(n9112) );
  OR2_X1 U7889 ( .A1(n9069), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U7890 ( .A1(n7512), .A2(n6596), .ZN(n7060) );
  OR2_X1 U7891 ( .A1(n9090), .A2(n15260), .ZN(n7512) );
  NAND2_X1 U7892 ( .A1(n7060), .A2(n7059), .ZN(n9140) );
  INV_X1 U7893 ( .A(n9142), .ZN(n7059) );
  XNOR2_X1 U7894 ( .A(n9295), .B(n9987), .ZN(n9101) );
  NAND2_X1 U7895 ( .A1(n9101), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9297) );
  AND2_X1 U7896 ( .A1(n9140), .A2(n9092), .ZN(n9291) );
  XNOR2_X1 U7897 ( .A(n9291), .B(n9987), .ZN(n9292) );
  XNOR2_X1 U7898 ( .A(n9611), .B(n10263), .ZN(n9442) );
  NAND2_X1 U7899 ( .A1(n9442), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U7900 ( .A1(n7509), .A2(n6595), .ZN(n7065) );
  OR2_X1 U7901 ( .A1(n9607), .A2(n9608), .ZN(n7509) );
  NAND2_X1 U7902 ( .A1(n14989), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n14988) );
  AOI21_X1 U7903 ( .B1(n7065), .B2(n7064), .A(n7514), .ZN(n9956) );
  AND2_X1 U7904 ( .A1(n10271), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7514) );
  INV_X1 U7905 ( .A(n9954), .ZN(n7064) );
  INV_X1 U7906 ( .A(n10522), .ZN(n10540) );
  NOR2_X1 U7907 ( .A1(n10521), .A2(n7515), .ZN(n10648) );
  AND2_X1 U7908 ( .A1(n10522), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U7909 ( .A1(n10658), .A2(n10659), .ZN(n10963) );
  NOR2_X1 U7910 ( .A1(n10955), .A2(n7500), .ZN(n12687) );
  NOR2_X1 U7911 ( .A1(n10654), .A2(n7501), .ZN(n7500) );
  INV_X1 U7912 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n7501) );
  XNOR2_X1 U7913 ( .A(n12692), .B(n12707), .ZN(n10965) );
  NAND2_X1 U7914 ( .A1(n10965), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12694) );
  NAND2_X1 U7915 ( .A1(n12756), .A2(n12757), .ZN(n12784) );
  NAND2_X1 U7916 ( .A1(n7510), .A2(n12752), .ZN(n12766) );
  XNOR2_X1 U7917 ( .A(n12787), .B(n12786), .ZN(n14528) );
  AOI21_X1 U7918 ( .B1(n12849), .B2(n12850), .A(n11256), .ZN(n12834) );
  AND4_X1 U7919 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n12961)
         );
  AND4_X1 U7920 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n11033) );
  NAND2_X1 U7921 ( .A1(n10911), .A2(n11888), .ZN(n14567) );
  NOR2_X1 U7922 ( .A1(n10696), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n10717) );
  OR2_X1 U7923 ( .A1(n10544), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10696) );
  INV_X1 U7924 ( .A(n14997), .ZN(n6708) );
  OR2_X1 U7925 ( .A1(n10257), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U7926 ( .A1(n10275), .A2(n10255), .ZN(n10257) );
  AOI21_X1 U7927 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(n10450) );
  AND3_X1 U7928 ( .A1(n10266), .A2(n10265), .A3(n10264), .ZN(n10457) );
  AND4_X1 U7929 ( .A1(n9999), .A2(n9998), .A3(n9997), .A4(n9996), .ZN(n10281)
         );
  NAND2_X1 U7930 ( .A1(n9902), .A2(n11850), .ZN(n10128) );
  INV_X1 U7931 ( .A(n9690), .ZN(n9890) );
  NAND2_X1 U7932 ( .A1(n11963), .A2(n11962), .ZN(n12015) );
  NOR2_X1 U7933 ( .A1(n7208), .A2(n6863), .ZN(n6862) );
  NAND2_X1 U7934 ( .A1(n6539), .A2(n15068), .ZN(n6863) );
  NAND2_X1 U7935 ( .A1(n11276), .A2(n11275), .ZN(n11278) );
  NAND2_X1 U7936 ( .A1(n12828), .A2(n15065), .ZN(n6929) );
  XNOR2_X1 U7937 ( .A(n13053), .B(n12837), .ZN(n12826) );
  NAND2_X1 U7938 ( .A1(n6882), .A2(n11288), .ZN(n12851) );
  OR2_X1 U7939 ( .A1(n6866), .A2(n11815), .ZN(n6865) );
  NAND2_X1 U7940 ( .A1(n6873), .A2(n6566), .ZN(n6872) );
  AOI21_X1 U7941 ( .B1(n12949), .B2(n11822), .A(n7263), .ZN(n7262) );
  NAND2_X1 U7942 ( .A1(n7261), .A2(n7259), .ZN(n12922) );
  NOR2_X1 U7943 ( .A1(n12919), .A2(n7260), .ZN(n7259) );
  INV_X1 U7944 ( .A(n7262), .ZN(n7260) );
  OAI21_X1 U7945 ( .B1(n11281), .B2(n6846), .A(n6844), .ZN(n12948) );
  NAND2_X1 U7946 ( .A1(n6848), .A2(n6545), .ZN(n6847) );
  NAND2_X1 U7947 ( .A1(n11163), .A2(n11915), .ZN(n12944) );
  NAND2_X1 U7948 ( .A1(n6702), .A2(n7245), .ZN(n12957) );
  AOI21_X1 U7949 ( .B1(n6574), .B2(n7249), .A(n7246), .ZN(n7245) );
  OAI21_X1 U7950 ( .B1(n11018), .B2(n11902), .A(n6552), .ZN(n6702) );
  INV_X1 U7951 ( .A(n11906), .ZN(n7249) );
  NAND2_X1 U7952 ( .A1(n11910), .A2(n11911), .ZN(n12002) );
  NAND2_X1 U7953 ( .A1(n6700), .A2(n11899), .ZN(n11038) );
  NAND2_X1 U7954 ( .A1(n11018), .A2(n11900), .ZN(n6700) );
  NAND2_X1 U7955 ( .A1(n7204), .A2(n12975), .ZN(n10933) );
  NAND2_X1 U7956 ( .A1(n12974), .A2(n7200), .ZN(n7204) );
  NAND2_X1 U7957 ( .A1(n9883), .A2(n11955), .ZN(n15046) );
  INV_X1 U7958 ( .A(n15062), .ZN(n15048) );
  AND4_X1 U7959 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(n10240)
         );
  NAND2_X1 U7960 ( .A1(n11828), .A2(n10134), .ZN(n15054) );
  NAND2_X1 U7961 ( .A1(n8565), .A2(n10800), .ZN(n9176) );
  AND2_X1 U7962 ( .A1(n8412), .A2(n7256), .ZN(n6710) );
  AND2_X1 U7963 ( .A1(n7257), .A2(n15338), .ZN(n7256) );
  NAND2_X1 U7964 ( .A1(n7357), .A2(n11145), .ZN(n11269) );
  NAND2_X1 U7965 ( .A1(n11144), .A2(n11143), .ZN(n7357) );
  NAND2_X1 U7966 ( .A1(n10765), .A2(n7092), .ZN(n10797) );
  NAND2_X1 U7967 ( .A1(n10587), .A2(n11801), .ZN(n7092) );
  OR2_X1 U7968 ( .A1(n10586), .A2(n10953), .ZN(n10765) );
  INV_X1 U7969 ( .A(n10368), .ZN(n7364) );
  NAND2_X1 U7970 ( .A1(n7362), .A2(n9835), .ZN(n10187) );
  INV_X1 U7971 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9178) );
  AND2_X1 U7972 ( .A1(n7047), .A2(n9053), .ZN(n7046) );
  NAND2_X1 U7973 ( .A1(n9346), .A2(n9345), .ZN(n9689) );
  NAND2_X1 U7974 ( .A1(n9037), .A2(n7081), .ZN(n7080) );
  NOR2_X1 U7975 ( .A1(n9210), .A2(n7082), .ZN(n7081) );
  INV_X1 U7976 ( .A(n9036), .ZN(n7082) );
  OAI21_X1 U7977 ( .B1(n8864), .B2(n8863), .A(n8865), .ZN(n9035) );
  NAND2_X1 U7978 ( .A1(n7094), .A2(n8620), .ZN(n8690) );
  NAND2_X1 U7979 ( .A1(n8618), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7094) );
  XNOR2_X1 U7980 ( .A(n8619), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U7981 ( .A1(n7345), .A2(n8533), .ZN(n8587) );
  NOR2_X1 U7982 ( .A1(n8515), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8536) );
  AND2_X1 U7983 ( .A1(n8471), .A2(n8470), .ZN(n8518) );
  OAI21_X1 U7984 ( .B1(n8464), .B2(n7085), .A(n7083), .ZN(n8521) );
  INV_X1 U7985 ( .A(n7084), .ZN(n7083) );
  OAI21_X1 U7986 ( .B1(n6569), .B2(n7085), .A(n7346), .ZN(n7084) );
  NAND2_X1 U7987 ( .A1(n8469), .A2(n8466), .ZN(n7085) );
  OR2_X1 U7988 ( .A1(n6562), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8515) );
  AND2_X1 U7989 ( .A1(n8469), .A2(n8468), .ZN(n8509) );
  INV_X1 U7990 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U7991 ( .A1(n8506), .A2(n8466), .ZN(n8510) );
  NAND2_X1 U7992 ( .A1(n8510), .A2(n8509), .ZN(n8512) );
  NAND2_X1 U7993 ( .A1(n8464), .A2(n6569), .ZN(n8506) );
  NAND2_X1 U7994 ( .A1(n7068), .A2(n7066), .ZN(n8547) );
  AOI21_X1 U7995 ( .B1(n7070), .B2(n7072), .A(n7067), .ZN(n7066) );
  INV_X1 U7996 ( .A(n8461), .ZN(n7067) );
  AND2_X1 U7997 ( .A1(n8461), .A2(n8460), .ZN(n8490) );
  AND2_X1 U7998 ( .A1(n8458), .A2(n8457), .ZN(n8482) );
  NAND2_X1 U7999 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8439) );
  INV_X1 U8000 ( .A(n12346), .ZN(n6698) );
  XNOR2_X1 U8001 ( .A(n7852), .B(n6529), .ZN(n9570) );
  INV_X1 U8002 ( .A(n7120), .ZN(n7119) );
  OAI21_X1 U8003 ( .B1(n12359), .B2(n7121), .A(n12399), .ZN(n7120) );
  INV_X1 U8004 ( .A(n12402), .ZN(n7118) );
  AND2_X1 U8005 ( .A1(n12357), .A2(n12355), .ZN(n13162) );
  INV_X1 U8006 ( .A(n9576), .ZN(n9566) );
  NAND2_X1 U8007 ( .A1(n13557), .A2(n12044), .ZN(n9574) );
  INV_X1 U8008 ( .A(n13207), .ZN(n7126) );
  INV_X1 U8009 ( .A(n12317), .ZN(n7128) );
  INV_X1 U8010 ( .A(n13247), .ZN(n13214) );
  NAND2_X1 U8011 ( .A1(n6989), .A2(n6558), .ZN(n7477) );
  XNOR2_X1 U8012 ( .A(n9371), .B(n7108), .ZN(n9317) );
  INV_X1 U8013 ( .A(n9376), .ZN(n7108) );
  OR2_X1 U8014 ( .A1(n8096), .A2(n8095), .ZN(n8117) );
  NOR2_X1 U8015 ( .A1(n9322), .A2(n14912), .ZN(n9336) );
  OR2_X1 U8016 ( .A1(n6525), .A2(n10166), .ZN(n7840) );
  AND2_X1 U8017 ( .A1(n14825), .A2(n14826), .ZN(n14823) );
  NOR2_X1 U8018 ( .A1(n14823), .A2(n7008), .ZN(n8957) );
  AND2_X1 U8019 ( .A1(n14829), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7008) );
  OR2_X1 U8020 ( .A1(n8957), .A2(n8956), .ZN(n7007) );
  OR2_X1 U8021 ( .A1(n8903), .A2(n8902), .ZN(n6995) );
  XNOR2_X1 U8022 ( .A(n11068), .B(n11081), .ZN(n13329) );
  NOR2_X1 U8023 ( .A1(n13316), .A2(n7009), .ZN(n11068) );
  AND2_X1 U8024 ( .A1(n11078), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7009) );
  NOR2_X1 U8025 ( .A1(n13329), .A2(n11069), .ZN(n13330) );
  AND3_X1 U8026 ( .A1(n7676), .A2(n7678), .A3(n7677), .ZN(n8087) );
  INV_X1 U8027 ( .A(n13616), .ZN(n7373) );
  NOR2_X1 U8028 ( .A1(n7439), .A2(n13432), .ZN(n7438) );
  NAND2_X1 U8029 ( .A1(n13436), .A2(n13714), .ZN(n13420) );
  NOR2_X1 U8030 ( .A1(n13464), .A2(n7295), .ZN(n7294) );
  INV_X1 U8031 ( .A(n12292), .ZN(n7295) );
  OR2_X1 U8032 ( .A1(n13477), .A2(n8193), .ZN(n7296) );
  INV_X1 U8033 ( .A(n7283), .ZN(n7282) );
  OAI21_X1 U8034 ( .B1(n8123), .B2(n6559), .A(n8140), .ZN(n7283) );
  NAND2_X1 U8035 ( .A1(n13535), .A2(n6565), .ZN(n13522) );
  INV_X1 U8036 ( .A(n7444), .ZN(n7443) );
  OAI21_X1 U8037 ( .B1(n7445), .B2(n8336), .A(n8339), .ZN(n7444) );
  INV_X1 U8038 ( .A(n12287), .ZN(n13567) );
  NAND2_X1 U8039 ( .A1(n8063), .A2(n8062), .ZN(n7287) );
  NAND2_X1 U8040 ( .A1(n7447), .A2(n11094), .ZN(n11099) );
  INV_X1 U8041 ( .A(n11098), .ZN(n7447) );
  AND2_X1 U8042 ( .A1(n12275), .A2(n8323), .ZN(n7457) );
  NAND2_X1 U8043 ( .A1(n6942), .A2(n7277), .ZN(n10401) );
  CLKBUF_X1 U8044 ( .A(n10299), .Z(n6942) );
  NAND2_X1 U8045 ( .A1(n10176), .A2(n10175), .ZN(n10174) );
  NAND2_X1 U8046 ( .A1(n8309), .A2(n12044), .ZN(n10068) );
  OR2_X1 U8047 ( .A1(n12053), .A2(n13269), .ZN(n6886) );
  NAND2_X1 U8048 ( .A1(n6889), .A2(n6888), .ZN(n6887) );
  INV_X1 U8049 ( .A(n9450), .ZN(n6888) );
  AND2_X1 U8050 ( .A1(n12042), .A2(n9467), .ZN(n9450) );
  NAND2_X1 U8051 ( .A1(n8160), .A2(n8159), .ZN(n13512) );
  OR2_X1 U8052 ( .A1(n11497), .A2(n8171), .ZN(n8160) );
  INV_X1 U8053 ( .A(n13557), .ZN(n14896) );
  INV_X1 U8054 ( .A(n13699), .ZN(n14927) );
  INV_X1 U8055 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7715) );
  AND2_X1 U8056 ( .A1(n7678), .A2(n7817), .ZN(n7243) );
  INV_X1 U8057 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8264) );
  AOI21_X1 U8058 ( .B1(n6643), .B2(P2_IR_REG_31__SCAN_IN), .A(n7485), .ZN(
        n7484) );
  INV_X1 U8059 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7487) );
  AND2_X2 U8060 ( .A1(n8087), .A2(n8086), .ZN(n8091) );
  AND2_X1 U8061 ( .A1(n7014), .A2(n7013), .ZN(n7844) );
  AND2_X1 U8062 ( .A1(n7614), .A2(n7615), .ZN(n7613) );
  INV_X1 U8063 ( .A(n10503), .ZN(n7614) );
  NAND2_X1 U8064 ( .A1(n13871), .A2(n13870), .ZN(n7643) );
  AND2_X1 U8065 ( .A1(n12532), .A2(n12531), .ZN(n13832) );
  AND2_X1 U8066 ( .A1(n12447), .A2(n7637), .ZN(n7636) );
  INV_X1 U8067 ( .A(n13842), .ZN(n7637) );
  AND2_X1 U8068 ( .A1(n13834), .A2(n12519), .ZN(n13862) );
  NAND2_X1 U8069 ( .A1(n6547), .A2(n6614), .ZN(n7192) );
  NAND2_X1 U8070 ( .A1(n7195), .A2(n12464), .ZN(n7194) );
  NAND2_X1 U8071 ( .A1(n13840), .A2(n13849), .ZN(n12463) );
  AOI21_X1 U8072 ( .B1(n7634), .B2(n7184), .A(n6638), .ZN(n7183) );
  INV_X1 U8073 ( .A(n14611), .ZN(n7184) );
  AOI22_X1 U8074 ( .A1(n7196), .A2(n7537), .B1(n9019), .B2(n13955), .ZN(n8880)
         );
  INV_X1 U8075 ( .A(n11564), .ZN(n11607) );
  NAND2_X1 U8076 ( .A1(n8723), .A2(n8724), .ZN(n8722) );
  NAND2_X1 U8077 ( .A1(n10487), .A2(n6833), .ZN(n10489) );
  OR2_X1 U8078 ( .A1(n10733), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6833) );
  INV_X1 U8079 ( .A(n7415), .ZN(n7414) );
  NOR2_X1 U8080 ( .A1(n14125), .A2(n7334), .ZN(n7333) );
  INV_X1 U8081 ( .A(n11713), .ZN(n7334) );
  NAND2_X1 U8082 ( .A1(n14174), .A2(n11710), .ZN(n14149) );
  INV_X1 U8083 ( .A(n11693), .ZN(n7385) );
  AND4_X1 U8084 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n12410) );
  OR2_X1 U8085 ( .A1(n10214), .A2(n10235), .ZN(n7408) );
  NAND2_X1 U8086 ( .A1(n7324), .A2(n7323), .ZN(n7322) );
  NAND2_X1 U8087 ( .A1(n11385), .A2(n11386), .ZN(n7321) );
  AND2_X1 U8088 ( .A1(n9516), .A2(n11385), .ZN(n6810) );
  CLKBUF_X1 U8089 ( .A(n9740), .Z(n6932) );
  NAND2_X1 U8090 ( .A1(n9648), .A2(n9231), .ZN(n9233) );
  INV_X1 U8091 ( .A(n11644), .ZN(n9655) );
  INV_X1 U8092 ( .A(n14221), .ZN(n14631) );
  INV_X1 U8093 ( .A(n11308), .ZN(n11633) );
  NAND2_X1 U8094 ( .A1(n8825), .A2(n8571), .ZN(n8835) );
  INV_X1 U8095 ( .A(n14039), .ZN(n14270) );
  NAND2_X1 U8096 ( .A1(n11615), .A2(n11614), .ZN(n14273) );
  OR2_X1 U8097 ( .A1(n11338), .A2(n11496), .ZN(n11340) );
  NAND2_X1 U8098 ( .A1(n11457), .A2(n11456), .ZN(n14343) );
  OR2_X1 U8099 ( .A1(n11516), .A2(n6931), .ZN(n8878) );
  AND2_X1 U8100 ( .A1(n7313), .A2(n8810), .ZN(n7311) );
  NAND2_X1 U8101 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7312) );
  INV_X1 U8102 ( .A(n7312), .ZN(n7310) );
  AND2_X1 U8103 ( .A1(n8251), .A2(n8237), .ZN(n8249) );
  AOI21_X1 U8104 ( .B1(n7601), .B2(n7812), .A(n6689), .ZN(n7600) );
  NAND2_X1 U8105 ( .A1(n7149), .A2(n6687), .ZN(n7813) );
  NAND2_X1 U8106 ( .A1(n8170), .A2(n7805), .ZN(n7165) );
  OR2_X1 U8107 ( .A1(n11514), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U8108 ( .A1(n7805), .A2(n7803), .ZN(n11514) );
  OR2_X1 U8109 ( .A1(n7802), .A2(SI_22_), .ZN(n7803) );
  NAND2_X1 U8110 ( .A1(n8156), .A2(n8155), .ZN(n8158) );
  INV_X1 U8111 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7577) );
  AND2_X2 U8112 ( .A1(n8611), .A2(n7199), .ZN(n8390) );
  AND2_X1 U8113 ( .A1(n8383), .A2(n8391), .ZN(n7578) );
  NOR2_X1 U8114 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8383) );
  NAND2_X1 U8115 ( .A1(n7797), .A2(n7606), .ZN(n7605) );
  INV_X1 U8116 ( .A(n8141), .ZN(n7606) );
  INV_X1 U8117 ( .A(n7798), .ZN(n7604) );
  INV_X1 U8118 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7490) );
  CLKBUF_X1 U8119 ( .A(n8429), .Z(n6916) );
  INV_X1 U8120 ( .A(n6753), .ZN(n14432) );
  NAND2_X1 U8121 ( .A1(n6979), .A2(n14441), .ZN(n14444) );
  NAND2_X1 U8122 ( .A1(n7470), .A2(n14448), .ZN(n14450) );
  INV_X1 U8123 ( .A(n6751), .ZN(n14456) );
  OAI21_X1 U8124 ( .B1(n14482), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6586), .ZN(
        n6751) );
  OAI21_X1 U8125 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14422) );
  AND2_X1 U8126 ( .A1(n7106), .A2(n7107), .ZN(n14467) );
  AOI22_X1 U8127 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14407), .B1(n14465), 
        .B2(n14406), .ZN(n14419) );
  NAND2_X1 U8128 ( .A1(n14704), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7101) );
  OAI21_X1 U8129 ( .B1(n14512), .B2(n14513), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n7464) );
  INV_X1 U8130 ( .A(n13053), .ZN(n12579) );
  NAND2_X1 U8131 ( .A1(n11224), .A2(n11223), .ZN(n13012) );
  NOR2_X1 U8132 ( .A1(n10555), .A2(n7029), .ZN(n10689) );
  OR2_X1 U8133 ( .A1(n10554), .A2(n10557), .ZN(n7029) );
  AND4_X1 U8134 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n12936) );
  AND4_X1 U8135 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10445) );
  MUX2_X1 U8136 ( .A(n15067), .B(n11832), .S(n11789), .Z(n9260) );
  NAND3_X1 U8137 ( .A1(n7023), .A2(n7017), .A3(n7016), .ZN(n10292) );
  NAND2_X1 U8138 ( .A1(n9543), .A2(n7019), .ZN(n7023) );
  NOR2_X1 U8139 ( .A1(n10293), .A2(n10294), .ZN(n10555) );
  NAND2_X1 U8140 ( .A1(n11189), .A2(n11188), .ZN(n13022) );
  XNOR2_X1 U8141 ( .A(n10709), .B(n10708), .ZN(n10710) );
  INV_X1 U8142 ( .A(n12872), .ZN(n12899) );
  INV_X1 U8143 ( .A(n12656), .ZN(n12951) );
  INV_X1 U8144 ( .A(n12961), .ZN(n12621) );
  INV_X1 U8145 ( .A(n15019), .ZN(n10919) );
  XNOR2_X1 U8146 ( .A(n9956), .B(n10254), .ZN(n14974) );
  NOR2_X1 U8147 ( .A1(n14974), .A2(n15030), .ZN(n14973) );
  XNOR2_X1 U8148 ( .A(n10648), .B(n10692), .ZN(n10523) );
  XNOR2_X1 U8149 ( .A(n12687), .B(n12707), .ZN(n10956) );
  OR2_X1 U8150 ( .A1(n12722), .A2(n12723), .ZN(n7511) );
  XNOR2_X1 U8151 ( .A(n12748), .B(n12755), .ZN(n12722) );
  NAND2_X1 U8152 ( .A1(n12796), .A2(n12795), .ZN(n6766) );
  XNOR2_X1 U8153 ( .A(n6768), .B(n12790), .ZN(n6767) );
  NAND2_X1 U8154 ( .A1(n14544), .A2(n6938), .ZN(n6768) );
  OR2_X1 U8155 ( .A1(n14542), .A2(n13028), .ZN(n6938) );
  INV_X1 U8156 ( .A(n12794), .ZN(n6765) );
  NAND2_X1 U8157 ( .A1(n11153), .A2(n11152), .ZN(n12381) );
  NAND2_X1 U8158 ( .A1(n6947), .A2(n6945), .ZN(n12992) );
  NOR2_X1 U8159 ( .A1(n6946), .A2(n6675), .ZN(n6945) );
  NAND2_X1 U8160 ( .A1(n11162), .A2(n11161), .ZN(n13033) );
  AND2_X1 U8161 ( .A1(n9690), .A2(n12771), .ZN(n15056) );
  OR2_X1 U8162 ( .A1(n11198), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U8163 ( .A1(n11973), .A2(n11972), .ZN(n12986) );
  OR2_X1 U8164 ( .A1(n15142), .A2(n11299), .ZN(n7211) );
  AOI21_X1 U8165 ( .B1(n12807), .B2(n6862), .A(n6858), .ZN(n12380) );
  OAI21_X1 U8166 ( .B1(n12807), .B2(n6861), .A(n6859), .ZN(n6858) );
  OR2_X1 U8167 ( .A1(n12383), .A2(n13107), .ZN(n6991) );
  INV_X1 U8168 ( .A(n6851), .ZN(n6857) );
  AOI21_X1 U8169 ( .B1(n12807), .B2(n6854), .A(n6852), .ZN(n6851) );
  NOR2_X1 U8170 ( .A1(n6855), .A2(n15125), .ZN(n6854) );
  OAI21_X1 U8171 ( .B1(n6855), .B2(n6853), .A(n6557), .ZN(n6852) );
  INV_X1 U8172 ( .A(n11278), .ZN(n13050) );
  OR2_X1 U8173 ( .A1(n15127), .A2(n13048), .ZN(n6952) );
  NAND2_X1 U8174 ( .A1(n11213), .A2(n11212), .ZN(n13073) );
  NAND2_X1 U8175 ( .A1(n11166), .A2(n11165), .ZN(n13096) );
  OAI22_X1 U8176 ( .A1(n9176), .A2(P3_D_REG_0__SCAN_IN), .B1(n10800), .B2(
        n10581), .ZN(n11730) );
  NAND2_X1 U8177 ( .A1(n9050), .A2(n7529), .ZN(n7528) );
  INV_X1 U8178 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U8179 ( .A1(n12395), .A2(n6567), .ZN(n13125) );
  OAI211_X1 U8180 ( .C1(n6560), .C2(n10563), .A(n6699), .B(n11135), .ZN(n11141) );
  NAND2_X1 U8181 ( .A1(n6637), .A2(n11813), .ZN(n6699) );
  INV_X1 U8182 ( .A(n10563), .ZN(n7475) );
  NAND2_X1 U8183 ( .A1(n10737), .A2(n12230), .ZN(n8054) );
  INV_X1 U8184 ( .A(n10418), .ZN(n12305) );
  OR2_X1 U8185 ( .A1(n8061), .A2(n8060), .ZN(n13254) );
  OR2_X1 U8186 ( .A1(n8999), .A2(n8998), .ZN(n6997) );
  NAND2_X1 U8187 ( .A1(n13384), .A2(n13383), .ZN(n7003) );
  OAI22_X1 U8188 ( .A1(n13381), .A2(n14858), .B1(n13382), .B2(n14851), .ZN(
        n6999) );
  OAI21_X1 U8189 ( .B1(n14873), .B2(n15392), .A(n13385), .ZN(n7001) );
  INV_X1 U8190 ( .A(n8369), .ZN(n7144) );
  OR2_X1 U8191 ( .A1(n13401), .A2(n13406), .ZN(n7132) );
  OR2_X1 U8192 ( .A1(n11482), .A2(n8171), .ZN(n8146) );
  AND2_X2 U8193 ( .A1(n10078), .A2(n9462), .ZN(n14972) );
  AND2_X1 U8194 ( .A1(n10685), .A2(n8283), .ZN(n14916) );
  NAND2_X1 U8195 ( .A1(n7586), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U8196 ( .A1(n14284), .A2(n14616), .ZN(n6901) );
  OAI21_X1 U8197 ( .B1(n10842), .B2(n10841), .A(n10840), .ZN(n12417) );
  NAND2_X1 U8198 ( .A1(n13911), .A2(n13912), .ZN(n13910) );
  INV_X1 U8199 ( .A(n9018), .ZN(n6818) );
  INV_X1 U8200 ( .A(n13932), .ZN(n14612) );
  AND2_X1 U8201 ( .A1(n8889), .A2(n8926), .ZN(n14221) );
  OR2_X1 U8202 ( .A1(n11630), .A2(n8813), .ZN(n8816) );
  NOR2_X1 U8203 ( .A1(n8680), .A2(n8681), .ZN(n8695) );
  NAND2_X1 U8204 ( .A1(n8740), .A2(n8739), .ZN(n8754) );
  XNOR2_X1 U8205 ( .A(n10489), .B(n14725), .ZN(n14723) );
  NAND2_X1 U8206 ( .A1(n14723), .A2(n15326), .ZN(n14722) );
  INV_X1 U8207 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7728) );
  NOR2_X1 U8208 ( .A1(n14018), .A2(n6828), .ZN(n14019) );
  INV_X1 U8209 ( .A(n6830), .ZN(n6828) );
  INV_X1 U8210 ( .A(n14022), .ZN(n6836) );
  OAI21_X1 U8211 ( .B1(n14023), .B2(n14021), .A(n14020), .ZN(n6835) );
  XNOR2_X1 U8212 ( .A(n14035), .B(n14032), .ZN(n14028) );
  AND2_X1 U8213 ( .A1(n7338), .A2(n7337), .ZN(n14076) );
  NAND2_X1 U8214 ( .A1(n14071), .A2(n14070), .ZN(n14072) );
  INV_X1 U8215 ( .A(n11719), .ZN(n6897) );
  NAND2_X1 U8216 ( .A1(n11720), .A2(n14494), .ZN(n6898) );
  AND2_X1 U8217 ( .A1(n11484), .A2(n11483), .ZN(n14325) );
  NAND2_X1 U8218 ( .A1(n14269), .A2(n6914), .ZN(n14349) );
  INV_X1 U8219 ( .A(n6915), .ZN(n6914) );
  OAI21_X1 U8220 ( .B1(n14270), .B2(n14793), .A(n14268), .ZN(n6915) );
  INV_X1 U8221 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n15251) );
  OR2_X1 U8222 ( .A1(n8802), .A2(n8801), .ZN(n6730) );
  INV_X1 U8223 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14434) );
  XNOR2_X1 U8224 ( .A(n14435), .B(n6980), .ZN(n15449) );
  INV_X1 U8225 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6980) );
  AOI21_X1 U8226 ( .B1(n14839), .B2(n14438), .A(n14476), .ZN(n15447) );
  XNOR2_X1 U8227 ( .A(n14467), .B(n14466), .ZN(n14696) );
  AND3_X1 U8228 ( .A1(n7460), .A2(n7462), .A3(n7459), .ZN(n14701) );
  INV_X1 U8229 ( .A(n14471), .ZN(n7459) );
  NOR2_X1 U8230 ( .A1(n14701), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n14472) );
  NAND2_X1 U8231 ( .A1(n7460), .A2(n7462), .ZN(n14470) );
  NOR2_X1 U8232 ( .A1(n7463), .A2(n6578), .ZN(n14516) );
  AND2_X1 U8233 ( .A1(n7463), .A2(n6578), .ZN(n14515) );
  INV_X1 U8234 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U8235 ( .A1(n7538), .A2(n7536), .ZN(n7540) );
  NAND2_X1 U8236 ( .A1(n11348), .A2(n11363), .ZN(n7538) );
  NAND2_X1 U8237 ( .A1(n11362), .A2(n11373), .ZN(n7536) );
  INV_X1 U8238 ( .A(n12061), .ZN(n7220) );
  NOR2_X1 U8239 ( .A1(n12069), .A2(n12066), .ZN(n7669) );
  INV_X1 U8240 ( .A(n7564), .ZN(n6735) );
  AOI21_X1 U8241 ( .B1(n7572), .B2(n7570), .A(n7569), .ZN(n7568) );
  OAI21_X1 U8242 ( .B1(n11400), .B2(n7572), .A(n6627), .ZN(n11407) );
  INV_X1 U8243 ( .A(n12087), .ZN(n7689) );
  NAND2_X1 U8244 ( .A1(n7565), .A2(n11410), .ZN(n7564) );
  NOR2_X1 U8245 ( .A1(n11408), .A2(n6735), .ZN(n6733) );
  OAI21_X1 U8246 ( .B1(n11407), .B2(n6735), .A(n7562), .ZN(n6734) );
  AOI21_X1 U8247 ( .B1(n7566), .B2(n7564), .A(n7563), .ZN(n7562) );
  NAND2_X1 U8248 ( .A1(n11408), .A2(n11407), .ZN(n11412) );
  NOR2_X1 U8249 ( .A1(n7565), .A2(n11410), .ZN(n7566) );
  INV_X1 U8250 ( .A(n6657), .ZN(n7684) );
  NAND2_X1 U8251 ( .A1(n7686), .A2(n7687), .ZN(n6783) );
  NAND2_X1 U8252 ( .A1(n12112), .A2(n6597), .ZN(n7687) );
  OR2_X1 U8253 ( .A1(n12105), .A2(n6920), .ZN(n7686) );
  NAND2_X1 U8254 ( .A1(n14260), .A2(n11427), .ZN(n11437) );
  NAND2_X1 U8255 ( .A1(n11422), .A2(n6738), .ZN(n6736) );
  NAND2_X1 U8256 ( .A1(n11419), .A2(n6739), .ZN(n6737) );
  NAND2_X1 U8257 ( .A1(n6783), .A2(n12117), .ZN(n6782) );
  INV_X1 U8258 ( .A(n12116), .ZN(n6781) );
  INV_X1 U8259 ( .A(n6783), .ZN(n6779) );
  NAND2_X1 U8260 ( .A1(n7582), .A2(n11452), .ZN(n7581) );
  NAND2_X1 U8261 ( .A1(n12145), .A2(n6917), .ZN(n12159) );
  NOR2_X1 U8262 ( .A1(n12146), .A2(n12147), .ZN(n6917) );
  NAND2_X1 U8263 ( .A1(n7659), .A2(n7658), .ZN(n7657) );
  INV_X1 U8264 ( .A(n12121), .ZN(n7658) );
  INV_X1 U8265 ( .A(n7654), .ZN(n7650) );
  INV_X1 U8266 ( .A(n6971), .ZN(n6970) );
  OAI21_X1 U8267 ( .B1(n14203), .B2(n11475), .A(n11474), .ZN(n6971) );
  NAND2_X1 U8268 ( .A1(n11485), .A2(n11486), .ZN(n6743) );
  NOR2_X1 U8269 ( .A1(n6962), .A2(n6891), .ZN(n6804) );
  NAND2_X1 U8270 ( .A1(n7674), .A2(n12180), .ZN(n7673) );
  NAND2_X1 U8271 ( .A1(n11517), .A2(n6977), .ZN(n6976) );
  INV_X1 U8272 ( .A(n11518), .ZN(n6977) );
  INV_X1 U8273 ( .A(n11549), .ZN(n6756) );
  NAND2_X1 U8274 ( .A1(n11563), .A2(n7542), .ZN(n7541) );
  INV_X1 U8275 ( .A(n11562), .ZN(n7542) );
  NAND2_X1 U8276 ( .A1(n6773), .A2(n6770), .ZN(n12189) );
  OAI21_X1 U8277 ( .B1(n6757), .B2(n6755), .A(n7543), .ZN(n11576) );
  NAND2_X1 U8278 ( .A1(n7544), .A2(n11562), .ZN(n7543) );
  OAI21_X1 U8279 ( .B1(n11550), .B2(n11551), .A(n7541), .ZN(n6757) );
  AOI21_X1 U8280 ( .B1(n11550), .B2(n11551), .A(n6756), .ZN(n6755) );
  INV_X1 U8281 ( .A(n12192), .ZN(n7664) );
  NAND2_X1 U8282 ( .A1(n12202), .A2(n12201), .ZN(n7680) );
  INV_X1 U8283 ( .A(n12229), .ZN(n7241) );
  NOR2_X1 U8284 ( .A1(n11287), .A2(n6884), .ZN(n6883) );
  INV_X1 U8285 ( .A(n11285), .ZN(n6884) );
  NAND2_X1 U8286 ( .A1(n6844), .A2(n6846), .ZN(n6842) );
  OR2_X1 U8287 ( .A1(n10926), .A2(n10925), .ZN(n12970) );
  AND2_X1 U8288 ( .A1(n10905), .A2(n11988), .ZN(n7251) );
  NAND2_X1 U8289 ( .A1(n7254), .A2(n10905), .ZN(n7253) );
  INV_X1 U8290 ( .A(n11867), .ZN(n7254) );
  OAI21_X1 U8291 ( .B1(n6686), .B2(n7077), .A(n10582), .ZN(n7076) );
  NAND2_X1 U8292 ( .A1(n6570), .A2(n7241), .ZN(n7239) );
  INV_X1 U8293 ( .A(n7819), .ZN(n7138) );
  INV_X1 U8294 ( .A(n7943), .ZN(n7276) );
  OAI21_X1 U8295 ( .B1(n7277), .B2(n7276), .A(n10463), .ZN(n7275) );
  INV_X1 U8296 ( .A(n7429), .ZN(n7428) );
  INV_X1 U8297 ( .A(n11603), .ZN(n6758) );
  NOR2_X1 U8298 ( .A1(n6969), .A2(n11603), .ZN(n6759) );
  NAND2_X1 U8299 ( .A1(n9028), .A2(n7537), .ZN(n11367) );
  INV_X1 U8300 ( .A(n8249), .ZN(n7598) );
  NOR2_X1 U8301 ( .A1(n7806), .A2(SI_23_), .ZN(n7170) );
  OAI21_X1 U8302 ( .B1(n6544), .B2(n11222), .A(n7168), .ZN(n7167) );
  OR2_X1 U8303 ( .A1(n7791), .A2(n8104), .ZN(n7796) );
  NAND2_X1 U8304 ( .A1(n8066), .A2(n8065), .ZN(n8083) );
  AOI21_X1 U8305 ( .B1(n7155), .B2(n7157), .A(n7594), .ZN(n7153) );
  NAND2_X1 U8306 ( .A1(n6642), .A2(n7774), .ZN(n7595) );
  INV_X1 U8307 ( .A(n7158), .ZN(n7157) );
  INV_X1 U8308 ( .A(n7156), .ZN(n7155) );
  OAI21_X1 U8309 ( .B1(n7763), .B2(n7157), .A(n7770), .ZN(n7156) );
  NAND2_X1 U8310 ( .A1(n7848), .A2(n7734), .ZN(n6723) );
  INV_X1 U8311 ( .A(n6760), .ZN(n14382) );
  OAI21_X1 U8312 ( .B1(n14439), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6573), .ZN(
        n6760) );
  INV_X1 U8313 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14383) );
  NAND2_X1 U8314 ( .A1(n10524), .A2(n6677), .ZN(n10655) );
  INV_X1 U8315 ( .A(n6883), .ZN(n6878) );
  NAND2_X1 U8316 ( .A1(n11903), .A2(n11906), .ZN(n7248) );
  INV_X1 U8317 ( .A(n11911), .ZN(n7246) );
  NAND2_X1 U8318 ( .A1(n9875), .A2(n11832), .ZN(n15045) );
  OR2_X1 U8319 ( .A1(n11967), .A2(n7354), .ZN(n7353) );
  INV_X1 U8320 ( .A(n11961), .ZN(n7354) );
  INV_X1 U8321 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7257) );
  AND2_X1 U8322 ( .A1(n6580), .A2(n15368), .ZN(n7047) );
  OR2_X1 U8323 ( .A1(n8616), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U8324 ( .A1(n7344), .A2(n8589), .ZN(n8619) );
  INV_X1 U8325 ( .A(n7347), .ZN(n7346) );
  OAI21_X1 U8326 ( .B1(n8509), .B2(n7348), .A(n8518), .ZN(n7347) );
  INV_X1 U8327 ( .A(n7071), .ZN(n7070) );
  OAI21_X1 U8328 ( .B1(n8482), .B2(n7072), .A(n8490), .ZN(n7071) );
  INV_X1 U8329 ( .A(n8458), .ZN(n7072) );
  INV_X1 U8330 ( .A(n7481), .ZN(n6906) );
  NAND2_X1 U8331 ( .A1(n11110), .A2(n11109), .ZN(n6955) );
  OR2_X1 U8332 ( .A1(n13409), .A2(n8368), .ZN(n8357) );
  INV_X1 U8333 ( .A(n8186), .ZN(n8200) );
  NOR2_X1 U8334 ( .A1(n13571), .A2(n13739), .ZN(n6911) );
  INV_X1 U8335 ( .A(n7369), .ZN(n7368) );
  NOR2_X1 U8336 ( .A1(n7989), .A2(n10393), .ZN(n8005) );
  OR2_X1 U8337 ( .A1(n10771), .A2(n10772), .ZN(n10770) );
  OR2_X1 U8338 ( .A1(n7969), .A2(n15377), .ZN(n7989) );
  NOR2_X1 U8339 ( .A1(n7923), .A2(n7922), .ZN(n7937) );
  NAND2_X1 U8340 ( .A1(n6911), .A2(n6910), .ZN(n13558) );
  OR2_X1 U8341 ( .A1(n7932), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7933) );
  INV_X1 U8342 ( .A(n10326), .ZN(n7611) );
  INV_X1 U8343 ( .A(n7613), .ZN(n7608) );
  INV_X1 U8344 ( .A(n13850), .ZN(n7195) );
  INV_X1 U8345 ( .A(n13811), .ZN(n7642) );
  INV_X1 U8346 ( .A(n7639), .ZN(n7188) );
  AOI21_X1 U8347 ( .B1(n6541), .B2(n7641), .A(n7640), .ZN(n7639) );
  INV_X1 U8348 ( .A(n13894), .ZN(n7640) );
  INV_X1 U8349 ( .A(n13870), .ZN(n7641) );
  INV_X1 U8350 ( .A(n11639), .ZN(n7560) );
  NAND2_X1 U8351 ( .A1(n7493), .A2(n6822), .ZN(n6821) );
  INV_X1 U8352 ( .A(n14273), .ZN(n7493) );
  NAND2_X1 U8353 ( .A1(n7499), .A2(n11641), .ZN(n6823) );
  NAND2_X1 U8354 ( .A1(n11487), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11507) );
  NAND2_X1 U8355 ( .A1(n7398), .A2(n7395), .ZN(n7394) );
  INV_X1 U8356 ( .A(n14163), .ZN(n7395) );
  NOR2_X1 U8357 ( .A1(n14253), .A2(n14258), .ZN(n7498) );
  INV_X1 U8358 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U8359 ( .A1(n11363), .A2(n11367), .ZN(n11362) );
  NAND2_X1 U8360 ( .A1(n6711), .A2(n6604), .ZN(n14138) );
  NAND2_X1 U8361 ( .A1(n14182), .A2(n7388), .ZN(n6711) );
  NOR2_X1 U8362 ( .A1(n7389), .A2(n7397), .ZN(n7388) );
  NOR2_X2 U8363 ( .A1(n14226), .A2(n14332), .ZN(n14209) );
  OR2_X1 U8364 ( .A1(n14487), .A2(n14666), .ZN(n14253) );
  OR2_X1 U8365 ( .A1(n13957), .A2(n9919), .ZN(n11363) );
  INV_X1 U8366 ( .A(n8222), .ZN(n7603) );
  INV_X1 U8367 ( .A(n8231), .ZN(n8232) );
  AND2_X1 U8368 ( .A1(n7152), .A2(n6687), .ZN(n7148) );
  NAND2_X1 U8369 ( .A1(n7799), .A2(SI_21_), .ZN(n7801) );
  INV_X1 U8370 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9281) );
  AND2_X1 U8371 ( .A1(n7774), .A2(n7773), .ZN(n8015) );
  OR2_X1 U8372 ( .A1(n8630), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8661) );
  OR2_X1 U8373 ( .A1(n7762), .A2(n7761), .ZN(n7977) );
  AND2_X1 U8374 ( .A1(n8594), .A2(n8593), .ZN(n8624) );
  NAND2_X1 U8375 ( .A1(n7915), .A2(n7752), .ZN(n6721) );
  NAND2_X1 U8376 ( .A1(n7741), .A2(n7740), .ZN(n7889) );
  NAND2_X1 U8377 ( .A1(n9159), .A2(n8445), .ZN(n6939) );
  INV_X1 U8378 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U8379 ( .A1(n14379), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7468) );
  XNOR2_X1 U8380 ( .A(n14382), .B(n14383), .ZN(n14428) );
  NOR2_X1 U8381 ( .A1(n14393), .A2(n14392), .ZN(n14427) );
  NOR2_X1 U8382 ( .A1(n14449), .A2(n14391), .ZN(n14392) );
  OAI21_X1 U8383 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14397), .A(n14396), .ZN(
        n14423) );
  XNOR2_X1 U8384 ( .A(n11789), .B(n9878), .ZN(n9664) );
  INV_X1 U8385 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U8386 ( .A1(n15061), .A2(n11831), .ZN(n9875) );
  NAND2_X1 U8387 ( .A1(n9252), .A2(n15074), .ZN(n11832) );
  NAND2_X1 U8388 ( .A1(n12634), .A2(n6607), .ZN(n12593) );
  NOR2_X1 U8389 ( .A1(n7021), .A2(n7020), .ZN(n7019) );
  INV_X1 U8390 ( .A(n7526), .ZN(n7020) );
  AND2_X1 U8391 ( .A1(n10934), .A2(n8845), .ZN(n11022) );
  AND3_X1 U8392 ( .A1(n10695), .A2(n10694), .A3(n10693), .ZN(n11881) );
  INV_X1 U8393 ( .A(n7028), .ZN(n10709) );
  NAND2_X1 U8394 ( .A1(n11981), .A2(n11980), .ZN(n12018) );
  OR2_X1 U8395 ( .A1(n11950), .A2(n11936), .ZN(n7091) );
  OR2_X1 U8396 ( .A1(n11951), .A2(n11955), .ZN(n7090) );
  AOI21_X1 U8397 ( .B1(n7089), .B2(n12007), .A(n7087), .ZN(n11965) );
  OAI21_X1 U8398 ( .B1(n7088), .B2(n11936), .A(n11291), .ZN(n7087) );
  NAND2_X1 U8399 ( .A1(n11957), .A2(n11952), .ZN(n7089) );
  INV_X1 U8400 ( .A(n11954), .ZN(n7088) );
  INV_X1 U8401 ( .A(n15047), .ZN(n12684) );
  OR2_X1 U8402 ( .A1(n9127), .A2(n9126), .ZN(n9129) );
  OAI21_X1 U8403 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n9071), .A(n9129), .ZN(n9115) );
  AND2_X1 U8404 ( .A1(n7503), .A2(n7502), .ZN(n9064) );
  AND2_X1 U8405 ( .A1(n9063), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7502) );
  NOR2_X1 U8406 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  XNOR2_X1 U8407 ( .A(n9089), .B(n7513), .ZN(n9090) );
  NAND2_X1 U8408 ( .A1(n9098), .A2(n9099), .ZN(n9146) );
  NAND2_X1 U8409 ( .A1(n9297), .A2(n9298), .ZN(n9301) );
  AND2_X1 U8410 ( .A1(n9439), .A2(n9438), .ZN(n9606) );
  NAND2_X1 U8411 ( .A1(n9613), .A2(n9614), .ZN(n9615) );
  NAND2_X1 U8412 ( .A1(n14988), .A2(n9974), .ZN(n9975) );
  NAND2_X1 U8413 ( .A1(n9975), .A2(n9976), .ZN(n10524) );
  NAND2_X1 U8414 ( .A1(n12694), .A2(n12695), .ZN(n12698) );
  NAND2_X1 U8415 ( .A1(n12698), .A2(n12712), .ZN(n12724) );
  NAND2_X1 U8416 ( .A1(n14527), .A2(n12788), .ZN(n14545) );
  NOR2_X1 U8417 ( .A1(n14524), .A2(n12768), .ZN(n14556) );
  AND2_X1 U8418 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U8419 ( .A1(n14545), .A2(n14546), .ZN(n14544) );
  NOR2_X1 U8420 ( .A1(n12809), .A2(n15046), .ZN(n6946) );
  OR2_X1 U8421 ( .A1(n11250), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n11261) );
  AND2_X1 U8422 ( .A1(n11226), .A2(n11225), .ZN(n11237) );
  OAI21_X1 U8423 ( .B1(n6873), .B2(n6870), .A(n6868), .ZN(n12880) );
  AOI21_X1 U8424 ( .B1(n6871), .B2(n6869), .A(n6612), .ZN(n6868) );
  INV_X1 U8425 ( .A(n6566), .ZN(n6869) );
  NOR2_X1 U8426 ( .A1(n11214), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11226) );
  OR2_X1 U8427 ( .A1(n11203), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n11214) );
  INV_X1 U8428 ( .A(n12898), .ZN(n12918) );
  NOR2_X1 U8429 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n11180), .ZN(n11191) );
  AND2_X1 U8430 ( .A1(n11888), .A2(n11889), .ZN(n12979) );
  INV_X1 U8431 ( .A(n10907), .ZN(n15009) );
  AND2_X1 U8432 ( .A1(n10273), .A2(n10272), .ZN(n10275) );
  INV_X1 U8433 ( .A(n11828), .ZN(n9891) );
  AND4_X1 U8434 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n15019)
         );
  NAND2_X1 U8435 ( .A1(n7255), .A2(n11867), .ZN(n15016) );
  NAND2_X1 U8436 ( .A1(n10904), .A2(n11988), .ZN(n7255) );
  NOR2_X1 U8437 ( .A1(n10120), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10273) );
  OR2_X1 U8438 ( .A1(n9993), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U8439 ( .A1(n6706), .A2(n11850), .ZN(n10200) );
  OAI21_X1 U8440 ( .B1(n9901), .B2(n6705), .A(n6626), .ZN(n6706) );
  NOR2_X1 U8441 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9676) );
  NOR2_X1 U8442 ( .A1(n11984), .A2(n7213), .ZN(n6839) );
  NAND2_X1 U8443 ( .A1(n9889), .A2(n9888), .ZN(n9894) );
  NAND2_X1 U8444 ( .A1(n7208), .A2(n15068), .ZN(n6861) );
  AOI21_X1 U8445 ( .B1(n7208), .B2(n6860), .A(n11298), .ZN(n6859) );
  NOR2_X1 U8446 ( .A1(n6539), .A2(n15053), .ZN(n6860) );
  NAND2_X1 U8447 ( .A1(n6861), .A2(n15127), .ZN(n6853) );
  INV_X1 U8448 ( .A(n6859), .ZN(n6855) );
  NAND2_X1 U8449 ( .A1(n11260), .A2(n11259), .ZN(n13000) );
  OR2_X1 U8450 ( .A1(n11274), .A2(n11258), .ZN(n11259) );
  NAND2_X1 U8451 ( .A1(n12922), .A2(n11197), .ZN(n12905) );
  OR2_X1 U8452 ( .A1(n13096), .A2(n12962), .ZN(n12928) );
  OR2_X1 U8453 ( .A1(n12944), .A2(n12949), .ZN(n12945) );
  INV_X1 U8454 ( .A(n15054), .ZN(n15073) );
  OAI22_X1 U8455 ( .A1(n7355), .A2(n7353), .B1(n11966), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n7352) );
  NOR2_X1 U8456 ( .A1(n11959), .A2(n7356), .ZN(n7355) );
  INV_X1 U8457 ( .A(n11150), .ZN(n7356) );
  NAND2_X1 U8458 ( .A1(n10797), .A2(n10796), .ZN(n7093) );
  XNOR2_X1 U8459 ( .A(n8415), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U8460 ( .A1(n9059), .A2(n9058), .ZN(n10134) );
  NAND2_X1 U8461 ( .A1(n9343), .A2(n9342), .ZN(n9346) );
  NAND2_X1 U8462 ( .A1(n8858), .A2(n8408), .ZN(n9052) );
  OR2_X1 U8463 ( .A1(n8584), .A2(n8713), .ZN(n8530) );
  NAND2_X1 U8464 ( .A1(n8475), .A2(n8474), .ZN(n8532) );
  NAND2_X1 U8465 ( .A1(n8540), .A2(n8473), .ZN(n8475) );
  AND2_X1 U8466 ( .A1(n8536), .A2(n8537), .ZN(n8529) );
  NAND2_X1 U8467 ( .A1(n8521), .A2(n8471), .ZN(n8540) );
  AND2_X1 U8468 ( .A1(n8450), .A2(n8449), .ZN(n8524) );
  INV_X1 U8469 ( .A(n6567), .ZN(n7121) );
  INV_X1 U8470 ( .A(n13152), .ZN(n7474) );
  INV_X1 U8471 ( .A(n7478), .ZN(n7476) );
  NAND2_X1 U8472 ( .A1(n8070), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8096) );
  OR2_X1 U8473 ( .A1(n7952), .A2(n11802), .ZN(n7969) );
  INV_X1 U8474 ( .A(n7479), .ZN(n7127) );
  NAND2_X1 U8475 ( .A1(n12315), .A2(n6958), .ZN(n12311) );
  OR2_X1 U8476 ( .A1(n12316), .A2(n12310), .ZN(n6958) );
  OR2_X1 U8477 ( .A1(n8024), .A2(n8023), .ZN(n8036) );
  OR2_X1 U8478 ( .A1(n8161), .A2(n13156), .ZN(n8174) );
  NOR2_X1 U8479 ( .A1(n8174), .A2(n13220), .ZN(n8187) );
  INV_X1 U8480 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10393) );
  AND3_X1 U8481 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n7907) );
  AND2_X1 U8482 ( .A1(n12301), .A2(n12305), .ZN(n9324) );
  NOR2_X1 U8483 ( .A1(n8036), .A2(n13312), .ZN(n8057) );
  AND2_X1 U8484 ( .A1(n8057), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8070) );
  XNOR2_X1 U8485 ( .A(n7588), .B(n6527), .ZN(n7587) );
  INV_X1 U8486 ( .A(n12260), .ZN(n6986) );
  NOR2_X1 U8487 ( .A1(n12257), .A2(n12258), .ZN(n7234) );
  INV_X1 U8488 ( .A(n6525), .ZN(n8255) );
  OR2_X1 U8489 ( .A1(n7857), .A2(n7822), .ZN(n7823) );
  NAND2_X1 U8490 ( .A1(n8964), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U8491 ( .A1(n8973), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U8492 ( .A1(n9628), .A2(n7011), .ZN(n14842) );
  AND2_X1 U8493 ( .A1(n9634), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U8494 ( .A1(n14842), .A2(n14841), .ZN(n14840) );
  NOR2_X1 U8495 ( .A1(n14840), .A2(n7010), .ZN(n13285) );
  AND2_X1 U8496 ( .A1(n9635), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U8497 ( .A1(n13285), .A2(n13284), .ZN(n13283) );
  INV_X1 U8498 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U8499 ( .A1(n9846), .A2(n7005), .ZN(n9849) );
  NOR2_X1 U8500 ( .A1(n9637), .A2(n9627), .ZN(n7005) );
  NOR2_X1 U8501 ( .A1(n9849), .A2(n9848), .ZN(n11065) );
  NOR2_X1 U8502 ( .A1(n11065), .A2(n7004), .ZN(n13298) );
  AND2_X1 U8503 ( .A1(n11066), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8504 ( .A1(n13298), .A2(n13299), .ZN(n13297) );
  INV_X1 U8505 ( .A(n7440), .ZN(n7432) );
  NAND2_X1 U8506 ( .A1(n7437), .A2(n7440), .ZN(n7433) );
  AOI21_X1 U8507 ( .B1(n7436), .B2(n7437), .A(n12261), .ZN(n7435) );
  AND2_X1 U8508 ( .A1(n13440), .A2(n13243), .ZN(n7289) );
  NAND2_X1 U8509 ( .A1(n13718), .A2(n7139), .ZN(n7290) );
  AOI21_X1 U8510 ( .B1(n7280), .B2(n6559), .A(n6551), .ZN(n7279) );
  NOR2_X1 U8511 ( .A1(n8117), .A2(n8116), .ZN(n8136) );
  OR2_X1 U8512 ( .A1(n13549), .A2(n8340), .ZN(n8342) );
  AOI21_X1 U8513 ( .B1(n12285), .B2(n7285), .A(n6678), .ZN(n7284) );
  INV_X1 U8514 ( .A(n6911), .ZN(n13572) );
  INV_X1 U8515 ( .A(n13191), .ZN(n13231) );
  NAND2_X1 U8516 ( .A1(n10818), .A2(n7369), .ZN(n10998) );
  NAND2_X1 U8517 ( .A1(n10818), .A2(n10897), .ZN(n10888) );
  AOI21_X1 U8518 ( .B1(n8326), .B2(n10772), .A(n7450), .ZN(n7449) );
  NAND2_X1 U8519 ( .A1(n10770), .A2(n8326), .ZN(n10821) );
  NOR2_X1 U8520 ( .A1(n6625), .A2(n7269), .ZN(n7268) );
  AOI21_X1 U8521 ( .B1(n7457), .B2(n8322), .A(n6622), .ZN(n7456) );
  NOR2_X1 U8522 ( .A1(n12269), .A2(n7273), .ZN(n7271) );
  NOR2_X2 U8523 ( .A1(n14898), .A2(n14936), .ZN(n10180) );
  AND2_X1 U8524 ( .A1(n8090), .A2(n7489), .ZN(n7488) );
  INV_X1 U8525 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7489) );
  INV_X1 U8526 ( .A(n9533), .ZN(n9453) );
  NAND2_X1 U8527 ( .A1(n12038), .A2(n8359), .ZN(n14892) );
  AND2_X1 U8528 ( .A1(n10068), .A2(n14955), .ZN(n13699) );
  NAND2_X1 U8529 ( .A1(n6942), .A2(n7929), .ZN(n10403) );
  INV_X2 U8530 ( .A(n8171), .ZN(n12230) );
  AND2_X1 U8531 ( .A1(n12304), .A2(n9323), .ZN(n14953) );
  INV_X1 U8532 ( .A(n11321), .ZN(n7586) );
  NOR2_X1 U8533 ( .A1(n11323), .A2(n11316), .ZN(n7585) );
  AND2_X1 U8534 ( .A1(n8263), .A2(n7297), .ZN(n7675) );
  AND2_X1 U8535 ( .A1(n7298), .A2(n6661), .ZN(n7297) );
  NAND2_X1 U8536 ( .A1(n8091), .A2(n8090), .ZN(n8130) );
  OR2_X1 U8537 ( .A1(n8001), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8032) );
  AND2_X1 U8538 ( .A1(n8804), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8571) );
  NAND2_X1 U8539 ( .A1(n7634), .A2(n13879), .ZN(n7182) );
  INV_X1 U8540 ( .A(n7180), .ZN(n7179) );
  INV_X1 U8541 ( .A(n11519), .ZN(n11520) );
  NAND2_X1 U8542 ( .A1(n11520), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11541) );
  AOI21_X1 U8543 ( .B1(n13771), .B2(n12540), .A(n12550), .ZN(n7632) );
  INV_X1 U8544 ( .A(n7632), .ZN(n7630) );
  NOR2_X1 U8545 ( .A1(n9775), .A2(n9774), .ZN(n9937) );
  NAND2_X1 U8546 ( .A1(n7617), .A2(n7616), .ZN(n7615) );
  NAND2_X1 U8547 ( .A1(n13923), .A2(n13922), .ZN(n7638) );
  AND3_X1 U8548 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U8549 ( .A1(n12463), .A2(n13850), .ZN(n13853) );
  OR2_X1 U8550 ( .A1(n11459), .A2(n11458), .ZN(n11461) );
  NAND2_X1 U8551 ( .A1(n13791), .A2(n13861), .ZN(n7621) );
  CLKBUF_X1 U8552 ( .A(n12543), .Z(n6907) );
  INV_X1 U8553 ( .A(n8824), .ZN(n6922) );
  AND2_X1 U8554 ( .A1(n11476), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U8555 ( .A1(n7643), .A2(n6541), .ZN(n13809) );
  INV_X1 U8556 ( .A(n11507), .ZN(n11508) );
  NOR2_X1 U8557 ( .A1(n10225), .A2(n10224), .ZN(n10349) );
  NAND2_X1 U8558 ( .A1(n13853), .A2(n12464), .ZN(n13901) );
  NAND2_X1 U8559 ( .A1(n11565), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11592) );
  NOR2_X1 U8560 ( .A1(n10618), .A2(n10617), .ZN(n10740) );
  NOR2_X1 U8561 ( .A1(n7558), .A2(n7556), .ZN(n7555) );
  NAND2_X1 U8562 ( .A1(n7557), .A2(n11679), .ZN(n7556) );
  INV_X1 U8563 ( .A(n11687), .ZN(n7557) );
  INV_X1 U8564 ( .A(n7558), .ZN(n7554) );
  INV_X1 U8565 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14378) );
  NAND2_X1 U8566 ( .A1(n9588), .A2(n6832), .ZN(n13998) );
  OR2_X1 U8567 ( .A1(n10346), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8568 ( .A1(n13998), .A2(n13999), .ZN(n13997) );
  OR2_X1 U8569 ( .A1(n10828), .A2(n10834), .ZN(n6830) );
  NAND2_X1 U8570 ( .A1(n14055), .A2(n14042), .ZN(n7337) );
  INV_X1 U8571 ( .A(n7412), .ZN(n6726) );
  NOR2_X1 U8572 ( .A1(n14101), .A2(n7414), .ZN(n6727) );
  NAND2_X1 U8573 ( .A1(n14289), .A2(n13934), .ZN(n7339) );
  NAND2_X1 U8574 ( .A1(n7417), .A2(n7418), .ZN(n14057) );
  NOR2_X1 U8575 ( .A1(n14106), .A2(n14289), .ZN(n14095) );
  NAND2_X1 U8576 ( .A1(n14294), .A2(n11716), .ZN(n14087) );
  NAND2_X1 U8577 ( .A1(n14128), .A2(n14107), .ZN(n14106) );
  NOR2_X1 U8578 ( .A1(n14117), .A2(n6961), .ZN(n14103) );
  AND2_X1 U8579 ( .A1(n14132), .A2(n13936), .ZN(n6961) );
  OAI22_X1 U8580 ( .A1(n14138), .A2(n14137), .B1(n7499), .B2(n13937), .ZN(
        n14118) );
  NOR2_X1 U8581 ( .A1(n14150), .A2(n7391), .ZN(n7390) );
  NAND2_X1 U8582 ( .A1(n7394), .A2(n7392), .ZN(n7391) );
  INV_X1 U8583 ( .A(n14151), .ZN(n7392) );
  NAND2_X1 U8584 ( .A1(n14182), .A2(n7396), .ZN(n7393) );
  NAND2_X1 U8585 ( .A1(n7393), .A2(n7394), .ZN(n14166) );
  NAND2_X1 U8586 ( .A1(n14182), .A2(n14181), .ZN(n14180) );
  AND2_X1 U8587 ( .A1(n11355), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11476) );
  INV_X1 U8588 ( .A(n14199), .ZN(n14203) );
  AND2_X1 U8589 ( .A1(n11473), .A2(n11698), .ZN(n14199) );
  AOI21_X1 U8590 ( .B1(n7342), .B2(n11705), .A(n6621), .ZN(n7340) );
  AND2_X1 U8591 ( .A1(n10740), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10744) );
  INV_X1 U8592 ( .A(n7498), .ZN(n14254) );
  AOI21_X1 U8593 ( .B1(n14248), .B2(n14260), .A(n10736), .ZN(n11695) );
  AOI21_X1 U8594 ( .B1(n11661), .B2(n7328), .A(n6618), .ZN(n7327) );
  INV_X1 U8595 ( .A(n13944), .ZN(n14249) );
  OR2_X1 U8596 ( .A1(n10603), .A2(n10602), .ZN(n10618) );
  NAND2_X1 U8597 ( .A1(n14488), .A2(n14506), .ZN(n14487) );
  AOI21_X1 U8598 ( .B1(n7302), .B2(n7305), .A(n6620), .ZN(n7299) );
  INV_X1 U8599 ( .A(n10343), .ZN(n7406) );
  OR2_X1 U8600 ( .A1(n10042), .A2(n10041), .ZN(n10225) );
  OR2_X1 U8601 ( .A1(n10030), .A2(n10029), .ZN(n10042) );
  NAND2_X1 U8602 ( .A1(n7317), .A2(n7320), .ZN(n7314) );
  NAND2_X1 U8603 ( .A1(n7421), .A2(n7423), .ZN(n9749) );
  NAND2_X1 U8604 ( .A1(n6635), .A2(n7424), .ZN(n7423) );
  INV_X1 U8605 ( .A(n6564), .ZN(n7424) );
  INV_X1 U8606 ( .A(n9652), .ZN(n6814) );
  OR2_X1 U8607 ( .A1(n14637), .A2(n11352), .ZN(n14496) );
  NAND2_X1 U8608 ( .A1(n9233), .A2(n9232), .ZN(n9384) );
  NAND2_X1 U8609 ( .A1(n14752), .A2(n9919), .ZN(n9652) );
  NOR2_X1 U8610 ( .A1(n11372), .A2(n9652), .ZN(n9395) );
  NAND2_X1 U8611 ( .A1(n9655), .A2(n6964), .ZN(n9648) );
  INV_X1 U8612 ( .A(n9650), .ZN(n6964) );
  CLKBUF_X1 U8613 ( .A(n11644), .Z(n6896) );
  INV_X1 U8614 ( .A(n11635), .ZN(n11309) );
  INV_X1 U8615 ( .A(n10051), .ZN(n10058) );
  NAND2_X1 U8616 ( .A1(n14496), .A2(n14764), .ZN(n14796) );
  NAND2_X1 U8617 ( .A1(n8600), .A2(n8384), .ZN(n8387) );
  INV_X1 U8618 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U8619 ( .A1(n7605), .A2(n7798), .ZN(n8156) );
  XNOR2_X1 U8620 ( .A(n8129), .B(n8128), .ZN(n11351) );
  XNOR2_X1 U8621 ( .A(n8124), .B(SI_18_), .ZN(n8109) );
  OAI21_X1 U8622 ( .B1(n8031), .B2(n6715), .A(n6714), .ZN(n6713) );
  NAND2_X1 U8623 ( .A1(n8031), .A2(n6716), .ZN(n6712) );
  NAND2_X1 U8624 ( .A1(n7160), .A2(n7158), .ZN(n7999) );
  AND2_X1 U8625 ( .A1(n7160), .A2(n7979), .ZN(n7997) );
  AND2_X1 U8626 ( .A1(n6762), .A2(n6761), .ZN(n15387) );
  NOR2_X1 U8627 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_REG2_REG_25__SCAN_IN), 
        .ZN(n6762) );
  NOR2_X1 U8628 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), 
        .ZN(n6761) );
  INV_X1 U8629 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9675) );
  AOI21_X1 U8630 ( .B1(n6753), .B2(n14433), .A(n7469), .ZN(n14431) );
  AND2_X1 U8631 ( .A1(n14378), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7469) );
  XOR2_X1 U8632 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14430) );
  XNOR2_X1 U8633 ( .A(n14428), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14429) );
  XNOR2_X1 U8634 ( .A(n14442), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14443) );
  NOR2_X1 U8635 ( .A1(n14387), .A2(n14386), .ZN(n14446) );
  NOR2_X1 U8636 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14442), .ZN(n14386) );
  NAND2_X1 U8637 ( .A1(n7098), .A2(n14451), .ZN(n14452) );
  NAND2_X1 U8638 ( .A1(n7465), .A2(n14458), .ZN(n14459) );
  AOI21_X1 U8639 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14402), .A(n14401), .ZN(
        n14461) );
  OAI21_X1 U8640 ( .B1(n7105), .B2(n6754), .A(n7461), .ZN(n7460) );
  NAND2_X1 U8641 ( .A1(n7042), .A2(n7041), .ZN(n12572) );
  AOI21_X1 U8642 ( .B1(n6540), .B2(n7045), .A(n7519), .ZN(n7041) );
  NAND2_X1 U8643 ( .A1(n9542), .A2(n7527), .ZN(n9665) );
  NAND2_X1 U8644 ( .A1(n11179), .A2(n11178), .ZN(n12940) );
  INV_X1 U8645 ( .A(n7518), .ZN(n7517) );
  NAND2_X1 U8646 ( .A1(n15063), .A2(n9432), .ZN(n15066) );
  NAND2_X1 U8647 ( .A1(n12634), .A2(n11766), .ZN(n12595) );
  INV_X1 U8648 ( .A(n12975), .ZN(n10976) );
  AOI21_X1 U8649 ( .B1(n10709), .B2(n7535), .A(n7534), .ZN(n10864) );
  NAND2_X1 U8650 ( .A1(n7043), .A2(n11780), .ZN(n12602) );
  NAND2_X1 U8651 ( .A1(n12627), .A2(n12628), .ZN(n7043) );
  NAND2_X1 U8652 ( .A1(n7038), .A2(n11752), .ZN(n12611) );
  OR2_X1 U8653 ( .A1(n11754), .A2(n11753), .ZN(n7038) );
  NAND2_X1 U8654 ( .A1(n7034), .A2(n7039), .ZN(n12609) );
  NAND2_X1 U8655 ( .A1(n11754), .A2(n11752), .ZN(n7034) );
  INV_X1 U8656 ( .A(n9542), .ZN(n7025) );
  NAND2_X1 U8657 ( .A1(n7015), .A2(n9984), .ZN(n7024) );
  NAND2_X1 U8658 ( .A1(n7033), .A2(n7031), .ZN(n12618) );
  AOI21_X1 U8659 ( .B1(n7035), .B2(n7037), .A(n7032), .ZN(n7031) );
  INV_X1 U8660 ( .A(n12619), .ZN(n7032) );
  NAND2_X1 U8661 ( .A1(n7030), .A2(n7035), .ZN(n12620) );
  OR2_X1 U8662 ( .A1(n11754), .A2(n7037), .ZN(n7030) );
  NAND2_X1 U8663 ( .A1(n9665), .A2(n7526), .ZN(n9674) );
  OAI21_X1 U8664 ( .B1(n10292), .B2(n10291), .A(n10290), .ZN(n10293) );
  NAND2_X1 U8665 ( .A1(n12636), .A2(n12635), .ZN(n12634) );
  AND4_X1 U8666 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n10974) );
  NAND2_X1 U8667 ( .A1(n7027), .A2(n7026), .ZN(n10980) );
  NAND2_X1 U8668 ( .A1(n7533), .A2(n10866), .ZN(n7026) );
  NAND2_X1 U8669 ( .A1(n7028), .A2(n6608), .ZN(n7027) );
  NAND2_X1 U8670 ( .A1(n10870), .A2(n10869), .ZN(n14568) );
  AND4_X1 U8671 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n14581) );
  INV_X1 U8672 ( .A(n11881), .ZN(n14583) );
  NAND2_X1 U8673 ( .A1(n9479), .A2(n9478), .ZN(n9543) );
  OR2_X1 U8674 ( .A1(n9477), .A2(n12685), .ZN(n9478) );
  NAND2_X1 U8675 ( .A1(n9543), .A2(n9544), .ZN(n9542) );
  INV_X1 U8676 ( .A(n12672), .ZN(n12651) );
  AND4_X1 U8677 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n12871) );
  NAND2_X1 U8678 ( .A1(n11783), .A2(n11782), .ZN(n12661) );
  NAND4_X1 U8679 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n12837) );
  INV_X1 U8680 ( .A(n12871), .ZN(n12838) );
  INV_X1 U8681 ( .A(n12962), .ZN(n12677) );
  INV_X1 U8682 ( .A(n11033), .ZN(n12678) );
  INV_X1 U8683 ( .A(n10974), .ZN(n14564) );
  INV_X1 U8684 ( .A(n14581), .ZN(n14563) );
  NAND4_X1 U8685 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n15000) );
  NAND4_X1 U8686 ( .A1(n10261), .A2(n10260), .A3(n10259), .A4(n10258), .ZN(
        n15001) );
  INV_X1 U8687 ( .A(n10445), .ZN(n12680) );
  INV_X1 U8688 ( .A(n10281), .ZN(n12681) );
  INV_X1 U8689 ( .A(n11847), .ZN(n12683) );
  CLKBUF_X1 U8690 ( .A(n12684), .Z(n6954) );
  NAND2_X1 U8691 ( .A1(n7503), .A2(n9063), .ZN(n9125) );
  NOR2_X1 U8692 ( .A1(n6763), .A2(n15181), .ZN(n9276) );
  INV_X1 U8693 ( .A(n9271), .ZN(n6763) );
  INV_X1 U8694 ( .A(n7060), .ZN(n9143) );
  OR2_X1 U8695 ( .A1(n9292), .A2(n9293), .ZN(n7508) );
  NAND2_X1 U8696 ( .A1(n7058), .A2(n6694), .ZN(n9439) );
  XNOR2_X1 U8697 ( .A(n9606), .B(n10263), .ZN(n9607) );
  INV_X1 U8698 ( .A(n7065), .ZN(n9955) );
  NOR2_X1 U8699 ( .A1(n14973), .A2(n9957), .ZN(n9959) );
  OAI21_X1 U8700 ( .B1(n10523), .B2(n7062), .A(n7061), .ZN(n10955) );
  NAND2_X1 U8701 ( .A1(n7063), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7062) );
  NOR2_X1 U8702 ( .A1(n10956), .A2(n10957), .ZN(n12688) );
  NOR2_X1 U8703 ( .A1(n12709), .A2(n10957), .ZN(n7057) );
  NOR2_X1 U8704 ( .A1(n12688), .A2(n12689), .ZN(n12691) );
  OR2_X1 U8705 ( .A1(n12765), .A2(n14529), .ZN(n7049) );
  NOR2_X1 U8706 ( .A1(n14525), .A2(n14526), .ZN(n14524) );
  NAND2_X1 U8707 ( .A1(n8858), .A2(n6580), .ZN(n9208) );
  OR2_X1 U8708 ( .A1(n12383), .A2(n12968), .ZN(n6990) );
  NAND2_X1 U8709 ( .A1(n11281), .A2(n11280), .ZN(n12959) );
  NAND2_X1 U8710 ( .A1(n11021), .A2(n11020), .ZN(n13037) );
  AND2_X1 U8711 ( .A1(n14999), .A2(n11878), .ZN(n10909) );
  NAND2_X1 U8712 ( .A1(n6703), .A2(n11841), .ZN(n10129) );
  NAND2_X1 U8713 ( .A1(n9901), .A2(n11984), .ZN(n6703) );
  AND2_X1 U8714 ( .A1(n9431), .A2(n15040), .ZN(n15083) );
  AND2_X1 U8715 ( .A1(n15028), .A2(n15073), .ZN(n15038) );
  AND2_X1 U8716 ( .A1(n15142), .A2(n15073), .ZN(n13029) );
  INV_X1 U8717 ( .A(n12986), .ZN(n13043) );
  INV_X1 U8718 ( .A(n12015), .ZN(n13046) );
  NAND2_X1 U8719 ( .A1(n11271), .A2(n11270), .ZN(n13053) );
  AOI21_X1 U8720 ( .B1(n12829), .B2(n15068), .A(n6927), .ZN(n13051) );
  NAND2_X1 U8721 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U8722 ( .A1(n12855), .A2(n15062), .ZN(n6928) );
  NAND2_X1 U8723 ( .A1(n11249), .A2(n11248), .ZN(n13060) );
  AND2_X1 U8724 ( .A1(n12857), .A2(n12856), .ZN(n13058) );
  NAND2_X1 U8725 ( .A1(n6872), .A2(n6875), .ZN(n12897) );
  AND2_X1 U8726 ( .A1(n6865), .A2(n11814), .ZN(n6875) );
  NAND2_X1 U8727 ( .A1(n6874), .A2(n11284), .ZN(n12906) );
  NAND2_X1 U8728 ( .A1(n12915), .A2(n12919), .ZN(n6874) );
  NAND2_X1 U8729 ( .A1(n7261), .A2(n7262), .ZN(n12920) );
  NAND2_X1 U8730 ( .A1(n6843), .A2(n6847), .ZN(n12950) );
  NAND2_X1 U8731 ( .A1(n11281), .A2(n6849), .ZN(n6843) );
  NAND2_X1 U8732 ( .A1(n7247), .A2(n11906), .ZN(n11159) );
  NAND2_X1 U8733 ( .A1(n11038), .A2(n11999), .ZN(n7247) );
  NAND2_X1 U8734 ( .A1(n11008), .A2(n11007), .ZN(n11049) );
  NAND2_X1 U8735 ( .A1(n10914), .A2(n10913), .ZN(n11029) );
  INV_X1 U8736 ( .A(n9061), .ZN(n11729) );
  INV_X1 U8737 ( .A(n7352), .ZN(n7351) );
  INV_X1 U8738 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U8739 ( .A1(n7350), .A2(n11961), .ZN(n11968) );
  OAI21_X1 U8740 ( .B1(n9049), .B2(P3_IR_REG_28__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U8741 ( .A1(n9049), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6709) );
  XNOR2_X1 U8742 ( .A(n8413), .B(P3_IR_REG_26__SCAN_IN), .ZN(n10800) );
  NAND2_X1 U8743 ( .A1(n7530), .A2(n7258), .ZN(n8710) );
  AND2_X1 U8744 ( .A1(n8543), .A2(n8412), .ZN(n7258) );
  NAND2_X1 U8745 ( .A1(n10765), .A2(n10587), .ZN(n10764) );
  NAND2_X1 U8746 ( .A1(n7074), .A2(n10370), .ZN(n10583) );
  NAND2_X1 U8747 ( .A1(n10187), .A2(n6686), .ZN(n7074) );
  NAND2_X1 U8748 ( .A1(n10187), .A2(n10186), .ZN(n10369) );
  INV_X1 U8749 ( .A(n10134), .ZN(n12034) );
  XNOR2_X1 U8750 ( .A(n9055), .B(n9054), .ZN(n11828) );
  OAI21_X1 U8751 ( .B1(n9177), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U8752 ( .A1(n9835), .A2(n9834), .ZN(n9838) );
  INV_X1 U8753 ( .A(SI_20_), .ZN(n11187) );
  XNOR2_X1 U8754 ( .A(n9178), .B(n9179), .ZN(n9690) );
  NAND2_X1 U8755 ( .A1(n7080), .A2(n9212), .ZN(n9215) );
  INV_X1 U8756 ( .A(SI_17_), .ZN(n9039) );
  NAND2_X1 U8757 ( .A1(n9037), .A2(n9036), .ZN(n9211) );
  INV_X1 U8758 ( .A(SI_16_), .ZN(n8867) );
  INV_X1 U8759 ( .A(SI_13_), .ZN(n8591) );
  INV_X1 U8760 ( .A(SI_12_), .ZN(n10712) );
  OR2_X1 U8761 ( .A1(n8536), .A2(n8713), .ZN(n8538) );
  NAND2_X1 U8762 ( .A1(n8512), .A2(n8469), .ZN(n8519) );
  NAND2_X1 U8763 ( .A1(n8464), .A2(n8463), .ZN(n8504) );
  NAND2_X1 U8764 ( .A1(n7069), .A2(n8458), .ZN(n8491) );
  NAND2_X1 U8765 ( .A1(n8483), .A2(n8482), .ZN(n7069) );
  INV_X1 U8766 ( .A(n9668), .ZN(n9094) );
  NAND2_X1 U8767 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7051) );
  NAND2_X1 U8768 ( .A1(n8713), .A2(n8523), .ZN(n7052) );
  NAND2_X1 U8769 ( .A1(n9065), .A2(n8523), .ZN(n7050) );
  NAND2_X1 U8770 ( .A1(n7505), .A2(n8441), .ZN(n9251) );
  INV_X1 U8771 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15181) );
  INV_X1 U8772 ( .A(n6956), .ZN(n11108) );
  INV_X1 U8773 ( .A(n6988), .ZN(n13133) );
  NAND2_X1 U8774 ( .A1(n6989), .A2(n7478), .ZN(n10381) );
  NAND2_X1 U8775 ( .A1(n9568), .A2(n9576), .ZN(n9569) );
  OR2_X1 U8776 ( .A1(n14813), .A2(n12345), .ZN(n13213) );
  AND2_X1 U8777 ( .A1(n7119), .A2(n7118), .ZN(n7113) );
  OAI21_X1 U8778 ( .B1(n7119), .B2(n12402), .A(n7115), .ZN(n7114) );
  NAND2_X1 U8779 ( .A1(n7119), .A2(n7116), .ZN(n7115) );
  NAND2_X1 U8780 ( .A1(n7121), .A2(n7118), .ZN(n7116) );
  OR2_X1 U8781 ( .A1(n7121), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U8782 ( .A1(n8899), .A2(n6601), .ZN(n7834) );
  NAND2_X1 U8783 ( .A1(n13212), .A2(n12337), .ZN(n13153) );
  NAND2_X1 U8784 ( .A1(n12311), .A2(n12317), .ZN(n12327) );
  CLKBUF_X1 U8785 ( .A(n11813), .Z(n6989) );
  NAND2_X1 U8786 ( .A1(n7122), .A2(n7125), .ZN(n13212) );
  OR2_X1 U8787 ( .A1(n12311), .A2(n7127), .ZN(n7122) );
  NAND2_X1 U8788 ( .A1(n11141), .A2(n7109), .ZN(n14814) );
  OR2_X1 U8789 ( .A1(n10564), .A2(n10565), .ZN(n7109) );
  NOR2_X1 U8790 ( .A1(n14814), .A2(n14815), .ZN(n14812) );
  NOR2_X1 U8791 ( .A1(n13214), .A2(n12345), .ZN(n7110) );
  AND2_X1 U8792 ( .A1(n7477), .A2(n6560), .ZN(n11137) );
  INV_X1 U8793 ( .A(n7477), .ZN(n10392) );
  XNOR2_X1 U8794 ( .A(n11134), .B(n10561), .ZN(n10397) );
  NAND2_X1 U8795 ( .A1(n9336), .A2(n9332), .ZN(n14811) );
  NAND2_X1 U8796 ( .A1(n12327), .A2(n7481), .ZN(n13228) );
  INV_X1 U8797 ( .A(n12308), .ZN(n6798) );
  OR2_X1 U8798 ( .A1(n8101), .A2(n8100), .ZN(n13252) );
  OR2_X1 U8799 ( .A1(n8256), .A2(n7839), .ZN(n7841) );
  OR2_X1 U8800 ( .A1(n7857), .A2(n9040), .ZN(n6890) );
  NAND2_X1 U8801 ( .A1(n6893), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7644) );
  INV_X1 U8802 ( .A(n7007), .ZN(n8955) );
  NAND2_X1 U8803 ( .A1(n9007), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6996) );
  INV_X1 U8804 ( .A(n6995), .ZN(n8972) );
  NOR2_X1 U8805 ( .A1(n11070), .A2(n13330), .ZN(n11072) );
  XNOR2_X1 U8806 ( .A(n13394), .B(n7372), .ZN(n13387) );
  NAND2_X1 U8807 ( .A1(n7434), .A2(n7437), .ZN(n13415) );
  NAND2_X1 U8808 ( .A1(n13444), .A2(n7438), .ZN(n7434) );
  AOI21_X1 U8809 ( .B1(n13444), .B2(n13457), .A(n8355), .ZN(n13429) );
  NAND2_X1 U8810 ( .A1(n7296), .A2(n7294), .ZN(n13465) );
  OR2_X1 U8811 ( .A1(n10416), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U8812 ( .A1(n13522), .A2(n8346), .ZN(n13507) );
  NAND2_X1 U8813 ( .A1(n7281), .A2(n7282), .ZN(n13526) );
  OR2_X1 U8814 ( .A1(n6967), .A2(n6559), .ZN(n7281) );
  NAND2_X1 U8815 ( .A1(n13535), .A2(n8344), .ZN(n13520) );
  NAND2_X1 U8816 ( .A1(n6967), .A2(n8123), .ZN(n13534) );
  NAND2_X1 U8817 ( .A1(n11099), .A2(n8336), .ZN(n13568) );
  NAND2_X1 U8818 ( .A1(n7287), .A2(n7285), .ZN(n11097) );
  NAND2_X1 U8819 ( .A1(n7287), .A2(n8064), .ZN(n11095) );
  NAND2_X1 U8820 ( .A1(n7270), .A2(n7976), .ZN(n10769) );
  NAND2_X1 U8821 ( .A1(n7458), .A2(n7457), .ZN(n10467) );
  NAND2_X1 U8822 ( .A1(n7458), .A2(n8323), .ZN(n10464) );
  NAND2_X1 U8823 ( .A1(n10401), .A2(n7943), .ZN(n10462) );
  NAND2_X1 U8824 ( .A1(n7272), .A2(n7896), .ZN(n10069) );
  NAND2_X1 U8825 ( .A1(n10174), .A2(n8315), .ZN(n10101) );
  INV_X1 U8826 ( .A(n13600), .ZN(n14879) );
  INV_X1 U8827 ( .A(n7852), .ZN(n10169) );
  INV_X1 U8828 ( .A(n14874), .ZN(n13578) );
  INV_X1 U8829 ( .A(n13396), .ZN(n13707) );
  INV_X1 U8830 ( .A(n13621), .ZN(n7163) );
  INV_X1 U8831 ( .A(n7718), .ZN(n12375) );
  NAND2_X1 U8832 ( .A1(n6796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U8833 ( .A1(n8263), .A2(n6795), .ZN(n6796) );
  AND2_X1 U8834 ( .A1(n7298), .A2(n6655), .ZN(n6795) );
  XNOR2_X1 U8835 ( .A(n8275), .B(n7713), .ZN(n13767) );
  OR2_X1 U8836 ( .A1(n8273), .A2(n8272), .ZN(n10954) );
  INV_X1 U8837 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10419) );
  INV_X1 U8838 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8303) );
  AOI21_X1 U8839 ( .B1(n7484), .B2(n7486), .A(n6641), .ZN(n7482) );
  NAND2_X1 U8840 ( .A1(n8091), .A2(n7484), .ZN(n7483) );
  INV_X1 U8841 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9286) );
  INV_X1 U8842 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9419) );
  INV_X1 U8843 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9315) );
  INV_X1 U8844 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n8874) );
  INV_X1 U8845 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8629) );
  INV_X1 U8846 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8628) );
  INV_X1 U8847 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8592) );
  INV_X1 U8848 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8560) );
  INV_X1 U8849 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8558) );
  INV_X1 U8850 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8555) );
  INV_X1 U8851 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8559) );
  INV_X1 U8852 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8556) );
  OAI22_X1 U8853 ( .A1(n7844), .A2(n7012), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        P2_IR_REG_2__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U8854 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7012) );
  INV_X1 U8855 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U8856 ( .A1(n10320), .A2(n7175), .ZN(n7174) );
  INV_X1 U8857 ( .A(n10322), .ZN(n7175) );
  NAND2_X1 U8858 ( .A1(n10327), .A2(n10326), .ZN(n10499) );
  NAND2_X1 U8859 ( .A1(n10499), .A2(n7615), .ZN(n10502) );
  NAND2_X1 U8860 ( .A1(n7643), .A2(n12483), .ZN(n13812) );
  NAND2_X1 U8861 ( .A1(n11499), .A2(n11498), .ZN(n14319) );
  OR2_X1 U8862 ( .A1(n11497), .A2(n11496), .ZN(n11499) );
  NAND2_X1 U8863 ( .A1(n14609), .A2(n7634), .ZN(n13821) );
  AND2_X1 U8864 ( .A1(n13832), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U8865 ( .A1(n7622), .A2(n7625), .ZN(n7620) );
  NAND2_X1 U8866 ( .A1(n7638), .A2(n12447), .ZN(n13841) );
  NAND2_X1 U8867 ( .A1(n11450), .A2(n11449), .ZN(n14645) );
  NAND2_X1 U8868 ( .A1(n7189), .A2(n7192), .ZN(n13871) );
  NAND2_X1 U8869 ( .A1(n7191), .A2(n7190), .ZN(n7189) );
  INV_X1 U8870 ( .A(n12463), .ZN(n7191) );
  INV_X1 U8871 ( .A(n14325), .ZN(n13876) );
  OAI21_X1 U8872 ( .B1(n14610), .B2(n7185), .A(n7183), .ZN(n13880) );
  NAND2_X1 U8873 ( .A1(n14610), .A2(n14611), .ZN(n14609) );
  XOR2_X1 U8874 ( .A(n9352), .B(n9351), .Z(n9354) );
  OR2_X1 U8875 ( .A1(n8837), .A2(n8830), .ZN(n13932) );
  INV_X1 U8876 ( .A(n11692), .ZN(n6746) );
  OR2_X1 U8877 ( .A1(n11607), .A2(n8838), .ZN(n8839) );
  NAND2_X1 U8878 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6834) );
  NAND2_X1 U8879 ( .A1(n8722), .A2(n6579), .ZN(n8680) );
  NOR2_X1 U8880 ( .A1(n8695), .A2(n6827), .ZN(n8697) );
  AND2_X1 U8881 ( .A1(n9768), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8882 ( .A1(n8754), .A2(n6674), .ZN(n8755) );
  NAND2_X1 U8883 ( .A1(n8755), .A2(n8756), .ZN(n8769) );
  NAND2_X1 U8884 ( .A1(n8769), .A2(n6826), .ZN(n8770) );
  OR2_X1 U8885 ( .A1(n10025), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6826) );
  NOR2_X1 U8886 ( .A1(n9589), .A2(n9590), .ZN(n9694) );
  NAND2_X1 U8887 ( .A1(n13997), .A2(n6831), .ZN(n9589) );
  OR2_X1 U8888 ( .A1(n14006), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8889 ( .A1(n14722), .A2(n10490), .ZN(n10493) );
  AND2_X1 U8890 ( .A1(n10829), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14018) );
  AND2_X1 U8891 ( .A1(n6830), .A2(n6829), .ZN(n10829) );
  NAND2_X1 U8892 ( .A1(n10828), .A2(n10834), .ZN(n6829) );
  NAND2_X1 U8893 ( .A1(n11625), .A2(n11624), .ZN(n14039) );
  NAND2_X1 U8894 ( .A1(n7410), .A2(n7409), .ZN(n14059) );
  NAND2_X1 U8895 ( .A1(n14309), .A2(n11713), .ZN(n14124) );
  NAND2_X1 U8896 ( .A1(n14192), .A2(n11709), .ZN(n14176) );
  NAND2_X1 U8897 ( .A1(n7343), .A2(n11706), .ZN(n14216) );
  OR2_X1 U8898 ( .A1(n14234), .A2(n11705), .ZN(n7343) );
  INV_X1 U8899 ( .A(n14343), .ZN(n14240) );
  NAND2_X1 U8900 ( .A1(n7383), .A2(n7384), .ZN(n14626) );
  NAND2_X1 U8901 ( .A1(n6959), .A2(n10754), .ZN(n10756) );
  CLKBUF_X1 U8902 ( .A(n14656), .Z(n6959) );
  NAND2_X1 U8903 ( .A1(n7330), .A2(n10597), .ZN(n10751) );
  NAND2_X1 U8904 ( .A1(n14486), .A2(n14491), .ZN(n7330) );
  NAND2_X1 U8905 ( .A1(n7408), .A2(n7407), .ZN(n10344) );
  NAND2_X1 U8906 ( .A1(n7408), .A2(n10213), .ZN(n10220) );
  NAND2_X1 U8907 ( .A1(n7301), .A2(n10237), .ZN(n10359) );
  NAND2_X1 U8908 ( .A1(n10236), .A2(n10235), .ZN(n7301) );
  NAND2_X1 U8909 ( .A1(n7316), .A2(n7321), .ZN(n9765) );
  NAND2_X1 U8910 ( .A1(n6932), .A2(n7322), .ZN(n7316) );
  OAI21_X1 U8911 ( .B1(n6810), .B2(n6809), .A(n8808), .ZN(n6808) );
  NAND2_X1 U8912 ( .A1(n6807), .A2(n6806), .ZN(n10008) );
  NAND2_X1 U8913 ( .A1(n7492), .A2(n7324), .ZN(n6806) );
  INV_X1 U8914 ( .A(n6810), .ZN(n6807) );
  NAND2_X1 U8915 ( .A1(n7426), .A2(n9525), .ZN(n9748) );
  NAND2_X1 U8916 ( .A1(n9524), .A2(n11646), .ZN(n7426) );
  OR2_X1 U8917 ( .A1(n14747), .A2(n14624), .ZN(n14738) );
  OR2_X1 U8918 ( .A1(n14747), .A2(n14637), .ZN(n14247) );
  OR2_X1 U8919 ( .A1(n9217), .A2(n8835), .ZN(n14642) );
  INV_X1 U8920 ( .A(n14247), .ZN(n14262) );
  INV_X2 U8921 ( .A(n14806), .ZN(n14808) );
  OR2_X1 U8922 ( .A1(n14283), .A2(n14663), .ZN(n6960) );
  OR3_X1 U8923 ( .A1(n14329), .A2(n14328), .A3(n14327), .ZN(n14359) );
  AOI21_X1 U8924 ( .B1(n7310), .B2(P1_IR_REG_29__SCAN_IN), .A(n6634), .ZN(
        n7308) );
  OR2_X1 U8925 ( .A1(n8809), .A2(n7312), .ZN(n7307) );
  NAND2_X1 U8926 ( .A1(n7494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U8927 ( .A1(n7596), .A2(n7600), .ZN(n8250) );
  NAND2_X1 U8928 ( .A1(n7813), .A2(n7601), .ZN(n7596) );
  NAND2_X1 U8929 ( .A1(n7171), .A2(n7172), .ZN(n8183) );
  NAND2_X1 U8930 ( .A1(n8170), .A2(n6544), .ZN(n7172) );
  NAND2_X1 U8931 ( .A1(n7165), .A2(n7806), .ZN(n7171) );
  NAND2_X1 U8932 ( .A1(n8604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U8933 ( .A1(n8390), .A2(n7578), .ZN(n8602) );
  OR2_X1 U8934 ( .A1(n7604), .A2(n7605), .ZN(n8144) );
  INV_X1 U8935 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n15420) );
  INV_X1 U8936 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9476) );
  INV_X1 U8937 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9284) );
  INV_X1 U8938 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9417) );
  INV_X1 U8939 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9313) );
  INV_X1 U8940 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8633) );
  INV_X1 U8941 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8626) );
  INV_X1 U8942 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8598) );
  INV_X1 U8943 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8582) );
  INV_X1 U8944 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n15259) );
  INV_X1 U8945 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8551) );
  INV_X1 U8946 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8459) );
  INV_X1 U8947 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8452) );
  INV_X1 U8948 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U8949 ( .A1(n7491), .A2(n7490), .ZN(n8425) );
  NAND2_X1 U8950 ( .A1(n14437), .A2(n14436), .ZN(n14478) );
  NAND2_X1 U8951 ( .A1(n15449), .A2(n15450), .ZN(n14436) );
  AOI21_X1 U8952 ( .B1(n8967), .B2(n14440), .A(n15445), .ZN(n15439) );
  XNOR2_X1 U8953 ( .A(n14429), .B(n6924), .ZN(n15440) );
  XNOR2_X1 U8954 ( .A(n14443), .B(n14444), .ZN(n15438) );
  INV_X1 U8955 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7471) );
  XNOR2_X1 U8956 ( .A(n14450), .B(n7099), .ZN(n15443) );
  INV_X1 U8957 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7099) );
  XNOR2_X1 U8958 ( .A(n14452), .B(n14453), .ZN(n14482) );
  XNOR2_X1 U8959 ( .A(n14456), .B(n7466), .ZN(n14483) );
  INV_X1 U8960 ( .A(n14457), .ZN(n7466) );
  OAI21_X1 U8961 ( .B1(n7097), .B2(n6731), .A(n6619), .ZN(n14693) );
  NOR2_X1 U8962 ( .A1(n14688), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6731) );
  NOR2_X1 U8963 ( .A1(n14693), .A2(n14692), .ZN(n14691) );
  AND2_X1 U8964 ( .A1(n7103), .A2(n7100), .ZN(n14512) );
  AOI21_X1 U8965 ( .B1(n14702), .B2(n7104), .A(n6553), .ZN(n7103) );
  NAND2_X1 U8966 ( .A1(n14704), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7104) );
  INV_X1 U8967 ( .A(n7511), .ZN(n12749) );
  INV_X1 U8968 ( .A(n6764), .ZN(n12797) );
  OAI211_X1 U8969 ( .C1(n6767), .C2(n12791), .A(n6766), .B(n6765), .ZN(n6764)
         );
  OAI21_X1 U8970 ( .B1(n12380), .B2(n15140), .A(n7209), .ZN(P3_U3488) );
  INV_X1 U8971 ( .A(n7210), .ZN(n7209) );
  OAI21_X1 U8972 ( .B1(n12383), .B2(n13040), .A(n6629), .ZN(n7210) );
  NAND2_X1 U8973 ( .A1(n12807), .A2(n6599), .ZN(n6856) );
  INV_X1 U8974 ( .A(n6951), .ZN(n6950) );
  OAI21_X1 U8975 ( .B1(n13050), .B2(n13049), .A(n6952), .ZN(n6951) );
  INV_X1 U8976 ( .A(n6904), .ZN(n6903) );
  OAI21_X1 U8977 ( .B1(n13714), .B2(n13238), .A(n13132), .ZN(n6904) );
  INV_X1 U8978 ( .A(n6997), .ZN(n8997) );
  INV_X1 U8979 ( .A(n7001), .ZN(n7000) );
  NAND2_X1 U8980 ( .A1(n6999), .A2(n12044), .ZN(n6998) );
  NAND2_X1 U8981 ( .A1(n7003), .A2(n6527), .ZN(n7002) );
  OAI211_X1 U8982 ( .C1(n13618), .C2(n13561), .A(n8375), .B(n7700), .ZN(
        P2_U3236) );
  AOI21_X1 U8983 ( .B1(n13615), .B2(n14874), .A(n8374), .ZN(n8375) );
  OR2_X1 U8984 ( .A1(n14972), .A2(n7141), .ZN(n7140) );
  NAND2_X1 U8985 ( .A1(n13708), .A2(n14972), .ZN(n7142) );
  INV_X1 U8986 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U8987 ( .A1(n14961), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8988 ( .A1(n13708), .A2(n14962), .ZN(n6895) );
  AND2_X1 U8989 ( .A1(n6901), .A2(n13776), .ZN(n6900) );
  AOI21_X1 U8990 ( .B1(n6836), .B2(n14727), .A(n6835), .ZN(n14025) );
  NAND2_X1 U8991 ( .A1(n6913), .A2(n6912), .ZN(P1_U3526) );
  NAND2_X1 U8992 ( .A1(n14797), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8993 ( .A1(n6983), .A2(n6982), .ZN(P1_U3523) );
  NAND2_X1 U8994 ( .A1(n14797), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8995 ( .A1(n8809), .A2(n8810), .ZN(n11736) );
  INV_X1 U8996 ( .A(n7097), .ZN(n14689) );
  INV_X1 U8997 ( .A(n7105), .ZN(n14699) );
  INV_X1 U8998 ( .A(n7462), .ZN(n14697) );
  NOR2_X1 U8999 ( .A1(n14472), .A2(n14702), .ZN(n14705) );
  NOR2_X1 U9000 ( .A1(n14516), .A2(n14515), .ZN(n14474) );
  OAI21_X1 U9001 ( .B1(n14515), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7096), .ZN(
        n7095) );
  OR2_X1 U9002 ( .A1(n13050), .A2(n12575), .ZN(n6539) );
  AND2_X1 U9003 ( .A1(n6546), .A2(n12662), .ZN(n6540) );
  AND2_X1 U9004 ( .A1(n7642), .A2(n12483), .ZN(n6541) );
  INV_X2 U9005 ( .A(n12242), .ZN(n12228) );
  AND2_X1 U9006 ( .A1(n7192), .A2(n6541), .ZN(n6542) );
  INV_X1 U9007 ( .A(n11661), .ZN(n7329) );
  OR2_X1 U9008 ( .A1(n10930), .A2(n12969), .ZN(n6543) );
  INV_X1 U9009 ( .A(n14164), .ZN(n7398) );
  INV_X1 U9010 ( .A(n9991), .ZN(n7022) );
  AND2_X1 U9011 ( .A1(n7805), .A2(n7173), .ZN(n6544) );
  AOI21_X1 U9012 ( .B1(n12662), .B2(n7521), .A(n6600), .ZN(n7520) );
  INV_X1 U9013 ( .A(n7520), .ZN(n7519) );
  NAND2_X1 U9014 ( .A1(n13033), .A2(n12951), .ZN(n6545) );
  AND2_X1 U9015 ( .A1(n7044), .A2(n12603), .ZN(n6546) );
  OR2_X1 U9016 ( .A1(n12478), .A2(n13802), .ZN(n6547) );
  OR2_X1 U9017 ( .A1(n11641), .A2(n13938), .ZN(n11700) );
  INV_X1 U9018 ( .A(n14704), .ZN(n7102) );
  AND2_X1 U9019 ( .A1(n14373), .A2(n11516), .ZN(n14314) );
  INV_X1 U9020 ( .A(n14688), .ZN(n6732) );
  INV_X1 U9021 ( .A(n12201), .ZN(n7683) );
  NAND2_X1 U9022 ( .A1(n8146), .A2(n8145), .ZN(n13529) );
  AND2_X1 U9023 ( .A1(n7367), .A2(n11123), .ZN(n6548) );
  INV_X1 U9024 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8810) );
  AND2_X1 U9025 ( .A1(n7665), .A2(n7664), .ZN(n6549) );
  OR2_X1 U9026 ( .A1(n12095), .A2(n12094), .ZN(n6550) );
  INV_X1 U9027 ( .A(n12331), .ZN(n7480) );
  AND2_X1 U9028 ( .A1(n13150), .A2(n12330), .ZN(n12331) );
  AND2_X1 U9029 ( .A1(n13529), .A2(n13249), .ZN(n6551) );
  AND2_X1 U9030 ( .A1(n6574), .A2(n6701), .ZN(n6552) );
  NOR2_X1 U9031 ( .A1(n7387), .A2(n11694), .ZN(n7386) );
  INV_X1 U9032 ( .A(n12100), .ZN(n7685) );
  AND2_X1 U9033 ( .A1(n7102), .A2(n11091), .ZN(n6553) );
  OR2_X1 U9034 ( .A1(n12112), .A2(n6597), .ZN(n6554) );
  INV_X1 U9035 ( .A(n12197), .ZN(n7218) );
  AND2_X1 U9036 ( .A1(n7587), .A2(n9915), .ZN(n6555) );
  AND2_X1 U9037 ( .A1(n6991), .A2(n12382), .ZN(n6556) );
  OR2_X1 U9038 ( .A1(n15127), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U9039 ( .A1(n12024), .A2(n9892), .ZN(n15068) );
  INV_X1 U9040 ( .A(n15068), .ZN(n15053) );
  AND2_X1 U9041 ( .A1(n9515), .A2(n9514), .ZN(n11385) );
  INV_X1 U9042 ( .A(n11385), .ZN(n7324) );
  INV_X1 U9043 ( .A(n9019), .ZN(n12545) );
  OAI211_X2 U9044 ( .C1(n8899), .C2(n8906), .A(n7851), .B(n7850), .ZN(n7852)
         );
  NOR2_X1 U9045 ( .A1(n10382), .A2(n7476), .ZN(n6558) );
  AND2_X1 U9046 ( .A1(n11841), .A2(n11842), .ZN(n11984) );
  INV_X1 U9047 ( .A(n7130), .ZN(n12043) );
  AND2_X1 U9048 ( .A1(n13672), .A2(n13250), .ZN(n6559) );
  INV_X1 U9049 ( .A(n11694), .ZN(n10755) );
  NAND2_X1 U9050 ( .A1(n11445), .A2(n11693), .ZN(n11694) );
  NOR2_X1 U9051 ( .A1(n10397), .A2(n10391), .ZN(n6560) );
  INV_X1 U9052 ( .A(n9097), .ZN(n7513) );
  INV_X1 U9053 ( .A(n14088), .ZN(n7419) );
  INV_X1 U9054 ( .A(n8875), .ZN(n7441) );
  NAND2_X1 U9055 ( .A1(n7677), .A2(n7678), .ZN(n7964) );
  AND2_X1 U9056 ( .A1(n12331), .A2(n13228), .ZN(n6561) );
  NAND2_X1 U9057 ( .A1(n7621), .A2(n13862), .ZN(n13831) );
  OR2_X1 U9058 ( .A1(n8500), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n6562) );
  AND3_X1 U9059 ( .A1(n9281), .A2(n8382), .A3(n8381), .ZN(n6563) );
  OR2_X2 U9060 ( .A1(n14145), .A2(n14144), .ZN(n14309) );
  AND2_X1 U9061 ( .A1(n11385), .A2(n7323), .ZN(n6564) );
  AND2_X1 U9062 ( .A1(n7454), .A2(n8344), .ZN(n6565) );
  NOR2_X1 U9063 ( .A1(n11815), .A2(n6876), .ZN(n6566) );
  AND2_X1 U9064 ( .A1(n12398), .A2(n12394), .ZN(n6567) );
  NAND2_X1 U9065 ( .A1(n15015), .A2(n10928), .ZN(n6568) );
  AND2_X1 U9066 ( .A1(n7086), .A2(n8463), .ZN(n6569) );
  AND2_X1 U9067 ( .A1(n12211), .A2(n12210), .ZN(n6570) );
  AND2_X1 U9068 ( .A1(n9727), .A2(n9726), .ZN(n6571) );
  OR2_X1 U9069 ( .A1(n14467), .A2(n14466), .ZN(n6572) );
  OR2_X1 U9070 ( .A1(n14380), .A2(n14381), .ZN(n6573) );
  AND2_X1 U9071 ( .A1(n11158), .A2(n7248), .ZN(n6574) );
  INV_X1 U9072 ( .A(n6719), .ZN(n7381) );
  NAND2_X1 U9073 ( .A1(n7384), .A2(n7382), .ZN(n6719) );
  OR2_X1 U9074 ( .A1(n12189), .A2(n12188), .ZN(n6575) );
  AND3_X1 U9075 ( .A1(n7843), .A2(n7842), .A3(n7840), .ZN(n6576) );
  XNOR2_X1 U9076 ( .A(n6834), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13960) );
  INV_X1 U9077 ( .A(n13960), .ZN(n6931) );
  OR2_X1 U9078 ( .A1(n14107), .A2(n13935), .ZN(n6577) );
  NAND2_X1 U9079 ( .A1(n11602), .A2(n11601), .ZN(n14280) );
  INV_X1 U9080 ( .A(n14280), .ZN(n6822) );
  NAND2_X1 U9081 ( .A1(n7722), .A2(n7718), .ZN(n7855) );
  XNOR2_X1 U9082 ( .A(n14519), .B(n14416), .ZN(n6578) );
  OR2_X1 U9083 ( .A1(n9742), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6579) );
  AND2_X1 U9084 ( .A1(n8408), .A2(n8409), .ZN(n6580) );
  INV_X1 U9085 ( .A(n7677), .ZN(n7846) );
  AND2_X1 U9086 ( .A1(n7420), .A2(n6577), .ZN(n6581) );
  AND2_X1 U9087 ( .A1(n6899), .A2(n7338), .ZN(n6582) );
  AND2_X1 U9088 ( .A1(n9069), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6583) );
  INV_X1 U9089 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U9090 ( .A1(n8022), .A2(n8021), .ZN(n14819) );
  XNOR2_X1 U9091 ( .A(n14284), .B(n14042), .ZN(n14056) );
  INV_X1 U9092 ( .A(n14056), .ZN(n7416) );
  INV_X1 U9093 ( .A(n12958), .ZN(n6848) );
  INV_X1 U9094 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13748) );
  XNOR2_X1 U9095 ( .A(n12381), .B(n12676), .ZN(n12009) );
  INV_X1 U9096 ( .A(n13440), .ZN(n13718) );
  NAND2_X1 U9097 ( .A1(n11528), .A2(n11527), .ZN(n14307) );
  INV_X1 U9098 ( .A(n14307), .ZN(n7499) );
  AND2_X1 U9099 ( .A1(n8716), .A2(n13118), .ZN(n9678) );
  OR2_X1 U9100 ( .A1(n14080), .A2(n14280), .ZN(n6584) );
  XNOR2_X1 U9101 ( .A(n14523), .B(n14522), .ZN(n6585) );
  OR2_X1 U9102 ( .A1(n14453), .A2(n14452), .ZN(n6586) );
  AND2_X1 U9103 ( .A1(n6995), .A2(n6994), .ZN(n6587) );
  INV_X1 U9104 ( .A(n11406), .ZN(n7569) );
  OR2_X1 U9105 ( .A1(n14169), .A2(n6823), .ZN(n6588) );
  NAND2_X1 U9106 ( .A1(n8416), .A2(n8414), .ZN(n6589) );
  INV_X1 U9107 ( .A(n11386), .ZN(n7323) );
  OR2_X1 U9108 ( .A1(n9987), .A2(n9291), .ZN(n6590) );
  INV_X1 U9109 ( .A(n11411), .ZN(n7565) );
  AND2_X1 U9110 ( .A1(n14075), .A2(n7337), .ZN(n6591) );
  AND2_X1 U9111 ( .A1(n12251), .A2(n12250), .ZN(n6592) );
  OR2_X1 U9112 ( .A1(n14581), .A2(n10865), .ZN(n6593) );
  AND3_X1 U9113 ( .A1(n9488), .A2(n9487), .A3(n9486), .ZN(n9903) );
  OR2_X1 U9114 ( .A1(n7751), .A2(n7750), .ZN(n6594) );
  OR2_X1 U9115 ( .A1(n10263), .A2(n9606), .ZN(n6595) );
  OR2_X1 U9116 ( .A1(n7513), .A2(n9089), .ZN(n6596) );
  AND2_X1 U9117 ( .A1(n12109), .A2(n12108), .ZN(n6597) );
  AND2_X1 U9118 ( .A1(n13643), .A2(n13245), .ZN(n6598) );
  AND2_X1 U9119 ( .A1(n6862), .A2(n6557), .ZN(n6599) );
  AND2_X1 U9120 ( .A1(n11785), .A2(n11784), .ZN(n6600) );
  INV_X1 U9121 ( .A(n11638), .ZN(n7561) );
  AND2_X1 U9122 ( .A1(n7441), .A2(n6536), .ZN(n6601) );
  AND2_X1 U9123 ( .A1(n7296), .A2(n12292), .ZN(n6602) );
  AND2_X1 U9124 ( .A1(n10908), .A2(n11878), .ZN(n6603) );
  INV_X1 U9125 ( .A(n7374), .ZN(n13408) );
  INV_X1 U9126 ( .A(n6909), .ZN(n13484) );
  NOR2_X1 U9127 ( .A1(n13499), .A2(n13648), .ZN(n6909) );
  OR2_X1 U9128 ( .A1(n7390), .A2(n7389), .ZN(n6604) );
  INV_X1 U9129 ( .A(n12174), .ZN(n6962) );
  AND2_X1 U9130 ( .A1(n6970), .A2(n6743), .ZN(n6605) );
  INV_X1 U9131 ( .A(n11425), .ZN(n7548) );
  NAND2_X1 U9132 ( .A1(n12755), .A2(n12748), .ZN(n6606) );
  INV_X1 U9133 ( .A(n7193), .ZN(n7190) );
  NAND2_X1 U9134 ( .A1(n6547), .A2(n12464), .ZN(n7193) );
  AND2_X1 U9135 ( .A1(n11767), .A2(n11766), .ZN(n6607) );
  AND2_X1 U9136 ( .A1(n7532), .A2(n10866), .ZN(n6608) );
  NAND3_X1 U9137 ( .A1(n15181), .A2(n8523), .A3(n8438), .ZN(n6609) );
  OR2_X1 U9138 ( .A1(n7480), .A2(n7128), .ZN(n6610) );
  OR2_X1 U9139 ( .A1(n7218), .A2(n12198), .ZN(n6611) );
  AND2_X1 U9140 ( .A1(n13073), .A2(n12909), .ZN(n6612) );
  NAND2_X1 U9141 ( .A1(n7511), .A2(n6606), .ZN(n7510) );
  NAND2_X1 U9142 ( .A1(n8069), .A2(n8068), .ZN(n13743) );
  AND2_X1 U9143 ( .A1(n10543), .A2(n10542), .ZN(n6613) );
  INV_X1 U9144 ( .A(n12261), .ZN(n13418) );
  NAND2_X1 U9145 ( .A1(n12479), .A2(n7194), .ZN(n6614) );
  AND2_X1 U9146 ( .A1(n12299), .A2(n13418), .ZN(n6615) );
  OR2_X1 U9147 ( .A1(n14444), .A2(n14443), .ZN(n6616) );
  NAND2_X1 U9148 ( .A1(n7393), .A2(n7390), .ZN(n6617) );
  NOR2_X1 U9149 ( .A1(n14666), .A2(n13944), .ZN(n6618) );
  OR2_X1 U9150 ( .A1(n6732), .A2(n9845), .ZN(n6619) );
  NOR2_X1 U9151 ( .A1(n14790), .A2(n13947), .ZN(n6620) );
  NOR2_X1 U9152 ( .A1(n14337), .A2(n13940), .ZN(n6621) );
  NOR2_X1 U9153 ( .A1(n12103), .A2(n8324), .ZN(n6622) );
  NOR2_X1 U9154 ( .A1(n13206), .A2(n12333), .ZN(n6623) );
  INV_X1 U9155 ( .A(n6850), .ZN(n6849) );
  NAND2_X1 U9156 ( .A1(n6545), .A2(n11280), .ZN(n6850) );
  AND2_X1 U9157 ( .A1(n12571), .A2(n12662), .ZN(n6624) );
  OAI21_X1 U9158 ( .B1(n7534), .B2(n7535), .A(n6593), .ZN(n7533) );
  AND2_X1 U9159 ( .A1(n12115), .A2(n13258), .ZN(n6625) );
  AND2_X1 U9160 ( .A1(n11990), .A2(n6704), .ZN(n6626) );
  INV_X1 U9161 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n15338) );
  INV_X1 U9162 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U9163 ( .A1(n7398), .A2(n14181), .ZN(n7397) );
  AND2_X1 U9164 ( .A1(n7570), .A2(n7569), .ZN(n6627) );
  NAND2_X1 U9165 ( .A1(n8858), .A2(n7047), .ZN(n6628) );
  AND2_X1 U9166 ( .A1(n11300), .A2(n7211), .ZN(n6629) );
  NOR2_X1 U9167 ( .A1(n11755), .A2(n12961), .ZN(n6630) );
  NOR2_X1 U9168 ( .A1(n14280), .A2(n14062), .ZN(n6631) );
  OR2_X1 U9169 ( .A1(n11278), .A2(n12575), .ZN(n11291) );
  OR2_X1 U9170 ( .A1(n13264), .A2(n13184), .ZN(n6632) );
  INV_X1 U9171 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8456) );
  INV_X1 U9172 ( .A(n7286), .ZN(n7285) );
  NAND2_X1 U9173 ( .A1(n12283), .A2(n8064), .ZN(n7286) );
  INV_X1 U9174 ( .A(n8469), .ZN(n7348) );
  INV_X1 U9175 ( .A(n7594), .ZN(n7593) );
  OAI21_X1 U9176 ( .B1(n7595), .B2(n8015), .A(n7780), .ZN(n7594) );
  NAND2_X1 U9177 ( .A1(n7796), .A2(n7795), .ZN(n6633) );
  AND2_X1 U9178 ( .A1(n7313), .A2(n7309), .ZN(n6634) );
  OR2_X1 U9179 ( .A1(n7425), .A2(n9747), .ZN(n6635) );
  AND2_X1 U9180 ( .A1(n13440), .A2(n7139), .ZN(n6636) );
  AND2_X1 U9181 ( .A1(n6558), .A2(n7475), .ZN(n6637) );
  NOR2_X1 U9182 ( .A1(n12423), .A2(n12424), .ZN(n6638) );
  INV_X1 U9183 ( .A(n6820), .ZN(n14045) );
  NOR2_X1 U9184 ( .A1(n14080), .A2(n6821), .ZN(n6820) );
  AND2_X1 U9185 ( .A1(n14284), .A2(n14042), .ZN(n6639) );
  NAND2_X1 U9186 ( .A1(n13512), .A2(n8347), .ZN(n6640) );
  AND2_X1 U9187 ( .A1(n7485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6641) );
  OR2_X1 U9188 ( .A1(n8045), .A2(SI_14_), .ZN(n6642) );
  INV_X1 U9189 ( .A(n12202), .ZN(n7682) );
  NAND2_X1 U9190 ( .A1(n7488), .A2(n7487), .ZN(n6643) );
  INV_X1 U9191 ( .A(n7634), .ZN(n7185) );
  AND2_X1 U9192 ( .A1(n13822), .A2(n13820), .ZN(n7634) );
  AND2_X1 U9193 ( .A1(n13060), .A2(n12838), .ZN(n6644) );
  INV_X1 U9194 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U9195 ( .A1(n7661), .A2(n7660), .ZN(n7659) );
  NAND2_X1 U9196 ( .A1(n11291), .A2(n11290), .ZN(n12812) );
  OR2_X1 U9197 ( .A1(n6822), .A2(n14058), .ZN(n6645) );
  INV_X1 U9198 ( .A(n11563), .ZN(n7544) );
  INV_X1 U9199 ( .A(n11415), .ZN(n7563) );
  OR2_X1 U9200 ( .A1(n13073), .A2(n12909), .ZN(n6646) );
  OR2_X1 U9201 ( .A1(n11029), .A2(n10974), .ZN(n11900) );
  OR2_X1 U9202 ( .A1(n12940), .A2(n12952), .ZN(n11923) );
  INV_X1 U9203 ( .A(n11923), .ZN(n7263) );
  INV_X1 U9204 ( .A(n12275), .ZN(n10463) );
  OR2_X1 U9205 ( .A1(n13529), .A2(n13249), .ZN(n6647) );
  OR2_X1 U9206 ( .A1(n10868), .A2(n9251), .ZN(n6648) );
  OR2_X1 U9207 ( .A1(n14460), .A2(n14459), .ZN(n6649) );
  OR2_X1 U9208 ( .A1(n14382), .A2(n14383), .ZN(n6650) );
  AND2_X1 U9209 ( .A1(n6882), .A2(n6880), .ZN(n6652) );
  INV_X1 U9210 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7014) );
  INV_X1 U9211 ( .A(n13771), .ZN(n7633) );
  AOI21_X1 U9212 ( .B1(n12549), .B2(n12548), .A(n12550), .ZN(n13771) );
  AND2_X1 U9213 ( .A1(n6990), .A2(n12378), .ZN(n6653) );
  NOR2_X1 U9214 ( .A1(n14705), .A2(n14704), .ZN(n6654) );
  AND2_X1 U9215 ( .A1(n11851), .A2(n11857), .ZN(n11989) );
  INV_X1 U9216 ( .A(n11989), .ZN(n7206) );
  AND2_X1 U9217 ( .A1(n7817), .A2(n7815), .ZN(n6655) );
  AND2_X1 U9218 ( .A1(n12928), .A2(n11825), .ZN(n12946) );
  OR2_X1 U9219 ( .A1(n12667), .A2(n11784), .ZN(n6656) );
  AND2_X1 U9220 ( .A1(n12097), .A2(n12096), .ZN(n6657) );
  AND2_X1 U9221 ( .A1(n11694), .A2(n10754), .ZN(n6658) );
  AND2_X1 U9222 ( .A1(n10690), .A2(n10919), .ZN(n6659) );
  INV_X1 U9223 ( .A(n11284), .ZN(n6876) );
  AND2_X1 U9224 ( .A1(n11446), .A2(n7581), .ZN(n6660) );
  AND2_X1 U9225 ( .A1(n6655), .A2(n7715), .ZN(n6661) );
  AND2_X1 U9226 ( .A1(n7578), .A2(n7577), .ZN(n6662) );
  INV_X1 U9227 ( .A(n7699), .ZN(n7612) );
  AND2_X1 U9228 ( .A1(n7680), .A2(n6611), .ZN(n6663) );
  NOR2_X1 U9229 ( .A1(n7528), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6664) );
  INV_X1 U9230 ( .A(n11590), .ZN(n7576) );
  NAND2_X1 U9231 ( .A1(n7684), .A2(n7685), .ZN(n6665) );
  INV_X1 U9232 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n15368) );
  INV_X1 U9233 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8613) );
  AND2_X1 U9234 ( .A1(n6842), .A2(n11282), .ZN(n6666) );
  OR2_X1 U9235 ( .A1(n13512), .A2(n13248), .ZN(n6667) );
  AND2_X1 U9236 ( .A1(n6857), .A2(n6856), .ZN(n6668) );
  INV_X1 U9237 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8801) );
  INV_X1 U9238 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7486) );
  INV_X1 U9239 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7309) );
  OR2_X1 U9240 ( .A1(n7560), .A2(n11638), .ZN(n6669) );
  NAND2_X1 U9241 ( .A1(n7474), .A2(n12337), .ZN(n6670) );
  OR2_X1 U9242 ( .A1(n7633), .A2(n7631), .ZN(n6671) );
  AND2_X1 U9243 ( .A1(n8612), .A2(n8613), .ZN(n6672) );
  INV_X1 U9244 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8553) );
  CLKBUF_X3 U9245 ( .A(n9484), .Z(n11274) );
  INV_X1 U9246 ( .A(n13243), .ZN(n7139) );
  INV_X1 U9247 ( .A(n14996), .ZN(n6707) );
  NAND2_X1 U9248 ( .A1(n10739), .A2(n10738), .ZN(n13930) );
  INV_X1 U9249 ( .A(n13930), .ZN(n7497) );
  AND2_X1 U9250 ( .A1(n10818), .A2(n7367), .ZN(n6673) );
  INV_X1 U9251 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U9252 ( .A1(n7583), .A2(n12217), .ZN(n13386) );
  INV_X1 U9253 ( .A(n13386), .ZN(n7372) );
  OR2_X1 U9254 ( .A1(n10019), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6674) );
  INV_X1 U9255 ( .A(n11622), .ZN(n11496) );
  INV_X1 U9256 ( .A(n13861), .ZN(n7624) );
  AND2_X1 U9257 ( .A1(n12837), .A2(n15062), .ZN(n6675) );
  NOR2_X1 U9258 ( .A1(n13192), .A2(n12345), .ZN(n6676) );
  NOR2_X1 U9259 ( .A1(n14235), .A2(n14337), .ZN(n6813) );
  INV_X1 U9260 ( .A(n7371), .ZN(n13511) );
  OR2_X1 U9261 ( .A1(n10540), .A2(n9965), .ZN(n6677) );
  AND2_X1 U9262 ( .A1(n13743), .A2(n13253), .ZN(n6678) );
  AND2_X1 U9263 ( .A1(n7383), .A2(n7381), .ZN(n6679) );
  AND2_X1 U9264 ( .A1(n7097), .A2(n6732), .ZN(n6680) );
  OR2_X1 U9265 ( .A1(n14169), .A2(n14314), .ZN(n6681) );
  NAND2_X1 U9266 ( .A1(n12429), .A2(n12430), .ZN(n6682) );
  OR2_X1 U9267 ( .A1(n13710), .A2(n13668), .ZN(n6683) );
  OR2_X1 U9268 ( .A1(n13710), .A2(n13730), .ZN(n6684) );
  AND2_X1 U9269 ( .A1(n12327), .A2(n12326), .ZN(n6685) );
  OR2_X1 U9270 ( .A1(n9244), .A2(n9243), .ZN(n14797) );
  AND2_X1 U9271 ( .A1(n9411), .A2(n9410), .ZN(n15125) );
  INV_X1 U9272 ( .A(n13735), .ZN(n6910) );
  NAND2_X1 U9273 ( .A1(n8263), .A2(n7712), .ZN(n8267) );
  AND2_X1 U9274 ( .A1(n7364), .A2(n10186), .ZN(n6686) );
  OR2_X1 U9275 ( .A1(n7810), .A2(SI_25_), .ZN(n6687) );
  NAND2_X1 U9276 ( .A1(n8173), .A2(n8172), .ZN(n13653) );
  INV_X1 U9277 ( .A(n13653), .ZN(n7370) );
  INV_X1 U9278 ( .A(n10654), .ZN(n10962) );
  AND2_X1 U9279 ( .A1(n9665), .A2(n7523), .ZN(n6688) );
  NOR2_X1 U9280 ( .A1(n8232), .A2(SI_27_), .ZN(n6689) );
  INV_X1 U9281 ( .A(n7496), .ZN(n10057) );
  NOR2_X1 U9282 ( .A1(n9948), .A2(n11403), .ZN(n7496) );
  INV_X1 U9283 ( .A(n7602), .ZN(n7601) );
  OR2_X1 U9284 ( .A1(n8233), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U9285 ( .A1(n7526), .A2(n7525), .ZN(n7524) );
  INV_X1 U9286 ( .A(n10370), .ZN(n7077) );
  AND2_X1 U9287 ( .A1(n10499), .A2(n7613), .ZN(n6690) );
  INV_X1 U9288 ( .A(n12084), .ZN(n7365) );
  INV_X1 U9289 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7713) );
  AND2_X2 U9290 ( .A1(n9560), .A2(n9559), .ZN(n15142) );
  NAND2_X1 U9291 ( .A1(n9336), .A2(n9325), .ZN(n14813) );
  INV_X1 U9292 ( .A(n14813), .ZN(n13227) );
  INV_X1 U9293 ( .A(n14758), .ZN(n6809) );
  NAND2_X1 U9294 ( .A1(n10021), .A2(n10020), .ZN(n11409) );
  INV_X1 U9295 ( .A(n11409), .ZN(n7495) );
  AND2_X2 U9296 ( .A1(n10078), .A2(n10077), .ZN(n14962) );
  XNOR2_X1 U9297 ( .A(n7816), .B(n7815), .ZN(n8360) );
  NAND2_X1 U9298 ( .A1(n10218), .A2(n10217), .ZN(n14790) );
  INV_X1 U9299 ( .A(n14790), .ZN(n6824) );
  AND2_X1 U9300 ( .A1(n12782), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U9301 ( .A1(n7508), .A2(n6590), .ZN(n7058) );
  AND2_X1 U9302 ( .A1(n12765), .A2(n14529), .ZN(n6692) );
  OR2_X1 U9303 ( .A1(n12307), .A2(n12306), .ZN(n6693) );
  INV_X1 U9304 ( .A(n7492), .ZN(n9516) );
  INV_X1 U9305 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7197) );
  INV_X1 U9306 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7013) );
  INV_X1 U9307 ( .A(n8306), .ZN(n12044) );
  INV_X1 U9308 ( .A(n9915), .ZN(n12301) );
  NAND2_X1 U9309 ( .A1(n8301), .A2(n8302), .ZN(n9915) );
  AND2_X1 U9310 ( .A1(n9438), .A2(n9294), .ZN(n6694) );
  OR2_X1 U9311 ( .A1(n9430), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6695) );
  INV_X1 U9312 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7313) );
  INV_X1 U9313 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7267) );
  INV_X1 U9314 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U9315 ( .A1(n14349), .A2(n6528), .ZN(n6913) );
  NAND2_X2 U9316 ( .A1(n6696), .A2(n13162), .ZN(n12360) );
  NAND2_X1 U9317 ( .A1(n12311), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U9318 ( .A1(n11116), .A2(n11115), .ZN(n12315) );
  NOR2_X2 U9319 ( .A1(n12391), .A2(n11114), .ZN(n11116) );
  AND4_X2 U9320 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7891), .ZN(n7678)
         );
  AOI21_X1 U9321 ( .B1(n13183), .B2(n9725), .A(n13182), .ZN(n13172) );
  NAND2_X1 U9322 ( .A1(n9861), .A2(n6697), .ZN(n10376) );
  NAND3_X1 U9323 ( .A1(n9855), .A2(n9854), .A3(n9857), .ZN(n6697) );
  XNOR2_X1 U9324 ( .A(n12356), .B(n9565), .ZN(n9576) );
  NAND3_X1 U9325 ( .A1(n7530), .A2(n6710), .A3(n8543), .ZN(n9049) );
  XNOR2_X2 U9326 ( .A(n6709), .B(n9050), .ZN(n11302) );
  INV_X1 U9327 ( .A(SI_14_), .ZN(n6716) );
  AND2_X1 U9328 ( .A1(n6721), .A2(n6594), .ZN(n7931) );
  NAND3_X1 U9329 ( .A1(n6721), .A2(n6594), .A3(n7753), .ZN(n6722) );
  OAI21_X1 U9330 ( .B1(n7849), .B2(n7848), .A(n7734), .ZN(n6725) );
  NAND3_X1 U9331 ( .A1(n6724), .A2(n7864), .A3(n6723), .ZN(n7737) );
  NAND2_X1 U9332 ( .A1(n7849), .A2(n7734), .ZN(n6724) );
  XNOR2_X1 U9333 ( .A(n6725), .B(n7864), .ZN(n9348) );
  NAND2_X1 U9334 ( .A1(n11400), .A2(n7570), .ZN(n7567) );
  NAND2_X1 U9335 ( .A1(n6729), .A2(n11391), .ZN(n6728) );
  NAND2_X1 U9336 ( .A1(n11390), .A2(n11392), .ZN(n6729) );
  INV_X1 U9337 ( .A(n7199), .ZN(n8606) );
  NAND2_X1 U9338 ( .A1(n14693), .A2(n14692), .ZN(n14463) );
  NAND3_X1 U9339 ( .A1(n7545), .A2(n6737), .A3(n6736), .ZN(n11444) );
  INV_X1 U9340 ( .A(n7547), .ZN(n6741) );
  NAND2_X1 U9341 ( .A1(n6745), .A2(n11691), .ZN(P1_U3242) );
  NAND2_X1 U9342 ( .A1(n6747), .A2(n6746), .ZN(n6745) );
  NAND2_X1 U9343 ( .A1(n6750), .A2(n6748), .ZN(n6747) );
  NAND2_X1 U9344 ( .A1(n6749), .A2(n11337), .ZN(n6748) );
  NAND2_X1 U9345 ( .A1(n7559), .A2(n7554), .ZN(n6749) );
  AOI21_X1 U9346 ( .B1(n7559), .B2(n7555), .A(n11685), .ZN(n6750) );
  NAND2_X1 U9347 ( .A1(n11616), .A2(n11617), .ZN(n11621) );
  INV_X1 U9348 ( .A(n7467), .ZN(n14380) );
  XNOR2_X1 U9349 ( .A(n7467), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14439) );
  MUX2_X1 U9350 ( .A(n14543), .B(n9272), .S(n15181), .Z(n9273) );
  NAND2_X1 U9351 ( .A1(n14528), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U9352 ( .A1(n12050), .A2(n12049), .ZN(n6769) );
  NAND2_X1 U9353 ( .A1(n12189), .A2(n12188), .ZN(n6937) );
  NAND2_X1 U9354 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  INV_X1 U9355 ( .A(n12184), .ZN(n6771) );
  INV_X1 U9356 ( .A(n6776), .ZN(n6772) );
  NAND2_X1 U9357 ( .A1(n6775), .A2(n6774), .ZN(n6773) );
  NAND2_X1 U9358 ( .A1(n6776), .A2(n12184), .ZN(n6775) );
  NAND2_X1 U9359 ( .A1(n7671), .A2(n7670), .ZN(n6776) );
  AND3_X1 U9360 ( .A1(n6785), .A2(n6786), .A3(n6784), .ZN(n12081) );
  NAND2_X1 U9361 ( .A1(n6788), .A2(n6787), .ZN(n6785) );
  AND3_X2 U9362 ( .A1(n7677), .A2(n7709), .A3(n6651), .ZN(n7244) );
  INV_X2 U9363 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8090) );
  AND3_X2 U9364 ( .A1(n6791), .A2(n6790), .A3(n6789), .ZN(n7677) );
  OAI21_X1 U9365 ( .B1(n12107), .B2(n12106), .A(n6554), .ZN(n6920) );
  NAND2_X1 U9366 ( .A1(n6792), .A2(n7227), .ZN(n12107) );
  NAND3_X1 U9367 ( .A1(n6793), .A2(n6550), .A3(n6665), .ZN(n6792) );
  INV_X1 U9368 ( .A(n12093), .ZN(n6793) );
  NAND2_X1 U9369 ( .A1(n8263), .A2(n7298), .ZN(n6794) );
  NAND2_X1 U9370 ( .A1(n6797), .A2(n6693), .ZN(P2_U3328) );
  NAND2_X1 U9371 ( .A1(n6799), .A2(n6798), .ZN(n6797) );
  NAND3_X1 U9372 ( .A1(n6802), .A2(n6801), .A3(n6800), .ZN(n6799) );
  OR2_X1 U9373 ( .A1(n12303), .A2(n6986), .ZN(n6800) );
  NAND2_X1 U9374 ( .A1(n12303), .A2(n12259), .ZN(n6801) );
  NAND2_X1 U9375 ( .A1(n6803), .A2(n6555), .ZN(n6802) );
  NAND2_X1 U9376 ( .A1(n12303), .A2(n12302), .ZN(n6803) );
  NOR2_X1 U9377 ( .A1(n14758), .A2(n7324), .ZN(n6805) );
  NOR2_X1 U9378 ( .A1(n6808), .A2(n9787), .ZN(n14757) );
  NAND2_X2 U9379 ( .A1(n11748), .A2(n14708), .ZN(n11516) );
  XNOR2_X2 U9380 ( .A(n6812), .B(n8613), .ZN(n11748) );
  INV_X1 U9381 ( .A(n6813), .ZN(n14226) );
  INV_X2 U9382 ( .A(n14737), .ZN(n11380) );
  NAND3_X1 U9383 ( .A1(n11374), .A2(n6814), .A3(n14737), .ZN(n7492) );
  NAND2_X2 U9384 ( .A1(n6816), .A2(n6817), .ZN(n11372) );
  AOI22_X1 U9385 ( .A1(n11455), .A2(n13988), .B1(n11613), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6815) );
  AOI22_X2 U9386 ( .A1(n11455), .A2(n13972), .B1(n11613), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U9387 ( .A1(n11622), .A2(n6818), .ZN(n6817) );
  AND2_X1 U9388 ( .A1(n8877), .A2(n8878), .ZN(n6819) );
  NOR3_X2 U9389 ( .A1(n14169), .A2(n14301), .A3(n6823), .ZN(n14128) );
  NOR2_X2 U9390 ( .A1(n10360), .A2(n14672), .ZN(n14488) );
  NAND2_X1 U9391 ( .A1(n11039), .A2(n11903), .ZN(n6837) );
  NAND2_X1 U9392 ( .A1(n11028), .A2(n11896), .ZN(n6838) );
  NAND2_X1 U9393 ( .A1(n9906), .A2(n10128), .ZN(n10109) );
  NAND2_X1 U9394 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  NAND2_X1 U9395 ( .A1(n9889), .A2(n6839), .ZN(n9905) );
  NAND3_X1 U9396 ( .A1(n7530), .A2(n7215), .A3(n8543), .ZN(n6840) );
  NAND2_X1 U9397 ( .A1(n6840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9398 ( .A1(n11281), .A2(n6844), .ZN(n6841) );
  NAND2_X1 U9399 ( .A1(n6666), .A2(n6841), .ZN(n12931) );
  NAND2_X1 U9400 ( .A1(n11284), .A2(n6867), .ZN(n6866) );
  INV_X1 U9401 ( .A(n12919), .ZN(n6867) );
  NAND2_X1 U9402 ( .A1(n11286), .A2(n11285), .ZN(n12869) );
  INV_X1 U9403 ( .A(n6885), .ZN(n12836) );
  NAND2_X1 U9404 ( .A1(n12974), .A2(n10931), .ZN(n14562) );
  NAND2_X1 U9405 ( .A1(n10451), .A2(n10427), .ZN(n10916) );
  NAND2_X1 U9406 ( .A1(n7207), .A2(n7206), .ZN(n10203) );
  OAI21_X1 U9407 ( .B1(n12836), .B2(n11289), .A(n6656), .ZN(n12825) );
  NOR2_X1 U9408 ( .A1(n12824), .A2(n7696), .ZN(n12808) );
  NAND2_X1 U9409 ( .A1(n10453), .A2(n10452), .ZN(n10451) );
  OAI21_X2 U9410 ( .B1(n8063), .B2(n7286), .A(n7284), .ZN(n13566) );
  NAND2_X1 U9411 ( .A1(n6966), .A2(n6632), .ZN(n7272) );
  OAI21_X1 U9412 ( .B1(n10299), .B2(n7276), .A(n7274), .ZN(n7959) );
  AOI21_X1 U9413 ( .B1(n7291), .B2(n7290), .A(n7289), .ZN(n13419) );
  NAND2_X1 U9414 ( .A1(n7143), .A2(n13618), .ZN(n13708) );
  NAND2_X1 U9415 ( .A1(n6895), .A2(n6894), .ZN(P2_U3496) );
  INV_X1 U9416 ( .A(n6889), .ZN(n12263) );
  NAND2_X1 U9417 ( .A1(n6887), .A2(n6886), .ZN(n10161) );
  NAND2_X1 U9418 ( .A1(n7835), .A2(n8311), .ZN(n6889) );
  NAND2_X1 U9419 ( .A1(n7229), .A2(n7233), .ZN(n12303) );
  OAI22_X2 U9420 ( .A1(n7688), .A2(n12082), .B1(n12083), .B2(n7689), .ZN(
        n12095) );
  OAI22_X1 U9421 ( .A1(n12067), .A2(n7669), .B1(n12068), .B2(n7668), .ZN(
        n12075) );
  NAND2_X1 U9422 ( .A1(n7663), .A2(n7652), .ZN(n7651) );
  NAND3_X1 U9423 ( .A1(n7646), .A2(n7644), .A3(n6890), .ZN(n12042) );
  NAND3_X1 U9424 ( .A1(n12171), .A2(n6918), .A3(n12170), .ZN(n12176) );
  NAND3_X1 U9425 ( .A1(n7224), .A2(n7226), .A3(n7223), .ZN(n7225) );
  OR3_X1 U9426 ( .A1(n12209), .A2(n12208), .A3(n7230), .ZN(n7229) );
  NAND3_X1 U9427 ( .A1(n6892), .A2(n12048), .A3(n12047), .ZN(n12046) );
  NAND2_X1 U9428 ( .A1(n12040), .A2(n12043), .ZN(n6892) );
  NAND2_X1 U9429 ( .A1(n8220), .A2(n12296), .ZN(n13454) );
  NAND2_X1 U9430 ( .A1(n8122), .A2(n8121), .ZN(n13555) );
  NAND2_X1 U9431 ( .A1(n7959), .A2(n7958), .ZN(n10673) );
  NAND2_X1 U9432 ( .A1(n7164), .A2(n7163), .ZN(n7162) );
  NAND2_X1 U9433 ( .A1(n14086), .A2(n7335), .ZN(n7338) );
  NAND2_X1 U9434 ( .A1(n11717), .A2(n7416), .ZN(n6899) );
  XNOR2_X1 U9435 ( .A(n14445), .B(n7471), .ZN(n14481) );
  NAND2_X1 U9436 ( .A1(n12931), .A2(n11283), .ZN(n12915) );
  XNOR2_X1 U9437 ( .A(n9252), .B(n15074), .ZN(n15067) );
  NAND2_X1 U9438 ( .A1(n10109), .A2(n10108), .ZN(n10201) );
  NAND2_X1 U9439 ( .A1(n10203), .A2(n10116), .ZN(n10426) );
  NAND2_X1 U9440 ( .A1(n6902), .A2(n6900), .ZN(P1_U3214) );
  NAND2_X1 U9441 ( .A1(n7176), .A2(n14612), .ZN(n6902) );
  NAND2_X1 U9442 ( .A1(n12510), .A2(n13789), .ZN(n13791) );
  NAND2_X1 U9443 ( .A1(n13777), .A2(n12440), .ZN(n12444) );
  NAND2_X1 U9444 ( .A1(n10154), .A2(n10153), .ZN(n10321) );
  NAND2_X1 U9445 ( .A1(n12500), .A2(n13892), .ZN(n13790) );
  NAND2_X1 U9446 ( .A1(n7618), .A2(n7619), .ZN(n13836) );
  OR2_X2 U9447 ( .A1(n9711), .A2(n9710), .ZN(n7635) );
  OAI22_X1 U9448 ( .A1(n9355), .A2(n9354), .B1(n9353), .B2(n9352), .ZN(n9356)
         );
  NAND2_X1 U9449 ( .A1(n7592), .A2(n7590), .ZN(n8066) );
  AOI21_X1 U9450 ( .B1(n7125), .B2(n7127), .A(n6670), .ZN(n7123) );
  NAND2_X1 U9451 ( .A1(n6905), .A2(n6903), .ZN(P2_U3186) );
  NAND3_X1 U9452 ( .A1(n6965), .A2(n13227), .A3(n13125), .ZN(n6905) );
  NAND3_X1 U9453 ( .A1(n10918), .A2(n10917), .A3(n6543), .ZN(n7203) );
  NAND2_X1 U9454 ( .A1(n12684), .A2(n9878), .ZN(n11842) );
  INV_X1 U9455 ( .A(n10930), .ZN(n10928) );
  NAND2_X2 U9456 ( .A1(n6534), .A2(n9161), .ZN(n11198) );
  NAND2_X1 U9457 ( .A1(n15047), .A2(n9903), .ZN(n11841) );
  NOR2_X1 U9458 ( .A1(n12825), .A2(n12826), .ZN(n12824) );
  NAND3_X1 U9459 ( .A1(n9249), .A2(n6648), .A3(n9250), .ZN(n15074) );
  NAND2_X1 U9460 ( .A1(n15067), .A2(n15066), .ZN(n7212) );
  NAND2_X1 U9461 ( .A1(n7131), .A2(n11187), .ZN(n7797) );
  NAND2_X1 U9462 ( .A1(n7809), .A2(n7808), .ZN(n8195) );
  NAND2_X1 U9463 ( .A1(n7154), .A2(n7153), .ZN(n7592) );
  NAND2_X1 U9464 ( .A1(n7146), .A2(n14892), .ZN(n7145) );
  NAND2_X1 U9465 ( .A1(n10327), .A2(n7610), .ZN(n7609) );
  INV_X1 U9466 ( .A(n12525), .ZN(n8819) );
  NAND2_X1 U9467 ( .A1(n8826), .A2(n8882), .ZN(n8881) );
  NAND2_X1 U9468 ( .A1(n9318), .A2(n9317), .ZN(n9378) );
  NAND2_X1 U9469 ( .A1(n9373), .A2(n9377), .ZN(n11742) );
  AND2_X2 U9470 ( .A1(n9323), .A2(n9718), .ZN(n13557) );
  INV_X1 U9471 ( .A(n6941), .ZN(n7143) );
  NAND2_X1 U9472 ( .A1(n10301), .A2(n10300), .ZN(n10299) );
  NAND2_X1 U9473 ( .A1(n13624), .A2(n6683), .ZN(P2_U3527) );
  NAND2_X1 U9474 ( .A1(n13709), .A2(n6684), .ZN(P2_U3495) );
  NAND2_X1 U9475 ( .A1(n10673), .A2(n7975), .ZN(n7270) );
  NAND2_X1 U9476 ( .A1(n7913), .A2(n7912), .ZN(n10301) );
  NAND2_X1 U9477 ( .A1(n13622), .A2(n14927), .ZN(n7164) );
  NAND2_X1 U9478 ( .A1(n7880), .A2(n7879), .ZN(n10098) );
  NOR2_X1 U9479 ( .A1(n13620), .A2(n7162), .ZN(n7161) );
  OAI21_X1 U9480 ( .B1(n13505), .B2(n13506), .A(n6667), .ZN(n6968) );
  NAND2_X1 U9481 ( .A1(n8391), .A2(n8390), .ZN(n8800) );
  OAI21_X1 U9482 ( .B1(n11389), .B2(n11388), .A(n11387), .ZN(n11396) );
  NAND2_X1 U9483 ( .A1(n11619), .A2(n11618), .ZN(n7552) );
  NAND2_X1 U9484 ( .A1(n14481), .A2(n14480), .ZN(n7470) );
  NAND2_X1 U9485 ( .A1(n15443), .A2(n15444), .ZN(n7098) );
  OAI21_X1 U9486 ( .B1(n14428), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6650), .ZN(
        n6930) );
  NAND2_X1 U9487 ( .A1(n14483), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7465) );
  OAI21_X1 U9488 ( .B1(n14484), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6649), .ZN(
        n7097) );
  OR2_X1 U9489 ( .A1(n10168), .A2(n7852), .ZN(n14897) );
  NAND2_X1 U9490 ( .A1(n7366), .A2(n7365), .ZN(n10302) );
  NOR2_X2 U9491 ( .A1(n13643), .A2(n13484), .ZN(n13472) );
  NOR2_X1 U9492 ( .A1(n7654), .A2(n7653), .ZN(n7652) );
  NAND2_X1 U9493 ( .A1(n12163), .A2(n12162), .ZN(n6918) );
  AOI21_X1 U9494 ( .B1(n12107), .B2(n12106), .A(n12104), .ZN(n12105) );
  NAND2_X1 U9495 ( .A1(n6935), .A2(n6934), .ZN(n7670) );
  NAND2_X1 U9496 ( .A1(n7656), .A2(n12165), .ZN(n7655) );
  OAI21_X1 U9497 ( .B1(n6549), .B2(n6919), .A(n6663), .ZN(n7679) );
  INV_X1 U9498 ( .A(n12066), .ZN(n7668) );
  CLKBUF_X3 U9499 ( .A(n12070), .Z(n12242) );
  NAND2_X1 U9500 ( .A1(n7228), .A2(n7649), .ZN(n6933) );
  INV_X1 U9501 ( .A(n7674), .ZN(n6935) );
  NAND3_X1 U9502 ( .A1(n7553), .A2(n7552), .A3(n6669), .ZN(n7559) );
  NAND2_X1 U9503 ( .A1(n7573), .A2(n7575), .ZN(n11605) );
  OR2_X1 U9504 ( .A1(n11583), .A2(n14707), .ZN(n8815) );
  AOI21_X2 U9505 ( .B1(n10147), .B2(n10146), .A(n7695), .ZN(n10154) );
  AOI21_X1 U9506 ( .B1(n8819), .B2(n13957), .A(n6922), .ZN(n8826) );
  INV_X1 U9507 ( .A(n7178), .ZN(n13778) );
  NAND2_X1 U9508 ( .A1(n13778), .A2(n13779), .ZN(n13777) );
  NAND2_X1 U9509 ( .A1(n10321), .A2(n7174), .ZN(n10327) );
  OAI21_X1 U9510 ( .B1(n14610), .B2(n7182), .A(n7179), .ZN(n7178) );
  NOR2_X1 U9511 ( .A1(n9356), .A2(n9357), .ZN(n9711) );
  NAND2_X1 U9512 ( .A1(n13910), .A2(n12541), .ZN(n7177) );
  XNOR2_X1 U9513 ( .A(n7177), .B(n13771), .ZN(n7176) );
  XNOR2_X1 U9515 ( .A(n8396), .B(n8395), .ZN(n14368) );
  NAND2_X1 U9516 ( .A1(n11621), .A2(n11620), .ZN(n7553) );
  INV_X1 U9517 ( .A(n11437), .ZN(n11434) );
  NAND2_X1 U9518 ( .A1(n6925), .A2(n6660), .ZN(n6975) );
  NAND4_X1 U9519 ( .A1(n11444), .A2(n11442), .A3(n11443), .A4(n11441), .ZN(
        n6925) );
  XNOR2_X1 U9520 ( .A(n14459), .B(n14460), .ZN(n14484) );
  NAND2_X1 U9521 ( .A1(n10593), .A2(n10592), .ZN(n14486) );
  NAND2_X1 U9522 ( .A1(n10023), .A2(n10022), .ZN(n10236) );
  NAND2_X1 U9523 ( .A1(n11704), .A2(n11703), .ZN(n14234) );
  NAND2_X1 U9524 ( .A1(n11712), .A2(n11711), .ZN(n14145) );
  NAND2_X1 U9525 ( .A1(n9927), .A2(n9926), .ZN(n10015) );
  NAND2_X1 U9526 ( .A1(n9511), .A2(n9510), .ZN(n9740) );
  NAND2_X1 U9527 ( .A1(n14656), .A2(n6658), .ZN(n11702) );
  NAND2_X1 U9528 ( .A1(n6933), .A2(n12166), .ZN(n12171) );
  OR2_X1 U9529 ( .A1(n6525), .A2(n7821), .ZN(n7825) );
  NAND2_X1 U9530 ( .A1(n7679), .A2(n7681), .ZN(n12207) );
  NAND2_X1 U9531 ( .A1(n6937), .A2(n6936), .ZN(n7667) );
  NAND2_X1 U9532 ( .A1(n12725), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12756) );
  NOR2_X1 U9533 ( .A1(n7699), .A2(n7611), .ZN(n7610) );
  INV_X1 U9534 ( .A(n7506), .ZN(n7505) );
  NAND2_X1 U9535 ( .A1(n7292), .A2(n7293), .ZN(n13456) );
  INV_X1 U9536 ( .A(n13433), .ZN(n7291) );
  OAI21_X1 U9537 ( .B1(n13619), .B2(n13699), .A(n13617), .ZN(n6941) );
  AOI21_X1 U9539 ( .B1(n12885), .B2(n11245), .A(n7697), .ZN(n12865) );
  XNOR2_X1 U9540 ( .A(n7264), .B(n12771), .ZN(n12026) );
  INV_X1 U9541 ( .A(n12020), .ZN(n7361) );
  AOI211_X2 U9542 ( .C1(n12030), .C2(n12029), .A(n12028), .B(n12027), .ZN(
        n12037) );
  XNOR2_X2 U9543 ( .A(n7214), .B(n15338), .ZN(n9051) );
  INV_X1 U9544 ( .A(n9888), .ZN(n7213) );
  NAND2_X1 U9545 ( .A1(n10426), .A2(n10425), .ZN(n10453) );
  NAND3_X1 U9546 ( .A1(n6948), .A2(n12807), .A3(n15068), .ZN(n6947) );
  NAND2_X1 U9547 ( .A1(n6949), .A2(n12007), .ZN(n6948) );
  INV_X1 U9548 ( .A(n12808), .ZN(n6949) );
  NAND2_X1 U9549 ( .A1(n6953), .A2(n6950), .ZN(P3_U3455) );
  OR2_X1 U9550 ( .A1(n13047), .A2(n15125), .ZN(n6953) );
  NAND2_X1 U9551 ( .A1(n7464), .A2(n14511), .ZN(n7463) );
  NAND2_X1 U9552 ( .A1(n14512), .A2(n14513), .ZN(n14511) );
  NAND2_X1 U9553 ( .A1(n14463), .A2(n14694), .ZN(n7106) );
  OAI21_X1 U9554 ( .B1(n14431), .B2(n14430), .A(n7468), .ZN(n7467) );
  NAND2_X1 U9555 ( .A1(n7655), .A2(n7651), .ZN(n12163) );
  XNOR2_X1 U9556 ( .A(n12115), .B(n6529), .ZN(n11134) );
  NAND2_X1 U9557 ( .A1(n10753), .A2(n10752), .ZN(n14656) );
  NAND2_X1 U9558 ( .A1(n6978), .A2(n6976), .ZN(n11531) );
  NAND2_X1 U9559 ( .A1(n6975), .A2(n6973), .ZN(n11469) );
  OAI21_X1 U9560 ( .B1(n11370), .B2(n7540), .A(n7539), .ZN(n11371) );
  NAND3_X1 U9561 ( .A1(n8610), .A2(n7199), .A3(n8611), .ZN(n8614) );
  NAND2_X2 U9562 ( .A1(n14109), .A2(n14108), .ZN(n14294) );
  NAND3_X1 U9563 ( .A1(n14282), .A2(n14281), .A3(n6960), .ZN(n14351) );
  NOR2_X2 U9564 ( .A1(n14202), .A2(n14203), .ZN(n14201) );
  NAND2_X1 U9565 ( .A1(n7431), .A2(n8318), .ZN(n10071) );
  XNOR2_X1 U9566 ( .A(n8358), .B(n7147), .ZN(n7146) );
  NAND3_X1 U9567 ( .A1(n7315), .A2(n9766), .A3(n7314), .ZN(n9925) );
  NAND2_X1 U9568 ( .A1(n7300), .A2(n7299), .ZN(n10591) );
  AOI21_X2 U9569 ( .B1(n14200), .B2(n14203), .A(n11708), .ZN(n14191) );
  NAND4_X1 U9570 ( .A1(n8611), .A2(n8610), .A3(n6672), .A4(n7199), .ZN(n7427)
         );
  NAND2_X1 U9571 ( .A1(n8809), .A2(n7311), .ZN(n7306) );
  NAND2_X1 U9572 ( .A1(n7663), .A2(n7650), .ZN(n7649) );
  INV_X1 U9573 ( .A(n10098), .ZN(n6966) );
  OR2_X1 U9574 ( .A1(n12081), .A2(n7690), .ZN(n7688) );
  NAND2_X1 U9575 ( .A1(n7278), .A2(n7279), .ZN(n13505) );
  INV_X1 U9576 ( .A(n6968), .ZN(n13495) );
  XNOR2_X1 U9577 ( .A(n12342), .B(n12343), .ZN(n13215) );
  AND3_X4 U9578 ( .A1(n7244), .A2(n7678), .A3(n7676), .ZN(n8263) );
  XNOR2_X1 U9579 ( .A(n13601), .B(n6529), .ZN(n10396) );
  NAND2_X1 U9580 ( .A1(n13124), .A2(n13123), .ZN(n6965) );
  NOR3_X2 U9581 ( .A1(n12384), .A2(n12345), .A3(n11111), .ZN(n12391) );
  NAND2_X1 U9582 ( .A1(n7142), .A2(n7140), .ZN(P2_U3528) );
  NAND2_X1 U9583 ( .A1(n7124), .A2(n7123), .ZN(n13154) );
  INV_X2 U9584 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15392) );
  XNOR2_X1 U9585 ( .A(n7731), .B(SI_1_), .ZN(n7831) );
  NAND4_X1 U9586 ( .A1(n11472), .A2(n11471), .A3(n14218), .A4(n14199), .ZN(
        n6972) );
  NAND3_X1 U9587 ( .A1(n11505), .A2(n7579), .A3(n11504), .ZN(n6978) );
  NAND2_X1 U9588 ( .A1(n15440), .A2(n15439), .ZN(n6979) );
  INV_X1 U9589 ( .A(n14516), .ZN(n7096) );
  INV_X1 U9590 ( .A(n14691), .ZN(n7107) );
  XNOR2_X1 U9591 ( .A(n7095), .B(n6585), .ZN(SUB_1596_U4) );
  NAND2_X1 U9592 ( .A1(n7212), .A2(n9886), .ZN(n15042) );
  NAND2_X1 U9593 ( .A1(n7374), .A2(n7373), .ZN(n13395) );
  NAND2_X1 U9594 ( .A1(n13540), .A2(n13731), .ZN(n13527) );
  NAND2_X1 U9595 ( .A1(n10180), .A2(n14947), .ZN(n10099) );
  INV_X1 U9596 ( .A(n10099), .ZN(n7366) );
  OR2_X1 U9597 ( .A1(n14897), .A2(n14901), .ZN(n14898) );
  NAND2_X1 U9598 ( .A1(n7371), .A2(n7370), .ZN(n13499) );
  NOR2_X2 U9599 ( .A1(n13447), .A2(n13440), .ZN(n13436) );
  NOR2_X4 U9600 ( .A1(n10815), .A2(n13587), .ZN(n10818) );
  NAND2_X1 U9601 ( .A1(n14352), .A2(n6528), .ZN(n6983) );
  OR2_X1 U9602 ( .A1(n6582), .A2(n14764), .ZN(n6985) );
  NAND2_X1 U9603 ( .A1(n7341), .A2(n7340), .ZN(n14200) );
  NAND2_X1 U9604 ( .A1(n7666), .A2(n12193), .ZN(n7665) );
  NAND2_X1 U9605 ( .A1(n12055), .A2(n12061), .ZN(n7224) );
  INV_X1 U9606 ( .A(n7656), .ZN(n7228) );
  OAI21_X1 U9607 ( .B1(n7855), .B2(n9538), .A(n7648), .ZN(n7647) );
  NAND2_X1 U9608 ( .A1(n8091), .A2(n7488), .ZN(n8297) );
  NAND2_X1 U9609 ( .A1(n7225), .A2(n7219), .ZN(n12067) );
  NAND2_X1 U9610 ( .A1(n12057), .A2(n12061), .ZN(n7223) );
  AND2_X2 U9611 ( .A1(n7496), .A2(n7495), .ZN(n10051) );
  INV_X1 U9612 ( .A(n14035), .ZN(n14036) );
  NAND2_X1 U9613 ( .A1(n12395), .A2(n12394), .ZN(n13124) );
  NAND2_X1 U9614 ( .A1(n11742), .A2(n9573), .ZN(n11743) );
  INV_X1 U9615 ( .A(n13215), .ZN(n7111) );
  NAND2_X1 U9616 ( .A1(n12379), .A2(n6653), .ZN(P3_U3204) );
  NAND2_X1 U9617 ( .A1(n6668), .A2(n6556), .ZN(P3_U3456) );
  NAND3_X1 U9618 ( .A1(n6993), .A2(n6992), .A3(n7574), .ZN(n7573) );
  NAND2_X1 U9619 ( .A1(n11579), .A2(n11578), .ZN(n6992) );
  NAND2_X1 U9620 ( .A1(n11575), .A2(n11574), .ZN(n6993) );
  NAND2_X1 U9621 ( .A1(n12880), .A2(n12879), .ZN(n11286) );
  INV_X1 U9622 ( .A(n10201), .ZN(n7207) );
  NAND3_X1 U9623 ( .A1(n7002), .A2(n7000), .A3(n6998), .ZN(P2_U3233) );
  INV_X1 U9624 ( .A(n9664), .ZN(n9666) );
  OR2_X1 U9625 ( .A1(n7527), .A2(n7524), .ZN(n7015) );
  NAND2_X1 U9626 ( .A1(n7022), .A2(n9985), .ZN(n7016) );
  NAND3_X1 U9627 ( .A1(n7018), .A2(n7523), .A3(n7022), .ZN(n7017) );
  NAND3_X1 U9628 ( .A1(n7525), .A2(n9544), .A3(n7022), .ZN(n7021) );
  AOI21_X1 U9629 ( .B1(n7025), .B2(n7523), .A(n7024), .ZN(n9992) );
  INV_X1 U9630 ( .A(n7524), .ZN(n7523) );
  NAND2_X1 U9631 ( .A1(n11754), .A2(n7035), .ZN(n7033) );
  NAND2_X1 U9632 ( .A1(n12627), .A2(n6540), .ZN(n7042) );
  OAI21_X1 U9633 ( .B1(n12627), .B2(n7045), .A(n6546), .ZN(n11783) );
  NAND2_X1 U9634 ( .A1(n8858), .A2(n7046), .ZN(n9177) );
  NAND2_X1 U9635 ( .A1(n12766), .A2(n6692), .ZN(n7048) );
  OAI211_X1 U9636 ( .C1(n12766), .C2(n14529), .A(n7049), .B(n7048), .ZN(n14525) );
  OAI211_X2 U9637 ( .C1(n9065), .C2(n7051), .A(n7052), .B(n7050), .ZN(n9069)
         );
  NAND2_X1 U9638 ( .A1(n7055), .A2(n7054), .ZN(n12720) );
  NAND2_X1 U9639 ( .A1(n12689), .A2(n12711), .ZN(n7054) );
  NAND2_X1 U9640 ( .A1(n7056), .A2(n7057), .ZN(n7055) );
  INV_X1 U9641 ( .A(n10956), .ZN(n7056) );
  NAND2_X1 U9642 ( .A1(n10650), .A2(n7063), .ZN(n7061) );
  NOR2_X1 U9643 ( .A1(n10649), .A2(n10650), .ZN(n10653) );
  NOR2_X1 U9644 ( .A1(n10523), .A2(n14586), .ZN(n10649) );
  INV_X1 U9645 ( .A(n10652), .ZN(n7063) );
  NAND2_X1 U9646 ( .A1(n8483), .A2(n7070), .ZN(n7068) );
  NAND2_X1 U9647 ( .A1(n7073), .A2(n7075), .ZN(n10585) );
  NAND3_X1 U9648 ( .A1(n7362), .A2(n10370), .A3(n9835), .ZN(n7073) );
  NAND2_X1 U9649 ( .A1(n7080), .A2(n7078), .ZN(n9343) );
  NAND3_X1 U9650 ( .A1(n7091), .A2(n7090), .A3(n12826), .ZN(n11957) );
  NAND2_X1 U9651 ( .A1(n14472), .A2(n7101), .ZN(n7100) );
  INV_X1 U9652 ( .A(n9317), .ZN(n9321) );
  AND2_X4 U9653 ( .A1(n10068), .A2(n7130), .ZN(n12356) );
  NAND2_X1 U9654 ( .A1(n12360), .A2(n7113), .ZN(n7112) );
  OAI211_X1 U9655 ( .C1(n12360), .C2(n7117), .A(n7114), .B(n7112), .ZN(n12407)
         );
  NAND2_X2 U9656 ( .A1(n12360), .A2(n12359), .ZN(n12395) );
  INV_X1 U9657 ( .A(n10418), .ZN(n7129) );
  XNOR2_X1 U9658 ( .A(n7130), .B(n7129), .ZN(n8309) );
  OAI22_X1 U9659 ( .A1(n7433), .A2(n13444), .B1(n7435), .B2(n7432), .ZN(n13401) );
  NAND3_X1 U9660 ( .A1(n7132), .A2(n13402), .A3(n14892), .ZN(n13404) );
  NAND2_X1 U9661 ( .A1(n7820), .A2(n7819), .ZN(n13440) );
  NAND2_X1 U9662 ( .A1(n7820), .A2(n7137), .ZN(n7136) );
  INV_X1 U9663 ( .A(n7812), .ZN(n7152) );
  NAND2_X1 U9664 ( .A1(n7978), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U9665 ( .A1(n7978), .A2(n7763), .ZN(n7160) );
  MUX2_X1 U9666 ( .A(n13623), .B(n7161), .S(n14972), .Z(n13624) );
  MUX2_X1 U9667 ( .A(n15376), .B(n7161), .S(n14962), .Z(n13709) );
  INV_X1 U9668 ( .A(n7806), .ZN(n7173) );
  NAND2_X1 U9669 ( .A1(n12463), .A2(n6542), .ZN(n7186) );
  NAND2_X1 U9670 ( .A1(n7186), .A2(n7187), .ZN(n12500) );
  INV_X1 U9671 ( .A(n14674), .ZN(n8808) );
  NAND2_X4 U9672 ( .A1(n7196), .A2(n14674), .ZN(n12525) );
  NAND2_X1 U9673 ( .A1(n10918), .A2(n10917), .ZN(n15018) );
  NAND2_X1 U9674 ( .A1(n7205), .A2(n9065), .ZN(n8479) );
  INV_X1 U9675 ( .A(n12198), .ZN(n7217) );
  INV_X1 U9676 ( .A(n12055), .ZN(n7222) );
  NAND3_X1 U9677 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(n7219) );
  INV_X1 U9678 ( .A(n12060), .ZN(n7226) );
  OAI21_X1 U9679 ( .B1(n12122), .B2(n7657), .A(n7703), .ZN(n7656) );
  NAND3_X1 U9680 ( .A1(n6592), .A2(n7236), .A3(n7231), .ZN(n7230) );
  AND2_X1 U9681 ( .A1(n7240), .A2(n7239), .ZN(n7232) );
  NAND2_X1 U9682 ( .A1(n7242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7816) );
  NAND4_X1 U9683 ( .A1(n7244), .A2(n7676), .A3(n7298), .A4(n7243), .ZN(n7242)
         );
  NAND2_X1 U9684 ( .A1(n10904), .A2(n7251), .ZN(n7250) );
  INV_X1 U9685 ( .A(n11017), .ZN(n11018) );
  NAND3_X1 U9686 ( .A1(n7265), .A2(n7359), .A3(n7358), .ZN(n7264) );
  NAND2_X1 U9688 ( .A1(n7270), .A2(n7268), .ZN(n7995) );
  NAND2_X1 U9689 ( .A1(n7272), .A2(n7271), .ZN(n7913) );
  AND2_X1 U9690 ( .A1(n12273), .A2(n7929), .ZN(n7277) );
  NAND2_X1 U9691 ( .A1(n13555), .A2(n7280), .ZN(n7278) );
  NAND2_X1 U9692 ( .A1(n13477), .A2(n7294), .ZN(n7292) );
  INV_X1 U9693 ( .A(n13456), .ZN(n8220) );
  AND2_X2 U9694 ( .A1(n7712), .A2(n7713), .ZN(n7298) );
  NAND2_X1 U9695 ( .A1(n10236), .A2(n7302), .ZN(n7300) );
  NOR2_X1 U9696 ( .A1(n7304), .A2(n7303), .ZN(n7302) );
  NOR2_X1 U9697 ( .A1(n10235), .A2(n7305), .ZN(n7303) );
  NAND2_X1 U9698 ( .A1(n9740), .A2(n7317), .ZN(n7315) );
  NAND2_X1 U9699 ( .A1(n7325), .A2(n7327), .ZN(n14261) );
  NAND2_X1 U9700 ( .A1(n14486), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U9701 ( .A1(n14086), .A2(n7339), .ZN(n11717) );
  NAND2_X1 U9702 ( .A1(n14234), .A2(n7342), .ZN(n7341) );
  XNOR2_X1 U9703 ( .A(n13954), .B(n11372), .ZN(n11645) );
  INV_X1 U9704 ( .A(n14261), .ZN(n10753) );
  NAND2_X1 U9705 ( .A1(n8587), .A2(n8586), .ZN(n7344) );
  NAND2_X1 U9706 ( .A1(n8532), .A2(n8531), .ZN(n7345) );
  OR2_X1 U9707 ( .A1(n11151), .A2(n7353), .ZN(n7349) );
  NAND2_X1 U9708 ( .A1(n11151), .A2(n7355), .ZN(n7350) );
  NAND2_X1 U9709 ( .A1(n7349), .A2(n7351), .ZN(n11970) );
  NAND2_X1 U9710 ( .A1(n11151), .A2(n11150), .ZN(n11960) );
  NAND2_X1 U9711 ( .A1(n12022), .A2(n12986), .ZN(n7358) );
  INV_X1 U9712 ( .A(n12021), .ZN(n7359) );
  NOR2_X2 U9713 ( .A1(n10302), .A2(n12091), .ZN(n10409) );
  NOR2_X2 U9714 ( .A1(n13558), .A2(n13672), .ZN(n13540) );
  NOR2_X2 U9715 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  INV_X1 U9716 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7378) );
  INV_X1 U9717 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7376) );
  NAND4_X1 U9718 ( .A1(n8433), .A2(n7380), .A3(n7379), .A4(n7378), .ZN(n7377)
         );
  INV_X1 U9719 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8433) );
  NOR2_X1 U9720 ( .A1(n14260), .A2(n10736), .ZN(n7387) );
  NAND2_X1 U9721 ( .A1(n14248), .A2(n7386), .ZN(n7383) );
  NAND2_X1 U9722 ( .A1(n7399), .A2(n7402), .ZN(n10613) );
  OR2_X1 U9723 ( .A1(n10214), .A2(n7404), .ZN(n7399) );
  INV_X1 U9724 ( .A(n10213), .ZN(n7400) );
  NAND2_X1 U9725 ( .A1(n7401), .A2(n7405), .ZN(n10611) );
  NAND2_X1 U9726 ( .A1(n10214), .A2(n7407), .ZN(n7401) );
  AOI21_X1 U9727 ( .B1(n7405), .B2(n7403), .A(n10590), .ZN(n7402) );
  INV_X1 U9728 ( .A(n7407), .ZN(n7403) );
  INV_X1 U9729 ( .A(n7405), .ZN(n7404) );
  NAND2_X1 U9730 ( .A1(n14101), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U9731 ( .A1(n14101), .A2(n6581), .ZN(n7417) );
  NAND2_X1 U9732 ( .A1(n14101), .A2(n6577), .ZN(n14089) );
  NAND2_X1 U9733 ( .A1(n9524), .A2(n7422), .ZN(n7421) );
  INV_X1 U9734 ( .A(n7427), .ZN(n8809) );
  NAND2_X1 U9735 ( .A1(n7427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8811) );
  OAI21_X1 U9736 ( .B1(n10176), .B2(n7430), .A(n7428), .ZN(n7431) );
  OAI21_X1 U9737 ( .B1(n10175), .B2(n7430), .A(n8316), .ZN(n7429) );
  INV_X1 U9738 ( .A(n8315), .ZN(n7430) );
  AOI21_X2 U9739 ( .B1(n7438), .B2(n8355), .A(n6636), .ZN(n7437) );
  NAND2_X1 U9740 ( .A1(n13401), .A2(n13406), .ZN(n13402) );
  INV_X1 U9741 ( .A(n8312), .ZN(n12265) );
  NAND2_X1 U9742 ( .A1(n7448), .A2(n7449), .ZN(n8327) );
  NAND2_X1 U9743 ( .A1(n10771), .A2(n8326), .ZN(n7448) );
  OAI21_X2 U9744 ( .B1(n13535), .B2(n7453), .A(n7451), .ZN(n13490) );
  NAND2_X1 U9745 ( .A1(n7455), .A2(n7456), .ZN(n10677) );
  NAND2_X1 U9746 ( .A1(n10405), .A2(n7457), .ZN(n7455) );
  INV_X1 U9747 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7461) );
  NOR2_X2 U9748 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7472) );
  NOR2_X2 U9749 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7473) );
  AND2_X2 U9750 ( .A1(n7473), .A2(n7472), .ZN(n8049) );
  NAND2_X1 U9751 ( .A1(n13154), .A2(n12341), .ZN(n12342) );
  OR2_X1 U9752 ( .A1(n10379), .A2(n10380), .ZN(n7478) );
  NAND4_X1 U9753 ( .A1(n8611), .A2(n8610), .A3(n7199), .A4(n8612), .ZN(n7494)
         );
  NAND2_X1 U9754 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
  AND2_X1 U9755 ( .A1(n8441), .A2(n6695), .ZN(n7504) );
  OAI21_X1 U9756 ( .B1(n8439), .B2(n8438), .A(n7507), .ZN(n7506) );
  NAND2_X1 U9757 ( .A1(n8438), .A2(n8713), .ZN(n7507) );
  INV_X1 U9758 ( .A(n11783), .ZN(n7516) );
  AOI21_X1 U9759 ( .B1(n7516), .B2(n6624), .A(n7517), .ZN(n11791) );
  AND2_X1 U9760 ( .A1(n8407), .A2(n8543), .ZN(n8858) );
  AND2_X1 U9761 ( .A1(n7530), .A2(n8543), .ZN(n8416) );
  AOI22_X1 U9762 ( .A1(n11368), .A2(n11348), .B1(n11373), .B2(n11369), .ZN(
        n7539) );
  AND2_X1 U9763 ( .A1(n7551), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U9764 ( .A1(n7567), .A2(n7568), .ZN(n11405) );
  NAND2_X1 U9765 ( .A1(n8390), .A2(n6662), .ZN(n8604) );
  INV_X1 U9766 ( .A(n8604), .ZN(n8600) );
  INV_X1 U9767 ( .A(n11517), .ZN(n7580) );
  INV_X1 U9768 ( .A(n11451), .ZN(n7582) );
  NAND3_X1 U9769 ( .A1(n7584), .A2(n11328), .A3(n11327), .ZN(n13753) );
  NAND3_X1 U9770 ( .A1(n12300), .A2(n12298), .A3(n7589), .ZN(n7588) );
  NAND2_X1 U9771 ( .A1(n8016), .A2(n8015), .ZN(n8018) );
  OAI21_X1 U9772 ( .B1(n7813), .B2(n7599), .A(n7597), .ZN(n8252) );
  NAND2_X1 U9773 ( .A1(n7798), .A2(n7797), .ZN(n8142) );
  INV_X1 U9774 ( .A(n10501), .ZN(n7616) );
  INV_X1 U9775 ( .A(n10500), .ZN(n7617) );
  NAND2_X1 U9776 ( .A1(n13791), .A2(n7622), .ZN(n7618) );
  OAI211_X1 U9777 ( .C1(n13910), .C2(n6671), .A(n7628), .B(n7626), .ZN(n12563)
         );
  OAI22_X1 U9778 ( .A1(n7630), .A2(n7627), .B1(n12557), .B2(n7632), .ZN(n7626)
         );
  NOR2_X1 U9779 ( .A1(n13771), .A2(n12557), .ZN(n7627) );
  NAND2_X1 U9780 ( .A1(n13910), .A2(n7629), .ZN(n7628) );
  NOR2_X1 U9781 ( .A1(n12557), .A2(n7630), .ZN(n7629) );
  INV_X1 U9782 ( .A(n12557), .ZN(n7631) );
  OAI22_X2 U9783 ( .A1(n9823), .A2(n9822), .B1(n7635), .B2(n9821), .ZN(n10147)
         );
  XNOR2_X2 U9784 ( .A(n7635), .B(n9821), .ZN(n9823) );
  XNOR2_X2 U9785 ( .A(n12444), .B(n12445), .ZN(n13923) );
  NAND3_X1 U9786 ( .A1(n7718), .A2(n12373), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7648) );
  INV_X1 U9787 ( .A(n7647), .ZN(n7646) );
  NAND2_X1 U9788 ( .A1(n12122), .A2(n12121), .ZN(n7663) );
  NAND2_X1 U9789 ( .A1(n7673), .A2(n7672), .ZN(n7671) );
  INV_X1 U9790 ( .A(n12179), .ZN(n7672) );
  INV_X1 U9791 ( .A(n7675), .ZN(n13747) );
  INV_X1 U9792 ( .A(n9252), .ZN(n12685) );
  NAND2_X2 U9793 ( .A1(n11005), .A2(n11004), .ZN(n11754) );
  AOI22_X1 U9794 ( .A1(n9019), .A2(n9230), .B1(n8823), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n8824) );
  AOI22_X2 U9795 ( .A1(n12417), .A2(n12416), .B1(n12415), .B2(n12414), .ZN(
        n14610) );
  NAND3_X1 U9796 ( .A1(n11743), .A2(n9578), .A3(n9575), .ZN(n13183) );
  INV_X1 U9797 ( .A(n8416), .ZN(n9056) );
  NAND2_X1 U9798 ( .A1(n14890), .A2(n14891), .ZN(n14889) );
  NAND2_X4 U9799 ( .A1(n8360), .A2(n13761), .ZN(n8899) );
  NAND4_X2 U9800 ( .A1(n7826), .A2(n7825), .A3(n7824), .A4(n7823), .ZN(n13269)
         );
  NAND2_X1 U9801 ( .A1(n8361), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U9802 ( .A1(n8014), .A2(n8013), .ZN(n10803) );
  NAND2_X1 U9803 ( .A1(n8320), .A2(n8319), .ZN(n10303) );
  OR2_X1 U9804 ( .A1(n11799), .A2(P1_B_REG_SCAN_IN), .ZN(n8573) );
  INV_X1 U9805 ( .A(n13552), .ZN(n8121) );
  NAND2_X2 U9806 ( .A1(n14051), .A2(n14642), .ZN(n14639) );
  INV_X1 U9807 ( .A(n14260), .ZN(n10752) );
  AND2_X1 U9808 ( .A1(n10696), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9809 ( .A1(n10718), .A2(n10872), .ZN(n7692) );
  AND2_X1 U9810 ( .A1(n10145), .A2(n10144), .ZN(n7695) );
  AND2_X1 U9811 ( .A1(n12579), .A2(n11788), .ZN(n7696) );
  INV_X1 U9812 ( .A(n14578), .ZN(n10908) );
  NOR2_X1 U9813 ( .A1(n12868), .A2(n12863), .ZN(n7697) );
  AND2_X1 U9814 ( .A1(n7989), .A2(n10393), .ZN(n7698) );
  INV_X1 U9815 ( .A(SI_15_), .ZN(n8694) );
  NAND2_X2 U9816 ( .A1(n8308), .A2(n13595), .ZN(n13598) );
  INV_X1 U9817 ( .A(n13582), .ZN(n14883) );
  AND2_X1 U9818 ( .A1(n10784), .A2(n10783), .ZN(n7699) );
  OR2_X1 U9819 ( .A1(n13619), .A2(n13582), .ZN(n7700) );
  NOR3_X1 U9820 ( .A1(n12297), .A2(n12296), .A3(n12295), .ZN(n7701) );
  INV_X1 U9821 ( .A(n12296), .ZN(n13457) );
  AND2_X1 U9822 ( .A1(n12145), .A2(n12144), .ZN(n7703) );
  OR2_X1 U9823 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  INV_X1 U9824 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8409) );
  INV_X1 U9825 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8410) );
  INV_X1 U9826 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8404) );
  CLKBUF_X3 U9827 ( .A(n12070), .Z(n12237) );
  INV_X1 U9828 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8381) );
  AND2_X1 U9829 ( .A1(n7977), .A2(n7980), .ZN(n7763) );
  AND2_X1 U9830 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  INV_X1 U9831 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7922) );
  INV_X1 U9832 ( .A(n13261), .ZN(n12099) );
  INV_X1 U9833 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10602) );
  INV_X1 U9834 ( .A(n14125), .ZN(n11714) );
  INV_X1 U9835 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U9836 ( .A1(n7771), .A2(n8591), .ZN(n7774) );
  INV_X1 U9837 ( .A(n12771), .ZN(n12023) );
  INV_X1 U9838 ( .A(n12569), .ZN(n8716) );
  NAND2_X1 U9839 ( .A1(n11237), .A2(n11236), .ZN(n11250) );
  NOR2_X1 U9840 ( .A1(n10935), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n10934) );
  INV_X1 U9841 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10255) );
  OR2_X1 U9842 ( .A1(n9176), .A2(n9175), .ZN(n9421) );
  INV_X1 U9843 ( .A(n9421), .ZN(n9186) );
  OR2_X1 U9844 ( .A1(n9833), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9834) );
  AND2_X1 U9845 ( .A1(n9865), .A2(n9860), .ZN(n9861) );
  NAND2_X1 U9846 ( .A1(n7720), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U9847 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8200), .ZN(n8212) );
  NAND2_X1 U9848 ( .A1(n8147), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8161) );
  NOR2_X1 U9849 ( .A1(n8280), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8269) );
  AND2_X1 U9850 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  INV_X1 U9851 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U9852 ( .A1(n15270), .A2(n11541), .ZN(n11553) );
  NAND2_X1 U9853 ( .A1(n11508), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11519) );
  INV_X1 U9854 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10617) );
  AND2_X1 U9855 ( .A1(n8889), .A2(n8827), .ZN(n8834) );
  OR2_X1 U9856 ( .A1(n8797), .A2(n8796), .ZN(n9218) );
  NAND2_X1 U9857 ( .A1(n7782), .A2(n8867), .ZN(n8082) );
  NOR2_X1 U9858 ( .A1(n14422), .A2(n14421), .ZN(n14401) );
  OAI21_X1 U9859 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15157), .A(n14408), .ZN(
        n14469) );
  NAND2_X1 U9860 ( .A1(n9260), .A2(n9257), .ZN(n9479) );
  AND2_X1 U9861 ( .A1(n11022), .A2(n15147), .ZN(n11168) );
  INV_X1 U9862 ( .A(n13000), .ZN(n12667) );
  AND4_X1 U9863 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n12575) );
  AND2_X1 U9864 ( .A1(n8567), .A2(n10581), .ZN(n8420) );
  NAND2_X1 U9865 ( .A1(n11167), .A2(n11168), .ZN(n11180) );
  OR2_X1 U9866 ( .A1(n10872), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10935) );
  INV_X1 U9867 ( .A(n11859), .ZN(n10420) );
  OR2_X1 U9868 ( .A1(n9556), .A2(n11730), .ZN(n9424) );
  NAND2_X1 U9869 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  OR2_X1 U9870 ( .A1(n11244), .A2(n12886), .ZN(n12863) );
  INV_X1 U9871 ( .A(n12946), .ZN(n12949) );
  NOR2_X1 U9872 ( .A1(n9423), .A2(n9186), .ZN(n9409) );
  AND2_X1 U9873 ( .A1(n9688), .A2(n9344), .ZN(n9345) );
  AND2_X1 U9874 ( .A1(n8865), .A2(n8692), .ZN(n8862) );
  AND2_X1 U9875 ( .A1(n8454), .A2(n8453), .ZN(n8496) );
  INV_X1 U9876 ( .A(n13123), .ZN(n12398) );
  OR2_X1 U9877 ( .A1(n11806), .A2(n10374), .ZN(n10375) );
  OR2_X1 U9878 ( .A1(n12325), .A2(n12324), .ZN(n12326) );
  AND2_X1 U9879 ( .A1(n8136), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8147) );
  INV_X1 U9880 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11802) );
  INV_X1 U9881 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n13312) );
  INV_X1 U9882 ( .A(n13246), .ZN(n13192) );
  INV_X1 U9883 ( .A(n14819), .ZN(n10897) );
  INV_X1 U9884 ( .A(n12273), .ZN(n10404) );
  INV_X1 U9885 ( .A(n14892), .ZN(n13509) );
  AND2_X1 U9886 ( .A1(n13861), .A2(n12509), .ZN(n13789) );
  NAND2_X1 U9887 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  INV_X1 U9888 ( .A(n13947), .ZN(n10846) );
  NOR2_X1 U9889 ( .A1(n11461), .A2(n11341), .ZN(n11355) );
  INV_X1 U9890 ( .A(n11630), .ZN(n11606) );
  INV_X1 U9891 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14379) );
  INV_X1 U9892 ( .A(n10642), .ZN(n11448) );
  NOR2_X1 U9893 ( .A1(n8835), .A2(n8834), .ZN(n11689) );
  INV_X1 U9894 ( .A(n11658), .ZN(n10590) );
  INV_X1 U9895 ( .A(n11332), .ZN(n8889) );
  INV_X1 U9896 ( .A(n11365), .ZN(n9746) );
  AND2_X1 U9897 ( .A1(n11364), .A2(n11362), .ZN(n9234) );
  INV_X1 U9898 ( .A(n14633), .ZN(n14222) );
  AND2_X1 U9899 ( .A1(n14043), .A2(n11640), .ZN(n14075) );
  INV_X1 U9900 ( .A(n14793), .ZN(n14759) );
  INV_X1 U9901 ( .A(n14494), .ZN(n14629) );
  INV_X1 U9902 ( .A(n11654), .ZN(n10059) );
  OR2_X1 U9903 ( .A1(n8797), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8799) );
  AND2_X1 U9904 ( .A1(n8082), .A2(n7784), .ZN(n8065) );
  OR2_X1 U9905 ( .A1(n12799), .A2(n10314), .ZN(n12814) );
  AND2_X1 U9906 ( .A1(n9409), .A2(n9262), .ZN(n12643) );
  INV_X1 U9907 ( .A(n12666), .ZN(n12648) );
  INV_X1 U9908 ( .A(n12575), .ZN(n12828) );
  AND4_X1 U9909 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n12872) );
  AND4_X1 U9910 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n12962) );
  INV_X1 U9911 ( .A(n9296), .ZN(n9987) );
  INV_X1 U9912 ( .A(n12791), .ZN(n14990) );
  AND2_X1 U9913 ( .A1(n10313), .A2(n10312), .ZN(n12799) );
  NOR2_X1 U9914 ( .A1(n9431), .A2(n15056), .ZN(n15028) );
  AND3_X1 U9915 ( .A1(n9424), .A2(n9423), .A3(n9422), .ZN(n9560) );
  INV_X1 U9916 ( .A(n12810), .ZN(n12821) );
  OR2_X1 U9917 ( .A1(n15050), .A2(n15118), .ZN(n14601) );
  AND2_X1 U9918 ( .A1(n15056), .A2(n10134), .ZN(n15118) );
  INV_X1 U9919 ( .A(n15046), .ZN(n15065) );
  AND2_X1 U9920 ( .A1(n9198), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9061) );
  INV_X1 U9921 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9050) );
  INV_X1 U9922 ( .A(n14821), .ZN(n13223) );
  AND2_X1 U9923 ( .A1(n10685), .A2(n8376), .ZN(n8897) );
  INV_X1 U9924 ( .A(n14865), .ZN(n13358) );
  AND2_X1 U9925 ( .A1(n8918), .A2(n8917), .ZN(n14865) );
  OR2_X1 U9926 ( .A1(n8914), .A2(n8901), .ZN(n14858) );
  INV_X1 U9927 ( .A(n14858), .ZN(n13380) );
  AND2_X1 U9928 ( .A1(n13598), .A2(n14900), .ZN(n13600) );
  AND2_X1 U9929 ( .A1(n13598), .A2(n12044), .ZN(n14874) );
  INV_X1 U9930 ( .A(n13668), .ZN(n13692) );
  AND2_X1 U9931 ( .A1(n8277), .A2(n8276), .ZN(n14908) );
  AND2_X1 U9932 ( .A1(n8002), .A2(n8032), .ZN(n11076) );
  AND2_X1 U9933 ( .A1(n7903), .A2(n7932), .ZN(n8973) );
  NAND2_X1 U9934 ( .A1(n8833), .A2(n14642), .ZN(n14616) );
  AND4_X1 U9935 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n14042) );
  AND2_X1 U9936 ( .A1(n11361), .A2(n11360), .ZN(n13905) );
  OR2_X1 U9937 ( .A1(n14718), .A2(n11688), .ZN(n10634) );
  INV_X1 U9938 ( .A(n14021), .ZN(n14728) );
  NAND2_X1 U9939 ( .A1(n10744), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11459) );
  INV_X1 U9940 ( .A(n14489), .ZN(n14743) );
  INV_X1 U9941 ( .A(n14738), .ZN(n14259) );
  INV_X1 U9942 ( .A(n9243), .ZN(n9646) );
  OR2_X1 U9943 ( .A1(n9227), .A2(n8828), .ZN(n14793) );
  INV_X1 U9944 ( .A(n14796), .ZN(n14663) );
  AND2_X1 U9945 ( .A1(n8799), .A2(n8798), .ZN(n9243) );
  INV_X1 U9946 ( .A(n14368), .ZN(n8574) );
  INV_X1 U9947 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8388) );
  AND2_X1 U9948 ( .A1(n9077), .A2(n9076), .ZN(n14987) );
  NAND2_X1 U9949 ( .A1(n9197), .A2(n9429), .ZN(n12666) );
  NAND2_X1 U9950 ( .A1(n9190), .A2(n9420), .ZN(n12672) );
  INV_X1 U9951 ( .A(n12936), .ZN(n12908) );
  INV_X1 U9952 ( .A(n12795), .ZN(n14983) );
  OR2_X1 U9953 ( .A1(n15083), .A2(n15034), .ZN(n12968) );
  NAND2_X1 U9954 ( .A1(n9429), .A2(n15056), .ZN(n15040) );
  INV_X2 U9955 ( .A(n15083), .ZN(n15080) );
  NAND2_X1 U9956 ( .A1(n15142), .A2(n14601), .ZN(n13040) );
  AOI21_X1 U9957 ( .B1(n12823), .B2(n12822), .A(n12821), .ZN(n13056) );
  OR2_X1 U9958 ( .A1(n15125), .A2(n10138), .ZN(n13107) );
  INV_X2 U9959 ( .A(n15125), .ZN(n15127) );
  INV_X1 U9960 ( .A(n8567), .ZN(n10768) );
  OR2_X1 U9961 ( .A1(n8861), .A2(n8860), .ZN(n12782) );
  INV_X1 U9962 ( .A(n9610), .ZN(n10271) );
  NAND2_X1 U9963 ( .A1(n9579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14821) );
  INV_X1 U9964 ( .A(n14818), .ZN(n13238) );
  OR2_X1 U9965 ( .A1(n8914), .A2(n13761), .ZN(n14851) );
  INV_X1 U9966 ( .A(n14809), .ZN(n14873) );
  NAND2_X1 U9967 ( .A1(n13598), .A2(n14888), .ZN(n13582) );
  NAND2_X1 U9968 ( .A1(n14972), .A2(n14953), .ZN(n13668) );
  INV_X1 U9969 ( .A(n14972), .ZN(n14970) );
  INV_X1 U9970 ( .A(n13424), .ZN(n13714) );
  INV_X1 U9971 ( .A(n13529), .ZN(n13731) );
  INV_X1 U9972 ( .A(n14962), .ZN(n14961) );
  NOR2_X1 U9973 ( .A1(n14913), .A2(n14908), .ZN(n14909) );
  NAND2_X1 U9974 ( .A1(n8296), .A2(n8295), .ZN(n14912) );
  INV_X1 U9975 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10953) );
  INV_X1 U9976 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9471) );
  INV_X1 U9977 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U9978 ( .A1(n9358), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14620) );
  INV_X1 U9979 ( .A(n14616), .ZN(n13921) );
  INV_X1 U9980 ( .A(n14042), .ZN(n14068) );
  INV_X1 U9981 ( .A(n12410), .ZN(n13945) );
  OR2_X1 U9982 ( .A1(n14718), .A2(n8926), .ZN(n14020) );
  OR2_X1 U9983 ( .A1(n14051), .A2(n11352), .ZN(n14489) );
  AOI211_X1 U9984 ( .C1(n14262), .C2(n14274), .A(n14065), .B(n14064), .ZN(
        n14066) );
  OR2_X1 U9985 ( .A1(n14747), .A2(n11334), .ZN(n14739) );
  OR2_X1 U9986 ( .A1(n9244), .A2(n9646), .ZN(n14806) );
  AND3_X1 U9987 ( .A1(n14680), .A2(n14679), .A3(n14678), .ZN(n14687) );
  NAND2_X1 U9988 ( .A1(n8831), .A2(n8797), .ZN(n14749) );
  NAND2_X1 U9989 ( .A1(n8126), .A2(n8112), .ZN(n11338) );
  INV_X1 U9990 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8872) );
  INV_X1 U9991 ( .A(n13268), .ZN(P2_U3947) );
  NOR2_X1 U9992 ( .A1(n8575), .A2(n8825), .ZN(P1_U4016) );
  NOR2_X1 U9993 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7706) );
  NOR2_X1 U9994 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7709) );
  NOR2_X1 U9995 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7711) );
  INV_X2 U9996 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8281) );
  XNOR2_X2 U9997 ( .A(n7714), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U9998 ( .A1(n8255), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7727) );
  INV_X1 U9999 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n7717) );
  OR2_X1 U10000 ( .A1(n8256), .A2(n7717), .ZN(n7726) );
  NAND2_X1 U10001 ( .A1(n7907), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10002 ( .A1(n7937), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10003 ( .A1(n8005), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8024) );
  INV_X1 U10004 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8023) );
  INV_X1 U10005 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8095) );
  INV_X1 U10006 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8116) );
  INV_X1 U10007 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13156) );
  INV_X1 U10008 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13220) );
  NAND2_X1 U10009 ( .A1(n8187), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8186) );
  INV_X1 U10010 ( .A(n8212), .ZN(n7719) );
  NAND2_X1 U10011 ( .A1(n7719), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8214) );
  INV_X1 U10012 ( .A(n8214), .ZN(n7720) );
  INV_X1 U10013 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15161) );
  NAND2_X1 U10014 ( .A1(n8214), .A2(n15161), .ZN(n7721) );
  NAND2_X1 U10015 ( .A1(n8240), .A2(n7721), .ZN(n13437) );
  OR2_X1 U10016 ( .A1(n8257), .A2(n13437), .ZN(n7725) );
  INV_X1 U10017 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7723) );
  OR2_X1 U10018 ( .A1(n6943), .A2(n7723), .ZN(n7724) );
  NAND4_X1 U10019 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n7724), .ZN(n13243) );
  INV_X1 U10020 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8876) );
  AND2_X1 U10021 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7729) );
  NAND2_X1 U10022 ( .A1(n9161), .A2(n7729), .ZN(n8822) );
  AND2_X1 U10023 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U10024 ( .A1(n6538), .A2(n7730), .ZN(n7837) );
  NAND2_X1 U10025 ( .A1(n8822), .A2(n7837), .ZN(n7830) );
  INV_X1 U10026 ( .A(SI_1_), .ZN(n9247) );
  NOR2_X1 U10027 ( .A1(n7731), .A2(n9247), .ZN(n7732) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n6538), .Z(n7733) );
  XNOR2_X1 U10029 ( .A(n7733), .B(SI_2_), .ZN(n7849) );
  NAND2_X1 U10030 ( .A1(n7733), .A2(SI_2_), .ZN(n7734) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6538), .Z(n7735) );
  INV_X1 U10032 ( .A(SI_3_), .ZN(n8499) );
  XNOR2_X1 U10033 ( .A(n7735), .B(n8499), .ZN(n7864) );
  NAND2_X1 U10034 ( .A1(n7735), .A2(SI_3_), .ZN(n7736) );
  NAND2_X1 U10035 ( .A1(n7737), .A2(n7736), .ZN(n7876) );
  XNOR2_X1 U10036 ( .A(n7739), .B(SI_4_), .ZN(n7875) );
  INV_X1 U10037 ( .A(n7875), .ZN(n7738) );
  NAND2_X1 U10038 ( .A1(n7876), .A2(n7738), .ZN(n7741) );
  NAND2_X1 U10039 ( .A1(n7739), .A2(SI_4_), .ZN(n7740) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6536), .Z(n7743) );
  XNOR2_X1 U10041 ( .A(n7743), .B(SI_5_), .ZN(n7888) );
  INV_X1 U10042 ( .A(n7888), .ZN(n7742) );
  NAND2_X1 U10043 ( .A1(n7889), .A2(n7742), .ZN(n7745) );
  NAND2_X1 U10044 ( .A1(n7743), .A2(SI_5_), .ZN(n7744) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6536), .Z(n7747) );
  XNOR2_X1 U10046 ( .A(n7747), .B(SI_6_), .ZN(n7897) );
  INV_X1 U10047 ( .A(n7897), .ZN(n7746) );
  NAND2_X1 U10048 ( .A1(n7747), .A2(SI_6_), .ZN(n7914) );
  MUX2_X1 U10049 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6536), .Z(n7749) );
  NAND2_X1 U10050 ( .A1(n7749), .A2(SI_7_), .ZN(n7748) );
  AND2_X1 U10051 ( .A1(n7914), .A2(n7748), .ZN(n7752) );
  INV_X1 U10052 ( .A(n7748), .ZN(n7751) );
  XNOR2_X1 U10053 ( .A(n7749), .B(SI_7_), .ZN(n7916) );
  INV_X1 U10054 ( .A(n7916), .ZN(n7750) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6536), .Z(n7754) );
  XNOR2_X1 U10056 ( .A(n7754), .B(SI_8_), .ZN(n7930) );
  INV_X1 U10057 ( .A(n7930), .ZN(n7753) );
  NAND2_X1 U10058 ( .A1(n7754), .A2(SI_8_), .ZN(n7755) );
  MUX2_X1 U10059 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6536), .Z(n7757) );
  XNOR2_X1 U10060 ( .A(n7757), .B(SI_9_), .ZN(n7944) );
  INV_X1 U10061 ( .A(n7944), .ZN(n7756) );
  NAND2_X1 U10062 ( .A1(n7757), .A2(SI_9_), .ZN(n7960) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6536), .Z(n7760) );
  NAND2_X1 U10064 ( .A1(n7760), .A2(SI_10_), .ZN(n7759) );
  AND2_X1 U10065 ( .A1(n7960), .A2(n7759), .ZN(n7758) );
  INV_X1 U10066 ( .A(n7759), .ZN(n7762) );
  XNOR2_X1 U10067 ( .A(n7760), .B(SI_10_), .ZN(n7962) );
  INV_X1 U10068 ( .A(n7962), .ZN(n7761) );
  MUX2_X1 U10069 ( .A(n8633), .B(n8629), .S(n6536), .Z(n7764) );
  INV_X1 U10070 ( .A(SI_11_), .ZN(n8478) );
  NAND2_X1 U10071 ( .A1(n7764), .A2(n8478), .ZN(n7980) );
  INV_X1 U10072 ( .A(n7764), .ZN(n7765) );
  NAND2_X1 U10073 ( .A1(n7765), .A2(SI_11_), .ZN(n7979) );
  INV_X1 U10074 ( .A(n7979), .ZN(n7766) );
  MUX2_X1 U10075 ( .A(n8588), .B(n8736), .S(n6536), .Z(n7767) );
  NAND2_X1 U10076 ( .A1(n7767), .A2(n10712), .ZN(n7770) );
  INV_X1 U10077 ( .A(n7767), .ZN(n7768) );
  NAND2_X1 U10078 ( .A1(n7768), .A2(SI_12_), .ZN(n7769) );
  MUX2_X1 U10079 ( .A(n8872), .B(n8874), .S(n6535), .Z(n7771) );
  INV_X1 U10080 ( .A(n7771), .ZN(n7772) );
  NAND2_X1 U10081 ( .A1(n7772), .A2(SI_13_), .ZN(n7773) );
  MUX2_X1 U10082 ( .A(n9313), .B(n9315), .S(n6536), .Z(n7778) );
  MUX2_X1 U10083 ( .A(n9417), .B(n9419), .S(n6535), .Z(n7775) );
  INV_X1 U10084 ( .A(n7775), .ZN(n7776) );
  NAND2_X1 U10085 ( .A1(n7776), .A2(SI_15_), .ZN(n7777) );
  NAND2_X1 U10086 ( .A1(n7781), .A2(n7777), .ZN(n8047) );
  NOR2_X1 U10087 ( .A1(n7778), .A2(n6716), .ZN(n7779) );
  MUX2_X1 U10088 ( .A(n9284), .B(n9286), .S(n6536), .Z(n7782) );
  INV_X1 U10089 ( .A(n7782), .ZN(n7783) );
  NAND2_X1 U10090 ( .A1(n7783), .A2(SI_16_), .ZN(n7784) );
  MUX2_X1 U10091 ( .A(n9476), .B(n9471), .S(n6535), .Z(n8084) );
  NAND2_X1 U10092 ( .A1(n8084), .A2(n9039), .ZN(n8106) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6535), .Z(n8108) );
  OAI21_X1 U10094 ( .B1(n8108), .B2(SI_18_), .A(SI_19_), .ZN(n7787) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6536), .Z(n8127) );
  INV_X1 U10096 ( .A(n8127), .ZN(n7786) );
  NOR2_X1 U10097 ( .A1(SI_18_), .A2(SI_19_), .ZN(n7785) );
  INV_X1 U10098 ( .A(n8108), .ZN(n8110) );
  INV_X1 U10099 ( .A(n7789), .ZN(n7791) );
  INV_X1 U10100 ( .A(n8084), .ZN(n7790) );
  NAND2_X1 U10101 ( .A1(n7790), .A2(SI_17_), .ZN(n8104) );
  INV_X1 U10102 ( .A(n7792), .ZN(n7794) );
  AOI22_X1 U10103 ( .A1(SI_18_), .A2(n8108), .B1(n8127), .B2(SI_19_), .ZN(
        n7793) );
  INV_X1 U10104 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9719) );
  MUX2_X1 U10105 ( .A(n15251), .B(n9719), .S(n6535), .Z(n8141) );
  MUX2_X1 U10106 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6535), .Z(n7799) );
  OAI21_X1 U10107 ( .B1(SI_21_), .B2(n7799), .A(n7801), .ZN(n7800) );
  INV_X1 U10108 ( .A(n7800), .ZN(n8155) );
  INV_X1 U10109 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7804) );
  MUX2_X1 U10110 ( .A(n7804), .B(n10419), .S(n6535), .Z(n8168) );
  MUX2_X1 U10111 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6536), .Z(n7806) );
  INV_X1 U10112 ( .A(SI_23_), .ZN(n11222) );
  INV_X1 U10113 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11801) );
  MUX2_X1 U10114 ( .A(n11801), .B(n10953), .S(n6535), .Z(n8194) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6535), .Z(n7810) );
  XNOR2_X1 U10116 ( .A(n7810), .B(SI_25_), .ZN(n8206) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n6535), .Z(n7811) );
  NAND2_X1 U10118 ( .A1(n7811), .A2(SI_26_), .ZN(n8222) );
  OAI21_X1 U10119 ( .B1(SI_26_), .B2(n7811), .A(n8222), .ZN(n7812) );
  NAND2_X1 U10120 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  INV_X1 U10121 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7817) );
  XNOR2_X2 U10122 ( .A(n7818), .B(n7817), .ZN(n13761) );
  NAND2_X1 U10123 ( .A1(n13763), .A2(n12230), .ZN(n7820) );
  INV_X1 U10125 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13765) );
  OR2_X1 U10126 ( .A1(n7832), .A2(n13765), .ZN(n7819) );
  INV_X1 U10127 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7821) );
  INV_X1 U10128 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13270) );
  OR2_X1 U10129 ( .A1(n7855), .A2(n13270), .ZN(n7824) );
  INV_X1 U10130 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U10131 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7827) );
  MUX2_X1 U10132 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7827), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7829) );
  INV_X1 U10133 ( .A(n7844), .ZN(n7828) );
  NAND2_X1 U10134 ( .A1(n7829), .A2(n7828), .ZN(n13271) );
  OAI211_X2 U10135 ( .C1(n8899), .C2(n13271), .A(n7834), .B(n7833), .ZN(n12053) );
  NAND2_X1 U10136 ( .A1(n13269), .A2(n9451), .ZN(n7835) );
  INV_X1 U10137 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9538) );
  INV_X1 U10138 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U10139 ( .A1(n6536), .A2(SI_0_), .ZN(n7836) );
  INV_X1 U10140 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10141 ( .A1(n7836), .A2(n8437), .ZN(n7838) );
  NAND2_X1 U10142 ( .A1(n7838), .A2(n7837), .ZN(n13769) );
  MUX2_X1 U10143 ( .A(n7014), .B(n13769), .S(n8899), .Z(n12041) );
  INV_X1 U10144 ( .A(n12041), .ZN(n9467) );
  INV_X2 U10145 ( .A(n7857), .ZN(n12218) );
  NAND2_X1 U10146 ( .A1(n12218), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7843) );
  INV_X1 U10147 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14827) );
  OR2_X1 U10148 ( .A1(n7855), .A2(n14827), .ZN(n7842) );
  INV_X1 U10149 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7839) );
  INV_X1 U10150 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10166) );
  INV_X1 U10151 ( .A(n7845), .ZN(n7847) );
  NAND2_X1 U10152 ( .A1(n7847), .A2(n7846), .ZN(n8906) );
  XNOR2_X1 U10153 ( .A(n7848), .B(n7849), .ZN(n9018) );
  OR2_X1 U10154 ( .A1(n8171), .A2(n9018), .ZN(n7851) );
  OR2_X1 U10155 ( .A1(n7832), .A2(n8556), .ZN(n7850) );
  NAND2_X1 U10156 ( .A1(n10161), .A2(n8312), .ZN(n7854) );
  OR2_X1 U10157 ( .A1(n13267), .A2(n7852), .ZN(n7853) );
  NAND2_X1 U10158 ( .A1(n7854), .A2(n7853), .ZN(n14887) );
  NAND2_X1 U10159 ( .A1(n8361), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7861) );
  OR2_X1 U10160 ( .A1(n7855), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7860) );
  INV_X1 U10161 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7856) );
  OR2_X1 U10162 ( .A1(n7857), .A2(n7856), .ZN(n7859) );
  INV_X1 U10163 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8907) );
  OR2_X1 U10164 ( .A1(n6525), .A2(n8907), .ZN(n7858) );
  NAND4_X1 U10165 ( .A1(n7861), .A2(n7860), .A3(n7859), .A4(n7858), .ZN(n13266) );
  NAND2_X1 U10166 ( .A1(n7846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7863) );
  INV_X1 U10167 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U10168 ( .A(n7863), .B(n7862), .ZN(n8908) );
  OR2_X1 U10169 ( .A1(n8171), .A2(n9348), .ZN(n7866) );
  OR2_X1 U10170 ( .A1(n7832), .A2(n8559), .ZN(n7865) );
  OAI211_X1 U10171 ( .C1(n8899), .C2(n8908), .A(n7866), .B(n7865), .ZN(n9565)
         );
  INV_X1 U10172 ( .A(n14901), .ZN(n14930) );
  OR2_X1 U10173 ( .A1(n13266), .A2(n14930), .ZN(n8314) );
  NAND2_X1 U10174 ( .A1(n13266), .A2(n14930), .ZN(n7867) );
  NAND2_X1 U10175 ( .A1(n8314), .A2(n7867), .ZN(n14886) );
  NAND2_X1 U10176 ( .A1(n14887), .A2(n14886), .ZN(n7869) );
  OR2_X1 U10177 ( .A1(n13266), .A2(n14901), .ZN(n7868) );
  NAND2_X1 U10178 ( .A1(n7869), .A2(n7868), .ZN(n10173) );
  NAND2_X1 U10179 ( .A1(n6893), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7873) );
  INV_X1 U10180 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10179) );
  OR2_X1 U10181 ( .A1(n6525), .A2(n10179), .ZN(n7872) );
  XNOR2_X1 U10182 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10181) );
  OR2_X1 U10183 ( .A1(n7855), .A2(n10181), .ZN(n7871) );
  OR2_X1 U10184 ( .A1(n7857), .A2(n14967), .ZN(n7870) );
  NAND4_X1 U10185 ( .A1(n7873), .A2(n7872), .A3(n7871), .A4(n7870), .ZN(n13265) );
  OR2_X1 U10186 ( .A1(n7846), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10187 ( .A1(n7890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7874) );
  XNOR2_X1 U10188 ( .A(n7874), .B(n7891), .ZN(n8909) );
  XNOR2_X1 U10189 ( .A(n7876), .B(n7875), .ZN(n9512) );
  NAND2_X1 U10190 ( .A1(n9512), .A2(n12230), .ZN(n7878) );
  OR2_X1 U10191 ( .A1(n7832), .A2(n8553), .ZN(n7877) );
  XNOR2_X1 U10192 ( .A(n13265), .B(n10182), .ZN(n12266) );
  NAND2_X1 U10193 ( .A1(n10173), .A2(n12266), .ZN(n7880) );
  OR2_X1 U10194 ( .A1(n13265), .A2(n14936), .ZN(n7879) );
  INV_X1 U10195 ( .A(n8257), .ZN(n8072) );
  AOI21_X1 U10196 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7881) );
  NOR2_X1 U10197 ( .A1(n7881), .A2(n7907), .ZN(n13173) );
  NAND2_X1 U10198 ( .A1(n8072), .A2(n13173), .ZN(n7887) );
  INV_X1 U10199 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8910) );
  OR2_X1 U10200 ( .A1(n6525), .A2(n8910), .ZN(n7886) );
  INV_X1 U10201 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10202 ( .A1(n8256), .A2(n7882), .ZN(n7885) );
  INV_X1 U10203 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7883) );
  OR2_X1 U10204 ( .A1(n6943), .A2(n7883), .ZN(n7884) );
  NAND4_X1 U10205 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n13264) );
  XNOR2_X1 U10206 ( .A(n7889), .B(n7888), .ZN(n9741) );
  NAND2_X1 U10207 ( .A1(n9741), .A2(n12230), .ZN(n7895) );
  INV_X1 U10208 ( .A(n7890), .ZN(n7892) );
  NAND2_X1 U10209 ( .A1(n7892), .A2(n7891), .ZN(n7899) );
  NAND2_X1 U10210 ( .A1(n7899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7893) );
  XNOR2_X1 U10211 ( .A(n7893), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9007) );
  AOI22_X1 U10212 ( .A1(n8133), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8132), .B2(
        n9007), .ZN(n7894) );
  NAND2_X1 U10213 ( .A1(n7895), .A2(n7894), .ZN(n13184) );
  NAND2_X1 U10214 ( .A1(n13264), .A2(n13184), .ZN(n7896) );
  XNOR2_X1 U10215 ( .A(n7898), .B(n7897), .ZN(n9767) );
  NAND2_X1 U10216 ( .A1(n9767), .A2(n12230), .ZN(n7905) );
  INV_X1 U10217 ( .A(n7899), .ZN(n7900) );
  INV_X1 U10218 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U10219 ( .A1(n7900), .A2(n15415), .ZN(n7902) );
  NAND2_X1 U10220 ( .A1(n7902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7901) );
  MUX2_X1 U10221 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7901), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n7903) );
  AOI22_X1 U10222 ( .A1(n8133), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8132), .B2(
        n8973), .ZN(n7904) );
  NAND2_X1 U10223 ( .A1(n7905), .A2(n7904), .ZN(n12084) );
  NAND2_X1 U10224 ( .A1(n8255), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7911) );
  INV_X1 U10225 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7906) );
  OR2_X1 U10226 ( .A1(n8256), .A2(n7906), .ZN(n7910) );
  OAI21_X1 U10227 ( .B1(n7907), .B2(P2_REG3_REG_6__SCAN_IN), .A(n7923), .ZN(
        n10194) );
  OR2_X1 U10228 ( .A1(n8257), .A2(n10194), .ZN(n7909) );
  INV_X1 U10229 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8896) );
  OR2_X1 U10230 ( .A1(n7857), .A2(n8896), .ZN(n7908) );
  NAND4_X1 U10231 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), .ZN(n13263) );
  XNOR2_X1 U10232 ( .A(n12084), .B(n13263), .ZN(n12269) );
  OR2_X1 U10233 ( .A1(n12084), .A2(n13263), .ZN(n7912) );
  NAND2_X1 U10234 ( .A1(n7915), .A2(n7914), .ZN(n7917) );
  XNOR2_X1 U10235 ( .A(n7917), .B(n7916), .ZN(n9928) );
  NAND2_X1 U10236 ( .A1(n9928), .A2(n12230), .ZN(n7920) );
  NAND2_X1 U10237 ( .A1(n7932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7918) );
  XNOR2_X1 U10238 ( .A(n7918), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9634) );
  AOI22_X1 U10239 ( .A1(n8133), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8132), .B2(
        n9634), .ZN(n7919) );
  NAND2_X1 U10240 ( .A1(n8361), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7928) );
  INV_X1 U10241 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7921) );
  OR2_X1 U10242 ( .A1(n6525), .A2(n7921), .ZN(n7927) );
  AND2_X1 U10243 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  OR2_X1 U10244 ( .A1(n7924), .A2(n7937), .ZN(n9811) );
  OR2_X1 U10245 ( .A1(n8257), .A2(n9811), .ZN(n7926) );
  INV_X1 U10246 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8974) );
  OR2_X1 U10247 ( .A1(n6943), .A2(n8974), .ZN(n7925) );
  NAND4_X1 U10248 ( .A1(n7928), .A2(n7927), .A3(n7926), .A4(n7925), .ZN(n13262) );
  XNOR2_X1 U10249 ( .A(n12091), .B(n13262), .ZN(n12270) );
  INV_X1 U10250 ( .A(n12270), .ZN(n10300) );
  OR2_X1 U10251 ( .A1(n12091), .A2(n13262), .ZN(n7929) );
  XNOR2_X1 U10252 ( .A(n7931), .B(n7930), .ZN(n10018) );
  NAND2_X1 U10253 ( .A1(n10018), .A2(n12230), .ZN(n7935) );
  NAND2_X1 U10254 ( .A1(n7933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7947) );
  XNOR2_X1 U10255 ( .A(n7947), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9635) );
  AOI22_X1 U10256 ( .A1(n8133), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8132), .B2(
        n9635), .ZN(n7934) );
  NAND2_X1 U10257 ( .A1(n7935), .A2(n7934), .ZN(n14952) );
  NAND2_X1 U10258 ( .A1(n8255), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7942) );
  INV_X1 U10259 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7936) );
  OR2_X1 U10260 ( .A1(n8256), .A2(n7936), .ZN(n7941) );
  OR2_X1 U10261 ( .A1(n7937), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10262 ( .A1(n7952), .A2(n7938), .ZN(n10411) );
  OR2_X1 U10263 ( .A1(n8257), .A2(n10411), .ZN(n7940) );
  INV_X1 U10264 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9629) );
  OR2_X1 U10265 ( .A1(n6943), .A2(n9629), .ZN(n7939) );
  NAND4_X1 U10266 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n13261) );
  XNOR2_X1 U10267 ( .A(n14952), .B(n12099), .ZN(n12273) );
  NAND2_X1 U10268 ( .A1(n14952), .A2(n13261), .ZN(n7943) );
  XNOR2_X1 U10269 ( .A(n7945), .B(n7944), .ZN(n10024) );
  NAND2_X1 U10270 ( .A1(n10024), .A2(n12230), .ZN(n7951) );
  INV_X1 U10271 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10272 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  NAND2_X1 U10273 ( .A1(n7948), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7949) );
  XNOR2_X1 U10274 ( .A(n7949), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9636) );
  AOI22_X1 U10275 ( .A1(n8133), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8132), .B2(
        n9636), .ZN(n7950) );
  NAND2_X1 U10276 ( .A1(n6893), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7957) );
  INV_X1 U10277 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10470) );
  OR2_X1 U10278 ( .A1(n6525), .A2(n10470), .ZN(n7956) );
  NAND2_X1 U10279 ( .A1(n7952), .A2(n11802), .ZN(n7953) );
  NAND2_X1 U10280 ( .A1(n7969), .A2(n7953), .ZN(n11805) );
  OR2_X1 U10281 ( .A1(n8257), .A2(n11805), .ZN(n7955) );
  INV_X1 U10282 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9630) );
  OR2_X1 U10283 ( .A1(n6943), .A2(n9630), .ZN(n7954) );
  NAND4_X1 U10284 ( .A1(n7957), .A2(n7956), .A3(n7955), .A4(n7954), .ZN(n13260) );
  XNOR2_X1 U10285 ( .A(n12103), .B(n13260), .ZN(n12275) );
  NAND2_X1 U10286 ( .A1(n12103), .A2(n13260), .ZN(n7958) );
  NAND2_X1 U10287 ( .A1(n7961), .A2(n7960), .ZN(n7963) );
  XNOR2_X1 U10288 ( .A(n7963), .B(n7962), .ZN(n10215) );
  NAND2_X1 U10289 ( .A1(n10215), .A2(n12230), .ZN(n7968) );
  NAND2_X1 U10290 ( .A1(n7964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7965) );
  MUX2_X1 U10291 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7965), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n7966) );
  NOR2_X1 U10292 ( .A1(n7964), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8050) );
  INV_X1 U10293 ( .A(n8050), .ZN(n7983) );
  NAND2_X1 U10294 ( .A1(n7966), .A2(n7983), .ZN(n9637) );
  INV_X1 U10295 ( .A(n9637), .ZN(n9847) );
  AOI22_X1 U10296 ( .A1(n8133), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8132), 
        .B2(n9847), .ZN(n7967) );
  NAND2_X1 U10297 ( .A1(n8361), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7974) );
  INV_X1 U10298 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n13597) );
  OR2_X1 U10299 ( .A1(n6525), .A2(n13597), .ZN(n7973) );
  NAND2_X1 U10300 ( .A1(n7969), .A2(n15377), .ZN(n7970) );
  NAND2_X1 U10301 ( .A1(n7989), .A2(n7970), .ZN(n13596) );
  OR2_X1 U10302 ( .A1(n8257), .A2(n13596), .ZN(n7972) );
  INV_X1 U10303 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9627) );
  OR2_X1 U10304 ( .A1(n6943), .A2(n9627), .ZN(n7971) );
  NAND4_X1 U10305 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(n13259) );
  XNOR2_X1 U10306 ( .A(n13601), .B(n13259), .ZN(n12278) );
  INV_X1 U10307 ( .A(n12278), .ZN(n7975) );
  NAND2_X1 U10308 ( .A1(n13601), .A2(n13259), .ZN(n7976) );
  NAND2_X1 U10309 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U10310 ( .A1(n10345), .A2(n12230), .ZN(n7988) );
  NAND2_X1 U10311 ( .A1(n7983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7984) );
  MUX2_X1 U10312 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7984), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n7986) );
  INV_X1 U10313 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10314 ( .A1(n8050), .A2(n7985), .ZN(n8001) );
  NAND2_X1 U10315 ( .A1(n7986), .A2(n8001), .ZN(n11075) );
  INV_X1 U10316 ( .A(n11075), .ZN(n11066) );
  AOI22_X1 U10317 ( .A1(n8133), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8132), 
        .B2(n11066), .ZN(n7987) );
  NAND2_X2 U10318 ( .A1(n7988), .A2(n7987), .ZN(n12115) );
  NAND2_X1 U10319 ( .A1(n8255), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7993) );
  INV_X1 U10320 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15413) );
  OR2_X1 U10321 ( .A1(n8256), .A2(n15413), .ZN(n7992) );
  OR2_X1 U10322 ( .A1(n7698), .A2(n8005), .ZN(n10777) );
  OR2_X1 U10323 ( .A1(n8257), .A2(n10777), .ZN(n7991) );
  INV_X1 U10324 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15381) );
  OR2_X1 U10325 ( .A1(n6943), .A2(n15381), .ZN(n7990) );
  NAND4_X1 U10326 ( .A1(n7993), .A2(n7992), .A3(n7991), .A4(n7990), .ZN(n13258) );
  OR2_X1 U10327 ( .A1(n12115), .A2(n13258), .ZN(n7994) );
  NAND2_X1 U10328 ( .A1(n7995), .A2(n7994), .ZN(n10814) );
  OR2_X1 U10329 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  NAND2_X1 U10330 ( .A1(n7999), .A2(n7998), .ZN(n10594) );
  NAND2_X1 U10331 ( .A1(n10594), .A2(n12230), .ZN(n8004) );
  NAND2_X1 U10332 ( .A1(n8001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8000) );
  MUX2_X1 U10333 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8000), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8002) );
  AOI22_X1 U10334 ( .A1(n8133), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8132), 
        .B2(n11076), .ZN(n8003) );
  NAND2_X2 U10335 ( .A1(n8004), .A2(n8003), .ZN(n13587) );
  NAND2_X1 U10336 ( .A1(n8361), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8010) );
  OR2_X1 U10337 ( .A1(n8005), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10338 ( .A1(n8024), .A2(n8006), .ZN(n13584) );
  OR2_X1 U10339 ( .A1(n8257), .A2(n13584), .ZN(n8009) );
  INV_X1 U10340 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11067) );
  OR2_X1 U10341 ( .A1(n6943), .A2(n11067), .ZN(n8008) );
  INV_X1 U10342 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13585) );
  OR2_X1 U10343 ( .A1(n6525), .A2(n13585), .ZN(n8007) );
  NAND4_X1 U10344 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n13257) );
  INV_X1 U10345 ( .A(n13257), .ZN(n8011) );
  OR2_X1 U10346 ( .A1(n13587), .A2(n8011), .ZN(n10804) );
  NAND2_X1 U10347 ( .A1(n13587), .A2(n8011), .ZN(n8012) );
  NAND2_X1 U10348 ( .A1(n10804), .A2(n8012), .ZN(n12277) );
  NAND2_X1 U10349 ( .A1(n10814), .A2(n12277), .ZN(n8014) );
  OR2_X1 U10350 ( .A1(n13587), .A2(n13257), .ZN(n8013) );
  OR2_X1 U10351 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  NAND2_X1 U10352 ( .A1(n8018), .A2(n8017), .ZN(n10598) );
  NAND2_X1 U10353 ( .A1(n10598), .A2(n12230), .ZN(n8022) );
  NAND2_X1 U10354 ( .A1(n8032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8020) );
  INV_X1 U10355 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8019) );
  XNOR2_X1 U10356 ( .A(n8020), .B(n8019), .ZN(n11077) );
  INV_X1 U10357 ( .A(n11077), .ZN(n14864) );
  AOI22_X1 U10358 ( .A1(n8133), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8132), 
        .B2(n14864), .ZN(n8021) );
  NAND2_X1 U10359 ( .A1(n12218), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8029) );
  INV_X1 U10360 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15398) );
  OR2_X1 U10361 ( .A1(n8256), .A2(n15398), .ZN(n8028) );
  NAND2_X1 U10362 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  NAND2_X1 U10363 ( .A1(n8036), .A2(n8025), .ZN(n14822) );
  OR2_X1 U10364 ( .A1(n8257), .A2(n14822), .ZN(n8027) );
  INV_X1 U10365 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11073) );
  OR2_X1 U10366 ( .A1(n6525), .A2(n11073), .ZN(n8026) );
  NAND4_X1 U10367 ( .A1(n8029), .A2(n8028), .A3(n8027), .A4(n8026), .ZN(n13256) );
  NOR2_X1 U10368 ( .A1(n14819), .A2(n13256), .ZN(n8030) );
  INV_X1 U10369 ( .A(n13256), .ZN(n10567) );
  NAND2_X1 U10370 ( .A1(n10732), .A2(n12230), .ZN(n8035) );
  OAI21_X1 U10371 ( .B1(n8032), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U10372 ( .A(n8033), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U10373 ( .A1(n8133), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8132), 
        .B2(n11078), .ZN(n8034) );
  AND2_X1 U10374 ( .A1(n8036), .A2(n13312), .ZN(n8037) );
  OR2_X1 U10375 ( .A1(n8037), .A2(n8057), .ZN(n10889) );
  OR2_X1 U10376 ( .A1(n8257), .A2(n10889), .ZN(n8041) );
  INV_X1 U10377 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11058) );
  OR2_X1 U10378 ( .A1(n8256), .A2(n11058), .ZN(n8040) );
  INV_X1 U10379 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10890) );
  OR2_X1 U10380 ( .A1(n6525), .A2(n10890), .ZN(n8039) );
  INV_X1 U10381 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15380) );
  OR2_X1 U10382 ( .A1(n6943), .A2(n15380), .ZN(n8038) );
  NAND4_X1 U10383 ( .A1(n8041), .A2(n8040), .A3(n8039), .A4(n8038), .ZN(n13255) );
  XNOR2_X1 U10384 ( .A(n12139), .B(n13255), .ZN(n12284) );
  INV_X1 U10385 ( .A(n12284), .ZN(n8042) );
  NAND2_X1 U10386 ( .A1(n10883), .A2(n8042), .ZN(n8044) );
  NAND2_X1 U10387 ( .A1(n12139), .A2(n13255), .ZN(n8043) );
  NAND2_X1 U10388 ( .A1(n8044), .A2(n8043), .ZN(n10991) );
  INV_X1 U10389 ( .A(n10991), .ZN(n8063) );
  INV_X1 U10390 ( .A(n8047), .ZN(n8048) );
  NAND2_X1 U10391 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U10392 ( .A1(n8051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8052) );
  XNOR2_X1 U10393 ( .A(n8052), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U10394 ( .A1(n8133), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8132), 
        .B2(n13328), .ZN(n8053) );
  INV_X1 U10395 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15332) );
  INV_X1 U10396 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8055) );
  OR2_X1 U10397 ( .A1(n8256), .A2(n8055), .ZN(n8056) );
  OAI21_X1 U10398 ( .B1(n6525), .B2(n15332), .A(n8056), .ZN(n8061) );
  NOR2_X1 U10399 ( .A1(n8057), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8058) );
  OR2_X1 U10400 ( .A1(n8070), .A2(n8058), .ZN(n12387) );
  INV_X1 U10401 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11069) );
  OR2_X1 U10402 ( .A1(n6943), .A2(n11069), .ZN(n8059) );
  OAI21_X1 U10403 ( .B1(n8257), .B2(n12387), .A(n8059), .ZN(n8060) );
  XNOR2_X1 U10404 ( .A(n13696), .B(n13254), .ZN(n12285) );
  INV_X1 U10405 ( .A(n12285), .ZN(n8062) );
  OR2_X1 U10406 ( .A1(n13696), .A2(n13254), .ZN(n8064) );
  XNOR2_X1 U10407 ( .A(n8066), .B(n8065), .ZN(n11447) );
  NAND2_X1 U10408 ( .A1(n11447), .A2(n12230), .ZN(n8069) );
  OR2_X1 U10409 ( .A1(n8087), .A2(n7486), .ZN(n8067) );
  XNOR2_X1 U10410 ( .A(n8067), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U10411 ( .A1(n8133), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8132), 
        .B2(n13345), .ZN(n8068) );
  OR2_X1 U10412 ( .A1(n8070), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8071) );
  AND2_X1 U10413 ( .A1(n8096), .A2(n8071), .ZN(n11120) );
  NAND2_X1 U10414 ( .A1(n8072), .A2(n11120), .ZN(n8079) );
  INV_X1 U10415 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8073) );
  OR2_X1 U10416 ( .A1(n8256), .A2(n8073), .ZN(n8078) );
  INV_X1 U10417 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8074) );
  OR2_X1 U10418 ( .A1(n6943), .A2(n8074), .ZN(n8077) );
  INV_X1 U10419 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8075) );
  OR2_X1 U10420 ( .A1(n6525), .A2(n8075), .ZN(n8076) );
  NAND4_X1 U10421 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n13253) );
  INV_X1 U10422 ( .A(n13253), .ZN(n8080) );
  OR2_X1 U10423 ( .A1(n13743), .A2(n8080), .ZN(n8336) );
  NAND2_X1 U10424 ( .A1(n13743), .A2(n8080), .ZN(n8081) );
  NAND2_X1 U10425 ( .A1(n8336), .A2(n8081), .ZN(n12283) );
  INV_X1 U10426 ( .A(n12283), .ZN(n11094) );
  NAND2_X1 U10427 ( .A1(n8083), .A2(n8082), .ZN(n8105) );
  XNOR2_X1 U10428 ( .A(n8084), .B(SI_17_), .ZN(n8085) );
  XNOR2_X1 U10429 ( .A(n8105), .B(n8085), .ZN(n11453) );
  NAND2_X1 U10430 ( .A1(n11453), .A2(n12230), .ZN(n8094) );
  INV_X1 U10431 ( .A(n8091), .ZN(n8088) );
  NAND2_X1 U10432 ( .A1(n8088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8089) );
  MUX2_X1 U10433 ( .A(n8089), .B(P2_IR_REG_31__SCAN_IN), .S(n8090), .Z(n8092)
         );
  NAND2_X1 U10434 ( .A1(n8092), .A2(n8130), .ZN(n13364) );
  INV_X1 U10435 ( .A(n13364), .ZN(n13346) );
  AOI22_X1 U10436 ( .A1(n8133), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8132), 
        .B2(n13346), .ZN(n8093) );
  NAND2_X1 U10437 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U10438 ( .A1(n8117), .A2(n8097), .ZN(n13574) );
  NAND2_X1 U10439 ( .A1(n12218), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8098) );
  OAI21_X1 U10440 ( .B1(n13574), .B2(n8257), .A(n8098), .ZN(n8101) );
  INV_X1 U10441 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U10442 ( .A1(n8361), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8099) );
  OAI21_X1 U10443 ( .B1(n13575), .B2(n6525), .A(n8099), .ZN(n8100) );
  XNOR2_X1 U10444 ( .A(n13739), .B(n13252), .ZN(n12287) );
  NAND2_X1 U10445 ( .A1(n13566), .A2(n13567), .ZN(n8103) );
  NAND2_X1 U10446 ( .A1(n13739), .A2(n13252), .ZN(n8102) );
  NAND2_X1 U10447 ( .A1(n8103), .A2(n8102), .ZN(n13553) );
  INV_X1 U10448 ( .A(n13553), .ZN(n8122) );
  NAND2_X1 U10449 ( .A1(n8105), .A2(n8104), .ZN(n8107) );
  NAND2_X1 U10450 ( .A1(n8107), .A2(n8106), .ZN(n8124) );
  NAND2_X1 U10451 ( .A1(n8109), .A2(n8108), .ZN(n8126) );
  INV_X1 U10452 ( .A(n8109), .ZN(n8111) );
  NAND2_X1 U10453 ( .A1(n8111), .A2(n8110), .ZN(n8112) );
  NAND2_X1 U10454 ( .A1(n8130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8113) );
  XNOR2_X1 U10455 ( .A(n8113), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U10456 ( .A1(n8133), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8132), 
        .B2(n13365), .ZN(n8114) );
  AND2_X1 U10457 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  OR2_X1 U10458 ( .A1(n8118), .A2(n8136), .ZN(n13559) );
  AOI22_X1 U10459 ( .A1(n8255), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n6893), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10460 ( .A1(n12218), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8119) );
  OAI211_X1 U10461 ( .C1(n13559), .C2(n8257), .A(n8120), .B(n8119), .ZN(n13251) );
  XNOR2_X1 U10462 ( .A(n13735), .B(n13251), .ZN(n13552) );
  OR2_X1 U10463 ( .A1(n13735), .A2(n13251), .ZN(n8123) );
  INV_X1 U10464 ( .A(SI_18_), .ZN(n15396) );
  OR2_X1 U10465 ( .A1(n8124), .A2(n15396), .ZN(n8125) );
  NAND2_X1 U10466 ( .A1(n8126), .A2(n8125), .ZN(n8129) );
  XNOR2_X1 U10467 ( .A(n8127), .B(SI_19_), .ZN(n8128) );
  NAND2_X1 U10468 ( .A1(n11351), .A2(n12230), .ZN(n8135) );
  NAND2_X1 U10469 ( .A1(n8297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8131) );
  AOI22_X1 U10470 ( .A1(n8133), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6527), 
        .B2(n8132), .ZN(n8134) );
  NAND2_X2 U10471 ( .A1(n8135), .A2(n8134), .ZN(n13672) );
  NOR2_X1 U10472 ( .A1(n8136), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8137) );
  OR2_X1 U10473 ( .A1(n8147), .A2(n8137), .ZN(n13544) );
  AOI22_X1 U10474 ( .A1(n8255), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8361), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n8139) );
  INV_X1 U10475 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13375) );
  OR2_X1 U10476 ( .A1(n6943), .A2(n13375), .ZN(n8138) );
  OAI211_X1 U10477 ( .C1(n13544), .C2(n8257), .A(n8139), .B(n8138), .ZN(n13250) );
  OR2_X1 U10478 ( .A1(n13672), .A2(n13250), .ZN(n8140) );
  NAND2_X1 U10479 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  NAND2_X1 U10480 ( .A1(n8144), .A2(n8143), .ZN(n11482) );
  OR2_X1 U10481 ( .A1(n7832), .A2(n9719), .ZN(n8145) );
  OR2_X1 U10482 ( .A1(n8147), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8148) );
  AND2_X1 U10483 ( .A1(n8161), .A2(n8148), .ZN(n13528) );
  NAND2_X1 U10484 ( .A1(n13528), .A2(n8072), .ZN(n8154) );
  INV_X1 U10485 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10486 ( .A1(n12218), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10487 ( .A1(n6893), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8149) );
  OAI211_X1 U10488 ( .C1(n6525), .C2(n8151), .A(n8150), .B(n8149), .ZN(n8152)
         );
  INV_X1 U10489 ( .A(n8152), .ZN(n8153) );
  NAND2_X1 U10490 ( .A1(n8154), .A2(n8153), .ZN(n13249) );
  INV_X1 U10491 ( .A(n13249), .ZN(n8345) );
  OR2_X1 U10492 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U10493 ( .A1(n8158), .A2(n8157), .ZN(n11497) );
  INV_X1 U10494 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9916) );
  OR2_X1 U10495 ( .A1(n7832), .A2(n9916), .ZN(n8159) );
  NAND2_X1 U10496 ( .A1(n8161), .A2(n13156), .ZN(n8162) );
  NAND2_X1 U10497 ( .A1(n8174), .A2(n8162), .ZN(n13514) );
  OR2_X1 U10498 ( .A1(n13514), .A2(n8257), .ZN(n8167) );
  INV_X1 U10499 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13513) );
  NAND2_X1 U10500 ( .A1(n12218), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10501 ( .A1(n8361), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U10502 ( .C1(n6525), .C2(n13513), .A(n8164), .B(n8163), .ZN(n8165)
         );
  INV_X1 U10503 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U10504 ( .A1(n8167), .A2(n8166), .ZN(n13248) );
  XNOR2_X1 U10505 ( .A(n13512), .B(n13248), .ZN(n13506) );
  NAND2_X1 U10506 ( .A1(n11514), .A2(n8168), .ZN(n8169) );
  NAND2_X1 U10507 ( .A1(n8170), .A2(n8169), .ZN(n10416) );
  OR2_X1 U10508 ( .A1(n7832), .A2(n10419), .ZN(n8172) );
  NAND2_X1 U10509 ( .A1(n8174), .A2(n13220), .ZN(n8176) );
  INV_X1 U10510 ( .A(n8187), .ZN(n8175) );
  NAND2_X1 U10511 ( .A1(n8176), .A2(n8175), .ZN(n13497) );
  OR2_X1 U10512 ( .A1(n13497), .A2(n8257), .ZN(n8181) );
  INV_X1 U10513 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U10514 ( .A1(n6893), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10515 ( .A1(n12218), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8177) );
  OAI211_X1 U10516 ( .C1(n13496), .C2(n6525), .A(n8178), .B(n8177), .ZN(n8179)
         );
  INV_X1 U10517 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U10518 ( .A1(n8181), .A2(n8180), .ZN(n13247) );
  XNOR2_X1 U10519 ( .A(n13653), .B(n13214), .ZN(n13494) );
  NAND2_X1 U10520 ( .A1(n13495), .A2(n13494), .ZN(n13493) );
  NAND2_X1 U10521 ( .A1(n13653), .A2(n13247), .ZN(n8182) );
  XNOR2_X1 U10522 ( .A(n8183), .B(SI_23_), .ZN(n11525) );
  NAND2_X1 U10523 ( .A1(n11525), .A2(n12230), .ZN(n8185) );
  INV_X1 U10524 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n15307) );
  OR2_X1 U10525 ( .A1(n7832), .A2(n15307), .ZN(n8184) );
  NAND2_X1 U10526 ( .A1(n8361), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8192) );
  INV_X1 U10527 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13485) );
  OR2_X1 U10528 ( .A1(n6525), .A2(n13485), .ZN(n8191) );
  OAI21_X1 U10529 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8187), .A(n8186), .ZN(
        n13482) );
  OR2_X1 U10530 ( .A1(n8257), .A2(n13482), .ZN(n8190) );
  INV_X1 U10531 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8188) );
  OR2_X1 U10532 ( .A1(n6943), .A2(n8188), .ZN(n8189) );
  NAND4_X1 U10533 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), .ZN(n13246) );
  NAND2_X1 U10534 ( .A1(n13648), .A2(n13246), .ZN(n12291) );
  INV_X1 U10535 ( .A(n12291), .ZN(n8193) );
  OR2_X1 U10536 ( .A1(n13648), .A2(n13246), .ZN(n12292) );
  NAND2_X1 U10537 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  NAND2_X1 U10538 ( .A1(n11537), .A2(n12230), .ZN(n8199) );
  OR2_X1 U10539 ( .A1(n7832), .A2(n10953), .ZN(n8198) );
  NAND2_X1 U10540 ( .A1(n6893), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8205) );
  INV_X1 U10541 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13468) );
  OR2_X1 U10542 ( .A1(n6525), .A2(n13468), .ZN(n8204) );
  OAI21_X1 U10543 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8200), .A(n8212), .ZN(
        n13467) );
  OR2_X1 U10544 ( .A1(n8257), .A2(n13467), .ZN(n8203) );
  INV_X1 U10545 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8201) );
  OR2_X1 U10546 ( .A1(n6943), .A2(n8201), .ZN(n8202) );
  NAND4_X1 U10547 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n13245) );
  XNOR2_X1 U10548 ( .A(n13643), .B(n13245), .ZN(n13464) );
  NAND2_X1 U10549 ( .A1(n11559), .A2(n12230), .ZN(n8209) );
  INV_X1 U10550 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11062) );
  OR2_X1 U10551 ( .A1(n7832), .A2(n11062), .ZN(n8208) );
  NAND2_X1 U10552 ( .A1(n8361), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8219) );
  INV_X1 U10553 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8210) );
  OR2_X1 U10554 ( .A1(n6525), .A2(n8210), .ZN(n8218) );
  INV_X1 U10555 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10556 ( .A1(n8212), .A2(n8211), .ZN(n8213) );
  NAND2_X1 U10557 ( .A1(n8214), .A2(n8213), .ZN(n13450) );
  OR2_X1 U10558 ( .A1(n8257), .A2(n13450), .ZN(n8217) );
  INV_X1 U10559 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8215) );
  OR2_X1 U10560 ( .A1(n6943), .A2(n8215), .ZN(n8216) );
  NAND4_X1 U10561 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n13244) );
  INV_X1 U10562 ( .A(n13244), .ZN(n13194) );
  XNOR2_X1 U10563 ( .A(n13638), .B(n13194), .ZN(n12296) );
  OR2_X1 U10564 ( .A1(n13638), .A2(n13244), .ZN(n8221) );
  NAND2_X1 U10565 ( .A1(n13454), .A2(n8221), .ZN(n13433) );
  INV_X1 U10566 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14367) );
  INV_X1 U10567 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13762) );
  MUX2_X1 U10568 ( .A(n14367), .B(n13762), .S(n6536), .Z(n8231) );
  XNOR2_X1 U10569 ( .A(n8232), .B(SI_27_), .ZN(n8224) );
  NAND2_X1 U10570 ( .A1(n13760), .A2(n12230), .ZN(n8226) );
  OR2_X1 U10571 ( .A1(n7832), .A2(n13762), .ZN(n8225) );
  NAND2_X1 U10572 ( .A1(n8255), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8230) );
  INV_X1 U10573 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13712) );
  OR2_X1 U10574 ( .A1(n8256), .A2(n13712), .ZN(n8229) );
  INV_X1 U10575 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13128) );
  XNOR2_X1 U10576 ( .A(n8240), .B(n13128), .ZN(n13421) );
  OR2_X1 U10577 ( .A1(n8257), .A2(n13421), .ZN(n8228) );
  INV_X1 U10578 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13629) );
  OR2_X1 U10579 ( .A1(n6943), .A2(n13629), .ZN(n8227) );
  NAND4_X1 U10580 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n13242) );
  INV_X1 U10581 ( .A(n13242), .ZN(n8356) );
  XNOR2_X1 U10582 ( .A(n13424), .B(n8356), .ZN(n12261) );
  INV_X1 U10583 ( .A(SI_27_), .ZN(n12565) );
  NOR2_X1 U10584 ( .A1(n8231), .A2(n12565), .ZN(n8233) );
  INV_X1 U10585 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11750) );
  INV_X1 U10586 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13759) );
  MUX2_X1 U10587 ( .A(n11750), .B(n13759), .S(n6535), .Z(n8235) );
  INV_X1 U10588 ( .A(SI_28_), .ZN(n11303) );
  NAND2_X1 U10589 ( .A1(n8235), .A2(n11303), .ZN(n8251) );
  INV_X1 U10590 ( .A(n8235), .ZN(n8236) );
  NAND2_X1 U10591 ( .A1(n8236), .A2(SI_28_), .ZN(n8237) );
  NAND2_X1 U10592 ( .A1(n13756), .A2(n12230), .ZN(n8239) );
  OR2_X1 U10593 ( .A1(n7832), .A2(n13759), .ZN(n8238) );
  NAND2_X1 U10594 ( .A1(n12218), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8247) );
  INV_X1 U10595 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13410) );
  OR2_X1 U10596 ( .A1(n6525), .A2(n13410), .ZN(n8246) );
  INV_X1 U10597 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15376) );
  OR2_X1 U10598 ( .A1(n8256), .A2(n15376), .ZN(n8245) );
  INV_X1 U10599 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12403) );
  OAI21_X1 U10600 ( .B1(n8240), .B2(n13128), .A(n12403), .ZN(n8243) );
  INV_X1 U10601 ( .A(n8240), .ZN(n8242) );
  AND2_X1 U10602 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8241) );
  NAND2_X1 U10603 ( .A1(n8242), .A2(n8241), .ZN(n8373) );
  NAND2_X1 U10604 ( .A1(n8243), .A2(n8373), .ZN(n13400) );
  OR2_X1 U10605 ( .A1(n8257), .A2(n13400), .ZN(n8244) );
  NAND4_X1 U10606 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(n13241) );
  INV_X1 U10607 ( .A(n13241), .ZN(n8368) );
  NAND2_X1 U10608 ( .A1(n13409), .A2(n8368), .ZN(n8248) );
  NAND2_X1 U10609 ( .A1(n8357), .A2(n8248), .ZN(n12297) );
  INV_X1 U10610 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14363) );
  INV_X1 U10611 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12372) );
  MUX2_X1 U10612 ( .A(n14363), .B(n12372), .S(n6536), .Z(n11126) );
  XNOR2_X1 U10613 ( .A(n11126), .B(SI_29_), .ZN(n11124) );
  NAND2_X1 U10614 ( .A1(n12371), .A2(n12230), .ZN(n8254) );
  OR2_X1 U10615 ( .A1(n7832), .A2(n12372), .ZN(n8253) );
  NAND2_X1 U10616 ( .A1(n8255), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10617 ( .A1(n12218), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8260) );
  INV_X1 U10618 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15268) );
  OR2_X1 U10619 ( .A1(n8256), .A2(n15268), .ZN(n8259) );
  OR2_X1 U10620 ( .A1(n8257), .A2(n8373), .ZN(n8258) );
  NAND4_X1 U10621 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8258), .ZN(n13240) );
  XNOR2_X1 U10622 ( .A(n13616), .B(n13240), .ZN(n12299) );
  XNOR2_X1 U10623 ( .A(n8262), .B(n12299), .ZN(n13619) );
  NAND2_X1 U10624 ( .A1(n8263), .A2(n8264), .ZN(n8302) );
  NAND2_X1 U10625 ( .A1(n8269), .A2(n8265), .ZN(n8271) );
  NAND2_X1 U10626 ( .A1(n8271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8266) );
  MUX2_X1 U10627 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8266), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8268) );
  NAND2_X1 U10628 ( .A1(n8268), .A2(n8267), .ZN(n11061) );
  NOR2_X1 U10629 ( .A1(n8269), .A2(n7486), .ZN(n8270) );
  MUX2_X1 U10630 ( .A(n7486), .B(n8270), .S(P2_IR_REG_24__SCAN_IN), .Z(n8273)
         );
  INV_X1 U10631 ( .A(n8271), .ZN(n8272) );
  XNOR2_X1 U10632 ( .A(P2_B_REG_SCAN_IN), .B(n10954), .ZN(n8274) );
  NAND2_X1 U10633 ( .A1(n11061), .A2(n8274), .ZN(n8277) );
  NAND2_X1 U10634 ( .A1(n8267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8275) );
  INV_X1 U10635 ( .A(n13767), .ZN(n8276) );
  INV_X1 U10636 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14914) );
  NAND2_X1 U10637 ( .A1(n14908), .A2(n14914), .ZN(n8279) );
  NAND2_X1 U10638 ( .A1(n11061), .A2(n13767), .ZN(n8278) );
  NAND2_X1 U10639 ( .A1(n8279), .A2(n8278), .ZN(n14915) );
  NAND2_X1 U10640 ( .A1(n8280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8282) );
  XNOR2_X1 U10641 ( .A(n8282), .B(n8281), .ZN(n10685) );
  AND2_X1 U10642 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9329), .ZN(n8283) );
  INV_X1 U10643 ( .A(n14916), .ZN(n14913) );
  NOR2_X1 U10644 ( .A1(n14915), .A2(n14913), .ZN(n8294) );
  NOR4_X1 U10645 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8287) );
  NOR4_X1 U10646 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8286) );
  NOR4_X1 U10647 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8285) );
  NOR4_X1 U10648 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8284) );
  NAND4_X1 U10649 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n8293)
         );
  NOR2_X1 U10650 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .ZN(
        n8291) );
  NOR4_X1 U10651 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8290) );
  NOR4_X1 U10652 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8289) );
  NOR4_X1 U10653 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8288) );
  NAND4_X1 U10654 ( .A1(n8291), .A2(n8290), .A3(n8289), .A4(n8288), .ZN(n8292)
         );
  OAI21_X1 U10655 ( .B1(n8293), .B2(n8292), .A(n14908), .ZN(n9460) );
  NAND2_X1 U10656 ( .A1(n8294), .A2(n9460), .ZN(n9322) );
  INV_X1 U10657 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U10658 ( .A1(n14908), .A2(n14911), .ZN(n8296) );
  NAND2_X1 U10659 ( .A1(n10954), .A2(n13767), .ZN(n8295) );
  INV_X1 U10660 ( .A(n8263), .ZN(n8299) );
  NAND2_X1 U10661 ( .A1(n9718), .A2(n12044), .ZN(n12304) );
  NAND2_X1 U10662 ( .A1(n8299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10663 ( .A1(n8302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10664 ( .A1(n12304), .A2(n9324), .ZN(n9461) );
  NAND2_X1 U10665 ( .A1(n14912), .A2(n9461), .ZN(n8305) );
  OR2_X1 U10666 ( .A1(n9322), .A2(n8305), .ZN(n8308) );
  NAND2_X1 U10667 ( .A1(n12302), .A2(n9323), .ZN(n9459) );
  INV_X1 U10668 ( .A(n9459), .ZN(n8307) );
  INV_X1 U10669 ( .A(n12302), .ZN(n9536) );
  NOR2_X1 U10670 ( .A1(n9536), .A2(n9915), .ZN(n9537) );
  INV_X1 U10671 ( .A(n9537), .ZN(n8310) );
  NAND2_X1 U10672 ( .A1(n10068), .A2(n8310), .ZN(n14888) );
  OR2_X1 U10673 ( .A1(n12042), .A2(n12041), .ZN(n9533) );
  NAND2_X1 U10674 ( .A1(n12263), .A2(n9453), .ZN(n9452) );
  NAND2_X1 U10675 ( .A1(n9452), .A2(n8311), .ZN(n10163) );
  NAND2_X1 U10676 ( .A1(n10163), .A2(n12265), .ZN(n10162) );
  NAND2_X1 U10677 ( .A1(n10162), .A2(n8313), .ZN(n14890) );
  INV_X1 U10678 ( .A(n14886), .ZN(n14891) );
  NAND2_X1 U10679 ( .A1(n14889), .A2(n8314), .ZN(n10176) );
  INV_X1 U10680 ( .A(n12266), .ZN(n10175) );
  OR2_X1 U10681 ( .A1(n13265), .A2(n10182), .ZN(n8315) );
  INV_X1 U10682 ( .A(n13184), .ZN(n14947) );
  NAND2_X1 U10683 ( .A1(n14947), .A2(n13264), .ZN(n8316) );
  INV_X1 U10684 ( .A(n13264), .ZN(n8317) );
  NAND2_X1 U10685 ( .A1(n8317), .A2(n13184), .ZN(n8318) );
  NAND2_X1 U10686 ( .A1(n10071), .A2(n12269), .ZN(n8320) );
  INV_X1 U10687 ( .A(n13263), .ZN(n12086) );
  NAND2_X1 U10688 ( .A1(n12084), .A2(n12086), .ZN(n8319) );
  INV_X1 U10689 ( .A(n13262), .ZN(n9863) );
  AND2_X1 U10690 ( .A1(n12091), .A2(n9863), .ZN(n8321) );
  NOR2_X1 U10691 ( .A1(n14952), .A2(n12099), .ZN(n8322) );
  NAND2_X1 U10692 ( .A1(n14952), .A2(n12099), .ZN(n8323) );
  INV_X1 U10693 ( .A(n13260), .ZN(n8324) );
  NAND2_X1 U10694 ( .A1(n10677), .A2(n12278), .ZN(n10676) );
  INV_X1 U10695 ( .A(n13259), .ZN(n12111) );
  OR2_X1 U10696 ( .A1(n13601), .A2(n12111), .ZN(n8325) );
  XNOR2_X1 U10697 ( .A(n12115), .B(n13258), .ZN(n12279) );
  INV_X1 U10698 ( .A(n12279), .ZN(n10772) );
  INV_X1 U10699 ( .A(n13258), .ZN(n10389) );
  AND2_X1 U10700 ( .A1(n12115), .A2(n10389), .ZN(n10819) );
  NOR2_X1 U10701 ( .A1(n12277), .A2(n10819), .ZN(n8326) );
  XNOR2_X1 U10702 ( .A(n14819), .B(n13256), .ZN(n12281) );
  NAND2_X1 U10703 ( .A1(n8327), .A2(n12281), .ZN(n10807) );
  OR2_X1 U10704 ( .A1(n14819), .A2(n10567), .ZN(n8328) );
  NAND2_X1 U10705 ( .A1(n10807), .A2(n8328), .ZN(n10884) );
  INV_X1 U10706 ( .A(n13255), .ZN(n8330) );
  NAND2_X1 U10707 ( .A1(n12139), .A2(n8330), .ZN(n8329) );
  NAND2_X1 U10708 ( .A1(n10884), .A2(n8329), .ZN(n8332) );
  OR2_X1 U10709 ( .A1(n12139), .A2(n8330), .ZN(n8331) );
  NAND2_X1 U10710 ( .A1(n8332), .A2(n8331), .ZN(n10992) );
  INV_X1 U10711 ( .A(n13254), .ZN(n11111) );
  NOR2_X1 U10712 ( .A1(n13696), .A2(n11111), .ZN(n8333) );
  NAND2_X1 U10713 ( .A1(n13696), .A2(n11111), .ZN(n8334) );
  NAND2_X1 U10714 ( .A1(n8335), .A2(n8334), .ZN(n11098) );
  INV_X1 U10715 ( .A(n13252), .ZN(n8338) );
  NAND2_X1 U10716 ( .A1(n13739), .A2(n8338), .ZN(n8337) );
  OR2_X1 U10717 ( .A1(n13739), .A2(n8338), .ZN(n8339) );
  INV_X1 U10718 ( .A(n13251), .ZN(n13140) );
  NOR2_X1 U10719 ( .A1(n13735), .A2(n13140), .ZN(n8340) );
  NAND2_X1 U10720 ( .A1(n13735), .A2(n13140), .ZN(n8341) );
  XNOR2_X1 U10721 ( .A(n13672), .B(n13250), .ZN(n13536) );
  INV_X1 U10722 ( .A(n13250), .ZN(n8343) );
  OR2_X1 U10723 ( .A1(n13672), .A2(n8343), .ZN(n8344) );
  XNOR2_X1 U10724 ( .A(n13529), .B(n8345), .ZN(n13525) );
  NAND2_X1 U10725 ( .A1(n13529), .A2(n8345), .ZN(n8346) );
  INV_X1 U10726 ( .A(n13248), .ZN(n8347) );
  INV_X1 U10727 ( .A(n13494), .ZN(n8348) );
  NAND2_X1 U10728 ( .A1(n13490), .A2(n8348), .ZN(n8350) );
  OR2_X1 U10729 ( .A1(n13653), .A2(n13214), .ZN(n8349) );
  NOR2_X1 U10730 ( .A1(n13648), .A2(n13192), .ZN(n8351) );
  NAND2_X1 U10731 ( .A1(n13648), .A2(n13192), .ZN(n8352) );
  INV_X1 U10732 ( .A(n13245), .ZN(n13167) );
  NAND2_X1 U10733 ( .A1(n13643), .A2(n13167), .ZN(n8353) );
  NAND2_X1 U10734 ( .A1(n8354), .A2(n8353), .ZN(n13444) );
  AND2_X1 U10735 ( .A1(n13638), .A2(n13194), .ZN(n8355) );
  NAND2_X1 U10736 ( .A1(n13402), .A2(n8357), .ZN(n8358) );
  INV_X1 U10737 ( .A(n9718), .ZN(n12262) );
  NAND2_X1 U10738 ( .A1(n12262), .A2(n12301), .ZN(n12038) );
  NAND2_X1 U10739 ( .A1(n6527), .A2(n12305), .ZN(n8359) );
  INV_X1 U10740 ( .A(n8360), .ZN(n14845) );
  NAND2_X1 U10741 ( .A1(n14845), .A2(n9324), .ZN(n13191) );
  INV_X1 U10742 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10743 ( .A1(n12218), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10744 ( .A1(n8361), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8362) );
  OAI211_X1 U10745 ( .C1(n6525), .C2(n8364), .A(n8363), .B(n8362), .ZN(n13239)
         );
  INV_X1 U10746 ( .A(n13239), .ZN(n8367) );
  NAND2_X1 U10747 ( .A1(n8360), .A2(n9324), .ZN(n13193) );
  INV_X1 U10748 ( .A(P2_B_REG_SCAN_IN), .ZN(n8365) );
  NOR2_X1 U10749 ( .A1(n13761), .A2(n8365), .ZN(n8366) );
  OR2_X1 U10750 ( .A1(n13193), .A2(n8366), .ZN(n13388) );
  OAI22_X1 U10751 ( .A1(n8368), .A2(n13191), .B1(n8367), .B2(n13388), .ZN(
        n8369) );
  INV_X1 U10752 ( .A(n13638), .ZN(n13453) );
  NAND2_X1 U10753 ( .A1(n9451), .A2(n12041), .ZN(n10168) );
  INV_X1 U10754 ( .A(n14952), .ZN(n10412) );
  AND2_X2 U10755 ( .A1(n10409), .A2(n10412), .ZN(n10469) );
  INV_X1 U10756 ( .A(n12103), .ZN(n10517) );
  NAND2_X1 U10757 ( .A1(n10469), .A2(n10517), .ZN(n10674) );
  OR2_X2 U10758 ( .A1(n10674), .A2(n13601), .ZN(n10775) );
  OR2_X2 U10759 ( .A1(n10775), .A2(n12115), .ZN(n10815) );
  INV_X1 U10760 ( .A(n13743), .ZN(n11123) );
  NAND2_X1 U10761 ( .A1(n13453), .A2(n13472), .ZN(n13447) );
  AOI21_X1 U10762 ( .B1(n13616), .B2(n13408), .A(n14896), .ZN(n8370) );
  AND2_X1 U10763 ( .A1(n13395), .A2(n8370), .ZN(n13615) );
  INV_X1 U10764 ( .A(n9323), .ZN(n9532) );
  NOR2_X1 U10765 ( .A1(n9532), .A2(n9718), .ZN(n14900) );
  NAND2_X1 U10766 ( .A1(n13616), .A2(n13600), .ZN(n8372) );
  NAND2_X1 U10767 ( .A1(n13561), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8371) );
  OAI211_X1 U10768 ( .C1(n13595), .C2(n8373), .A(n8372), .B(n8371), .ZN(n8374)
         );
  INV_X1 U10769 ( .A(n9329), .ZN(n8376) );
  NAND2_X2 U10770 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8897), .ZN(n13268) );
  NOR2_X1 U10771 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8380) );
  NAND2_X1 U10772 ( .A1(n8387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8386) );
  INV_X1 U10773 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8385) );
  XNOR2_X1 U10774 ( .A(n8386), .B(n8385), .ZN(n8804) );
  INV_X1 U10775 ( .A(n8571), .ZN(n8575) );
  INV_X1 U10776 ( .A(n8390), .ZN(n9624) );
  NOR2_X1 U10777 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8394) );
  NOR2_X1 U10778 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n8393) );
  NAND4_X1 U10779 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n8607)
         );
  OR2_X2 U10780 ( .A1(n9624), .A2(n8607), .ZN(n8397) );
  INV_X1 U10781 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10782 ( .A1(n8397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8399) );
  INV_X1 U10783 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8398) );
  XNOR2_X1 U10784 ( .A(n8399), .B(n8398), .ZN(n11063) );
  NAND4_X1 U10785 ( .A1(n8402), .A2(n8401), .A3(n8516), .A4(n8544), .ZN(n8406)
         );
  NAND4_X1 U10786 ( .A1(n8583), .A2(n8537), .A3(n8404), .A4(n8403), .ZN(n8405)
         );
  NAND2_X1 U10787 ( .A1(n8710), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10788 ( .A1(n6589), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U10789 ( .A1(n8421), .A2(n8417), .ZN(n8423) );
  NAND2_X1 U10790 ( .A1(n8423), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U10791 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8418), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8419) );
  NAND2_X1 U10792 ( .A1(n10800), .A2(n8420), .ZN(n9199) );
  INV_X1 U10793 ( .A(n8421), .ZN(n9058) );
  NAND2_X1 U10794 ( .A1(n9058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8422) );
  MUX2_X1 U10795 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8422), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8424) );
  NAND2_X1 U10796 ( .A1(n8424), .A2(n8423), .ZN(n9198) );
  OR2_X2 U10797 ( .A1(n9199), .A2(n11729), .ZN(n12686) );
  NAND2_X1 U10798 ( .A1(n6536), .A2(P1_U3086), .ZN(n14372) );
  AND2_X1 U10799 ( .A1(n9161), .A2(P1_U3086), .ZN(n11731) );
  INV_X2 U10800 ( .A(n11731), .ZN(n14370) );
  INV_X1 U10801 ( .A(n14372), .ZN(n11732) );
  INV_X1 U10802 ( .A(n11732), .ZN(n11751) );
  NAND2_X1 U10803 ( .A1(n8425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8426) );
  MUX2_X1 U10804 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8426), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8427) );
  NAND2_X1 U10805 ( .A1(n8427), .A2(n6916), .ZN(n8679) );
  OAI222_X1 U10806 ( .A1(n11751), .A2(n8448), .B1(n14370), .B2(n9018), .C1(
        P1_U3086), .C2(n8679), .ZN(P1_U3353) );
  NAND2_X1 U10807 ( .A1(n6916), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8428) );
  MUX2_X1 U10808 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8428), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8430) );
  OR2_X1 U10809 ( .A1(n6916), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8432) );
  AND2_X1 U10810 ( .A1(n8430), .A2(n8432), .ZN(n13988) );
  INV_X1 U10811 ( .A(n13988), .ZN(n13982) );
  OAI222_X1 U10812 ( .A1(n11751), .A2(n8452), .B1(n14370), .B2(n9348), .C1(
        P1_U3086), .C2(n13982), .ZN(P1_U3352) );
  NAND2_X1 U10813 ( .A1(n9161), .A2(P2_U3088), .ZN(n13764) );
  NAND2_X1 U10814 ( .A1(n6535), .A2(P2_U3088), .ZN(n13766) );
  INV_X1 U10815 ( .A(n9512), .ZN(n8552) );
  NAND2_X1 U10816 ( .A1(n8432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8431) );
  MUX2_X1 U10817 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8431), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8435) );
  INV_X1 U10818 ( .A(n8432), .ZN(n8434) );
  NAND2_X1 U10819 ( .A1(n8434), .A2(n8433), .ZN(n8548) );
  NAND2_X1 U10820 ( .A1(n8435), .A2(n8548), .ZN(n8936) );
  OAI222_X1 U10821 ( .A1(n11751), .A2(n8456), .B1(n14370), .B2(n8552), .C1(
        P1_U3086), .C2(n8936), .ZN(P1_U3351) );
  INV_X1 U10822 ( .A(n9741), .ZN(n8554) );
  NAND2_X1 U10823 ( .A1(n8548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8436) );
  XNOR2_X1 U10824 ( .A(n8436), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9742) );
  INV_X1 U10825 ( .A(n9742), .ZN(n8734) );
  OAI222_X1 U10826 ( .A1(n11751), .A2(n8459), .B1(n14370), .B2(n8554), .C1(
        P1_U3086), .C2(n8734), .ZN(P1_U3350) );
  NOR2_X1 U10827 ( .A1(n6535), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13109) );
  INV_X2 U10828 ( .A(n13109), .ZN(n13120) );
  XNOR2_X1 U10829 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8444) );
  NAND2_X1 U10830 ( .A1(n8437), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8535) );
  XNOR2_X1 U10831 ( .A(n8444), .B(n8535), .ZN(n9248) );
  NAND2_X1 U10832 ( .A1(n6536), .A2(P3_U3151), .ZN(n13122) );
  CLKBUF_X1 U10833 ( .A(n13122), .Z(n13115) );
  INV_X1 U10834 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8438) );
  INV_X1 U10835 ( .A(n9065), .ZN(n8441) );
  OAI222_X1 U10836 ( .A1(n13120), .A2(n9248), .B1(n13115), .B2(n9247), .C1(
        P3_U3151), .C2(n9251), .ZN(P3_U3294) );
  NAND2_X1 U10837 ( .A1(n8543), .A2(n8544), .ZN(n8500) );
  OR2_X1 U10838 ( .A1(n8529), .A2(n8713), .ZN(n8442) );
  INV_X1 U10839 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8528) );
  XNOR2_X1 U10840 ( .A(n8442), .B(n8528), .ZN(n10662) );
  INV_X1 U10841 ( .A(n8535), .ZN(n8443) );
  NAND2_X1 U10842 ( .A1(n8444), .A2(n8443), .ZN(n8447) );
  NAND2_X1 U10843 ( .A1(n8445), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10844 ( .A1(n8447), .A2(n8446), .ZN(n8525) );
  NAND2_X1 U10845 ( .A1(n8556), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10846 ( .A1(n8448), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10847 ( .A1(n8525), .A2(n8524), .ZN(n8451) );
  NAND2_X1 U10848 ( .A1(n8451), .A2(n8450), .ZN(n8497) );
  NAND2_X1 U10849 ( .A1(n8559), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10850 ( .A1(n8452), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10851 ( .A1(n8497), .A2(n8496), .ZN(n8455) );
  NAND2_X1 U10852 ( .A1(n8455), .A2(n8454), .ZN(n8483) );
  NAND2_X1 U10853 ( .A1(n8456), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10854 ( .A1(n8459), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10855 ( .A1(n8551), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10856 ( .A1(n8547), .A2(n8462), .ZN(n8464) );
  NAND2_X1 U10857 ( .A1(n8558), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10858 ( .A1(n8560), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10859 ( .A1(n8466), .A2(n8465), .ZN(n8503) );
  NAND2_X1 U10860 ( .A1(n8582), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10861 ( .A1(n8467), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10862 ( .A1(n8592), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10863 ( .A1(n8628), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10864 ( .A1(n8474), .A2(n8472), .ZN(n8539) );
  INV_X1 U10865 ( .A(n8539), .ZN(n8473) );
  XNOR2_X1 U10866 ( .A(n8629), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8476) );
  XNOR2_X1 U10867 ( .A(n8532), .B(n8476), .ZN(n10691) );
  INV_X1 U10868 ( .A(n10691), .ZN(n8477) );
  OAI222_X1 U10869 ( .A1(P3_U3151), .A2(n10662), .B1(n13115), .B2(n8478), .C1(
        n13120), .C2(n8477), .ZN(P3_U3284) );
  NAND2_X1 U10870 ( .A1(n8479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8480) );
  MUX2_X1 U10871 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8480), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8481) );
  AND2_X1 U10872 ( .A1(n8486), .A2(n8481), .ZN(n9668) );
  INV_X1 U10873 ( .A(SI_4_), .ZN(n8485) );
  XNOR2_X1 U10874 ( .A(n8483), .B(n8482), .ZN(n9667) );
  INV_X1 U10875 ( .A(n9667), .ZN(n8484) );
  OAI222_X1 U10876 ( .A1(P3_U3151), .A2(n9094), .B1(n13115), .B2(n8485), .C1(
        n13120), .C2(n8484), .ZN(P3_U3291) );
  INV_X1 U10877 ( .A(n8543), .ZN(n8489) );
  NAND2_X1 U10878 ( .A1(n8486), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8487) );
  MUX2_X1 U10879 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8487), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8488) );
  NAND2_X1 U10880 ( .A1(n8489), .A2(n8488), .ZN(n9296) );
  INV_X1 U10881 ( .A(SI_5_), .ZN(n8493) );
  XNOR2_X1 U10882 ( .A(n8491), .B(n8490), .ZN(n9986) );
  INV_X1 U10883 ( .A(n9986), .ZN(n8492) );
  OAI222_X1 U10884 ( .A1(P3_U3151), .A2(n9296), .B1(n13115), .B2(n8493), .C1(
        n13120), .C2(n8492), .ZN(P3_U3290) );
  INV_X1 U10885 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10886 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6609), .ZN(n8494) );
  XNOR2_X1 U10887 ( .A(n8495), .B(n8494), .ZN(n9097) );
  XNOR2_X1 U10888 ( .A(n8497), .B(n8496), .ZN(n9485) );
  INV_X1 U10889 ( .A(n9485), .ZN(n8498) );
  OAI222_X1 U10890 ( .A1(P3_U3151), .A2(n9097), .B1(n13115), .B2(n8499), .C1(
        n13120), .C2(n8498), .ZN(P3_U3292) );
  NAND2_X1 U10891 ( .A1(n8500), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8502) );
  INV_X1 U10892 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8501) );
  XNOR2_X1 U10893 ( .A(n8502), .B(n8501), .ZN(n9612) );
  INV_X1 U10894 ( .A(SI_7_), .ZN(n8508) );
  NAND2_X1 U10895 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  AND2_X1 U10896 ( .A1(n8506), .A2(n8505), .ZN(n10262) );
  INV_X1 U10897 ( .A(n10262), .ZN(n8507) );
  OAI222_X1 U10898 ( .A1(P3_U3151), .A2(n9612), .B1(n13115), .B2(n8508), .C1(
        n13120), .C2(n8507), .ZN(P3_U3288) );
  OR2_X1 U10899 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10900 ( .A1(n8512), .A2(n8511), .ZN(n10268) );
  INV_X1 U10901 ( .A(SI_8_), .ZN(n10267) );
  NAND2_X1 U10902 ( .A1(n6562), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8513) );
  MUX2_X1 U10903 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8513), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8514) );
  AND2_X1 U10904 ( .A1(n8514), .A2(n8515), .ZN(n9610) );
  OAI222_X1 U10905 ( .A1(n13120), .A2(n10268), .B1(n13115), .B2(n10267), .C1(
        P3_U3151), .C2(n10271), .ZN(P3_U3287) );
  NAND2_X1 U10906 ( .A1(n8515), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U10907 ( .A(n8517), .B(n8516), .ZN(n14982) );
  INV_X1 U10908 ( .A(SI_9_), .ZN(n15215) );
  OR2_X1 U10909 ( .A1(n8519), .A2(n8518), .ZN(n8520) );
  AND2_X1 U10910 ( .A1(n8521), .A2(n8520), .ZN(n10251) );
  INV_X1 U10911 ( .A(n10251), .ZN(n8522) );
  OAI222_X1 U10912 ( .A1(P3_U3151), .A2(n14982), .B1(n13115), .B2(n15215), 
        .C1(n13120), .C2(n8522), .ZN(P3_U3286) );
  INV_X1 U10913 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8523) );
  INV_X1 U10914 ( .A(SI_2_), .ZN(n8527) );
  XNOR2_X1 U10915 ( .A(n8525), .B(n8524), .ZN(n9480) );
  INV_X1 U10916 ( .A(n9480), .ZN(n8526) );
  OAI222_X1 U10917 ( .A1(P3_U3151), .A2(n9069), .B1(n13115), .B2(n8527), .C1(
        n13120), .C2(n8526), .ZN(P3_U3293) );
  XNOR2_X1 U10918 ( .A(n8530), .B(P3_IR_REG_12__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U10919 ( .A1(n8629), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10920 ( .A1(n8633), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8533) );
  XNOR2_X1 U10921 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8586) );
  XNOR2_X1 U10922 ( .A(n8587), .B(n8586), .ZN(n10711) );
  OAI222_X1 U10923 ( .A1(P3_U3151), .A2(n10962), .B1(n13115), .B2(n10712), 
        .C1(n13120), .C2(n10711), .ZN(P3_U3283) );
  INV_X1 U10924 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10925 ( .A1(n8820), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8534) );
  AND2_X1 U10926 ( .A1(n8535), .A2(n8534), .ZN(n9162) );
  INV_X1 U10927 ( .A(SI_0_), .ZN(n9160) );
  OAI222_X1 U10928 ( .A1(P3_U3151), .A2(n15181), .B1(n13120), .B2(n9162), .C1(
        n9160), .C2(n13115), .ZN(P3_U3295) );
  XNOR2_X1 U10929 ( .A(n8538), .B(n8537), .ZN(n10522) );
  XNOR2_X1 U10930 ( .A(n8540), .B(n8539), .ZN(n10539) );
  INV_X1 U10931 ( .A(n10539), .ZN(n8542) );
  INV_X1 U10932 ( .A(SI_10_), .ZN(n8541) );
  OAI222_X1 U10933 ( .A1(n10522), .A2(P3_U3151), .B1(n13120), .B2(n8542), .C1(
        n8541), .C2(n13115), .ZN(P3_U3285) );
  OR2_X1 U10934 ( .A1(n8543), .A2(n8713), .ZN(n8545) );
  XNOR2_X1 U10935 ( .A(n8545), .B(n8544), .ZN(n10115) );
  XNOR2_X1 U10936 ( .A(n8558), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8546) );
  XNOR2_X1 U10937 ( .A(n8547), .B(n8546), .ZN(n10112) );
  INV_X1 U10938 ( .A(SI_6_), .ZN(n10111) );
  OAI222_X1 U10939 ( .A1(P3_U3151), .A2(n10115), .B1(n13120), .B2(n10112), 
        .C1(n10111), .C2(n13115), .ZN(P3_U3289) );
  INV_X1 U10940 ( .A(n9767), .ZN(n8557) );
  OAI21_X1 U10941 ( .B1(n8548), .B2(P1_IR_REG_5__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8549) );
  MUX2_X1 U10942 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8549), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8550) );
  AND2_X1 U10943 ( .A1(n8550), .A2(n8606), .ZN(n9768) );
  INV_X1 U10944 ( .A(n9768), .ZN(n8683) );
  OAI222_X1 U10945 ( .A1(n11751), .A2(n8551), .B1(n14370), .B2(n8557), .C1(
        P1_U3086), .C2(n8683), .ZN(P1_U3349) );
  INV_X1 U10946 ( .A(n13764), .ZN(n8577) );
  INV_X1 U10947 ( .A(n8577), .ZN(n13749) );
  INV_X1 U10948 ( .A(n13766), .ZN(n13755) );
  INV_X1 U10949 ( .A(n13755), .ZN(n10417) );
  OAI222_X1 U10950 ( .A1(n13749), .A2(n8553), .B1(n10417), .B2(n8552), .C1(
        P2_U3088), .C2(n8909), .ZN(P2_U3323) );
  INV_X1 U10951 ( .A(n9007), .ZN(n8911) );
  OAI222_X1 U10952 ( .A1(n13749), .A2(n8555), .B1(n10417), .B2(n8554), .C1(
        P2_U3088), .C2(n8911), .ZN(P2_U3322) );
  OAI222_X1 U10953 ( .A1(n13749), .A2(n8556), .B1(n10417), .B2(n9018), .C1(
        P2_U3088), .C2(n8906), .ZN(P2_U3325) );
  INV_X1 U10954 ( .A(n8973), .ZN(n8920) );
  OAI222_X1 U10955 ( .A1(n13749), .A2(n8558), .B1(n10417), .B2(n8557), .C1(
        P2_U3088), .C2(n8920), .ZN(P2_U3321) );
  OAI222_X1 U10956 ( .A1(n13749), .A2(n8559), .B1(n10417), .B2(n9348), .C1(
        P2_U3088), .C2(n8908), .ZN(P2_U3324) );
  INV_X1 U10957 ( .A(n9928), .ZN(n8562) );
  INV_X1 U10958 ( .A(n9634), .ZN(n8977) );
  OAI222_X1 U10959 ( .A1(n13749), .A2(n8560), .B1(n10417), .B2(n8562), .C1(
        P2_U3088), .C2(n8977), .ZN(P2_U3320) );
  NAND2_X1 U10960 ( .A1(n8606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U10961 ( .A(n8561), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9929) );
  INV_X1 U10962 ( .A(n9929), .ZN(n8707) );
  OAI222_X1 U10963 ( .A1(n11751), .A2(n15259), .B1(n14370), .B2(n8562), .C1(
        P1_U3086), .C2(n8707), .ZN(P1_U3348) );
  INV_X1 U10964 ( .A(P3_B_REG_SCAN_IN), .ZN(n8563) );
  XNOR2_X1 U10965 ( .A(n10581), .B(n8563), .ZN(n8564) );
  NAND2_X1 U10966 ( .A1(n8564), .A2(n10768), .ZN(n8565) );
  INV_X1 U10967 ( .A(n9176), .ZN(n8634) );
  INV_X1 U10968 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10969 ( .A1(n8634), .A2(n8566), .ZN(n8569) );
  OR2_X1 U10970 ( .A1(n10800), .A2(n8567), .ZN(n8568) );
  NAND2_X1 U10971 ( .A1(n8569), .A2(n8568), .ZN(n9556) );
  NAND2_X1 U10972 ( .A1(n11729), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8570) );
  OAI21_X1 U10973 ( .B1(n9556), .B2(n11729), .A(n8570), .ZN(P3_U3377) );
  INV_X1 U10974 ( .A(n8835), .ZN(n8831) );
  NAND3_X1 U10975 ( .A1(n11799), .A2(P1_B_REG_SCAN_IN), .A3(n11063), .ZN(n8572) );
  NAND3_X1 U10976 ( .A1(n8573), .A2(n8572), .A3(n8574), .ZN(n8797) );
  INV_X1 U10977 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8576) );
  NOR2_X1 U10978 ( .A1(n8575), .A2(n8574), .ZN(n11797) );
  AOI22_X1 U10979 ( .A1(n14749), .A2(n8576), .B1(n11797), .B2(n11063), .ZN(
        P1_U3446) );
  INV_X1 U10980 ( .A(n10018), .ZN(n8581) );
  NAND2_X1 U10981 ( .A1(n8577), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10982 ( .A1(n9635), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14844) );
  OAI211_X1 U10983 ( .C1(n8581), .C2(n10417), .A(n8578), .B(n14844), .ZN(
        P2_U3319) );
  NOR2_X1 U10984 ( .A1(n8606), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8594) );
  INV_X1 U10985 ( .A(n8594), .ZN(n8579) );
  NAND2_X1 U10986 ( .A1(n8579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8580) );
  XNOR2_X1 U10987 ( .A(n8580), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10019) );
  INV_X1 U10988 ( .A(n10019), .ZN(n8750) );
  OAI222_X1 U10989 ( .A1(n11751), .A2(n8582), .B1(n14370), .B2(n8581), .C1(
        P1_U3086), .C2(n8750), .ZN(P1_U3347) );
  NAND2_X1 U10990 ( .A1(n8584), .A2(n8583), .ZN(n8616) );
  NAND2_X1 U10991 ( .A1(n8616), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U10992 ( .A(n8585), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12707) );
  INV_X1 U10993 ( .A(n12707), .ZN(n12693) );
  NAND2_X1 U10994 ( .A1(n8588), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10995 ( .A(n8618), .B(n8874), .ZN(n10867) );
  INV_X1 U10996 ( .A(n10867), .ZN(n8590) );
  OAI222_X1 U10997 ( .A1(P3_U3151), .A2(n12693), .B1(n13115), .B2(n8591), .C1(
        n13120), .C2(n8590), .ZN(P3_U3282) );
  INV_X1 U10998 ( .A(n10024), .ZN(n8597) );
  INV_X1 U10999 ( .A(n9636), .ZN(n13287) );
  OAI222_X1 U11000 ( .A1(n13749), .A2(n8592), .B1(n10417), .B2(n8597), .C1(
        P2_U3088), .C2(n13287), .ZN(P2_U3318) );
  INV_X1 U11001 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8593) );
  INV_X1 U11002 ( .A(n8624), .ZN(n8595) );
  NAND2_X1 U11003 ( .A1(n8595), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8596) );
  XNOR2_X1 U11004 ( .A(n8596), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10025) );
  INV_X1 U11005 ( .A(n10025), .ZN(n8773) );
  OAI222_X1 U11006 ( .A1(n11751), .A2(n8598), .B1(n14370), .B2(n8597), .C1(
        P1_U3086), .C2(n8773), .ZN(P1_U3346) );
  INV_X1 U11007 ( .A(n8804), .ZN(n8599) );
  NAND2_X1 U11008 ( .A1(n8599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11692) );
  NAND2_X1 U11009 ( .A1(n8835), .A2(n11692), .ZN(n8664) );
  NAND2_X1 U11010 ( .A1(n8602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8603) );
  MUX2_X1 U11011 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8603), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8605) );
  NAND2_X1 U11012 ( .A1(n8605), .A2(n8604), .ZN(n11308) );
  NAND2_X1 U11013 ( .A1(n14374), .A2(n11633), .ZN(n11332) );
  INV_X1 U11014 ( .A(n8607), .ZN(n8609) );
  NOR2_X1 U11015 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8608) );
  AND2_X2 U11016 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  INV_X1 U11017 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8612) );
  AOI21_X1 U11018 ( .B1(n8889), .B2(n8804), .A(n11455), .ZN(n8663) );
  INV_X1 U11019 ( .A(n8663), .ZN(n8615) );
  AND2_X1 U11020 ( .A1(n8664), .A2(n8615), .ZN(n14715) );
  CLKBUF_X2 U11021 ( .A(P1_U4016), .Z(n13956) );
  NOR2_X1 U11022 ( .A1(n14715), .A2(n13956), .ZN(P1_U3085) );
  NAND2_X1 U11023 ( .A1(n8687), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U11024 ( .A(n8617), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12699) );
  INV_X1 U11025 ( .A(n12699), .ZN(n12690) );
  NAND2_X1 U11026 ( .A1(n8619), .A2(n8872), .ZN(n8620) );
  XNOR2_X1 U11027 ( .A(n9315), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U11028 ( .A(n8690), .B(n8621), .ZN(n10912) );
  INV_X1 U11029 ( .A(n10912), .ZN(n8622) );
  OAI222_X1 U11030 ( .A1(P3_U3151), .A2(n12690), .B1(n13115), .B2(n6716), .C1(
        n13120), .C2(n8622), .ZN(P3_U3281) );
  INV_X1 U11031 ( .A(n10215), .ZN(n8627) );
  INV_X1 U11032 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11033 ( .A1(n8624), .A2(n8623), .ZN(n8630) );
  NAND2_X1 U11034 ( .A1(n8630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8625) );
  XNOR2_X1 U11035 ( .A(n8625), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10216) );
  INV_X1 U11036 ( .A(n10216), .ZN(n8781) );
  OAI222_X1 U11037 ( .A1(n11751), .A2(n8626), .B1(n14370), .B2(n8627), .C1(
        P1_U3086), .C2(n8781), .ZN(P1_U3345) );
  OAI222_X1 U11038 ( .A1(n13749), .A2(n8628), .B1(n10417), .B2(n8627), .C1(
        P2_U3088), .C2(n9637), .ZN(P2_U3317) );
  INV_X1 U11039 ( .A(n10345), .ZN(n8632) );
  OAI222_X1 U11040 ( .A1(n13749), .A2(n8629), .B1(n10417), .B2(n8632), .C1(
        P2_U3088), .C2(n11075), .ZN(P2_U3316) );
  NAND2_X1 U11041 ( .A1(n8661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8631) );
  XNOR2_X1 U11042 ( .A(n8631), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10346) );
  INV_X1 U11043 ( .A(n10346), .ZN(n8949) );
  OAI222_X1 U11044 ( .A1(n11751), .A2(n8633), .B1(n14370), .B2(n8632), .C1(
        P1_U3086), .C2(n8949), .ZN(P1_U3344) );
  NOR2_X1 U11045 ( .A1(n8634), .A2(n11729), .ZN(n8636) );
  CLKBUF_X1 U11046 ( .A(n8636), .Z(n8660) );
  INV_X1 U11047 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n15186) );
  NOR2_X1 U11048 ( .A1(n8660), .A2(n15186), .ZN(P3_U3256) );
  INV_X1 U11049 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n8635) );
  NOR2_X1 U11050 ( .A1(n8660), .A2(n8635), .ZN(P3_U3257) );
  INV_X1 U11051 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n8637) );
  NOR2_X1 U11052 ( .A1(n8660), .A2(n8637), .ZN(P3_U3258) );
  INV_X1 U11053 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n8638) );
  NOR2_X1 U11054 ( .A1(n8660), .A2(n8638), .ZN(P3_U3259) );
  INV_X1 U11055 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n15253) );
  NOR2_X1 U11056 ( .A1(n8660), .A2(n15253), .ZN(P3_U3263) );
  INV_X1 U11057 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n8639) );
  NOR2_X1 U11058 ( .A1(n8636), .A2(n8639), .ZN(P3_U3239) );
  INV_X1 U11059 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n8640) );
  NOR2_X1 U11060 ( .A1(n8636), .A2(n8640), .ZN(P3_U3238) );
  INV_X1 U11061 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n8641) );
  NOR2_X1 U11062 ( .A1(n8636), .A2(n8641), .ZN(P3_U3237) );
  INV_X1 U11063 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n8642) );
  NOR2_X1 U11064 ( .A1(n8636), .A2(n8642), .ZN(P3_U3236) );
  INV_X1 U11065 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n8643) );
  NOR2_X1 U11066 ( .A1(n8636), .A2(n8643), .ZN(P3_U3235) );
  INV_X1 U11067 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15290) );
  NOR2_X1 U11068 ( .A1(n8636), .A2(n15290), .ZN(P3_U3234) );
  INV_X1 U11069 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15159) );
  NOR2_X1 U11070 ( .A1(n8636), .A2(n15159), .ZN(P3_U3260) );
  INV_X1 U11071 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n8644) );
  NOR2_X1 U11072 ( .A1(n8660), .A2(n8644), .ZN(P3_U3261) );
  INV_X1 U11073 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n15361) );
  NOR2_X1 U11074 ( .A1(n8636), .A2(n15361), .ZN(P3_U3262) );
  INV_X1 U11075 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n8645) );
  NOR2_X1 U11076 ( .A1(n8636), .A2(n8645), .ZN(P3_U3242) );
  INV_X1 U11077 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n8646) );
  NOR2_X1 U11078 ( .A1(n8636), .A2(n8646), .ZN(P3_U3241) );
  INV_X1 U11079 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n8647) );
  NOR2_X1 U11080 ( .A1(n8636), .A2(n8647), .ZN(P3_U3240) );
  INV_X1 U11081 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n8648) );
  NOR2_X1 U11082 ( .A1(n8660), .A2(n8648), .ZN(P3_U3254) );
  INV_X1 U11083 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n8649) );
  NOR2_X1 U11084 ( .A1(n8660), .A2(n8649), .ZN(P3_U3253) );
  INV_X1 U11085 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n8650) );
  NOR2_X1 U11086 ( .A1(n8660), .A2(n8650), .ZN(P3_U3252) );
  INV_X1 U11087 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U11088 ( .A1(n8660), .A2(n15362), .ZN(P3_U3251) );
  INV_X1 U11089 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n8651) );
  NOR2_X1 U11090 ( .A1(n8660), .A2(n8651), .ZN(P3_U3250) );
  INV_X1 U11091 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n8652) );
  NOR2_X1 U11092 ( .A1(n8660), .A2(n8652), .ZN(P3_U3249) );
  INV_X1 U11093 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n8653) );
  NOR2_X1 U11094 ( .A1(n8660), .A2(n8653), .ZN(P3_U3248) );
  INV_X1 U11095 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n8654) );
  NOR2_X1 U11096 ( .A1(n8660), .A2(n8654), .ZN(P3_U3247) );
  INV_X1 U11097 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n8655) );
  NOR2_X1 U11098 ( .A1(n8660), .A2(n8655), .ZN(P3_U3246) );
  INV_X1 U11099 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n8656) );
  NOR2_X1 U11100 ( .A1(n8660), .A2(n8656), .ZN(P3_U3245) );
  INV_X1 U11101 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n8657) );
  NOR2_X1 U11102 ( .A1(n8660), .A2(n8657), .ZN(P3_U3244) );
  INV_X1 U11103 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n8658) );
  NOR2_X1 U11104 ( .A1(n8660), .A2(n8658), .ZN(P3_U3243) );
  INV_X1 U11105 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n8659) );
  NOR2_X1 U11106 ( .A1(n8660), .A2(n8659), .ZN(P3_U3255) );
  INV_X1 U11107 ( .A(n10594), .ZN(n8735) );
  OAI21_X1 U11108 ( .B1(n8661), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8870) );
  XNOR2_X1 U11109 ( .A(n8870), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U11110 ( .A1(n14006), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11732), .ZN(n8662) );
  OAI21_X1 U11111 ( .B1(n8735), .B2(n14370), .A(n8662), .ZN(P1_U3343) );
  NAND2_X1 U11112 ( .A1(n8664), .A2(n8663), .ZN(n14718) );
  OR3_X1 U11113 ( .A1(n14718), .A2(n6526), .A3(n11748), .ZN(n14021) );
  INV_X1 U11114 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8883) );
  MUX2_X1 U11115 ( .A(n8883), .B(P1_REG2_REG_2__SCAN_IN), .S(n8679), .Z(n13974) );
  INV_X1 U11116 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U11117 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9661), .S(n13960), .Z(
        n13966) );
  AND2_X1 U11118 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8665) );
  NAND2_X1 U11119 ( .A1(n13966), .A2(n8665), .ZN(n13965) );
  NAND2_X1 U11120 ( .A1(n13960), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11121 ( .A1(n13965), .A2(n8666), .ZN(n13973) );
  NAND2_X1 U11122 ( .A1(n13974), .A2(n13973), .ZN(n13990) );
  INV_X1 U11123 ( .A(n8679), .ZN(n13972) );
  NAND2_X1 U11124 ( .A1(n13972), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13989) );
  NAND2_X1 U11125 ( .A1(n13990), .A2(n13989), .ZN(n8668) );
  INV_X1 U11126 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9022) );
  MUX2_X1 U11127 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9022), .S(n13988), .Z(n8667) );
  NAND2_X1 U11128 ( .A1(n8668), .A2(n8667), .ZN(n13993) );
  NAND2_X1 U11129 ( .A1(n13988), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11130 ( .A1(n13993), .A2(n8932), .ZN(n8670) );
  INV_X1 U11131 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9360) );
  MUX2_X1 U11132 ( .A(n9360), .B(P1_REG2_REG_4__SCAN_IN), .S(n8936), .Z(n8669)
         );
  NAND2_X1 U11133 ( .A1(n8670), .A2(n8669), .ZN(n8934) );
  INV_X1 U11134 ( .A(n8936), .ZN(n9513) );
  NAND2_X1 U11135 ( .A1(n9513), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11136 ( .A1(n8934), .A2(n8726), .ZN(n8672) );
  INV_X1 U11137 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U11138 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9760), .S(n9742), .Z(n8671)
         );
  NAND2_X1 U11139 ( .A1(n8672), .A2(n8671), .ZN(n8728) );
  NAND2_X1 U11140 ( .A1(n9742), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11141 ( .A1(n8728), .A2(n8676), .ZN(n8674) );
  INV_X1 U11142 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9786) );
  MUX2_X1 U11143 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9786), .S(n9768), .Z(n8673)
         );
  NAND2_X1 U11144 ( .A1(n8674), .A2(n8673), .ZN(n8702) );
  MUX2_X1 U11145 ( .A(n9786), .B(P1_REG2_REG_6__SCAN_IN), .S(n9768), .Z(n8675)
         );
  NAND3_X1 U11146 ( .A1(n8728), .A2(n8676), .A3(n8675), .ZN(n8677) );
  AND3_X1 U11147 ( .A1(n14728), .A2(n8702), .A3(n8677), .ZN(n8686) );
  MUX2_X1 U11148 ( .A(n14800), .B(P1_REG1_REG_6__SCAN_IN), .S(n9768), .Z(n8681) );
  INV_X1 U11149 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9023) );
  INV_X1 U11150 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8884) );
  INV_X1 U11151 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8678) );
  XOR2_X1 U11152 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n13960), .Z(n13963) );
  NAND3_X1 U11153 ( .A1(n13963), .A2(P1_REG1_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n13961) );
  OAI21_X1 U11154 ( .B1(n6931), .B2(n8678), .A(n13961), .ZN(n13976) );
  MUX2_X1 U11155 ( .A(n8884), .B(P1_REG1_REG_2__SCAN_IN), .S(n8679), .Z(n13977) );
  NAND2_X1 U11156 ( .A1(n13976), .A2(n13977), .ZN(n13975) );
  OAI21_X1 U11157 ( .B1(n8679), .B2(n8884), .A(n13975), .ZN(n13986) );
  MUX2_X1 U11158 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9023), .S(n13988), .Z(
        n13987) );
  NAND2_X1 U11159 ( .A1(n13986), .A2(n13987), .ZN(n13985) );
  OAI21_X1 U11160 ( .B1(n9023), .B2(n13982), .A(n13985), .ZN(n8928) );
  INV_X1 U11161 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9529) );
  MUX2_X1 U11162 ( .A(n9529), .B(P1_REG1_REG_4__SCAN_IN), .S(n8936), .Z(n8929)
         );
  AOI22_X1 U11163 ( .A1(n8928), .A2(n8929), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n9513), .ZN(n8723) );
  INV_X1 U11164 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9518) );
  XNOR2_X1 U11165 ( .A(n9742), .B(n9518), .ZN(n8724) );
  INV_X1 U11166 ( .A(n6526), .ZN(n11688) );
  AOI211_X1 U11167 ( .C1(n8681), .C2(n8680), .A(n8695), .B(n10634), .ZN(n8685)
         );
  INV_X1 U11168 ( .A(n11748), .ZN(n8926) );
  NAND2_X1 U11169 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U11170 ( .A1(n14715), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8682) );
  OAI211_X1 U11171 ( .C1(n14020), .C2(n8683), .A(n10156), .B(n8682), .ZN(n8684) );
  OR3_X1 U11172 ( .A1(n8686), .A2(n8685), .A3(n8684), .ZN(P1_U3249) );
  OAI21_X1 U11173 ( .B1(n8687), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8688) );
  XNOR2_X1 U11174 ( .A(n8688), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12742) );
  INV_X1 U11175 ( .A(n12742), .ZN(n12755) );
  AND2_X1 U11176 ( .A1(n9313), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11177 ( .A1(n9315), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11178 ( .A1(n9417), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U11179 ( .A1(n9419), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U11180 ( .A(n8864), .B(n8862), .ZN(n11006) );
  INV_X1 U11181 ( .A(n11006), .ZN(n8693) );
  OAI222_X1 U11182 ( .A1(P3_U3151), .A2(n12755), .B1(n13122), .B2(n8694), .C1(
        n13120), .C2(n8693), .ZN(P3_U3280) );
  MUX2_X1 U11183 ( .A(n14802), .B(P1_REG1_REG_7__SCAN_IN), .S(n9929), .Z(n8696) );
  NOR2_X1 U11184 ( .A1(n8697), .A2(n8696), .ZN(n8738) );
  AOI211_X1 U11185 ( .C1(n8697), .C2(n8696), .A(n10634), .B(n8738), .ZN(n8709)
         );
  NAND2_X1 U11186 ( .A1(n9768), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11187 ( .A1(n8702), .A2(n8701), .ZN(n8699) );
  INV_X1 U11188 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9947) );
  MUX2_X1 U11189 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9947), .S(n9929), .Z(n8698)
         );
  NAND2_X1 U11190 ( .A1(n8699), .A2(n8698), .ZN(n8745) );
  MUX2_X1 U11191 ( .A(n9947), .B(P1_REG2_REG_7__SCAN_IN), .S(n9929), .Z(n8700)
         );
  NAND3_X1 U11192 ( .A1(n8702), .A2(n8701), .A3(n8700), .ZN(n8703) );
  NAND3_X1 U11193 ( .A1(n14728), .A2(n8745), .A3(n8703), .ZN(n8706) );
  NAND2_X1 U11194 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10329) );
  INV_X1 U11195 ( .A(n10329), .ZN(n8704) );
  AOI21_X1 U11196 ( .B1(n14715), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n8704), .ZN(
        n8705) );
  OAI211_X1 U11197 ( .C1(n14020), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8708)
         );
  OR2_X1 U11198 ( .A1(n8709), .A2(n8708), .ZN(P1_U3250) );
  INV_X1 U11199 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15316) );
  MUX2_X1 U11200 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8711), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8712) );
  INV_X1 U11201 ( .A(n8714), .ZN(n13111) );
  XNOR2_X2 U11202 ( .A(n7702), .B(n13112), .ZN(n12569) );
  AND2_X2 U11203 ( .A1(n8715), .A2(n12569), .ZN(n10084) );
  NAND2_X1 U11204 ( .A1(n6530), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8720) );
  AND2_X4 U11205 ( .A1(n8716), .A2(n8715), .ZN(n11154) );
  NAND2_X1 U11206 ( .A1(n11154), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11207 ( .A1(n6532), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11208 ( .A1(n9678), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11209 ( .A1(n15064), .A2(P3_U3897), .ZN(n8721) );
  OAI21_X1 U11210 ( .B1(P3_U3897), .B2(n15316), .A(n8721), .ZN(P3_U3493) );
  INV_X1 U11211 ( .A(n10634), .ZN(n14727) );
  OAI21_X1 U11212 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8730) );
  MUX2_X1 U11213 ( .A(n9760), .B(P1_REG2_REG_5__SCAN_IN), .S(n9742), .Z(n8725)
         );
  NAND3_X1 U11214 ( .A1(n8934), .A2(n8726), .A3(n8725), .ZN(n8727) );
  AND3_X1 U11215 ( .A1(n14728), .A2(n8728), .A3(n8727), .ZN(n8729) );
  AOI21_X1 U11216 ( .B1(n14727), .B2(n8730), .A(n8729), .ZN(n8733) );
  NAND2_X1 U11217 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9825) );
  INV_X1 U11218 ( .A(n9825), .ZN(n8731) );
  AOI21_X1 U11219 ( .B1(n14715), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n8731), .ZN(
        n8732) );
  OAI211_X1 U11220 ( .C1(n8734), .C2(n14020), .A(n8733), .B(n8732), .ZN(
        P1_U3248) );
  INV_X1 U11221 ( .A(n11076), .ZN(n13302) );
  OAI222_X1 U11222 ( .A1(n13749), .A2(n8736), .B1(n10417), .B2(n8735), .C1(
        P2_U3088), .C2(n13302), .ZN(P2_U3315) );
  NAND2_X1 U11223 ( .A1(n12042), .A2(P2_U3947), .ZN(n8737) );
  OAI21_X1 U11224 ( .B1(n8820), .B2(P2_U3947), .A(n8737), .ZN(P2_U3531) );
  AOI21_X1 U11225 ( .B1(n9929), .B2(P1_REG1_REG_7__SCAN_IN), .A(n8738), .ZN(
        n8740) );
  INV_X1 U11226 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9936) );
  MUX2_X1 U11227 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9936), .S(n10019), .Z(n8739) );
  OAI21_X1 U11228 ( .B1(n8740), .B2(n8739), .A(n8754), .ZN(n8752) );
  NAND2_X1 U11229 ( .A1(n9929), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11230 ( .A1(n8745), .A2(n8744), .ZN(n8742) );
  INV_X1 U11231 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10063) );
  MUX2_X1 U11232 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10063), .S(n10019), .Z(
        n8741) );
  NAND2_X1 U11233 ( .A1(n8742), .A2(n8741), .ZN(n8759) );
  MUX2_X1 U11234 ( .A(n10063), .B(P1_REG2_REG_8__SCAN_IN), .S(n10019), .Z(
        n8743) );
  NAND3_X1 U11235 ( .A1(n8745), .A2(n8744), .A3(n8743), .ZN(n8746) );
  NAND3_X1 U11236 ( .A1(n14728), .A2(n8759), .A3(n8746), .ZN(n8749) );
  NAND2_X1 U11237 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10504) );
  INV_X1 U11238 ( .A(n10504), .ZN(n8747) );
  AOI21_X1 U11239 ( .B1(n14715), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n8747), .ZN(
        n8748) );
  OAI211_X1 U11240 ( .C1(n14020), .C2(n8750), .A(n8749), .B(n8748), .ZN(n8751)
         );
  AOI21_X1 U11241 ( .B1(n8752), .B2(n14727), .A(n8751), .ZN(n8753) );
  INV_X1 U11242 ( .A(n8753), .ZN(P1_U3251) );
  INV_X1 U11243 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10028) );
  MUX2_X1 U11244 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10028), .S(n10025), .Z(
        n8756) );
  OAI21_X1 U11245 ( .B1(n8756), .B2(n8755), .A(n8769), .ZN(n8766) );
  NAND2_X1 U11246 ( .A1(n10019), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8758) );
  INV_X1 U11247 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8772) );
  MUX2_X1 U11248 ( .A(n8772), .B(P1_REG2_REG_9__SCAN_IN), .S(n10025), .Z(n8757) );
  AOI21_X1 U11249 ( .B1(n8759), .B2(n8758), .A(n8757), .ZN(n8776) );
  INV_X1 U11250 ( .A(n8776), .ZN(n8761) );
  NAND3_X1 U11251 ( .A1(n8759), .A2(n8758), .A3(n8757), .ZN(n8760) );
  NAND3_X1 U11252 ( .A1(n8761), .A2(n14728), .A3(n8760), .ZN(n8764) );
  NAND2_X1 U11253 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10791) );
  INV_X1 U11254 ( .A(n10791), .ZN(n8762) );
  AOI21_X1 U11255 ( .B1(n14715), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8762), .ZN(
        n8763) );
  OAI211_X1 U11256 ( .C1(n14020), .C2(n8773), .A(n8764), .B(n8763), .ZN(n8765)
         );
  AOI21_X1 U11257 ( .B1(n8766), .B2(n14727), .A(n8765), .ZN(n8767) );
  INV_X1 U11258 ( .A(n8767), .ZN(P1_U3252) );
  INV_X1 U11259 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8768) );
  MUX2_X1 U11260 ( .A(n8768), .B(P1_REG1_REG_10__SCAN_IN), .S(n10216), .Z(
        n8771) );
  NOR2_X1 U11261 ( .A1(n8770), .A2(n8771), .ZN(n8945) );
  AOI211_X1 U11262 ( .C1(n8771), .C2(n8770), .A(n10634), .B(n8945), .ZN(n8784)
         );
  NOR2_X1 U11263 ( .A1(n8773), .A2(n8772), .ZN(n8775) );
  INV_X1 U11264 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U11265 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10222), .S(n10216), .Z(
        n8774) );
  OAI21_X1 U11266 ( .B1(n8776), .B2(n8775), .A(n8774), .ZN(n8943) );
  INV_X1 U11267 ( .A(n8943), .ZN(n8778) );
  NOR3_X1 U11268 ( .A1(n8776), .A2(n8775), .A3(n8774), .ZN(n8777) );
  NOR3_X1 U11269 ( .A1(n8778), .A2(n8777), .A3(n14021), .ZN(n8783) );
  NAND2_X1 U11270 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10849)
         );
  INV_X1 U11271 ( .A(n10849), .ZN(n8779) );
  AOI21_X1 U11272 ( .B1(n14715), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8779), .ZN(
        n8780) );
  OAI21_X1 U11273 ( .B1(n14020), .B2(n8781), .A(n8780), .ZN(n8782) );
  OR3_X1 U11274 ( .A1(n8784), .A2(n8783), .A3(n8782), .ZN(P1_U3253) );
  OR2_X1 U11275 ( .A1(n8797), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11276 ( .A1(n14368), .A2(n11063), .ZN(n8785) );
  AND2_X1 U11277 ( .A1(n8786), .A2(n8785), .ZN(n9220) );
  NOR4_X1 U11278 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n8795) );
  NOR4_X1 U11279 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8794) );
  INV_X1 U11280 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15182) );
  INV_X1 U11281 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15199) );
  INV_X1 U11282 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15239) );
  INV_X1 U11283 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15360) );
  NAND4_X1 U11284 ( .A1(n15182), .A2(n15199), .A3(n15239), .A4(n15360), .ZN(
        n8792) );
  NOR4_X1 U11285 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n8790) );
  NOR4_X1 U11286 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8789) );
  NOR4_X1 U11287 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8788) );
  NOR4_X1 U11288 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8787) );
  NAND4_X1 U11289 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n8791)
         );
  NOR4_X1 U11290 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8792), .A4(n8791), .ZN(n8793) );
  AND3_X1 U11291 ( .A1(n8795), .A2(n8794), .A3(n8793), .ZN(n8796) );
  AND2_X1 U11292 ( .A1(n9220), .A2(n9218), .ZN(n9647) );
  NAND2_X1 U11293 ( .A1(n11799), .A2(n14368), .ZN(n8798) );
  NAND2_X1 U11294 ( .A1(n9647), .A2(n9243), .ZN(n8837) );
  NAND2_X1 U11295 ( .A1(n11305), .A2(n11635), .ZN(n11331) );
  NAND2_X1 U11296 ( .A1(n8808), .A2(n11352), .ZN(n9217) );
  NAND2_X1 U11297 ( .A1(n8837), .A2(n9217), .ZN(n8807) );
  NAND2_X1 U11298 ( .A1(n11635), .A2(n14635), .ZN(n8827) );
  INV_X1 U11299 ( .A(n8834), .ZN(n8805) );
  AND3_X1 U11300 ( .A1(n8805), .A2(n8825), .A3(n8804), .ZN(n8806) );
  NAND2_X1 U11301 ( .A1(n8807), .A2(n8806), .ZN(n9358) );
  NOR2_X1 U11302 ( .A1(n9358), .A2(P1_U3086), .ZN(n9031) );
  INV_X1 U11303 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U11304 ( .A1(n11564), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8818) );
  OR2_X1 U11305 ( .A1(n11608), .A2(n9917), .ZN(n8817) );
  INV_X1 U11306 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8813) );
  INV_X1 U11307 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14707) );
  OAI21_X1 U11308 ( .B1(n6535), .B2(n9160), .A(n8820), .ZN(n8821) );
  NAND2_X1 U11309 ( .A1(n8822), .A2(n8821), .ZN(n14375) );
  MUX2_X1 U11310 ( .A(n7491), .B(n14375), .S(n11516), .Z(n9919) );
  INV_X1 U11311 ( .A(n9919), .ZN(n9230) );
  INV_X1 U11312 ( .A(n8825), .ZN(n8823) );
  INV_X1 U11313 ( .A(n13957), .ZN(n9654) );
  OAI222_X1 U11314 ( .A1(n9919), .A2(n12543), .B1(n12545), .B2(n9654), .C1(
        n8825), .C2(n14707), .ZN(n8882) );
  OAI21_X1 U11315 ( .B1(n8826), .B2(n8882), .A(n8881), .ZN(n8924) );
  NAND2_X1 U11316 ( .A1(n11305), .A2(n11308), .ZN(n9227) );
  INV_X1 U11317 ( .A(n8827), .ZN(n8828) );
  NAND2_X1 U11318 ( .A1(n14793), .A2(n11332), .ZN(n8829) );
  OR2_X1 U11319 ( .A1(n8829), .A2(n8835), .ZN(n8830) );
  INV_X1 U11320 ( .A(n8837), .ZN(n8832) );
  NAND2_X1 U11321 ( .A1(n11309), .A2(n11308), .ZN(n11683) );
  NOR2_X1 U11322 ( .A1(n11683), .A2(n14374), .ZN(n9651) );
  NAND3_X1 U11323 ( .A1(n8832), .A2(n8831), .A3(n9651), .ZN(n8833) );
  AOI22_X1 U11324 ( .A1(n8924), .A2(n14612), .B1(n9230), .B2(n14616), .ZN(
        n8844) );
  INV_X1 U11325 ( .A(n11689), .ZN(n8836) );
  OR2_X1 U11326 ( .A1(n8837), .A2(n8836), .ZN(n13915) );
  NAND2_X1 U11327 ( .A1(n8889), .A2(n11748), .ZN(n14633) );
  NOR2_X1 U11328 ( .A1(n13915), .A2(n14633), .ZN(n12558) );
  INV_X1 U11329 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13958) );
  OR2_X1 U11330 ( .A1(n11608), .A2(n13958), .ZN(n8841) );
  OR2_X1 U11331 ( .A1(n11630), .A2(n9661), .ZN(n8840) );
  INV_X1 U11332 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U11333 ( .A1(n12558), .A2(n13955), .ZN(n8843) );
  OAI211_X1 U11334 ( .C1(n9031), .C2(n9917), .A(n8844), .B(n8843), .ZN(
        P1_U3232) );
  INV_X1 U11335 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n15378) );
  NAND2_X1 U11336 ( .A1(n9676), .A2(n9675), .ZN(n9993) );
  INV_X1 U11337 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U11338 ( .A1(n10717), .A2(n10716), .ZN(n10872) );
  INV_X1 U11339 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8845) );
  NOR2_X1 U11340 ( .A1(n10934), .A2(n8845), .ZN(n8846) );
  OR2_X1 U11341 ( .A1(n11022), .A2(n8846), .ZN(n12614) );
  NAND2_X1 U11342 ( .A1(n11154), .A2(n12614), .ZN(n8850) );
  NAND2_X1 U11343 ( .A1(n6530), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U11344 ( .A1(n6533), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U11345 ( .A1(n11216), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U11346 ( .A1(n12621), .A2(P3_U3897), .ZN(n8851) );
  OAI21_X1 U11347 ( .B1(P3_U3897), .B2(n15378), .A(n8851), .ZN(P3_U3507) );
  INV_X1 U11348 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15379) );
  NAND2_X1 U11349 ( .A1(n10257), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U11350 ( .A1(n10544), .A2(n8852), .ZN(n15010) );
  NAND2_X1 U11351 ( .A1(n11154), .A2(n15010), .ZN(n8856) );
  NAND2_X1 U11352 ( .A1(n6530), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11353 ( .A1(n6531), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11354 ( .A1(n11216), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11355 ( .A1(n10919), .A2(P3_U3897), .ZN(n8857) );
  OAI21_X1 U11356 ( .B1(P3_U3897), .B2(n15379), .A(n8857), .ZN(P3_U3501) );
  NOR2_X1 U11357 ( .A1(n8858), .A2(n8713), .ZN(n8859) );
  MUX2_X1 U11358 ( .A(n8713), .B(n8859), .S(P3_IR_REG_16__SCAN_IN), .Z(n8861)
         );
  INV_X1 U11359 ( .A(n9052), .ZN(n8860) );
  INV_X1 U11360 ( .A(n8862), .ZN(n8863) );
  NAND2_X1 U11361 ( .A1(n9284), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11362 ( .A1(n9286), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U11363 ( .A1(n9036), .A2(n8866), .ZN(n9033) );
  XNOR2_X1 U11364 ( .A(n9035), .B(n9033), .ZN(n11019) );
  INV_X1 U11365 ( .A(n11019), .ZN(n8868) );
  OAI222_X1 U11366 ( .A1(n12782), .A2(P3_U3151), .B1(n13120), .B2(n8868), .C1(
        n8867), .C2(n13115), .ZN(P3_U3279) );
  INV_X1 U11367 ( .A(n10598), .ZN(n8873) );
  INV_X1 U11368 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11369 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  NAND2_X1 U11370 ( .A1(n8871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9310) );
  XNOR2_X1 U11371 ( .A(n9310), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10599) );
  INV_X1 U11372 ( .A(n10599), .ZN(n9598) );
  OAI222_X1 U11373 ( .A1(n11751), .A2(n8872), .B1(n14370), .B2(n8873), .C1(
        P1_U3086), .C2(n9598), .ZN(P1_U3342) );
  OAI222_X1 U11374 ( .A1(n13749), .A2(n8874), .B1(n10417), .B2(n8873), .C1(
        P2_U3088), .C2(n11077), .ZN(P2_U3314) );
  AND2_X4 U11375 ( .A1(n11516), .A2(n9161), .ZN(n11622) );
  NAND2_X1 U11376 ( .A1(n11622), .A2(n7441), .ZN(n8879) );
  OR2_X1 U11377 ( .A1(n11623), .A2(n8876), .ZN(n8877) );
  AND2_X2 U11378 ( .A1(n11307), .A2(n11365), .ZN(n12522) );
  INV_X4 U11379 ( .A(n12522), .ZN(n12551) );
  XNOR2_X1 U11380 ( .A(n8880), .B(n12551), .ZN(n9015) );
  INV_X1 U11381 ( .A(n13955), .ZN(n9028) );
  OAI22_X1 U11382 ( .A1(n12525), .A2(n9028), .B1(n14752), .B2(n12542), .ZN(
        n9013) );
  XNOR2_X1 U11383 ( .A(n9015), .B(n9013), .ZN(n9016) );
  OAI21_X1 U11384 ( .B1(n12522), .B2(n8882), .A(n8881), .ZN(n9017) );
  XOR2_X1 U11385 ( .A(n9016), .B(n9017), .Z(n8894) );
  NAND2_X1 U11386 ( .A1(n11582), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8888) );
  INV_X1 U11387 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9792) );
  OR2_X1 U11388 ( .A1(n11608), .A2(n9792), .ZN(n8887) );
  OR2_X1 U11389 ( .A1(n11630), .A2(n8883), .ZN(n8886) );
  OR2_X1 U11390 ( .A1(n11583), .A2(n8884), .ZN(n8885) );
  NAND4_X2 U11391 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n13954) );
  AOI22_X1 U11392 ( .A1(n12558), .A2(n13954), .B1(n7537), .B2(n14616), .ZN(
        n8893) );
  INV_X1 U11393 ( .A(n9031), .ZN(n8891) );
  AOI22_X1 U11394 ( .A1(n8891), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n8890), .B2(
        n13957), .ZN(n8892) );
  OAI211_X1 U11395 ( .C1(n8894), .C2(n13932), .A(n8893), .B(n8892), .ZN(
        P1_U3222) );
  INV_X1 U11396 ( .A(n8909), .ZN(n8994) );
  INV_X1 U11397 ( .A(n8908), .ZN(n8964) );
  INV_X1 U11398 ( .A(n8906), .ZN(n14829) );
  XNOR2_X1 U11399 ( .A(n8906), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14826) );
  XNOR2_X1 U11400 ( .A(n13271), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n13279) );
  AND2_X1 U11401 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13278) );
  NAND2_X1 U11402 ( .A1(n13279), .A2(n13278), .ZN(n13277) );
  INV_X1 U11403 ( .A(n13271), .ZN(n8905) );
  NAND2_X1 U11404 ( .A1(n8905), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11405 ( .A1(n13277), .A2(n8895), .ZN(n14825) );
  XOR2_X1 U11406 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8908), .Z(n8956) );
  XOR2_X1 U11407 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n8909), .Z(n8984) );
  NOR2_X1 U11408 ( .A1(n8985), .A2(n8984), .ZN(n8983) );
  AOI21_X1 U11409 ( .B1(n8994), .B2(P2_REG1_REG_4__SCAN_IN), .A(n8983), .ZN(
        n8999) );
  XNOR2_X1 U11410 ( .A(n9007), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n8998) );
  MUX2_X1 U11411 ( .A(n8896), .B(P2_REG1_REG_6__SCAN_IN), .S(n8973), .Z(n8902)
         );
  NAND2_X1 U11412 ( .A1(n9324), .A2(n10685), .ZN(n8898) );
  AOI21_X1 U11413 ( .B1(n8899), .B2(n8898), .A(n8897), .ZN(n14846) );
  INV_X1 U11414 ( .A(n14846), .ZN(n8918) );
  OR2_X1 U11415 ( .A1(n8360), .A2(P2_U3088), .ZN(n13757) );
  INV_X1 U11416 ( .A(n13757), .ZN(n8900) );
  NAND2_X1 U11417 ( .A1(n8918), .A2(n8900), .ZN(n8914) );
  INV_X1 U11418 ( .A(n13761), .ZN(n8901) );
  AOI211_X1 U11419 ( .C1(n8903), .C2(n8902), .A(n14858), .B(n8972), .ZN(n8923)
         );
  MUX2_X1 U11420 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7821), .S(n13271), .Z(
        n13274) );
  INV_X1 U11421 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8904) );
  NOR3_X1 U11422 ( .A1(n13274), .A2(n8904), .A3(n7014), .ZN(n13273) );
  AOI21_X1 U11423 ( .B1(n8905), .B2(P2_REG2_REG_1__SCAN_IN), .A(n13273), .ZN(
        n14834) );
  MUX2_X1 U11424 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10166), .S(n8906), .Z(
        n14833) );
  OR2_X1 U11425 ( .A1(n14834), .A2(n14833), .ZN(n14836) );
  NAND2_X1 U11426 ( .A1(n14829), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8959) );
  MUX2_X1 U11427 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n8907), .S(n8908), .Z(n8958)
         );
  AOI21_X1 U11428 ( .B1(n14836), .B2(n8959), .A(n8958), .ZN(n8988) );
  NOR2_X1 U11429 ( .A1(n8908), .A2(n8907), .ZN(n8987) );
  MUX2_X1 U11430 ( .A(n10179), .B(P2_REG2_REG_4__SCAN_IN), .S(n8909), .Z(n8986) );
  OAI21_X1 U11431 ( .B1(n8988), .B2(n8987), .A(n8986), .ZN(n9003) );
  NAND2_X1 U11432 ( .A1(n8994), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9002) );
  MUX2_X1 U11433 ( .A(n8910), .B(P2_REG2_REG_5__SCAN_IN), .S(n9007), .Z(n9001)
         );
  AOI21_X1 U11434 ( .B1(n9003), .B2(n9002), .A(n9001), .ZN(n9000) );
  NOR2_X1 U11435 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  INV_X1 U11436 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10193) );
  MUX2_X1 U11437 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10193), .S(n8973), .Z(n8912) );
  OAI21_X1 U11438 ( .B1(n9000), .B2(n8913), .A(n8912), .ZN(n8970) );
  INV_X1 U11439 ( .A(n8970), .ZN(n8916) );
  NOR3_X1 U11440 ( .A1(n9000), .A2(n8913), .A3(n8912), .ZN(n8915) );
  NOR3_X1 U11441 ( .A1(n8916), .A2(n8915), .A3(n14851), .ZN(n8922) );
  AND2_X1 U11442 ( .A1(n8360), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11443 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9735) );
  AND2_X1 U11444 ( .A1(n14846), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14809) );
  NAND2_X1 U11445 ( .A1(n14809), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8919) );
  OAI211_X1 U11446 ( .C1(n13358), .C2(n8920), .A(n9735), .B(n8919), .ZN(n8921)
         );
  OR3_X1 U11447 ( .A1(n8923), .A2(n8922), .A3(n8921), .ZN(P2_U3220) );
  NAND2_X1 U11448 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13964) );
  MUX2_X1 U11449 ( .A(n13964), .B(n8924), .S(n6526), .Z(n8927) );
  OR2_X1 U11450 ( .A1(n6526), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11451 ( .A1(n8926), .A2(n8925), .ZN(n14709) );
  NAND2_X1 U11452 ( .A1(n14709), .A2(n7491), .ZN(n14712) );
  OAI211_X1 U11453 ( .C1(n8927), .C2(n11748), .A(n13956), .B(n14712), .ZN(
        n13981) );
  XOR2_X1 U11454 ( .A(n8929), .B(n8928), .Z(n8939) );
  INV_X1 U11455 ( .A(n14715), .ZN(n14732) );
  INV_X1 U11456 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U11457 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9712) );
  OAI21_X1 U11458 ( .B1(n14732), .B2(n8930), .A(n9712), .ZN(n8938) );
  MUX2_X1 U11459 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9360), .S(n8936), .Z(n8931)
         );
  NAND3_X1 U11460 ( .A1(n13993), .A2(n8932), .A3(n8931), .ZN(n8933) );
  NAND3_X1 U11461 ( .A1(n14728), .A2(n8934), .A3(n8933), .ZN(n8935) );
  OAI21_X1 U11462 ( .B1(n14020), .B2(n8936), .A(n8935), .ZN(n8937) );
  AOI211_X1 U11463 ( .C1(n14727), .C2(n8939), .A(n8938), .B(n8937), .ZN(n8940)
         );
  NAND2_X1 U11464 ( .A1(n13981), .A2(n8940), .ZN(P1_U3247) );
  NAND2_X1 U11465 ( .A1(n10216), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8942) );
  INV_X1 U11466 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10362) );
  MUX2_X1 U11467 ( .A(n10362), .B(P1_REG2_REG_11__SCAN_IN), .S(n10346), .Z(
        n8941) );
  AOI21_X1 U11468 ( .B1(n8943), .B2(n8942), .A(n8941), .ZN(n9591) );
  NAND3_X1 U11469 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n8944) );
  NAND2_X1 U11470 ( .A1(n8944), .A2(n14728), .ZN(n8954) );
  AOI21_X1 U11471 ( .B1(n10216), .B2(P1_REG1_REG_10__SCAN_IN), .A(n8945), .ZN(
        n8947) );
  INV_X1 U11472 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10227) );
  MUX2_X1 U11473 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10227), .S(n10346), .Z(
        n8946) );
  NAND2_X1 U11474 ( .A1(n8947), .A2(n8946), .ZN(n9588) );
  OAI21_X1 U11475 ( .B1(n8947), .B2(n8946), .A(n9588), .ZN(n8948) );
  NAND2_X1 U11476 ( .A1(n8948), .A2(n14727), .ZN(n8953) );
  NAND2_X1 U11477 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14617)
         );
  INV_X1 U11478 ( .A(n14617), .ZN(n8951) );
  NOR2_X1 U11479 ( .A1(n14020), .A2(n8949), .ZN(n8950) );
  AOI211_X1 U11480 ( .C1(n14715), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8951), .B(
        n8950), .ZN(n8952) );
  OAI211_X1 U11481 ( .C1(n9591), .C2(n8954), .A(n8953), .B(n8952), .ZN(
        P1_U3254) );
  INV_X1 U11482 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8967) );
  AOI211_X1 U11483 ( .C1(n8957), .C2(n8956), .A(n8955), .B(n14858), .ZN(n8962)
         );
  AND3_X1 U11484 ( .A1(n14836), .A2(n8959), .A3(n8958), .ZN(n8960) );
  NOR3_X1 U11485 ( .A1(n14851), .A2(n8988), .A3(n8960), .ZN(n8961) );
  NOR2_X1 U11486 ( .A1(n8962), .A2(n8961), .ZN(n8966) );
  INV_X1 U11487 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U11488 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14903), .ZN(n8963) );
  AOI21_X1 U11489 ( .B1(n14865), .B2(n8964), .A(n8963), .ZN(n8965) );
  OAI211_X1 U11490 ( .C1(n14873), .C2(n8967), .A(n8966), .B(n8965), .ZN(
        P2_U3217) );
  NAND2_X1 U11491 ( .A1(n8973), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U11492 ( .A(n7921), .B(P2_REG2_REG_7__SCAN_IN), .S(n9634), .Z(n8968)
         );
  AOI21_X1 U11493 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n9633) );
  NAND3_X1 U11494 ( .A1(n8970), .A2(n8969), .A3(n8968), .ZN(n8971) );
  INV_X1 U11495 ( .A(n14851), .ZN(n14867) );
  NAND2_X1 U11496 ( .A1(n8971), .A2(n14867), .ZN(n8982) );
  MUX2_X1 U11497 ( .A(n8974), .B(P2_REG1_REG_7__SCAN_IN), .S(n9634), .Z(n8975)
         );
  NOR2_X1 U11498 ( .A1(n6587), .A2(n8975), .ZN(n9628) );
  AOI211_X1 U11499 ( .C1(n6587), .C2(n8975), .A(n14858), .B(n9628), .ZN(n8976)
         );
  INV_X1 U11500 ( .A(n8976), .ZN(n8981) );
  NOR2_X1 U11501 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7922), .ZN(n8979) );
  NOR2_X1 U11502 ( .A1(n13358), .A2(n8977), .ZN(n8978) );
  AOI211_X1 U11503 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n14809), .A(n8979), .B(
        n8978), .ZN(n8980) );
  OAI211_X1 U11504 ( .C1(n9633), .C2(n8982), .A(n8981), .B(n8980), .ZN(
        P2_U3221) );
  AOI211_X1 U11505 ( .C1(n8985), .C2(n8984), .A(n14858), .B(n8983), .ZN(n8992)
         );
  INV_X1 U11506 ( .A(n9003), .ZN(n8990) );
  NOR3_X1 U11507 ( .A1(n8988), .A2(n8987), .A3(n8986), .ZN(n8989) );
  NOR3_X1 U11508 ( .A1(n14851), .A2(n8990), .A3(n8989), .ZN(n8991) );
  NOR2_X1 U11509 ( .A1(n8992), .A2(n8991), .ZN(n8996) );
  AND2_X1 U11510 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8993) );
  AOI21_X1 U11511 ( .B1(n14865), .B2(n8994), .A(n8993), .ZN(n8995) );
  OAI211_X1 U11512 ( .C1(n14873), .C2(n6924), .A(n8996), .B(n8995), .ZN(
        P2_U3218) );
  AOI211_X1 U11513 ( .C1(n8999), .C2(n8998), .A(n14858), .B(n8997), .ZN(n9012)
         );
  INV_X1 U11514 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9010) );
  INV_X1 U11515 ( .A(n9000), .ZN(n9005) );
  NAND3_X1 U11516 ( .A1(n9003), .A2(n9002), .A3(n9001), .ZN(n9004) );
  NAND3_X1 U11517 ( .A1(n9005), .A2(n14867), .A3(n9004), .ZN(n9009) );
  AND2_X1 U11518 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9006) );
  AOI21_X1 U11519 ( .B1(n14865), .B2(n9007), .A(n9006), .ZN(n9008) );
  OAI211_X1 U11520 ( .C1(n14873), .C2(n9010), .A(n9009), .B(n9008), .ZN(n9011)
         );
  OR2_X1 U11521 ( .A1(n9012), .A2(n9011), .ZN(P2_U3219) );
  INV_X1 U11522 ( .A(n9013), .ZN(n9014) );
  AOI22_X1 U11523 ( .A1(n9017), .A2(n9016), .B1(n9015), .B2(n9014), .ZN(n9355)
         );
  INV_X1 U11524 ( .A(n13954), .ZN(n9386) );
  INV_X2 U11525 ( .A(n11623), .ZN(n11613) );
  OAI22_X1 U11526 ( .A1(n12525), .A2(n9386), .B1(n11374), .B2(n12542), .ZN(
        n9352) );
  AOI22_X1 U11527 ( .A1(n7196), .A2(n11372), .B1(n9019), .B2(n13954), .ZN(
        n9020) );
  XNOR2_X1 U11528 ( .A(n9020), .B(n12551), .ZN(n9351) );
  XNOR2_X1 U11529 ( .A(n9355), .B(n9354), .ZN(n9021) );
  NAND2_X1 U11530 ( .A1(n9021), .A2(n14612), .ZN(n9030) );
  INV_X1 U11531 ( .A(n13915), .ZN(n14614) );
  NAND2_X1 U11532 ( .A1(n11582), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9027) );
  OR2_X1 U11533 ( .A1(n11608), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9026) );
  OR2_X1 U11534 ( .A1(n11630), .A2(n9022), .ZN(n9025) );
  OR2_X1 U11535 ( .A1(n11583), .A2(n9023), .ZN(n9024) );
  NAND4_X1 U11536 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(n13953) );
  INV_X1 U11537 ( .A(n13953), .ZN(n11379) );
  OAI22_X1 U11538 ( .A1(n9028), .A2(n14631), .B1(n11379), .B2(n14633), .ZN(
        n9235) );
  AOI22_X1 U11539 ( .A1(n11372), .A2(n14616), .B1(n14614), .B2(n9235), .ZN(
        n9029) );
  OAI211_X1 U11540 ( .C1(n9031), .C2(n9792), .A(n9030), .B(n9029), .ZN(
        P1_U3237) );
  NAND2_X1 U11541 ( .A1(n9052), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9032) );
  XNOR2_X1 U11542 ( .A(n9032), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14529) );
  INV_X1 U11543 ( .A(n14529), .ZN(n12786) );
  INV_X1 U11544 ( .A(n9033), .ZN(n9034) );
  XNOR2_X1 U11545 ( .A(n9471), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U11546 ( .A(n9211), .B(n9210), .ZN(n11160) );
  INV_X1 U11547 ( .A(n11160), .ZN(n9038) );
  OAI222_X1 U11548 ( .A1(P3_U3151), .A2(n12786), .B1(n13115), .B2(n9039), .C1(
        n13120), .C2(n9038), .ZN(P3_U3278) );
  OAI22_X1 U11549 ( .A1(n9040), .A2(n14858), .B1(n14851), .B2(n8904), .ZN(
        n9043) );
  AOI21_X1 U11550 ( .B1(n13380), .B2(n9040), .A(n14865), .ZN(n9041) );
  OAI21_X1 U11551 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14851), .A(n9041), .ZN(
        n9042) );
  MUX2_X1 U11552 ( .A(n9043), .B(n9042), .S(P2_IR_REG_0__SCAN_IN), .Z(n9045)
         );
  INV_X1 U11553 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15441) );
  OAI22_X1 U11554 ( .A1(n14873), .A2(n15441), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9538), .ZN(n9044) );
  OR2_X1 U11555 ( .A1(n9045), .A2(n9044), .ZN(P2_U3214) );
  MUX2_X1 U11556 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12777), .Z(n9084) );
  XNOR2_X1 U11557 ( .A(n9084), .B(n7513), .ZN(n9086) );
  MUX2_X1 U11558 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9051), .Z(n9046) );
  XOR2_X1 U11559 ( .A(n9251), .B(n9046), .Z(n9124) );
  INV_X1 U11560 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9430) );
  INV_X1 U11561 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9562) );
  MUX2_X1 U11562 ( .A(n9430), .B(n9562), .S(n9051), .Z(n9271) );
  INV_X1 U11563 ( .A(n9251), .ZN(n9135) );
  INV_X1 U11564 ( .A(n9046), .ZN(n9047) );
  AOI22_X1 U11565 ( .A1(n9124), .A2(n9276), .B1(n9135), .B2(n9047), .ZN(n9109)
         );
  MUX2_X1 U11566 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n9051), .Z(n9048) );
  XNOR2_X1 U11567 ( .A(n9048), .B(n9069), .ZN(n9110) );
  OAI22_X1 U11568 ( .A1(n9109), .A2(n9110), .B1(n9048), .B2(n9069), .ZN(n9087)
         );
  XOR2_X1 U11569 ( .A(n9086), .B(n9087), .Z(n9083) );
  AND2_X1 U11570 ( .A1(n11302), .A2(P3_U3897), .ZN(n12795) );
  NAND2_X1 U11571 ( .A1(n9056), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9057) );
  MUX2_X1 U11572 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9057), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9059) );
  NAND2_X2 U11573 ( .A1(n9891), .A2(n12034), .ZN(n11936) );
  INV_X1 U11574 ( .A(n9198), .ZN(n9062) );
  OR2_X1 U11575 ( .A1(n11936), .A2(n9062), .ZN(n9060) );
  NAND2_X1 U11576 ( .A1(n10868), .A2(n9060), .ZN(n9077) );
  NAND2_X1 U11577 ( .A1(n9199), .A2(n9061), .ZN(n9405) );
  NAND2_X1 U11578 ( .A1(n9062), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12036) );
  AND2_X1 U11579 ( .A1(n9405), .A2(n12036), .ZN(n9075) );
  OR2_X1 U11580 ( .A1(n9077), .A2(n9075), .ZN(n9068) );
  INV_X1 U11581 ( .A(n11302), .ZN(n12031) );
  MUX2_X1 U11582 ( .A(n9068), .B(n12686), .S(n12031), .Z(n14981) );
  INV_X1 U11583 ( .A(n14981), .ZN(n14543) );
  NAND2_X1 U11584 ( .A1(n12031), .A2(n12710), .ZN(n9195) );
  OR2_X1 U11585 ( .A1(n9068), .A2(n9195), .ZN(n14994) );
  INV_X1 U11586 ( .A(n14994), .ZN(n14554) );
  INV_X1 U11587 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U11588 ( .A1(n9065), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9063) );
  INV_X1 U11589 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15082) );
  AOI21_X1 U11590 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n9065), .A(n9064), .ZN(
        n9113) );
  NAND2_X1 U11591 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n9069), .ZN(n9066) );
  XNOR2_X1 U11592 ( .A(n15260), .B(n9090), .ZN(n9067) );
  NAND2_X1 U11593 ( .A1(n14554), .A2(n9067), .ZN(n9080) );
  OR2_X1 U11594 ( .A1(n9068), .A2(n12710), .ZN(n12791) );
  NAND2_X1 U11595 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n9069), .ZN(n9072) );
  INV_X1 U11596 ( .A(n9069), .ZN(n9483) );
  INV_X1 U11597 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U11598 ( .A1(n9483), .A2(n15129), .B1(P3_REG1_REG_2__SCAN_IN), .B2(
        n9069), .ZN(n9116) );
  NAND2_X1 U11599 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15181), .ZN(n9071) );
  INV_X1 U11600 ( .A(n9071), .ZN(n9268) );
  OR2_X1 U11601 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9071), .ZN(n9070) );
  OAI21_X1 U11602 ( .B1(n9251), .B2(n9268), .A(n9070), .ZN(n9127) );
  INV_X1 U11603 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11604 ( .A1(n9116), .A2(n9115), .ZN(n9114) );
  NAND2_X1 U11605 ( .A1(n9072), .A2(n9114), .ZN(n9096) );
  XNOR2_X1 U11606 ( .A(n9096), .B(n7513), .ZN(n9073) );
  NAND2_X1 U11607 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n9073), .ZN(n9098) );
  OAI21_X1 U11608 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n9073), .A(n9098), .ZN(
        n9074) );
  NAND2_X1 U11609 ( .A1(n14990), .A2(n9074), .ZN(n9079) );
  INV_X1 U11610 ( .A(n9075), .ZN(n9076) );
  INV_X1 U11611 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U11612 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9897), .ZN(n9503) );
  AOI21_X1 U11613 ( .B1(n14987), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n9503), .ZN(
        n9078) );
  NAND3_X1 U11614 ( .A1(n9080), .A2(n9079), .A3(n9078), .ZN(n9081) );
  AOI21_X1 U11615 ( .B1(n7513), .B2(n14543), .A(n9081), .ZN(n9082) );
  OAI21_X1 U11616 ( .B1(n9083), .B2(n14983), .A(n9082), .ZN(P3_U3185) );
  MUX2_X1 U11617 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12777), .Z(n9287) );
  XNOR2_X1 U11618 ( .A(n9287), .B(n9987), .ZN(n9289) );
  INV_X1 U11619 ( .A(n9084), .ZN(n9085) );
  AOI22_X1 U11620 ( .A1(n9087), .A2(n9086), .B1(n7513), .B2(n9085), .ZN(n9138)
         );
  INV_X2 U11621 ( .A(n12710), .ZN(n12777) );
  MUX2_X1 U11622 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12777), .Z(n9088) );
  XOR2_X1 U11623 ( .A(n9668), .B(n9088), .Z(n9139) );
  OAI22_X1 U11624 ( .A1(n9138), .A2(n9139), .B1(n9088), .B2(n9094), .ZN(n9290)
         );
  XOR2_X1 U11625 ( .A(n9289), .B(n9290), .Z(n9108) );
  INV_X1 U11626 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11627 ( .A1(n9094), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9092) );
  INV_X1 U11628 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U11629 ( .A1(n9668), .A2(n9910), .ZN(n9091) );
  NAND2_X1 U11630 ( .A1(n9092), .A2(n9091), .ZN(n9142) );
  XNOR2_X1 U11631 ( .A(n9293), .B(n9292), .ZN(n9093) );
  NAND2_X1 U11632 ( .A1(n14554), .A2(n9093), .ZN(n9105) );
  NAND2_X1 U11633 ( .A1(n9094), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9100) );
  INV_X1 U11634 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9095) );
  MUX2_X1 U11635 ( .A(n9095), .B(P3_REG1_REG_4__SCAN_IN), .S(n9668), .Z(n9145)
         );
  NAND2_X1 U11636 ( .A1(n9097), .A2(n9096), .ZN(n9099) );
  NAND2_X1 U11637 ( .A1(n9145), .A2(n9146), .ZN(n9144) );
  OAI21_X1 U11638 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n9101), .A(n9297), .ZN(
        n9102) );
  NAND2_X1 U11639 ( .A1(n14990), .A2(n9102), .ZN(n9104) );
  NOR2_X1 U11640 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9675), .ZN(n10001) );
  AOI21_X1 U11641 ( .B1(n14987), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10001), .ZN(
        n9103) );
  NAND3_X1 U11642 ( .A1(n9105), .A2(n9104), .A3(n9103), .ZN(n9106) );
  AOI21_X1 U11643 ( .B1(n9987), .B2(n14543), .A(n9106), .ZN(n9107) );
  OAI21_X1 U11644 ( .B1(n9108), .B2(n14983), .A(n9107), .ZN(P3_U3187) );
  XOR2_X1 U11645 ( .A(n9110), .B(n9109), .Z(n9123) );
  AOI21_X1 U11646 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9120) );
  OAI21_X1 U11647 ( .B1(n9116), .B2(n9115), .A(n9114), .ZN(n9117) );
  NAND2_X1 U11648 ( .A1(n14990), .A2(n9117), .ZN(n9119) );
  AOI22_X1 U11649 ( .A1(n14987), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9118) );
  OAI211_X1 U11650 ( .C1(n9120), .C2(n14994), .A(n9119), .B(n9118), .ZN(n9121)
         );
  AOI21_X1 U11651 ( .B1(n9483), .B2(n14543), .A(n9121), .ZN(n9122) );
  OAI21_X1 U11652 ( .B1(n9123), .B2(n14983), .A(n9122), .ZN(P3_U3184) );
  XOR2_X1 U11653 ( .A(n9276), .B(n9124), .Z(n9137) );
  XNOR2_X1 U11654 ( .A(n9125), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11655 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11656 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U11657 ( .A1(n14990), .A2(n9130), .ZN(n9132) );
  AOI22_X1 U11658 ( .A1(n14987), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9131) );
  OAI211_X1 U11659 ( .C1(n9133), .C2(n14994), .A(n9132), .B(n9131), .ZN(n9134)
         );
  AOI21_X1 U11660 ( .B1(n9135), .B2(n14543), .A(n9134), .ZN(n9136) );
  OAI21_X1 U11661 ( .B1(n9137), .B2(n14983), .A(n9136), .ZN(P3_U3183) );
  XOR2_X1 U11662 ( .A(n9139), .B(n9138), .Z(n9154) );
  INV_X1 U11663 ( .A(n9140), .ZN(n9141) );
  AOI21_X1 U11664 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9151) );
  OAI21_X1 U11665 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9147) );
  NAND2_X1 U11666 ( .A1(n14990), .A2(n9147), .ZN(n9150) );
  INV_X1 U11667 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9148) );
  NOR2_X1 U11668 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9148), .ZN(n9684) );
  AOI21_X1 U11669 ( .B1(n14987), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n9684), .ZN(
        n9149) );
  OAI211_X1 U11670 ( .C1(n9151), .C2(n14994), .A(n9150), .B(n9149), .ZN(n9152)
         );
  AOI21_X1 U11671 ( .B1(n9668), .B2(n14543), .A(n9152), .ZN(n9153) );
  OAI21_X1 U11672 ( .B1(n9154), .B2(n14983), .A(n9153), .ZN(P3_U3186) );
  NAND2_X1 U11673 ( .A1(n6530), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U11674 ( .A1(n11154), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11675 ( .A1(n6532), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11676 ( .A1(n9678), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9155) );
  OR2_X1 U11677 ( .A1(n9484), .A2(n9160), .ZN(n9164) );
  OAI211_X1 U11678 ( .C1(n15181), .C2(n10868), .A(n9164), .B(n9163), .ZN(n9432) );
  NAND2_X1 U11679 ( .A1(n15063), .A2(n9564), .ZN(n11826) );
  INV_X1 U11680 ( .A(n11826), .ZN(n11827) );
  NOR2_X1 U11681 ( .A1(n15061), .A2(n11827), .ZN(n11987) );
  NOR2_X1 U11682 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .ZN(
        n9168) );
  NOR4_X1 U11683 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_3__SCAN_IN), .ZN(n9167) );
  NOR4_X1 U11684 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9166) );
  NOR4_X1 U11685 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9165) );
  NAND4_X1 U11686 ( .A1(n9168), .A2(n9167), .A3(n9166), .A4(n9165), .ZN(n9174)
         );
  NOR4_X1 U11687 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9172) );
  NOR4_X1 U11688 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9171) );
  NOR4_X1 U11689 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9170) );
  NOR4_X1 U11690 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n9169) );
  NAND4_X1 U11691 ( .A1(n9172), .A2(n9171), .A3(n9170), .A4(n9169), .ZN(n9173)
         );
  NOR2_X1 U11692 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  NOR2_X1 U11693 ( .A1(n9424), .A2(n9186), .ZN(n9408) );
  NAND2_X1 U11694 ( .A1(n9177), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11695 ( .A1(n11828), .A2(n9690), .ZN(n9180) );
  NAND2_X1 U11696 ( .A1(n9180), .A2(n10134), .ZN(n9185) );
  NAND2_X1 U11697 ( .A1(n9690), .A2(n12034), .ZN(n9182) );
  NAND2_X1 U11698 ( .A1(n6628), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11699 ( .A1(n9182), .A2(n12771), .ZN(n9183) );
  NAND2_X1 U11700 ( .A1(n9183), .A2(n11828), .ZN(n9184) );
  NAND2_X1 U11701 ( .A1(n9185), .A2(n9184), .ZN(n9880) );
  NAND3_X1 U11702 ( .A1(n9408), .A2(n15054), .A3(n9880), .ZN(n9189) );
  NAND2_X1 U11703 ( .A1(n11730), .A2(n9556), .ZN(n9423) );
  NAND2_X1 U11704 ( .A1(n11828), .A2(n9890), .ZN(n12014) );
  NAND2_X1 U11705 ( .A1(n12034), .A2(n12771), .ZN(n9892) );
  OR2_X1 U11706 ( .A1(n12014), .A2(n9892), .ZN(n9406) );
  INV_X1 U11707 ( .A(n9406), .ZN(n9187) );
  NAND2_X1 U11708 ( .A1(n9409), .A2(n9187), .ZN(n9188) );
  NAND2_X1 U11709 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  INV_X1 U11710 ( .A(n9405), .ZN(n9420) );
  NAND2_X1 U11711 ( .A1(n9678), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U11712 ( .A1(n6530), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11713 ( .A1(n6531), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9192) );
  NAND2_X1 U11714 ( .A1(n11154), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11715 ( .A1(n6534), .A2(n9195), .ZN(n9883) );
  AND2_X1 U11716 ( .A1(n9690), .A2(n12023), .ZN(n12030) );
  INV_X1 U11717 ( .A(n12030), .ZN(n9554) );
  OR2_X1 U11718 ( .A1(n9554), .A2(n11936), .ZN(n9401) );
  OR2_X1 U11719 ( .A1(n9405), .A2(n9401), .ZN(n9404) );
  INV_X1 U11720 ( .A(n9404), .ZN(n12032) );
  AND2_X1 U11721 ( .A1(n9883), .A2(n12032), .ZN(n9196) );
  NAND2_X1 U11722 ( .A1(n9409), .A2(n9196), .ZN(n12646) );
  INV_X1 U11723 ( .A(n12646), .ZN(n12663) );
  OR2_X1 U11724 ( .A1(n9408), .A2(n15056), .ZN(n9197) );
  NOR2_X1 U11725 ( .A1(n9405), .A2(n15054), .ZN(n9429) );
  AOI22_X1 U11726 ( .A1(n12685), .A2(n12663), .B1(n12648), .B2(n9432), .ZN(
        n9207) );
  INV_X1 U11727 ( .A(n9880), .ZN(n9202) );
  OR2_X1 U11728 ( .A1(n9409), .A2(n9406), .ZN(n9201) );
  OR2_X1 U11729 ( .A1(n11936), .A2(n12030), .ZN(n9426) );
  AND3_X1 U11730 ( .A1(n9199), .A2(n9198), .A3(n9426), .ZN(n9200) );
  OAI211_X1 U11731 ( .C1(n9408), .C2(n9202), .A(n9201), .B(n9200), .ZN(n9203)
         );
  NAND2_X1 U11732 ( .A1(n9203), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9205) );
  OR2_X1 U11733 ( .A1(n9409), .A2(n9404), .ZN(n9204) );
  NAND2_X2 U11734 ( .A1(n9205), .A2(n9204), .ZN(n12670) );
  OR2_X1 U11735 ( .A1(n12670), .A2(P3_U3151), .ZN(n9546) );
  NAND2_X1 U11736 ( .A1(n9546), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9206) );
  OAI211_X1 U11737 ( .C1(n11987), .C2(n12672), .A(n9207), .B(n9206), .ZN(
        P3_U3172) );
  NAND2_X1 U11738 ( .A1(n9208), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9209) );
  XNOR2_X1 U11739 ( .A(n9209), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14542) );
  INV_X1 U11740 ( .A(n14542), .ZN(n12781) );
  NAND2_X1 U11741 ( .A1(n9471), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11742 ( .A1(n15420), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9342) );
  INV_X1 U11743 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U11744 ( .A1(n9626), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U11745 ( .A1(n9342), .A2(n9213), .ZN(n9214) );
  NAND2_X1 U11746 ( .A1(n9215), .A2(n9214), .ZN(n9216) );
  NAND2_X1 U11747 ( .A1(n9343), .A2(n9216), .ZN(n11164) );
  OAI222_X1 U11748 ( .A1(P3_U3151), .A2(n12781), .B1(n13115), .B2(n15396), 
        .C1(n13120), .C2(n11164), .ZN(P3_U3277) );
  NAND3_X1 U11749 ( .A1(n11689), .A2(n9218), .A3(n9217), .ZN(n9219) );
  OR2_X1 U11750 ( .A1(n9220), .A2(n9219), .ZN(n9244) );
  INV_X1 U11751 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9229) );
  INV_X1 U11752 ( .A(n11307), .ZN(n9221) );
  NAND2_X1 U11753 ( .A1(n9221), .A2(n9746), .ZN(n9222) );
  NAND2_X1 U11754 ( .A1(n12551), .A2(n9222), .ZN(n14637) );
  OR2_X1 U11755 ( .A1(n11331), .A2(n14635), .ZN(n14764) );
  NAND2_X1 U11756 ( .A1(n11633), .A2(n11309), .ZN(n9224) );
  NAND2_X1 U11757 ( .A1(n14374), .A2(n11352), .ZN(n9223) );
  NAND2_X1 U11758 ( .A1(n13957), .A2(n9919), .ZN(n9225) );
  NAND2_X1 U11759 ( .A1(n11363), .A2(n9225), .ZN(n11366) );
  OAI21_X1 U11760 ( .B1(n14796), .B2(n14494), .A(n11366), .ZN(n9226) );
  NAND2_X1 U11761 ( .A1(n13955), .A2(n14222), .ZN(n9918) );
  OAI211_X1 U11762 ( .C1(n9227), .C2(n9919), .A(n9226), .B(n9918), .ZN(n14347)
         );
  NAND2_X1 U11763 ( .A1(n6528), .A2(n14347), .ZN(n9228) );
  OAI21_X1 U11764 ( .B1(n6528), .B2(n9229), .A(n9228), .ZN(P1_U3459) );
  INV_X1 U11765 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9242) );
  AND2_X1 U11766 ( .A1(n13957), .A2(n9230), .ZN(n9650) );
  OR2_X1 U11767 ( .A1(n13955), .A2(n7537), .ZN(n9231) );
  INV_X1 U11768 ( .A(n11645), .ZN(n9232) );
  OAI21_X1 U11769 ( .B1(n9233), .B2(n9232), .A(n9384), .ZN(n9798) );
  INV_X1 U11770 ( .A(n9798), .ZN(n9240) );
  AND2_X1 U11771 ( .A1(n13955), .A2(n14752), .ZN(n11369) );
  INV_X1 U11772 ( .A(n11369), .ZN(n11364) );
  NAND2_X1 U11773 ( .A1(n9234), .A2(n11645), .ZN(n9388) );
  OAI21_X1 U11774 ( .B1(n9234), .B2(n11645), .A(n9388), .ZN(n9236) );
  AOI21_X1 U11775 ( .B1(n9236), .B2(n14494), .A(n9235), .ZN(n9800) );
  NAND2_X1 U11776 ( .A1(n9652), .A2(n11372), .ZN(n9237) );
  NAND2_X1 U11777 ( .A1(n9237), .A2(n8808), .ZN(n9238) );
  NOR2_X1 U11778 ( .A1(n9395), .A2(n9238), .ZN(n9794) );
  AOI21_X1 U11779 ( .B1(n14759), .B2(n11372), .A(n9794), .ZN(n9239) );
  OAI211_X1 U11780 ( .C1(n9240), .C2(n14663), .A(n9800), .B(n9239), .ZN(n9245)
         );
  NAND2_X1 U11781 ( .A1(n9245), .A2(n6528), .ZN(n9241) );
  OAI21_X1 U11782 ( .B1(n6528), .B2(n9242), .A(n9241), .ZN(P1_U3465) );
  NAND2_X1 U11783 ( .A1(n9245), .A2(n14808), .ZN(n9246) );
  OAI21_X1 U11784 ( .B1(n14808), .B2(n8884), .A(n9246), .ZN(P1_U3530) );
  OR2_X1 U11785 ( .A1(n9484), .A2(n9247), .ZN(n9250) );
  OR2_X2 U11786 ( .A1(n11730), .A2(n12014), .ZN(n9255) );
  NAND2_X1 U11787 ( .A1(n11828), .A2(n12771), .ZN(n9253) );
  NAND2_X1 U11788 ( .A1(n9253), .A2(n9690), .ZN(n9254) );
  INV_X1 U11789 ( .A(n15074), .ZN(n9885) );
  NAND2_X1 U11790 ( .A1(n12685), .A2(n9885), .ZN(n11831) );
  NAND2_X1 U11791 ( .A1(n15066), .A2(n9489), .ZN(n9256) );
  NAND2_X1 U11792 ( .A1(n9875), .A2(n9256), .ZN(n9257) );
  INV_X1 U11793 ( .A(n15061), .ZN(n9258) );
  NAND3_X1 U11794 ( .A1(n9258), .A2(n15067), .A3(n11786), .ZN(n9259) );
  OAI211_X1 U11795 ( .C1(n9260), .C2(n15066), .A(n9479), .B(n9259), .ZN(n9261)
         );
  NAND2_X1 U11796 ( .A1(n9261), .A2(n12651), .ZN(n9267) );
  NAND2_X1 U11797 ( .A1(n15064), .A2(n12663), .ZN(n9264) );
  NOR2_X1 U11798 ( .A1(n9883), .A2(n9404), .ZN(n9262) );
  NAND2_X1 U11799 ( .A1(n15063), .A2(n12643), .ZN(n9263) );
  OAI211_X1 U11800 ( .C1(n9885), .C2(n12666), .A(n9264), .B(n9263), .ZN(n9265)
         );
  AOI21_X1 U11801 ( .B1(n9546), .B2(P3_REG3_REG_1__SCAN_IN), .A(n9265), .ZN(
        n9266) );
  NAND2_X1 U11802 ( .A1(n9267), .A2(n9266), .ZN(P3_U3162) );
  NAND3_X1 U11803 ( .A1(n14994), .A2(n12791), .A3(n14983), .ZN(n9275) );
  NAND2_X1 U11804 ( .A1(n14990), .A2(n9268), .ZN(n9270) );
  AOI22_X1 U11805 ( .A1(n14987), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9269) );
  OAI211_X1 U11806 ( .C1(n6695), .C2(n14994), .A(n9270), .B(n9269), .ZN(n9274)
         );
  NOR2_X1 U11807 ( .A1(n14983), .A2(n9271), .ZN(n9272) );
  AOI211_X1 U11808 ( .C1(n9276), .C2(n9275), .A(n9274), .B(n9273), .ZN(n9277)
         );
  INV_X1 U11809 ( .A(n9277), .ZN(P3_U3182) );
  INV_X1 U11810 ( .A(n11447), .ZN(n9285) );
  NAND2_X1 U11811 ( .A1(n7199), .A2(n9278), .ZN(n9415) );
  OR2_X1 U11812 ( .A1(n9415), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11813 ( .A1(n9280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9279) );
  MUX2_X1 U11814 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9279), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9283) );
  INV_X1 U11815 ( .A(n9280), .ZN(n9282) );
  NAND2_X1 U11816 ( .A1(n9282), .A2(n9281), .ZN(n9472) );
  NAND2_X1 U11817 ( .A1(n9283), .A2(n9472), .ZN(n10642) );
  OAI222_X1 U11818 ( .A1(n14372), .A2(n9284), .B1(n14370), .B2(n9285), .C1(
        n10642), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U11819 ( .A(n13345), .ZN(n11085) );
  OAI222_X1 U11820 ( .A1(n13764), .A2(n9286), .B1(n13766), .B2(n9285), .C1(
        n11085), .C2(P2_U3088), .ZN(P2_U3311) );
  MUX2_X1 U11821 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12777), .Z(n9435) );
  XNOR2_X1 U11822 ( .A(n9435), .B(n10115), .ZN(n9436) );
  INV_X1 U11823 ( .A(n9287), .ZN(n9288) );
  AOI22_X1 U11824 ( .A1(n9290), .A2(n9289), .B1(n9987), .B2(n9288), .ZN(n9437)
         );
  XOR2_X1 U11825 ( .A(n9436), .B(n9437), .Z(n9308) );
  NAND2_X1 U11826 ( .A1(n10115), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9438) );
  OR2_X1 U11827 ( .A1(n10115), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9294) );
  OAI21_X1 U11828 ( .B1(n7058), .B2(n6694), .A(n9439), .ZN(n9306) );
  INV_X1 U11829 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U11830 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15331), .ZN(n10247) );
  AOI21_X1 U11831 ( .B1(n14987), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10247), .ZN(
        n9304) );
  NAND2_X1 U11832 ( .A1(n9296), .A2(n9295), .ZN(n9298) );
  INV_X1 U11833 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9299) );
  MUX2_X1 U11834 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n9299), .S(n10115), .Z(n9300) );
  NAND2_X1 U11835 ( .A1(n9300), .A2(n9301), .ZN(n9440) );
  OAI21_X1 U11836 ( .B1(n9301), .B2(n9300), .A(n9440), .ZN(n9302) );
  NAND2_X1 U11837 ( .A1(n14990), .A2(n9302), .ZN(n9303) );
  OAI211_X1 U11838 ( .C1(n14981), .C2(n10115), .A(n9304), .B(n9303), .ZN(n9305) );
  AOI21_X1 U11839 ( .B1(n9306), .B2(n14554), .A(n9305), .ZN(n9307) );
  OAI21_X1 U11840 ( .B1(n9308), .B2(n14983), .A(n9307), .ZN(P3_U3188) );
  INV_X1 U11841 ( .A(n10732), .ZN(n9314) );
  INV_X1 U11842 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11843 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND2_X1 U11844 ( .A1(n9311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9312) );
  XNOR2_X1 U11845 ( .A(n9312), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10733) );
  INV_X1 U11846 ( .A(n10733), .ZN(n9698) );
  OAI222_X1 U11847 ( .A1(n14372), .A2(n9313), .B1(n14370), .B2(n9314), .C1(
        n9698), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U11848 ( .A(n11078), .ZN(n13313) );
  OAI222_X1 U11849 ( .A1(n13764), .A2(n9315), .B1(n13766), .B2(n9314), .C1(
        n13313), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U11850 ( .A1(n13269), .A2(n9574), .ZN(n9371) );
  NAND2_X1 U11851 ( .A1(n9450), .A2(n9574), .ZN(n9464) );
  NAND2_X1 U11852 ( .A1(n12356), .A2(n12041), .ZN(n9316) );
  NAND2_X1 U11853 ( .A1(n9464), .A2(n9316), .ZN(n9320) );
  INV_X1 U11854 ( .A(n9320), .ZN(n9318) );
  INV_X1 U11855 ( .A(n9378), .ZN(n9319) );
  AOI21_X1 U11856 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9341) );
  NOR2_X1 U11857 ( .A1(n14953), .A2(n9324), .ZN(n9325) );
  INV_X1 U11858 ( .A(n14912), .ZN(n9327) );
  INV_X1 U11859 ( .A(n14915), .ZN(n9326) );
  NAND3_X1 U11860 ( .A1(n9327), .A2(n9326), .A3(n9460), .ZN(n9328) );
  NAND2_X1 U11861 ( .A1(n9328), .A2(n9459), .ZN(n9331) );
  AND3_X1 U11862 ( .A1(n9461), .A2(n9329), .A3(n10685), .ZN(n9330) );
  NAND2_X1 U11863 ( .A1(n9331), .A2(n9330), .ZN(n9579) );
  NOR2_X1 U11864 ( .A1(n9579), .A2(P2_U3088), .ZN(n9465) );
  INV_X1 U11865 ( .A(n9465), .ZN(n9335) );
  INV_X1 U11866 ( .A(n12304), .ZN(n9332) );
  INV_X1 U11867 ( .A(n14811), .ZN(n13235) );
  NAND2_X1 U11868 ( .A1(n12042), .A2(n13231), .ZN(n9334) );
  INV_X2 U11869 ( .A(n13193), .ZN(n13230) );
  NAND2_X1 U11870 ( .A1(n13267), .A2(n13230), .ZN(n9333) );
  NAND2_X1 U11871 ( .A1(n9334), .A2(n9333), .ZN(n9454) );
  AOI22_X1 U11872 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n9335), .B1(n13235), .B2(
        n9454), .ZN(n9340) );
  INV_X1 U11873 ( .A(n9336), .ZN(n9338) );
  INV_X1 U11874 ( .A(n14900), .ZN(n9337) );
  OAI21_X2 U11875 ( .B1(n9338), .B2(n9337), .A(n13595), .ZN(n14818) );
  NAND2_X1 U11876 ( .A1(n14818), .A2(n12053), .ZN(n9339) );
  OAI211_X1 U11877 ( .C1(n9341), .C2(n14813), .A(n9340), .B(n9339), .ZN(
        P2_U3194) );
  INV_X1 U11878 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U11879 ( .A1(n9720), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9688) );
  INV_X1 U11880 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U11881 ( .A1(n9722), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9344) );
  OR2_X1 U11882 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U11883 ( .A1(n9689), .A2(n9347), .ZN(n11174) );
  INV_X1 U11884 ( .A(SI_19_), .ZN(n11176) );
  OAI222_X1 U11885 ( .A1(n13120), .A2(n11174), .B1(n13122), .B2(n11176), .C1(
        P3_U3151), .C2(n12023), .ZN(P3_U3276) );
  OR2_X1 U11886 ( .A1(n9348), .A2(n11496), .ZN(n9349) );
  AOI22_X1 U11887 ( .A1(n7196), .A2(n11380), .B1(n9019), .B2(n13953), .ZN(
        n9350) );
  XNOR2_X1 U11888 ( .A(n9350), .B(n12551), .ZN(n9707) );
  AOI22_X1 U11889 ( .A1(n12553), .A2(n13953), .B1(n12554), .B2(n11380), .ZN(
        n9706) );
  XNOR2_X1 U11890 ( .A(n9707), .B(n9706), .ZN(n9357) );
  INV_X1 U11891 ( .A(n9351), .ZN(n9353) );
  AOI211_X1 U11892 ( .C1(n9357), .C2(n9356), .A(n13932), .B(n9711), .ZN(n9370)
         );
  INV_X1 U11893 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U11894 ( .A1(n6963), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9364) );
  INV_X1 U11895 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9359) );
  OR2_X1 U11896 ( .A1(n11607), .A2(n9359), .ZN(n9363) );
  XNOR2_X1 U11897 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10005) );
  OR2_X1 U11898 ( .A1(n11608), .A2(n10005), .ZN(n9362) );
  OR2_X1 U11899 ( .A1(n11630), .A2(n9360), .ZN(n9361) );
  OR2_X1 U11900 ( .A1(n11386), .A2(n14633), .ZN(n9366) );
  NAND2_X1 U11901 ( .A1(n13954), .A2(n14221), .ZN(n9365) );
  NAND2_X1 U11902 ( .A1(n9366), .A2(n9365), .ZN(n9392) );
  AOI22_X1 U11903 ( .A1(n14614), .A2(n9392), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n9368) );
  NAND2_X1 U11904 ( .A1(n14616), .A2(n11380), .ZN(n9367) );
  OAI211_X1 U11905 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14620), .A(n9368), .B(
        n9367), .ZN(n9369) );
  OR2_X1 U11906 ( .A1(n9370), .A2(n9369), .ZN(P1_U3218) );
  NAND2_X1 U11907 ( .A1(n9376), .A2(n9371), .ZN(n9372) );
  NAND2_X1 U11908 ( .A1(n9378), .A2(n9372), .ZN(n9373) );
  NAND2_X1 U11909 ( .A1(n13267), .A2(n9574), .ZN(n9571) );
  XNOR2_X1 U11910 ( .A(n9570), .B(n9571), .ZN(n9377) );
  INV_X1 U11911 ( .A(n13266), .ZN(n9577) );
  OAI22_X1 U11912 ( .A1(n6940), .A2(n13191), .B1(n9577), .B2(n13193), .ZN(
        n10164) );
  INV_X1 U11913 ( .A(n10164), .ZN(n9374) );
  OAI22_X1 U11914 ( .A1(n9374), .A2(n14811), .B1(n9465), .B2(n14827), .ZN(
        n9375) );
  AOI21_X1 U11915 ( .B1(n7852), .B2(n14818), .A(n9375), .ZN(n9382) );
  INV_X1 U11916 ( .A(n9574), .ZN(n12345) );
  OAI22_X1 U11917 ( .A1(n13213), .A2(n6940), .B1(n9376), .B2(n14813), .ZN(
        n9380) );
  INV_X1 U11918 ( .A(n9377), .ZN(n9379) );
  NAND3_X1 U11919 ( .A1(n9380), .A2(n9379), .A3(n9378), .ZN(n9381) );
  OAI211_X1 U11920 ( .C1(n14813), .C2(n11742), .A(n9382), .B(n9381), .ZN(
        P2_U3209) );
  NAND2_X1 U11921 ( .A1(n9386), .A2(n11374), .ZN(n9383) );
  NAND2_X1 U11922 ( .A1(n9384), .A2(n9383), .ZN(n9385) );
  XNOR2_X1 U11923 ( .A(n11380), .B(n13953), .ZN(n11646) );
  INV_X1 U11924 ( .A(n11646), .ZN(n9389) );
  NAND2_X1 U11925 ( .A1(n9385), .A2(n9389), .ZN(n9511) );
  OAI21_X1 U11926 ( .B1(n9385), .B2(n9389), .A(n9511), .ZN(n9393) );
  INV_X1 U11927 ( .A(n9393), .ZN(n14740) );
  INV_X1 U11928 ( .A(n14496), .ZN(n9394) );
  NAND2_X1 U11929 ( .A1(n9386), .A2(n11372), .ZN(n9387) );
  NAND2_X1 U11930 ( .A1(n9388), .A2(n9387), .ZN(n9524) );
  XNOR2_X1 U11931 ( .A(n9524), .B(n9389), .ZN(n9390) );
  NOR2_X1 U11932 ( .A1(n9390), .A2(n14629), .ZN(n9391) );
  AOI211_X1 U11933 ( .C1(n9394), .C2(n9393), .A(n9392), .B(n9391), .ZN(n14746)
         );
  INV_X1 U11934 ( .A(n9395), .ZN(n9396) );
  AOI211_X1 U11935 ( .C1(n11380), .C2(n9396), .A(n14674), .B(n9516), .ZN(
        n14744) );
  AOI21_X1 U11936 ( .B1(n14759), .B2(n11380), .A(n14744), .ZN(n9397) );
  OAI211_X1 U11937 ( .C1(n14740), .C2(n14764), .A(n14746), .B(n9397), .ZN(
        n9399) );
  NAND2_X1 U11938 ( .A1(n9399), .A2(n14808), .ZN(n9398) );
  OAI21_X1 U11939 ( .B1(n14808), .B2(n9023), .A(n9398), .ZN(P1_U3531) );
  INV_X1 U11940 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U11941 ( .A1(n9399), .A2(n6528), .ZN(n9400) );
  OAI21_X1 U11942 ( .B1(n6528), .B2(n15363), .A(n9400), .ZN(P1_U3468) );
  INV_X1 U11943 ( .A(n9401), .ZN(n9402) );
  NOR3_X1 U11944 ( .A1(n11987), .A2(n15073), .A3(n9402), .ZN(n9403) );
  AOI21_X1 U11945 ( .B1(n15065), .B2(n12685), .A(n9403), .ZN(n9561) );
  OAI21_X1 U11946 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9407) );
  NAND2_X1 U11947 ( .A1(n9408), .A2(n9407), .ZN(n9411) );
  NAND3_X1 U11948 ( .A1(n9409), .A2(n9420), .A3(n9880), .ZN(n9410) );
  OR2_X1 U11949 ( .A1(n15125), .A2(n15054), .ZN(n13049) );
  INV_X1 U11950 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9412) );
  OAI22_X1 U11951 ( .A1(n9564), .A2(n13049), .B1(n15127), .B2(n9412), .ZN(
        n9413) );
  INV_X1 U11952 ( .A(n9413), .ZN(n9414) );
  OAI21_X1 U11953 ( .B1(n9561), .B2(n15125), .A(n9414), .ZN(P3_U3390) );
  INV_X1 U11954 ( .A(n10737), .ZN(n9418) );
  NAND2_X1 U11955 ( .A1(n9415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9416) );
  XNOR2_X1 U11956 ( .A(n9416), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14725) );
  INV_X1 U11957 ( .A(n14725), .ZN(n10488) );
  OAI222_X1 U11958 ( .A1(n14372), .A2(n9417), .B1(n14370), .B2(n9418), .C1(
        n10488), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U11959 ( .A(n13328), .ZN(n11081) );
  OAI222_X1 U11960 ( .A1(n13764), .A2(n9419), .B1(n13766), .B2(n9418), .C1(
        n11081), .C2(P2_U3088), .ZN(P2_U3312) );
  AND2_X1 U11961 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  NOR2_X1 U11962 ( .A1(n12771), .A2(n10134), .ZN(n9552) );
  NAND2_X1 U11963 ( .A1(n9890), .A2(n9552), .ZN(n9881) );
  NAND2_X1 U11964 ( .A1(n11936), .A2(n9881), .ZN(n9425) );
  INV_X1 U11965 ( .A(n9425), .ZN(n9427) );
  AND2_X1 U11966 ( .A1(n9426), .A2(n9425), .ZN(n9558) );
  MUX2_X1 U11967 ( .A(n9427), .B(n9558), .S(n9556), .Z(n9428) );
  NAND2_X1 U11968 ( .A1(n9560), .A2(n9428), .ZN(n9431) );
  MUX2_X1 U11969 ( .A(n9430), .B(n9561), .S(n15080), .Z(n9434) );
  INV_X2 U11970 ( .A(n15040), .ZN(n15075) );
  AOI22_X1 U11971 ( .A1(n15038), .A2(n9432), .B1(n15075), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11972 ( .A1(n9434), .A2(n9433), .ZN(P3_U3233) );
  MUX2_X1 U11973 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12777), .Z(n9602) );
  INV_X1 U11974 ( .A(n9612), .ZN(n10263) );
  XNOR2_X1 U11975 ( .A(n9602), .B(n10263), .ZN(n9604) );
  OAI22_X1 U11976 ( .A1(n9437), .A2(n9436), .B1(n9435), .B2(n10115), .ZN(n9605) );
  XOR2_X1 U11977 ( .A(n9604), .B(n9605), .Z(n9449) );
  INV_X1 U11978 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9608) );
  XNOR2_X1 U11979 ( .A(n9608), .B(n9607), .ZN(n9447) );
  NAND2_X1 U11980 ( .A1(n10115), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9441) );
  OAI21_X1 U11981 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n9442), .A(n9613), .ZN(
        n9443) );
  NAND2_X1 U11982 ( .A1(n9443), .A2(n14990), .ZN(n9445) );
  AND2_X1 U11983 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10339) );
  AOI21_X1 U11984 ( .B1(n14987), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10339), .ZN(
        n9444) );
  OAI211_X1 U11985 ( .C1(n14981), .C2(n9612), .A(n9445), .B(n9444), .ZN(n9446)
         );
  AOI21_X1 U11986 ( .B1(n9447), .B2(n14554), .A(n9446), .ZN(n9448) );
  OAI21_X1 U11987 ( .B1(n9449), .B2(n14983), .A(n9448), .ZN(P3_U3189) );
  XNOR2_X1 U11988 ( .A(n12263), .B(n9450), .ZN(n10095) );
  INV_X1 U11989 ( .A(n14953), .ZN(n14946) );
  OAI211_X1 U11990 ( .C1(n9451), .C2(n12041), .A(n13557), .B(n10168), .ZN(
        n10091) );
  OAI21_X1 U11991 ( .B1(n9451), .B2(n14946), .A(n10091), .ZN(n9458) );
  OAI21_X1 U11992 ( .B1(n12263), .B2(n9453), .A(n9452), .ZN(n9455) );
  AOI21_X1 U11993 ( .B1(n9455), .B2(n14892), .A(n9454), .ZN(n9457) );
  INV_X1 U11994 ( .A(n10068), .ZN(n14960) );
  NAND2_X1 U11995 ( .A1(n10095), .A2(n14960), .ZN(n9456) );
  NAND2_X1 U11996 ( .A1(n9457), .A2(n9456), .ZN(n10092) );
  AOI211_X1 U11997 ( .C1(n14943), .C2(n10095), .A(n9458), .B(n10092), .ZN(
        n14920) );
  AND3_X1 U11998 ( .A1(n9460), .A2(n14915), .A3(n9459), .ZN(n10078) );
  NAND2_X1 U11999 ( .A1(n9461), .A2(n14916), .ZN(n10075) );
  NOR2_X1 U12000 ( .A1(n14912), .A2(n10075), .ZN(n9462) );
  NAND2_X1 U12001 ( .A1(n14970), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9463) );
  OAI21_X1 U12002 ( .B1(n14920), .B2(n14970), .A(n9463), .ZN(P2_U3500) );
  INV_X1 U12003 ( .A(n13213), .ZN(n13205) );
  AOI22_X1 U12004 ( .A1(n13205), .A2(n12042), .B1(n9467), .B2(n13227), .ZN(
        n9470) );
  INV_X1 U12005 ( .A(n9464), .ZN(n9469) );
  NAND2_X1 U12006 ( .A1(n13269), .A2(n13230), .ZN(n9534) );
  OAI22_X1 U12007 ( .A1(n9465), .A2(n9538), .B1(n14811), .B2(n9534), .ZN(n9466) );
  AOI21_X1 U12008 ( .B1(n9467), .B2(n14818), .A(n9466), .ZN(n9468) );
  OAI21_X1 U12009 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(P2_U3204) );
  INV_X1 U12010 ( .A(n11453), .ZN(n9475) );
  OAI222_X1 U12011 ( .A1(P2_U3088), .A2(n13364), .B1(n13766), .B2(n9475), .C1(
        n9471), .C2(n13749), .ZN(P2_U3310) );
  NAND2_X1 U12012 ( .A1(n9472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9473) );
  MUX2_X1 U12013 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9473), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9474) );
  AND2_X1 U12014 ( .A1(n9624), .A2(n9474), .ZN(n11454) );
  INV_X1 U12015 ( .A(n11454), .ZN(n10832) );
  OAI222_X1 U12016 ( .A1(n14372), .A2(n9476), .B1(n14370), .B2(n9475), .C1(
        n10832), .C2(P1_U3086), .ZN(P1_U3338) );
  XNOR2_X1 U12017 ( .A(n9885), .B(n11789), .ZN(n9477) );
  INV_X1 U12018 ( .A(n15064), .ZN(n9887) );
  OR2_X1 U12019 ( .A1(n11198), .A2(n9480), .ZN(n9482) );
  OR2_X1 U12020 ( .A1(n9484), .A2(SI_2_), .ZN(n9481) );
  OAI211_X1 U12021 ( .C1(n9483), .C2(n10868), .A(n9482), .B(n9481), .ZN(n9876)
         );
  XNOR2_X1 U12022 ( .A(n9876), .B(n11789), .ZN(n9494) );
  XNOR2_X1 U12023 ( .A(n9887), .B(n9494), .ZN(n9544) );
  OR2_X1 U12024 ( .A1(n9484), .A2(SI_3_), .ZN(n9488) );
  OR2_X1 U12025 ( .A1(n11198), .A2(n9485), .ZN(n9487) );
  OR2_X1 U12026 ( .A1(n10868), .A2(n7513), .ZN(n9486) );
  NAND2_X1 U12027 ( .A1(n6530), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U12028 ( .A1(n11154), .A2(n9897), .ZN(n9492) );
  NAND2_X1 U12029 ( .A1(n6531), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U12030 ( .A1(n9678), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9490) );
  XNOR2_X1 U12031 ( .A(n9664), .B(n15047), .ZN(n9496) );
  INV_X1 U12032 ( .A(n9494), .ZN(n9495) );
  NAND2_X1 U12033 ( .A1(n9495), .A2(n9887), .ZN(n9497) );
  NAND2_X1 U12034 ( .A1(n9665), .A2(n12651), .ZN(n9509) );
  AOI21_X1 U12035 ( .B1(n9542), .B2(n9497), .A(n9496), .ZN(n9508) );
  NAND2_X1 U12036 ( .A1(n6530), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9502) );
  AND2_X1 U12037 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9498) );
  OR2_X1 U12038 ( .A1(n9498), .A2(n9676), .ZN(n9912) );
  NAND2_X1 U12039 ( .A1(n11154), .A2(n9912), .ZN(n9501) );
  NAND2_X1 U12040 ( .A1(n6533), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U12041 ( .A1(n11216), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9499) );
  AOI21_X1 U12042 ( .B1(n15064), .B2(n12643), .A(n9503), .ZN(n9505) );
  NAND2_X1 U12043 ( .A1(n12648), .A2(n9903), .ZN(n9504) );
  OAI211_X1 U12044 ( .C1(n11847), .C2(n12646), .A(n9505), .B(n9504), .ZN(n9506) );
  AOI21_X1 U12045 ( .B1(n9897), .B2(n12670), .A(n9506), .ZN(n9507) );
  OAI21_X1 U12046 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(P3_U3158) );
  NAND2_X1 U12047 ( .A1(n14737), .A2(n11379), .ZN(n9510) );
  NAND2_X1 U12048 ( .A1(n9512), .A2(n11622), .ZN(n9515) );
  AOI22_X1 U12049 ( .A1(n11613), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11455), 
        .B2(n9513), .ZN(n9514) );
  XNOR2_X1 U12050 ( .A(n7324), .B(n11386), .ZN(n11649) );
  XNOR2_X1 U12051 ( .A(n6932), .B(n11649), .ZN(n10012) );
  OAI22_X1 U12052 ( .A1(n10008), .A2(n14674), .B1(n11385), .B2(n14793), .ZN(
        n9527) );
  AOI21_X1 U12053 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9517) );
  NOR2_X1 U12054 ( .A1(n9517), .A2(n9752), .ZN(n9827) );
  NAND2_X1 U12055 ( .A1(n11489), .A2(n9827), .ZN(n9523) );
  OR2_X1 U12056 ( .A1(n11583), .A2(n9518), .ZN(n9522) );
  INV_X1 U12057 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9519) );
  OR2_X1 U12058 ( .A1(n11607), .A2(n9519), .ZN(n9521) );
  OR2_X1 U12059 ( .A1(n11630), .A2(n9760), .ZN(n9520) );
  NAND4_X1 U12060 ( .A1(n9523), .A2(n9522), .A3(n9521), .A4(n9520), .ZN(n13952) );
  NAND2_X1 U12061 ( .A1(n11379), .A2(n11380), .ZN(n9525) );
  XNOR2_X1 U12062 ( .A(n9748), .B(n11649), .ZN(n9526) );
  OAI222_X1 U12063 ( .A1(n14631), .A2(n11379), .B1(n14633), .B2(n9781), .C1(
        n14629), .C2(n9526), .ZN(n10009) );
  AOI211_X1 U12064 ( .C1(n10012), .C2(n14796), .A(n9527), .B(n10009), .ZN(
        n9530) );
  OR2_X1 U12065 ( .A1(n9530), .A2(n14806), .ZN(n9528) );
  OAI21_X1 U12066 ( .B1(n14808), .B2(n9529), .A(n9528), .ZN(P1_U3532) );
  OR2_X1 U12067 ( .A1(n9530), .A2(n14797), .ZN(n9531) );
  OAI21_X1 U12068 ( .B1(n6528), .B2(n9359), .A(n9531), .ZN(P1_U3471) );
  NOR2_X1 U12069 ( .A1(n12041), .A2(n9532), .ZN(n14918) );
  NAND2_X1 U12070 ( .A1(n12042), .A2(n12041), .ZN(n12040) );
  AND2_X1 U12071 ( .A1(n12040), .A2(n9533), .ZN(n12264) );
  NOR2_X1 U12072 ( .A1(n14960), .A2(n14892), .ZN(n9535) );
  OAI21_X1 U12073 ( .B1(n12264), .B2(n9535), .A(n9534), .ZN(n14917) );
  AOI21_X1 U12074 ( .B1(n14918), .B2(n9536), .A(n14917), .ZN(n9541) );
  AND2_X1 U12075 ( .A1(n13598), .A2(n9537), .ZN(n10096) );
  INV_X1 U12076 ( .A(n12264), .ZN(n14919) );
  OAI22_X1 U12077 ( .A1(n13598), .A2(n8904), .B1(n9538), .B2(n13595), .ZN(
        n9539) );
  AOI21_X1 U12078 ( .B1(n10096), .B2(n14919), .A(n9539), .ZN(n9540) );
  OAI21_X1 U12079 ( .B1(n9541), .B2(n13561), .A(n9540), .ZN(P2_U3265) );
  OAI21_X1 U12080 ( .B1(n9544), .B2(n9543), .A(n9542), .ZN(n9550) );
  INV_X1 U12081 ( .A(n12643), .ZN(n12665) );
  OAI22_X1 U12082 ( .A1(n9252), .A2(n12665), .B1(n15047), .B2(n12646), .ZN(
        n9545) );
  INV_X1 U12083 ( .A(n9545), .ZN(n9548) );
  NAND2_X1 U12084 ( .A1(n9546), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9547) );
  OAI211_X1 U12085 ( .C1(n12666), .C2(n9876), .A(n9548), .B(n9547), .ZN(n9549)
         );
  AOI21_X1 U12086 ( .B1(n9550), .B2(n12651), .A(n9549), .ZN(n9551) );
  INV_X1 U12087 ( .A(n9551), .ZN(P3_U3177) );
  INV_X1 U12088 ( .A(n9552), .ZN(n9553) );
  OAI21_X1 U12089 ( .B1(n15054), .B2(n9890), .A(n9553), .ZN(n9555) );
  AOI21_X1 U12090 ( .B1(n9555), .B2(n9554), .A(n11955), .ZN(n9557) );
  MUX2_X1 U12091 ( .A(n9558), .B(n9557), .S(n9556), .Z(n9559) );
  INV_X1 U12092 ( .A(n13029), .ZN(n12996) );
  MUX2_X1 U12093 ( .A(n9562), .B(n9561), .S(n15142), .Z(n9563) );
  OAI21_X1 U12094 ( .B1(n9564), .B2(n12996), .A(n9563), .ZN(P3_U3459) );
  NAND2_X1 U12095 ( .A1(n9567), .A2(n9566), .ZN(n9575) );
  INV_X1 U12096 ( .A(n9567), .ZN(n9568) );
  AND2_X1 U12097 ( .A1(n9575), .A2(n9569), .ZN(n11744) );
  INV_X1 U12098 ( .A(n9570), .ZN(n9572) );
  NAND2_X1 U12099 ( .A1(n9572), .A2(n9571), .ZN(n11741) );
  AND2_X1 U12100 ( .A1(n11744), .A2(n11741), .ZN(n9573) );
  XNOR2_X1 U12101 ( .A(n14936), .B(n6529), .ZN(n9723) );
  NAND2_X1 U12102 ( .A1(n13265), .A2(n13542), .ZN(n9724) );
  XNOR2_X1 U12103 ( .A(n9723), .B(n9724), .ZN(n9578) );
  OAI21_X1 U12104 ( .B1(n11743), .B2(n9578), .A(n13183), .ZN(n9586) );
  NOR4_X1 U12105 ( .A1(n13213), .A2(n9578), .A3(n9577), .A4(n9576), .ZN(n9585)
         );
  NAND2_X1 U12106 ( .A1(n13266), .A2(n13231), .ZN(n9581) );
  NAND2_X1 U12107 ( .A1(n13264), .A2(n13230), .ZN(n9580) );
  NAND2_X1 U12108 ( .A1(n9581), .A2(n9580), .ZN(n10177) );
  AOI22_X1 U12109 ( .A1(n13235), .A2(n10177), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9583) );
  NAND2_X1 U12110 ( .A1(n14818), .A2(n14936), .ZN(n9582) );
  OAI211_X1 U12111 ( .C1(n14821), .C2(n10181), .A(n9583), .B(n9582), .ZN(n9584) );
  AOI211_X1 U12112 ( .C1(n9586), .C2(n13227), .A(n9585), .B(n9584), .ZN(n9587)
         );
  INV_X1 U12113 ( .A(n9587), .ZN(P2_U3202) );
  INV_X1 U12114 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10606) );
  MUX2_X1 U12115 ( .A(n10606), .B(P1_REG1_REG_13__SCAN_IN), .S(n10599), .Z(
        n9590) );
  INV_X1 U12116 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10351) );
  MUX2_X1 U12117 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10351), .S(n14006), .Z(
        n13999) );
  AOI211_X1 U12118 ( .C1(n9590), .C2(n9589), .A(n10634), .B(n9694), .ZN(n9601)
         );
  AOI21_X1 U12119 ( .B1(n10346), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9591), .ZN(
        n14003) );
  INV_X1 U12120 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U12121 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9592), .S(n14006), .Z(
        n14004) );
  NAND2_X1 U12122 ( .A1(n14003), .A2(n14004), .ZN(n14002) );
  OAI21_X1 U12123 ( .B1(n14006), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14002), 
        .ZN(n9595) );
  INV_X1 U12124 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9593) );
  MUX2_X1 U12125 ( .A(n9593), .B(P1_REG2_REG_13__SCAN_IN), .S(n10599), .Z(
        n9594) );
  NOR2_X1 U12126 ( .A1(n9595), .A2(n9594), .ZN(n9692) );
  AOI211_X1 U12127 ( .C1(n9595), .C2(n9594), .A(n14021), .B(n9692), .ZN(n9600)
         );
  NAND2_X1 U12128 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13881)
         );
  INV_X1 U12129 ( .A(n13881), .ZN(n9596) );
  AOI21_X1 U12130 ( .B1(n14715), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9596), .ZN(
        n9597) );
  OAI21_X1 U12131 ( .B1(n14020), .B2(n9598), .A(n9597), .ZN(n9599) );
  OR3_X1 U12132 ( .A1(n9601), .A2(n9600), .A3(n9599), .ZN(P1_U3256) );
  MUX2_X1 U12133 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12777), .Z(n9960) );
  XNOR2_X1 U12134 ( .A(n9960), .B(n10271), .ZN(n9961) );
  INV_X1 U12135 ( .A(n9602), .ZN(n9603) );
  AOI22_X1 U12136 ( .A1(n9605), .A2(n9604), .B1(n10263), .B2(n9603), .ZN(n9962) );
  XOR2_X1 U12137 ( .A(n9961), .B(n9962), .Z(n9623) );
  NAND2_X1 U12138 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10271), .ZN(n9609) );
  OAI21_X1 U12139 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10271), .A(n9609), .ZN(
        n9954) );
  XNOR2_X1 U12140 ( .A(n9955), .B(n9954), .ZN(n9621) );
  INV_X1 U12141 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U12142 ( .A1(n9610), .A2(n15136), .B1(P3_REG1_REG_8__SCAN_IN), .B2(
        n10271), .ZN(n9616) );
  NAND2_X1 U12143 ( .A1(n9612), .A2(n9611), .ZN(n9614) );
  NAND2_X1 U12144 ( .A1(n9616), .A2(n9615), .ZN(n9971) );
  OAI21_X1 U12145 ( .B1(n9616), .B2(n9615), .A(n9971), .ZN(n9617) );
  NAND2_X1 U12146 ( .A1(n9617), .A2(n14990), .ZN(n9619) );
  NOR2_X1 U12147 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10272), .ZN(n10442) );
  AOI21_X1 U12148 ( .B1(n14987), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10442), .ZN(
        n9618) );
  OAI211_X1 U12149 ( .C1(n14981), .C2(n10271), .A(n9619), .B(n9618), .ZN(n9620) );
  AOI21_X1 U12150 ( .B1(n9621), .B2(n14554), .A(n9620), .ZN(n9622) );
  OAI21_X1 U12151 ( .B1(n9623), .B2(n14983), .A(n9622), .ZN(P3_U3190) );
  NAND2_X1 U12152 ( .A1(n9624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9625) );
  XNOR2_X1 U12153 ( .A(n9625), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14011) );
  INV_X1 U12154 ( .A(n14011), .ZN(n10834) );
  OAI222_X1 U12155 ( .A1(n14372), .A2(n15420), .B1(n14370), .B2(n11338), .C1(
        n10834), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U12156 ( .A(n13365), .ZN(n13357) );
  OAI222_X1 U12157 ( .A1(P2_U3088), .A2(n13357), .B1(n13766), .B2(n11338), 
        .C1(n9626), .C2(n13749), .ZN(P2_U3309) );
  MUX2_X1 U12158 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9627), .S(n9637), .Z(n9632) );
  MUX2_X1 U12159 ( .A(n9629), .B(P2_REG1_REG_8__SCAN_IN), .S(n9635), .Z(n14841) );
  MUX2_X1 U12160 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9630), .S(n9636), .Z(n13284) );
  OAI21_X1 U12161 ( .B1(n9636), .B2(P2_REG1_REG_9__SCAN_IN), .A(n13283), .ZN(
        n9631) );
  NOR2_X1 U12162 ( .A1(n9631), .A2(n9632), .ZN(n9846) );
  AOI211_X1 U12163 ( .C1(n9632), .C2(n9631), .A(n14858), .B(n9846), .ZN(n9645)
         );
  AOI21_X1 U12164 ( .B1(n9634), .B2(P2_REG2_REG_7__SCAN_IN), .A(n9633), .ZN(
        n14853) );
  INV_X1 U12165 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n15205) );
  MUX2_X1 U12166 ( .A(n15205), .B(P2_REG2_REG_8__SCAN_IN), .S(n9635), .Z(
        n14852) );
  NOR2_X1 U12167 ( .A1(n14853), .A2(n14852), .ZN(n14850) );
  AOI21_X1 U12168 ( .B1(n9635), .B2(P2_REG2_REG_8__SCAN_IN), .A(n14850), .ZN(
        n13292) );
  MUX2_X1 U12169 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10470), .S(n9636), .Z(
        n13291) );
  NAND2_X1 U12170 ( .A1(n13292), .A2(n13291), .ZN(n13290) );
  OAI21_X1 U12171 ( .B1(n9636), .B2(P2_REG2_REG_9__SCAN_IN), .A(n13290), .ZN(
        n9639) );
  MUX2_X1 U12172 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n13597), .S(n9637), .Z(
        n9638) );
  NOR2_X1 U12173 ( .A1(n9639), .A2(n9638), .ZN(n9840) );
  AOI211_X1 U12174 ( .C1(n9639), .C2(n9638), .A(n14851), .B(n9840), .ZN(n9644)
         );
  INV_X1 U12175 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9642) );
  NOR2_X1 U12176 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15377), .ZN(n9640) );
  AOI21_X1 U12177 ( .B1(n14865), .B2(n9847), .A(n9640), .ZN(n9641) );
  OAI21_X1 U12178 ( .B1(n14873), .B2(n9642), .A(n9641), .ZN(n9643) );
  OR3_X1 U12179 ( .A1(n9645), .A2(n9644), .A3(n9643), .ZN(P2_U3224) );
  OAI222_X1 U12180 ( .A1(n14372), .A2(n15251), .B1(n14370), .B2(n11482), .C1(
        n11635), .C2(P1_U3086), .ZN(P1_U3335) );
  NAND3_X1 U12181 ( .A1(n9647), .A2(n11689), .A3(n9646), .ZN(n14051) );
  INV_X2 U12182 ( .A(n14639), .ZN(n14747) );
  INV_X1 U12183 ( .A(n9648), .ZN(n9649) );
  AOI21_X1 U12184 ( .B1(n9650), .B2(n6896), .A(n9649), .ZN(n14750) );
  INV_X1 U12185 ( .A(n9651), .ZN(n14624) );
  OAI21_X1 U12186 ( .B1(n14752), .B2(n9919), .A(n9652), .ZN(n9656) );
  OR2_X1 U12187 ( .A1(n9656), .A2(n14674), .ZN(n14751) );
  OAI22_X1 U12188 ( .A1(n14489), .A2(n14751), .B1(n13958), .B2(n14642), .ZN(
        n9653) );
  AOI21_X1 U12189 ( .B1(n14259), .B2(n7537), .A(n9653), .ZN(n9663) );
  OAI21_X1 U12190 ( .B1(n9655), .B2(n9654), .A(n14494), .ZN(n9659) );
  XNOR2_X1 U12191 ( .A(n9656), .B(n13955), .ZN(n9657) );
  AOI21_X1 U12192 ( .B1(n9657), .B2(n14494), .A(n13957), .ZN(n9658) );
  AOI21_X1 U12193 ( .B1(n9659), .B2(n14631), .A(n9658), .ZN(n9660) );
  AOI21_X1 U12194 ( .B1(n14222), .B2(n13954), .A(n9660), .ZN(n14753) );
  MUX2_X1 U12195 ( .A(n9661), .B(n14753), .S(n14639), .Z(n9662) );
  OAI211_X1 U12196 ( .C1(n14247), .C2(n14750), .A(n9663), .B(n9662), .ZN(
        P1_U3292) );
  OR2_X1 U12197 ( .A1(n11274), .A2(SI_4_), .ZN(n9671) );
  OR2_X1 U12198 ( .A1(n11198), .A2(n9667), .ZN(n9670) );
  OR2_X1 U12199 ( .A1(n10868), .A2(n9668), .ZN(n9669) );
  AND3_X2 U12200 ( .A1(n9671), .A2(n9670), .A3(n9669), .ZN(n11846) );
  XNOR2_X1 U12201 ( .A(n11846), .B(n11789), .ZN(n9672) );
  NAND2_X1 U12202 ( .A1(n9672), .A2(n11847), .ZN(n9984) );
  OAI21_X1 U12203 ( .B1(n9672), .B2(n11847), .A(n9984), .ZN(n9673) );
  AOI21_X1 U12204 ( .B1(n9674), .B2(n9673), .A(n6688), .ZN(n9687) );
  NAND2_X1 U12205 ( .A1(n6530), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9682) );
  OR2_X1 U12206 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  NAND2_X1 U12207 ( .A1(n9993), .A2(n9677), .ZN(n10210) );
  NAND2_X1 U12208 ( .A1(n11154), .A2(n10210), .ZN(n9681) );
  NAND2_X1 U12209 ( .A1(n6531), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U12210 ( .A1(n11216), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9679) );
  INV_X1 U12211 ( .A(n11846), .ZN(n9911) );
  OAI22_X1 U12212 ( .A1(n10240), .A2(n12646), .B1(n9911), .B2(n12666), .ZN(
        n9683) );
  AOI211_X1 U12213 ( .C1(n12643), .C2(n6954), .A(n9684), .B(n9683), .ZN(n9686)
         );
  NAND2_X1 U12214 ( .A1(n12670), .A2(n9912), .ZN(n9685) );
  OAI211_X1 U12215 ( .C1(n9687), .C2(n12672), .A(n9686), .B(n9685), .ZN(
        P3_U3170) );
  XNOR2_X1 U12216 ( .A(n9831), .B(n15251), .ZN(n11186) );
  INV_X1 U12217 ( .A(n11186), .ZN(n9691) );
  OAI222_X1 U12218 ( .A1(n13120), .A2(n9691), .B1(n13122), .B2(n11187), .C1(
        P3_U3151), .C2(n9690), .ZN(P3_U3275) );
  AOI21_X1 U12219 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10599), .A(n9692), .ZN(
        n10477) );
  INV_X1 U12220 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U12221 ( .A(n9693), .B(P1_REG2_REG_14__SCAN_IN), .S(n10733), .Z(
        n10476) );
  XNOR2_X1 U12222 ( .A(n10477), .B(n10476), .ZN(n9702) );
  AOI21_X1 U12223 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10599), .A(n9694), .ZN(
        n9696) );
  INV_X1 U12224 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10621) );
  MUX2_X1 U12225 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10621), .S(n10733), .Z(
        n9695) );
  NAND2_X1 U12226 ( .A1(n9696), .A2(n9695), .ZN(n10487) );
  OAI21_X1 U12227 ( .B1(n9696), .B2(n9695), .A(n10487), .ZN(n9697) );
  NAND2_X1 U12228 ( .A1(n9697), .A2(n14727), .ZN(n9701) );
  AND2_X1 U12229 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n13781) );
  NOR2_X1 U12230 ( .A1(n14020), .A2(n9698), .ZN(n9699) );
  AOI211_X1 U12231 ( .C1(n14715), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n13781), 
        .B(n9699), .ZN(n9700) );
  OAI211_X1 U12232 ( .C1(n14021), .C2(n9702), .A(n9701), .B(n9700), .ZN(
        P1_U3257) );
  OAI22_X1 U12233 ( .A1(n11385), .A2(n6907), .B1(n11386), .B2(n12542), .ZN(
        n9703) );
  XNOR2_X1 U12234 ( .A(n9703), .B(n12551), .ZN(n9822) );
  OR2_X1 U12235 ( .A1(n11385), .A2(n12542), .ZN(n9705) );
  NAND2_X1 U12236 ( .A1(n12553), .A2(n7323), .ZN(n9704) );
  NAND2_X1 U12237 ( .A1(n9705), .A2(n9704), .ZN(n9821) );
  INV_X1 U12238 ( .A(n9706), .ZN(n9709) );
  INV_X1 U12239 ( .A(n9707), .ZN(n9708) );
  XOR2_X1 U12240 ( .A(n9823), .B(n9822), .Z(n9717) );
  INV_X1 U12241 ( .A(n12558), .ZN(n13925) );
  OAI21_X1 U12242 ( .B1(n13925), .B2(n9781), .A(n9712), .ZN(n9713) );
  AOI21_X1 U12243 ( .B1(n8890), .B2(n13953), .A(n9713), .ZN(n9714) );
  OAI21_X1 U12244 ( .B1(n10005), .B2(n14620), .A(n9714), .ZN(n9715) );
  AOI21_X1 U12245 ( .B1(n7324), .B2(n14616), .A(n9715), .ZN(n9716) );
  OAI21_X1 U12246 ( .B1(n9717), .B2(n13932), .A(n9716), .ZN(P1_U3230) );
  OAI222_X1 U12247 ( .A1(n13764), .A2(n9719), .B1(P2_U3088), .B2(n9718), .C1(
        n10417), .C2(n11482), .ZN(P2_U3307) );
  INV_X1 U12248 ( .A(n11351), .ZN(n9721) );
  OAI222_X1 U12249 ( .A1(n14372), .A2(n9720), .B1(n14370), .B2(n9721), .C1(
        P1_U3086), .C2(n14635), .ZN(P1_U3336) );
  OAI222_X1 U12250 ( .A1(n13764), .A2(n9722), .B1(n13766), .B2(n9721), .C1(
        n12044), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U12251 ( .A(n13184), .B(n12356), .ZN(n9727) );
  NAND2_X1 U12252 ( .A1(n13264), .A2(n13542), .ZN(n9726) );
  INV_X1 U12253 ( .A(n9723), .ZN(n13179) );
  NAND2_X1 U12254 ( .A1(n13179), .A2(n9724), .ZN(n9725) );
  XNOR2_X1 U12255 ( .A(n9727), .B(n9726), .ZN(n13182) );
  XNOR2_X1 U12256 ( .A(n12084), .B(n12356), .ZN(n9806) );
  INV_X1 U12257 ( .A(n9806), .ZN(n9729) );
  NAND2_X1 U12258 ( .A1(n13263), .A2(n13542), .ZN(n9730) );
  INV_X1 U12259 ( .A(n9730), .ZN(n9728) );
  AND2_X1 U12260 ( .A1(n9729), .A2(n9728), .ZN(n9856) );
  INV_X1 U12261 ( .A(n9856), .ZN(n9731) );
  NAND2_X1 U12262 ( .A1(n9806), .A2(n9730), .ZN(n9854) );
  NAND2_X1 U12263 ( .A1(n9731), .A2(n9854), .ZN(n9732) );
  INV_X1 U12264 ( .A(n9732), .ZN(n9734) );
  INV_X1 U12265 ( .A(n9855), .ZN(n9733) );
  NOR2_X1 U12266 ( .A1(n9733), .A2(n9732), .ZN(n9808) );
  INV_X1 U12267 ( .A(n9808), .ZN(n9805) );
  OAI211_X1 U12268 ( .C1(n9855), .C2(n9734), .A(n9805), .B(n13227), .ZN(n9739)
         );
  INV_X1 U12269 ( .A(n10194), .ZN(n9737) );
  AOI22_X1 U12270 ( .A1(n13230), .A2(n13262), .B1(n13264), .B2(n13231), .ZN(
        n10072) );
  OAI21_X1 U12271 ( .B1(n14811), .B2(n10072), .A(n9735), .ZN(n9736) );
  AOI21_X1 U12272 ( .B1(n9737), .B2(n13223), .A(n9736), .ZN(n9738) );
  OAI211_X1 U12273 ( .C1(n7365), .C2(n13238), .A(n9739), .B(n9738), .ZN(
        P2_U3211) );
  NAND2_X1 U12274 ( .A1(n9741), .A2(n11622), .ZN(n9744) );
  AOI22_X1 U12275 ( .A1(n11613), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11455), 
        .B2(n9742), .ZN(n9743) );
  NAND2_X1 U12276 ( .A1(n14758), .A2(n9781), .ZN(n9771) );
  OR2_X1 U12277 ( .A1(n14758), .A2(n9781), .ZN(n9745) );
  NAND2_X1 U12278 ( .A1(n9771), .A2(n9745), .ZN(n11650) );
  INV_X1 U12279 ( .A(n11650), .ZN(n9750) );
  XNOR2_X1 U12280 ( .A(n9765), .B(n9750), .ZN(n14762) );
  NAND2_X1 U12281 ( .A1(n9746), .A2(n11352), .ZN(n11334) );
  NOR2_X1 U12282 ( .A1(n11385), .A2(n7323), .ZN(n9747) );
  NAND2_X1 U12283 ( .A1(n9749), .A2(n9750), .ZN(n9772) );
  OAI21_X1 U12284 ( .B1(n9750), .B2(n9749), .A(n9772), .ZN(n9759) );
  NAND2_X1 U12285 ( .A1(n6963), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9756) );
  INV_X1 U12286 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9751) );
  OR2_X1 U12287 ( .A1(n11607), .A2(n9751), .ZN(n9755) );
  NAND2_X1 U12288 ( .A1(n9752), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9775) );
  OAI21_X1 U12289 ( .B1(n9752), .B2(P1_REG3_REG_6__SCAN_IN), .A(n9775), .ZN(
        n10155) );
  OR2_X1 U12290 ( .A1(n11608), .A2(n10155), .ZN(n9754) );
  OR2_X1 U12291 ( .A1(n11630), .A2(n9786), .ZN(n9753) );
  NAND4_X1 U12292 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(n13951) );
  INV_X1 U12293 ( .A(n13951), .ZN(n10151) );
  OAI22_X1 U12294 ( .A1(n10151), .A2(n14633), .B1(n11386), .B2(n14631), .ZN(
        n9758) );
  NOR2_X1 U12295 ( .A1(n14762), .A2(n14496), .ZN(n9757) );
  AOI211_X1 U12296 ( .C1(n14494), .C2(n9759), .A(n9758), .B(n9757), .ZN(n14761) );
  MUX2_X1 U12297 ( .A(n9760), .B(n14761), .S(n14639), .Z(n9764) );
  INV_X1 U12298 ( .A(n9827), .ZN(n9761) );
  OAI22_X1 U12299 ( .A1(n14738), .A2(n6809), .B1(n9761), .B2(n14642), .ZN(
        n9762) );
  AOI21_X1 U12300 ( .B1(n14757), .B2(n14743), .A(n9762), .ZN(n9763) );
  OAI211_X1 U12301 ( .C1(n14762), .C2(n14739), .A(n9764), .B(n9763), .ZN(
        P1_U3288) );
  OR2_X1 U12302 ( .A1(n14758), .A2(n13952), .ZN(n9766) );
  NAND2_X1 U12303 ( .A1(n9767), .A2(n11622), .ZN(n9770) );
  AOI22_X1 U12304 ( .A1(n11613), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11455), 
        .B2(n9768), .ZN(n9769) );
  NAND2_X1 U12305 ( .A1(n9770), .A2(n9769), .ZN(n11398) );
  XNOR2_X1 U12306 ( .A(n11398), .B(n13951), .ZN(n11651) );
  XNOR2_X1 U12307 ( .A(n9925), .B(n11651), .ZN(n14765) );
  NAND2_X1 U12308 ( .A1(n9772), .A2(n9771), .ZN(n9933) );
  XNOR2_X1 U12309 ( .A(n9933), .B(n11651), .ZN(n9783) );
  NAND2_X1 U12310 ( .A1(n6963), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9780) );
  INV_X1 U12311 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9773) );
  OR2_X1 U12312 ( .A1(n11607), .A2(n9773), .ZN(n9779) );
  AND2_X1 U12313 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  OR2_X1 U12314 ( .A1(n9776), .A2(n9937), .ZN(n10328) );
  OR2_X1 U12315 ( .A1(n11608), .A2(n10328), .ZN(n9778) );
  OR2_X1 U12316 ( .A1(n11630), .A2(n9947), .ZN(n9777) );
  NAND4_X1 U12317 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n13950) );
  INV_X1 U12318 ( .A(n13950), .ZN(n10323) );
  OAI22_X1 U12319 ( .A1(n9781), .A2(n14631), .B1(n10323), .B2(n14633), .ZN(
        n9782) );
  AOI21_X1 U12320 ( .B1(n9783), .B2(n14494), .A(n9782), .ZN(n9784) );
  OAI21_X1 U12321 ( .B1(n14765), .B2(n14496), .A(n9784), .ZN(n14768) );
  INV_X1 U12322 ( .A(n14768), .ZN(n9785) );
  MUX2_X1 U12323 ( .A(n9786), .B(n9785), .S(n14639), .Z(n9791) );
  INV_X1 U12324 ( .A(n11398), .ZN(n14767) );
  NAND2_X1 U12325 ( .A1(n14767), .A2(n9787), .ZN(n9948) );
  OAI211_X1 U12326 ( .C1(n14767), .C2(n9787), .A(n8808), .B(n9948), .ZN(n14766) );
  INV_X1 U12327 ( .A(n14766), .ZN(n9789) );
  OAI22_X1 U12328 ( .A1(n14738), .A2(n14767), .B1(n10155), .B2(n14642), .ZN(
        n9788) );
  AOI21_X1 U12329 ( .B1(n14743), .B2(n9789), .A(n9788), .ZN(n9790) );
  OAI211_X1 U12330 ( .C1(n14765), .C2(n14739), .A(n9791), .B(n9790), .ZN(
        P1_U3287) );
  NOR2_X1 U12331 ( .A1(n14642), .A2(n9792), .ZN(n9793) );
  AOI21_X1 U12332 ( .B1(n14747), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9793), .ZN(
        n9796) );
  NAND2_X1 U12333 ( .A1(n14743), .A2(n9794), .ZN(n9795) );
  OAI211_X1 U12334 ( .C1(n14738), .C2(n11374), .A(n9796), .B(n9795), .ZN(n9797) );
  AOI21_X1 U12335 ( .B1(n14262), .B2(n9798), .A(n9797), .ZN(n9799) );
  OAI21_X1 U12336 ( .B1(n14747), .B2(n9800), .A(n9799), .ZN(P1_U3291) );
  INV_X1 U12337 ( .A(n12091), .ZN(n14880) );
  XNOR2_X1 U12338 ( .A(n12091), .B(n12356), .ZN(n9864) );
  NAND2_X1 U12339 ( .A1(n13262), .A2(n13542), .ZN(n9801) );
  NAND2_X1 U12340 ( .A1(n9864), .A2(n9801), .ZN(n9857) );
  INV_X1 U12341 ( .A(n9864), .ZN(n9803) );
  INV_X1 U12342 ( .A(n9801), .ZN(n9802) );
  NAND2_X1 U12343 ( .A1(n9803), .A2(n9802), .ZN(n9858) );
  AND2_X1 U12344 ( .A1(n9857), .A2(n9858), .ZN(n9807) );
  INV_X1 U12345 ( .A(n9807), .ZN(n9804) );
  AOI21_X1 U12346 ( .B1(n9805), .B2(n9804), .A(n14813), .ZN(n9810) );
  NOR3_X1 U12347 ( .A1(n13213), .A2(n12086), .A3(n9806), .ZN(n9809) );
  OAI21_X1 U12348 ( .B1(n9808), .B2(n9856), .A(n9807), .ZN(n9862) );
  OAI21_X1 U12349 ( .B1(n9810), .B2(n9809), .A(n9862), .ZN(n9817) );
  INV_X1 U12350 ( .A(n9811), .ZN(n14876) );
  NAND2_X1 U12351 ( .A1(n13263), .A2(n13231), .ZN(n9813) );
  NAND2_X1 U12352 ( .A1(n13261), .A2(n13230), .ZN(n9812) );
  NAND2_X1 U12353 ( .A1(n9813), .A2(n9812), .ZN(n10304) );
  INV_X1 U12354 ( .A(n10304), .ZN(n9814) );
  OAI22_X1 U12355 ( .A1(n14811), .A2(n9814), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7922), .ZN(n9815) );
  AOI21_X1 U12356 ( .B1(n14876), .B2(n13223), .A(n9815), .ZN(n9816) );
  OAI211_X1 U12357 ( .C1(n14880), .C2(n13238), .A(n9817), .B(n9816), .ZN(
        P2_U3185) );
  NAND2_X1 U12358 ( .A1(n14758), .A2(n6923), .ZN(n9819) );
  NAND2_X1 U12359 ( .A1(n12554), .A2(n13952), .ZN(n9818) );
  NAND2_X1 U12360 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  XNOR2_X1 U12361 ( .A(n9820), .B(n12551), .ZN(n10143) );
  AOI22_X1 U12362 ( .A1(n14758), .A2(n12554), .B1(n12553), .B2(n13952), .ZN(
        n10144) );
  XNOR2_X1 U12363 ( .A(n10143), .B(n10144), .ZN(n10146) );
  XOR2_X1 U12364 ( .A(n10146), .B(n10147), .Z(n9830) );
  INV_X1 U12365 ( .A(n14620), .ZN(n13918) );
  NAND2_X1 U12366 ( .A1(n8890), .A2(n7323), .ZN(n9824) );
  OAI211_X1 U12367 ( .C1(n13925), .C2(n10151), .A(n9825), .B(n9824), .ZN(n9826) );
  AOI21_X1 U12368 ( .B1(n9827), .B2(n13918), .A(n9826), .ZN(n9829) );
  NAND2_X1 U12369 ( .A1(n14616), .A2(n14758), .ZN(n9828) );
  OAI211_X1 U12370 ( .C1(n9830), .C2(n13932), .A(n9829), .B(n9828), .ZN(
        P1_U3227) );
  INV_X1 U12371 ( .A(SI_21_), .ZN(n11200) );
  INV_X1 U12372 ( .A(n9831), .ZN(n9832) );
  NAND2_X1 U12373 ( .A1(n9832), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9835) );
  INV_X1 U12374 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U12375 ( .A1(n15252), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12376 ( .A1(n9916), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U12377 ( .A1(n10186), .A2(n9836), .ZN(n9837) );
  NAND2_X1 U12378 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  NAND2_X1 U12379 ( .A1(n10187), .A2(n9839), .ZN(n11199) );
  OAI222_X1 U12380 ( .A1(P3_U3151), .A2(n11828), .B1(n13122), .B2(n11200), 
        .C1(n13120), .C2(n11199), .ZN(P3_U3274) );
  AOI21_X1 U12381 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n9847), .A(n9840), .ZN(
        n9842) );
  INV_X1 U12382 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11074) );
  MUX2_X1 U12383 ( .A(n11074), .B(P2_REG2_REG_11__SCAN_IN), .S(n11075), .Z(
        n9841) );
  NAND2_X1 U12384 ( .A1(n9842), .A2(n9841), .ZN(n13306) );
  OAI21_X1 U12385 ( .B1(n9842), .B2(n9841), .A(n13306), .ZN(n9852) );
  INV_X1 U12386 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9845) );
  AND2_X1 U12387 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9843) );
  AOI21_X1 U12388 ( .B1(n14865), .B2(n11066), .A(n9843), .ZN(n9844) );
  OAI21_X1 U12389 ( .B1(n14873), .B2(n9845), .A(n9844), .ZN(n9851) );
  XNOR2_X1 U12390 ( .A(n11066), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n9848) );
  AOI211_X1 U12391 ( .C1(n9849), .C2(n9848), .A(n14858), .B(n11065), .ZN(n9850) );
  AOI211_X1 U12392 ( .C1(n14867), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9853)
         );
  INV_X1 U12393 ( .A(n9853), .ZN(P2_U3225) );
  XNOR2_X1 U12394 ( .A(n14952), .B(n6529), .ZN(n11806) );
  NAND2_X1 U12395 ( .A1(n13261), .A2(n13542), .ZN(n10373) );
  XNOR2_X1 U12396 ( .A(n11806), .B(n10373), .ZN(n9865) );
  NAND2_X1 U12397 ( .A1(n9857), .A2(n9856), .ZN(n9859) );
  OAI21_X1 U12398 ( .B1(n9862), .B2(n9865), .A(n10376), .ZN(n9873) );
  OR4_X1 U12399 ( .A1(n9865), .A2(n9864), .A3(n13213), .A4(n9863), .ZN(n9871)
         );
  NAND2_X1 U12400 ( .A1(n13262), .A2(n13231), .ZN(n9867) );
  NAND2_X1 U12401 ( .A1(n13260), .A2(n13230), .ZN(n9866) );
  AND2_X1 U12402 ( .A1(n9867), .A2(n9866), .ZN(n10406) );
  OR2_X1 U12403 ( .A1(n14821), .A2(n10411), .ZN(n9868) );
  NAND2_X1 U12404 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14843) );
  OAI211_X1 U12405 ( .C1(n14811), .C2(n10406), .A(n9868), .B(n14843), .ZN(
        n9869) );
  INV_X1 U12406 ( .A(n9869), .ZN(n9870) );
  OAI211_X1 U12407 ( .C1(n10412), .C2(n13238), .A(n9871), .B(n9870), .ZN(n9872) );
  AOI21_X1 U12408 ( .B1(n9873), .B2(n13227), .A(n9872), .ZN(n9874) );
  INV_X1 U12409 ( .A(n9874), .ZN(P2_U3193) );
  INV_X1 U12410 ( .A(n9876), .ZN(n9877) );
  NAND2_X1 U12411 ( .A1(n9887), .A2(n9877), .ZN(n11838) );
  NAND2_X1 U12412 ( .A1(n15043), .A2(n11838), .ZN(n9901) );
  INV_X1 U12413 ( .A(n9903), .ZN(n9878) );
  XNOR2_X1 U12414 ( .A(n9901), .B(n11984), .ZN(n15095) );
  INV_X1 U12415 ( .A(n15095), .ZN(n9900) );
  AND2_X1 U12416 ( .A1(n9891), .A2(n15056), .ZN(n15025) );
  INV_X1 U12417 ( .A(n15025), .ZN(n15078) );
  NOR2_X1 U12418 ( .A1(n15083), .A2(n15078), .ZN(n12846) );
  INV_X1 U12419 ( .A(n12846), .ZN(n10461) );
  AND2_X1 U12420 ( .A1(n15054), .A2(n12030), .ZN(n9879) );
  NAND2_X1 U12421 ( .A1(n9880), .A2(n9879), .ZN(n9882) );
  NAND2_X1 U12422 ( .A1(n9882), .A2(n9881), .ZN(n15050) );
  INV_X1 U12423 ( .A(n9883), .ZN(n9884) );
  OAI22_X1 U12424 ( .A1(n9887), .A2(n15048), .B1(n11847), .B2(n15046), .ZN(
        n9896) );
  NAND2_X1 U12425 ( .A1(n9252), .A2(n9885), .ZN(n9886) );
  NAND2_X1 U12426 ( .A1(n9887), .A2(n9876), .ZN(n9888) );
  NAND2_X1 U12427 ( .A1(n9891), .A2(n9890), .ZN(n12024) );
  INV_X1 U12428 ( .A(n9905), .ZN(n9893) );
  AOI211_X1 U12429 ( .C1(n11984), .C2(n9894), .A(n15053), .B(n9893), .ZN(n9895) );
  AOI211_X1 U12430 ( .C1(n15095), .C2(n15050), .A(n9896), .B(n9895), .ZN(
        n15092) );
  MUX2_X1 U12431 ( .A(n15260), .B(n15092), .S(n15080), .Z(n9899) );
  AND2_X1 U12432 ( .A1(n9903), .A2(n15073), .ZN(n15094) );
  AOI22_X1 U12433 ( .A1(n15028), .A2(n15094), .B1(n15075), .B2(n9897), .ZN(
        n9898) );
  OAI211_X1 U12434 ( .C1(n9900), .C2(n10461), .A(n9899), .B(n9898), .ZN(
        P3_U3230) );
  NAND2_X1 U12435 ( .A1(n11847), .A2(n11846), .ZN(n11850) );
  NAND2_X1 U12436 ( .A1(n12683), .A2(n9911), .ZN(n9902) );
  XNOR2_X1 U12437 ( .A(n10129), .B(n10128), .ZN(n15096) );
  INV_X1 U12438 ( .A(n15050), .ZN(n15072) );
  INV_X1 U12439 ( .A(n10240), .ZN(n12682) );
  AOI22_X1 U12440 ( .A1(n15065), .A2(n12682), .B1(n6954), .B2(n15062), .ZN(
        n9908) );
  NAND2_X1 U12441 ( .A1(n6954), .A2(n9903), .ZN(n9904) );
  OAI211_X1 U12442 ( .C1(n9906), .C2(n10128), .A(n10109), .B(n15068), .ZN(
        n9907) );
  OAI211_X1 U12443 ( .C1(n15096), .C2(n15072), .A(n9908), .B(n9907), .ZN(
        n15097) );
  INV_X1 U12444 ( .A(n15097), .ZN(n9909) );
  MUX2_X1 U12445 ( .A(n9910), .B(n9909), .S(n15080), .Z(n9914) );
  NOR2_X1 U12446 ( .A1(n9911), .A2(n15054), .ZN(n15098) );
  AOI22_X1 U12447 ( .A1(n15098), .A2(n15028), .B1(n15075), .B2(n9912), .ZN(
        n9913) );
  OAI211_X1 U12448 ( .C1(n15096), .C2(n10461), .A(n9914), .B(n9913), .ZN(
        P3_U3229) );
  OAI222_X1 U12449 ( .A1(n14372), .A2(n15252), .B1(n14370), .B2(n11497), .C1(
        n11308), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U12450 ( .A1(n13764), .A2(n9916), .B1(P2_U3088), .B2(n9915), .C1(
        n10417), .C2(n11497), .ZN(P2_U3306) );
  INV_X1 U12451 ( .A(n11366), .ZN(n11647) );
  AOI21_X1 U12452 ( .B1(n14494), .B2(n14639), .A(n14262), .ZN(n9923) );
  OAI22_X1 U12453 ( .A1(n14747), .A2(n9918), .B1(n9917), .B2(n14642), .ZN(
        n9921) );
  NOR2_X1 U12454 ( .A1(n14489), .A2(n14674), .ZN(n14195) );
  INV_X1 U12455 ( .A(n14195), .ZN(n10365) );
  AOI21_X1 U12456 ( .B1(n10365), .B2(n14738), .A(n9919), .ZN(n9920) );
  AOI211_X1 U12457 ( .C1(n14747), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9921), .B(
        n9920), .ZN(n9922) );
  OAI21_X1 U12458 ( .B1(n11647), .B2(n9923), .A(n9922), .ZN(P1_U3293) );
  INV_X1 U12459 ( .A(n11651), .ZN(n9924) );
  NAND2_X1 U12460 ( .A1(n9925), .A2(n9924), .ZN(n9927) );
  OR2_X1 U12461 ( .A1(n11398), .A2(n13951), .ZN(n9926) );
  NAND2_X1 U12462 ( .A1(n9928), .A2(n11622), .ZN(n9931) );
  AOI22_X1 U12463 ( .A1(n11613), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11455), 
        .B2(n9929), .ZN(n9930) );
  NAND2_X1 U12464 ( .A1(n9931), .A2(n9930), .ZN(n11403) );
  XNOR2_X1 U12465 ( .A(n11403), .B(n13950), .ZN(n11652) );
  XNOR2_X1 U12466 ( .A(n10015), .B(n11652), .ZN(n14771) );
  OR2_X1 U12467 ( .A1(n11398), .A2(n10151), .ZN(n9932) );
  NAND2_X1 U12468 ( .A1(n9933), .A2(n9932), .ZN(n9935) );
  NAND2_X1 U12469 ( .A1(n11398), .A2(n10151), .ZN(n9934) );
  NAND2_X1 U12470 ( .A1(n9935), .A2(n9934), .ZN(n10037) );
  XNOR2_X1 U12471 ( .A(n10037), .B(n11652), .ZN(n9944) );
  NAND2_X1 U12472 ( .A1(n11582), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9942) );
  OR2_X1 U12473 ( .A1(n11583), .A2(n9936), .ZN(n9941) );
  NAND2_X1 U12474 ( .A1(n9937), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10030) );
  OR2_X1 U12475 ( .A1(n9937), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12476 ( .A1(n10030), .A2(n9938), .ZN(n10507) );
  OR2_X1 U12477 ( .A1(n11608), .A2(n10507), .ZN(n9940) );
  OR2_X1 U12478 ( .A1(n11630), .A2(n10063), .ZN(n9939) );
  NAND4_X1 U12479 ( .A1(n9942), .A2(n9941), .A3(n9940), .A4(n9939), .ZN(n13949) );
  INV_X1 U12480 ( .A(n13949), .ZN(n10330) );
  OAI22_X1 U12481 ( .A1(n10151), .A2(n14631), .B1(n10330), .B2(n14633), .ZN(
        n9943) );
  AOI21_X1 U12482 ( .B1(n9944), .B2(n14494), .A(n9943), .ZN(n9945) );
  OAI21_X1 U12483 ( .B1(n14771), .B2(n14496), .A(n9945), .ZN(n14774) );
  INV_X1 U12484 ( .A(n14774), .ZN(n9946) );
  MUX2_X1 U12485 ( .A(n9947), .B(n9946), .S(n14639), .Z(n9953) );
  AOI21_X1 U12486 ( .B1(n9948), .B2(n11403), .A(n14674), .ZN(n9949) );
  NAND2_X1 U12487 ( .A1(n9949), .A2(n10057), .ZN(n14772) );
  INV_X1 U12488 ( .A(n14772), .ZN(n9951) );
  INV_X1 U12489 ( .A(n11403), .ZN(n14773) );
  OAI22_X1 U12490 ( .A1(n14738), .A2(n14773), .B1(n10328), .B2(n14642), .ZN(
        n9950) );
  AOI21_X1 U12491 ( .B1(n14743), .B2(n9951), .A(n9950), .ZN(n9952) );
  OAI211_X1 U12492 ( .C1(n14771), .C2(n14739), .A(n9953), .B(n9952), .ZN(
        P1_U3286) );
  INV_X1 U12493 ( .A(n14982), .ZN(n10254) );
  NOR2_X1 U12494 ( .A1(n10254), .A2(n9956), .ZN(n9957) );
  INV_X1 U12495 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15030) );
  INV_X1 U12496 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U12497 ( .A1(n10540), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15013), 
        .B2(n10522), .ZN(n9958) );
  NOR2_X1 U12498 ( .A1(n9959), .A2(n9958), .ZN(n10521) );
  AOI21_X1 U12499 ( .B1(n9959), .B2(n9958), .A(n10521), .ZN(n9983) );
  OAI22_X1 U12500 ( .A1(n9962), .A2(n9961), .B1(n9960), .B2(n10271), .ZN(
        n14976) );
  MUX2_X1 U12501 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12777), .Z(n9963) );
  NAND2_X1 U12502 ( .A1(n9963), .A2(n14982), .ZN(n14977) );
  NAND2_X1 U12503 ( .A1(n14976), .A2(n14977), .ZN(n14975) );
  INV_X1 U12504 ( .A(n9963), .ZN(n9964) );
  NAND2_X1 U12505 ( .A1(n9964), .A2(n10254), .ZN(n14979) );
  INV_X1 U12506 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U12507 ( .A(n15013), .B(n9965), .S(n12777), .Z(n9966) );
  NAND2_X1 U12508 ( .A1(n9966), .A2(n10540), .ZN(n10527) );
  INV_X1 U12509 ( .A(n9966), .ZN(n9967) );
  NAND2_X1 U12510 ( .A1(n9967), .A2(n10522), .ZN(n9968) );
  NAND2_X1 U12511 ( .A1(n10527), .A2(n9968), .ZN(n9969) );
  AOI21_X1 U12512 ( .B1(n14975), .B2(n14979), .A(n9969), .ZN(n10529) );
  AND3_X1 U12513 ( .A1(n14975), .A2(n14979), .A3(n9969), .ZN(n9970) );
  OAI21_X1 U12514 ( .B1(n10529), .B2(n9970), .A(n12795), .ZN(n9982) );
  AOI22_X1 U12515 ( .A1(n10540), .A2(n9965), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n10522), .ZN(n9976) );
  NAND2_X1 U12516 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10271), .ZN(n9972) );
  NAND2_X1 U12517 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  NAND2_X1 U12518 ( .A1(n14982), .A2(n9973), .ZN(n9974) );
  XNOR2_X1 U12519 ( .A(n9973), .B(n10254), .ZN(n14989) );
  OAI21_X1 U12520 ( .B1(n9976), .B2(n9975), .A(n10524), .ZN(n9980) );
  INV_X1 U12521 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U12522 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9977), .ZN(n10538) );
  AOI21_X1 U12523 ( .B1(n14987), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n10538), 
        .ZN(n9978) );
  OAI21_X1 U12524 ( .B1(n14981), .B2(n10522), .A(n9978), .ZN(n9979) );
  AOI21_X1 U12525 ( .B1(n9980), .B2(n14990), .A(n9979), .ZN(n9981) );
  OAI211_X1 U12526 ( .C1(n9983), .C2(n14994), .A(n9982), .B(n9981), .ZN(
        P3_U3192) );
  INV_X1 U12527 ( .A(n9984), .ZN(n9985) );
  OR2_X1 U12528 ( .A1(n11274), .A2(SI_5_), .ZN(n9990) );
  OR2_X1 U12529 ( .A1(n11198), .A2(n9986), .ZN(n9989) );
  OR2_X1 U12530 ( .A1(n10868), .A2(n9987), .ZN(n9988) );
  XNOR2_X1 U12531 ( .A(n10110), .B(n11789), .ZN(n10241) );
  XNOR2_X1 U12532 ( .A(n10241), .B(n10240), .ZN(n9991) );
  AOI21_X1 U12533 ( .B1(n9992), .B2(n9991), .A(n10292), .ZN(n10004) );
  NAND2_X1 U12534 ( .A1(n6530), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U12535 ( .A1(n9993), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9994) );
  AND2_X1 U12536 ( .A1(n10120), .A2(n9994), .ZN(n15041) );
  INV_X1 U12537 ( .A(n15041), .ZN(n9995) );
  NAND2_X1 U12538 ( .A1(n11154), .A2(n9995), .ZN(n9998) );
  NAND2_X1 U12539 ( .A1(n6532), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U12540 ( .A1(n11216), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9996) );
  INV_X1 U12541 ( .A(n10110), .ZN(n10209) );
  OAI22_X1 U12542 ( .A1(n10281), .A2(n12646), .B1(n10209), .B2(n12666), .ZN(
        n10000) );
  AOI211_X1 U12543 ( .C1(n12643), .C2(n12683), .A(n10001), .B(n10000), .ZN(
        n10003) );
  NAND2_X1 U12544 ( .A1(n12670), .A2(n10210), .ZN(n10002) );
  OAI211_X1 U12545 ( .C1(n10004), .C2(n12672), .A(n10003), .B(n10002), .ZN(
        P3_U3167) );
  INV_X1 U12546 ( .A(n10005), .ZN(n10006) );
  INV_X1 U12547 ( .A(n14642), .ZN(n14735) );
  AOI22_X1 U12548 ( .A1(n14259), .A2(n7324), .B1(n10006), .B2(n14735), .ZN(
        n10007) );
  OAI21_X1 U12549 ( .B1(n10365), .B2(n10008), .A(n10007), .ZN(n10011) );
  MUX2_X1 U12550 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10009), .S(n14639), .Z(
        n10010) );
  AOI211_X1 U12551 ( .C1(n14262), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10013) );
  INV_X1 U12552 ( .A(n10013), .ZN(P1_U3289) );
  INV_X1 U12553 ( .A(n11652), .ZN(n10014) );
  NAND2_X1 U12554 ( .A1(n10015), .A2(n10014), .ZN(n10017) );
  OR2_X1 U12555 ( .A1(n11403), .A2(n13950), .ZN(n10016) );
  NAND2_X1 U12556 ( .A1(n10017), .A2(n10016), .ZN(n10056) );
  NAND2_X1 U12557 ( .A1(n10018), .A2(n11622), .ZN(n10021) );
  AOI22_X1 U12558 ( .A1(n11613), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11455), 
        .B2(n10019), .ZN(n10020) );
  XNOR2_X1 U12559 ( .A(n11409), .B(n13949), .ZN(n11654) );
  NAND2_X1 U12560 ( .A1(n10056), .A2(n10059), .ZN(n10023) );
  OR2_X1 U12561 ( .A1(n11409), .A2(n13949), .ZN(n10022) );
  NAND2_X1 U12562 ( .A1(n10024), .A2(n11622), .ZN(n10027) );
  AOI22_X1 U12563 ( .A1(n11613), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11455), 
        .B2(n10025), .ZN(n10026) );
  NAND2_X1 U12564 ( .A1(n11582), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10035) );
  OR2_X1 U12565 ( .A1(n11583), .A2(n10028), .ZN(n10034) );
  INV_X1 U12566 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U12567 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NAND2_X1 U12568 ( .A1(n10042), .A2(n10031), .ZN(n10790) );
  OR2_X1 U12569 ( .A1(n11608), .A2(n10790), .ZN(n10033) );
  OR2_X1 U12570 ( .A1(n11630), .A2(n8772), .ZN(n10032) );
  NAND4_X1 U12571 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n13948) );
  XNOR2_X1 U12572 ( .A(n11413), .B(n13948), .ZN(n11657) );
  XNOR2_X1 U12573 ( .A(n10236), .B(n11657), .ZN(n14782) );
  AND2_X1 U12574 ( .A1(n11403), .A2(n10323), .ZN(n10036) );
  OAI22_X1 U12575 ( .A1(n10037), .A2(n10036), .B1(n10323), .B2(n11403), .ZN(
        n10060) );
  NAND2_X1 U12576 ( .A1(n10060), .A2(n11654), .ZN(n10039) );
  OR2_X1 U12577 ( .A1(n11409), .A2(n10330), .ZN(n10038) );
  NAND2_X1 U12578 ( .A1(n10039), .A2(n10038), .ZN(n10214) );
  INV_X1 U12579 ( .A(n11657), .ZN(n10235) );
  XNOR2_X1 U12580 ( .A(n10214), .B(n10235), .ZN(n10049) );
  NAND2_X1 U12581 ( .A1(n6963), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10047) );
  INV_X1 U12582 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10040) );
  OR2_X1 U12583 ( .A1(n11607), .A2(n10040), .ZN(n10046) );
  NAND2_X1 U12584 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  NAND2_X1 U12585 ( .A1(n10225), .A2(n10043), .ZN(n10852) );
  OR2_X1 U12586 ( .A1(n11608), .A2(n10852), .ZN(n10045) );
  OR2_X1 U12587 ( .A1(n11630), .A2(n10222), .ZN(n10044) );
  NAND4_X1 U12588 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n13947) );
  OAI22_X1 U12589 ( .A1(n10846), .A2(n14633), .B1(n10330), .B2(n14631), .ZN(
        n10048) );
  AOI21_X1 U12590 ( .B1(n10049), .B2(n14494), .A(n10048), .ZN(n10050) );
  OAI21_X1 U12591 ( .B1(n14782), .B2(n14496), .A(n10050), .ZN(n14785) );
  NAND2_X1 U12592 ( .A1(n14785), .A2(n14639), .ZN(n10055) );
  OAI22_X1 U12593 ( .A1(n14639), .A2(n8772), .B1(n10790), .B2(n14642), .ZN(
        n10053) );
  INV_X1 U12594 ( .A(n11413), .ZN(n14784) );
  OAI211_X1 U12595 ( .C1(n14784), .C2(n10051), .A(n8808), .B(n10223), .ZN(
        n14783) );
  NOR2_X1 U12596 ( .A1(n14783), .A2(n14489), .ZN(n10052) );
  AOI211_X1 U12597 ( .C1(n14259), .C2(n11413), .A(n10053), .B(n10052), .ZN(
        n10054) );
  OAI211_X1 U12598 ( .C1(n14782), .C2(n14739), .A(n10055), .B(n10054), .ZN(
        P1_U3284) );
  XNOR2_X1 U12599 ( .A(n10056), .B(n10059), .ZN(n14780) );
  INV_X1 U12600 ( .A(n14780), .ZN(n10067) );
  OAI211_X1 U12601 ( .C1(n7495), .C2(n7496), .A(n8808), .B(n10058), .ZN(n14777) );
  XNOR2_X1 U12602 ( .A(n10060), .B(n10059), .ZN(n10061) );
  AOI222_X1 U12603 ( .A1(n14494), .A2(n10061), .B1(n13948), .B2(n14222), .C1(
        n13950), .C2(n14221), .ZN(n14778) );
  OAI21_X1 U12604 ( .B1(n11352), .B2(n14777), .A(n14778), .ZN(n10062) );
  NAND2_X1 U12605 ( .A1(n10062), .A2(n14639), .ZN(n10066) );
  OAI22_X1 U12606 ( .A1(n14639), .A2(n10063), .B1(n10507), .B2(n14642), .ZN(
        n10064) );
  AOI21_X1 U12607 ( .B1(n14259), .B2(n11409), .A(n10064), .ZN(n10065) );
  OAI211_X1 U12608 ( .C1(n14247), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        P1_U3285) );
  INV_X1 U12609 ( .A(n14943), .ZN(n14955) );
  XNOR2_X1 U12610 ( .A(n10069), .B(n12269), .ZN(n10190) );
  AOI21_X1 U12611 ( .B1(n10099), .B2(n12084), .A(n14896), .ZN(n10070) );
  AND2_X1 U12612 ( .A1(n10070), .A2(n10302), .ZN(n10196) );
  XOR2_X1 U12613 ( .A(n10071), .B(n12269), .Z(n10073) );
  OAI21_X1 U12614 ( .B1(n10073), .B2(n13509), .A(n10072), .ZN(n10191) );
  AOI211_X1 U12615 ( .C1(n14927), .C2(n10190), .A(n10196), .B(n10191), .ZN(
        n10081) );
  AOI22_X1 U12616 ( .A1(n13692), .A2(n12084), .B1(n14970), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10074) );
  OAI21_X1 U12617 ( .B1(n10081), .B2(n14970), .A(n10074), .ZN(P2_U3505) );
  INV_X1 U12618 ( .A(n10075), .ZN(n10076) );
  AND2_X1 U12619 ( .A1(n14912), .A2(n10076), .ZN(n10077) );
  NAND2_X1 U12620 ( .A1(n14962), .A2(n14953), .ZN(n13730) );
  INV_X1 U12621 ( .A(n13730), .ZN(n13744) );
  NOR2_X1 U12622 ( .A1(n14962), .A2(n7906), .ZN(n10079) );
  AOI21_X1 U12623 ( .B1(n13744), .B2(n12084), .A(n10079), .ZN(n10080) );
  OAI21_X1 U12624 ( .B1(n10081), .B2(n14961), .A(n10080), .ZN(P2_U3448) );
  INV_X1 U12625 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n15242) );
  INV_X1 U12626 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n11167) );
  INV_X1 U12627 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15147) );
  INV_X1 U12628 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U12629 ( .A1(n11191), .A2(n11190), .ZN(n11203) );
  INV_X1 U12630 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n11225) );
  INV_X1 U12631 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n11236) );
  INV_X1 U12632 ( .A(n10313), .ZN(n10083) );
  NAND2_X1 U12633 ( .A1(n11263), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U12634 ( .A1(n10083), .A2(n10082), .ZN(n12830) );
  NAND2_X1 U12635 ( .A1(n11154), .A2(n12830), .ZN(n10088) );
  NAND2_X1 U12636 ( .A1(n6530), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12637 ( .A1(n6531), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U12638 ( .A1(n6944), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U12639 ( .A1(n12837), .A2(P3_U3897), .ZN(n10089) );
  OAI21_X1 U12640 ( .B1(P3_U3897), .B2(n15242), .A(n10089), .ZN(P3_U3518) );
  INV_X1 U12641 ( .A(n13595), .ZN(n14902) );
  AOI22_X1 U12642 ( .A1(n13600), .A2(n12053), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14902), .ZN(n10090) );
  OAI21_X1 U12643 ( .B1(n13578), .B2(n10091), .A(n10090), .ZN(n10094) );
  MUX2_X1 U12644 ( .A(n10092), .B(P2_REG2_REG_1__SCAN_IN), .S(n13561), .Z(
        n10093) );
  AOI211_X1 U12645 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10097) );
  INV_X1 U12646 ( .A(n10097), .ZN(P2_U3264) );
  XNOR2_X1 U12647 ( .A(n13264), .B(n13184), .ZN(n12268) );
  XOR2_X1 U12648 ( .A(n10098), .B(n12268), .Z(n14950) );
  OAI211_X1 U12649 ( .C1(n10180), .C2(n14947), .A(n13557), .B(n10099), .ZN(
        n14944) );
  AOI22_X1 U12650 ( .A1(n13600), .A2(n13184), .B1(n14902), .B2(n13173), .ZN(
        n10100) );
  OAI21_X1 U12651 ( .B1(n14944), .B2(n13578), .A(n10100), .ZN(n10106) );
  XOR2_X1 U12652 ( .A(n10101), .B(n12268), .Z(n10104) );
  NAND2_X1 U12653 ( .A1(n13265), .A2(n13231), .ZN(n10103) );
  NAND2_X1 U12654 ( .A1(n13263), .A2(n13230), .ZN(n10102) );
  AND2_X1 U12655 ( .A1(n10103), .A2(n10102), .ZN(n13177) );
  OAI21_X1 U12656 ( .B1(n10104), .B2(n13509), .A(n13177), .ZN(n14949) );
  MUX2_X1 U12657 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14949), .S(n13598), .Z(
        n10105) );
  AOI211_X1 U12658 ( .C1(n14950), .C2(n14883), .A(n10106), .B(n10105), .ZN(
        n10107) );
  INV_X1 U12659 ( .A(n10107), .ZN(P2_U3260) );
  NAND2_X1 U12660 ( .A1(n12683), .A2(n11846), .ZN(n10108) );
  NAND2_X1 U12661 ( .A1(n10240), .A2(n10110), .ZN(n11851) );
  NAND2_X1 U12662 ( .A1(n12682), .A2(n10209), .ZN(n11857) );
  OR2_X1 U12663 ( .A1(n11274), .A2(n10111), .ZN(n10114) );
  OR2_X1 U12664 ( .A1(n11198), .A2(n10112), .ZN(n10113) );
  OAI211_X1 U12665 ( .C1(n6534), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n15037) );
  NAND2_X1 U12666 ( .A1(n10281), .A2(n15037), .ZN(n11861) );
  INV_X1 U12667 ( .A(n15037), .ZN(n10245) );
  NAND2_X1 U12668 ( .A1(n12681), .A2(n10245), .ZN(n11859) );
  NAND2_X1 U12669 ( .A1(n11861), .A2(n11859), .ZN(n10130) );
  NAND2_X1 U12670 ( .A1(n10240), .A2(n10209), .ZN(n10117) );
  AND2_X1 U12671 ( .A1(n10130), .A2(n10117), .ZN(n10116) );
  INV_X1 U12672 ( .A(n10426), .ZN(n10119) );
  AOI21_X1 U12673 ( .B1(n10203), .B2(n10117), .A(n10130), .ZN(n10118) );
  NOR3_X1 U12674 ( .A1(n10119), .A2(n10118), .A3(n15053), .ZN(n10127) );
  NAND2_X1 U12675 ( .A1(n6530), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10125) );
  AND2_X1 U12676 ( .A1(n10120), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10121) );
  OR2_X1 U12677 ( .A1(n10121), .A2(n10273), .ZN(n10458) );
  NAND2_X1 U12678 ( .A1(n11154), .A2(n10458), .ZN(n10124) );
  NAND2_X1 U12679 ( .A1(n6533), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12680 ( .A1(n6944), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10122) );
  OAI22_X1 U12681 ( .A1(n10445), .A2(n15046), .B1(n10240), .B2(n15048), .ZN(
        n10126) );
  NOR2_X1 U12682 ( .A1(n10127), .A2(n10126), .ZN(n15032) );
  INV_X1 U12683 ( .A(n15142), .ZN(n15140) );
  INV_X1 U12684 ( .A(n10128), .ZN(n11990) );
  NAND2_X1 U12685 ( .A1(n10200), .A2(n11989), .ZN(n10422) );
  NAND2_X1 U12686 ( .A1(n10422), .A2(n11851), .ZN(n10131) );
  INV_X1 U12687 ( .A(n10130), .ZN(n11985) );
  NAND2_X1 U12688 ( .A1(n10131), .A2(n11985), .ZN(n10133) );
  OR2_X1 U12689 ( .A1(n10131), .A2(n11985), .ZN(n10132) );
  AND2_X1 U12690 ( .A1(n10133), .A2(n10132), .ZN(n15033) );
  INV_X1 U12691 ( .A(n15033), .ZN(n10141) );
  INV_X1 U12692 ( .A(n13040), .ZN(n10136) );
  OAI22_X1 U12693 ( .A1(n12996), .A2(n10245), .B1(n15142), .B2(n9299), .ZN(
        n10135) );
  AOI21_X1 U12694 ( .B1(n10141), .B2(n10136), .A(n10135), .ZN(n10137) );
  OAI21_X1 U12695 ( .B1(n15032), .B2(n15140), .A(n10137), .ZN(P3_U3465) );
  INV_X1 U12696 ( .A(n14601), .ZN(n10138) );
  INV_X1 U12697 ( .A(n13107), .ZN(n10140) );
  INV_X1 U12698 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15145) );
  OAI22_X1 U12699 ( .A1(n10245), .A2(n13049), .B1(n15127), .B2(n15145), .ZN(
        n10139) );
  AOI21_X1 U12700 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10142) );
  OAI21_X1 U12701 ( .B1(n15032), .B2(n15125), .A(n10142), .ZN(P3_U3408) );
  INV_X1 U12702 ( .A(n10143), .ZN(n10145) );
  NAND2_X1 U12703 ( .A1(n11398), .A2(n6923), .ZN(n10149) );
  NAND2_X1 U12704 ( .A1(n12554), .A2(n13951), .ZN(n10148) );
  NAND2_X1 U12705 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  XNOR2_X1 U12706 ( .A(n10150), .B(n12551), .ZN(n10320) );
  NOR2_X1 U12707 ( .A1(n12525), .A2(n10151), .ZN(n10152) );
  AOI21_X1 U12708 ( .B1(n11398), .B2(n12554), .A(n10152), .ZN(n10322) );
  XNOR2_X1 U12709 ( .A(n10320), .B(n10322), .ZN(n10153) );
  OAI211_X1 U12710 ( .C1(n10154), .C2(n10153), .A(n10321), .B(n14612), .ZN(
        n10160) );
  NOR2_X1 U12711 ( .A1(n14620), .A2(n10155), .ZN(n10158) );
  OAI21_X1 U12712 ( .B1(n13925), .B2(n10323), .A(n10156), .ZN(n10157) );
  AOI211_X1 U12713 ( .C1(n8890), .C2(n13952), .A(n10158), .B(n10157), .ZN(
        n10159) );
  OAI211_X1 U12714 ( .C1(n14767), .C2(n13921), .A(n10160), .B(n10159), .ZN(
        P1_U3239) );
  XNOR2_X1 U12715 ( .A(n10161), .B(n12265), .ZN(n14924) );
  OAI21_X1 U12716 ( .B1(n12265), .B2(n10163), .A(n10162), .ZN(n10165) );
  AOI21_X1 U12717 ( .B1(n10165), .B2(n14892), .A(n10164), .ZN(n14922) );
  MUX2_X1 U12718 ( .A(n14922), .B(n10166), .S(n13561), .Z(n10172) );
  INV_X1 U12719 ( .A(n14897), .ZN(n10167) );
  AOI211_X1 U12720 ( .C1(n7852), .C2(n10168), .A(n14896), .B(n10167), .ZN(
        n14921) );
  OAI22_X1 U12721 ( .A1(n14879), .A2(n10169), .B1(n13595), .B2(n14827), .ZN(
        n10170) );
  AOI21_X1 U12722 ( .B1(n14874), .B2(n14921), .A(n10170), .ZN(n10171) );
  OAI211_X1 U12723 ( .C1(n13582), .C2(n14924), .A(n10172), .B(n10171), .ZN(
        P2_U3263) );
  XNOR2_X1 U12724 ( .A(n10173), .B(n10175), .ZN(n14939) );
  OAI21_X1 U12725 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10178) );
  AOI21_X1 U12726 ( .B1(n10178), .B2(n14892), .A(n10177), .ZN(n14938) );
  MUX2_X1 U12727 ( .A(n10179), .B(n14938), .S(n13598), .Z(n10185) );
  AOI211_X1 U12728 ( .C1(n14936), .C2(n14898), .A(n14896), .B(n10180), .ZN(
        n14935) );
  OAI22_X1 U12729 ( .A1(n14879), .A2(n10182), .B1(n10181), .B2(n13595), .ZN(
        n10183) );
  AOI21_X1 U12730 ( .B1(n14935), .B2(n14874), .A(n10183), .ZN(n10184) );
  OAI211_X1 U12731 ( .C1(n13582), .C2(n14939), .A(n10185), .B(n10184), .ZN(
        P2_U3261) );
  XNOR2_X1 U12732 ( .A(n10419), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n10368) );
  XNOR2_X1 U12733 ( .A(n10369), .B(n10368), .ZN(n11210) );
  INV_X1 U12734 ( .A(n11210), .ZN(n10189) );
  OAI22_X1 U12735 ( .A1(n12034), .A2(P3_U3151), .B1(SI_22_), .B2(n13115), .ZN(
        n10188) );
  AOI21_X1 U12736 ( .B1(n10189), .B2(n13109), .A(n10188), .ZN(P3_U3273) );
  INV_X1 U12737 ( .A(n10190), .ZN(n10199) );
  INV_X1 U12738 ( .A(n10191), .ZN(n10192) );
  MUX2_X1 U12739 ( .A(n10193), .B(n10192), .S(n13598), .Z(n10198) );
  OAI22_X1 U12740 ( .A1(n14879), .A2(n7365), .B1(n10194), .B2(n13595), .ZN(
        n10195) );
  AOI21_X1 U12741 ( .B1(n14874), .B2(n10196), .A(n10195), .ZN(n10197) );
  OAI211_X1 U12742 ( .C1(n10199), .C2(n13582), .A(n10198), .B(n10197), .ZN(
        P2_U3259) );
  XNOR2_X1 U12743 ( .A(n10200), .B(n7206), .ZN(n15101) );
  NAND2_X1 U12744 ( .A1(n10201), .A2(n11989), .ZN(n10202) );
  NAND2_X1 U12745 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  NAND2_X1 U12746 ( .A1(n10204), .A2(n15068), .ZN(n10207) );
  OAI22_X1 U12747 ( .A1(n10281), .A2(n15046), .B1(n11847), .B2(n15048), .ZN(
        n10205) );
  INV_X1 U12748 ( .A(n10205), .ZN(n10206) );
  OAI211_X1 U12749 ( .C1(n15101), .C2(n15072), .A(n10207), .B(n10206), .ZN(
        n15102) );
  MUX2_X1 U12750 ( .A(n15102), .B(P3_REG2_REG_5__SCAN_IN), .S(n15083), .Z(
        n10208) );
  INV_X1 U12751 ( .A(n10208), .ZN(n10212) );
  NOR2_X1 U12752 ( .A1(n10209), .A2(n15054), .ZN(n15103) );
  AOI22_X1 U12753 ( .A1(n15103), .A2(n15028), .B1(n15075), .B2(n10210), .ZN(
        n10211) );
  OAI211_X1 U12754 ( .C1(n15101), .C2(n10461), .A(n10212), .B(n10211), .ZN(
        P3_U3228) );
  INV_X1 U12755 ( .A(n13948), .ZN(n10785) );
  NAND2_X1 U12756 ( .A1(n11413), .A2(n10785), .ZN(n10213) );
  NAND2_X1 U12757 ( .A1(n10215), .A2(n11622), .ZN(n10218) );
  AOI22_X1 U12758 ( .A1(n11613), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11455), 
        .B2(n10216), .ZN(n10217) );
  OR2_X1 U12759 ( .A1(n14790), .A2(n10846), .ZN(n10343) );
  NAND2_X1 U12760 ( .A1(n14790), .A2(n10846), .ZN(n10219) );
  NAND2_X1 U12761 ( .A1(n10343), .A2(n10219), .ZN(n11656) );
  AOI21_X1 U12762 ( .B1(n10220), .B2(n11656), .A(n14629), .ZN(n10221) );
  AOI22_X1 U12763 ( .A1(n10221), .A2(n10344), .B1(n14221), .B2(n13948), .ZN(
        n14792) );
  OAI22_X1 U12764 ( .A1(n14639), .A2(n10222), .B1(n10852), .B2(n14642), .ZN(
        n10234) );
  AOI21_X1 U12765 ( .B1(n10223), .B2(n14790), .A(n14674), .ZN(n10232) );
  NAND2_X1 U12766 ( .A1(n11582), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10231) );
  INV_X1 U12767 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10224) );
  AND2_X1 U12768 ( .A1(n10225), .A2(n10224), .ZN(n10226) );
  OR2_X1 U12769 ( .A1(n10226), .A2(n10349), .ZN(n14619) );
  OR2_X1 U12770 ( .A1(n11608), .A2(n14619), .ZN(n10230) );
  OR2_X1 U12771 ( .A1(n11630), .A2(n10362), .ZN(n10229) );
  OR2_X1 U12772 ( .A1(n11583), .A2(n10227), .ZN(n10228) );
  NAND4_X1 U12773 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n13946) );
  AOI22_X1 U12774 ( .A1(n10232), .A2(n10360), .B1(n14222), .B2(n13946), .ZN(
        n14791) );
  NOR2_X1 U12775 ( .A1(n14791), .A2(n14489), .ZN(n10233) );
  AOI211_X1 U12776 ( .C1(n14259), .C2(n14790), .A(n10234), .B(n10233), .ZN(
        n10239) );
  OR2_X1 U12777 ( .A1(n11413), .A2(n13948), .ZN(n10237) );
  XNOR2_X1 U12778 ( .A(n10359), .B(n11656), .ZN(n14795) );
  NAND2_X1 U12779 ( .A1(n14795), .A2(n14262), .ZN(n10238) );
  OAI211_X1 U12780 ( .C1(n14792), .C2(n14747), .A(n10239), .B(n10238), .ZN(
        P1_U3283) );
  INV_X1 U12781 ( .A(n12670), .ZN(n10250) );
  NAND2_X1 U12782 ( .A1(n10241), .A2(n10240), .ZN(n10283) );
  INV_X1 U12783 ( .A(n10283), .ZN(n10242) );
  NOR2_X1 U12784 ( .A1(n10292), .A2(n10242), .ZN(n10244) );
  XNOR2_X1 U12785 ( .A(n15037), .B(n9489), .ZN(n10284) );
  XNOR2_X1 U12786 ( .A(n10281), .B(n10284), .ZN(n10243) );
  NAND2_X1 U12787 ( .A1(n10244), .A2(n10243), .ZN(n10336) );
  OAI211_X1 U12788 ( .C1(n10244), .C2(n10243), .A(n10336), .B(n12651), .ZN(
        n10249) );
  OAI22_X1 U12789 ( .A1(n10445), .A2(n12646), .B1(n10245), .B2(n12666), .ZN(
        n10246) );
  AOI211_X1 U12790 ( .C1(n12643), .C2(n12682), .A(n10247), .B(n10246), .ZN(
        n10248) );
  OAI211_X1 U12791 ( .C1(n15041), .C2(n10250), .A(n10249), .B(n10248), .ZN(
        P3_U3179) );
  OR2_X1 U12792 ( .A1(n11274), .A2(SI_9_), .ZN(n10253) );
  OR2_X1 U12793 ( .A1(n11198), .A2(n10251), .ZN(n10252) );
  OAI211_X1 U12794 ( .C1(n10254), .C2(n6534), .A(n10253), .B(n10252), .ZN(
        n15026) );
  XNOR2_X1 U12795 ( .A(n15026), .B(n11786), .ZN(n10553) );
  NAND2_X1 U12796 ( .A1(n6530), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n10261) );
  OR2_X1 U12797 ( .A1(n10275), .A2(n10255), .ZN(n10256) );
  NAND2_X1 U12798 ( .A1(n10257), .A2(n10256), .ZN(n15027) );
  NAND2_X1 U12799 ( .A1(n11154), .A2(n15027), .ZN(n10260) );
  NAND2_X1 U12800 ( .A1(n6533), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12801 ( .A1(n6944), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n10258) );
  XNOR2_X1 U12802 ( .A(n10553), .B(n15001), .ZN(n10294) );
  OR2_X1 U12803 ( .A1(n11274), .A2(SI_7_), .ZN(n10266) );
  OR2_X1 U12804 ( .A1(n11198), .A2(n10262), .ZN(n10265) );
  OR2_X1 U12805 ( .A1(n6534), .A2(n10263), .ZN(n10264) );
  NAND2_X1 U12806 ( .A1(n10445), .A2(n10457), .ZN(n11862) );
  INV_X1 U12807 ( .A(n10457), .ZN(n10337) );
  NAND2_X1 U12808 ( .A1(n12680), .A2(n10337), .ZN(n11863) );
  NAND2_X1 U12809 ( .A1(n11862), .A2(n11863), .ZN(n10452) );
  XNOR2_X1 U12810 ( .A(n10452), .B(n9489), .ZN(n10438) );
  OR2_X1 U12811 ( .A1(n11274), .A2(n10267), .ZN(n10270) );
  OR2_X1 U12812 ( .A1(n11198), .A2(n10268), .ZN(n10269) );
  OAI211_X1 U12813 ( .C1(n10868), .C2(n10271), .A(n10270), .B(n10269), .ZN(
        n10915) );
  XNOR2_X1 U12814 ( .A(n10915), .B(n11770), .ZN(n10287) );
  NAND2_X1 U12815 ( .A1(n6530), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10279) );
  NOR2_X1 U12816 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  OR2_X1 U12817 ( .A1(n10275), .A2(n10274), .ZN(n10447) );
  NAND2_X1 U12818 ( .A1(n11154), .A2(n10447), .ZN(n10278) );
  NAND2_X1 U12819 ( .A1(n6533), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U12820 ( .A1(n6944), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10276) );
  NAND4_X1 U12821 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n12679) );
  INV_X1 U12822 ( .A(n10286), .ZN(n10440) );
  INV_X1 U12823 ( .A(n10284), .ZN(n10280) );
  NAND2_X1 U12824 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND4_X1 U12825 ( .A1(n10438), .A2(n10440), .A3(n10283), .A4(n10282), .ZN(
        n10291) );
  NAND2_X1 U12826 ( .A1(n12681), .A2(n10284), .ZN(n10335) );
  OAI21_X1 U12827 ( .B1(n10286), .B2(n10335), .A(n10438), .ZN(n10289) );
  INV_X1 U12828 ( .A(n10438), .ZN(n10285) );
  OAI21_X1 U12829 ( .B1(n10286), .B2(n10445), .A(n10285), .ZN(n10288) );
  AOI22_X1 U12830 ( .A1(n10289), .A2(n10288), .B1(n10287), .B2(n12679), .ZN(
        n10290) );
  AOI21_X1 U12831 ( .B1(n10294), .B2(n10293), .A(n10555), .ZN(n10298) );
  AND2_X1 U12832 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n14986) );
  INV_X1 U12833 ( .A(n12679), .ZN(n15020) );
  OAI22_X1 U12834 ( .A1(n15020), .A2(n12665), .B1(n15026), .B2(n12666), .ZN(
        n10295) );
  AOI211_X1 U12835 ( .C1(n12663), .C2(n10919), .A(n14986), .B(n10295), .ZN(
        n10297) );
  NAND2_X1 U12836 ( .A1(n12670), .A2(n15027), .ZN(n10296) );
  OAI211_X1 U12837 ( .C1(n10298), .C2(n12672), .A(n10297), .B(n10296), .ZN(
        P3_U3171) );
  OAI21_X1 U12838 ( .B1(n10301), .B2(n10300), .A(n6942), .ZN(n14882) );
  AOI211_X1 U12839 ( .C1(n12091), .C2(n10302), .A(n14896), .B(n10409), .ZN(
        n14875) );
  XNOR2_X1 U12840 ( .A(n10303), .B(n12270), .ZN(n10305) );
  AOI21_X1 U12841 ( .B1(n10305), .B2(n14892), .A(n10304), .ZN(n14885) );
  INV_X1 U12842 ( .A(n14885), .ZN(n10306) );
  AOI211_X1 U12843 ( .C1(n14927), .C2(n14882), .A(n14875), .B(n10306), .ZN(
        n10311) );
  INV_X1 U12844 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10307) );
  NOR2_X1 U12845 ( .A1(n14962), .A2(n10307), .ZN(n10308) );
  AOI21_X1 U12846 ( .B1(n13744), .B2(n12091), .A(n10308), .ZN(n10309) );
  OAI21_X1 U12847 ( .B1(n10311), .B2(n14961), .A(n10309), .ZN(P2_U3451) );
  AOI22_X1 U12848 ( .A1(n13692), .A2(n12091), .B1(n14970), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10310) );
  OAI21_X1 U12849 ( .B1(n10311), .B2(n14970), .A(n10310), .ZN(P2_U3506) );
  INV_X1 U12850 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15375) );
  INV_X1 U12851 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n10312) );
  NOR2_X1 U12852 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  NAND2_X1 U12853 ( .A1(n11154), .A2(n12814), .ZN(n10318) );
  NAND2_X1 U12854 ( .A1(n6530), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U12855 ( .A1(n6532), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U12856 ( .A1(n6944), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U12857 ( .A1(n12828), .A2(P3_U3897), .ZN(n10319) );
  OAI21_X1 U12858 ( .B1(P3_U3897), .B2(n15375), .A(n10319), .ZN(P3_U3519) );
  NOR2_X1 U12859 ( .A1(n12525), .A2(n10323), .ZN(n10324) );
  AOI21_X1 U12860 ( .B1(n11403), .B2(n12554), .A(n10324), .ZN(n10501) );
  AOI22_X1 U12861 ( .A1(n11403), .A2(n6923), .B1(n12554), .B2(n13950), .ZN(
        n10325) );
  XNOR2_X1 U12862 ( .A(n10325), .B(n12551), .ZN(n10500) );
  XOR2_X1 U12863 ( .A(n10501), .B(n10500), .Z(n10326) );
  OAI211_X1 U12864 ( .C1(n10327), .C2(n10326), .A(n10499), .B(n14612), .ZN(
        n10334) );
  NOR2_X1 U12865 ( .A1(n14620), .A2(n10328), .ZN(n10332) );
  OAI21_X1 U12866 ( .B1(n13925), .B2(n10330), .A(n10329), .ZN(n10331) );
  AOI211_X1 U12867 ( .C1(n8890), .C2(n13951), .A(n10332), .B(n10331), .ZN(
        n10333) );
  OAI211_X1 U12868 ( .C1(n14773), .C2(n13921), .A(n10334), .B(n10333), .ZN(
        P1_U3213) );
  NAND2_X1 U12869 ( .A1(n10336), .A2(n10335), .ZN(n10439) );
  XNOR2_X1 U12870 ( .A(n10439), .B(n10438), .ZN(n10342) );
  OAI22_X1 U12871 ( .A1(n15020), .A2(n12646), .B1(n12666), .B2(n10337), .ZN(
        n10338) );
  AOI211_X1 U12872 ( .C1(n12643), .C2(n12681), .A(n10339), .B(n10338), .ZN(
        n10341) );
  NAND2_X1 U12873 ( .A1(n12670), .A2(n10458), .ZN(n10340) );
  OAI211_X1 U12874 ( .C1(n10342), .C2(n12672), .A(n10341), .B(n10340), .ZN(
        P3_U3153) );
  NAND2_X1 U12875 ( .A1(n10345), .A2(n11622), .ZN(n10348) );
  AOI22_X1 U12876 ( .A1(n11613), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10346), 
        .B2(n11455), .ZN(n10347) );
  XNOR2_X1 U12877 ( .A(n14672), .B(n13946), .ZN(n11658) );
  XNOR2_X1 U12878 ( .A(n10611), .B(n10590), .ZN(n10358) );
  NAND2_X1 U12879 ( .A1(n11582), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10355) );
  OR2_X1 U12880 ( .A1(n11630), .A2(n9592), .ZN(n10354) );
  NAND2_X1 U12881 ( .A1(n10349), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10603) );
  OR2_X1 U12882 ( .A1(n10349), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U12883 ( .A1(n10603), .A2(n10350), .ZN(n14497) );
  OR2_X1 U12884 ( .A1(n11608), .A2(n14497), .ZN(n10353) );
  OR2_X1 U12885 ( .A1(n11583), .A2(n10351), .ZN(n10352) );
  OR2_X1 U12886 ( .A1(n12410), .A2(n14633), .ZN(n10357) );
  NAND2_X1 U12887 ( .A1(n13947), .A2(n14221), .ZN(n10356) );
  NAND2_X1 U12888 ( .A1(n10357), .A2(n10356), .ZN(n14615) );
  AOI21_X1 U12889 ( .B1(n10358), .B2(n14494), .A(n14615), .ZN(n14680) );
  XNOR2_X1 U12890 ( .A(n10591), .B(n10590), .ZN(n14677) );
  AND2_X1 U12891 ( .A1(n10360), .A2(n14672), .ZN(n10361) );
  OR2_X1 U12892 ( .A1(n10361), .A2(n14488), .ZN(n14675) );
  OAI22_X1 U12893 ( .A1(n14639), .A2(n10362), .B1(n14619), .B2(n14642), .ZN(
        n10363) );
  AOI21_X1 U12894 ( .B1(n14672), .B2(n14259), .A(n10363), .ZN(n10364) );
  OAI21_X1 U12895 ( .B1(n14675), .B2(n10365), .A(n10364), .ZN(n10366) );
  AOI21_X1 U12896 ( .B1(n14677), .B2(n14262), .A(n10366), .ZN(n10367) );
  OAI21_X1 U12897 ( .B1(n14680), .B2(n14747), .A(n10367), .ZN(P1_U3282) );
  NAND2_X1 U12898 ( .A1(n10419), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10370) );
  XNOR2_X1 U12899 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n10582) );
  XNOR2_X1 U12900 ( .A(n10583), .B(n10582), .ZN(n11221) );
  NAND2_X1 U12901 ( .A1(n11221), .A2(n13109), .ZN(n10371) );
  OAI211_X1 U12902 ( .C1(n11222), .C2(n13115), .A(n10371), .B(n12036), .ZN(
        P3_U3272) );
  INV_X1 U12903 ( .A(n13601), .ZN(n10388) );
  AND2_X1 U12904 ( .A1(n13259), .A2(n13542), .ZN(n10372) );
  NAND2_X1 U12905 ( .A1(n10396), .A2(n10372), .ZN(n10390) );
  OAI21_X1 U12906 ( .B1(n10396), .B2(n10372), .A(n10390), .ZN(n10382) );
  NAND2_X1 U12907 ( .A1(n13260), .A2(n13542), .ZN(n10377) );
  INV_X1 U12908 ( .A(n10377), .ZN(n10380) );
  XNOR2_X1 U12909 ( .A(n12103), .B(n6529), .ZN(n10379) );
  INV_X1 U12910 ( .A(n10373), .ZN(n10374) );
  NAND2_X1 U12911 ( .A1(n10376), .A2(n10375), .ZN(n10378) );
  XNOR2_X1 U12912 ( .A(n10379), .B(n10377), .ZN(n11807) );
  AOI211_X1 U12913 ( .C1(n10382), .C2(n10381), .A(n14813), .B(n10392), .ZN(
        n10383) );
  INV_X1 U12914 ( .A(n10383), .ZN(n10387) );
  INV_X1 U12915 ( .A(n13596), .ZN(n10385) );
  AOI22_X1 U12916 ( .A1(n13231), .A2(n13260), .B1(n13258), .B2(n13230), .ZN(
        n10678) );
  OAI22_X1 U12917 ( .A1(n14811), .A2(n10678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15377), .ZN(n10384) );
  AOI21_X1 U12918 ( .B1(n10385), .B2(n13223), .A(n10384), .ZN(n10386) );
  OAI211_X1 U12919 ( .C1(n10388), .C2(n13238), .A(n10387), .B(n10386), .ZN(
        P2_U3189) );
  NOR2_X1 U12920 ( .A1(n10389), .A2(n12345), .ZN(n10561) );
  INV_X1 U12921 ( .A(n10390), .ZN(n10391) );
  AOI21_X1 U12922 ( .B1(n10392), .B2(n10397), .A(n11137), .ZN(n10400) );
  NOR2_X1 U12923 ( .A1(n14821), .A2(n10777), .ZN(n10395) );
  AOI22_X1 U12924 ( .A1(n13231), .A2(n13259), .B1(n13257), .B2(n13230), .ZN(
        n10773) );
  OAI22_X1 U12925 ( .A1(n14811), .A2(n10773), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10393), .ZN(n10394) );
  AOI211_X1 U12926 ( .C1(n12115), .C2(n14818), .A(n10395), .B(n10394), .ZN(
        n10399) );
  NAND4_X1 U12927 ( .A1(n10397), .A2(n13205), .A3(n13259), .A4(n10396), .ZN(
        n10398) );
  OAI211_X1 U12928 ( .C1(n10400), .C2(n14813), .A(n10399), .B(n10398), .ZN(
        P2_U3208) );
  INV_X1 U12929 ( .A(n10401), .ZN(n10402) );
  AOI21_X1 U12930 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n14959) );
  INV_X1 U12931 ( .A(n14959), .ZN(n14956) );
  XNOR2_X1 U12932 ( .A(n10405), .B(n10404), .ZN(n10407) );
  OAI21_X1 U12933 ( .B1(n10407), .B2(n13509), .A(n10406), .ZN(n14958) );
  INV_X1 U12934 ( .A(n14958), .ZN(n10408) );
  MUX2_X1 U12935 ( .A(n15205), .B(n10408), .S(n13598), .Z(n10415) );
  INV_X1 U12936 ( .A(n10409), .ZN(n10410) );
  AOI211_X1 U12937 ( .C1(n14952), .C2(n10410), .A(n14896), .B(n10469), .ZN(
        n14951) );
  OAI22_X1 U12938 ( .A1(n14879), .A2(n10412), .B1(n10411), .B2(n13595), .ZN(
        n10413) );
  AOI21_X1 U12939 ( .B1(n14951), .B2(n14874), .A(n10413), .ZN(n10414) );
  OAI211_X1 U12940 ( .C1(n13582), .C2(n14956), .A(n10415), .B(n10414), .ZN(
        P2_U3257) );
  OAI222_X1 U12941 ( .A1(n13764), .A2(n10419), .B1(P2_U3088), .B2(n10418), 
        .C1(n10417), .C2(n10416), .ZN(P2_U3305) );
  AND2_X1 U12942 ( .A1(n11851), .A2(n11861), .ZN(n10421) );
  INV_X1 U12943 ( .A(n10452), .ZN(n11991) );
  NAND2_X1 U12944 ( .A1(n10450), .A2(n11991), .ZN(n10423) );
  NAND2_X1 U12945 ( .A1(n15020), .A2(n10915), .ZN(n11867) );
  INV_X1 U12946 ( .A(n10915), .ZN(n10424) );
  NAND2_X1 U12947 ( .A1(n12679), .A2(n10424), .ZN(n11868) );
  XNOR2_X1 U12948 ( .A(n10904), .B(n11988), .ZN(n10429) );
  INV_X1 U12949 ( .A(n10429), .ZN(n15112) );
  NAND2_X1 U12950 ( .A1(n12681), .A2(n15037), .ZN(n10425) );
  NAND2_X1 U12951 ( .A1(n12680), .A2(n10457), .ZN(n10427) );
  XNOR2_X1 U12952 ( .A(n10916), .B(n11988), .ZN(n10428) );
  NAND2_X1 U12953 ( .A1(n10428), .A2(n15068), .ZN(n10432) );
  NAND2_X1 U12954 ( .A1(n10429), .A2(n15050), .ZN(n10431) );
  AOI22_X1 U12955 ( .A1(n12680), .A2(n15062), .B1(n15065), .B2(n15001), .ZN(
        n10430) );
  NAND3_X1 U12956 ( .A1(n10432), .A2(n10431), .A3(n10430), .ZN(n15114) );
  NAND2_X1 U12957 ( .A1(n15114), .A2(n15080), .ZN(n10437) );
  INV_X1 U12958 ( .A(n15028), .ZN(n10434) );
  NAND2_X1 U12959 ( .A1(n10915), .A2(n15073), .ZN(n15111) );
  INV_X1 U12960 ( .A(n10447), .ZN(n10433) );
  OAI22_X1 U12961 ( .A1(n10434), .A2(n15111), .B1(n10433), .B2(n15040), .ZN(
        n10435) );
  AOI21_X1 U12962 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15083), .A(n10435), .ZN(
        n10436) );
  OAI211_X1 U12963 ( .C1(n15112), .C2(n10461), .A(n10437), .B(n10436), .ZN(
        P3_U3225) );
  MUX2_X1 U12964 ( .A(n12680), .B(n10439), .S(n10438), .Z(n10441) );
  XNOR2_X1 U12965 ( .A(n10441), .B(n10440), .ZN(n10449) );
  AOI22_X1 U12966 ( .A1(n12648), .A2(n10915), .B1(n15001), .B2(n12663), .ZN(
        n10444) );
  INV_X1 U12967 ( .A(n10442), .ZN(n10443) );
  OAI211_X1 U12968 ( .C1(n10445), .C2(n12665), .A(n10444), .B(n10443), .ZN(
        n10446) );
  AOI21_X1 U12969 ( .B1(n10447), .B2(n12670), .A(n10446), .ZN(n10448) );
  OAI21_X1 U12970 ( .B1(n10449), .B2(n12672), .A(n10448), .ZN(P3_U3161) );
  XNOR2_X1 U12971 ( .A(n10450), .B(n10452), .ZN(n15106) );
  AOI22_X1 U12972 ( .A1(n12681), .A2(n15062), .B1(n15065), .B2(n12679), .ZN(
        n10455) );
  OAI211_X1 U12973 ( .C1(n10453), .C2(n10452), .A(n10451), .B(n15068), .ZN(
        n10454) );
  OAI211_X1 U12974 ( .C1(n15106), .C2(n15072), .A(n10455), .B(n10454), .ZN(
        n15107) );
  INV_X1 U12975 ( .A(n15107), .ZN(n10456) );
  MUX2_X1 U12976 ( .A(n9608), .B(n10456), .S(n15080), .Z(n10460) );
  AND2_X1 U12977 ( .A1(n10457), .A2(n15073), .ZN(n15108) );
  AOI22_X1 U12978 ( .A1(n15028), .A2(n15108), .B1(n15075), .B2(n10458), .ZN(
        n10459) );
  OAI211_X1 U12979 ( .C1(n15106), .C2(n10461), .A(n10460), .B(n10459), .ZN(
        P3_U3226) );
  XNOR2_X1 U12980 ( .A(n10462), .B(n10463), .ZN(n10513) );
  AOI21_X1 U12981 ( .B1(n10464), .B2(n10463), .A(n13509), .ZN(n10468) );
  NAND2_X1 U12982 ( .A1(n13261), .A2(n13231), .ZN(n10466) );
  NAND2_X1 U12983 ( .A1(n13259), .A2(n13230), .ZN(n10465) );
  NAND2_X1 U12984 ( .A1(n10466), .A2(n10465), .ZN(n11803) );
  AOI21_X1 U12985 ( .B1(n10468), .B2(n10467), .A(n11803), .ZN(n10512) );
  INV_X1 U12986 ( .A(n10512), .ZN(n10474) );
  OAI211_X1 U12987 ( .C1(n10469), .C2(n10517), .A(n13557), .B(n10674), .ZN(
        n10511) );
  OAI22_X1 U12988 ( .A1(n13598), .A2(n10470), .B1(n11805), .B2(n13595), .ZN(
        n10471) );
  AOI21_X1 U12989 ( .B1(n12103), .B2(n13600), .A(n10471), .ZN(n10472) );
  OAI21_X1 U12990 ( .B1(n10511), .B2(n13578), .A(n10472), .ZN(n10473) );
  AOI21_X1 U12991 ( .B1(n10474), .B2(n13598), .A(n10473), .ZN(n10475) );
  OAI21_X1 U12992 ( .B1(n13582), .B2(n10513), .A(n10475), .ZN(P2_U3256) );
  INV_X1 U12993 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10641) );
  NOR2_X1 U12994 ( .A1(n11448), .A2(n10641), .ZN(n10482) );
  NAND2_X1 U12995 ( .A1(n10733), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10479) );
  OR2_X1 U12996 ( .A1(n10477), .A2(n10476), .ZN(n10478) );
  NAND2_X1 U12997 ( .A1(n10479), .A2(n10478), .ZN(n10480) );
  NOR2_X1 U12998 ( .A1(n14725), .A2(n10480), .ZN(n10481) );
  XOR2_X1 U12999 ( .A(n10488), .B(n10480), .Z(n14720) );
  NOR2_X1 U13000 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14720), .ZN(n14719) );
  NOR2_X1 U13001 ( .A1(n10481), .A2(n14719), .ZN(n10484) );
  AOI211_X1 U13002 ( .C1(n11448), .C2(n10641), .A(n10482), .B(n10484), .ZN(
        n10486) );
  NAND2_X1 U13003 ( .A1(n10642), .A2(n10641), .ZN(n10483) );
  OAI211_X1 U13004 ( .C1(n10642), .C2(n10641), .A(n10484), .B(n10483), .ZN(
        n10640) );
  INV_X1 U13005 ( .A(n10640), .ZN(n10485) );
  NOR3_X1 U13006 ( .A1(n10486), .A2(n10485), .A3(n14021), .ZN(n10497) );
  NAND2_X1 U13007 ( .A1(n10488), .A2(n10489), .ZN(n10490) );
  INV_X1 U13008 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15326) );
  INV_X1 U13009 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14649) );
  NOR2_X1 U13010 ( .A1(n11448), .A2(n14649), .ZN(n10491) );
  AOI21_X1 U13011 ( .B1(n11448), .B2(n14649), .A(n10491), .ZN(n10492) );
  NOR2_X1 U13012 ( .A1(n10493), .A2(n10492), .ZN(n10633) );
  AOI211_X1 U13013 ( .C1(n10493), .C2(n10492), .A(n10634), .B(n10633), .ZN(
        n10496) );
  NAND2_X1 U13014 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13843)
         );
  NAND2_X1 U13015 ( .A1(n14715), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n10494) );
  OAI211_X1 U13016 ( .C1(n14020), .C2(n10642), .A(n13843), .B(n10494), .ZN(
        n10495) );
  OR3_X1 U13017 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(P1_U3259) );
  AOI22_X1 U13018 ( .A1(n11409), .A2(n6923), .B1(n12554), .B2(n13949), .ZN(
        n10498) );
  XNOR2_X1 U13019 ( .A(n10498), .B(n12551), .ZN(n10784) );
  AOI22_X1 U13020 ( .A1(n11409), .A2(n12554), .B1(n12553), .B2(n13949), .ZN(
        n10783) );
  XNOR2_X1 U13021 ( .A(n10784), .B(n10783), .ZN(n10503) );
  AOI21_X1 U13022 ( .B1(n10503), .B2(n10502), .A(n6690), .ZN(n10510) );
  OAI21_X1 U13023 ( .B1(n13925), .B2(n10785), .A(n10504), .ZN(n10505) );
  AOI21_X1 U13024 ( .B1(n8890), .B2(n13950), .A(n10505), .ZN(n10506) );
  OAI21_X1 U13025 ( .B1(n10507), .B2(n14620), .A(n10506), .ZN(n10508) );
  AOI21_X1 U13026 ( .B1(n11409), .B2(n14616), .A(n10508), .ZN(n10509) );
  OAI21_X1 U13027 ( .B1(n10510), .B2(n13932), .A(n10509), .ZN(P1_U3221) );
  OAI211_X1 U13028 ( .C1(n13699), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        n10519) );
  INV_X1 U13029 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10514) );
  OAI22_X1 U13030 ( .A1(n10517), .A2(n13730), .B1(n14962), .B2(n10514), .ZN(
        n10515) );
  AOI21_X1 U13031 ( .B1(n10519), .B2(n14962), .A(n10515), .ZN(n10516) );
  INV_X1 U13032 ( .A(n10516), .ZN(P2_U3457) );
  OAI22_X1 U13033 ( .A1(n10517), .A2(n13668), .B1(n14972), .B2(n9630), .ZN(
        n10518) );
  AOI21_X1 U13034 ( .B1(n10519), .B2(n14972), .A(n10518), .ZN(n10520) );
  INV_X1 U13035 ( .A(n10520), .ZN(P2_U3508) );
  INV_X1 U13036 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14586) );
  AOI21_X1 U13037 ( .B1(n14586), .B2(n10523), .A(n10649), .ZN(n10537) );
  INV_X1 U13038 ( .A(n10662), .ZN(n10692) );
  XNOR2_X1 U13039 ( .A(n10655), .B(n10692), .ZN(n10525) );
  NAND2_X1 U13040 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10525), .ZN(n10656) );
  OAI21_X1 U13041 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10525), .A(n10656), 
        .ZN(n10535) );
  AND2_X1 U13042 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10701) );
  AOI21_X1 U13043 ( .B1(n14987), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n10701), 
        .ZN(n10526) );
  OAI21_X1 U13044 ( .B1(n14981), .B2(n10662), .A(n10526), .ZN(n10534) );
  INV_X1 U13045 ( .A(n10527), .ZN(n10528) );
  NOR2_X1 U13046 ( .A1(n10529), .A2(n10528), .ZN(n10531) );
  MUX2_X1 U13047 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12777), .Z(n10663) );
  XNOR2_X1 U13048 ( .A(n10663), .B(n10662), .ZN(n10530) );
  NOR2_X1 U13049 ( .A1(n10531), .A2(n10530), .ZN(n10665) );
  AOI21_X1 U13050 ( .B1(n10531), .B2(n10530), .A(n10665), .ZN(n10532) );
  NOR2_X1 U13051 ( .A1(n10532), .A2(n14983), .ZN(n10533) );
  AOI211_X1 U13052 ( .C1(n14990), .C2(n10535), .A(n10534), .B(n10533), .ZN(
        n10536) );
  OAI21_X1 U13053 ( .B1(n10537), .B2(n14994), .A(n10536), .ZN(P3_U3193) );
  AOI21_X1 U13054 ( .B1(n15001), .B2(n12643), .A(n10538), .ZN(n10552) );
  OR2_X1 U13055 ( .A1(n11198), .A2(n10539), .ZN(n10543) );
  OR2_X1 U13056 ( .A1(n11274), .A2(SI_10_), .ZN(n10542) );
  OR2_X1 U13057 ( .A1(n10868), .A2(n10540), .ZN(n10541) );
  NAND2_X1 U13058 ( .A1(n12648), .A2(n15009), .ZN(n10551) );
  NAND2_X1 U13059 ( .A1(n6530), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13060 ( .A1(n10544), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U13061 ( .A1(n10696), .A2(n10545), .ZN(n14584) );
  NAND2_X1 U13062 ( .A1(n11154), .A2(n14584), .ZN(n10548) );
  NAND2_X1 U13063 ( .A1(n6532), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13064 ( .A1(n11216), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U13065 ( .A1(n15000), .A2(n12663), .ZN(n10550) );
  NAND3_X1 U13066 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n10559) );
  XNOR2_X1 U13067 ( .A(n15009), .B(n11786), .ZN(n10688) );
  XNOR2_X1 U13068 ( .A(n10688), .B(n15019), .ZN(n10557) );
  NOR2_X1 U13069 ( .A1(n10553), .A2(n15001), .ZN(n10554) );
  OR2_X1 U13070 ( .A1(n10555), .A2(n10554), .ZN(n10556) );
  AOI211_X1 U13071 ( .C1(n10557), .C2(n10556), .A(n12672), .B(n10689), .ZN(
        n10558) );
  AOI211_X1 U13072 ( .C1(n15010), .C2(n12670), .A(n10559), .B(n10558), .ZN(
        n10560) );
  INV_X1 U13073 ( .A(n10560), .ZN(P3_U3157) );
  NAND2_X1 U13074 ( .A1(n13257), .A2(n13542), .ZN(n10562) );
  INV_X1 U13075 ( .A(n10562), .ZN(n10565) );
  XNOR2_X1 U13076 ( .A(n13587), .B(n6529), .ZN(n10564) );
  NOR2_X1 U13077 ( .A1(n11134), .A2(n10561), .ZN(n10563) );
  XNOR2_X1 U13078 ( .A(n10564), .B(n10562), .ZN(n11135) );
  XNOR2_X1 U13079 ( .A(n14819), .B(n6529), .ZN(n10568) );
  AND2_X1 U13080 ( .A1(n13256), .A2(n13542), .ZN(n10566) );
  NAND2_X1 U13081 ( .A1(n10568), .A2(n10566), .ZN(n10570) );
  OAI21_X1 U13082 ( .B1(n10568), .B2(n10566), .A(n10570), .ZN(n14815) );
  NOR2_X1 U13083 ( .A1(n13213), .A2(n10567), .ZN(n10569) );
  AOI22_X1 U13084 ( .A1(n14812), .A2(n13227), .B1(n10569), .B2(n10568), .ZN(
        n10580) );
  XNOR2_X1 U13085 ( .A(n12139), .B(n12356), .ZN(n11110) );
  NAND2_X1 U13086 ( .A1(n13255), .A2(n13542), .ZN(n11109) );
  XNOR2_X1 U13087 ( .A(n11110), .B(n11109), .ZN(n10572) );
  INV_X1 U13088 ( .A(n10572), .ZN(n10579) );
  INV_X1 U13089 ( .A(n10570), .ZN(n10571) );
  NAND2_X1 U13090 ( .A1(n11108), .A2(n13227), .ZN(n10578) );
  NOR2_X1 U13091 ( .A1(n14821), .A2(n10889), .ZN(n10576) );
  NAND2_X1 U13092 ( .A1(n13254), .A2(n13230), .ZN(n10574) );
  NAND2_X1 U13093 ( .A1(n13256), .A2(n13231), .ZN(n10573) );
  AND2_X1 U13094 ( .A1(n10574), .A2(n10573), .ZN(n10885) );
  OAI22_X1 U13095 ( .A1(n14811), .A2(n10885), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13312), .ZN(n10575) );
  AOI211_X1 U13096 ( .C1(n12139), .C2(n14818), .A(n10576), .B(n10575), .ZN(
        n10577) );
  OAI211_X1 U13097 ( .C1(n10580), .C2(n10579), .A(n10578), .B(n10577), .ZN(
        P2_U3187) );
  INV_X1 U13098 ( .A(n10581), .ZN(n10589) );
  NAND2_X1 U13099 ( .A1(n15307), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13100 ( .A1(n10586), .A2(n10953), .ZN(n10587) );
  XNOR2_X1 U13101 ( .A(n10764), .B(n11801), .ZN(n11232) );
  INV_X1 U13102 ( .A(n11232), .ZN(n10588) );
  INV_X1 U13103 ( .A(SI_24_), .ZN(n11233) );
  OAI222_X1 U13104 ( .A1(P3_U3151), .A2(n10589), .B1(n13120), .B2(n10588), 
        .C1(n11233), .C2(n13115), .ZN(P3_U3271) );
  NAND2_X1 U13105 ( .A1(n10591), .A2(n10590), .ZN(n10593) );
  OR2_X1 U13106 ( .A1(n14672), .A2(n13946), .ZN(n10592) );
  NAND2_X1 U13107 ( .A1(n10594), .A2(n11622), .ZN(n10596) );
  AOI22_X1 U13108 ( .A1(n14006), .A2(n11455), .B1(n11613), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10595) );
  INV_X1 U13109 ( .A(n14506), .ZN(n11428) );
  XNOR2_X1 U13110 ( .A(n11428), .B(n13945), .ZN(n14485) );
  INV_X1 U13111 ( .A(n14485), .ZN(n14491) );
  NAND2_X1 U13112 ( .A1(n14506), .A2(n12410), .ZN(n10597) );
  NAND2_X1 U13113 ( .A1(n10598), .A2(n11622), .ZN(n10601) );
  AOI22_X1 U13114 ( .A1(n10599), .A2(n11455), .B1(n11613), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13115 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  NAND2_X1 U13116 ( .A1(n10618), .A2(n10604), .ZN(n13885) );
  OR2_X1 U13117 ( .A1(n13885), .A2(n11608), .ZN(n10610) );
  INV_X1 U13118 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10605) );
  OR2_X1 U13119 ( .A1(n11607), .A2(n10605), .ZN(n10609) );
  OR2_X1 U13120 ( .A1(n11630), .A2(n9593), .ZN(n10608) );
  OR2_X1 U13121 ( .A1(n11583), .A2(n10606), .ZN(n10607) );
  NAND4_X1 U13122 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n13944) );
  XNOR2_X1 U13123 ( .A(n14666), .B(n14249), .ZN(n11661) );
  XNOR2_X1 U13124 ( .A(n10751), .B(n7329), .ZN(n14664) );
  INV_X1 U13125 ( .A(n13946), .ZN(n13824) );
  OR2_X1 U13126 ( .A1(n14672), .A2(n13824), .ZN(n10612) );
  NAND2_X1 U13127 ( .A1(n10613), .A2(n10612), .ZN(n14492) );
  NAND2_X1 U13128 ( .A1(n14492), .A2(n14485), .ZN(n10615) );
  NAND2_X1 U13129 ( .A1(n14506), .A2(n13945), .ZN(n10614) );
  NAND2_X1 U13130 ( .A1(n10615), .A2(n10614), .ZN(n10729) );
  XNOR2_X1 U13131 ( .A(n10729), .B(n11661), .ZN(n10616) );
  NAND2_X1 U13132 ( .A1(n10616), .A2(n14494), .ZN(n10627) );
  AND2_X1 U13133 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  OR2_X1 U13134 ( .A1(n10619), .A2(n10740), .ZN(n14252) );
  INV_X1 U13135 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10620) );
  OR2_X1 U13136 ( .A1(n11607), .A2(n10620), .ZN(n10623) );
  OR2_X1 U13137 ( .A1(n11583), .A2(n10621), .ZN(n10622) );
  AND2_X1 U13138 ( .A1(n10623), .A2(n10622), .ZN(n10625) );
  OR2_X1 U13139 ( .A1(n11630), .A2(n9693), .ZN(n10624) );
  OAI211_X1 U13140 ( .C1(n14252), .C2(n11608), .A(n10625), .B(n10624), .ZN(
        n13943) );
  NAND2_X1 U13141 ( .A1(n13943), .A2(n14222), .ZN(n10626) );
  NAND2_X1 U13142 ( .A1(n10627), .A2(n10626), .ZN(n14671) );
  NOR2_X1 U13143 ( .A1(n12410), .A2(n14631), .ZN(n14665) );
  OAI21_X1 U13144 ( .B1(n14671), .B2(n14665), .A(n14639), .ZN(n10632) );
  OAI22_X1 U13145 ( .A1(n14639), .A2(n9593), .B1(n13885), .B2(n14642), .ZN(
        n10630) );
  NAND2_X1 U13146 ( .A1(n14666), .A2(n14487), .ZN(n10628) );
  NAND3_X1 U13147 ( .A1(n14253), .A2(n8808), .A3(n10628), .ZN(n14668) );
  NOR2_X1 U13148 ( .A1(n14668), .A2(n14489), .ZN(n10629) );
  AOI211_X1 U13149 ( .C1(n14259), .C2(n14666), .A(n10630), .B(n10629), .ZN(
        n10631) );
  OAI211_X1 U13150 ( .C1(n14247), .C2(n14664), .A(n10632), .B(n10631), .ZN(
        P1_U3280) );
  AOI21_X1 U13151 ( .B1(n11448), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10633), 
        .ZN(n10636) );
  XNOR2_X1 U13152 ( .A(n11454), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10635) );
  NOR2_X1 U13153 ( .A1(n10636), .A2(n10635), .ZN(n10827) );
  AOI211_X1 U13154 ( .C1(n10636), .C2(n10635), .A(n10634), .B(n10827), .ZN(
        n10639) );
  NAND2_X1 U13155 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13857)
         );
  NAND2_X1 U13156 ( .A1(n14715), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n10637) );
  OAI211_X1 U13157 ( .C1(n14020), .C2(n10832), .A(n13857), .B(n10637), .ZN(
        n10638) );
  NOR2_X1 U13158 ( .A1(n10639), .A2(n10638), .ZN(n10647) );
  OAI21_X1 U13159 ( .B1(n10642), .B2(n10641), .A(n10640), .ZN(n10645) );
  INV_X1 U13160 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13161 ( .A1(n10832), .A2(n10831), .ZN(n10643) );
  AOI21_X1 U13162 ( .B1(n10831), .B2(n10832), .A(n10643), .ZN(n10644) );
  NAND2_X1 U13163 ( .A1(n10644), .A2(n10645), .ZN(n10830) );
  OAI211_X1 U13164 ( .C1(n10645), .C2(n10644), .A(n10830), .B(n14728), .ZN(
        n10646) );
  NAND2_X1 U13165 ( .A1(n10647), .A2(n10646), .ZN(P1_U3260) );
  NOR2_X1 U13166 ( .A1(n10692), .A2(n10648), .ZN(n10650) );
  NAND2_X1 U13167 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n10962), .ZN(n10651) );
  OAI21_X1 U13168 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n10962), .A(n10651), 
        .ZN(n10652) );
  AOI21_X1 U13169 ( .B1(n10653), .B2(n10652), .A(n10955), .ZN(n10672) );
  INV_X1 U13170 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U13171 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10962), .B1(n10654), 
        .B2(n14597), .ZN(n10659) );
  NAND2_X1 U13172 ( .A1(n10662), .A2(n10655), .ZN(n10657) );
  NAND2_X1 U13173 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  OAI21_X1 U13174 ( .B1(n10659), .B2(n10658), .A(n10963), .ZN(n10670) );
  INV_X1 U13175 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10660) );
  NOR2_X1 U13176 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10660), .ZN(n10723) );
  AOI21_X1 U13177 ( .B1(n14987), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n10723), 
        .ZN(n10661) );
  OAI21_X1 U13178 ( .B1(n14981), .B2(n10962), .A(n10661), .ZN(n10669) );
  MUX2_X1 U13179 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12777), .Z(n10959) );
  XNOR2_X1 U13180 ( .A(n10959), .B(n10962), .ZN(n10667) );
  NOR2_X1 U13181 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  OR2_X1 U13182 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  NOR3_X1 U13183 ( .A1(n10665), .A2(n10664), .A3(n10667), .ZN(n10958) );
  AOI211_X1 U13184 ( .C1(n10667), .C2(n10666), .A(n14983), .B(n10958), .ZN(
        n10668) );
  AOI211_X1 U13185 ( .C1(n14990), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10671) );
  OAI21_X1 U13186 ( .B1(n10672), .B2(n14994), .A(n10671), .ZN(P3_U3194) );
  XNOR2_X1 U13187 ( .A(n10673), .B(n12278), .ZN(n13602) );
  AOI21_X1 U13188 ( .B1(n10674), .B2(n13601), .A(n14896), .ZN(n10675) );
  AND2_X1 U13189 ( .A1(n10675), .A2(n10775), .ZN(n13603) );
  OAI211_X1 U13190 ( .C1(n10677), .C2(n12278), .A(n10676), .B(n14892), .ZN(
        n10679) );
  NAND2_X1 U13191 ( .A1(n10679), .A2(n10678), .ZN(n13594) );
  AOI211_X1 U13192 ( .C1(n14927), .C2(n13602), .A(n13603), .B(n13594), .ZN(
        n10684) );
  INV_X1 U13193 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10680) );
  NOR2_X1 U13194 ( .A1(n14962), .A2(n10680), .ZN(n10681) );
  AOI21_X1 U13195 ( .B1(n13601), .B2(n13744), .A(n10681), .ZN(n10682) );
  OAI21_X1 U13196 ( .B1(n10684), .B2(n14961), .A(n10682), .ZN(P2_U3460) );
  AOI22_X1 U13197 ( .A1(n13601), .A2(n13692), .B1(n14970), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n10683) );
  OAI21_X1 U13198 ( .B1(n10684), .B2(n14970), .A(n10683), .ZN(P2_U3509) );
  NAND2_X1 U13199 ( .A1(n11525), .A2(n13755), .ZN(n10686) );
  OR2_X1 U13200 ( .A1(n10685), .A2(P2_U3088), .ZN(n12308) );
  OAI211_X1 U13201 ( .C1(n15307), .C2(n13749), .A(n10686), .B(n12308), .ZN(
        P2_U3304) );
  INV_X1 U13202 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U13203 ( .A1(n11525), .A2(n11731), .ZN(n10687) );
  OAI211_X1 U13204 ( .C1(n11526), .C2(n11751), .A(n10687), .B(n11692), .ZN(
        P1_U3332) );
  INV_X1 U13205 ( .A(n10688), .ZN(n10690) );
  OR2_X1 U13206 ( .A1(n11198), .A2(n10691), .ZN(n10695) );
  OR2_X1 U13207 ( .A1(n11274), .A2(SI_11_), .ZN(n10694) );
  OR2_X1 U13208 ( .A1(n10868), .A2(n10692), .ZN(n10693) );
  XNOR2_X1 U13209 ( .A(n11881), .B(n11786), .ZN(n10708) );
  XNOR2_X1 U13210 ( .A(n10710), .B(n15000), .ZN(n10706) );
  NOR2_X1 U13211 ( .A1(n12666), .A2(n14583), .ZN(n10705) );
  NAND2_X1 U13212 ( .A1(n6530), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n10700) );
  OR2_X1 U13213 ( .A1(n7691), .A2(n10717), .ZN(n12978) );
  NAND2_X1 U13214 ( .A1(n11154), .A2(n12978), .ZN(n10699) );
  NAND2_X1 U13215 ( .A1(n6531), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U13216 ( .A1(n11216), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10697) );
  AOI21_X1 U13217 ( .B1(n10919), .B2(n12643), .A(n10701), .ZN(n10703) );
  NAND2_X1 U13218 ( .A1(n12670), .A2(n14584), .ZN(n10702) );
  OAI211_X1 U13219 ( .C1(n14581), .C2(n12646), .A(n10703), .B(n10702), .ZN(
        n10704) );
  AOI211_X1 U13220 ( .C1(n10706), .C2(n12651), .A(n10705), .B(n10704), .ZN(
        n10707) );
  INV_X1 U13221 ( .A(n10707), .ZN(P3_U3176) );
  OR2_X1 U13222 ( .A1(n10711), .A2(n11198), .ZN(n10714) );
  OR2_X1 U13223 ( .A1(n11274), .A2(n10712), .ZN(n10713) );
  OAI211_X1 U13224 ( .C1(n10868), .C2(n10962), .A(n10714), .B(n10713), .ZN(
        n12981) );
  XNOR2_X1 U13225 ( .A(n12981), .B(n11786), .ZN(n10865) );
  XNOR2_X1 U13226 ( .A(n14563), .B(n10865), .ZN(n10715) );
  XNOR2_X1 U13227 ( .A(n10864), .B(n10715), .ZN(n10728) );
  OR2_X1 U13228 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  NAND2_X1 U13229 ( .A1(n11154), .A2(n7692), .ZN(n10722) );
  NAND2_X1 U13230 ( .A1(n6530), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U13231 ( .A1(n6532), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n10720) );
  NAND2_X1 U13232 ( .A1(n11216), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13233 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n12975) );
  NAND2_X1 U13234 ( .A1(n12670), .A2(n12978), .ZN(n10725) );
  AOI21_X1 U13235 ( .B1(n15000), .B2(n12643), .A(n10723), .ZN(n10724) );
  OAI211_X1 U13236 ( .C1(n10976), .C2(n12646), .A(n10725), .B(n10724), .ZN(
        n10726) );
  AOI21_X1 U13237 ( .B1(n12648), .B2(n12981), .A(n10726), .ZN(n10727) );
  OAI21_X1 U13238 ( .B1(n10728), .B2(n12672), .A(n10727), .ZN(P3_U3164) );
  NAND2_X1 U13239 ( .A1(n10729), .A2(n7329), .ZN(n10731) );
  OR2_X1 U13240 ( .A1(n14666), .A2(n14249), .ZN(n10730) );
  NAND2_X1 U13241 ( .A1(n10731), .A2(n10730), .ZN(n14248) );
  NAND2_X1 U13242 ( .A1(n10732), .A2(n11622), .ZN(n10735) );
  AOI22_X1 U13243 ( .A1(n10733), .A2(n11455), .B1(n11613), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10734) );
  INV_X1 U13244 ( .A(n13943), .ZN(n13882) );
  NAND2_X1 U13245 ( .A1(n14258), .A2(n13882), .ZN(n11431) );
  INV_X1 U13246 ( .A(n11430), .ZN(n10736) );
  NAND2_X1 U13247 ( .A1(n10737), .A2(n11622), .ZN(n10739) );
  AOI22_X1 U13248 ( .A1(n11613), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11455), 
        .B2(n14725), .ZN(n10738) );
  NOR2_X1 U13249 ( .A1(n10740), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10741) );
  OR2_X1 U13250 ( .A1(n10744), .A2(n10741), .ZN(n13928) );
  AOI22_X1 U13251 ( .A1(n6963), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n11582), 
        .B2(P1_REG0_REG_15__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13252 ( .A1(n11606), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n10742) );
  OAI211_X1 U13253 ( .C1(n13928), .C2(n11608), .A(n10743), .B(n10742), .ZN(
        n13942) );
  INV_X1 U13254 ( .A(n13942), .ZN(n14630) );
  NAND2_X1 U13255 ( .A1(n13930), .A2(n14630), .ZN(n11445) );
  XNOR2_X1 U13256 ( .A(n11695), .B(n10755), .ZN(n10750) );
  OR2_X1 U13257 ( .A1(n10744), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U13258 ( .A1(n11459), .A2(n10745), .ZN(n14641) );
  AOI22_X1 U13259 ( .A1(n6963), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n11606), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13260 ( .A1(n11582), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n10746) );
  OAI211_X1 U13261 ( .C1(n14641), .C2(n11608), .A(n10747), .B(n10746), .ZN(
        n13941) );
  NAND2_X1 U13262 ( .A1(n13941), .A2(n14222), .ZN(n10748) );
  OAI21_X1 U13263 ( .B1(n13882), .B2(n14631), .A(n10748), .ZN(n10749) );
  AOI21_X1 U13264 ( .B1(n10750), .B2(n14494), .A(n10749), .ZN(n14654) );
  NAND2_X1 U13265 ( .A1(n14258), .A2(n13943), .ZN(n10754) );
  NAND2_X1 U13266 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  NAND2_X1 U13267 ( .A1(n11702), .A2(n10757), .ZN(n14652) );
  AOI21_X1 U13268 ( .B1(n13930), .B2(n14254), .A(n14674), .ZN(n10758) );
  NAND2_X1 U13269 ( .A1(n10758), .A2(n14623), .ZN(n14650) );
  INV_X1 U13270 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10759) );
  OAI22_X1 U13271 ( .A1(n14639), .A2(n10759), .B1(n13928), .B2(n14642), .ZN(
        n10760) );
  AOI21_X1 U13272 ( .B1(n13930), .B2(n14259), .A(n10760), .ZN(n10761) );
  OAI21_X1 U13273 ( .B1(n14650), .B2(n14489), .A(n10761), .ZN(n10762) );
  AOI21_X1 U13274 ( .B1(n14652), .B2(n14262), .A(n10762), .ZN(n10763) );
  OAI21_X1 U13275 ( .B1(n14654), .B2(n14747), .A(n10763), .ZN(P1_U3278) );
  INV_X1 U13276 ( .A(SI_25_), .ZN(n11247) );
  XNOR2_X1 U13277 ( .A(n11062), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n10766) );
  XNOR2_X1 U13278 ( .A(n10797), .B(n10766), .ZN(n11246) );
  INV_X1 U13279 ( .A(n11246), .ZN(n10767) );
  OAI222_X1 U13280 ( .A1(n13122), .A2(n11247), .B1(P3_U3151), .B2(n10768), 
        .C1(n13120), .C2(n10767), .ZN(P3_U3270) );
  XNOR2_X1 U13281 ( .A(n10769), .B(n12279), .ZN(n10860) );
  INV_X1 U13282 ( .A(n10860), .ZN(n10782) );
  INV_X1 U13283 ( .A(n10770), .ZN(n10820) );
  AOI21_X1 U13284 ( .B1(n10772), .B2(n10771), .A(n10820), .ZN(n10774) );
  OAI21_X1 U13285 ( .B1(n10774), .B2(n13509), .A(n10773), .ZN(n10858) );
  AOI21_X1 U13286 ( .B1(n10775), .B2(n12115), .A(n14896), .ZN(n10776) );
  NAND2_X1 U13287 ( .A1(n10776), .A2(n10815), .ZN(n10856) );
  OAI22_X1 U13288 ( .A1(n13598), .A2(n11074), .B1(n10777), .B2(n13595), .ZN(
        n10778) );
  AOI21_X1 U13289 ( .B1(n12115), .B2(n13600), .A(n10778), .ZN(n10779) );
  OAI21_X1 U13290 ( .B1(n10856), .B2(n13578), .A(n10779), .ZN(n10780) );
  AOI21_X1 U13291 ( .B1(n10858), .B2(n13598), .A(n10780), .ZN(n10781) );
  OAI21_X1 U13292 ( .B1(n13582), .B2(n10782), .A(n10781), .ZN(P2_U3254) );
  NOR2_X1 U13293 ( .A1(n12525), .A2(n10785), .ZN(n10786) );
  AOI21_X1 U13294 ( .B1(n11413), .B2(n12554), .A(n10786), .ZN(n10842) );
  XNOR2_X1 U13295 ( .A(n10839), .B(n10842), .ZN(n10789) );
  AOI22_X1 U13296 ( .A1(n11413), .A2(n6923), .B1(n12554), .B2(n13948), .ZN(
        n10787) );
  XOR2_X1 U13297 ( .A(n12551), .B(n10787), .Z(n10788) );
  NAND2_X1 U13298 ( .A1(n10789), .A2(n10788), .ZN(n10840) );
  OAI211_X1 U13299 ( .C1(n10789), .C2(n10788), .A(n10840), .B(n14612), .ZN(
        n10795) );
  NOR2_X1 U13300 ( .A1(n14620), .A2(n10790), .ZN(n10793) );
  OAI21_X1 U13301 ( .B1(n13925), .B2(n10846), .A(n10791), .ZN(n10792) );
  AOI211_X1 U13302 ( .C1(n8890), .C2(n13949), .A(n10793), .B(n10792), .ZN(
        n10794) );
  OAI211_X1 U13303 ( .C1(n14784), .C2(n13921), .A(n10795), .B(n10794), .ZN(
        P1_U3231) );
  NAND2_X1 U13304 ( .A1(n11062), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10796) );
  INV_X1 U13305 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U13306 ( .A1(n15281), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10798) );
  XNOR2_X1 U13307 ( .A(n13765), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n10799) );
  XNOR2_X1 U13308 ( .A(n11142), .B(n10799), .ZN(n11257) );
  INV_X1 U13309 ( .A(n11257), .ZN(n10802) );
  INV_X1 U13310 ( .A(SI_26_), .ZN(n11258) );
  INV_X1 U13311 ( .A(n10800), .ZN(n10801) );
  OAI222_X1 U13312 ( .A1(n13120), .A2(n10802), .B1(n13122), .B2(n11258), .C1(
        P3_U3151), .C2(n10801), .ZN(P3_U3269) );
  XOR2_X1 U13313 ( .A(n10803), .B(n12281), .Z(n10900) );
  INV_X1 U13314 ( .A(n10900), .ZN(n10813) );
  INV_X1 U13315 ( .A(n12281), .ZN(n10805) );
  NAND3_X1 U13316 ( .A1(n10821), .A2(n10805), .A3(n10804), .ZN(n10806) );
  NAND3_X1 U13317 ( .A1(n10807), .A2(n14892), .A3(n10806), .ZN(n10808) );
  AOI22_X1 U13318 ( .A1(n13231), .A2(n13257), .B1(n13255), .B2(n13230), .ZN(
        n14810) );
  NAND2_X1 U13319 ( .A1(n10808), .A2(n14810), .ZN(n10898) );
  OAI211_X1 U13320 ( .C1(n10818), .C2(n10897), .A(n13557), .B(n10888), .ZN(
        n10896) );
  OAI22_X1 U13321 ( .A1(n13598), .A2(n11073), .B1(n14822), .B2(n13595), .ZN(
        n10809) );
  AOI21_X1 U13322 ( .B1(n14819), .B2(n13600), .A(n10809), .ZN(n10810) );
  OAI21_X1 U13323 ( .B1(n10896), .B2(n13578), .A(n10810), .ZN(n10811) );
  AOI21_X1 U13324 ( .B1(n10898), .B2(n13598), .A(n10811), .ZN(n10812) );
  OAI21_X1 U13325 ( .B1(n10813), .B2(n13582), .A(n10812), .ZN(P2_U3252) );
  XNOR2_X1 U13326 ( .A(n10814), .B(n12277), .ZN(n13588) );
  NAND2_X1 U13327 ( .A1(n10815), .A2(n13587), .ZN(n10816) );
  NAND2_X1 U13328 ( .A1(n10816), .A2(n13557), .ZN(n10817) );
  NOR2_X1 U13329 ( .A1(n10818), .A2(n10817), .ZN(n13589) );
  OAI21_X1 U13330 ( .B1(n10820), .B2(n10819), .A(n12277), .ZN(n10822) );
  NAND3_X1 U13331 ( .A1(n10822), .A2(n14892), .A3(n10821), .ZN(n10823) );
  AOI22_X1 U13332 ( .A1(n13231), .A2(n13258), .B1(n13256), .B2(n13230), .ZN(
        n11133) );
  NAND2_X1 U13333 ( .A1(n10823), .A2(n11133), .ZN(n13583) );
  AOI211_X1 U13334 ( .C1(n14927), .C2(n13588), .A(n13589), .B(n13583), .ZN(
        n10826) );
  AOI22_X1 U13335 ( .A1(n13587), .A2(n13692), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n14970), .ZN(n10824) );
  OAI21_X1 U13336 ( .B1(n10826), .B2(n14970), .A(n10824), .ZN(P2_U3511) );
  AOI22_X1 U13337 ( .A1(n13587), .A2(n13744), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n14961), .ZN(n10825) );
  OAI21_X1 U13338 ( .B1(n10826), .B2(n14961), .A(n10825), .ZN(P2_U3466) );
  AOI21_X1 U13339 ( .B1(n11454), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10827), 
        .ZN(n10828) );
  OAI21_X1 U13340 ( .B1(n10829), .B2(P1_REG1_REG_18__SCAN_IN), .A(n14727), 
        .ZN(n10838) );
  OAI21_X1 U13341 ( .B1(n10832), .B2(n10831), .A(n10830), .ZN(n14012) );
  XNOR2_X1 U13342 ( .A(n14012), .B(n14011), .ZN(n14013) );
  XNOR2_X1 U13343 ( .A(n14013), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13344 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13904)
         );
  NAND2_X1 U13345 ( .A1(n14715), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n10833) );
  OAI211_X1 U13346 ( .C1(n14020), .C2(n10834), .A(n13904), .B(n10833), .ZN(
        n10835) );
  AOI21_X1 U13347 ( .B1(n14728), .B2(n10836), .A(n10835), .ZN(n10837) );
  OAI21_X1 U13348 ( .B1(n10838), .B2(n14018), .A(n10837), .ZN(P1_U3261) );
  INV_X1 U13349 ( .A(n10839), .ZN(n10841) );
  NAND2_X1 U13350 ( .A1(n14790), .A2(n6923), .ZN(n10844) );
  NAND2_X1 U13351 ( .A1(n12554), .A2(n13947), .ZN(n10843) );
  NAND2_X1 U13352 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  XNOR2_X1 U13353 ( .A(n10845), .B(n12522), .ZN(n12413) );
  NOR2_X1 U13354 ( .A1(n12525), .A2(n10846), .ZN(n10847) );
  AOI21_X1 U13355 ( .B1(n14790), .B2(n12554), .A(n10847), .ZN(n12412) );
  INV_X1 U13356 ( .A(n12412), .ZN(n12414) );
  XNOR2_X1 U13357 ( .A(n12413), .B(n12414), .ZN(n10848) );
  XNOR2_X1 U13358 ( .A(n12417), .B(n10848), .ZN(n10855) );
  OAI21_X1 U13359 ( .B1(n13925), .B2(n13824), .A(n10849), .ZN(n10850) );
  AOI21_X1 U13360 ( .B1(n8890), .B2(n13948), .A(n10850), .ZN(n10851) );
  OAI21_X1 U13361 ( .B1(n10852), .B2(n14620), .A(n10851), .ZN(n10853) );
  AOI21_X1 U13362 ( .B1(n14790), .B2(n14616), .A(n10853), .ZN(n10854) );
  OAI21_X1 U13363 ( .B1(n10855), .B2(n13932), .A(n10854), .ZN(P1_U3217) );
  INV_X1 U13364 ( .A(n12115), .ZN(n10857) );
  OAI21_X1 U13365 ( .B1(n10857), .B2(n14946), .A(n10856), .ZN(n10859) );
  AOI211_X1 U13366 ( .C1(n14927), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        n10863) );
  NAND2_X1 U13367 ( .A1(n14961), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10861) );
  OAI21_X1 U13368 ( .B1(n10863), .B2(n14961), .A(n10861), .ZN(P2_U3463) );
  NAND2_X1 U13369 ( .A1(n14970), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10862) );
  OAI21_X1 U13370 ( .B1(n10863), .B2(n14970), .A(n10862), .ZN(P2_U3510) );
  NAND2_X1 U13371 ( .A1(n14581), .A2(n10865), .ZN(n10866) );
  NAND2_X1 U13372 ( .A1(n10867), .A2(n11971), .ZN(n10870) );
  INV_X1 U13373 ( .A(n11274), .ZN(n11177) );
  INV_X1 U13374 ( .A(n10868), .ZN(n11175) );
  AOI22_X1 U13375 ( .A1(n11177), .A2(SI_13_), .B1(n11175), .B2(n12707), .ZN(
        n10869) );
  XNOR2_X1 U13376 ( .A(n14568), .B(n11786), .ZN(n10977) );
  XNOR2_X1 U13377 ( .A(n10977), .B(n12975), .ZN(n10871) );
  XNOR2_X1 U13378 ( .A(n10980), .B(n10871), .ZN(n10882) );
  NAND2_X1 U13379 ( .A1(n10872), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10873) );
  NAND2_X1 U13380 ( .A1(n10935), .A2(n10873), .ZN(n10987) );
  NAND2_X1 U13381 ( .A1(n11154), .A2(n10987), .ZN(n10877) );
  NAND2_X1 U13382 ( .A1(n6530), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13383 ( .A1(n6532), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U13384 ( .A1(n11216), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n10874) );
  AND2_X1 U13385 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n10967) );
  AOI21_X1 U13386 ( .B1(n14563), .B2(n12643), .A(n10967), .ZN(n10879) );
  NAND2_X1 U13387 ( .A1(n12670), .A2(n7692), .ZN(n10878) );
  OAI211_X1 U13388 ( .C1(n10974), .C2(n12646), .A(n10879), .B(n10878), .ZN(
        n10880) );
  AOI21_X1 U13389 ( .B1(n12648), .B2(n14568), .A(n10880), .ZN(n10881) );
  OAI21_X1 U13390 ( .B1(n10882), .B2(n12672), .A(n10881), .ZN(P3_U3174) );
  XNOR2_X1 U13391 ( .A(n10883), .B(n12284), .ZN(n11055) );
  INV_X1 U13392 ( .A(n11055), .ZN(n10895) );
  XNOR2_X1 U13393 ( .A(n10884), .B(n12284), .ZN(n10886) );
  OAI21_X1 U13394 ( .B1(n10886), .B2(n13509), .A(n10885), .ZN(n11053) );
  NAND2_X1 U13395 ( .A1(n11053), .A2(n13598), .ZN(n10894) );
  INV_X1 U13396 ( .A(n10998), .ZN(n10887) );
  AOI211_X1 U13397 ( .C1(n12139), .C2(n10888), .A(n14896), .B(n10887), .ZN(
        n11054) );
  INV_X1 U13398 ( .A(n12139), .ZN(n11060) );
  NOR2_X1 U13399 ( .A1(n11060), .A2(n14879), .ZN(n10892) );
  OAI22_X1 U13400 ( .A1(n13598), .A2(n10890), .B1(n10889), .B2(n13595), .ZN(
        n10891) );
  AOI211_X1 U13401 ( .C1(n11054), .C2(n14874), .A(n10892), .B(n10891), .ZN(
        n10893) );
  OAI211_X1 U13402 ( .C1(n10895), .C2(n13582), .A(n10894), .B(n10893), .ZN(
        P2_U3251) );
  OAI21_X1 U13403 ( .B1(n10897), .B2(n14946), .A(n10896), .ZN(n10899) );
  AOI211_X1 U13404 ( .C1(n10900), .C2(n14927), .A(n10899), .B(n10898), .ZN(
        n10903) );
  NAND2_X1 U13405 ( .A1(n14961), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10901) );
  OAI21_X1 U13406 ( .B1(n10903), .B2(n14961), .A(n10901), .ZN(P2_U3469) );
  NAND2_X1 U13407 ( .A1(n14970), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10902) );
  OAI21_X1 U13408 ( .B1(n10903), .B2(n14970), .A(n10902), .ZN(P2_U3512) );
  NAND2_X1 U13409 ( .A1(n15001), .A2(n15026), .ZN(n10905) );
  INV_X1 U13410 ( .A(n15001), .ZN(n11871) );
  INV_X1 U13411 ( .A(n15026), .ZN(n11872) );
  NAND2_X1 U13412 ( .A1(n11871), .A2(n11872), .ZN(n10906) );
  NAND2_X1 U13413 ( .A1(n15019), .A2(n15009), .ZN(n11877) );
  NAND2_X1 U13414 ( .A1(n10919), .A2(n10907), .ZN(n11878) );
  NAND2_X1 U13415 ( .A1(n11877), .A2(n11878), .ZN(n14996) );
  XNOR2_X1 U13416 ( .A(n15000), .B(n14583), .ZN(n14578) );
  NAND2_X1 U13417 ( .A1(n11882), .A2(n11881), .ZN(n11887) );
  NAND2_X1 U13418 ( .A1(n14581), .A2(n12981), .ZN(n11888) );
  INV_X1 U13419 ( .A(n12981), .ZN(n10910) );
  NAND2_X1 U13420 ( .A1(n14563), .A2(n10910), .ZN(n11889) );
  NAND2_X1 U13421 ( .A1(n12980), .A2(n12979), .ZN(n10911) );
  NAND2_X1 U13422 ( .A1(n10912), .A2(n11971), .ZN(n10914) );
  AOI22_X1 U13423 ( .A1(n11177), .A2(SI_14_), .B1(n11175), .B2(n12699), .ZN(
        n10913) );
  NAND2_X1 U13424 ( .A1(n11029), .A2(n10974), .ZN(n11899) );
  NAND2_X1 U13425 ( .A1(n11900), .A2(n11899), .ZN(n11896) );
  INV_X1 U13426 ( .A(n11896), .ZN(n11998) );
  XNOR2_X1 U13427 ( .A(n11017), .B(n11998), .ZN(n10952) );
  NOR2_X1 U13428 ( .A1(n15050), .A2(n15025), .ZN(n15034) );
  INV_X1 U13429 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U13430 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  XNOR2_X1 U13431 ( .A(n15001), .B(n15026), .ZN(n15015) );
  NAND2_X1 U13432 ( .A1(n11882), .A2(n14583), .ZN(n10924) );
  INV_X1 U13433 ( .A(n10924), .ZN(n10923) );
  AND2_X1 U13434 ( .A1(n15000), .A2(n11881), .ZN(n10921) );
  NAND2_X1 U13435 ( .A1(n10919), .A2(n15009), .ZN(n14576) );
  INV_X1 U13436 ( .A(n14576), .ZN(n10920) );
  NOR2_X1 U13437 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  INV_X1 U13438 ( .A(n10929), .ZN(n10926) );
  AND2_X1 U13439 ( .A1(n14996), .A2(n10924), .ZN(n10925) );
  INV_X1 U13440 ( .A(n12979), .ZN(n10927) );
  NAND2_X1 U13441 ( .A1(n15001), .A2(n11872), .ZN(n14574) );
  AND2_X1 U13442 ( .A1(n14574), .A2(n10929), .ZN(n12969) );
  NAND2_X1 U13443 ( .A1(n14563), .A2(n12981), .ZN(n10931) );
  NAND2_X1 U13444 ( .A1(n14562), .A2(n14568), .ZN(n10932) );
  NAND2_X1 U13445 ( .A1(n10933), .A2(n10932), .ZN(n11028) );
  XNOR2_X1 U13446 ( .A(n11028), .B(n11998), .ZN(n10942) );
  INV_X1 U13447 ( .A(n10934), .ZN(n10937) );
  NAND2_X1 U13448 ( .A1(n10935), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U13449 ( .A1(n10937), .A2(n10936), .ZN(n11041) );
  NAND2_X1 U13450 ( .A1(n11154), .A2(n11041), .ZN(n10941) );
  NAND2_X1 U13451 ( .A1(n6530), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U13452 ( .A1(n6531), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U13453 ( .A1(n11216), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n10938) );
  AOI222_X1 U13454 ( .A1(n15068), .A2(n10942), .B1(n12678), .B2(n15065), .C1(
        n12975), .C2(n15062), .ZN(n10949) );
  MUX2_X1 U13455 ( .A(n10943), .B(n10949), .S(n15080), .Z(n10945) );
  AOI22_X1 U13456 ( .A1(n11029), .A2(n15038), .B1(n15075), .B2(n10987), .ZN(
        n10944) );
  OAI211_X1 U13457 ( .C1(n10952), .C2(n12968), .A(n10945), .B(n10944), .ZN(
        P3_U3219) );
  INV_X1 U13458 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n10946) );
  MUX2_X1 U13459 ( .A(n10946), .B(n10949), .S(n15127), .Z(n10948) );
  INV_X1 U13460 ( .A(n13049), .ZN(n13095) );
  NAND2_X1 U13461 ( .A1(n11029), .A2(n13095), .ZN(n10947) );
  OAI211_X1 U13462 ( .C1(n10952), .C2(n13107), .A(n10948), .B(n10947), .ZN(
        P3_U3432) );
  INV_X1 U13463 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12696) );
  MUX2_X1 U13464 ( .A(n12696), .B(n10949), .S(n15142), .Z(n10951) );
  NAND2_X1 U13465 ( .A1(n11029), .A2(n13029), .ZN(n10950) );
  OAI211_X1 U13466 ( .C1(n10952), .C2(n13040), .A(n10951), .B(n10950), .ZN(
        P3_U3473) );
  INV_X1 U13467 ( .A(n11537), .ZN(n11800) );
  OAI222_X1 U13468 ( .A1(P2_U3088), .A2(n10954), .B1(n13766), .B2(n11800), 
        .C1(n10953), .C2(n13749), .ZN(P2_U3303) );
  INV_X1 U13469 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n10957) );
  AOI21_X1 U13470 ( .B1(n10957), .B2(n10956), .A(n12688), .ZN(n10973) );
  AOI21_X1 U13471 ( .B1(n10959), .B2(n10962), .A(n10958), .ZN(n10961) );
  MUX2_X1 U13472 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12777), .Z(n12706) );
  XNOR2_X1 U13473 ( .A(n12706), .B(n12707), .ZN(n10960) );
  NAND2_X1 U13474 ( .A1(n10961), .A2(n10960), .ZN(n12714) );
  OAI21_X1 U13475 ( .B1(n10961), .B2(n10960), .A(n12714), .ZN(n10971) );
  NAND2_X1 U13476 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10962), .ZN(n10964) );
  OAI21_X1 U13477 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n10965), .A(n12694), 
        .ZN(n10966) );
  NAND2_X1 U13478 ( .A1(n10966), .A2(n14990), .ZN(n10969) );
  AOI21_X1 U13479 ( .B1(n14987), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n10967), 
        .ZN(n10968) );
  OAI211_X1 U13480 ( .C1(n14981), .C2(n12693), .A(n10969), .B(n10968), .ZN(
        n10970) );
  AOI21_X1 U13481 ( .B1(n10971), .B2(n12795), .A(n10970), .ZN(n10972) );
  OAI21_X1 U13482 ( .B1(n10973), .B2(n14994), .A(n10972), .ZN(P3_U3195) );
  INV_X1 U13483 ( .A(n11029), .ZN(n10990) );
  XNOR2_X1 U13484 ( .A(n11029), .B(n9489), .ZN(n10975) );
  NOR2_X1 U13485 ( .A1(n10975), .A2(n14564), .ZN(n11003) );
  AOI21_X1 U13486 ( .B1(n10975), .B2(n14564), .A(n11003), .ZN(n10982) );
  NAND2_X1 U13487 ( .A1(n10977), .A2(n10976), .ZN(n10979) );
  NOR2_X1 U13488 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13489 ( .A1(n10981), .A2(n10982), .ZN(n11005) );
  OAI21_X1 U13490 ( .B1(n10982), .B2(n10981), .A(n11005), .ZN(n10983) );
  NAND2_X1 U13491 ( .A1(n10983), .A2(n12651), .ZN(n10989) );
  INV_X1 U13492 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n10984) );
  NOR2_X1 U13493 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10984), .ZN(n12700) );
  AOI21_X1 U13494 ( .B1(n12975), .B2(n12643), .A(n12700), .ZN(n10985) );
  OAI21_X1 U13495 ( .B1(n11033), .B2(n12646), .A(n10985), .ZN(n10986) );
  AOI21_X1 U13496 ( .B1(n10987), .B2(n12670), .A(n10986), .ZN(n10988) );
  OAI211_X1 U13497 ( .C1(n10990), .C2(n12666), .A(n10989), .B(n10988), .ZN(
        P3_U3155) );
  XOR2_X1 U13498 ( .A(n10991), .B(n12285), .Z(n13700) );
  XOR2_X1 U13499 ( .A(n12285), .B(n10992), .Z(n10993) );
  NAND2_X1 U13500 ( .A1(n10993), .A2(n14892), .ZN(n13697) );
  NAND2_X1 U13501 ( .A1(n13253), .A2(n13230), .ZN(n10995) );
  NAND2_X1 U13502 ( .A1(n13255), .A2(n13231), .ZN(n10994) );
  NAND2_X1 U13503 ( .A1(n10995), .A2(n10994), .ZN(n13695) );
  INV_X1 U13504 ( .A(n13695), .ZN(n10996) );
  OAI211_X1 U13505 ( .C1(n13595), .C2(n12387), .A(n13697), .B(n10996), .ZN(
        n10997) );
  NAND2_X1 U13506 ( .A1(n10997), .A2(n13598), .ZN(n11002) );
  AOI211_X1 U13507 ( .C1(n13696), .C2(n10998), .A(n14896), .B(n6673), .ZN(
        n13694) );
  INV_X1 U13508 ( .A(n13696), .ZN(n10999) );
  OAI22_X1 U13509 ( .A1(n10999), .A2(n14879), .B1(n13598), .B2(n15332), .ZN(
        n11000) );
  AOI21_X1 U13510 ( .B1(n13694), .B2(n14874), .A(n11000), .ZN(n11001) );
  OAI211_X1 U13511 ( .C1(n13700), .C2(n13582), .A(n11002), .B(n11001), .ZN(
        P2_U3250) );
  INV_X1 U13512 ( .A(n11003), .ZN(n11004) );
  NAND2_X1 U13513 ( .A1(n11006), .A2(n11971), .ZN(n11008) );
  AOI22_X1 U13514 ( .A1(n11177), .A2(SI_15_), .B1(n11175), .B2(n12742), .ZN(
        n11007) );
  XNOR2_X1 U13515 ( .A(n11049), .B(n9489), .ZN(n11009) );
  NOR2_X1 U13516 ( .A1(n11009), .A2(n12678), .ZN(n11753) );
  INV_X1 U13517 ( .A(n11753), .ZN(n11010) );
  NAND2_X1 U13518 ( .A1(n11009), .A2(n12678), .ZN(n11752) );
  NAND2_X1 U13519 ( .A1(n11010), .A2(n11752), .ZN(n11011) );
  XNOR2_X1 U13520 ( .A(n11754), .B(n11011), .ZN(n11016) );
  NAND2_X1 U13521 ( .A1(n14564), .A2(n12643), .ZN(n11012) );
  NAND2_X1 U13522 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12726)
         );
  OAI211_X1 U13523 ( .C1(n12961), .C2(n12646), .A(n11012), .B(n12726), .ZN(
        n11013) );
  AOI21_X1 U13524 ( .B1(n11041), .B2(n12670), .A(n11013), .ZN(n11015) );
  NAND2_X1 U13525 ( .A1(n11049), .A2(n12648), .ZN(n11014) );
  OAI211_X1 U13526 ( .C1(n11016), .C2(n12672), .A(n11015), .B(n11014), .ZN(
        P3_U3181) );
  OR2_X1 U13527 ( .A1(n11049), .A2(n11033), .ZN(n11907) );
  NAND2_X1 U13528 ( .A1(n11049), .A2(n11033), .ZN(n11906) );
  NAND2_X1 U13529 ( .A1(n11907), .A2(n11906), .ZN(n11903) );
  INV_X1 U13530 ( .A(n11903), .ZN(n11999) );
  NAND2_X1 U13531 ( .A1(n11019), .A2(n11971), .ZN(n11021) );
  INV_X1 U13532 ( .A(n12782), .ZN(n12744) );
  AOI22_X1 U13533 ( .A1(n11177), .A2(SI_16_), .B1(n11175), .B2(n12744), .ZN(
        n11020) );
  OR2_X1 U13534 ( .A1(n13037), .A2(n12961), .ZN(n11910) );
  NAND2_X1 U13535 ( .A1(n13037), .A2(n12961), .ZN(n11911) );
  XNOR2_X1 U13536 ( .A(n11159), .B(n12002), .ZN(n13108) );
  NOR2_X1 U13537 ( .A1(n11022), .A2(n15147), .ZN(n11023) );
  OR2_X1 U13538 ( .A1(n11168), .A2(n11023), .ZN(n12963) );
  NAND2_X1 U13539 ( .A1(n11154), .A2(n12963), .ZN(n11027) );
  NAND2_X1 U13540 ( .A1(n6530), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U13541 ( .A1(n6533), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U13542 ( .A1(n11216), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U13543 ( .A1(n11029), .A2(n14564), .ZN(n11030) );
  NAND2_X1 U13544 ( .A1(n11049), .A2(n12678), .ZN(n11031) );
  XNOR2_X1 U13545 ( .A(n11279), .B(n12002), .ZN(n11032) );
  OAI222_X1 U13546 ( .A1(n15046), .A2(n12656), .B1(n15048), .B2(n11033), .C1(
        n11032), .C2(n15053), .ZN(n13036) );
  NAND2_X1 U13547 ( .A1(n13036), .A2(n15080), .ZN(n11037) );
  INV_X1 U13548 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12751) );
  INV_X1 U13549 ( .A(n12614), .ZN(n11034) );
  OAI22_X1 U13550 ( .A1(n15080), .A2(n12751), .B1(n11034), .B2(n15040), .ZN(
        n11035) );
  AOI21_X1 U13551 ( .B1(n13037), .B2(n15038), .A(n11035), .ZN(n11036) );
  OAI211_X1 U13552 ( .C1(n13108), .C2(n12968), .A(n11037), .B(n11036), .ZN(
        P3_U3217) );
  XNOR2_X1 U13553 ( .A(n11038), .B(n11903), .ZN(n11052) );
  INV_X1 U13554 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12723) );
  XNOR2_X1 U13555 ( .A(n11039), .B(n11999), .ZN(n11040) );
  AOI222_X1 U13556 ( .A1(n15068), .A2(n11040), .B1(n12621), .B2(n15065), .C1(
        n14564), .C2(n15062), .ZN(n11047) );
  MUX2_X1 U13557 ( .A(n12723), .B(n11047), .S(n15080), .Z(n11043) );
  AOI22_X1 U13558 ( .A1(n11049), .A2(n15038), .B1(n15075), .B2(n11041), .ZN(
        n11042) );
  OAI211_X1 U13559 ( .C1(n11052), .C2(n12968), .A(n11043), .B(n11042), .ZN(
        P3_U3218) );
  INV_X1 U13560 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11044) );
  MUX2_X1 U13561 ( .A(n11044), .B(n11047), .S(n15127), .Z(n11046) );
  NAND2_X1 U13562 ( .A1(n11049), .A2(n13095), .ZN(n11045) );
  OAI211_X1 U13563 ( .C1(n11052), .C2(n13107), .A(n11046), .B(n11045), .ZN(
        P3_U3435) );
  INV_X1 U13564 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n11048) );
  MUX2_X1 U13565 ( .A(n11048), .B(n11047), .S(n15142), .Z(n11051) );
  NAND2_X1 U13566 ( .A1(n11049), .A2(n13029), .ZN(n11050) );
  OAI211_X1 U13567 ( .C1(n13040), .C2(n11052), .A(n11051), .B(n11050), .ZN(
        P3_U3474) );
  AOI211_X1 U13568 ( .C1(n14927), .C2(n11055), .A(n11054), .B(n11053), .ZN(
        n11057) );
  MUX2_X1 U13569 ( .A(n15380), .B(n11057), .S(n14972), .Z(n11056) );
  OAI21_X1 U13570 ( .B1(n11060), .B2(n13668), .A(n11056), .ZN(P2_U3513) );
  MUX2_X1 U13571 ( .A(n11058), .B(n11057), .S(n14962), .Z(n11059) );
  OAI21_X1 U13572 ( .B1(n11060), .B2(n13730), .A(n11059), .ZN(P2_U3472) );
  INV_X1 U13573 ( .A(n11559), .ZN(n11064) );
  OAI222_X1 U13574 ( .A1(n13764), .A2(n11062), .B1(n13766), .B2(n11064), .C1(
        P2_U3088), .C2(n11061), .ZN(P2_U3302) );
  OAI222_X1 U13575 ( .A1(n14372), .A2(n15281), .B1(n14370), .B2(n11064), .C1(
        P1_U3086), .C2(n11063), .ZN(P1_U3330) );
  XNOR2_X1 U13576 ( .A(n11076), .B(n11067), .ZN(n13299) );
  OAI21_X1 U13577 ( .B1(n11076), .B2(P2_REG1_REG_12__SCAN_IN), .A(n13297), 
        .ZN(n14861) );
  XNOR2_X1 U13578 ( .A(n14864), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14860) );
  NOR2_X1 U13579 ( .A1(n14861), .A2(n14860), .ZN(n14859) );
  AOI21_X1 U13580 ( .B1(n14864), .B2(P2_REG1_REG_13__SCAN_IN), .A(n14859), 
        .ZN(n13318) );
  XNOR2_X1 U13581 ( .A(n11078), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n13317) );
  NOR2_X1 U13582 ( .A1(n13318), .A2(n13317), .ZN(n13316) );
  NOR2_X1 U13583 ( .A1(n11068), .A2(n11081), .ZN(n11070) );
  XNOR2_X1 U13584 ( .A(n13345), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11071) );
  NOR2_X1 U13585 ( .A1(n11072), .A2(n11071), .ZN(n13344) );
  AOI211_X1 U13586 ( .C1(n11072), .C2(n11071), .A(n13344), .B(n14858), .ZN(
        n11093) );
  INV_X1 U13587 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n11091) );
  MUX2_X1 U13588 ( .A(n11073), .B(P2_REG2_REG_13__SCAN_IN), .S(n11077), .Z(
        n14868) );
  NAND2_X1 U13589 ( .A1(n11075), .A2(n11074), .ZN(n13304) );
  MUX2_X1 U13590 ( .A(n13585), .B(P2_REG2_REG_12__SCAN_IN), .S(n11076), .Z(
        n13305) );
  AOI21_X1 U13591 ( .B1(n13306), .B2(n13304), .A(n13305), .ZN(n13308) );
  AOI21_X1 U13592 ( .B1(n13585), .B2(n13302), .A(n13308), .ZN(n14869) );
  NAND2_X1 U13593 ( .A1(n14868), .A2(n14869), .ZN(n14866) );
  OAI21_X1 U13594 ( .B1(n11073), .B2(n11077), .A(n14866), .ZN(n11079) );
  NAND2_X1 U13595 ( .A1(n11078), .A2(n11079), .ZN(n11080) );
  XNOR2_X1 U13596 ( .A(n13313), .B(n11079), .ZN(n13321) );
  NAND2_X1 U13597 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n13321), .ZN(n13320) );
  NAND2_X1 U13598 ( .A1(n11080), .A2(n13320), .ZN(n11082) );
  NAND2_X1 U13599 ( .A1(n13328), .A2(n11082), .ZN(n11083) );
  XNOR2_X1 U13600 ( .A(n11082), .B(n11081), .ZN(n13326) );
  NAND2_X1 U13601 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13326), .ZN(n13325) );
  NAND2_X1 U13602 ( .A1(n11083), .A2(n13325), .ZN(n11087) );
  NAND2_X1 U13603 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n13345), .ZN(n13338) );
  INV_X1 U13604 ( .A(n13338), .ZN(n11084) );
  AOI21_X1 U13605 ( .B1(n8075), .B2(n11085), .A(n11084), .ZN(n11086) );
  NAND2_X1 U13606 ( .A1(n11086), .A2(n11087), .ZN(n13337) );
  OAI211_X1 U13607 ( .C1(n11087), .C2(n11086), .A(n14867), .B(n13337), .ZN(
        n11090) );
  INV_X1 U13608 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11118) );
  NOR2_X1 U13609 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11118), .ZN(n11088) );
  AOI21_X1 U13610 ( .B1(n14865), .B2(n13345), .A(n11088), .ZN(n11089) );
  OAI211_X1 U13611 ( .C1(n14873), .C2(n11091), .A(n11090), .B(n11089), .ZN(
        n11092) );
  OR2_X1 U13612 ( .A1(n11093), .A2(n11092), .ZN(P2_U3230) );
  NAND2_X1 U13613 ( .A1(n11095), .A2(n11094), .ZN(n11096) );
  NAND2_X1 U13614 ( .A1(n11097), .A2(n11096), .ZN(n13690) );
  INV_X1 U13615 ( .A(n11120), .ZN(n11103) );
  AOI21_X1 U13616 ( .B1(n11098), .B2(n12283), .A(n13509), .ZN(n11100) );
  NAND2_X1 U13617 ( .A1(n11100), .A2(n11099), .ZN(n13688) );
  NAND2_X1 U13618 ( .A1(n13252), .A2(n13230), .ZN(n11102) );
  NAND2_X1 U13619 ( .A1(n13254), .A2(n13231), .ZN(n11101) );
  AND2_X1 U13620 ( .A1(n11102), .A2(n11101), .ZN(n13686) );
  OAI211_X1 U13621 ( .C1(n13595), .C2(n11103), .A(n13688), .B(n13686), .ZN(
        n11106) );
  OAI211_X1 U13622 ( .C1(n6673), .C2(n11123), .A(n13557), .B(n13571), .ZN(
        n13687) );
  AOI22_X1 U13623 ( .A1(n13743), .A2(n13600), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n13561), .ZN(n11104) );
  OAI21_X1 U13624 ( .B1(n13687), .B2(n13578), .A(n11104), .ZN(n11105) );
  AOI21_X1 U13625 ( .B1(n11106), .B2(n13598), .A(n11105), .ZN(n11107) );
  OAI21_X1 U13626 ( .B1(n13582), .B2(n13690), .A(n11107), .ZN(P2_U3249) );
  XNOR2_X1 U13627 ( .A(n13696), .B(n6529), .ZN(n11112) );
  AND2_X1 U13628 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  XNOR2_X1 U13629 ( .A(n13743), .B(n6529), .ZN(n12316) );
  NAND2_X1 U13630 ( .A1(n13253), .A2(n13542), .ZN(n12309) );
  XNOR2_X1 U13631 ( .A(n12316), .B(n12309), .ZN(n11115) );
  OAI21_X1 U13632 ( .B1(n11116), .B2(n11115), .A(n12315), .ZN(n11117) );
  NAND2_X1 U13633 ( .A1(n11117), .A2(n13227), .ZN(n11122) );
  OAI22_X1 U13634 ( .A1(n14811), .A2(n13686), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11118), .ZN(n11119) );
  AOI21_X1 U13635 ( .B1(n11120), .B2(n13223), .A(n11119), .ZN(n11121) );
  OAI211_X1 U13636 ( .C1(n11123), .C2(n13238), .A(n11122), .B(n11121), .ZN(
        P2_U3198) );
  INV_X1 U13637 ( .A(SI_29_), .ZN(n13121) );
  NAND2_X1 U13638 ( .A1(n11126), .A2(n13121), .ZN(n11317) );
  NAND2_X1 U13639 ( .A1(n11321), .A2(n11317), .ZN(n11129) );
  INV_X1 U13640 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11966) );
  INV_X1 U13641 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12374) );
  MUX2_X1 U13642 ( .A(n11966), .B(n12374), .S(n6536), .Z(n11127) );
  INV_X1 U13643 ( .A(SI_30_), .ZN(n12570) );
  NOR2_X1 U13644 ( .A1(n11127), .A2(n12570), .ZN(n11316) );
  INV_X1 U13645 ( .A(n11316), .ZN(n11322) );
  NAND2_X1 U13646 ( .A1(n11127), .A2(n12570), .ZN(n11318) );
  AND2_X1 U13647 ( .A1(n11322), .A2(n11318), .ZN(n11128) );
  INV_X1 U13648 ( .A(n12231), .ZN(n12376) );
  OAI222_X1 U13649 ( .A1(n14370), .A2(n12376), .B1(P1_U3086), .B2(n11130), 
        .C1(n11966), .C2(n14372), .ZN(P1_U3325) );
  INV_X1 U13650 ( .A(n13584), .ZN(n11131) );
  NAND2_X1 U13651 ( .A1(n13223), .A2(n11131), .ZN(n11132) );
  NAND2_X1 U13652 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13301)
         );
  OAI211_X1 U13653 ( .C1(n11133), .C2(n14811), .A(n11132), .B(n13301), .ZN(
        n11139) );
  AOI22_X1 U13654 ( .A1(n11134), .A2(n13227), .B1(n13205), .B2(n13258), .ZN(
        n11136) );
  NOR3_X1 U13655 ( .A1(n11137), .A2(n11136), .A3(n11135), .ZN(n11138) );
  AOI211_X1 U13656 ( .C1(n13587), .C2(n14818), .A(n11139), .B(n11138), .ZN(
        n11140) );
  OAI21_X1 U13657 ( .B1(n11141), .B2(n14813), .A(n11140), .ZN(P2_U3196) );
  INV_X1 U13658 ( .A(n11142), .ZN(n11144) );
  INV_X1 U13659 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U13660 ( .A1(n14371), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U13661 ( .A1(n13765), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11145) );
  AND2_X1 U13662 ( .A1(n13762), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U13663 ( .A1(n14367), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11147) );
  INV_X1 U13664 ( .A(n11273), .ZN(n11149) );
  NAND2_X1 U13665 ( .A1(n11750), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U13666 ( .A1(n11149), .A2(n11148), .ZN(n11151) );
  NAND2_X1 U13667 ( .A1(n13759), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11150) );
  XNOR2_X1 U13668 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11958) );
  XNOR2_X1 U13669 ( .A(n11960), .B(n11958), .ZN(n13117) );
  NAND2_X1 U13670 ( .A1(n13117), .A2(n11971), .ZN(n11153) );
  OR2_X1 U13671 ( .A1(n11274), .A2(n13121), .ZN(n11152) );
  NAND2_X1 U13672 ( .A1(n11154), .A2(n12799), .ZN(n11978) );
  NAND2_X1 U13673 ( .A1(n6530), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n11157) );
  NAND2_X1 U13674 ( .A1(n6533), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U13675 ( .A1(n6944), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n11155) );
  NAND4_X1 U13676 ( .A1(n11978), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(
        n12676) );
  INV_X1 U13677 ( .A(n12002), .ZN(n11158) );
  NAND2_X1 U13678 ( .A1(n11160), .A2(n11971), .ZN(n11162) );
  AOI22_X1 U13679 ( .A1(n11177), .A2(SI_17_), .B1(n11175), .B2(n14529), .ZN(
        n11161) );
  OR2_X1 U13680 ( .A1(n13033), .A2(n12656), .ZN(n11823) );
  NAND2_X1 U13681 ( .A1(n13033), .A2(n12656), .ZN(n11915) );
  NAND2_X1 U13682 ( .A1(n11823), .A2(n11915), .ZN(n12958) );
  NAND2_X1 U13683 ( .A1(n12957), .A2(n6848), .ZN(n11163) );
  OR2_X1 U13684 ( .A1(n11164), .A2(n11198), .ZN(n11166) );
  AOI22_X1 U13685 ( .A1(n11177), .A2(SI_18_), .B1(n11175), .B2(n14542), .ZN(
        n11165) );
  OR2_X1 U13686 ( .A1(n11168), .A2(n11167), .ZN(n11169) );
  NAND2_X1 U13687 ( .A1(n11169), .A2(n11180), .ZN(n12954) );
  NAND2_X1 U13688 ( .A1(n11154), .A2(n12954), .ZN(n11173) );
  NAND2_X1 U13689 ( .A1(n6530), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U13690 ( .A1(n6531), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U13691 ( .A1(n11216), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U13692 ( .A1(n13096), .A2(n12962), .ZN(n11825) );
  NAND2_X1 U13693 ( .A1(n11174), .A2(n11971), .ZN(n11179) );
  AOI22_X1 U13694 ( .A1(n11177), .A2(n11176), .B1(n11175), .B2(n12023), .ZN(
        n11178) );
  AND2_X1 U13695 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n11180), .ZN(n11181) );
  OR2_X1 U13696 ( .A1(n11181), .A2(n11191), .ZN(n12941) );
  NAND2_X1 U13697 ( .A1(n11154), .A2(n12941), .ZN(n11185) );
  NAND2_X1 U13698 ( .A1(n6530), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U13699 ( .A1(n6532), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U13700 ( .A1(n11216), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n11182) );
  NAND4_X1 U13701 ( .A1(n11185), .A2(n11184), .A3(n11183), .A4(n11182), .ZN(
        n12952) );
  NAND2_X1 U13702 ( .A1(n12940), .A2(n12952), .ZN(n11922) );
  AND2_X1 U13703 ( .A1(n11922), .A2(n12928), .ZN(n11822) );
  NAND2_X1 U13704 ( .A1(n11186), .A2(n11971), .ZN(n11189) );
  OR2_X1 U13705 ( .A1(n11274), .A2(n11187), .ZN(n11188) );
  NAND2_X1 U13706 ( .A1(n6530), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n11196) );
  OR2_X1 U13707 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  NAND2_X1 U13708 ( .A1(n11203), .A2(n11192), .ZN(n12923) );
  NAND2_X1 U13709 ( .A1(n11154), .A2(n12923), .ZN(n11195) );
  NAND2_X1 U13710 ( .A1(n6533), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n11194) );
  NAND2_X1 U13711 ( .A1(n11216), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n11193) );
  XNOR2_X1 U13712 ( .A(n13022), .B(n12936), .ZN(n12919) );
  OR2_X1 U13713 ( .A1(n13022), .A2(n12936), .ZN(n11197) );
  OR2_X1 U13714 ( .A1(n11199), .A2(n11198), .ZN(n11202) );
  OR2_X1 U13715 ( .A1(n11274), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U13716 ( .A1(n6530), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U13717 ( .A1(n11203), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U13718 ( .A1(n11214), .A2(n11204), .ZN(n12912) );
  NAND2_X1 U13719 ( .A1(n11154), .A2(n12912), .ZN(n11207) );
  NAND2_X1 U13720 ( .A1(n6531), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U13721 ( .A1(n11216), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n11205) );
  NAND4_X1 U13722 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n12898) );
  NAND2_X1 U13723 ( .A1(n13079), .A2(n12918), .ZN(n11819) );
  NAND2_X1 U13724 ( .A1(n12905), .A2(n11819), .ZN(n11209) );
  OR2_X1 U13725 ( .A1(n13079), .A2(n12918), .ZN(n11818) );
  NAND2_X1 U13726 ( .A1(n11209), .A2(n11818), .ZN(n12895) );
  NAND2_X1 U13727 ( .A1(n11210), .A2(n11971), .ZN(n11213) );
  INV_X1 U13728 ( .A(SI_22_), .ZN(n11211) );
  OR2_X1 U13729 ( .A1(n11274), .A2(n11211), .ZN(n11212) );
  AND2_X1 U13730 ( .A1(n11214), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11215) );
  OR2_X1 U13731 ( .A1(n11215), .A2(n11226), .ZN(n12902) );
  NAND2_X1 U13732 ( .A1(n11154), .A2(n12902), .ZN(n11220) );
  NAND2_X1 U13733 ( .A1(n6530), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U13734 ( .A1(n6532), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U13735 ( .A1(n11216), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n11217) );
  NAND4_X1 U13736 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(
        n12909) );
  NAND2_X1 U13737 ( .A1(n13073), .A2(n12883), .ZN(n11927) );
  NAND2_X1 U13738 ( .A1(n12895), .A2(n11927), .ZN(n12885) );
  NAND2_X1 U13739 ( .A1(n11221), .A2(n11971), .ZN(n11224) );
  OR2_X1 U13740 ( .A1(n11274), .A2(n11222), .ZN(n11223) );
  NAND2_X1 U13741 ( .A1(n6530), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n11231) );
  NOR2_X1 U13742 ( .A1(n11226), .A2(n11225), .ZN(n11227) );
  OR2_X1 U13743 ( .A1(n11237), .A2(n11227), .ZN(n12890) );
  NAND2_X1 U13744 ( .A1(n11154), .A2(n12890), .ZN(n11230) );
  NAND2_X1 U13745 ( .A1(n6533), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U13746 ( .A1(n6944), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n11228) );
  OR2_X1 U13747 ( .A1(n13012), .A2(n12872), .ZN(n11933) );
  AND2_X1 U13748 ( .A1(n12884), .A2(n11933), .ZN(n12862) );
  NAND2_X1 U13749 ( .A1(n11232), .A2(n11971), .ZN(n11235) );
  OR2_X1 U13750 ( .A1(n11274), .A2(n11233), .ZN(n11234) );
  NAND2_X1 U13751 ( .A1(n6530), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n11242) );
  OR2_X1 U13752 ( .A1(n11237), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U13753 ( .A1(n11250), .A2(n11238), .ZN(n12873) );
  NAND2_X1 U13754 ( .A1(n11154), .A2(n12873), .ZN(n11241) );
  NAND2_X1 U13755 ( .A1(n6531), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U13756 ( .A1(n6944), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U13757 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n12854) );
  OR2_X1 U13758 ( .A1(n13008), .A2(n12882), .ZN(n11934) );
  NAND2_X1 U13759 ( .A1(n13008), .A2(n12882), .ZN(n11938) );
  INV_X1 U13760 ( .A(n12868), .ZN(n11243) );
  AND2_X1 U13761 ( .A1(n12862), .A2(n11243), .ZN(n11245) );
  INV_X1 U13762 ( .A(n11933), .ZN(n11244) );
  NAND2_X1 U13763 ( .A1(n12865), .A2(n11938), .ZN(n12849) );
  NAND2_X1 U13764 ( .A1(n11246), .A2(n11971), .ZN(n11249) );
  OR2_X1 U13765 ( .A1(n11274), .A2(n11247), .ZN(n11248) );
  NAND2_X1 U13766 ( .A1(n6530), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U13767 ( .A1(n11250), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n11251) );
  NAND2_X1 U13768 ( .A1(n11261), .A2(n11251), .ZN(n12859) );
  NAND2_X1 U13769 ( .A1(n11154), .A2(n12859), .ZN(n11254) );
  NAND2_X1 U13770 ( .A1(n6532), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U13771 ( .A1(n6944), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n11252) );
  OR2_X1 U13772 ( .A1(n13060), .A2(n12871), .ZN(n11946) );
  NAND2_X1 U13773 ( .A1(n13060), .A2(n12871), .ZN(n11942) );
  INV_X1 U13774 ( .A(n11942), .ZN(n11256) );
  NAND2_X1 U13775 ( .A1(n11257), .A2(n11971), .ZN(n11260) );
  NAND2_X1 U13776 ( .A1(n6530), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n11267) );
  NAND2_X1 U13777 ( .A1(n11261), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U13778 ( .A1(n11263), .A2(n11262), .ZN(n12842) );
  NAND2_X1 U13779 ( .A1(n11154), .A2(n12842), .ZN(n11266) );
  NAND2_X1 U13780 ( .A1(n6533), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U13781 ( .A1(n6944), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n11264) );
  NAND2_X1 U13782 ( .A1(n13000), .A2(n11784), .ZN(n11948) );
  XNOR2_X1 U13783 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n11268) );
  XNOR2_X1 U13784 ( .A(n11269), .B(n11268), .ZN(n12564) );
  NAND2_X1 U13785 ( .A1(n12564), .A2(n11971), .ZN(n11271) );
  OR2_X1 U13786 ( .A1(n11274), .A2(n12565), .ZN(n11270) );
  XNOR2_X1 U13787 ( .A(n13759), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n11272) );
  XNOR2_X1 U13788 ( .A(n11273), .B(n11272), .ZN(n11301) );
  NAND2_X1 U13789 ( .A1(n11301), .A2(n11971), .ZN(n11276) );
  OR2_X1 U13790 ( .A1(n11274), .A2(n11303), .ZN(n11275) );
  NAND2_X1 U13791 ( .A1(n11278), .A2(n12575), .ZN(n11290) );
  INV_X1 U13792 ( .A(n11290), .ZN(n11277) );
  NOR2_X1 U13793 ( .A1(n12579), .A2(n12837), .ZN(n12811) );
  NOR2_X1 U13794 ( .A1(n11277), .A2(n12811), .ZN(n11954) );
  INV_X1 U13795 ( .A(n11291), .ZN(n11953) );
  XOR2_X1 U13796 ( .A(n12009), .B(n12020), .Z(n12383) );
  INV_X1 U13797 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U13798 ( .A1(n11279), .A2(n12002), .ZN(n11281) );
  NAND2_X1 U13799 ( .A1(n13037), .A2(n12621), .ZN(n11280) );
  NAND2_X1 U13800 ( .A1(n11923), .A2(n11922), .ZN(n12932) );
  OR2_X1 U13801 ( .A1(n13096), .A2(n12677), .ZN(n12933) );
  AND2_X1 U13802 ( .A1(n12932), .A2(n12933), .ZN(n11282) );
  INV_X1 U13803 ( .A(n12952), .ZN(n12917) );
  OR2_X1 U13804 ( .A1(n12940), .A2(n12917), .ZN(n11283) );
  NAND2_X1 U13805 ( .A1(n13022), .A2(n12908), .ZN(n11284) );
  AND2_X1 U13806 ( .A1(n13079), .A2(n12898), .ZN(n11815) );
  OR2_X1 U13807 ( .A1(n13079), .A2(n12898), .ZN(n11814) );
  NAND2_X1 U13808 ( .A1(n13012), .A2(n12899), .ZN(n11285) );
  AND2_X1 U13809 ( .A1(n13008), .A2(n12854), .ZN(n11287) );
  OR2_X1 U13810 ( .A1(n13008), .A2(n12854), .ZN(n11288) );
  NOR2_X1 U13811 ( .A1(n13000), .A2(n12855), .ZN(n11289) );
  INV_X1 U13812 ( .A(n12837), .ZN(n11788) );
  NAND2_X1 U13813 ( .A1(n12828), .A2(n15062), .ZN(n11297) );
  NAND2_X1 U13814 ( .A1(n6530), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n11294) );
  NAND2_X1 U13815 ( .A1(n6531), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U13816 ( .A1(n6944), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n11292) );
  NAND4_X1 U13817 ( .A1(n11978), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n12675) );
  AND2_X1 U13818 ( .A1(n12031), .A2(P3_B_REG_SCAN_IN), .ZN(n11295) );
  NOR2_X1 U13819 ( .A1(n15046), .A2(n11295), .ZN(n12800) );
  NAND2_X1 U13820 ( .A1(n12675), .A2(n12800), .ZN(n11296) );
  NAND2_X1 U13821 ( .A1(n12381), .A2(n13029), .ZN(n11300) );
  INV_X1 U13822 ( .A(n11301), .ZN(n11304) );
  OAI222_X1 U13823 ( .A1(n13120), .A2(n11304), .B1(n13122), .B2(n11303), .C1(
        P3_U3151), .C2(n11302), .ZN(P3_U3267) );
  NAND2_X1 U13824 ( .A1(n11305), .A2(n11352), .ZN(n11306) );
  NAND2_X1 U13825 ( .A1(n11307), .A2(n11306), .ZN(n11631) );
  MUX2_X1 U13826 ( .A(n11309), .B(n11308), .S(n11631), .Z(n11348) );
  INV_X1 U13827 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15233) );
  OR2_X1 U13828 ( .A1(n11583), .A2(n15233), .ZN(n11314) );
  INV_X1 U13829 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n11310) );
  OR2_X1 U13830 ( .A1(n11630), .A2(n11310), .ZN(n11313) );
  INV_X1 U13831 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11311) );
  OR2_X1 U13832 ( .A1(n11607), .A2(n11311), .ZN(n11312) );
  AND3_X1 U13833 ( .A1(n11314), .A2(n11313), .A3(n11312), .ZN(n11673) );
  NAND2_X1 U13834 ( .A1(n11636), .A2(n11673), .ZN(n11678) );
  INV_X1 U13835 ( .A(n11678), .ZN(n11336) );
  MUX2_X1 U13836 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6535), .Z(n11315) );
  XNOR2_X1 U13837 ( .A(n11315), .B(SI_31_), .ZN(n11323) );
  NAND2_X1 U13838 ( .A1(n11318), .A2(n11317), .ZN(n11324) );
  INV_X1 U13839 ( .A(n11323), .ZN(n11319) );
  NOR2_X1 U13840 ( .A1(n11324), .A2(n11319), .ZN(n11320) );
  NAND2_X1 U13841 ( .A1(n11321), .A2(n11320), .ZN(n11328) );
  XNOR2_X1 U13842 ( .A(n11323), .B(n11322), .ZN(n11326) );
  NOR2_X1 U13843 ( .A1(n11324), .A2(n11323), .ZN(n11325) );
  OR2_X1 U13844 ( .A1(n11326), .A2(n11325), .ZN(n11327) );
  NAND2_X1 U13845 ( .A1(n13753), .A2(n11622), .ZN(n11330) );
  NAND2_X1 U13846 ( .A1(n11613), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U13847 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  NAND2_X1 U13848 ( .A1(n11334), .A2(n11333), .ZN(n11686) );
  NAND2_X1 U13849 ( .A1(n11686), .A2(n11683), .ZN(n11676) );
  INV_X1 U13850 ( .A(n11673), .ZN(n14031) );
  NAND2_X1 U13851 ( .A1(n11373), .A2(n14031), .ZN(n11675) );
  NOR2_X1 U13852 ( .A1(n14032), .A2(n11675), .ZN(n11335) );
  AOI211_X1 U13853 ( .C1(n11336), .C2(n14032), .A(n11676), .B(n11335), .ZN(
        n11337) );
  AOI22_X1 U13854 ( .A1(n11613), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11455), 
        .B2(n14011), .ZN(n11339) );
  INV_X1 U13855 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11458) );
  INV_X1 U13856 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11341) );
  AND2_X1 U13857 ( .A1(n11461), .A2(n11341), .ZN(n11342) );
  OR2_X1 U13858 ( .A1(n11342), .A2(n11355), .ZN(n14227) );
  INV_X1 U13859 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11345) );
  NAND2_X1 U13860 ( .A1(n11606), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11344) );
  NAND2_X1 U13861 ( .A1(n11582), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11343) );
  OAI211_X1 U13862 ( .C1(n11583), .C2(n11345), .A(n11344), .B(n11343), .ZN(
        n11346) );
  INV_X1 U13863 ( .A(n11346), .ZN(n11347) );
  OAI21_X1 U13864 ( .B1(n14227), .B2(n11608), .A(n11347), .ZN(n13940) );
  INV_X1 U13865 ( .A(n13940), .ZN(n14206) );
  OR3_X1 U13866 ( .A1(n14337), .A2(n14206), .A3(n11636), .ZN(n11350) );
  NAND3_X1 U13867 ( .A1(n14337), .A2(n14206), .A3(n11348), .ZN(n11349) );
  AND2_X1 U13868 ( .A1(n11350), .A2(n11349), .ZN(n11475) );
  NAND2_X1 U13869 ( .A1(n11351), .A2(n11622), .ZN(n11354) );
  AOI22_X1 U13870 ( .A1(n11613), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11352), 
        .B2(n11455), .ZN(n11353) );
  NOR2_X1 U13871 ( .A1(n11355), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11356) );
  NOR2_X1 U13872 ( .A1(n11476), .A2(n11356), .ZN(n14210) );
  NAND2_X1 U13873 ( .A1(n14210), .A2(n11489), .ZN(n11361) );
  INV_X1 U13874 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U13875 ( .A1(n11582), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11358) );
  NAND2_X1 U13876 ( .A1(n11606), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11357) );
  OAI211_X1 U13877 ( .C1(n15222), .C2(n11583), .A(n11358), .B(n11357), .ZN(
        n11359) );
  INV_X1 U13878 ( .A(n11359), .ZN(n11360) );
  OR2_X1 U13879 ( .A1(n14332), .A2(n13905), .ZN(n11473) );
  NAND2_X1 U13880 ( .A1(n14332), .A2(n13905), .ZN(n11698) );
  OAI21_X1 U13881 ( .B1(n11366), .B2(n11365), .A(n11364), .ZN(n11370) );
  INV_X1 U13882 ( .A(n11367), .ZN(n11368) );
  NAND2_X1 U13883 ( .A1(n11371), .A2(n11645), .ZN(n11378) );
  NAND2_X1 U13884 ( .A1(n11348), .A2(n11372), .ZN(n11376) );
  NAND2_X1 U13885 ( .A1(n11373), .A2(n11374), .ZN(n11375) );
  MUX2_X1 U13886 ( .A(n11376), .B(n11375), .S(n13954), .Z(n11377) );
  NAND3_X1 U13887 ( .A1(n11378), .A2(n11646), .A3(n11377), .ZN(n11384) );
  NAND2_X1 U13888 ( .A1(n11348), .A2(n13953), .ZN(n11382) );
  NAND2_X1 U13889 ( .A1(n11379), .A2(n11373), .ZN(n11381) );
  MUX2_X1 U13890 ( .A(n11382), .B(n11381), .S(n11380), .Z(n11383) );
  NAND2_X1 U13891 ( .A1(n11384), .A2(n11383), .ZN(n11389) );
  MUX2_X1 U13892 ( .A(n11386), .B(n11385), .S(n11348), .Z(n11388) );
  MUX2_X1 U13893 ( .A(n7323), .B(n7324), .S(n11373), .Z(n11387) );
  NAND2_X1 U13894 ( .A1(n11389), .A2(n11388), .ZN(n11394) );
  NAND2_X1 U13895 ( .A1(n11396), .A2(n11394), .ZN(n11390) );
  BUF_X1 U13896 ( .A(n11373), .Z(n11423) );
  MUX2_X1 U13897 ( .A(n13952), .B(n14758), .S(n11423), .Z(n11392) );
  MUX2_X1 U13898 ( .A(n13952), .B(n14758), .S(n11348), .Z(n11391) );
  INV_X1 U13899 ( .A(n11392), .ZN(n11393) );
  AND2_X1 U13900 ( .A1(n11394), .A2(n11393), .ZN(n11395) );
  NAND2_X1 U13901 ( .A1(n11396), .A2(n11395), .ZN(n11397) );
  MUX2_X1 U13902 ( .A(n13951), .B(n11398), .S(n11348), .Z(n11401) );
  MUX2_X1 U13903 ( .A(n13951), .B(n11398), .S(n11423), .Z(n11399) );
  INV_X1 U13904 ( .A(n11401), .ZN(n11402) );
  MUX2_X1 U13905 ( .A(n13950), .B(n11403), .S(n11423), .Z(n11406) );
  MUX2_X1 U13906 ( .A(n13950), .B(n11403), .S(n11348), .Z(n11404) );
  NAND2_X1 U13907 ( .A1(n11405), .A2(n11404), .ZN(n11408) );
  MUX2_X1 U13908 ( .A(n13949), .B(n11409), .S(n11348), .Z(n11411) );
  MUX2_X1 U13909 ( .A(n13949), .B(n11409), .S(n11423), .Z(n11410) );
  MUX2_X1 U13910 ( .A(n13948), .B(n11413), .S(n11423), .Z(n11415) );
  MUX2_X1 U13911 ( .A(n13948), .B(n11413), .S(n11348), .Z(n11414) );
  NAND2_X1 U13912 ( .A1(n11417), .A2(n11416), .ZN(n11420) );
  MUX2_X1 U13913 ( .A(n13947), .B(n14790), .S(n11348), .Z(n11421) );
  NAND2_X1 U13914 ( .A1(n11420), .A2(n11421), .ZN(n11419) );
  MUX2_X1 U13915 ( .A(n13947), .B(n14790), .S(n11423), .Z(n11418) );
  INV_X1 U13916 ( .A(n11420), .ZN(n11422) );
  MUX2_X1 U13917 ( .A(n13946), .B(n14672), .S(n11423), .Z(n11425) );
  INV_X1 U13918 ( .A(n11423), .ZN(n11636) );
  MUX2_X1 U13919 ( .A(n13946), .B(n14672), .S(n11636), .Z(n11424) );
  MUX2_X1 U13920 ( .A(n13944), .B(n14666), .S(n11373), .Z(n11440) );
  NAND2_X1 U13921 ( .A1(n14666), .A2(n11636), .ZN(n11426) );
  OAI211_X1 U13922 ( .C1(n14249), .C2(n11636), .A(n11440), .B(n11426), .ZN(
        n11427) );
  MUX2_X1 U13923 ( .A(n12410), .B(n14506), .S(n11636), .Z(n11436) );
  MUX2_X1 U13924 ( .A(n13945), .B(n11428), .S(n11373), .Z(n11435) );
  NAND2_X1 U13925 ( .A1(n11436), .A2(n11435), .ZN(n11429) );
  AOI21_X1 U13926 ( .B1(n11693), .B2(n11430), .A(n11636), .ZN(n11433) );
  AOI21_X1 U13927 ( .B1(n11445), .B2(n11431), .A(n11423), .ZN(n11432) );
  NOR2_X1 U13928 ( .A1(n11433), .A2(n11432), .ZN(n11443) );
  OR3_X1 U13929 ( .A1(n11437), .A2(n11436), .A3(n11435), .ZN(n11442) );
  NAND2_X1 U13930 ( .A1(n14249), .A2(n11373), .ZN(n11438) );
  OAI21_X1 U13931 ( .B1(n14666), .B2(n11373), .A(n11438), .ZN(n11439) );
  OR3_X1 U13932 ( .A1(n10752), .A2(n11440), .A3(n11439), .ZN(n11441) );
  MUX2_X1 U13933 ( .A(n11445), .B(n11693), .S(n11636), .Z(n11446) );
  NAND2_X1 U13934 ( .A1(n11447), .A2(n11622), .ZN(n11450) );
  AOI22_X1 U13935 ( .A1(n11613), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11455), 
        .B2(n11448), .ZN(n11449) );
  MUX2_X1 U13936 ( .A(n13941), .B(n14645), .S(n11373), .Z(n11452) );
  MUX2_X1 U13937 ( .A(n13941), .B(n14645), .S(n11636), .Z(n11451) );
  NAND2_X1 U13938 ( .A1(n11453), .A2(n11622), .ZN(n11457) );
  AOI22_X1 U13939 ( .A1(n11613), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11455), 
        .B2(n11454), .ZN(n11456) );
  NAND2_X1 U13940 ( .A1(n11459), .A2(n11458), .ZN(n11460) );
  AND2_X1 U13941 ( .A1(n11461), .A2(n11460), .ZN(n14238) );
  NAND2_X1 U13942 ( .A1(n14238), .A2(n11489), .ZN(n11466) );
  NAND2_X1 U13943 ( .A1(n6963), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U13944 ( .A1(n11582), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11462) );
  OAI211_X1 U13945 ( .C1(n10831), .C2(n11630), .A(n11463), .B(n11462), .ZN(
        n11464) );
  INV_X1 U13946 ( .A(n11464), .ZN(n11465) );
  NAND2_X1 U13947 ( .A1(n11466), .A2(n11465), .ZN(n14220) );
  NOR2_X1 U13948 ( .A1(n14343), .A2(n14220), .ZN(n11705) );
  NAND2_X1 U13949 ( .A1(n11469), .A2(n11705), .ZN(n11468) );
  INV_X1 U13950 ( .A(n14220), .ZN(n14632) );
  MUX2_X1 U13951 ( .A(n14632), .B(n14240), .S(n11636), .Z(n11467) );
  NAND2_X1 U13952 ( .A1(n11468), .A2(n11467), .ZN(n11472) );
  INV_X1 U13953 ( .A(n11469), .ZN(n11470) );
  AND2_X1 U13954 ( .A1(n14343), .A2(n14220), .ZN(n11663) );
  NAND2_X1 U13955 ( .A1(n11470), .A2(n11663), .ZN(n11471) );
  XNOR2_X1 U13956 ( .A(n14337), .B(n13940), .ZN(n14218) );
  MUX2_X1 U13957 ( .A(n11698), .B(n11473), .S(n11423), .Z(n11474) );
  NOR2_X1 U13958 ( .A1(n11476), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11477) );
  OR2_X1 U13959 ( .A1(n11487), .A2(n11477), .ZN(n13874) );
  INV_X1 U13960 ( .A(n13874), .ZN(n14186) );
  INV_X1 U13961 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U13962 ( .A1(n11582), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U13963 ( .A1(n11606), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11478) );
  OAI211_X1 U13964 ( .C1(n11480), .C2(n11583), .A(n11479), .B(n11478), .ZN(
        n11481) );
  AOI21_X1 U13965 ( .B1(n14186), .B2(n11489), .A(n11481), .ZN(n14205) );
  OR2_X1 U13966 ( .A1(n11482), .A2(n11496), .ZN(n11484) );
  OR2_X1 U13967 ( .A1(n6987), .A2(n15251), .ZN(n11483) );
  MUX2_X1 U13968 ( .A(n14205), .B(n14325), .S(n11423), .Z(n11486) );
  INV_X1 U13969 ( .A(n14205), .ZN(n13939) );
  MUX2_X1 U13970 ( .A(n13939), .B(n13876), .S(n11636), .Z(n11485) );
  OR2_X1 U13971 ( .A1(n11487), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11488) );
  AND2_X1 U13972 ( .A1(n11488), .A2(n11507), .ZN(n14171) );
  NAND2_X1 U13973 ( .A1(n14171), .A2(n11489), .ZN(n11495) );
  INV_X1 U13974 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U13975 ( .A1(n11582), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11491) );
  NAND2_X1 U13976 ( .A1(n11606), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11490) );
  OAI211_X1 U13977 ( .C1(n11492), .C2(n11583), .A(n11491), .B(n11490), .ZN(
        n11493) );
  INV_X1 U13978 ( .A(n11493), .ZN(n11494) );
  NAND2_X1 U13979 ( .A1(n11495), .A2(n11494), .ZN(n14183) );
  OR2_X1 U13980 ( .A1(n6987), .A2(n15252), .ZN(n11498) );
  MUX2_X1 U13981 ( .A(n14183), .B(n14319), .S(n11636), .Z(n11502) );
  MUX2_X1 U13982 ( .A(n14183), .B(n14319), .S(n11423), .Z(n11500) );
  NAND2_X1 U13983 ( .A1(n11501), .A2(n11500), .ZN(n11505) );
  NAND2_X1 U13984 ( .A1(n6963), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11513) );
  INV_X1 U13985 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11506) );
  OR2_X1 U13986 ( .A1(n11607), .A2(n11506), .ZN(n11512) );
  OAI21_X1 U13987 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11508), .A(n11519), 
        .ZN(n14156) );
  OR2_X1 U13988 ( .A1(n11608), .A2(n14156), .ZN(n11511) );
  INV_X1 U13989 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11509) );
  OR2_X1 U13990 ( .A1(n11630), .A2(n11509), .ZN(n11510) );
  NAND4_X1 U13991 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n13938) );
  OR2_X1 U13992 ( .A1(n11514), .A2(n6536), .ZN(n11515) );
  XNOR2_X1 U13993 ( .A(n11515), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14373) );
  MUX2_X1 U13994 ( .A(n13938), .B(n14314), .S(n11373), .Z(n11518) );
  MUX2_X1 U13995 ( .A(n13938), .B(n14314), .S(n11636), .Z(n11517) );
  NAND2_X1 U13996 ( .A1(n11582), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11524) );
  INV_X1 U13997 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15223) );
  OR2_X1 U13998 ( .A1(n11583), .A2(n15223), .ZN(n11523) );
  OAI21_X1 U13999 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11520), .A(n11541), 
        .ZN(n14136) );
  OR2_X1 U14000 ( .A1(n11608), .A2(n14136), .ZN(n11522) );
  OR2_X1 U14001 ( .A1(n11630), .A2(n15417), .ZN(n11521) );
  NAND4_X1 U14002 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n13937) );
  NAND2_X1 U14003 ( .A1(n11525), .A2(n11622), .ZN(n11528) );
  OR2_X1 U14004 ( .A1(n6987), .A2(n11526), .ZN(n11527) );
  MUX2_X1 U14005 ( .A(n13937), .B(n14307), .S(n11636), .Z(n11532) );
  NAND2_X1 U14006 ( .A1(n11531), .A2(n11532), .ZN(n11530) );
  MUX2_X1 U14007 ( .A(n13937), .B(n14307), .S(n11423), .Z(n11529) );
  NAND2_X1 U14008 ( .A1(n11530), .A2(n11529), .ZN(n11536) );
  INV_X1 U14009 ( .A(n11531), .ZN(n11534) );
  INV_X1 U14010 ( .A(n11532), .ZN(n11533) );
  NAND2_X1 U14011 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  NAND2_X1 U14012 ( .A1(n11536), .A2(n11535), .ZN(n11550) );
  NAND2_X1 U14013 ( .A1(n11537), .A2(n11622), .ZN(n11539) );
  NAND2_X1 U14014 ( .A1(n11613), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11538) );
  NAND2_X1 U14015 ( .A1(n11564), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11548) );
  INV_X1 U14016 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11540) );
  OR2_X1 U14017 ( .A1(n11583), .A2(n11540), .ZN(n11547) );
  INV_X1 U14018 ( .A(n11541), .ZN(n11543) );
  INV_X1 U14019 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15270) );
  INV_X1 U14020 ( .A(n11553), .ZN(n11542) );
  OAI21_X1 U14021 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11543), .A(n11542), 
        .ZN(n13866) );
  OR2_X1 U14022 ( .A1(n11608), .A2(n13866), .ZN(n11546) );
  INV_X1 U14023 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n11544) );
  OR2_X1 U14024 ( .A1(n11630), .A2(n11544), .ZN(n11545) );
  NAND4_X1 U14025 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n13936) );
  MUX2_X1 U14026 ( .A(n14301), .B(n13936), .S(n11636), .Z(n11551) );
  MUX2_X1 U14027 ( .A(n13936), .B(n14301), .S(n11636), .Z(n11549) );
  NAND2_X1 U14028 ( .A1(n11582), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11558) );
  INV_X1 U14029 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11552) );
  OR2_X1 U14030 ( .A1(n11583), .A2(n11552), .ZN(n11557) );
  NAND2_X1 U14031 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11553), .ZN(n11566) );
  OAI21_X1 U14032 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11553), .A(n11566), 
        .ZN(n14111) );
  OR2_X1 U14033 ( .A1(n11608), .A2(n14111), .ZN(n11556) );
  INV_X1 U14034 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11554) );
  OR2_X1 U14035 ( .A1(n11630), .A2(n11554), .ZN(n11555) );
  NAND4_X1 U14036 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n13935) );
  NAND2_X1 U14037 ( .A1(n11559), .A2(n11622), .ZN(n11561) );
  OR2_X1 U14038 ( .A1(n6987), .A2(n15281), .ZN(n11560) );
  MUX2_X1 U14039 ( .A(n13935), .B(n14293), .S(n11636), .Z(n11563) );
  MUX2_X1 U14040 ( .A(n14293), .B(n13935), .S(n11636), .Z(n11562) );
  NAND2_X1 U14041 ( .A1(n11564), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11571) );
  INV_X1 U14042 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15329) );
  OR2_X1 U14043 ( .A1(n11583), .A2(n15329), .ZN(n11570) );
  INV_X1 U14044 ( .A(n11566), .ZN(n11565) );
  INV_X1 U14045 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13914) );
  NAND2_X1 U14046 ( .A1(n11566), .A2(n13914), .ZN(n11567) );
  NAND2_X1 U14047 ( .A1(n11592), .A2(n11567), .ZN(n14093) );
  OR2_X1 U14048 ( .A1(n11608), .A2(n14093), .ZN(n11569) );
  INV_X1 U14049 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14096) );
  OR2_X1 U14050 ( .A1(n11630), .A2(n14096), .ZN(n11568) );
  NAND4_X1 U14051 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n13934) );
  NAND2_X1 U14052 ( .A1(n13763), .A2(n11622), .ZN(n11573) );
  OR2_X1 U14053 ( .A1(n6987), .A2(n14371), .ZN(n11572) );
  NAND2_X2 U14054 ( .A1(n11573), .A2(n11572), .ZN(n14289) );
  MUX2_X1 U14055 ( .A(n13934), .B(n14289), .S(n11423), .Z(n11577) );
  NAND2_X1 U14056 ( .A1(n11576), .A2(n11577), .ZN(n11575) );
  MUX2_X1 U14057 ( .A(n14289), .B(n13934), .S(n11423), .Z(n11574) );
  INV_X1 U14058 ( .A(n11576), .ZN(n11579) );
  INV_X1 U14059 ( .A(n11577), .ZN(n11578) );
  NAND2_X1 U14060 ( .A1(n13760), .A2(n11622), .ZN(n11581) );
  OR2_X1 U14061 ( .A1(n6987), .A2(n14367), .ZN(n11580) );
  NAND2_X1 U14062 ( .A1(n11582), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11588) );
  INV_X1 U14063 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15185) );
  OR2_X1 U14064 ( .A1(n11583), .A2(n15185), .ZN(n11587) );
  INV_X1 U14065 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13773) );
  XNOR2_X1 U14066 ( .A(n11592), .B(n13773), .ZN(n13772) );
  OR2_X1 U14067 ( .A1(n11608), .A2(n13772), .ZN(n11586) );
  INV_X1 U14068 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11584) );
  OR2_X1 U14069 ( .A1(n11630), .A2(n11584), .ZN(n11585) );
  MUX2_X1 U14070 ( .A(n14055), .B(n14042), .S(n11636), .Z(n11590) );
  MUX2_X1 U14071 ( .A(n14055), .B(n14042), .S(n11373), .Z(n11589) );
  NAND2_X1 U14072 ( .A1(n6963), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11600) );
  INV_X1 U14073 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15292) );
  OR2_X1 U14074 ( .A1(n11607), .A2(n15292), .ZN(n11599) );
  INV_X1 U14075 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11591) );
  OAI21_X1 U14076 ( .B1(n11592), .B2(n13773), .A(n11591), .ZN(n11595) );
  INV_X1 U14077 ( .A(n11592), .ZN(n11594) );
  AND2_X1 U14078 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n11593) );
  NAND2_X1 U14079 ( .A1(n11594), .A2(n11593), .ZN(n14049) );
  NAND2_X1 U14080 ( .A1(n11595), .A2(n14049), .ZN(n14078) );
  OR2_X1 U14081 ( .A1(n11608), .A2(n14078), .ZN(n11598) );
  INV_X1 U14082 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11596) );
  OR2_X1 U14083 ( .A1(n11630), .A2(n11596), .ZN(n11597) );
  NAND4_X1 U14084 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n14058) );
  NAND2_X1 U14085 ( .A1(n13756), .A2(n11622), .ZN(n11602) );
  OR2_X1 U14086 ( .A1(n6987), .A2(n11750), .ZN(n11601) );
  MUX2_X1 U14087 ( .A(n14058), .B(n14280), .S(n11423), .Z(n11604) );
  MUX2_X1 U14088 ( .A(n14058), .B(n14280), .S(n11636), .Z(n11603) );
  NAND2_X1 U14089 ( .A1(n6963), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11612) );
  NAND2_X1 U14090 ( .A1(n11606), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11611) );
  INV_X1 U14091 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15149) );
  OR2_X1 U14092 ( .A1(n11607), .A2(n15149), .ZN(n11610) );
  OR2_X1 U14093 ( .A1(n11608), .A2(n14049), .ZN(n11609) );
  NAND4_X1 U14094 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n14069) );
  NAND2_X1 U14095 ( .A1(n12371), .A2(n11622), .ZN(n11615) );
  NAND2_X1 U14096 ( .A1(n11613), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11614) );
  MUX2_X1 U14097 ( .A(n14069), .B(n14273), .S(n11636), .Z(n11617) );
  MUX2_X1 U14098 ( .A(n14273), .B(n14069), .S(n11348), .Z(n11620) );
  INV_X1 U14099 ( .A(n11616), .ZN(n11619) );
  INV_X1 U14100 ( .A(n11617), .ZN(n11618) );
  NAND2_X1 U14101 ( .A1(n12231), .A2(n11622), .ZN(n11625) );
  OR2_X1 U14102 ( .A1(n6987), .A2(n11966), .ZN(n11624) );
  INV_X1 U14103 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U14104 ( .A1(n6963), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14105 ( .A1(n11582), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11627) );
  OAI211_X1 U14106 ( .C1(n11630), .C2(n11629), .A(n11628), .B(n11627), .ZN(
        n14047) );
  INV_X1 U14107 ( .A(n11631), .ZN(n11632) );
  OAI22_X1 U14108 ( .A1(n11373), .A2(n11673), .B1(n11633), .B2(n11632), .ZN(
        n11634) );
  AOI22_X1 U14109 ( .A1(n14039), .A2(n11373), .B1(n14047), .B2(n11634), .ZN(
        n11638) );
  OAI21_X1 U14110 ( .B1(n14031), .B2(n11635), .A(n14047), .ZN(n11637) );
  MUX2_X1 U14111 ( .A(n11637), .B(n14270), .S(n11636), .Z(n11639) );
  XOR2_X1 U14112 ( .A(n14031), .B(n14032), .Z(n11687) );
  NAND2_X1 U14113 ( .A1(n14280), .A2(n14058), .ZN(n14043) );
  OR2_X1 U14114 ( .A1(n14280), .A2(n14058), .ZN(n11640) );
  XNOR2_X1 U14115 ( .A(n14289), .B(n13934), .ZN(n14088) );
  INV_X1 U14116 ( .A(n13937), .ZN(n13889) );
  XNOR2_X1 U14117 ( .A(n14307), .B(n13889), .ZN(n14137) );
  INV_X1 U14118 ( .A(n14314), .ZN(n11641) );
  NAND2_X1 U14119 ( .A1(n11641), .A2(n13938), .ZN(n11642) );
  NAND2_X1 U14120 ( .A1(n11700), .A2(n11642), .ZN(n14150) );
  INV_X1 U14121 ( .A(n14183), .ZN(n13890) );
  XNOR2_X1 U14122 ( .A(n14319), .B(n13890), .ZN(n14164) );
  XNOR2_X1 U14123 ( .A(n13876), .B(n13939), .ZN(n14181) );
  INV_X1 U14124 ( .A(n13941), .ZN(n13924) );
  NAND2_X1 U14125 ( .A1(n14645), .A2(n13924), .ZN(n11696) );
  OR2_X1 U14126 ( .A1(n14645), .A2(n13924), .ZN(n11643) );
  NAND2_X1 U14127 ( .A1(n11696), .A2(n11643), .ZN(n14627) );
  NAND4_X1 U14128 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n6896), .ZN(
        n11648) );
  NOR3_X1 U14129 ( .A1(n11650), .A2(n11649), .A3(n11648), .ZN(n11653) );
  NAND4_X1 U14130 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  NOR2_X1 U14131 ( .A1(n11656), .A2(n11655), .ZN(n11659) );
  NAND4_X1 U14132 ( .A1(n14485), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11660) );
  OR4_X1 U14133 ( .A1(n14627), .A2(n10752), .A3(n11661), .A4(n11660), .ZN(
        n11662) );
  NOR2_X1 U14134 ( .A1(n11694), .A2(n11662), .ZN(n11665) );
  INV_X1 U14135 ( .A(n11705), .ZN(n11664) );
  INV_X1 U14136 ( .A(n11663), .ZN(n11706) );
  NAND2_X1 U14137 ( .A1(n11664), .A2(n11706), .ZN(n14241) );
  NAND4_X1 U14138 ( .A1(n14181), .A2(n11665), .A3(n14218), .A4(n14241), .ZN(
        n11666) );
  OR4_X1 U14139 ( .A1(n14150), .A2(n14164), .A3(n14203), .A4(n11666), .ZN(
        n11667) );
  NOR2_X1 U14140 ( .A1(n14137), .A2(n11667), .ZN(n11668) );
  XNOR2_X1 U14141 ( .A(n14293), .B(n13935), .ZN(n14102) );
  XNOR2_X1 U14142 ( .A(n14301), .B(n13936), .ZN(n14125) );
  NAND4_X1 U14143 ( .A1(n14088), .A2(n11668), .A3(n14102), .A4(n14125), .ZN(
        n11669) );
  NOR4_X1 U14144 ( .A1(n11687), .A2(n14056), .A3(n14075), .A4(n11669), .ZN(
        n11671) );
  XNOR2_X1 U14145 ( .A(n14039), .B(n14047), .ZN(n11670) );
  XNOR2_X1 U14146 ( .A(n14273), .B(n14069), .ZN(n14060) );
  NAND3_X1 U14147 ( .A1(n11671), .A2(n11670), .A3(n14060), .ZN(n11672) );
  XNOR2_X1 U14148 ( .A(n11672), .B(n14635), .ZN(n11684) );
  INV_X1 U14149 ( .A(n11686), .ZN(n11679) );
  OAI21_X1 U14150 ( .B1(n11673), .B2(n11676), .A(n11675), .ZN(n11674) );
  OAI21_X1 U14151 ( .B1(n11679), .B2(n11675), .A(n11674), .ZN(n11681) );
  OAI21_X1 U14152 ( .B1(n14031), .B2(n11676), .A(n11678), .ZN(n11677) );
  OAI21_X1 U14153 ( .B1(n11679), .B2(n11678), .A(n11677), .ZN(n11680) );
  MUX2_X1 U14154 ( .A(n11681), .B(n11680), .S(n14032), .Z(n11682) );
  OAI21_X1 U14155 ( .B1(n11684), .B2(n11683), .A(n11682), .ZN(n11685) );
  NAND3_X1 U14156 ( .A1(n11689), .A2(n11688), .A3(n14221), .ZN(n11690) );
  OAI211_X1 U14157 ( .C1(n14374), .C2(n11692), .A(n11690), .B(P1_B_REG_SCAN_IN), .ZN(n11691) );
  INV_X1 U14158 ( .A(n14293), .ZN(n14107) );
  INV_X1 U14159 ( .A(n14301), .ZN(n14132) );
  NAND2_X1 U14160 ( .A1(n14240), .A2(n14220), .ZN(n11697) );
  AOI22_X1 U14161 ( .A1(n14242), .A2(n11697), .B1(n14632), .B2(n14343), .ZN(
        n14219) );
  NAND2_X1 U14162 ( .A1(n14219), .A2(n14218), .ZN(n14217) );
  OAI21_X1 U14163 ( .B1(n14206), .B2(n14337), .A(n14217), .ZN(n14202) );
  INV_X1 U14164 ( .A(n11698), .ZN(n11699) );
  NAND2_X1 U14165 ( .A1(n14325), .A2(n13939), .ZN(n14163) );
  NOR2_X1 U14166 ( .A1(n14319), .A2(n13890), .ZN(n14151) );
  INV_X1 U14167 ( .A(n13934), .ZN(n13828) );
  XNOR2_X1 U14168 ( .A(n14057), .B(n14056), .ZN(n11720) );
  INV_X1 U14169 ( .A(n14289), .ZN(n14097) );
  OR2_X1 U14170 ( .A1(n13930), .A2(n13942), .ZN(n11701) );
  NAND2_X1 U14171 ( .A1(n11702), .A2(n11701), .ZN(n14621) );
  NAND2_X1 U14172 ( .A1(n14621), .A2(n14627), .ZN(n11704) );
  OR2_X1 U14173 ( .A1(n14645), .A2(n13941), .ZN(n11703) );
  AND2_X1 U14174 ( .A1(n14337), .A2(n13940), .ZN(n11707) );
  INV_X1 U14175 ( .A(n13905), .ZN(n14223) );
  NOR2_X1 U14176 ( .A1(n14332), .A2(n14223), .ZN(n11708) );
  INV_X1 U14177 ( .A(n14181), .ZN(n14190) );
  OR2_X1 U14178 ( .A1(n14325), .A2(n14205), .ZN(n11709) );
  OR2_X1 U14179 ( .A1(n14319), .A2(n14183), .ZN(n11710) );
  NAND2_X1 U14180 ( .A1(n14149), .A2(n14150), .ZN(n11712) );
  OR2_X1 U14181 ( .A1(n14314), .A2(n13938), .ZN(n11711) );
  INV_X1 U14182 ( .A(n14137), .ZN(n14144) );
  NAND2_X1 U14183 ( .A1(n14307), .A2(n13937), .ZN(n11713) );
  OR2_X1 U14184 ( .A1(n14301), .A2(n13936), .ZN(n11715) );
  INV_X1 U14185 ( .A(n14102), .ZN(n14108) );
  NAND2_X1 U14186 ( .A1(n14293), .A2(n13935), .ZN(n11716) );
  NAND2_X1 U14187 ( .A1(n7419), .A2(n14087), .ZN(n14086) );
  AOI22_X1 U14188 ( .A1(n14222), .A2(n14058), .B1(n13934), .B2(n14221), .ZN(
        n11718) );
  OAI21_X1 U14189 ( .B1(n6582), .B2(n14496), .A(n11718), .ZN(n11719) );
  OR2_X2 U14190 ( .A1(n14188), .A2(n14319), .ZN(n14169) );
  INV_X1 U14191 ( .A(n14095), .ZN(n11722) );
  NAND2_X1 U14192 ( .A1(n14055), .A2(n14095), .ZN(n14080) );
  INV_X1 U14193 ( .A(n14080), .ZN(n11721) );
  AOI21_X1 U14194 ( .B1(n14284), .B2(n11722), .A(n11721), .ZN(n14285) );
  INV_X1 U14195 ( .A(n13772), .ZN(n11723) );
  AOI22_X1 U14196 ( .A1(n14747), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n11723), 
        .B2(n14735), .ZN(n11724) );
  OAI21_X1 U14197 ( .B1(n14055), .B2(n14738), .A(n11724), .ZN(n11726) );
  NOR2_X1 U14198 ( .A1(n6582), .A2(n14739), .ZN(n11725) );
  AOI211_X1 U14199 ( .C1(n14285), .C2(n14195), .A(n11726), .B(n11725), .ZN(
        n11727) );
  OAI21_X1 U14200 ( .B1(n14287), .B2(n14747), .A(n11727), .ZN(P1_U3266) );
  NAND2_X1 U14201 ( .A1(n11729), .A2(P3_D_REG_0__SCAN_IN), .ZN(n11728) );
  OAI21_X1 U14202 ( .B1(n11730), .B2(n11729), .A(n11728), .ZN(P3_U3376) );
  NAND3_X1 U14203 ( .A1(n7313), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n11735) );
  NAND2_X1 U14204 ( .A1(n13753), .A2(n11731), .ZN(n11734) );
  NAND2_X1 U14205 ( .A1(n11732), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11733) );
  OAI211_X1 U14206 ( .C1(n11736), .C2(n11735), .A(n11734), .B(n11733), .ZN(
        P1_U3324) );
  NAND2_X1 U14207 ( .A1(n13267), .A2(n13231), .ZN(n11738) );
  NAND2_X1 U14208 ( .A1(n13265), .A2(n13230), .ZN(n11737) );
  AND2_X1 U14209 ( .A1(n11738), .A2(n11737), .ZN(n14894) );
  OAI22_X1 U14210 ( .A1(n14811), .A2(n14894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14903), .ZN(n11740) );
  NOR2_X1 U14211 ( .A1(n13238), .A2(n14930), .ZN(n11739) );
  AOI211_X1 U14212 ( .C1(n14903), .C2(n13223), .A(n11740), .B(n11739), .ZN(
        n11747) );
  AND2_X1 U14213 ( .A1(n11742), .A2(n11741), .ZN(n11745) );
  OAI211_X1 U14214 ( .C1(n11745), .C2(n11744), .A(n11743), .B(n13227), .ZN(
        n11746) );
  NAND2_X1 U14215 ( .A1(n11747), .A2(n11746), .ZN(P2_U3190) );
  INV_X1 U14216 ( .A(n13756), .ZN(n11749) );
  OAI222_X1 U14217 ( .A1(n11751), .A2(n11750), .B1(n14370), .B2(n11749), .C1(
        n11748), .C2(P1_U3086), .ZN(P1_U3327) );
  XNOR2_X1 U14218 ( .A(n13037), .B(n11786), .ZN(n11755) );
  XNOR2_X1 U14219 ( .A(n11755), .B(n12621), .ZN(n12610) );
  XNOR2_X1 U14220 ( .A(n13033), .B(n11786), .ZN(n11756) );
  XNOR2_X1 U14221 ( .A(n11756), .B(n12951), .ZN(n12619) );
  INV_X1 U14222 ( .A(n11756), .ZN(n11757) );
  NAND2_X1 U14223 ( .A1(n11757), .A2(n12951), .ZN(n11758) );
  NAND2_X1 U14224 ( .A1(n12618), .A2(n11758), .ZN(n12654) );
  XNOR2_X1 U14225 ( .A(n13096), .B(n11786), .ZN(n11759) );
  XNOR2_X1 U14226 ( .A(n11759), .B(n12677), .ZN(n12653) );
  NAND2_X1 U14227 ( .A1(n12654), .A2(n12653), .ZN(n12652) );
  INV_X1 U14228 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14229 ( .A1(n11760), .A2(n12677), .ZN(n11761) );
  NAND2_X1 U14230 ( .A1(n12652), .A2(n11761), .ZN(n12588) );
  XNOR2_X1 U14231 ( .A(n12940), .B(n11786), .ZN(n11762) );
  XNOR2_X1 U14232 ( .A(n11762), .B(n12917), .ZN(n12587) );
  NAND2_X1 U14233 ( .A1(n12588), .A2(n12587), .ZN(n12586) );
  NAND2_X1 U14234 ( .A1(n11762), .A2(n12952), .ZN(n11763) );
  NAND2_X1 U14235 ( .A1(n12586), .A2(n11763), .ZN(n12636) );
  XNOR2_X1 U14236 ( .A(n13022), .B(n11786), .ZN(n11764) );
  XNOR2_X1 U14237 ( .A(n11764), .B(n12908), .ZN(n12635) );
  INV_X1 U14238 ( .A(n11764), .ZN(n11765) );
  NAND2_X1 U14239 ( .A1(n11765), .A2(n12908), .ZN(n11766) );
  XNOR2_X1 U14240 ( .A(n13079), .B(n11786), .ZN(n11768) );
  XNOR2_X1 U14241 ( .A(n11768), .B(n12918), .ZN(n12596) );
  INV_X1 U14242 ( .A(n12596), .ZN(n11767) );
  NAND2_X1 U14243 ( .A1(n11768), .A2(n12918), .ZN(n11769) );
  NAND2_X1 U14244 ( .A1(n12593), .A2(n11769), .ZN(n11773) );
  XNOR2_X1 U14245 ( .A(n13073), .B(n9489), .ZN(n11771) );
  INV_X1 U14246 ( .A(n11771), .ZN(n11772) );
  AOI22_X1 U14247 ( .A1(n12642), .A2(n12883), .B1(n11773), .B2(n11772), .ZN(
        n11776) );
  XNOR2_X1 U14248 ( .A(n13012), .B(n11786), .ZN(n11774) );
  XNOR2_X1 U14249 ( .A(n11776), .B(n11774), .ZN(n12580) );
  NAND2_X1 U14250 ( .A1(n12580), .A2(n12872), .ZN(n11778) );
  INV_X1 U14251 ( .A(n11774), .ZN(n11775) );
  OR2_X1 U14252 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  NAND2_X1 U14253 ( .A1(n11778), .A2(n11777), .ZN(n12627) );
  XNOR2_X1 U14254 ( .A(n13008), .B(n11786), .ZN(n11779) );
  XNOR2_X1 U14255 ( .A(n11779), .B(n12854), .ZN(n12628) );
  NAND2_X1 U14256 ( .A1(n11779), .A2(n12882), .ZN(n11780) );
  XNOR2_X1 U14257 ( .A(n13060), .B(n11786), .ZN(n11781) );
  XNOR2_X1 U14258 ( .A(n11781), .B(n12838), .ZN(n12603) );
  NAND2_X1 U14259 ( .A1(n11781), .A2(n12871), .ZN(n11782) );
  XNOR2_X1 U14260 ( .A(n13000), .B(n11786), .ZN(n11785) );
  XNOR2_X1 U14261 ( .A(n11785), .B(n12855), .ZN(n12662) );
  XNOR2_X1 U14262 ( .A(n13053), .B(n11786), .ZN(n11787) );
  XNOR2_X1 U14263 ( .A(n11787), .B(n12837), .ZN(n12571) );
  XOR2_X1 U14264 ( .A(n11786), .B(n12812), .Z(n11790) );
  XNOR2_X1 U14265 ( .A(n11791), .B(n11790), .ZN(n11796) );
  INV_X1 U14266 ( .A(n12676), .ZN(n12809) );
  AOI22_X1 U14267 ( .A1(n12837), .A2(n12643), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11792) );
  OAI21_X1 U14268 ( .B1(n12809), .B2(n12646), .A(n11792), .ZN(n11794) );
  NOR2_X1 U14269 ( .A1(n13050), .A2(n12666), .ZN(n11793) );
  AOI211_X1 U14270 ( .C1(n12814), .C2(n12670), .A(n11794), .B(n11793), .ZN(
        n11795) );
  OAI21_X1 U14271 ( .B1(n11796), .B2(n12672), .A(n11795), .ZN(P3_U3160) );
  INV_X1 U14272 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14273 ( .A1(n14749), .A2(n11798), .B1(n11797), .B2(n11799), .ZN(
        P1_U3445) );
  OAI222_X1 U14274 ( .A1(n14372), .A2(n11801), .B1(n14370), .B2(n11800), .C1(
        n11799), .C2(P1_U3086), .ZN(P1_U3331) );
  NOR2_X1 U14275 ( .A1(n11802), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13289) );
  AOI21_X1 U14276 ( .B1(n13235), .B2(n11803), .A(n13289), .ZN(n11804) );
  OAI21_X1 U14277 ( .B1(n11805), .B2(n14821), .A(n11804), .ZN(n11811) );
  INV_X1 U14278 ( .A(n10376), .ZN(n11809) );
  AOI22_X1 U14279 ( .A1(n11806), .A2(n13227), .B1(n13205), .B2(n13261), .ZN(
        n11808) );
  NOR3_X1 U14280 ( .A1(n11809), .A2(n11808), .A3(n11807), .ZN(n11810) );
  AOI211_X1 U14281 ( .C1(n12103), .C2(n14818), .A(n11811), .B(n11810), .ZN(
        n11812) );
  OAI21_X1 U14282 ( .B1(n6989), .B2(n14813), .A(n11812), .ZN(P2_U3203) );
  NAND2_X1 U14283 ( .A1(n12884), .A2(n11927), .ZN(n12896) );
  INV_X1 U14284 ( .A(n11814), .ZN(n11816) );
  MUX2_X1 U14285 ( .A(n11955), .B(n12908), .S(n13022), .Z(n11817) );
  AOI21_X1 U14286 ( .B1(n12936), .B2(n11936), .A(n11817), .ZN(n11821) );
  MUX2_X1 U14287 ( .A(n11819), .B(n11818), .S(n11955), .Z(n11820) );
  OAI21_X1 U14288 ( .B1(n12907), .B2(n11821), .A(n11820), .ZN(n11930) );
  INV_X1 U14289 ( .A(n11825), .ZN(n11824) );
  OAI211_X1 U14290 ( .C1(n11824), .C2(n11823), .A(n11822), .B(n11955), .ZN(
        n11921) );
  NAND3_X1 U14291 ( .A1(n11923), .A2(n11936), .A3(n11825), .ZN(n11920) );
  INV_X1 U14292 ( .A(n15067), .ZN(n11986) );
  NAND3_X1 U14293 ( .A1(n11986), .A2(n12034), .A3(n11826), .ZN(n11830) );
  OAI211_X1 U14294 ( .C1(n11827), .C2(n11828), .A(n11936), .B(n11832), .ZN(
        n11829) );
  AOI22_X1 U14295 ( .A1(n11830), .A2(n11829), .B1(n15061), .B2(n11828), .ZN(
        n11836) );
  INV_X1 U14296 ( .A(n11831), .ZN(n11834) );
  INV_X1 U14297 ( .A(n11832), .ZN(n11833) );
  MUX2_X1 U14298 ( .A(n11834), .B(n11833), .S(n11955), .Z(n11835) );
  NOR3_X1 U14299 ( .A1(n11836), .A2(n11835), .A3(n11994), .ZN(n11845) );
  NAND2_X1 U14300 ( .A1(n15064), .A2(n9876), .ZN(n11837) );
  NAND2_X1 U14301 ( .A1(n11842), .A2(n11837), .ZN(n11840) );
  NAND2_X1 U14302 ( .A1(n11841), .A2(n11838), .ZN(n11839) );
  MUX2_X1 U14303 ( .A(n11840), .B(n11839), .S(n11936), .Z(n11844) );
  MUX2_X1 U14304 ( .A(n11842), .B(n11841), .S(n11955), .Z(n11843) );
  OAI21_X1 U14305 ( .B1(n11845), .B2(n11844), .A(n11843), .ZN(n11849) );
  NOR3_X1 U14306 ( .A1(n11847), .A2(n11846), .A3(n11955), .ZN(n11848) );
  AOI21_X1 U14307 ( .B1(n11849), .B2(n11990), .A(n11848), .ZN(n11856) );
  INV_X1 U14308 ( .A(n11850), .ZN(n11854) );
  INV_X1 U14309 ( .A(n11851), .ZN(n11853) );
  INV_X1 U14310 ( .A(n11861), .ZN(n11852) );
  AOI211_X1 U14311 ( .C1(n11989), .C2(n11854), .A(n11853), .B(n11852), .ZN(
        n11855) );
  OAI22_X1 U14312 ( .A1(n11856), .A2(n7206), .B1(n11855), .B2(n11936), .ZN(
        n11860) );
  AOI21_X1 U14313 ( .B1(n11859), .B2(n11857), .A(n11955), .ZN(n11858) );
  AOI21_X1 U14314 ( .B1(n11860), .B2(n11859), .A(n11858), .ZN(n11866) );
  OAI21_X1 U14315 ( .B1(n11955), .B2(n11861), .A(n11991), .ZN(n11865) );
  MUX2_X1 U14316 ( .A(n11863), .B(n11862), .S(n11955), .Z(n11864) );
  OAI211_X1 U14317 ( .C1(n11866), .C2(n11865), .A(n11988), .B(n11864), .ZN(
        n11870) );
  INV_X1 U14318 ( .A(n15015), .ZN(n15017) );
  MUX2_X1 U14319 ( .A(n11868), .B(n11867), .S(n11936), .Z(n11869) );
  NAND3_X1 U14320 ( .A1(n11870), .A2(n15017), .A3(n11869), .ZN(n11876) );
  NAND2_X1 U14321 ( .A1(n15001), .A2(n11936), .ZN(n11874) );
  NAND2_X1 U14322 ( .A1(n11871), .A2(n11955), .ZN(n11873) );
  MUX2_X1 U14323 ( .A(n11874), .B(n11873), .S(n11872), .Z(n11875) );
  AND2_X1 U14324 ( .A1(n11876), .A2(n11875), .ZN(n11880) );
  MUX2_X1 U14325 ( .A(n11878), .B(n11877), .S(n11955), .Z(n11879) );
  OAI211_X1 U14326 ( .C1(n11880), .C2(n14996), .A(n10908), .B(n11879), .ZN(
        n11886) );
  OAI21_X1 U14327 ( .B1(n11882), .B2(n11881), .A(n11889), .ZN(n11883) );
  NAND2_X1 U14328 ( .A1(n11883), .A2(n11955), .ZN(n11885) );
  INV_X1 U14329 ( .A(n11888), .ZN(n11884) );
  AOI21_X1 U14330 ( .B1(n11886), .B2(n11885), .A(n11884), .ZN(n11891) );
  AOI21_X1 U14331 ( .B1(n11888), .B2(n11887), .A(n11955), .ZN(n11890) );
  OAI22_X1 U14332 ( .A1(n11891), .A2(n11890), .B1(n11955), .B2(n11889), .ZN(
        n11898) );
  INV_X1 U14333 ( .A(n11895), .ZN(n11892) );
  AND2_X1 U14334 ( .A1(n11892), .A2(n11893), .ZN(n14566) );
  INV_X1 U14335 ( .A(n11893), .ZN(n11894) );
  MUX2_X1 U14336 ( .A(n11895), .B(n11894), .S(n11936), .Z(n11897) );
  AOI211_X1 U14337 ( .C1(n11898), .C2(n14566), .A(n11897), .B(n11896), .ZN(
        n11905) );
  INV_X1 U14338 ( .A(n11899), .ZN(n11902) );
  INV_X1 U14339 ( .A(n11900), .ZN(n11901) );
  MUX2_X1 U14340 ( .A(n11902), .B(n11901), .S(n11955), .Z(n11904) );
  NOR3_X1 U14341 ( .A1(n11905), .A2(n11904), .A3(n11903), .ZN(n11914) );
  NAND2_X1 U14342 ( .A1(n11911), .A2(n11906), .ZN(n11909) );
  NAND2_X1 U14343 ( .A1(n11910), .A2(n11907), .ZN(n11908) );
  MUX2_X1 U14344 ( .A(n11909), .B(n11908), .S(n11936), .Z(n11913) );
  MUX2_X1 U14345 ( .A(n11911), .B(n11910), .S(n11955), .Z(n11912) );
  OAI21_X1 U14346 ( .B1(n11914), .B2(n11913), .A(n11912), .ZN(n11917) );
  INV_X1 U14347 ( .A(n11915), .ZN(n11916) );
  AOI22_X1 U14348 ( .A1(n11917), .A2(n6848), .B1(n11916), .B2(n11921), .ZN(
        n11918) );
  NOR2_X1 U14349 ( .A1(n11918), .A2(n12949), .ZN(n11919) );
  AOI21_X1 U14350 ( .B1(n11921), .B2(n11920), .A(n11919), .ZN(n11926) );
  INV_X1 U14351 ( .A(n11922), .ZN(n11924) );
  MUX2_X1 U14352 ( .A(n11924), .B(n7263), .S(n11955), .Z(n11925) );
  NOR3_X1 U14353 ( .A1(n12896), .A2(n12907), .A3(n12919), .ZN(n12004) );
  OAI21_X1 U14354 ( .B1(n11926), .B2(n11925), .A(n12004), .ZN(n11929) );
  MUX2_X1 U14355 ( .A(n11927), .B(n12884), .S(n11936), .Z(n11928) );
  OAI211_X1 U14356 ( .C1(n12896), .C2(n11930), .A(n11929), .B(n11928), .ZN(
        n11932) );
  NOR2_X1 U14357 ( .A1(n12899), .A2(n11936), .ZN(n11931) );
  AOI22_X1 U14358 ( .A1(n11932), .A2(n12886), .B1(n11931), .B2(n13012), .ZN(
        n11940) );
  NAND2_X1 U14359 ( .A1(n11934), .A2(n11933), .ZN(n11935) );
  NAND2_X1 U14360 ( .A1(n11935), .A2(n11938), .ZN(n11937) );
  MUX2_X1 U14361 ( .A(n11938), .B(n11937), .S(n11936), .Z(n11939) );
  OAI211_X1 U14362 ( .C1(n11940), .C2(n12868), .A(n12850), .B(n11939), .ZN(
        n11947) );
  INV_X1 U14363 ( .A(n11948), .ZN(n11941) );
  INV_X1 U14364 ( .A(n12833), .ZN(n12835) );
  NAND3_X1 U14365 ( .A1(n11947), .A2(n12835), .A3(n11942), .ZN(n11945) );
  INV_X1 U14366 ( .A(n11943), .ZN(n11944) );
  NAND2_X1 U14367 ( .A1(n11945), .A2(n11944), .ZN(n11951) );
  NAND3_X1 U14368 ( .A1(n11947), .A2(n12835), .A3(n11946), .ZN(n11949) );
  NAND2_X1 U14369 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  NAND2_X1 U14370 ( .A1(n12579), .A2(n12837), .ZN(n11952) );
  INV_X1 U14371 ( .A(n12812), .ZN(n12007) );
  NAND2_X1 U14372 ( .A1(n12007), .A2(n11955), .ZN(n11956) );
  NAND2_X1 U14373 ( .A1(n12381), .A2(n12809), .ZN(n12016) );
  OAI21_X1 U14374 ( .B1(n11957), .B2(n11956), .A(n12016), .ZN(n11964) );
  OR2_X1 U14375 ( .A1(n12381), .A2(n12809), .ZN(n12019) );
  INV_X1 U14376 ( .A(n11958), .ZN(n11959) );
  NAND2_X1 U14377 ( .A1(n14363), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11961) );
  XNOR2_X1 U14378 ( .A(n12374), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11967) );
  XNOR2_X1 U14379 ( .A(n11968), .B(n11967), .ZN(n12567) );
  NAND2_X1 U14380 ( .A1(n12567), .A2(n11971), .ZN(n11963) );
  OR2_X1 U14381 ( .A1(n11274), .A2(n12570), .ZN(n11962) );
  INV_X1 U14382 ( .A(n12675), .ZN(n11979) );
  NOR2_X1 U14383 ( .A1(n12015), .A2(n11979), .ZN(n12022) );
  INV_X1 U14384 ( .A(n12022), .ZN(n12008) );
  OAI211_X1 U14385 ( .C1(n11965), .C2(n11964), .A(n12019), .B(n12008), .ZN(
        n11983) );
  XNOR2_X1 U14386 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11969) );
  XNOR2_X1 U14387 ( .A(n11970), .B(n11969), .ZN(n13110) );
  NAND2_X1 U14388 ( .A1(n13110), .A2(n11971), .ZN(n11973) );
  INV_X1 U14389 ( .A(SI_31_), .ZN(n13116) );
  OR2_X1 U14390 ( .A1(n11274), .A2(n13116), .ZN(n11972) );
  NAND2_X1 U14391 ( .A1(n6530), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11977) );
  NAND2_X1 U14392 ( .A1(n6532), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U14393 ( .A1(n6944), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11975) );
  AND4_X1 U14394 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n12802) );
  OR2_X1 U14395 ( .A1(n12986), .A2(n12802), .ZN(n11981) );
  NAND2_X1 U14396 ( .A1(n12015), .A2(n11979), .ZN(n11980) );
  INV_X1 U14397 ( .A(n12018), .ZN(n11982) );
  INV_X1 U14398 ( .A(n12802), .ZN(n12674) );
  NOR2_X1 U14399 ( .A1(n13043), .A2(n12674), .ZN(n12021) );
  AOI21_X1 U14400 ( .B1(n11983), .B2(n11982), .A(n12021), .ZN(n12029) );
  INV_X1 U14401 ( .A(n15056), .ZN(n15076) );
  INV_X1 U14402 ( .A(n12850), .ZN(n12848) );
  INV_X1 U14403 ( .A(n12932), .ZN(n12929) );
  NAND4_X1 U14404 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11993) );
  NAND4_X1 U14405 ( .A1(n11989), .A2(n11990), .A3(n11991), .A4(n11988), .ZN(
        n11992) );
  NOR2_X1 U14406 ( .A1(n11993), .A2(n11992), .ZN(n11996) );
  NOR2_X1 U14407 ( .A1(n11994), .A2(n15015), .ZN(n11995) );
  NAND4_X1 U14408 ( .A1(n11996), .A2(n12979), .A3(n6707), .A4(n11995), .ZN(
        n11997) );
  NOR2_X1 U14409 ( .A1(n11997), .A2(n14578), .ZN(n12000) );
  NAND4_X1 U14410 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n14566), .ZN(
        n12001) );
  NOR4_X1 U14411 ( .A1(n12949), .A2(n12958), .A3(n12002), .A4(n12001), .ZN(
        n12003) );
  NAND4_X1 U14412 ( .A1(n12004), .A2(n12929), .A3(n12003), .A4(n12886), .ZN(
        n12005) );
  NOR4_X1 U14413 ( .A1(n12833), .A2(n12848), .A3(n12868), .A4(n12005), .ZN(
        n12006) );
  NAND4_X1 U14414 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12826), .ZN(
        n12011) );
  INV_X1 U14415 ( .A(n12009), .ZN(n12010) );
  XNOR2_X1 U14416 ( .A(n12012), .B(n12771), .ZN(n12013) );
  OAI22_X1 U14417 ( .A1(n12029), .A2(n15076), .B1(n12014), .B2(n12013), .ZN(
        n12028) );
  OAI21_X1 U14418 ( .B1(n13046), .B2(n12674), .A(n12016), .ZN(n12017) );
  INV_X1 U14419 ( .A(n12024), .ZN(n12025) );
  AND2_X2 U14420 ( .A1(n12026), .A2(n12025), .ZN(n12027) );
  NAND3_X1 U14421 ( .A1(n12032), .A2(n12031), .A3(n12777), .ZN(n12033) );
  OAI211_X1 U14422 ( .C1(n12034), .C2(n12036), .A(n12033), .B(P3_B_REG_SCAN_IN), .ZN(n12035) );
  OAI21_X1 U14423 ( .B1(n12037), .B2(n12036), .A(n12035), .ZN(P3_U3296) );
  NAND2_X1 U14424 ( .A1(n12302), .A2(n12305), .ZN(n12234) );
  OAI21_X1 U14425 ( .B1(n12038), .B2(n12044), .A(n12234), .ZN(n12260) );
  NAND2_X1 U14426 ( .A1(n12301), .A2(n12044), .ZN(n12039) );
  OAI211_X1 U14427 ( .C1(n7130), .C2(n12305), .A(n12304), .B(n12039), .ZN(
        n12259) );
  NAND2_X1 U14428 ( .A1(n12041), .A2(n12213), .ZN(n12047) );
  OAI21_X1 U14429 ( .B1(n12305), .B2(n12044), .A(n12043), .ZN(n12045) );
  NAND2_X1 U14430 ( .A1(n12046), .A2(n12045), .ZN(n12050) );
  NAND2_X1 U14431 ( .A1(n13269), .A2(n12213), .ZN(n12052) );
  NAND2_X1 U14432 ( .A1(n12053), .A2(n12070), .ZN(n12051) );
  NAND2_X1 U14433 ( .A1(n12052), .A2(n12051), .ZN(n12056) );
  AOI22_X1 U14434 ( .A1(n13269), .A2(n12070), .B1(n12053), .B2(n12213), .ZN(
        n12054) );
  NAND2_X1 U14435 ( .A1(n13267), .A2(n12070), .ZN(n12059) );
  NAND2_X1 U14436 ( .A1(n7852), .A2(n12213), .ZN(n12058) );
  NAND2_X1 U14437 ( .A1(n12059), .A2(n12058), .ZN(n12061) );
  AOI22_X1 U14438 ( .A1(n13267), .A2(n12213), .B1(n12070), .B2(n7852), .ZN(
        n12060) );
  NAND2_X1 U14439 ( .A1(n13266), .A2(n12213), .ZN(n12063) );
  NAND2_X1 U14440 ( .A1(n14901), .A2(n12070), .ZN(n12062) );
  NAND2_X1 U14441 ( .A1(n12063), .A2(n12062), .ZN(n12068) );
  NAND2_X1 U14442 ( .A1(n13266), .A2(n12242), .ZN(n12065) );
  NAND2_X1 U14443 ( .A1(n14901), .A2(n12213), .ZN(n12064) );
  NAND2_X1 U14444 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  INV_X1 U14445 ( .A(n12068), .ZN(n12069) );
  NAND2_X1 U14446 ( .A1(n13265), .A2(n12237), .ZN(n12072) );
  NAND2_X1 U14447 ( .A1(n14936), .A2(n12228), .ZN(n12071) );
  NAND2_X1 U14448 ( .A1(n12072), .A2(n12071), .ZN(n12074) );
  AOI22_X1 U14449 ( .A1(n13265), .A2(n12213), .B1(n12242), .B2(n14936), .ZN(
        n12073) );
  NAND2_X1 U14450 ( .A1(n13264), .A2(n12228), .ZN(n12077) );
  NAND2_X1 U14451 ( .A1(n13184), .A2(n12237), .ZN(n12076) );
  NAND2_X1 U14452 ( .A1(n12077), .A2(n12076), .ZN(n12079) );
  AOI22_X1 U14453 ( .A1(n12237), .A2(n13264), .B1(n13184), .B2(n12228), .ZN(
        n12078) );
  AOI21_X1 U14454 ( .B1(n12080), .B2(n12079), .A(n12078), .ZN(n12082) );
  AOI22_X1 U14455 ( .A1(n12084), .A2(n12228), .B1(n12237), .B2(n13263), .ZN(
        n12088) );
  INV_X1 U14456 ( .A(n12088), .ZN(n12083) );
  NAND2_X1 U14457 ( .A1(n12084), .A2(n12237), .ZN(n12085) );
  OAI21_X1 U14458 ( .B1(n12086), .B2(n12242), .A(n12085), .ZN(n12087) );
  NAND2_X1 U14459 ( .A1(n12091), .A2(n12237), .ZN(n12090) );
  NAND2_X1 U14460 ( .A1(n13262), .A2(n12228), .ZN(n12089) );
  NAND2_X1 U14461 ( .A1(n12090), .A2(n12089), .ZN(n12094) );
  AOI22_X1 U14462 ( .A1(n12091), .A2(n12213), .B1(n12237), .B2(n13262), .ZN(
        n12092) );
  AOI21_X1 U14463 ( .B1(n12095), .B2(n12094), .A(n12092), .ZN(n12093) );
  NAND2_X1 U14464 ( .A1(n14952), .A2(n12213), .ZN(n12097) );
  NAND2_X1 U14465 ( .A1(n13261), .A2(n12237), .ZN(n12096) );
  NAND2_X1 U14466 ( .A1(n14952), .A2(n12237), .ZN(n12098) );
  OAI21_X1 U14467 ( .B1(n12099), .B2(n12242), .A(n12098), .ZN(n12100) );
  NAND2_X1 U14468 ( .A1(n12103), .A2(n12237), .ZN(n12102) );
  NAND2_X1 U14469 ( .A1(n13260), .A2(n12213), .ZN(n12101) );
  NAND2_X1 U14470 ( .A1(n12102), .A2(n12101), .ZN(n12106) );
  AOI22_X1 U14471 ( .A1(n12103), .A2(n12213), .B1(n12237), .B2(n13260), .ZN(
        n12104) );
  NAND2_X1 U14472 ( .A1(n13601), .A2(n12213), .ZN(n12109) );
  NAND2_X1 U14473 ( .A1(n13259), .A2(n12237), .ZN(n12108) );
  NAND2_X1 U14474 ( .A1(n13601), .A2(n12237), .ZN(n12110) );
  OAI21_X1 U14475 ( .B1(n12111), .B2(n12242), .A(n12110), .ZN(n12112) );
  NAND2_X1 U14476 ( .A1(n12115), .A2(n12237), .ZN(n12114) );
  NAND2_X1 U14477 ( .A1(n13258), .A2(n12228), .ZN(n12113) );
  NAND2_X1 U14478 ( .A1(n12114), .A2(n12113), .ZN(n12117) );
  AOI22_X1 U14479 ( .A1(n12115), .A2(n12213), .B1(n12237), .B2(n13258), .ZN(
        n12116) );
  NAND2_X1 U14480 ( .A1(n13587), .A2(n12213), .ZN(n12119) );
  NAND2_X1 U14481 ( .A1(n13257), .A2(n12237), .ZN(n12118) );
  NAND2_X1 U14482 ( .A1(n12119), .A2(n12118), .ZN(n12121) );
  AOI22_X1 U14483 ( .A1(n13587), .A2(n12237), .B1(n13257), .B2(n12228), .ZN(
        n12120) );
  AND2_X1 U14484 ( .A1(n13256), .A2(n12237), .ZN(n12123) );
  AOI21_X1 U14485 ( .B1(n14819), .B2(n12228), .A(n12123), .ZN(n12143) );
  NAND2_X1 U14486 ( .A1(n14819), .A2(n12237), .ZN(n12125) );
  NAND2_X1 U14487 ( .A1(n13256), .A2(n12228), .ZN(n12124) );
  NAND2_X1 U14488 ( .A1(n12125), .A2(n12124), .ZN(n12142) );
  AOI22_X1 U14489 ( .A1(n13739), .A2(n12228), .B1(n12237), .B2(n13252), .ZN(
        n12128) );
  NAND2_X1 U14490 ( .A1(n13739), .A2(n12237), .ZN(n12127) );
  NAND2_X1 U14491 ( .A1(n13252), .A2(n12228), .ZN(n12126) );
  NAND2_X1 U14492 ( .A1(n12127), .A2(n12126), .ZN(n12154) );
  NAND2_X1 U14493 ( .A1(n12128), .A2(n12154), .ZN(n12133) );
  AND2_X1 U14494 ( .A1(n13253), .A2(n12237), .ZN(n12129) );
  AOI21_X1 U14495 ( .B1(n13743), .B2(n12213), .A(n12129), .ZN(n12150) );
  NAND2_X1 U14496 ( .A1(n13743), .A2(n12237), .ZN(n12131) );
  NAND2_X1 U14497 ( .A1(n13253), .A2(n12213), .ZN(n12130) );
  NAND2_X1 U14498 ( .A1(n12131), .A2(n12130), .ZN(n12149) );
  NAND2_X1 U14499 ( .A1(n12150), .A2(n12149), .ZN(n12132) );
  NAND2_X1 U14500 ( .A1(n12133), .A2(n12132), .ZN(n12148) );
  AND2_X1 U14501 ( .A1(n13254), .A2(n12237), .ZN(n12134) );
  AOI21_X1 U14502 ( .B1(n13696), .B2(n12213), .A(n12134), .ZN(n12152) );
  NAND2_X1 U14503 ( .A1(n13696), .A2(n12237), .ZN(n12136) );
  NAND2_X1 U14504 ( .A1(n13254), .A2(n12213), .ZN(n12135) );
  NAND2_X1 U14505 ( .A1(n12136), .A2(n12135), .ZN(n12151) );
  AND2_X1 U14506 ( .A1(n12152), .A2(n12151), .ZN(n12137) );
  AND2_X1 U14507 ( .A1(n13255), .A2(n12237), .ZN(n12138) );
  AOI21_X1 U14508 ( .B1(n12139), .B2(n12213), .A(n12138), .ZN(n12147) );
  NAND2_X1 U14509 ( .A1(n12139), .A2(n12237), .ZN(n12141) );
  NAND2_X1 U14510 ( .A1(n13255), .A2(n12213), .ZN(n12140) );
  NAND2_X1 U14511 ( .A1(n12141), .A2(n12140), .ZN(n12146) );
  AOI22_X1 U14512 ( .A1(n12147), .A2(n12146), .B1(n12143), .B2(n12142), .ZN(
        n12144) );
  INV_X1 U14513 ( .A(n12148), .ZN(n12157) );
  OAI22_X1 U14514 ( .A1(n12152), .A2(n12151), .B1(n12150), .B2(n12149), .ZN(
        n12156) );
  NOR2_X1 U14515 ( .A1(n13739), .A2(n13252), .ZN(n12153) );
  NOR2_X1 U14516 ( .A1(n12154), .A2(n12153), .ZN(n12155) );
  AOI21_X1 U14517 ( .B1(n12157), .B2(n12156), .A(n12155), .ZN(n12158) );
  AND2_X1 U14518 ( .A1(n12159), .A2(n12158), .ZN(n12165) );
  NAND2_X1 U14519 ( .A1(n13735), .A2(n12228), .ZN(n12161) );
  NAND2_X1 U14520 ( .A1(n13251), .A2(n12237), .ZN(n12160) );
  NAND2_X1 U14521 ( .A1(n12161), .A2(n12160), .ZN(n12168) );
  INV_X1 U14522 ( .A(n12168), .ZN(n12162) );
  NAND2_X1 U14523 ( .A1(n13735), .A2(n12237), .ZN(n12164) );
  OAI21_X1 U14524 ( .B1(n13140), .B2(n12242), .A(n12164), .ZN(n12167) );
  AND2_X1 U14525 ( .A1(n12165), .A2(n12167), .ZN(n12166) );
  INV_X1 U14526 ( .A(n12167), .ZN(n12169) );
  OR2_X1 U14527 ( .A1(n12169), .A2(n12168), .ZN(n12170) );
  NAND2_X1 U14528 ( .A1(n13672), .A2(n12237), .ZN(n12173) );
  NAND2_X1 U14529 ( .A1(n13250), .A2(n12213), .ZN(n12172) );
  NAND2_X1 U14530 ( .A1(n12173), .A2(n12172), .ZN(n12175) );
  AOI22_X1 U14531 ( .A1(n13672), .A2(n12213), .B1(n12237), .B2(n13250), .ZN(
        n12174) );
  NAND2_X1 U14532 ( .A1(n13529), .A2(n12213), .ZN(n12178) );
  NAND2_X1 U14533 ( .A1(n13249), .A2(n12237), .ZN(n12177) );
  NAND2_X1 U14534 ( .A1(n12178), .A2(n12177), .ZN(n12180) );
  AOI22_X1 U14535 ( .A1(n13529), .A2(n12237), .B1(n13249), .B2(n12213), .ZN(
        n12179) );
  NAND2_X1 U14536 ( .A1(n13512), .A2(n12237), .ZN(n12182) );
  NAND2_X1 U14537 ( .A1(n13248), .A2(n12213), .ZN(n12181) );
  NAND2_X1 U14538 ( .A1(n12182), .A2(n12181), .ZN(n12184) );
  AOI22_X1 U14539 ( .A1(n13512), .A2(n12213), .B1(n12237), .B2(n13248), .ZN(
        n12183) );
  NAND2_X1 U14540 ( .A1(n13653), .A2(n12213), .ZN(n12186) );
  NAND2_X1 U14541 ( .A1(n13247), .A2(n12237), .ZN(n12185) );
  NAND2_X1 U14542 ( .A1(n12186), .A2(n12185), .ZN(n12188) );
  AOI22_X1 U14543 ( .A1(n13653), .A2(n12237), .B1(n13247), .B2(n12228), .ZN(
        n12187) );
  NAND2_X1 U14544 ( .A1(n13648), .A2(n12237), .ZN(n12191) );
  NAND2_X1 U14545 ( .A1(n13246), .A2(n12228), .ZN(n12190) );
  NAND2_X1 U14546 ( .A1(n12191), .A2(n12190), .ZN(n12193) );
  AOI22_X1 U14547 ( .A1(n13648), .A2(n12213), .B1(n12237), .B2(n13246), .ZN(
        n12192) );
  NAND2_X1 U14548 ( .A1(n13643), .A2(n12228), .ZN(n12195) );
  NAND2_X1 U14549 ( .A1(n13245), .A2(n12237), .ZN(n12194) );
  NAND2_X1 U14550 ( .A1(n12195), .A2(n12194), .ZN(n12198) );
  NAND2_X1 U14551 ( .A1(n13643), .A2(n12237), .ZN(n12196) );
  OAI21_X1 U14552 ( .B1(n13167), .B2(n12242), .A(n12196), .ZN(n12197) );
  NAND2_X1 U14553 ( .A1(n13638), .A2(n12237), .ZN(n12200) );
  NAND2_X1 U14554 ( .A1(n13244), .A2(n12213), .ZN(n12199) );
  NAND2_X1 U14555 ( .A1(n12200), .A2(n12199), .ZN(n12202) );
  AOI22_X1 U14556 ( .A1(n13638), .A2(n12213), .B1(n12237), .B2(n13244), .ZN(
        n12201) );
  NAND2_X1 U14557 ( .A1(n13440), .A2(n12228), .ZN(n12204) );
  NAND2_X1 U14558 ( .A1(n13243), .A2(n12242), .ZN(n12203) );
  NAND2_X1 U14559 ( .A1(n12204), .A2(n12203), .ZN(n12206) );
  AOI22_X1 U14560 ( .A1(n13440), .A2(n12242), .B1(n13243), .B2(n12213), .ZN(
        n12205) );
  AOI21_X1 U14561 ( .B1(n12207), .B2(n12206), .A(n12205), .ZN(n12209) );
  NOR2_X1 U14562 ( .A1(n12207), .A2(n12206), .ZN(n12208) );
  NAND2_X1 U14563 ( .A1(n13424), .A2(n12237), .ZN(n12211) );
  NAND2_X1 U14564 ( .A1(n13242), .A2(n12213), .ZN(n12210) );
  AND2_X1 U14565 ( .A1(n13241), .A2(n12237), .ZN(n12212) );
  AOI21_X1 U14566 ( .B1(n13409), .B2(n12213), .A(n12212), .ZN(n12248) );
  NAND2_X1 U14567 ( .A1(n13409), .A2(n12242), .ZN(n12215) );
  NAND2_X1 U14568 ( .A1(n13241), .A2(n12228), .ZN(n12214) );
  NAND2_X1 U14569 ( .A1(n12215), .A2(n12214), .ZN(n12247) );
  INV_X1 U14570 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13750) );
  OR2_X1 U14571 ( .A1(n7832), .A2(n13750), .ZN(n12217) );
  INV_X1 U14572 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U14573 ( .A1(n12218), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12220) );
  NAND2_X1 U14574 ( .A1(n8361), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12219) );
  OAI211_X1 U14575 ( .C1(n6525), .C2(n12221), .A(n12220), .B(n12219), .ZN(
        n13390) );
  XNOR2_X1 U14576 ( .A(n13386), .B(n13390), .ZN(n12298) );
  AND2_X1 U14577 ( .A1(n13240), .A2(n12228), .ZN(n12223) );
  AOI21_X1 U14578 ( .B1(n13616), .B2(n12242), .A(n12223), .ZN(n12241) );
  NAND2_X1 U14579 ( .A1(n13616), .A2(n12213), .ZN(n12225) );
  NAND2_X1 U14580 ( .A1(n13240), .A2(n12237), .ZN(n12224) );
  NAND2_X1 U14581 ( .A1(n12225), .A2(n12224), .ZN(n12240) );
  NAND2_X1 U14582 ( .A1(n12241), .A2(n12240), .ZN(n12249) );
  OAI211_X1 U14583 ( .C1(n12248), .C2(n12247), .A(n12298), .B(n12249), .ZN(
        n12226) );
  INV_X1 U14584 ( .A(n12226), .ZN(n12227) );
  AOI22_X1 U14585 ( .A1(n13424), .A2(n12228), .B1(n12237), .B2(n13242), .ZN(
        n12229) );
  NAND2_X1 U14586 ( .A1(n12231), .A2(n12230), .ZN(n12233) );
  OR2_X1 U14587 ( .A1(n7832), .A2(n12374), .ZN(n12232) );
  NAND2_X1 U14588 ( .A1(n13390), .A2(n12213), .ZN(n12254) );
  NAND4_X1 U14589 ( .A1(n12254), .A2(n12301), .A3(n12234), .A4(n12304), .ZN(
        n12235) );
  AND2_X1 U14590 ( .A1(n12235), .A2(n13239), .ZN(n12236) );
  AOI21_X1 U14591 ( .B1(n13396), .B2(n12242), .A(n12236), .ZN(n12253) );
  NAND2_X1 U14592 ( .A1(n13396), .A2(n12213), .ZN(n12239) );
  NAND2_X1 U14593 ( .A1(n13239), .A2(n12237), .ZN(n12238) );
  NAND2_X1 U14594 ( .A1(n12239), .A2(n12238), .ZN(n12252) );
  OAI22_X1 U14595 ( .A1(n12253), .A2(n12252), .B1(n12241), .B2(n12240), .ZN(
        n12246) );
  MUX2_X1 U14596 ( .A(n13390), .B(n12242), .S(n13386), .Z(n12244) );
  NAND2_X1 U14597 ( .A1(n13390), .A2(n12242), .ZN(n12243) );
  NAND2_X1 U14598 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  NAND2_X1 U14599 ( .A1(n12246), .A2(n12245), .ZN(n12251) );
  NAND4_X1 U14600 ( .A1(n12249), .A2(n12298), .A3(n12248), .A4(n12247), .ZN(
        n12250) );
  NAND2_X1 U14601 ( .A1(n12253), .A2(n12252), .ZN(n12258) );
  AND2_X1 U14602 ( .A1(n13390), .A2(n12242), .ZN(n12256) );
  AND2_X1 U14603 ( .A1(n12254), .A2(n12213), .ZN(n12255) );
  MUX2_X1 U14604 ( .A(n12256), .B(n12255), .S(n13386), .Z(n12257) );
  NAND4_X1 U14605 ( .A1(n12265), .A2(n12264), .A3(n12263), .A4(n12262), .ZN(
        n12267) );
  NOR3_X1 U14606 ( .A1(n12267), .A2(n12266), .A3(n14886), .ZN(n12271) );
  NAND4_X1 U14607 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  NOR2_X1 U14608 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  NAND2_X1 U14609 ( .A1(n12275), .A2(n12274), .ZN(n12276) );
  NOR2_X1 U14610 ( .A1(n12277), .A2(n12276), .ZN(n12280) );
  NAND4_X1 U14611 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NOR2_X1 U14612 ( .A1(n12283), .A2(n12282), .ZN(n12286) );
  NAND4_X1 U14613 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  NOR2_X1 U14614 ( .A1(n13525), .A2(n12288), .ZN(n12289) );
  NAND4_X1 U14615 ( .A1(n13506), .A2(n12289), .A3(n13536), .A4(n13552), .ZN(
        n12290) );
  NOR2_X1 U14616 ( .A1(n13494), .A2(n12290), .ZN(n12293) );
  NAND2_X1 U14617 ( .A1(n12292), .A2(n12291), .ZN(n13478) );
  NAND4_X1 U14618 ( .A1(n12294), .A2(n12293), .A3(n13464), .A4(n13478), .ZN(
        n12295) );
  XOR2_X1 U14619 ( .A(n13239), .B(n13707), .Z(n12300) );
  NOR4_X1 U14620 ( .A1(n13191), .A2(n14913), .A3(n12304), .A4(n13761), .ZN(
        n12307) );
  OAI21_X1 U14621 ( .B1(n12308), .B2(n12305), .A(P2_B_REG_SCAN_IN), .ZN(n12306) );
  INV_X1 U14622 ( .A(n12309), .ZN(n12310) );
  XNOR2_X1 U14623 ( .A(n13739), .B(n6529), .ZN(n12325) );
  NAND2_X1 U14624 ( .A1(n13252), .A2(n13542), .ZN(n12323) );
  XNOR2_X1 U14625 ( .A(n12325), .B(n12323), .ZN(n12317) );
  NAND2_X1 U14626 ( .A1(n13251), .A2(n13230), .ZN(n12313) );
  NAND2_X1 U14627 ( .A1(n13253), .A2(n13231), .ZN(n12312) );
  NAND2_X1 U14628 ( .A1(n12313), .A2(n12312), .ZN(n13569) );
  AOI22_X1 U14629 ( .A1(n13235), .A2(n13569), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12314) );
  OAI21_X1 U14630 ( .B1(n13574), .B2(n14821), .A(n12314), .ZN(n12321) );
  INV_X1 U14631 ( .A(n12315), .ZN(n12319) );
  AOI22_X1 U14632 ( .A1(n12316), .A2(n13227), .B1(n13205), .B2(n13253), .ZN(
        n12318) );
  NOR3_X1 U14633 ( .A1(n12319), .A2(n12318), .A3(n12317), .ZN(n12320) );
  AOI211_X1 U14634 ( .C1(n13739), .C2(n14818), .A(n12321), .B(n12320), .ZN(
        n12322) );
  OAI21_X1 U14635 ( .B1(n12327), .B2(n14813), .A(n12322), .ZN(P2_U3200) );
  INV_X1 U14636 ( .A(n12323), .ZN(n12324) );
  XNOR2_X1 U14637 ( .A(n13735), .B(n12356), .ZN(n13141) );
  NAND2_X1 U14638 ( .A1(n13251), .A2(n13542), .ZN(n12328) );
  NOR2_X1 U14639 ( .A1(n13141), .A2(n12328), .ZN(n12329) );
  AOI21_X1 U14640 ( .B1(n13141), .B2(n12328), .A(n12329), .ZN(n13229) );
  NAND2_X1 U14641 ( .A1(n13250), .A2(n13542), .ZN(n12332) );
  XNOR2_X1 U14642 ( .A(n13206), .B(n12332), .ZN(n13150) );
  INV_X1 U14643 ( .A(n12329), .ZN(n12330) );
  INV_X1 U14644 ( .A(n12332), .ZN(n12333) );
  XNOR2_X1 U14645 ( .A(n13529), .B(n6529), .ZN(n12334) );
  NAND2_X1 U14646 ( .A1(n13249), .A2(n13542), .ZN(n12335) );
  XNOR2_X1 U14647 ( .A(n12334), .B(n12335), .ZN(n13207) );
  INV_X1 U14648 ( .A(n12334), .ZN(n12336) );
  NAND2_X1 U14649 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  NAND2_X1 U14650 ( .A1(n13248), .A2(n13542), .ZN(n12338) );
  XNOR2_X1 U14651 ( .A(n13512), .B(n6529), .ZN(n12340) );
  XOR2_X1 U14652 ( .A(n12338), .B(n12340), .Z(n13152) );
  INV_X1 U14653 ( .A(n12338), .ZN(n12339) );
  NAND2_X1 U14654 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  XNOR2_X1 U14655 ( .A(n13653), .B(n6529), .ZN(n12343) );
  NAND2_X1 U14656 ( .A1(n12342), .A2(n12343), .ZN(n12344) );
  XNOR2_X1 U14657 ( .A(n13648), .B(n6529), .ZN(n12346) );
  NAND2_X1 U14658 ( .A1(n12347), .A2(n12346), .ZN(n12348) );
  XNOR2_X1 U14659 ( .A(n13643), .B(n12356), .ZN(n13164) );
  NAND2_X1 U14660 ( .A1(n13245), .A2(n13542), .ZN(n12349) );
  NOR2_X1 U14661 ( .A1(n13164), .A2(n12349), .ZN(n12350) );
  AOI21_X1 U14662 ( .B1(n13164), .B2(n12349), .A(n12350), .ZN(n13190) );
  INV_X1 U14663 ( .A(n12350), .ZN(n12351) );
  XNOR2_X1 U14664 ( .A(n13638), .B(n6529), .ZN(n12352) );
  AND2_X1 U14665 ( .A1(n13244), .A2(n13542), .ZN(n12353) );
  NAND2_X1 U14666 ( .A1(n12352), .A2(n12353), .ZN(n12357) );
  INV_X1 U14667 ( .A(n12352), .ZN(n12361) );
  INV_X1 U14668 ( .A(n12353), .ZN(n12354) );
  NAND2_X1 U14669 ( .A1(n12361), .A2(n12354), .ZN(n12355) );
  XNOR2_X1 U14670 ( .A(n13440), .B(n12356), .ZN(n12393) );
  NAND2_X1 U14671 ( .A1(n13243), .A2(n13542), .ZN(n12392) );
  XNOR2_X1 U14672 ( .A(n12393), .B(n12392), .ZN(n12362) );
  INV_X1 U14673 ( .A(n12357), .ZN(n12358) );
  NOR2_X1 U14674 ( .A1(n12362), .A2(n12358), .ZN(n12359) );
  NOR2_X1 U14675 ( .A1(n12360), .A2(n14813), .ZN(n12364) );
  NOR3_X1 U14676 ( .A1(n12361), .A2(n13194), .A3(n13213), .ZN(n12363) );
  OAI21_X1 U14677 ( .B1(n12364), .B2(n12363), .A(n12362), .ZN(n12370) );
  NAND2_X1 U14678 ( .A1(n13244), .A2(n13231), .ZN(n12366) );
  NAND2_X1 U14679 ( .A1(n13242), .A2(n13230), .ZN(n12365) );
  NAND2_X1 U14680 ( .A1(n12366), .A2(n12365), .ZN(n13430) );
  AOI22_X1 U14681 ( .A1(n13235), .A2(n13430), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12367) );
  OAI21_X1 U14682 ( .B1(n13437), .B2(n14821), .A(n12367), .ZN(n12368) );
  AOI21_X1 U14683 ( .B1(n13440), .B2(n14818), .A(n12368), .ZN(n12369) );
  OAI211_X1 U14684 ( .C1(n14813), .C2(n12395), .A(n12370), .B(n12369), .ZN(
        P2_U3212) );
  INV_X1 U14685 ( .A(n12371), .ZN(n14365) );
  OAI222_X1 U14686 ( .A1(n13766), .A2(n14365), .B1(P2_U3088), .B2(n12373), 
        .C1(n12372), .C2(n13764), .ZN(P2_U3298) );
  OAI222_X1 U14687 ( .A1(n13766), .A2(n12376), .B1(P2_U3088), .B2(n12375), 
        .C1(n12374), .C2(n13764), .ZN(P2_U3297) );
  INV_X1 U14688 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12377) );
  MUX2_X1 U14689 ( .A(n12377), .B(n12380), .S(n15080), .Z(n12379) );
  AOI22_X1 U14690 ( .A1(n12381), .A2(n15038), .B1(n12799), .B2(n15075), .ZN(
        n12378) );
  INV_X1 U14691 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n15305) );
  NAND2_X1 U14692 ( .A1(n12381), .A2(n13095), .ZN(n12382) );
  INV_X1 U14693 ( .A(n12384), .ZN(n12385) );
  AOI22_X1 U14694 ( .A1(n12385), .A2(n13227), .B1(n13205), .B2(n13254), .ZN(
        n12390) );
  AOI22_X1 U14695 ( .A1(n13235), .A2(n13695), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12386) );
  OAI21_X1 U14696 ( .B1(n12387), .B2(n14821), .A(n12386), .ZN(n12388) );
  AOI21_X1 U14697 ( .B1(n13696), .B2(n14818), .A(n12388), .ZN(n12389) );
  OAI21_X1 U14698 ( .B1(n12391), .B2(n12390), .A(n12389), .ZN(P2_U3213) );
  NAND2_X1 U14699 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  XNOR2_X1 U14700 ( .A(n13424), .B(n6529), .ZN(n12397) );
  AND2_X1 U14701 ( .A1(n13242), .A2(n13542), .ZN(n12396) );
  NAND2_X1 U14702 ( .A1(n12397), .A2(n12396), .ZN(n12399) );
  OAI21_X1 U14703 ( .B1(n12397), .B2(n12396), .A(n12399), .ZN(n13123) );
  NAND2_X1 U14704 ( .A1(n13241), .A2(n13542), .ZN(n12400) );
  XNOR2_X1 U14705 ( .A(n12400), .B(n6529), .ZN(n12401) );
  XNOR2_X1 U14706 ( .A(n13409), .B(n12401), .ZN(n12402) );
  NOR2_X1 U14707 ( .A1(n14821), .A2(n13400), .ZN(n12405) );
  AOI22_X1 U14708 ( .A1(n13230), .A2(n13240), .B1(n13242), .B2(n13231), .ZN(
        n13403) );
  OAI22_X1 U14709 ( .A1(n14811), .A2(n13403), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12403), .ZN(n12404) );
  AOI211_X1 U14710 ( .C1(n13409), .C2(n14818), .A(n12405), .B(n12404), .ZN(
        n12406) );
  OAI21_X1 U14711 ( .B1(n12407), .B2(n14813), .A(n12406), .ZN(P2_U3192) );
  OR2_X1 U14712 ( .A1(n14506), .A2(n12545), .ZN(n12409) );
  NAND2_X1 U14713 ( .A1(n12553), .A2(n13945), .ZN(n12408) );
  NAND2_X1 U14714 ( .A1(n12409), .A2(n12408), .ZN(n12420) );
  INV_X1 U14715 ( .A(n12420), .ZN(n12424) );
  OAI22_X1 U14716 ( .A1(n14506), .A2(n6907), .B1(n12410), .B2(n12542), .ZN(
        n12411) );
  XNOR2_X1 U14717 ( .A(n12411), .B(n12551), .ZN(n12419) );
  INV_X1 U14718 ( .A(n12419), .ZN(n12423) );
  NAND2_X1 U14719 ( .A1(n12413), .A2(n12412), .ZN(n12416) );
  INV_X1 U14720 ( .A(n12413), .ZN(n12415) );
  AOI22_X1 U14721 ( .A1(n14672), .A2(n12554), .B1(n12553), .B2(n13946), .ZN(
        n12421) );
  AOI22_X1 U14722 ( .A1(n14672), .A2(n6923), .B1(n12554), .B2(n13946), .ZN(
        n12418) );
  XNOR2_X1 U14723 ( .A(n12418), .B(n12551), .ZN(n12422) );
  XOR2_X1 U14724 ( .A(n12421), .B(n12422), .Z(n14611) );
  XOR2_X1 U14725 ( .A(n12420), .B(n12419), .Z(n13822) );
  NAND2_X1 U14726 ( .A1(n12422), .A2(n12421), .ZN(n13820) );
  NAND2_X1 U14727 ( .A1(n14666), .A2(n6923), .ZN(n12426) );
  NAND2_X1 U14728 ( .A1(n12554), .A2(n13944), .ZN(n12425) );
  NAND2_X1 U14729 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  XNOR2_X1 U14730 ( .A(n12427), .B(n12551), .ZN(n12429) );
  AOI22_X1 U14731 ( .A1(n14666), .A2(n12554), .B1(n12553), .B2(n13944), .ZN(
        n12428) );
  XNOR2_X1 U14732 ( .A(n12429), .B(n12428), .ZN(n13879) );
  INV_X1 U14733 ( .A(n12428), .ZN(n12430) );
  NAND2_X1 U14734 ( .A1(n14258), .A2(n6923), .ZN(n12432) );
  NAND2_X1 U14735 ( .A1(n12554), .A2(n13943), .ZN(n12431) );
  NAND2_X1 U14736 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  XNOR2_X1 U14737 ( .A(n12433), .B(n12522), .ZN(n12436) );
  INV_X1 U14738 ( .A(n12436), .ZN(n12438) );
  NOR2_X1 U14739 ( .A1(n13882), .A2(n12525), .ZN(n12434) );
  AOI21_X1 U14740 ( .B1(n14258), .B2(n12554), .A(n12434), .ZN(n12435) );
  INV_X1 U14741 ( .A(n12435), .ZN(n12437) );
  AND2_X1 U14742 ( .A1(n12436), .A2(n12435), .ZN(n12439) );
  AOI21_X1 U14743 ( .B1(n12438), .B2(n12437), .A(n12439), .ZN(n13779) );
  INV_X1 U14744 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14745 ( .A1(n13930), .A2(n6923), .ZN(n12442) );
  NAND2_X1 U14746 ( .A1(n13942), .A2(n12554), .ZN(n12441) );
  NAND2_X1 U14747 ( .A1(n12442), .A2(n12441), .ZN(n12443) );
  XNOR2_X1 U14748 ( .A(n12443), .B(n12551), .ZN(n12445) );
  OAI22_X1 U14749 ( .A1(n7497), .A2(n12542), .B1(n14630), .B2(n12525), .ZN(
        n13922) );
  INV_X1 U14750 ( .A(n12444), .ZN(n12446) );
  NAND2_X1 U14751 ( .A1(n14645), .A2(n6923), .ZN(n12449) );
  NAND2_X1 U14752 ( .A1(n13941), .A2(n12554), .ZN(n12448) );
  NAND2_X1 U14753 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  XNOR2_X1 U14754 ( .A(n12450), .B(n12522), .ZN(n12453) );
  AND2_X1 U14755 ( .A1(n13941), .A2(n12553), .ZN(n12451) );
  AOI21_X1 U14756 ( .B1(n14645), .B2(n12554), .A(n12451), .ZN(n12452) );
  NAND2_X1 U14757 ( .A1(n12453), .A2(n12452), .ZN(n13849) );
  OAI21_X1 U14758 ( .B1(n12453), .B2(n12452), .A(n13849), .ZN(n13842) );
  NAND2_X1 U14759 ( .A1(n14343), .A2(n6923), .ZN(n12455) );
  NAND2_X1 U14760 ( .A1(n14220), .A2(n12554), .ZN(n12454) );
  NAND2_X1 U14761 ( .A1(n12455), .A2(n12454), .ZN(n12456) );
  XNOR2_X1 U14762 ( .A(n12456), .B(n12522), .ZN(n12458) );
  AND2_X1 U14763 ( .A1(n14220), .A2(n12553), .ZN(n12457) );
  AOI21_X1 U14764 ( .B1(n14343), .B2(n12554), .A(n12457), .ZN(n12459) );
  NAND2_X1 U14765 ( .A1(n12458), .A2(n12459), .ZN(n12464) );
  INV_X1 U14766 ( .A(n12458), .ZN(n12461) );
  INV_X1 U14767 ( .A(n12459), .ZN(n12460) );
  NAND2_X1 U14768 ( .A1(n12461), .A2(n12460), .ZN(n12462) );
  AND2_X1 U14769 ( .A1(n12464), .A2(n12462), .ZN(n13850) );
  NAND2_X1 U14770 ( .A1(n14337), .A2(n6923), .ZN(n12466) );
  NAND2_X1 U14771 ( .A1(n13940), .A2(n12554), .ZN(n12465) );
  NAND2_X1 U14772 ( .A1(n12466), .A2(n12465), .ZN(n12467) );
  XNOR2_X1 U14773 ( .A(n12467), .B(n12551), .ZN(n12477) );
  AOI22_X1 U14774 ( .A1(n14337), .A2(n12554), .B1(n12553), .B2(n13940), .ZN(
        n12475) );
  XNOR2_X1 U14775 ( .A(n12477), .B(n12475), .ZN(n13902) );
  NAND2_X1 U14776 ( .A1(n14332), .A2(n6923), .ZN(n12469) );
  OR2_X1 U14777 ( .A1(n13905), .A2(n12542), .ZN(n12468) );
  NAND2_X1 U14778 ( .A1(n12469), .A2(n12468), .ZN(n12470) );
  XNOR2_X1 U14779 ( .A(n12470), .B(n12522), .ZN(n12474) );
  NOR2_X1 U14780 ( .A1(n13905), .A2(n12525), .ZN(n12471) );
  AOI21_X1 U14781 ( .B1(n14332), .B2(n12554), .A(n12471), .ZN(n12473) );
  OR2_X1 U14782 ( .A1(n12474), .A2(n12473), .ZN(n12472) );
  AND2_X1 U14783 ( .A1(n13902), .A2(n12472), .ZN(n12479) );
  INV_X1 U14784 ( .A(n12472), .ZN(n12478) );
  XNOR2_X1 U14785 ( .A(n12474), .B(n12473), .ZN(n13799) );
  INV_X1 U14786 ( .A(n12475), .ZN(n12476) );
  NOR2_X1 U14787 ( .A1(n12477), .A2(n12476), .ZN(n13800) );
  NOR2_X1 U14788 ( .A1(n13799), .A2(n13800), .ZN(n13802) );
  OAI22_X1 U14789 ( .A1(n14325), .A2(n12545), .B1(n14205), .B2(n12525), .ZN(
        n12481) );
  OAI22_X1 U14790 ( .A1(n14325), .A2(n6907), .B1(n14205), .B2(n12545), .ZN(
        n12480) );
  XNOR2_X1 U14791 ( .A(n12480), .B(n12551), .ZN(n12482) );
  XOR2_X1 U14792 ( .A(n12481), .B(n12482), .Z(n13870) );
  NAND2_X1 U14793 ( .A1(n12482), .A2(n12481), .ZN(n12483) );
  NAND2_X1 U14794 ( .A1(n14319), .A2(n6923), .ZN(n12485) );
  NAND2_X1 U14795 ( .A1(n14183), .A2(n12554), .ZN(n12484) );
  NAND2_X1 U14796 ( .A1(n12485), .A2(n12484), .ZN(n12486) );
  XNOR2_X1 U14797 ( .A(n12486), .B(n12522), .ZN(n12489) );
  AND2_X1 U14798 ( .A1(n14183), .A2(n12553), .ZN(n12487) );
  AOI21_X1 U14799 ( .B1(n14319), .B2(n12554), .A(n12487), .ZN(n12488) );
  NAND2_X1 U14800 ( .A1(n12489), .A2(n12488), .ZN(n13894) );
  OAI21_X1 U14801 ( .B1(n12489), .B2(n12488), .A(n13894), .ZN(n13811) );
  NAND2_X1 U14802 ( .A1(n14314), .A2(n6923), .ZN(n12491) );
  NAND2_X1 U14803 ( .A1(n12554), .A2(n13938), .ZN(n12490) );
  NAND2_X1 U14804 ( .A1(n12491), .A2(n12490), .ZN(n12492) );
  XNOR2_X1 U14805 ( .A(n12492), .B(n12522), .ZN(n12495) );
  INV_X1 U14806 ( .A(n13938), .ZN(n12493) );
  NOR2_X1 U14807 ( .A1(n12525), .A2(n12493), .ZN(n12494) );
  AOI21_X1 U14808 ( .B1(n14314), .B2(n12554), .A(n12494), .ZN(n12496) );
  NAND2_X1 U14809 ( .A1(n12495), .A2(n12496), .ZN(n13787) );
  INV_X1 U14810 ( .A(n12495), .ZN(n12498) );
  INV_X1 U14811 ( .A(n12496), .ZN(n12497) );
  NAND2_X1 U14812 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  AND2_X1 U14813 ( .A1(n13787), .A2(n12499), .ZN(n13892) );
  NAND2_X1 U14814 ( .A1(n13790), .A2(n13787), .ZN(n12510) );
  NAND2_X1 U14815 ( .A1(n14307), .A2(n6923), .ZN(n12502) );
  NAND2_X1 U14816 ( .A1(n12554), .A2(n13937), .ZN(n12501) );
  NAND2_X1 U14817 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  XNOR2_X1 U14818 ( .A(n12503), .B(n12522), .ZN(n12505) );
  NOR2_X1 U14819 ( .A1(n12525), .A2(n13889), .ZN(n12504) );
  AOI21_X1 U14820 ( .B1(n14307), .B2(n12554), .A(n12504), .ZN(n12506) );
  NAND2_X1 U14821 ( .A1(n12505), .A2(n12506), .ZN(n13861) );
  INV_X1 U14822 ( .A(n12505), .ZN(n12508) );
  INV_X1 U14823 ( .A(n12506), .ZN(n12507) );
  NAND2_X1 U14824 ( .A1(n12508), .A2(n12507), .ZN(n12509) );
  NAND2_X1 U14825 ( .A1(n14301), .A2(n6923), .ZN(n12512) );
  NAND2_X1 U14826 ( .A1(n12554), .A2(n13936), .ZN(n12511) );
  NAND2_X1 U14827 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  XNOR2_X1 U14828 ( .A(n12513), .B(n12522), .ZN(n12515) );
  INV_X1 U14829 ( .A(n13936), .ZN(n13829) );
  NOR2_X1 U14830 ( .A1(n12525), .A2(n13829), .ZN(n12514) );
  AOI21_X1 U14831 ( .B1(n14301), .B2(n12554), .A(n12514), .ZN(n12516) );
  NAND2_X1 U14832 ( .A1(n12515), .A2(n12516), .ZN(n13834) );
  INV_X1 U14833 ( .A(n12515), .ZN(n12518) );
  INV_X1 U14834 ( .A(n12516), .ZN(n12517) );
  NAND2_X1 U14835 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U14836 ( .A1(n14293), .A2(n6923), .ZN(n12521) );
  NAND2_X1 U14837 ( .A1(n12554), .A2(n13935), .ZN(n12520) );
  NAND2_X1 U14838 ( .A1(n12521), .A2(n12520), .ZN(n12523) );
  XNOR2_X1 U14839 ( .A(n12523), .B(n12522), .ZN(n12527) );
  INV_X1 U14840 ( .A(n13935), .ZN(n12524) );
  NOR2_X1 U14841 ( .A1(n12525), .A2(n12524), .ZN(n12526) );
  AOI21_X1 U14842 ( .B1(n14293), .B2(n12554), .A(n12526), .ZN(n12528) );
  NAND2_X1 U14843 ( .A1(n12527), .A2(n12528), .ZN(n12532) );
  INV_X1 U14844 ( .A(n12527), .ZN(n12530) );
  INV_X1 U14845 ( .A(n12528), .ZN(n12529) );
  NAND2_X1 U14846 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  NAND2_X1 U14847 ( .A1(n13836), .A2(n12532), .ZN(n13911) );
  NAND2_X1 U14848 ( .A1(n14289), .A2(n6923), .ZN(n12534) );
  NAND2_X1 U14849 ( .A1(n12554), .A2(n13934), .ZN(n12533) );
  NAND2_X1 U14850 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  XNOR2_X1 U14851 ( .A(n12535), .B(n12551), .ZN(n12539) );
  NAND2_X1 U14852 ( .A1(n14289), .A2(n12554), .ZN(n12537) );
  NAND2_X1 U14853 ( .A1(n12553), .A2(n13934), .ZN(n12536) );
  NAND2_X1 U14854 ( .A1(n12537), .A2(n12536), .ZN(n12538) );
  NOR2_X1 U14855 ( .A1(n12539), .A2(n12538), .ZN(n12540) );
  AOI21_X1 U14856 ( .B1(n12539), .B2(n12538), .A(n12540), .ZN(n13912) );
  INV_X1 U14857 ( .A(n12540), .ZN(n12541) );
  OAI22_X1 U14858 ( .A1(n14055), .A2(n6907), .B1(n14042), .B2(n12542), .ZN(
        n12544) );
  XNOR2_X1 U14859 ( .A(n12544), .B(n12551), .ZN(n12549) );
  OR2_X1 U14860 ( .A1(n14055), .A2(n12545), .ZN(n12547) );
  NAND2_X1 U14861 ( .A1(n12553), .A2(n14068), .ZN(n12546) );
  NAND2_X1 U14862 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  NOR2_X1 U14863 ( .A1(n12549), .A2(n12548), .ZN(n12550) );
  AOI22_X1 U14864 ( .A1(n14280), .A2(n6923), .B1(n12554), .B2(n14058), .ZN(
        n12552) );
  XNOR2_X1 U14865 ( .A(n12552), .B(n12551), .ZN(n12556) );
  AOI22_X1 U14866 ( .A1(n14280), .A2(n12554), .B1(n12553), .B2(n14058), .ZN(
        n12555) );
  XNOR2_X1 U14867 ( .A(n12556), .B(n12555), .ZN(n12557) );
  AOI22_X1 U14868 ( .A1(n8890), .A2(n14068), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12560) );
  NAND2_X1 U14869 ( .A1(n12558), .A2(n14069), .ZN(n12559) );
  OAI211_X1 U14870 ( .C1(n14620), .C2(n14078), .A(n12560), .B(n12559), .ZN(
        n12561) );
  AOI21_X1 U14871 ( .B1(n14280), .B2(n14616), .A(n12561), .ZN(n12562) );
  OAI21_X1 U14872 ( .B1(n12563), .B2(n13932), .A(n12562), .ZN(P1_U3220) );
  INV_X1 U14873 ( .A(n12564), .ZN(n12566) );
  OAI222_X1 U14874 ( .A1(P3_U3151), .A2(n12777), .B1(n13120), .B2(n12566), 
        .C1(n12565), .C2(n13122), .ZN(P3_U3268) );
  INV_X1 U14875 ( .A(n12567), .ZN(n12568) );
  OAI222_X1 U14876 ( .A1(n13122), .A2(n12570), .B1(P3_U3151), .B2(n12569), 
        .C1(n13120), .C2(n12568), .ZN(P3_U3265) );
  XNOR2_X1 U14877 ( .A(n12572), .B(n12571), .ZN(n12573) );
  NAND2_X1 U14878 ( .A1(n12573), .A2(n12651), .ZN(n12578) );
  AOI22_X1 U14879 ( .A1(n12855), .A2(n12643), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12574) );
  OAI21_X1 U14880 ( .B1(n12575), .B2(n12646), .A(n12574), .ZN(n12576) );
  AOI21_X1 U14881 ( .B1(n12830), .B2(n12670), .A(n12576), .ZN(n12577) );
  OAI211_X1 U14882 ( .C1(n12579), .C2(n12666), .A(n12578), .B(n12577), .ZN(
        P3_U3154) );
  XNOR2_X1 U14883 ( .A(n12580), .B(n12899), .ZN(n12585) );
  NAND2_X1 U14884 ( .A1(n12670), .A2(n12890), .ZN(n12582) );
  AOI22_X1 U14885 ( .A1(n12854), .A2(n12663), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12581) );
  OAI211_X1 U14886 ( .C1(n12883), .C2(n12665), .A(n12582), .B(n12581), .ZN(
        n12583) );
  AOI21_X1 U14887 ( .B1(n13012), .B2(n12648), .A(n12583), .ZN(n12584) );
  OAI21_X1 U14888 ( .B1(n12585), .B2(n12672), .A(n12584), .ZN(P3_U3156) );
  OAI211_X1 U14889 ( .C1(n12588), .C2(n12587), .A(n12586), .B(n12651), .ZN(
        n12592) );
  NAND2_X1 U14890 ( .A1(n12677), .A2(n12643), .ZN(n12589) );
  NAND2_X1 U14891 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12793)
         );
  OAI211_X1 U14892 ( .C1(n12936), .C2(n12646), .A(n12589), .B(n12793), .ZN(
        n12590) );
  AOI21_X1 U14893 ( .B1(n12941), .B2(n12670), .A(n12590), .ZN(n12591) );
  OAI211_X1 U14894 ( .C1(n12666), .C2(n12940), .A(n12592), .B(n12591), .ZN(
        P3_U3159) );
  INV_X1 U14895 ( .A(n12593), .ZN(n12594) );
  AOI21_X1 U14896 ( .B1(n12596), .B2(n12595), .A(n12594), .ZN(n12601) );
  AOI22_X1 U14897 ( .A1(n12908), .A2(n12643), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12598) );
  NAND2_X1 U14898 ( .A1(n12670), .A2(n12912), .ZN(n12597) );
  OAI211_X1 U14899 ( .C1(n12883), .C2(n12646), .A(n12598), .B(n12597), .ZN(
        n12599) );
  AOI21_X1 U14900 ( .B1(n13079), .B2(n12648), .A(n12599), .ZN(n12600) );
  OAI21_X1 U14901 ( .B1(n12601), .B2(n12672), .A(n12600), .ZN(P3_U3163) );
  XOR2_X1 U14902 ( .A(n12603), .B(n12602), .Z(n12608) );
  NAND2_X1 U14903 ( .A1(n12670), .A2(n12859), .ZN(n12605) );
  AOI22_X1 U14904 ( .A1(n12855), .A2(n12663), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12604) );
  OAI211_X1 U14905 ( .C1(n12882), .C2(n12665), .A(n12605), .B(n12604), .ZN(
        n12606) );
  AOI21_X1 U14906 ( .B1(n13060), .B2(n12648), .A(n12606), .ZN(n12607) );
  OAI21_X1 U14907 ( .B1(n12608), .B2(n12672), .A(n12607), .ZN(P3_U3165) );
  INV_X1 U14908 ( .A(n13037), .ZN(n12617) );
  OAI211_X1 U14909 ( .C1(n12611), .C2(n12610), .A(n12609), .B(n12651), .ZN(
        n12616) );
  NAND2_X1 U14910 ( .A1(n12678), .A2(n12643), .ZN(n12612) );
  NAND2_X1 U14911 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12758)
         );
  OAI211_X1 U14912 ( .C1(n12656), .C2(n12646), .A(n12612), .B(n12758), .ZN(
        n12613) );
  AOI21_X1 U14913 ( .B1(n12614), .B2(n12670), .A(n12613), .ZN(n12615) );
  OAI211_X1 U14914 ( .C1(n12617), .C2(n12666), .A(n12616), .B(n12615), .ZN(
        P3_U3166) );
  INV_X1 U14915 ( .A(n13033), .ZN(n12626) );
  OAI211_X1 U14916 ( .C1(n12620), .C2(n12619), .A(n12618), .B(n12651), .ZN(
        n12625) );
  NAND2_X1 U14917 ( .A1(n12621), .A2(n12643), .ZN(n12622) );
  NAND2_X1 U14918 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14530)
         );
  OAI211_X1 U14919 ( .C1(n12962), .C2(n12646), .A(n12622), .B(n14530), .ZN(
        n12623) );
  AOI21_X1 U14920 ( .B1(n12963), .B2(n12670), .A(n12623), .ZN(n12624) );
  OAI211_X1 U14921 ( .C1(n12626), .C2(n12666), .A(n12625), .B(n12624), .ZN(
        P3_U3168) );
  XOR2_X1 U14922 ( .A(n12628), .B(n12627), .Z(n12633) );
  AOI22_X1 U14923 ( .A1(n12838), .A2(n12663), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12630) );
  NAND2_X1 U14924 ( .A1(n12670), .A2(n12873), .ZN(n12629) );
  OAI211_X1 U14925 ( .C1(n12872), .C2(n12665), .A(n12630), .B(n12629), .ZN(
        n12631) );
  AOI21_X1 U14926 ( .B1(n13008), .B2(n12648), .A(n12631), .ZN(n12632) );
  OAI21_X1 U14927 ( .B1(n12633), .B2(n12672), .A(n12632), .ZN(P3_U3169) );
  INV_X1 U14928 ( .A(n13022), .ZN(n12641) );
  OAI211_X1 U14929 ( .C1(n12636), .C2(n12635), .A(n12634), .B(n12651), .ZN(
        n12640) );
  AOI22_X1 U14930 ( .A1(n12898), .A2(n12663), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12637) );
  OAI21_X1 U14931 ( .B1(n12917), .B2(n12665), .A(n12637), .ZN(n12638) );
  AOI21_X1 U14932 ( .B1(n12923), .B2(n12670), .A(n12638), .ZN(n12639) );
  OAI211_X1 U14933 ( .C1(n12641), .C2(n12666), .A(n12640), .B(n12639), .ZN(
        P3_U3173) );
  XNOR2_X1 U14934 ( .A(n12642), .B(n12909), .ZN(n12650) );
  NAND2_X1 U14935 ( .A1(n12670), .A2(n12902), .ZN(n12645) );
  AOI22_X1 U14936 ( .A1(n12898), .A2(n12643), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12644) );
  OAI211_X1 U14937 ( .C1(n12872), .C2(n12646), .A(n12645), .B(n12644), .ZN(
        n12647) );
  AOI21_X1 U14938 ( .B1(n13073), .B2(n12648), .A(n12647), .ZN(n12649) );
  OAI21_X1 U14939 ( .B1(n12650), .B2(n12672), .A(n12649), .ZN(P3_U3175) );
  INV_X1 U14940 ( .A(n13096), .ZN(n12660) );
  OAI211_X1 U14941 ( .C1(n12654), .C2(n12653), .A(n12652), .B(n12651), .ZN(
        n12659) );
  AND2_X1 U14942 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14553) );
  AOI21_X1 U14943 ( .B1(n12952), .B2(n12663), .A(n14553), .ZN(n12655) );
  OAI21_X1 U14944 ( .B1(n12656), .B2(n12665), .A(n12655), .ZN(n12657) );
  AOI21_X1 U14945 ( .B1(n12954), .B2(n12670), .A(n12657), .ZN(n12658) );
  OAI211_X1 U14946 ( .C1(n12660), .C2(n12666), .A(n12659), .B(n12658), .ZN(
        P3_U3178) );
  XOR2_X1 U14947 ( .A(n12662), .B(n12661), .Z(n12673) );
  AOI22_X1 U14948 ( .A1(n12837), .A2(n12663), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12664) );
  OAI21_X1 U14949 ( .B1(n12871), .B2(n12665), .A(n12664), .ZN(n12669) );
  NOR2_X1 U14950 ( .A1(n12667), .A2(n12666), .ZN(n12668) );
  AOI211_X1 U14951 ( .C1(n12842), .C2(n12670), .A(n12669), .B(n12668), .ZN(
        n12671) );
  OAI21_X1 U14952 ( .B1(n12673), .B2(n12672), .A(n12671), .ZN(P3_U3180) );
  MUX2_X1 U14953 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12674), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14954 ( .A(n12675), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12686), .Z(
        P3_U3521) );
  MUX2_X1 U14955 ( .A(n12676), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12686), .Z(
        P3_U3520) );
  MUX2_X1 U14956 ( .A(n12855), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12686), .Z(
        P3_U3517) );
  MUX2_X1 U14957 ( .A(n12838), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12686), .Z(
        P3_U3516) );
  MUX2_X1 U14958 ( .A(n12854), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12686), .Z(
        P3_U3515) );
  MUX2_X1 U14959 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12899), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14960 ( .A(n12909), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12686), .Z(
        P3_U3513) );
  MUX2_X1 U14961 ( .A(n12898), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12686), .Z(
        P3_U3512) );
  MUX2_X1 U14962 ( .A(n12908), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12686), .Z(
        P3_U3511) );
  MUX2_X1 U14963 ( .A(n12952), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12686), .Z(
        P3_U3510) );
  MUX2_X1 U14964 ( .A(n12677), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12686), .Z(
        P3_U3509) );
  MUX2_X1 U14965 ( .A(n12951), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12686), .Z(
        P3_U3508) );
  MUX2_X1 U14966 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12678), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14967 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14564), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14968 ( .A(n12975), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12686), .Z(
        P3_U3504) );
  MUX2_X1 U14969 ( .A(n14563), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12686), .Z(
        P3_U3503) );
  MUX2_X1 U14970 ( .A(n15000), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12686), .Z(
        P3_U3502) );
  MUX2_X1 U14971 ( .A(n15001), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12686), .Z(
        P3_U3500) );
  MUX2_X1 U14972 ( .A(n12679), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12686), .Z(
        P3_U3499) );
  MUX2_X1 U14973 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12680), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14974 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12681), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14975 ( .A(n12682), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12686), .Z(
        P3_U3496) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12683), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14977 ( .A(n6954), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12686), .Z(
        P3_U3494) );
  MUX2_X1 U14978 ( .A(n12685), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12686), .Z(
        P3_U3492) );
  MUX2_X1 U14979 ( .A(n15063), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12686), .Z(
        P3_U3491) );
  NOR2_X1 U14980 ( .A1(n12707), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U14981 ( .A1(n12690), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12729) );
  OAI21_X1 U14982 ( .B1(n12690), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12729), 
        .ZN(n12709) );
  AOI21_X1 U14983 ( .B1(n12691), .B2(n12709), .A(n12720), .ZN(n12719) );
  NAND2_X1 U14984 ( .A1(n12693), .A2(n12692), .ZN(n12695) );
  OR2_X1 U14985 ( .A1(n12699), .A2(n12696), .ZN(n12728) );
  NAND2_X1 U14986 ( .A1(n12699), .A2(n12696), .ZN(n12697) );
  AND2_X1 U14987 ( .A1(n12728), .A2(n12697), .ZN(n12712) );
  OAI21_X1 U14988 ( .B1(n12698), .B2(n12712), .A(n12724), .ZN(n12705) );
  INV_X1 U14989 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12703) );
  INV_X1 U14990 ( .A(n14987), .ZN(n14532) );
  NAND2_X1 U14991 ( .A1(n14543), .A2(n12699), .ZN(n12702) );
  INV_X1 U14992 ( .A(n12700), .ZN(n12701) );
  OAI211_X1 U14993 ( .C1(n12703), .C2(n14532), .A(n12702), .B(n12701), .ZN(
        n12704) );
  AOI21_X1 U14994 ( .B1(n12705), .B2(n14990), .A(n12704), .ZN(n12718) );
  INV_X1 U14995 ( .A(n12706), .ZN(n12708) );
  NAND2_X1 U14996 ( .A1(n12708), .A2(n12707), .ZN(n12713) );
  AND2_X1 U14997 ( .A1(n12714), .A2(n12713), .ZN(n12716) );
  INV_X1 U14998 ( .A(n12709), .ZN(n12711) );
  MUX2_X1 U14999 ( .A(n12712), .B(n12711), .S(n12710), .Z(n12715) );
  NAND3_X1 U15000 ( .A1(n12714), .A2(n12715), .A3(n12713), .ZN(n12731) );
  OAI211_X1 U15001 ( .C1(n12716), .C2(n12715), .A(n12795), .B(n12731), .ZN(
        n12717) );
  OAI211_X1 U15002 ( .C1(n12719), .C2(n14994), .A(n12718), .B(n12717), .ZN(
        P3_U3196) );
  INV_X1 U15003 ( .A(n12720), .ZN(n12721) );
  NAND2_X1 U15004 ( .A1(n12729), .A2(n12721), .ZN(n12748) );
  AOI21_X1 U15005 ( .B1(n12723), .B2(n12722), .A(n12749), .ZN(n12739) );
  NAND2_X1 U15006 ( .A1(n12728), .A2(n12724), .ZN(n12754) );
  XOR2_X1 U15007 ( .A(n12755), .B(n12754), .Z(n12725) );
  OAI21_X1 U15008 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12725), .A(n12756), 
        .ZN(n12737) );
  INV_X1 U15009 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U15010 ( .A1(n14543), .A2(n12742), .ZN(n12727) );
  OAI211_X1 U15011 ( .C1(n14409), .C2(n14532), .A(n12727), .B(n12726), .ZN(
        n12736) );
  MUX2_X1 U15012 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12777), .Z(n12733) );
  MUX2_X1 U15013 ( .A(n12729), .B(n12728), .S(n12777), .Z(n12730) );
  NAND2_X1 U15014 ( .A1(n12731), .A2(n12730), .ZN(n12740) );
  XNOR2_X1 U15015 ( .A(n12740), .B(n12755), .ZN(n12732) );
  NOR2_X1 U15016 ( .A1(n12732), .A2(n12733), .ZN(n12741) );
  AOI21_X1 U15017 ( .B1(n12733), .B2(n12732), .A(n12741), .ZN(n12734) );
  NOR2_X1 U15018 ( .A1(n12734), .A2(n14983), .ZN(n12735) );
  AOI211_X1 U15019 ( .C1(n14990), .C2(n12737), .A(n12736), .B(n12735), .ZN(
        n12738) );
  OAI21_X1 U15020 ( .B1(n12739), .B2(n14994), .A(n12738), .ZN(P3_U3197) );
  INV_X1 U15021 ( .A(n12740), .ZN(n12743) );
  AOI21_X1 U15022 ( .B1(n12743), .B2(n12742), .A(n12741), .ZN(n12775) );
  INV_X1 U15023 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13038) );
  MUX2_X1 U15024 ( .A(n12751), .B(n13038), .S(n12777), .Z(n12745) );
  NOR2_X1 U15025 ( .A1(n12745), .A2(n12744), .ZN(n12774) );
  NAND2_X1 U15026 ( .A1(n12745), .A2(n12744), .ZN(n12773) );
  INV_X1 U15027 ( .A(n12773), .ZN(n12746) );
  NOR2_X1 U15028 ( .A1(n12774), .A2(n12746), .ZN(n12747) );
  XNOR2_X1 U15029 ( .A(n12775), .B(n12747), .ZN(n12764) );
  NAND2_X1 U15030 ( .A1(n12782), .A2(n12751), .ZN(n12750) );
  OAI21_X1 U15031 ( .B1(n12782), .B2(n12751), .A(n12750), .ZN(n12752) );
  OAI21_X1 U15032 ( .B1(n7510), .B2(n12752), .A(n12766), .ZN(n12753) );
  NAND2_X1 U15033 ( .A1(n12753), .A2(n14554), .ZN(n12763) );
  NAND2_X1 U15034 ( .A1(n12755), .A2(n12754), .ZN(n12757) );
  XNOR2_X1 U15035 ( .A(n12782), .B(n13038), .ZN(n12783) );
  XNOR2_X1 U15036 ( .A(n12784), .B(n12783), .ZN(n12761) );
  NOR2_X1 U15037 ( .A1(n14981), .A2(n12782), .ZN(n12760) );
  INV_X1 U15038 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U15039 ( .B1(n14532), .B2(n14377), .A(n12758), .ZN(n12759) );
  AOI211_X1 U15040 ( .C1(n12761), .C2(n14990), .A(n12760), .B(n12759), .ZN(
        n12762) );
  OAI211_X1 U15041 ( .C1(n14983), .C2(n12764), .A(n12763), .B(n12762), .ZN(
        P3_U3198) );
  NAND2_X1 U15042 ( .A1(n12782), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12765) );
  NOR2_X1 U15043 ( .A1(n14529), .A2(n12767), .ZN(n12768) );
  INV_X1 U15044 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14526) );
  INV_X1 U15045 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15046 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14542), .B1(n12781), 
        .B2(n12769), .ZN(n14555) );
  NOR2_X1 U15047 ( .A1(n14556), .A2(n14555), .ZN(n14557) );
  AOI21_X1 U15048 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n12781), .A(n14557), 
        .ZN(n12770) );
  XNOR2_X1 U15049 ( .A(n12771), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12772) );
  XNOR2_X1 U15050 ( .A(n12770), .B(n12772), .ZN(n12798) );
  XNOR2_X1 U15051 ( .A(n12771), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12789) );
  MUX2_X1 U15052 ( .A(n12772), .B(n12789), .S(n12777), .Z(n12780) );
  MUX2_X1 U15053 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12777), .Z(n12776) );
  OAI21_X1 U15054 ( .B1(n12775), .B2(n12774), .A(n12773), .ZN(n14535) );
  XNOR2_X1 U15055 ( .A(n12776), .B(n12786), .ZN(n14536) );
  NOR2_X1 U15056 ( .A1(n14535), .A2(n14536), .ZN(n14534) );
  AOI21_X1 U15057 ( .B1(n12776), .B2(n12786), .A(n14534), .ZN(n12778) );
  XNOR2_X1 U15058 ( .A(n12778), .B(n14542), .ZN(n14548) );
  MUX2_X1 U15059 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12777), .Z(n14549) );
  NOR2_X1 U15060 ( .A1(n14548), .A2(n14549), .ZN(n14547) );
  AOI21_X1 U15061 ( .B1(n12778), .B2(n14542), .A(n14547), .ZN(n12779) );
  XOR2_X1 U15062 ( .A(n12780), .B(n12779), .Z(n12796) );
  INV_X1 U15063 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U15064 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12781), .B1(n14542), 
        .B2(n13028), .ZN(n14546) );
  INV_X1 U15065 ( .A(n12787), .ZN(n12785) );
  NAND2_X1 U15066 ( .A1(n12786), .A2(n12785), .ZN(n12788) );
  INV_X1 U15067 ( .A(n12789), .ZN(n12790) );
  NAND2_X1 U15068 ( .A1(n14987), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12792) );
  OAI211_X1 U15069 ( .C1(n14981), .C2(n12023), .A(n12793), .B(n12792), .ZN(
        n12794) );
  OAI21_X1 U15070 ( .B1(n12798), .B2(n14994), .A(n12797), .ZN(P3_U3201) );
  INV_X1 U15071 ( .A(n15038), .ZN(n12816) );
  NAND2_X1 U15072 ( .A1(n12799), .A2(n15075), .ZN(n12803) );
  INV_X1 U15073 ( .A(n12800), .ZN(n12801) );
  OR2_X1 U15074 ( .A1(n12802), .A2(n12801), .ZN(n13041) );
  AOI21_X1 U15075 ( .B1(n12803), .B2(n13041), .A(n15083), .ZN(n12805) );
  AOI21_X1 U15076 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15083), .A(n12805), 
        .ZN(n12804) );
  OAI21_X1 U15077 ( .B1(n13043), .B2(n12816), .A(n12804), .ZN(P3_U3202) );
  AOI21_X1 U15078 ( .B1(n15083), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12805), 
        .ZN(n12806) );
  OAI21_X1 U15079 ( .B1(n13046), .B2(n12816), .A(n12806), .ZN(P3_U3203) );
  INV_X1 U15080 ( .A(n12992), .ZN(n12819) );
  NOR2_X1 U15081 ( .A1(n12821), .A2(n12811), .ZN(n12813) );
  XNOR2_X1 U15082 ( .A(n12813), .B(n12812), .ZN(n12993) );
  INV_X1 U15083 ( .A(n12968), .ZN(n14570) );
  AOI22_X1 U15084 ( .A1(n15083), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15075), 
        .B2(n12814), .ZN(n12815) );
  OAI21_X1 U15085 ( .B1(n13050), .B2(n12816), .A(n12815), .ZN(n12817) );
  AOI21_X1 U15086 ( .B1(n12993), .B2(n14570), .A(n12817), .ZN(n12818) );
  OAI21_X1 U15087 ( .B1(n12819), .B2(n15083), .A(n12818), .ZN(P3_U3205) );
  INV_X1 U15088 ( .A(n12820), .ZN(n12823) );
  INV_X1 U15089 ( .A(n12826), .ZN(n12822) );
  AOI21_X1 U15090 ( .B1(n12826), .B2(n12825), .A(n12824), .ZN(n12827) );
  INV_X1 U15091 ( .A(n12827), .ZN(n12829) );
  MUX2_X1 U15092 ( .A(n15240), .B(n13051), .S(n15080), .Z(n12832) );
  AOI22_X1 U15093 ( .A1(n13053), .A2(n15038), .B1(n15075), .B2(n12830), .ZN(
        n12831) );
  OAI211_X1 U15094 ( .C1(n13056), .C2(n12968), .A(n12832), .B(n12831), .ZN(
        P3_U3206) );
  XNOR2_X1 U15095 ( .A(n12834), .B(n12833), .ZN(n13001) );
  XNOR2_X1 U15096 ( .A(n12836), .B(n12835), .ZN(n12840) );
  AOI22_X1 U15097 ( .A1(n12838), .A2(n15062), .B1(n12837), .B2(n15065), .ZN(
        n12839) );
  OAI21_X1 U15098 ( .B1(n12840), .B2(n15053), .A(n12839), .ZN(n12841) );
  AOI21_X1 U15099 ( .B1(n13001), .B2(n15050), .A(n12841), .ZN(n13003) );
  NAND2_X1 U15100 ( .A1(n13000), .A2(n15038), .ZN(n12844) );
  AOI22_X1 U15101 ( .A1(n15083), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15075), 
        .B2(n12842), .ZN(n12843) );
  NAND2_X1 U15102 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  AOI21_X1 U15103 ( .B1(n13001), .B2(n12846), .A(n12845), .ZN(n12847) );
  OAI21_X1 U15104 ( .B1(n13003), .B2(n15083), .A(n12847), .ZN(P3_U3207) );
  XNOR2_X1 U15105 ( .A(n12849), .B(n12848), .ZN(n13063) );
  INV_X1 U15106 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12858) );
  NAND2_X1 U15107 ( .A1(n12851), .A2(n12850), .ZN(n12852) );
  NAND2_X1 U15108 ( .A1(n12852), .A2(n15068), .ZN(n12853) );
  OR2_X1 U15109 ( .A1(n6652), .A2(n12853), .ZN(n12857) );
  AOI22_X1 U15110 ( .A1(n15065), .A2(n12855), .B1(n12854), .B2(n15062), .ZN(
        n12856) );
  MUX2_X1 U15111 ( .A(n12858), .B(n13058), .S(n15080), .Z(n12861) );
  AOI22_X1 U15112 ( .A1(n13060), .A2(n15038), .B1(n15075), .B2(n12859), .ZN(
        n12860) );
  OAI211_X1 U15113 ( .C1(n13063), .C2(n12968), .A(n12861), .B(n12860), .ZN(
        P3_U3208) );
  NAND2_X1 U15114 ( .A1(n12885), .A2(n12862), .ZN(n12864) );
  AND2_X1 U15115 ( .A1(n12864), .A2(n12863), .ZN(n12867) );
  INV_X1 U15116 ( .A(n12865), .ZN(n12866) );
  AOI21_X1 U15117 ( .B1(n12867), .B2(n12868), .A(n12866), .ZN(n13067) );
  XNOR2_X1 U15118 ( .A(n12869), .B(n12868), .ZN(n12870) );
  OAI222_X1 U15119 ( .A1(n15048), .A2(n12872), .B1(n15046), .B2(n12871), .C1(
        n12870), .C2(n15053), .ZN(n13007) );
  NAND2_X1 U15120 ( .A1(n13007), .A2(n15080), .ZN(n12878) );
  INV_X1 U15121 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12875) );
  INV_X1 U15122 ( .A(n12873), .ZN(n12874) );
  OAI22_X1 U15123 ( .A1(n15080), .A2(n12875), .B1(n12874), .B2(n15040), .ZN(
        n12876) );
  AOI21_X1 U15124 ( .B1(n13008), .B2(n15038), .A(n12876), .ZN(n12877) );
  OAI211_X1 U15125 ( .C1(n13067), .C2(n12968), .A(n12878), .B(n12877), .ZN(
        P3_U3209) );
  XNOR2_X1 U15126 ( .A(n12880), .B(n12879), .ZN(n12881) );
  OAI222_X1 U15127 ( .A1(n15048), .A2(n12883), .B1(n15046), .B2(n12882), .C1(
        n15053), .C2(n12881), .ZN(n13011) );
  NAND2_X1 U15128 ( .A1(n12885), .A2(n12884), .ZN(n12887) );
  NAND2_X1 U15129 ( .A1(n12887), .A2(n12886), .ZN(n12889) );
  OR2_X1 U15130 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  NAND2_X1 U15131 ( .A1(n12889), .A2(n12888), .ZN(n13071) );
  AOI22_X1 U15132 ( .A1(n15083), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15075), 
        .B2(n12890), .ZN(n12892) );
  NAND2_X1 U15133 ( .A1(n13012), .A2(n15038), .ZN(n12891) );
  OAI211_X1 U15134 ( .C1(n13071), .C2(n12968), .A(n12892), .B(n12891), .ZN(
        n12893) );
  AOI21_X1 U15135 ( .B1(n13011), .B2(n15080), .A(n12893), .ZN(n12894) );
  INV_X1 U15136 ( .A(n12894), .ZN(P3_U3210) );
  XOR2_X1 U15137 ( .A(n12896), .B(n12895), .Z(n13076) );
  INV_X1 U15138 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12901) );
  XNOR2_X1 U15139 ( .A(n12897), .B(n12896), .ZN(n12900) );
  AOI222_X1 U15140 ( .A1(n15068), .A2(n12900), .B1(n12899), .B2(n15065), .C1(
        n12898), .C2(n15062), .ZN(n13072) );
  MUX2_X1 U15141 ( .A(n12901), .B(n13072), .S(n15080), .Z(n12904) );
  AOI22_X1 U15142 ( .A1(n13073), .A2(n15038), .B1(n15075), .B2(n12902), .ZN(
        n12903) );
  OAI211_X1 U15143 ( .C1(n13076), .C2(n12968), .A(n12904), .B(n12903), .ZN(
        P3_U3211) );
  XOR2_X1 U15144 ( .A(n12905), .B(n12907), .Z(n13082) );
  INV_X1 U15145 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12911) );
  XOR2_X1 U15146 ( .A(n12906), .B(n12907), .Z(n12910) );
  AOI222_X1 U15147 ( .A1(n15068), .A2(n12910), .B1(n12909), .B2(n15065), .C1(
        n12908), .C2(n15062), .ZN(n13077) );
  MUX2_X1 U15148 ( .A(n12911), .B(n13077), .S(n15080), .Z(n12914) );
  AOI22_X1 U15149 ( .A1(n13079), .A2(n15038), .B1(n15075), .B2(n12912), .ZN(
        n12913) );
  OAI211_X1 U15150 ( .C1(n13082), .C2(n12968), .A(n12914), .B(n12913), .ZN(
        P3_U3212) );
  XNOR2_X1 U15151 ( .A(n12915), .B(n12919), .ZN(n12916) );
  OAI222_X1 U15152 ( .A1(n15046), .A2(n12918), .B1(n15048), .B2(n12917), .C1(
        n15053), .C2(n12916), .ZN(n13021) );
  NAND2_X1 U15153 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  NAND2_X1 U15154 ( .A1(n12922), .A2(n12921), .ZN(n13086) );
  AOI22_X1 U15155 ( .A1(n15083), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15075), 
        .B2(n12923), .ZN(n12925) );
  NAND2_X1 U15156 ( .A1(n13022), .A2(n15038), .ZN(n12924) );
  OAI211_X1 U15157 ( .C1(n13086), .C2(n12968), .A(n12925), .B(n12924), .ZN(
        n12926) );
  AOI21_X1 U15158 ( .B1(n13021), .B2(n15080), .A(n12926), .ZN(n12927) );
  INV_X1 U15159 ( .A(n12927), .ZN(P3_U3213) );
  NAND2_X1 U15160 ( .A1(n12945), .A2(n12928), .ZN(n12930) );
  XNOR2_X1 U15161 ( .A(n12930), .B(n12929), .ZN(n13092) );
  INV_X1 U15162 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12939) );
  INV_X1 U15163 ( .A(n12931), .ZN(n12935) );
  AOI21_X1 U15164 ( .B1(n12948), .B2(n12933), .A(n12932), .ZN(n12934) );
  NOR3_X1 U15165 ( .A1(n12935), .A2(n12934), .A3(n15053), .ZN(n12938) );
  OAI22_X1 U15166 ( .A1(n12962), .A2(n15048), .B1(n12936), .B2(n15046), .ZN(
        n12937) );
  NOR2_X1 U15167 ( .A1(n12938), .A2(n12937), .ZN(n13087) );
  MUX2_X1 U15168 ( .A(n12939), .B(n13087), .S(n15080), .Z(n12943) );
  INV_X1 U15169 ( .A(n12940), .ZN(n13089) );
  AOI22_X1 U15170 ( .A1(n13089), .A2(n15038), .B1(n15075), .B2(n12941), .ZN(
        n12942) );
  OAI211_X1 U15171 ( .C1(n13092), .C2(n12968), .A(n12943), .B(n12942), .ZN(
        P3_U3214) );
  INV_X1 U15172 ( .A(n12944), .ZN(n12947) );
  OAI21_X1 U15173 ( .B1(n12947), .B2(n12946), .A(n12945), .ZN(n13099) );
  OAI21_X1 U15174 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(n12953) );
  AOI222_X1 U15175 ( .A1(n15068), .A2(n12953), .B1(n12952), .B2(n15065), .C1(
        n12951), .C2(n15062), .ZN(n13093) );
  MUX2_X1 U15176 ( .A(n12769), .B(n13093), .S(n15080), .Z(n12956) );
  AOI22_X1 U15177 ( .A1(n13096), .A2(n15038), .B1(n15075), .B2(n12954), .ZN(
        n12955) );
  OAI211_X1 U15178 ( .C1(n13099), .C2(n12968), .A(n12956), .B(n12955), .ZN(
        P3_U3215) );
  XNOR2_X1 U15179 ( .A(n12957), .B(n12958), .ZN(n13103) );
  XNOR2_X1 U15180 ( .A(n12959), .B(n12958), .ZN(n12960) );
  OAI222_X1 U15181 ( .A1(n15046), .A2(n12962), .B1(n15048), .B2(n12961), .C1(
        n12960), .C2(n15053), .ZN(n13032) );
  NAND2_X1 U15182 ( .A1(n13032), .A2(n15080), .ZN(n12967) );
  INV_X1 U15183 ( .A(n12963), .ZN(n12964) );
  OAI22_X1 U15184 ( .A1(n15080), .A2(n14526), .B1(n12964), .B2(n15040), .ZN(
        n12965) );
  AOI21_X1 U15185 ( .B1(n13033), .B2(n15038), .A(n12965), .ZN(n12966) );
  OAI211_X1 U15186 ( .C1(n13103), .C2(n12968), .A(n12967), .B(n12966), .ZN(
        P3_U3216) );
  NAND2_X1 U15187 ( .A1(n15018), .A2(n15015), .ZN(n14575) );
  NAND2_X1 U15188 ( .A1(n14575), .A2(n12969), .ZN(n12971) );
  NAND2_X1 U15189 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  NAND2_X1 U15190 ( .A1(n12972), .A2(n12979), .ZN(n12973) );
  NAND3_X1 U15191 ( .A1(n12974), .A2(n15068), .A3(n12973), .ZN(n12977) );
  AOI22_X1 U15192 ( .A1(n15062), .A2(n15000), .B1(n12975), .B2(n15065), .ZN(
        n12976) );
  NAND2_X1 U15193 ( .A1(n12977), .A2(n12976), .ZN(n14596) );
  NAND2_X1 U15194 ( .A1(n14596), .A2(n15080), .ZN(n12985) );
  AOI22_X1 U15195 ( .A1(n15083), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15075), 
        .B2(n12978), .ZN(n12984) );
  XNOR2_X1 U15196 ( .A(n12980), .B(n12979), .ZN(n14593) );
  NAND2_X1 U15197 ( .A1(n14593), .A2(n14570), .ZN(n12983) );
  AND2_X1 U15198 ( .A1(n12981), .A2(n15073), .ZN(n14594) );
  NAND2_X1 U15199 ( .A1(n15028), .A2(n14594), .ZN(n12982) );
  NAND4_X1 U15200 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        P3_U3221) );
  INV_X1 U15201 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U15202 ( .A1(n12986), .A2(n13029), .ZN(n12988) );
  INV_X1 U15203 ( .A(n13041), .ZN(n12987) );
  NAND2_X1 U15204 ( .A1(n12987), .A2(n15142), .ZN(n12991) );
  OAI211_X1 U15205 ( .C1(n15142), .C2(n12989), .A(n12988), .B(n12991), .ZN(
        P3_U3490) );
  NAND2_X1 U15206 ( .A1(n15140), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12990) );
  OAI211_X1 U15207 ( .C1(n13046), .C2(n12996), .A(n12991), .B(n12990), .ZN(
        P3_U3489) );
  INV_X1 U15208 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12994) );
  AOI21_X1 U15209 ( .B1(n12993), .B2(n14601), .A(n12992), .ZN(n13047) );
  MUX2_X1 U15210 ( .A(n12994), .B(n13047), .S(n15142), .Z(n12995) );
  OAI21_X1 U15211 ( .B1(n13050), .B2(n12996), .A(n12995), .ZN(P3_U3487) );
  INV_X1 U15212 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12997) );
  MUX2_X1 U15213 ( .A(n12997), .B(n13051), .S(n15142), .Z(n12999) );
  NAND2_X1 U15214 ( .A1(n13053), .A2(n13029), .ZN(n12998) );
  OAI211_X1 U15215 ( .C1(n13056), .C2(n13040), .A(n12999), .B(n12998), .ZN(
        P3_U3486) );
  AOI22_X1 U15216 ( .A1(n13001), .A2(n15118), .B1(n15073), .B2(n13000), .ZN(
        n13002) );
  NAND2_X1 U15217 ( .A1(n13003), .A2(n13002), .ZN(n13057) );
  MUX2_X1 U15218 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13057), .S(n15142), .Z(
        P3_U3485) );
  INV_X1 U15219 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13004) );
  MUX2_X1 U15220 ( .A(n13004), .B(n13058), .S(n15142), .Z(n13006) );
  NAND2_X1 U15221 ( .A1(n13060), .A2(n13029), .ZN(n13005) );
  OAI211_X1 U15222 ( .C1(n13040), .C2(n13063), .A(n13006), .B(n13005), .ZN(
        P3_U3484) );
  INV_X1 U15223 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13009) );
  AOI21_X1 U15224 ( .B1(n15073), .B2(n13008), .A(n13007), .ZN(n13064) );
  MUX2_X1 U15225 ( .A(n13009), .B(n13064), .S(n15142), .Z(n13010) );
  OAI21_X1 U15226 ( .B1(n13067), .B2(n13040), .A(n13010), .ZN(P3_U3483) );
  INV_X1 U15227 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13013) );
  AOI21_X1 U15228 ( .B1(n15073), .B2(n13012), .A(n13011), .ZN(n13068) );
  MUX2_X1 U15229 ( .A(n13013), .B(n13068), .S(n15142), .Z(n13014) );
  OAI21_X1 U15230 ( .B1(n13040), .B2(n13071), .A(n13014), .ZN(P3_U3482) );
  INV_X1 U15231 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13015) );
  MUX2_X1 U15232 ( .A(n13015), .B(n13072), .S(n15142), .Z(n13017) );
  NAND2_X1 U15233 ( .A1(n13073), .A2(n13029), .ZN(n13016) );
  OAI211_X1 U15234 ( .C1(n13076), .C2(n13040), .A(n13017), .B(n13016), .ZN(
        P3_U3481) );
  INV_X1 U15235 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13018) );
  MUX2_X1 U15236 ( .A(n13018), .B(n13077), .S(n15142), .Z(n13020) );
  NAND2_X1 U15237 ( .A1(n13079), .A2(n13029), .ZN(n13019) );
  OAI211_X1 U15238 ( .C1(n13040), .C2(n13082), .A(n13020), .B(n13019), .ZN(
        P3_U3480) );
  INV_X1 U15239 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13023) );
  AOI21_X1 U15240 ( .B1(n15073), .B2(n13022), .A(n13021), .ZN(n13083) );
  MUX2_X1 U15241 ( .A(n13023), .B(n13083), .S(n15142), .Z(n13024) );
  OAI21_X1 U15242 ( .B1(n13040), .B2(n13086), .A(n13024), .ZN(P3_U3479) );
  INV_X1 U15243 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13025) );
  MUX2_X1 U15244 ( .A(n13025), .B(n13087), .S(n15142), .Z(n13027) );
  NAND2_X1 U15245 ( .A1(n13089), .A2(n13029), .ZN(n13026) );
  OAI211_X1 U15246 ( .C1(n13092), .C2(n13040), .A(n13027), .B(n13026), .ZN(
        P3_U3478) );
  MUX2_X1 U15247 ( .A(n13028), .B(n13093), .S(n15142), .Z(n13031) );
  NAND2_X1 U15248 ( .A1(n13096), .A2(n13029), .ZN(n13030) );
  OAI211_X1 U15249 ( .C1(n13040), .C2(n13099), .A(n13031), .B(n13030), .ZN(
        P3_U3477) );
  INV_X1 U15250 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13034) );
  AOI21_X1 U15251 ( .B1(n15073), .B2(n13033), .A(n13032), .ZN(n13100) );
  MUX2_X1 U15252 ( .A(n13034), .B(n13100), .S(n15142), .Z(n13035) );
  OAI21_X1 U15253 ( .B1(n13040), .B2(n13103), .A(n13035), .ZN(P3_U3476) );
  AOI21_X1 U15254 ( .B1(n15073), .B2(n13037), .A(n13036), .ZN(n13104) );
  MUX2_X1 U15255 ( .A(n13038), .B(n13104), .S(n15142), .Z(n13039) );
  OAI21_X1 U15256 ( .B1(n13040), .B2(n13108), .A(n13039), .ZN(P3_U3475) );
  NOR2_X1 U15257 ( .A1(n13041), .A2(n15125), .ZN(n13044) );
  AOI21_X1 U15258 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15125), .A(n13044), 
        .ZN(n13042) );
  OAI21_X1 U15259 ( .B1(n13043), .B2(n13049), .A(n13042), .ZN(P3_U3458) );
  AOI21_X1 U15260 ( .B1(n15125), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13044), 
        .ZN(n13045) );
  OAI21_X1 U15261 ( .B1(n13046), .B2(n13049), .A(n13045), .ZN(P3_U3457) );
  INV_X1 U15262 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13048) );
  INV_X1 U15263 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13052) );
  MUX2_X1 U15264 ( .A(n13052), .B(n13051), .S(n15127), .Z(n13055) );
  NAND2_X1 U15265 ( .A1(n13053), .A2(n13095), .ZN(n13054) );
  OAI211_X1 U15266 ( .C1(n13056), .C2(n13107), .A(n13055), .B(n13054), .ZN(
        P3_U3454) );
  MUX2_X1 U15267 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13057), .S(n15127), .Z(
        P3_U3453) );
  INV_X1 U15268 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13059) );
  MUX2_X1 U15269 ( .A(n13059), .B(n13058), .S(n15127), .Z(n13062) );
  NAND2_X1 U15270 ( .A1(n13060), .A2(n13095), .ZN(n13061) );
  OAI211_X1 U15271 ( .C1(n13063), .C2(n13107), .A(n13062), .B(n13061), .ZN(
        P3_U3452) );
  INV_X1 U15272 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13065) );
  MUX2_X1 U15273 ( .A(n13065), .B(n13064), .S(n15127), .Z(n13066) );
  OAI21_X1 U15274 ( .B1(n13067), .B2(n13107), .A(n13066), .ZN(P3_U3451) );
  INV_X1 U15275 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13069) );
  MUX2_X1 U15276 ( .A(n13069), .B(n13068), .S(n15127), .Z(n13070) );
  OAI21_X1 U15277 ( .B1(n13071), .B2(n13107), .A(n13070), .ZN(P3_U3450) );
  INV_X1 U15278 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n15419) );
  MUX2_X1 U15279 ( .A(n15419), .B(n13072), .S(n15127), .Z(n13075) );
  NAND2_X1 U15280 ( .A1(n13073), .A2(n13095), .ZN(n13074) );
  OAI211_X1 U15281 ( .C1(n13076), .C2(n13107), .A(n13075), .B(n13074), .ZN(
        P3_U3449) );
  INV_X1 U15282 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13078) );
  MUX2_X1 U15283 ( .A(n13078), .B(n13077), .S(n15127), .Z(n13081) );
  NAND2_X1 U15284 ( .A1(n13079), .A2(n13095), .ZN(n13080) );
  OAI211_X1 U15285 ( .C1(n13082), .C2(n13107), .A(n13081), .B(n13080), .ZN(
        P3_U3448) );
  INV_X1 U15286 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13084) );
  MUX2_X1 U15287 ( .A(n13084), .B(n13083), .S(n15127), .Z(n13085) );
  OAI21_X1 U15288 ( .B1(n13086), .B2(n13107), .A(n13085), .ZN(P3_U3447) );
  INV_X1 U15289 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13088) );
  MUX2_X1 U15290 ( .A(n13088), .B(n13087), .S(n15127), .Z(n13091) );
  NAND2_X1 U15291 ( .A1(n13089), .A2(n13095), .ZN(n13090) );
  OAI211_X1 U15292 ( .C1(n13092), .C2(n13107), .A(n13091), .B(n13090), .ZN(
        P3_U3446) );
  INV_X1 U15293 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U15294 ( .A(n13094), .B(n13093), .S(n15127), .Z(n13098) );
  NAND2_X1 U15295 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  OAI211_X1 U15296 ( .C1(n13099), .C2(n13107), .A(n13098), .B(n13097), .ZN(
        P3_U3444) );
  INV_X1 U15297 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13101) );
  MUX2_X1 U15298 ( .A(n13101), .B(n13100), .S(n15127), .Z(n13102) );
  OAI21_X1 U15299 ( .B1(n13103), .B2(n13107), .A(n13102), .ZN(P3_U3441) );
  INV_X1 U15300 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13105) );
  MUX2_X1 U15301 ( .A(n13105), .B(n13104), .S(n15127), .Z(n13106) );
  OAI21_X1 U15302 ( .B1(n13108), .B2(n13107), .A(n13106), .ZN(P3_U3438) );
  NAND2_X1 U15303 ( .A1(n13110), .A2(n13109), .ZN(n13114) );
  NAND4_X1 U15304 ( .A1(n8714), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n13112), .ZN(n13113) );
  OAI211_X1 U15305 ( .C1(n13116), .C2(n13115), .A(n13114), .B(n13113), .ZN(
        P3_U3264) );
  INV_X1 U15306 ( .A(n13117), .ZN(n13119) );
  OAI222_X1 U15307 ( .A1(n13122), .A2(n13121), .B1(n13120), .B2(n13119), .C1(
        n13118), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15308 ( .A(n13421), .ZN(n13131) );
  NAND2_X1 U15309 ( .A1(n13241), .A2(n13230), .ZN(n13127) );
  NAND2_X1 U15310 ( .A1(n13243), .A2(n13231), .ZN(n13126) );
  NAND2_X1 U15311 ( .A1(n13127), .A2(n13126), .ZN(n13416) );
  INV_X1 U15312 ( .A(n13416), .ZN(n13129) );
  OAI22_X1 U15313 ( .A1(n14811), .A2(n13129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13128), .ZN(n13130) );
  AOI21_X1 U15314 ( .B1(n13131), .B2(n13223), .A(n13130), .ZN(n13132) );
  INV_X1 U15315 ( .A(n13648), .ZN(n13486) );
  OAI22_X1 U15316 ( .A1(n13133), .A2(n14813), .B1(n13192), .B2(n13213), .ZN(
        n13135) );
  NAND2_X1 U15317 ( .A1(n13135), .A2(n13134), .ZN(n13139) );
  OAI22_X1 U15318 ( .A1(n13214), .A2(n13191), .B1(n13167), .B2(n13193), .ZN(
        n13480) );
  INV_X1 U15319 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13136) );
  OAI22_X1 U15320 ( .A1(n14821), .A2(n13482), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13136), .ZN(n13137) );
  AOI21_X1 U15321 ( .B1(n13480), .B2(n13235), .A(n13137), .ZN(n13138) );
  OAI211_X1 U15322 ( .C1(n13486), .C2(n13238), .A(n13139), .B(n13138), .ZN(
        P2_U3188) );
  INV_X1 U15323 ( .A(n13228), .ZN(n13143) );
  NOR3_X1 U15324 ( .A1(n13141), .A2(n13140), .A3(n13213), .ZN(n13142) );
  AOI21_X1 U15325 ( .B1(n13143), .B2(n13227), .A(n13142), .ZN(n13151) );
  NAND2_X1 U15326 ( .A1(n13672), .A2(n14818), .ZN(n13147) );
  AND2_X1 U15327 ( .A1(n13251), .A2(n13231), .ZN(n13144) );
  AOI21_X1 U15328 ( .B1(n13249), .B2(n13230), .A(n13144), .ZN(n13538) );
  INV_X1 U15329 ( .A(n13538), .ZN(n13145) );
  AOI22_X1 U15330 ( .A1(n13145), .A2(n13235), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13146) );
  OAI211_X1 U15331 ( .C1(n14821), .C2(n13544), .A(n13147), .B(n13146), .ZN(
        n13148) );
  AOI21_X1 U15332 ( .B1(n6561), .B2(n13227), .A(n13148), .ZN(n13149) );
  OAI21_X1 U15333 ( .B1(n13151), .B2(n13150), .A(n13149), .ZN(P2_U3191) );
  INV_X1 U15334 ( .A(n13512), .ZN(n13726) );
  AOI21_X1 U15335 ( .B1(n13153), .B2(n13152), .A(n14813), .ZN(n13155) );
  NAND2_X1 U15336 ( .A1(n13155), .A2(n13154), .ZN(n13160) );
  AOI22_X1 U15337 ( .A1(n13247), .A2(n13230), .B1(n13231), .B2(n13249), .ZN(
        n13508) );
  INV_X1 U15338 ( .A(n13508), .ZN(n13158) );
  OAI22_X1 U15339 ( .A1(n14821), .A2(n13514), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13156), .ZN(n13157) );
  AOI21_X1 U15340 ( .B1(n13158), .B2(n13235), .A(n13157), .ZN(n13159) );
  OAI211_X1 U15341 ( .C1(n13726), .C2(n13238), .A(n13160), .B(n13159), .ZN(
        P2_U3195) );
  INV_X1 U15342 ( .A(n13162), .ZN(n13163) );
  AOI21_X1 U15343 ( .B1(n13161), .B2(n13163), .A(n14813), .ZN(n13166) );
  NOR3_X1 U15344 ( .A1(n13164), .A2(n13167), .A3(n13213), .ZN(n13165) );
  OAI21_X1 U15345 ( .B1(n13166), .B2(n13165), .A(n12360), .ZN(n13171) );
  OAI22_X1 U15346 ( .A1(n7139), .A2(n13193), .B1(n13167), .B2(n13191), .ZN(
        n13445) );
  AOI22_X1 U15347 ( .A1(n13235), .A2(n13445), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13168) );
  OAI21_X1 U15348 ( .B1(n13450), .B2(n14821), .A(n13168), .ZN(n13169) );
  AOI21_X1 U15349 ( .B1(n13638), .B2(n14818), .A(n13169), .ZN(n13170) );
  NAND2_X1 U15350 ( .A1(n13171), .A2(n13170), .ZN(P2_U3197) );
  NAND2_X1 U15351 ( .A1(n13172), .A2(n13227), .ZN(n13188) );
  INV_X1 U15352 ( .A(n13173), .ZN(n13174) );
  OR2_X1 U15353 ( .A1(n14821), .A2(n13174), .ZN(n13176) );
  NAND2_X1 U15354 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13175) );
  OAI211_X1 U15355 ( .C1(n14811), .C2(n13177), .A(n13176), .B(n13175), .ZN(
        n13178) );
  INV_X1 U15356 ( .A(n13178), .ZN(n13187) );
  INV_X1 U15357 ( .A(n13265), .ZN(n13180) );
  OAI22_X1 U15358 ( .A1(n13213), .A2(n13180), .B1(n13179), .B2(n14813), .ZN(
        n13181) );
  NAND3_X1 U15359 ( .A1(n13183), .A2(n13182), .A3(n13181), .ZN(n13186) );
  NAND2_X1 U15360 ( .A1(n14818), .A2(n13184), .ZN(n13185) );
  NAND4_X1 U15361 ( .A1(n13188), .A2(n13187), .A3(n13186), .A4(n13185), .ZN(
        P2_U3199) );
  INV_X1 U15362 ( .A(n13643), .ZN(n13200) );
  OAI211_X1 U15363 ( .C1(n13190), .C2(n13189), .A(n13161), .B(n13227), .ZN(
        n13199) );
  INV_X1 U15364 ( .A(n13467), .ZN(n13197) );
  OAI22_X1 U15365 ( .A1(n13194), .A2(n13193), .B1(n13192), .B2(n13191), .ZN(
        n13462) );
  INV_X1 U15366 ( .A(n13462), .ZN(n13195) );
  INV_X1 U15367 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15226) );
  OAI22_X1 U15368 ( .A1(n13195), .A2(n14811), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15226), .ZN(n13196) );
  AOI21_X1 U15369 ( .B1(n13197), .B2(n13223), .A(n13196), .ZN(n13198) );
  OAI211_X1 U15370 ( .C1(n13200), .C2(n13238), .A(n13199), .B(n13198), .ZN(
        P2_U3201) );
  INV_X1 U15371 ( .A(n13528), .ZN(n13204) );
  NAND2_X1 U15372 ( .A1(n13248), .A2(n13230), .ZN(n13202) );
  NAND2_X1 U15373 ( .A1(n13250), .A2(n13231), .ZN(n13201) );
  NAND2_X1 U15374 ( .A1(n13202), .A2(n13201), .ZN(n13523) );
  AOI22_X1 U15375 ( .A1(n13523), .A2(n13235), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13203) );
  OAI21_X1 U15376 ( .B1(n13204), .B2(n14821), .A(n13203), .ZN(n13210) );
  AOI22_X1 U15377 ( .A1(n13206), .A2(n13227), .B1(n13205), .B2(n13250), .ZN(
        n13208) );
  NOR3_X1 U15378 ( .A1(n6561), .A2(n13208), .A3(n13207), .ZN(n13209) );
  AOI211_X1 U15379 ( .C1(n13529), .C2(n14818), .A(n13210), .B(n13209), .ZN(
        n13211) );
  OAI21_X1 U15380 ( .B1(n13212), .B2(n14813), .A(n13211), .ZN(P2_U3205) );
  OAI22_X1 U15381 ( .A1(n13215), .A2(n14813), .B1(n13214), .B2(n13213), .ZN(
        n13217) );
  NAND2_X1 U15382 ( .A1(n13217), .A2(n13216), .ZN(n13226) );
  INV_X1 U15383 ( .A(n13497), .ZN(n13224) );
  NAND2_X1 U15384 ( .A1(n13248), .A2(n13231), .ZN(n13219) );
  NAND2_X1 U15385 ( .A1(n13246), .A2(n13230), .ZN(n13218) );
  NAND2_X1 U15386 ( .A1(n13219), .A2(n13218), .ZN(n13491) );
  INV_X1 U15387 ( .A(n13491), .ZN(n13221) );
  OAI22_X1 U15388 ( .A1(n13221), .A2(n14811), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13220), .ZN(n13222) );
  AOI21_X1 U15389 ( .B1(n13224), .B2(n13223), .A(n13222), .ZN(n13225) );
  OAI211_X1 U15390 ( .C1(n7370), .C2(n13238), .A(n13226), .B(n13225), .ZN(
        P2_U3207) );
  OAI211_X1 U15391 ( .C1(n6685), .C2(n13229), .A(n13228), .B(n13227), .ZN(
        n13237) );
  NAND2_X1 U15392 ( .A1(n13250), .A2(n13230), .ZN(n13233) );
  NAND2_X1 U15393 ( .A1(n13252), .A2(n13231), .ZN(n13232) );
  NAND2_X1 U15394 ( .A1(n13233), .A2(n13232), .ZN(n13550) );
  AND2_X1 U15395 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13360) );
  NOR2_X1 U15396 ( .A1(n14821), .A2(n13559), .ZN(n13234) );
  AOI211_X1 U15397 ( .C1(n13235), .C2(n13550), .A(n13360), .B(n13234), .ZN(
        n13236) );
  OAI211_X1 U15398 ( .C1(n6910), .C2(n13238), .A(n13237), .B(n13236), .ZN(
        P2_U3210) );
  MUX2_X1 U15399 ( .A(n13390), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13268), .Z(
        P2_U3562) );
  MUX2_X1 U15400 ( .A(n13239), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13268), .Z(
        P2_U3561) );
  MUX2_X1 U15401 ( .A(n13240), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13268), .Z(
        P2_U3560) );
  MUX2_X1 U15402 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13241), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15403 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13242), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15404 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13243), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15405 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13244), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15406 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13245), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15407 ( .A(n13246), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13268), .Z(
        P2_U3554) );
  MUX2_X1 U15408 ( .A(n13247), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13268), .Z(
        P2_U3553) );
  MUX2_X1 U15409 ( .A(n13248), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13268), .Z(
        P2_U3552) );
  MUX2_X1 U15410 ( .A(n13249), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13268), .Z(
        P2_U3551) );
  MUX2_X1 U15411 ( .A(n13250), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13268), .Z(
        P2_U3550) );
  MUX2_X1 U15412 ( .A(n13251), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13268), .Z(
        P2_U3549) );
  MUX2_X1 U15413 ( .A(n13252), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13268), .Z(
        P2_U3548) );
  MUX2_X1 U15414 ( .A(n13253), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13268), .Z(
        P2_U3547) );
  MUX2_X1 U15415 ( .A(n13254), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13268), .Z(
        P2_U3546) );
  MUX2_X1 U15416 ( .A(n13255), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13268), .Z(
        P2_U3545) );
  MUX2_X1 U15417 ( .A(n13256), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13268), .Z(
        P2_U3544) );
  MUX2_X1 U15418 ( .A(n13257), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13268), .Z(
        P2_U3543) );
  MUX2_X1 U15419 ( .A(n13258), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13268), .Z(
        P2_U3542) );
  MUX2_X1 U15420 ( .A(n13259), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13268), .Z(
        P2_U3541) );
  MUX2_X1 U15421 ( .A(n13260), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13268), .Z(
        P2_U3540) );
  MUX2_X1 U15422 ( .A(n13261), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13268), .Z(
        P2_U3539) );
  MUX2_X1 U15423 ( .A(n13262), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13268), .Z(
        P2_U3538) );
  MUX2_X1 U15424 ( .A(n13263), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13268), .Z(
        P2_U3537) );
  MUX2_X1 U15425 ( .A(n13264), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13268), .Z(
        P2_U3536) );
  MUX2_X1 U15426 ( .A(n13265), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13268), .Z(
        P2_U3535) );
  MUX2_X1 U15427 ( .A(n13266), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13268), .Z(
        P2_U3534) );
  MUX2_X1 U15428 ( .A(n13267), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13268), .Z(
        P2_U3533) );
  MUX2_X1 U15429 ( .A(n13269), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13268), .Z(
        P2_U3532) );
  OAI22_X1 U15430 ( .A1(n13358), .A2(n13271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13270), .ZN(n13272) );
  AOI21_X1 U15431 ( .B1(n14809), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n13272), .ZN(
        n13282) );
  INV_X1 U15432 ( .A(n13273), .ZN(n13276) );
  OAI21_X1 U15433 ( .B1(n8904), .B2(n7014), .A(n13274), .ZN(n13275) );
  NAND3_X1 U15434 ( .A1(n14867), .A2(n13276), .A3(n13275), .ZN(n13281) );
  OAI211_X1 U15435 ( .C1(n13279), .C2(n13278), .A(n13380), .B(n13277), .ZN(
        n13280) );
  NAND3_X1 U15436 ( .A1(n13282), .A2(n13281), .A3(n13280), .ZN(P2_U3215) );
  OAI21_X1 U15437 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n13286) );
  NAND2_X1 U15438 ( .A1(n13286), .A2(n13380), .ZN(n13296) );
  NOR2_X1 U15439 ( .A1(n13358), .A2(n13287), .ZN(n13288) );
  AOI211_X1 U15440 ( .C1(n14809), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n13289), .B(
        n13288), .ZN(n13295) );
  OAI21_X1 U15441 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13293) );
  NAND2_X1 U15442 ( .A1(n13293), .A2(n14867), .ZN(n13294) );
  NAND3_X1 U15443 ( .A1(n13296), .A2(n13295), .A3(n13294), .ZN(P2_U3223) );
  OAI21_X1 U15444 ( .B1(n13299), .B2(n13298), .A(n13297), .ZN(n13300) );
  NAND2_X1 U15445 ( .A1(n13300), .A2(n13380), .ZN(n13311) );
  OAI21_X1 U15446 ( .B1(n13358), .B2(n13302), .A(n13301), .ZN(n13303) );
  AOI21_X1 U15447 ( .B1(n14809), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n13303), 
        .ZN(n13310) );
  AND3_X1 U15448 ( .A1(n13306), .A2(n13305), .A3(n13304), .ZN(n13307) );
  OAI21_X1 U15449 ( .B1(n13308), .B2(n13307), .A(n14867), .ZN(n13309) );
  NAND3_X1 U15450 ( .A1(n13311), .A2(n13310), .A3(n13309), .ZN(P2_U3226) );
  NOR2_X1 U15451 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13312), .ZN(n13315) );
  NOR2_X1 U15452 ( .A1(n13358), .A2(n13313), .ZN(n13314) );
  AOI211_X1 U15453 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n14809), .A(n13315), 
        .B(n13314), .ZN(n13324) );
  AOI211_X1 U15454 ( .C1(n13318), .C2(n13317), .A(n13316), .B(n14858), .ZN(
        n13319) );
  INV_X1 U15455 ( .A(n13319), .ZN(n13323) );
  OAI211_X1 U15456 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n13321), .A(n14867), 
        .B(n13320), .ZN(n13322) );
  NAND3_X1 U15457 ( .A1(n13324), .A2(n13323), .A3(n13322), .ZN(P2_U3228) );
  OAI211_X1 U15458 ( .C1(n13326), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14867), 
        .B(n13325), .ZN(n13336) );
  INV_X1 U15459 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n15184) );
  NOR2_X1 U15460 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15184), .ZN(n13327) );
  AOI21_X1 U15461 ( .B1(n14865), .B2(n13328), .A(n13327), .ZN(n13335) );
  INV_X1 U15462 ( .A(n13329), .ZN(n13332) );
  INV_X1 U15463 ( .A(n13330), .ZN(n13331) );
  OAI211_X1 U15464 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n13332), .A(n13380), 
        .B(n13331), .ZN(n13334) );
  NAND2_X1 U15465 ( .A1(n14809), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n13333) );
  NAND4_X1 U15466 ( .A1(n13336), .A2(n13335), .A3(n13334), .A4(n13333), .ZN(
        P2_U3229) );
  NAND2_X1 U15467 ( .A1(n13338), .A2(n13337), .ZN(n13341) );
  NOR2_X1 U15468 ( .A1(n13364), .A2(n13575), .ZN(n13339) );
  AOI21_X1 U15469 ( .B1(n13575), .B2(n13364), .A(n13339), .ZN(n13340) );
  NAND2_X1 U15470 ( .A1(n13340), .A2(n13341), .ZN(n13353) );
  OAI211_X1 U15471 ( .C1(n13341), .C2(n13340), .A(n14867), .B(n13353), .ZN(
        n13352) );
  AND2_X1 U15472 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13342) );
  AOI21_X1 U15473 ( .B1(n14865), .B2(n13346), .A(n13342), .ZN(n13343) );
  INV_X1 U15474 ( .A(n13343), .ZN(n13350) );
  AOI21_X1 U15475 ( .B1(n13345), .B2(P2_REG1_REG_16__SCAN_IN), .A(n13344), 
        .ZN(n13348) );
  XNOR2_X1 U15476 ( .A(n13346), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13347) );
  NOR2_X1 U15477 ( .A1(n13348), .A2(n13347), .ZN(n13361) );
  AOI211_X1 U15478 ( .C1(n13348), .C2(n13347), .A(n13361), .B(n14858), .ZN(
        n13349) );
  AOI211_X1 U15479 ( .C1(n14809), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n13350), 
        .B(n13349), .ZN(n13351) );
  NAND2_X1 U15480 ( .A1(n13352), .A2(n13351), .ZN(P2_U3231) );
  OAI21_X1 U15481 ( .B1(n13364), .B2(n13575), .A(n13353), .ZN(n13354) );
  AND2_X1 U15482 ( .A1(n13354), .A2(n13365), .ZN(n13355) );
  NOR2_X1 U15483 ( .A1(n13354), .A2(n13365), .ZN(n13378) );
  OR2_X1 U15484 ( .A1(n13355), .A2(n13378), .ZN(n13356) );
  NOR2_X1 U15485 ( .A1(n13356), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13377) );
  AOI21_X1 U15486 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13356), .A(n13377), 
        .ZN(n13372) );
  NOR2_X1 U15487 ( .A1(n13358), .A2(n13357), .ZN(n13359) );
  AOI211_X1 U15488 ( .C1(n14809), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13360), 
        .B(n13359), .ZN(n13371) );
  INV_X1 U15489 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13363) );
  INV_X1 U15490 ( .A(n13361), .ZN(n13362) );
  OAI21_X1 U15491 ( .B1(n13364), .B2(n13363), .A(n13362), .ZN(n13366) );
  AND2_X1 U15492 ( .A1(n13366), .A2(n13365), .ZN(n13373) );
  NOR2_X1 U15493 ( .A1(n13366), .A2(n13365), .ZN(n13367) );
  NOR2_X1 U15494 ( .A1(n13373), .A2(n13367), .ZN(n13369) );
  AND2_X1 U15495 ( .A1(n13369), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13374) );
  INV_X1 U15496 ( .A(n13374), .ZN(n13368) );
  OAI211_X1 U15497 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13369), .A(n13380), 
        .B(n13368), .ZN(n13370) );
  OAI211_X1 U15498 ( .C1(n13372), .C2(n14851), .A(n13371), .B(n13370), .ZN(
        P2_U3232) );
  NOR2_X1 U15499 ( .A1(n13374), .A2(n13373), .ZN(n13376) );
  XNOR2_X1 U15500 ( .A(n13376), .B(n13375), .ZN(n13381) );
  NOR2_X1 U15501 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  XNOR2_X1 U15502 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13379), .ZN(n13382) );
  NAND2_X1 U15503 ( .A1(n13381), .A2(n13380), .ZN(n13384) );
  AOI21_X1 U15504 ( .B1(n13382), .B2(n14867), .A(n14865), .ZN(n13383) );
  NAND2_X1 U15505 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13385)
         );
  NOR2_X2 U15506 ( .A1(n13387), .A2(n14896), .ZN(n13608) );
  NAND2_X1 U15507 ( .A1(n13608), .A2(n14874), .ZN(n13393) );
  INV_X1 U15508 ( .A(n13388), .ZN(n13389) );
  AND2_X1 U15509 ( .A1(n13390), .A2(n13389), .ZN(n13611) );
  INV_X1 U15510 ( .A(n13611), .ZN(n13391) );
  NOR2_X1 U15511 ( .A1(n13561), .A2(n13391), .ZN(n13397) );
  AOI21_X1 U15512 ( .B1(n13561), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13397), 
        .ZN(n13392) );
  OAI211_X1 U15513 ( .C1(n7372), .C2(n14879), .A(n13393), .B(n13392), .ZN(
        P2_U3234) );
  AOI211_X1 U15514 ( .C1(n13396), .C2(n13395), .A(n14896), .B(n13394), .ZN(
        n13612) );
  NAND2_X1 U15515 ( .A1(n13612), .A2(n14874), .ZN(n13399) );
  AOI21_X1 U15516 ( .B1(n13561), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13397), 
        .ZN(n13398) );
  OAI211_X1 U15517 ( .C1(n13707), .C2(n14879), .A(n13399), .B(n13398), .ZN(
        P2_U3235) );
  INV_X1 U15518 ( .A(n13400), .ZN(n13405) );
  NAND2_X1 U15519 ( .A1(n13404), .A2(n13403), .ZN(n13620) );
  AOI21_X1 U15520 ( .B1(n13405), .B2(n14902), .A(n13620), .ZN(n13414) );
  XNOR2_X1 U15521 ( .A(n13407), .B(n13406), .ZN(n13622) );
  NAND2_X1 U15522 ( .A1(n13622), .A2(n14883), .ZN(n13413) );
  AOI211_X1 U15523 ( .C1(n13409), .C2(n13420), .A(n14896), .B(n7374), .ZN(
        n13621) );
  INV_X1 U15524 ( .A(n13409), .ZN(n13710) );
  OAI22_X1 U15525 ( .A1(n13710), .A2(n14879), .B1(n13598), .B2(n13410), .ZN(
        n13411) );
  AOI21_X1 U15526 ( .B1(n13621), .B2(n14874), .A(n13411), .ZN(n13412) );
  OAI211_X1 U15527 ( .C1(n13561), .C2(n13414), .A(n13413), .B(n13412), .ZN(
        P2_U3237) );
  XNOR2_X1 U15528 ( .A(n13415), .B(n13418), .ZN(n13417) );
  AOI21_X1 U15529 ( .B1(n13417), .B2(n14892), .A(n13416), .ZN(n13626) );
  XNOR2_X1 U15530 ( .A(n13419), .B(n13418), .ZN(n13627) );
  INV_X1 U15531 ( .A(n13627), .ZN(n13427) );
  OAI211_X1 U15532 ( .C1(n13714), .C2(n13436), .A(n13557), .B(n13420), .ZN(
        n13625) );
  INV_X1 U15533 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13422) );
  OAI22_X1 U15534 ( .A1(n13598), .A2(n13422), .B1(n13421), .B2(n13595), .ZN(
        n13423) );
  AOI21_X1 U15535 ( .B1(n13424), .B2(n13600), .A(n13423), .ZN(n13425) );
  OAI21_X1 U15536 ( .B1(n13625), .B2(n13578), .A(n13425), .ZN(n13426) );
  AOI21_X1 U15537 ( .B1(n13427), .B2(n14883), .A(n13426), .ZN(n13428) );
  OAI21_X1 U15538 ( .B1(n13626), .B2(n13561), .A(n13428), .ZN(P2_U3238) );
  XNOR2_X1 U15539 ( .A(n13429), .B(n13432), .ZN(n13431) );
  AOI21_X1 U15540 ( .B1(n13431), .B2(n14892), .A(n13430), .ZN(n13634) );
  XNOR2_X1 U15541 ( .A(n13433), .B(n13432), .ZN(n13631) );
  NAND2_X1 U15542 ( .A1(n13440), .A2(n13447), .ZN(n13434) );
  NAND2_X1 U15543 ( .A1(n13434), .A2(n13557), .ZN(n13435) );
  OR2_X1 U15544 ( .A1(n13436), .A2(n13435), .ZN(n13632) );
  INV_X1 U15545 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13438) );
  OAI22_X1 U15546 ( .A1(n13598), .A2(n13438), .B1(n13437), .B2(n13595), .ZN(
        n13439) );
  AOI21_X1 U15547 ( .B1(n13440), .B2(n13600), .A(n13439), .ZN(n13441) );
  OAI21_X1 U15548 ( .B1(n13632), .B2(n13578), .A(n13441), .ZN(n13442) );
  AOI21_X1 U15549 ( .B1(n13631), .B2(n14883), .A(n13442), .ZN(n13443) );
  OAI21_X1 U15550 ( .B1(n13634), .B2(n13561), .A(n13443), .ZN(P2_U3239) );
  XNOR2_X1 U15551 ( .A(n13457), .B(n13444), .ZN(n13446) );
  AOI21_X1 U15552 ( .B1(n13446), .B2(n14892), .A(n13445), .ZN(n13640) );
  INV_X1 U15553 ( .A(n13472), .ZN(n13449) );
  INV_X1 U15554 ( .A(n13447), .ZN(n13448) );
  AOI211_X1 U15555 ( .C1(n13638), .C2(n13449), .A(n14896), .B(n13448), .ZN(
        n13637) );
  INV_X1 U15556 ( .A(n13598), .ZN(n13561) );
  INV_X1 U15557 ( .A(n13450), .ZN(n13451) );
  AOI22_X1 U15558 ( .A1(n13561), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13451), 
        .B2(n14902), .ZN(n13452) );
  OAI21_X1 U15559 ( .B1(n13453), .B2(n14879), .A(n13452), .ZN(n13459) );
  INV_X1 U15560 ( .A(n13454), .ZN(n13455) );
  AOI21_X1 U15561 ( .B1(n13457), .B2(n13456), .A(n13455), .ZN(n13641) );
  NOR2_X1 U15562 ( .A1(n13641), .A2(n13582), .ZN(n13458) );
  AOI211_X1 U15563 ( .C1(n13637), .C2(n14874), .A(n13459), .B(n13458), .ZN(
        n13460) );
  OAI21_X1 U15564 ( .B1(n13561), .B2(n13640), .A(n13460), .ZN(P2_U3240) );
  XNOR2_X1 U15565 ( .A(n13461), .B(n13464), .ZN(n13463) );
  AOI21_X1 U15566 ( .B1(n13463), .B2(n14892), .A(n13462), .ZN(n13645) );
  INV_X1 U15567 ( .A(n13464), .ZN(n13466) );
  OAI21_X1 U15568 ( .B1(n6602), .B2(n13466), .A(n13465), .ZN(n13646) );
  OAI22_X1 U15569 ( .A1(n13598), .A2(n13468), .B1(n13467), .B2(n13595), .ZN(
        n13469) );
  AOI21_X1 U15570 ( .B1(n13643), .B2(n13600), .A(n13469), .ZN(n13474) );
  NAND2_X1 U15571 ( .A1(n13643), .A2(n13484), .ZN(n13470) );
  NAND2_X1 U15572 ( .A1(n13470), .A2(n13557), .ZN(n13471) );
  NOR2_X1 U15573 ( .A1(n13472), .A2(n13471), .ZN(n13642) );
  NAND2_X1 U15574 ( .A1(n13642), .A2(n14874), .ZN(n13473) );
  OAI211_X1 U15575 ( .C1(n13646), .C2(n13582), .A(n13474), .B(n13473), .ZN(
        n13475) );
  INV_X1 U15576 ( .A(n13475), .ZN(n13476) );
  OAI21_X1 U15577 ( .B1(n13561), .B2(n13645), .A(n13476), .ZN(P2_U3241) );
  XOR2_X1 U15578 ( .A(n13477), .B(n13478), .Z(n13651) );
  XOR2_X1 U15579 ( .A(n13479), .B(n13478), .Z(n13481) );
  AOI21_X1 U15580 ( .B1(n13481), .B2(n14892), .A(n13480), .ZN(n13650) );
  OAI21_X1 U15581 ( .B1(n13482), .B2(n13595), .A(n13650), .ZN(n13483) );
  NAND2_X1 U15582 ( .A1(n13483), .A2(n13598), .ZN(n13489) );
  AOI211_X1 U15583 ( .C1(n13648), .C2(n13499), .A(n14896), .B(n6909), .ZN(
        n13647) );
  OAI22_X1 U15584 ( .A1(n13486), .A2(n14879), .B1(n13598), .B2(n13485), .ZN(
        n13487) );
  AOI21_X1 U15585 ( .B1(n13647), .B2(n14874), .A(n13487), .ZN(n13488) );
  OAI211_X1 U15586 ( .C1(n13651), .C2(n13582), .A(n13489), .B(n13488), .ZN(
        P2_U3242) );
  XNOR2_X1 U15587 ( .A(n13490), .B(n13494), .ZN(n13492) );
  AOI21_X1 U15588 ( .B1(n13492), .B2(n14892), .A(n13491), .ZN(n13655) );
  OAI21_X1 U15589 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(n13656) );
  OAI22_X1 U15590 ( .A1(n13497), .A2(n13595), .B1(n13598), .B2(n13496), .ZN(
        n13498) );
  AOI21_X1 U15591 ( .B1(n13653), .B2(n13600), .A(n13498), .ZN(n13502) );
  AOI21_X1 U15592 ( .B1(n13653), .B2(n13511), .A(n14896), .ZN(n13500) );
  AND2_X1 U15593 ( .A1(n13500), .A2(n13499), .ZN(n13652) );
  NAND2_X1 U15594 ( .A1(n13652), .A2(n14874), .ZN(n13501) );
  OAI211_X1 U15595 ( .C1(n13656), .C2(n13582), .A(n13502), .B(n13501), .ZN(
        n13503) );
  INV_X1 U15596 ( .A(n13503), .ZN(n13504) );
  OAI21_X1 U15597 ( .B1(n13655), .B2(n13561), .A(n13504), .ZN(P2_U3243) );
  XNOR2_X1 U15598 ( .A(n13505), .B(n13506), .ZN(n13659) );
  INV_X1 U15599 ( .A(n13659), .ZN(n13519) );
  XOR2_X1 U15600 ( .A(n13507), .B(n13506), .Z(n13510) );
  OAI21_X1 U15601 ( .B1(n13510), .B2(n13509), .A(n13508), .ZN(n13657) );
  NAND2_X1 U15602 ( .A1(n13657), .A2(n13598), .ZN(n13518) );
  AOI211_X1 U15603 ( .C1(n13512), .C2(n13527), .A(n14896), .B(n7371), .ZN(
        n13658) );
  NOR2_X1 U15604 ( .A1(n13726), .A2(n14879), .ZN(n13516) );
  OAI22_X1 U15605 ( .A1(n13514), .A2(n13595), .B1(n13598), .B2(n13513), .ZN(
        n13515) );
  AOI211_X1 U15606 ( .C1(n13658), .C2(n14874), .A(n13516), .B(n13515), .ZN(
        n13517) );
  OAI211_X1 U15607 ( .C1(n13519), .C2(n13582), .A(n13518), .B(n13517), .ZN(
        P2_U3244) );
  NAND2_X1 U15608 ( .A1(n13520), .A2(n13525), .ZN(n13521) );
  NAND2_X1 U15609 ( .A1(n13522), .A2(n13521), .ZN(n13524) );
  AOI21_X1 U15610 ( .B1(n13524), .B2(n14892), .A(n13523), .ZN(n13665) );
  XNOR2_X1 U15611 ( .A(n13526), .B(n13525), .ZN(n13662) );
  OAI211_X1 U15612 ( .C1(n13540), .C2(n13731), .A(n13557), .B(n13527), .ZN(
        n13663) );
  AOI22_X1 U15613 ( .A1(n13561), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13528), 
        .B2(n14902), .ZN(n13531) );
  NAND2_X1 U15614 ( .A1(n13529), .A2(n13600), .ZN(n13530) );
  OAI211_X1 U15615 ( .C1(n13663), .C2(n13578), .A(n13531), .B(n13530), .ZN(
        n13532) );
  AOI21_X1 U15616 ( .B1(n13662), .B2(n14883), .A(n13532), .ZN(n13533) );
  OAI21_X1 U15617 ( .B1(n13665), .B2(n13561), .A(n13533), .ZN(P2_U3245) );
  XNOR2_X1 U15618 ( .A(n13534), .B(n13536), .ZN(n13674) );
  OAI211_X1 U15619 ( .C1(n13537), .C2(n13536), .A(n13535), .B(n14892), .ZN(
        n13539) );
  NAND2_X1 U15620 ( .A1(n13539), .A2(n13538), .ZN(n13670) );
  AND2_X1 U15621 ( .A1(n13672), .A2(n13558), .ZN(n13541) );
  OR2_X1 U15622 ( .A1(n13541), .A2(n13540), .ZN(n13669) );
  NOR2_X1 U15623 ( .A1(n13669), .A2(n13542), .ZN(n13543) );
  OAI21_X1 U15624 ( .B1(n13670), .B2(n13543), .A(n13598), .ZN(n13548) );
  INV_X1 U15625 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13545) );
  OAI22_X1 U15626 ( .A1(n13598), .A2(n13545), .B1(n13544), .B2(n13595), .ZN(
        n13546) );
  AOI21_X1 U15627 ( .B1(n13672), .B2(n13600), .A(n13546), .ZN(n13547) );
  OAI211_X1 U15628 ( .C1(n13674), .C2(n13582), .A(n13548), .B(n13547), .ZN(
        P2_U3246) );
  XNOR2_X1 U15629 ( .A(n13549), .B(n8121), .ZN(n13551) );
  AOI21_X1 U15630 ( .B1(n13551), .B2(n14892), .A(n13550), .ZN(n13678) );
  NAND2_X1 U15631 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U15632 ( .A1(n6967), .A2(n13554), .ZN(n13676) );
  NAND2_X1 U15633 ( .A1(n13572), .A2(n13735), .ZN(n13556) );
  AND3_X1 U15634 ( .A1(n13558), .A2(n13557), .A3(n13556), .ZN(n13675) );
  NAND2_X1 U15635 ( .A1(n13675), .A2(n14874), .ZN(n13563) );
  INV_X1 U15636 ( .A(n13559), .ZN(n13560) );
  AOI22_X1 U15637 ( .A1(n13561), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13560), 
        .B2(n14902), .ZN(n13562) );
  OAI211_X1 U15638 ( .C1(n6910), .C2(n14879), .A(n13563), .B(n13562), .ZN(
        n13564) );
  AOI21_X1 U15639 ( .B1(n13676), .B2(n14883), .A(n13564), .ZN(n13565) );
  OAI21_X1 U15640 ( .B1(n13678), .B2(n13561), .A(n13565), .ZN(P2_U3247) );
  XNOR2_X1 U15641 ( .A(n13566), .B(n13567), .ZN(n13683) );
  XNOR2_X1 U15642 ( .A(n13568), .B(n13567), .ZN(n13570) );
  AOI21_X1 U15643 ( .B1(n13570), .B2(n14892), .A(n13569), .ZN(n13682) );
  INV_X1 U15644 ( .A(n13682), .ZN(n13580) );
  AOI21_X1 U15645 ( .B1(n13571), .B2(n13739), .A(n14896), .ZN(n13573) );
  NAND2_X1 U15646 ( .A1(n13573), .A2(n13572), .ZN(n13681) );
  OAI22_X1 U15647 ( .A1(n13598), .A2(n13575), .B1(n13574), .B2(n13595), .ZN(
        n13576) );
  AOI21_X1 U15648 ( .B1(n13739), .B2(n13600), .A(n13576), .ZN(n13577) );
  OAI21_X1 U15649 ( .B1(n13681), .B2(n13578), .A(n13577), .ZN(n13579) );
  AOI21_X1 U15650 ( .B1(n13580), .B2(n13598), .A(n13579), .ZN(n13581) );
  OAI21_X1 U15651 ( .B1(n13683), .B2(n13582), .A(n13581), .ZN(P2_U3248) );
  NAND2_X1 U15652 ( .A1(n13583), .A2(n13598), .ZN(n13593) );
  OAI22_X1 U15653 ( .A1(n13598), .A2(n13585), .B1(n13584), .B2(n13595), .ZN(
        n13586) );
  AOI21_X1 U15654 ( .B1(n13587), .B2(n13600), .A(n13586), .ZN(n13592) );
  NAND2_X1 U15655 ( .A1(n13588), .A2(n14883), .ZN(n13591) );
  NAND2_X1 U15656 ( .A1(n13589), .A2(n14874), .ZN(n13590) );
  NAND4_X1 U15657 ( .A1(n13593), .A2(n13592), .A3(n13591), .A4(n13590), .ZN(
        P2_U3253) );
  NAND2_X1 U15658 ( .A1(n13594), .A2(n13598), .ZN(n13607) );
  OAI22_X1 U15659 ( .A1(n13598), .A2(n13597), .B1(n13596), .B2(n13595), .ZN(
        n13599) );
  AOI21_X1 U15660 ( .B1(n13601), .B2(n13600), .A(n13599), .ZN(n13606) );
  NAND2_X1 U15661 ( .A1(n13602), .A2(n14883), .ZN(n13605) );
  NAND2_X1 U15662 ( .A1(n13603), .A2(n14874), .ZN(n13604) );
  NAND4_X1 U15663 ( .A1(n13607), .A2(n13606), .A3(n13605), .A4(n13604), .ZN(
        P2_U3255) );
  INV_X1 U15664 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13609) );
  NOR2_X1 U15665 ( .A1(n13608), .A2(n13611), .ZN(n13701) );
  MUX2_X1 U15666 ( .A(n13609), .B(n13701), .S(n14972), .Z(n13610) );
  OAI21_X1 U15667 ( .B1(n7372), .B2(n13668), .A(n13610), .ZN(P2_U3530) );
  INV_X1 U15668 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13613) );
  NOR2_X1 U15669 ( .A1(n13612), .A2(n13611), .ZN(n13704) );
  MUX2_X1 U15670 ( .A(n13613), .B(n13704), .S(n14972), .Z(n13614) );
  OAI21_X1 U15671 ( .B1(n13707), .B2(n13668), .A(n13614), .ZN(P2_U3529) );
  AOI21_X1 U15672 ( .B1(n14953), .B2(n13616), .A(n13615), .ZN(n13617) );
  INV_X1 U15673 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13623) );
  OAI211_X1 U15674 ( .C1(n13627), .C2(n13699), .A(n13626), .B(n13625), .ZN(
        n13628) );
  INV_X1 U15675 ( .A(n13628), .ZN(n13711) );
  MUX2_X1 U15676 ( .A(n13629), .B(n13711), .S(n14972), .Z(n13630) );
  OAI21_X1 U15677 ( .B1(n13714), .B2(n13668), .A(n13630), .ZN(P2_U3526) );
  NAND2_X1 U15678 ( .A1(n13631), .A2(n14927), .ZN(n13633) );
  NAND3_X1 U15679 ( .A1(n13634), .A2(n13633), .A3(n13632), .ZN(n13715) );
  MUX2_X1 U15680 ( .A(n13715), .B(P2_REG1_REG_26__SCAN_IN), .S(n14970), .Z(
        n13635) );
  INV_X1 U15681 ( .A(n13635), .ZN(n13636) );
  OAI21_X1 U15682 ( .B1(n13718), .B2(n13668), .A(n13636), .ZN(P2_U3525) );
  AOI21_X1 U15683 ( .B1(n14953), .B2(n13638), .A(n13637), .ZN(n13639) );
  OAI211_X1 U15684 ( .C1(n13641), .C2(n13699), .A(n13640), .B(n13639), .ZN(
        n13719) );
  MUX2_X1 U15685 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13719), .S(n14972), .Z(
        P2_U3524) );
  AOI21_X1 U15686 ( .B1(n14953), .B2(n13643), .A(n13642), .ZN(n13644) );
  OAI211_X1 U15687 ( .C1(n13646), .C2(n13699), .A(n13645), .B(n13644), .ZN(
        n13720) );
  MUX2_X1 U15688 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13720), .S(n14972), .Z(
        P2_U3523) );
  AOI21_X1 U15689 ( .B1(n14953), .B2(n13648), .A(n13647), .ZN(n13649) );
  OAI211_X1 U15690 ( .C1(n13651), .C2(n13699), .A(n13650), .B(n13649), .ZN(
        n13721) );
  MUX2_X1 U15691 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13721), .S(n14972), .Z(
        P2_U3522) );
  AOI21_X1 U15692 ( .B1(n14953), .B2(n13653), .A(n13652), .ZN(n13654) );
  OAI211_X1 U15693 ( .C1(n13699), .C2(n13656), .A(n13655), .B(n13654), .ZN(
        n13722) );
  MUX2_X1 U15694 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13722), .S(n14972), .Z(
        P2_U3521) );
  INV_X1 U15695 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13660) );
  AOI211_X1 U15696 ( .C1(n14927), .C2(n13659), .A(n13658), .B(n13657), .ZN(
        n13723) );
  MUX2_X1 U15697 ( .A(n13660), .B(n13723), .S(n14972), .Z(n13661) );
  OAI21_X1 U15698 ( .B1(n13726), .B2(n13668), .A(n13661), .ZN(P2_U3520) );
  NAND2_X1 U15699 ( .A1(n13662), .A2(n14927), .ZN(n13664) );
  NAND3_X1 U15700 ( .A1(n13665), .A2(n13664), .A3(n13663), .ZN(n13727) );
  MUX2_X1 U15701 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13727), .S(n14972), .Z(
        n13666) );
  INV_X1 U15702 ( .A(n13666), .ZN(n13667) );
  OAI21_X1 U15703 ( .B1(n13731), .B2(n13668), .A(n13667), .ZN(P2_U3519) );
  NOR2_X1 U15704 ( .A1(n13669), .A2(n14896), .ZN(n13671) );
  AOI211_X1 U15705 ( .C1(n14953), .C2(n13672), .A(n13671), .B(n13670), .ZN(
        n13673) );
  OAI21_X1 U15706 ( .B1(n13699), .B2(n13674), .A(n13673), .ZN(n13732) );
  MUX2_X1 U15707 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13732), .S(n14972), .Z(
        P2_U3518) );
  AOI21_X1 U15708 ( .B1(n13676), .B2(n14927), .A(n13675), .ZN(n13677) );
  NAND2_X1 U15709 ( .A1(n13678), .A2(n13677), .ZN(n13733) );
  MUX2_X1 U15710 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13733), .S(n14972), .Z(
        n13679) );
  AOI21_X1 U15711 ( .B1(n13692), .B2(n13735), .A(n13679), .ZN(n13680) );
  INV_X1 U15712 ( .A(n13680), .ZN(P2_U3517) );
  OAI211_X1 U15713 ( .C1(n13699), .C2(n13683), .A(n13682), .B(n13681), .ZN(
        n13737) );
  MUX2_X1 U15714 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13737), .S(n14972), .Z(
        n13684) );
  AOI21_X1 U15715 ( .B1(n13692), .B2(n13739), .A(n13684), .ZN(n13685) );
  INV_X1 U15716 ( .A(n13685), .ZN(P2_U3516) );
  AND2_X1 U15717 ( .A1(n13687), .A2(n13686), .ZN(n13689) );
  OAI211_X1 U15718 ( .C1(n13690), .C2(n13699), .A(n13689), .B(n13688), .ZN(
        n13741) );
  MUX2_X1 U15719 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13741), .S(n14972), .Z(
        n13691) );
  AOI21_X1 U15720 ( .B1(n13692), .B2(n13743), .A(n13691), .ZN(n13693) );
  INV_X1 U15721 ( .A(n13693), .ZN(P2_U3515) );
  AOI211_X1 U15722 ( .C1(n14953), .C2(n13696), .A(n13695), .B(n13694), .ZN(
        n13698) );
  OAI211_X1 U15723 ( .C1(n13700), .C2(n13699), .A(n13698), .B(n13697), .ZN(
        n13746) );
  MUX2_X1 U15724 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13746), .S(n14972), .Z(
        P2_U3514) );
  INV_X1 U15725 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13702) );
  MUX2_X1 U15726 ( .A(n13702), .B(n13701), .S(n14962), .Z(n13703) );
  OAI21_X1 U15727 ( .B1(n7372), .B2(n13730), .A(n13703), .ZN(P2_U3498) );
  INV_X1 U15728 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13705) );
  MUX2_X1 U15729 ( .A(n13705), .B(n13704), .S(n14962), .Z(n13706) );
  OAI21_X1 U15730 ( .B1(n13707), .B2(n13730), .A(n13706), .ZN(P2_U3497) );
  MUX2_X1 U15731 ( .A(n13712), .B(n13711), .S(n14962), .Z(n13713) );
  OAI21_X1 U15732 ( .B1(n13714), .B2(n13730), .A(n13713), .ZN(P2_U3494) );
  MUX2_X1 U15733 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13715), .S(n14962), .Z(
        n13716) );
  INV_X1 U15734 ( .A(n13716), .ZN(n13717) );
  OAI21_X1 U15735 ( .B1(n13718), .B2(n13730), .A(n13717), .ZN(P2_U3493) );
  MUX2_X1 U15736 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13719), .S(n14962), .Z(
        P2_U3492) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13720), .S(n14962), .Z(
        P2_U3491) );
  MUX2_X1 U15738 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13721), .S(n14962), .Z(
        P2_U3490) );
  MUX2_X1 U15739 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13722), .S(n14962), .Z(
        P2_U3489) );
  INV_X1 U15740 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13724) );
  MUX2_X1 U15741 ( .A(n13724), .B(n13723), .S(n14962), .Z(n13725) );
  OAI21_X1 U15742 ( .B1(n13726), .B2(n13730), .A(n13725), .ZN(P2_U3488) );
  MUX2_X1 U15743 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13727), .S(n14962), .Z(
        n13728) );
  INV_X1 U15744 ( .A(n13728), .ZN(n13729) );
  OAI21_X1 U15745 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(P2_U3487) );
  MUX2_X1 U15746 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13732), .S(n14962), .Z(
        P2_U3486) );
  MUX2_X1 U15747 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13733), .S(n14962), .Z(
        n13734) );
  AOI21_X1 U15748 ( .B1(n13744), .B2(n13735), .A(n13734), .ZN(n13736) );
  INV_X1 U15749 ( .A(n13736), .ZN(P2_U3484) );
  MUX2_X1 U15750 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13737), .S(n14962), .Z(
        n13738) );
  AOI21_X1 U15751 ( .B1(n13744), .B2(n13739), .A(n13738), .ZN(n13740) );
  INV_X1 U15752 ( .A(n13740), .ZN(P2_U3481) );
  MUX2_X1 U15753 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13741), .S(n14962), .Z(
        n13742) );
  AOI21_X1 U15754 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13745) );
  INV_X1 U15755 ( .A(n13745), .ZN(P2_U3478) );
  MUX2_X1 U15756 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13746), .S(n14962), .Z(
        P2_U3475) );
  NAND3_X1 U15757 ( .A1(n13748), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13751) );
  OAI22_X1 U15758 ( .A1(n13747), .A2(n13751), .B1(n13750), .B2(n13749), .ZN(
        n13752) );
  AOI21_X1 U15759 ( .B1(n13753), .B2(n13755), .A(n13752), .ZN(n13754) );
  INV_X1 U15760 ( .A(n13754), .ZN(P2_U3296) );
  NAND2_X1 U15761 ( .A1(n13756), .A2(n13755), .ZN(n13758) );
  OAI211_X1 U15762 ( .C1(n13764), .C2(n13759), .A(n13758), .B(n13757), .ZN(
        P2_U3299) );
  INV_X1 U15763 ( .A(n13760), .ZN(n14366) );
  OAI222_X1 U15764 ( .A1(n13764), .A2(n13762), .B1(n13766), .B2(n14366), .C1(
        P2_U3088), .C2(n13761), .ZN(P2_U3300) );
  INV_X1 U15765 ( .A(n13763), .ZN(n14369) );
  OAI222_X1 U15766 ( .A1(P2_U3088), .A2(n13767), .B1(n13766), .B2(n14369), 
        .C1(n13765), .C2(n13764), .ZN(P2_U3301) );
  INV_X1 U15767 ( .A(n13769), .ZN(n13770) );
  MUX2_X1 U15768 ( .A(n13770), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NOR2_X1 U15769 ( .A1(n14620), .A2(n13772), .ZN(n13775) );
  INV_X1 U15770 ( .A(n14058), .ZN(n14062) );
  OAI22_X1 U15771 ( .A1(n13925), .A2(n14062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13773), .ZN(n13774) );
  AOI211_X1 U15772 ( .C1(n8890), .C2(n13934), .A(n13775), .B(n13774), .ZN(
        n13776) );
  INV_X1 U15773 ( .A(n14258), .ZN(n14659) );
  OAI21_X1 U15774 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n13780) );
  NAND2_X1 U15775 ( .A1(n13780), .A2(n14612), .ZN(n13786) );
  NAND2_X1 U15776 ( .A1(n13942), .A2(n14222), .ZN(n14657) );
  INV_X1 U15777 ( .A(n13781), .ZN(n13782) );
  OAI21_X1 U15778 ( .B1(n13915), .B2(n14657), .A(n13782), .ZN(n13784) );
  NOR2_X1 U15779 ( .A1(n14620), .A2(n14252), .ZN(n13783) );
  AOI211_X1 U15780 ( .C1(n8890), .C2(n13944), .A(n13784), .B(n13783), .ZN(
        n13785) );
  OAI211_X1 U15781 ( .C1(n14659), .C2(n13921), .A(n13786), .B(n13785), .ZN(
        P1_U3215) );
  INV_X1 U15782 ( .A(n13787), .ZN(n13788) );
  NOR2_X1 U15783 ( .A1(n13789), .A2(n13788), .ZN(n13792) );
  INV_X1 U15784 ( .A(n13791), .ZN(n13863) );
  AOI21_X1 U15785 ( .B1(n13792), .B2(n13896), .A(n13863), .ZN(n13798) );
  NAND2_X1 U15786 ( .A1(n13938), .A2(n14221), .ZN(n13794) );
  NAND2_X1 U15787 ( .A1(n13936), .A2(n14222), .ZN(n13793) );
  NAND2_X1 U15788 ( .A1(n13794), .A2(n13793), .ZN(n14306) );
  AOI22_X1 U15789 ( .A1(n14614), .A2(n14306), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13795) );
  OAI21_X1 U15790 ( .B1(n14136), .B2(n14620), .A(n13795), .ZN(n13796) );
  AOI21_X1 U15791 ( .B1(n14307), .B2(n14616), .A(n13796), .ZN(n13797) );
  OAI21_X1 U15792 ( .B1(n13798), .B2(n13932), .A(n13797), .ZN(P1_U3216) );
  INV_X1 U15793 ( .A(n14332), .ZN(n14213) );
  NAND2_X1 U15794 ( .A1(n13901), .A2(n13902), .ZN(n13900) );
  INV_X1 U15795 ( .A(n13900), .ZN(n13801) );
  OAI21_X1 U15796 ( .B1(n13801), .B2(n13800), .A(n13799), .ZN(n13804) );
  NAND2_X1 U15797 ( .A1(n13900), .A2(n13802), .ZN(n13803) );
  NAND3_X1 U15798 ( .A1(n13804), .A2(n14612), .A3(n13803), .ZN(n13808) );
  NAND2_X1 U15799 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14026)
         );
  NAND2_X1 U15800 ( .A1(n8890), .A2(n13940), .ZN(n13805) );
  OAI211_X1 U15801 ( .C1(n14205), .C2(n13925), .A(n14026), .B(n13805), .ZN(
        n13806) );
  AOI21_X1 U15802 ( .B1(n14210), .B2(n13918), .A(n13806), .ZN(n13807) );
  OAI211_X1 U15803 ( .C1(n14213), .C2(n13921), .A(n13808), .B(n13807), .ZN(
        P1_U3219) );
  INV_X1 U15804 ( .A(n13809), .ZN(n13810) );
  AOI21_X1 U15805 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n13819) );
  INV_X1 U15806 ( .A(n14171), .ZN(n13816) );
  OR2_X1 U15807 ( .A1(n14205), .A2(n14631), .ZN(n13814) );
  NAND2_X1 U15808 ( .A1(n13938), .A2(n14222), .ZN(n13813) );
  NAND2_X1 U15809 ( .A1(n13814), .A2(n13813), .ZN(n14167) );
  AOI22_X1 U15810 ( .A1(n14167), .A2(n14614), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13815) );
  OAI21_X1 U15811 ( .B1(n13816), .B2(n14620), .A(n13815), .ZN(n13817) );
  AOI21_X1 U15812 ( .B1(n14319), .B2(n14616), .A(n13817), .ZN(n13818) );
  OAI21_X1 U15813 ( .B1(n13819), .B2(n13932), .A(n13818), .ZN(P1_U3223) );
  AND2_X1 U15814 ( .A1(n14609), .A2(n13820), .ZN(n13823) );
  OAI211_X1 U15815 ( .C1(n13823), .C2(n13822), .A(n14612), .B(n13821), .ZN(
        n13827) );
  OAI22_X1 U15816 ( .A1(n14249), .A2(n14633), .B1(n13824), .B2(n14631), .ZN(
        n14493) );
  AND2_X1 U15817 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14001) );
  NOR2_X1 U15818 ( .A1(n14620), .A2(n14497), .ZN(n13825) );
  AOI211_X1 U15819 ( .C1(n14614), .C2(n14493), .A(n14001), .B(n13825), .ZN(
        n13826) );
  OAI211_X1 U15820 ( .C1(n14506), .C2(n13921), .A(n13827), .B(n13826), .ZN(
        P1_U3224) );
  OAI22_X1 U15821 ( .A1(n13829), .A2(n14631), .B1(n13828), .B2(n14633), .ZN(
        n14104) );
  AOI22_X1 U15822 ( .A1(n14614), .A2(n14104), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13830) );
  OAI21_X1 U15823 ( .B1(n14111), .B2(n14620), .A(n13830), .ZN(n13838) );
  INV_X1 U15824 ( .A(n13832), .ZN(n13833) );
  NAND3_X1 U15825 ( .A1(n13831), .A2(n13834), .A3(n13833), .ZN(n13835) );
  AOI21_X1 U15826 ( .B1(n13836), .B2(n13835), .A(n13932), .ZN(n13837) );
  AOI211_X1 U15827 ( .C1(n14293), .C2(n14616), .A(n13838), .B(n13837), .ZN(
        n13839) );
  INV_X1 U15828 ( .A(n13839), .ZN(P1_U3225) );
  INV_X1 U15829 ( .A(n13840), .ZN(n13852) );
  AOI21_X1 U15830 ( .B1(n13842), .B2(n13841), .A(n13852), .ZN(n13848) );
  OAI21_X1 U15831 ( .B1(n13925), .B2(n14632), .A(n13843), .ZN(n13844) );
  AOI21_X1 U15832 ( .B1(n8890), .B2(n13942), .A(n13844), .ZN(n13845) );
  OAI21_X1 U15833 ( .B1(n14641), .B2(n14620), .A(n13845), .ZN(n13846) );
  AOI21_X1 U15834 ( .B1(n14645), .B2(n14616), .A(n13846), .ZN(n13847) );
  OAI21_X1 U15835 ( .B1(n13848), .B2(n13932), .A(n13847), .ZN(P1_U3226) );
  INV_X1 U15836 ( .A(n13849), .ZN(n13851) );
  NOR3_X1 U15837 ( .A1(n13852), .A2(n13851), .A3(n13850), .ZN(n13855) );
  INV_X1 U15838 ( .A(n13853), .ZN(n13854) );
  OAI21_X1 U15839 ( .B1(n13855), .B2(n13854), .A(n14612), .ZN(n13860) );
  AND2_X1 U15840 ( .A1(n13941), .A2(n14221), .ZN(n13856) );
  AOI21_X1 U15841 ( .B1(n13940), .B2(n14222), .A(n13856), .ZN(n14340) );
  OAI21_X1 U15842 ( .B1(n14340), .B2(n13915), .A(n13857), .ZN(n13858) );
  AOI21_X1 U15843 ( .B1(n14238), .B2(n13918), .A(n13858), .ZN(n13859) );
  OAI211_X1 U15844 ( .C1(n14240), .C2(n13921), .A(n13860), .B(n13859), .ZN(
        P1_U3228) );
  NOR3_X1 U15845 ( .A1(n13863), .A2(n7624), .A3(n13862), .ZN(n13865) );
  INV_X1 U15846 ( .A(n13831), .ZN(n13864) );
  OAI21_X1 U15847 ( .B1(n13865), .B2(n13864), .A(n14612), .ZN(n13869) );
  INV_X1 U15848 ( .A(n13866), .ZN(n14129) );
  AOI22_X1 U15849 ( .A1(n14221), .A2(n13937), .B1(n13935), .B2(n14222), .ZN(
        n14119) );
  OAI22_X1 U15850 ( .A1(n13915), .A2(n14119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15270), .ZN(n13867) );
  AOI21_X1 U15851 ( .B1(n13918), .B2(n14129), .A(n13867), .ZN(n13868) );
  OAI211_X1 U15852 ( .C1(n14132), .C2(n13921), .A(n13869), .B(n13868), .ZN(
        P1_U3229) );
  XNOR2_X1 U15853 ( .A(n13871), .B(n13870), .ZN(n13878) );
  INV_X1 U15854 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15397) );
  OAI22_X1 U15855 ( .A1(n13890), .A2(n13925), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15397), .ZN(n13872) );
  AOI21_X1 U15856 ( .B1(n8890), .B2(n14223), .A(n13872), .ZN(n13873) );
  OAI21_X1 U15857 ( .B1(n13874), .B2(n14620), .A(n13873), .ZN(n13875) );
  AOI21_X1 U15858 ( .B1(n13876), .B2(n14616), .A(n13875), .ZN(n13877) );
  OAI21_X1 U15859 ( .B1(n13878), .B2(n13932), .A(n13877), .ZN(P1_U3233) );
  XNOR2_X1 U15860 ( .A(n13880), .B(n13879), .ZN(n13888) );
  OAI21_X1 U15861 ( .B1(n13925), .B2(n13882), .A(n13881), .ZN(n13883) );
  AOI21_X1 U15862 ( .B1(n8890), .B2(n13945), .A(n13883), .ZN(n13884) );
  OAI21_X1 U15863 ( .B1(n13885), .B2(n14620), .A(n13884), .ZN(n13886) );
  AOI21_X1 U15864 ( .B1(n14666), .B2(n14616), .A(n13886), .ZN(n13887) );
  OAI21_X1 U15865 ( .B1(n13888), .B2(n13932), .A(n13887), .ZN(P1_U3234) );
  OAI22_X1 U15866 ( .A1(n13890), .A2(n14631), .B1(n13889), .B2(n14633), .ZN(
        n14153) );
  AOI22_X1 U15867 ( .A1(n14153), .A2(n14614), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13891) );
  OAI21_X1 U15868 ( .B1(n14156), .B2(n14620), .A(n13891), .ZN(n13898) );
  INV_X1 U15869 ( .A(n13892), .ZN(n13893) );
  NAND3_X1 U15870 ( .A1(n13809), .A2(n13894), .A3(n13893), .ZN(n13895) );
  AOI21_X1 U15871 ( .B1(n13896), .B2(n13895), .A(n13932), .ZN(n13897) );
  AOI211_X1 U15872 ( .C1(n14314), .C2(n14616), .A(n13898), .B(n13897), .ZN(
        n13899) );
  INV_X1 U15873 ( .A(n13899), .ZN(P1_U3235) );
  INV_X1 U15874 ( .A(n14337), .ZN(n14231) );
  OAI21_X1 U15875 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13903) );
  NAND2_X1 U15876 ( .A1(n13903), .A2(n14612), .ZN(n13909) );
  NOR2_X1 U15877 ( .A1(n14620), .A2(n14227), .ZN(n13907) );
  OAI21_X1 U15878 ( .B1(n13925), .B2(n13905), .A(n13904), .ZN(n13906) );
  AOI211_X1 U15879 ( .C1(n8890), .C2(n14220), .A(n13907), .B(n13906), .ZN(
        n13908) );
  OAI211_X1 U15880 ( .C1(n14231), .C2(n13921), .A(n13909), .B(n13908), .ZN(
        P1_U3238) );
  OAI21_X1 U15881 ( .B1(n13912), .B2(n13911), .A(n13910), .ZN(n13913) );
  NAND2_X1 U15882 ( .A1(n13913), .A2(n14612), .ZN(n13920) );
  INV_X1 U15883 ( .A(n14093), .ZN(n13917) );
  AOI22_X1 U15884 ( .A1(n14068), .A2(n14222), .B1(n14221), .B2(n13935), .ZN(
        n14090) );
  OAI22_X1 U15885 ( .A1(n13915), .A2(n14090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13914), .ZN(n13916) );
  AOI21_X1 U15886 ( .B1(n13918), .B2(n13917), .A(n13916), .ZN(n13919) );
  OAI211_X1 U15887 ( .C1(n14097), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        P1_U3240) );
  XNOR2_X1 U15888 ( .A(n13923), .B(n13922), .ZN(n13933) );
  NAND2_X1 U15889 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14730)
         );
  OAI21_X1 U15890 ( .B1(n13925), .B2(n13924), .A(n14730), .ZN(n13926) );
  AOI21_X1 U15891 ( .B1(n8890), .B2(n13943), .A(n13926), .ZN(n13927) );
  OAI21_X1 U15892 ( .B1(n13928), .B2(n14620), .A(n13927), .ZN(n13929) );
  AOI21_X1 U15893 ( .B1(n13930), .B2(n14616), .A(n13929), .ZN(n13931) );
  OAI21_X1 U15894 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(P1_U3241) );
  MUX2_X1 U15895 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14031), .S(n13956), .Z(
        P1_U3591) );
  MUX2_X1 U15896 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14047), .S(n13956), .Z(
        P1_U3590) );
  MUX2_X1 U15897 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14069), .S(n13956), .Z(
        P1_U3589) );
  MUX2_X1 U15898 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14058), .S(n13956), .Z(
        P1_U3588) );
  MUX2_X1 U15899 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14068), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15900 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13934), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15901 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13935), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15902 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13936), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15903 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13937), .S(n13956), .Z(
        P1_U3583) );
  MUX2_X1 U15904 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13938), .S(n13956), .Z(
        P1_U3582) );
  MUX2_X1 U15905 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14183), .S(n13956), .Z(
        P1_U3581) );
  MUX2_X1 U15906 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13939), .S(n13956), .Z(
        P1_U3580) );
  MUX2_X1 U15907 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14223), .S(n13956), .Z(
        P1_U3579) );
  MUX2_X1 U15908 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13940), .S(n13956), .Z(
        P1_U3578) );
  MUX2_X1 U15909 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14220), .S(n13956), .Z(
        P1_U3577) );
  MUX2_X1 U15910 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13941), .S(n13956), .Z(
        P1_U3576) );
  MUX2_X1 U15911 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13942), .S(n13956), .Z(
        P1_U3575) );
  MUX2_X1 U15912 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13943), .S(n13956), .Z(
        P1_U3574) );
  MUX2_X1 U15913 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13944), .S(n13956), .Z(
        P1_U3573) );
  MUX2_X1 U15914 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13945), .S(n13956), .Z(
        P1_U3572) );
  MUX2_X1 U15915 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13946), .S(n13956), .Z(
        P1_U3571) );
  MUX2_X1 U15916 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13947), .S(n13956), .Z(
        P1_U3570) );
  MUX2_X1 U15917 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13948), .S(n13956), .Z(
        P1_U3569) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13949), .S(n13956), .Z(
        P1_U3568) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13950), .S(n13956), .Z(
        P1_U3567) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13951), .S(n13956), .Z(
        P1_U3566) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13952), .S(n13956), .Z(
        P1_U3565) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n7323), .S(n13956), .Z(
        P1_U3564) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13953), .S(n13956), .Z(
        P1_U3563) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13954), .S(n13956), .Z(
        P1_U3562) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13955), .S(n13956), .Z(
        P1_U3561) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13957), .S(n13956), .Z(
        P1_U3560) );
  INV_X1 U15927 ( .A(n14020), .ZN(n14724) );
  OAI22_X1 U15928 ( .A1(n14732), .A2(n14378), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13958), .ZN(n13959) );
  AOI21_X1 U15929 ( .B1(n13960), .B2(n14724), .A(n13959), .ZN(n13970) );
  AND2_X1 U15930 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13962) );
  OAI211_X1 U15931 ( .C1(n13963), .C2(n13962), .A(n14727), .B(n13961), .ZN(
        n13969) );
  INV_X1 U15932 ( .A(n13964), .ZN(n13967) );
  OAI211_X1 U15933 ( .C1(n13967), .C2(n13966), .A(n14728), .B(n13965), .ZN(
        n13968) );
  NAND3_X1 U15934 ( .A1(n13970), .A2(n13969), .A3(n13968), .ZN(P1_U3244) );
  OAI22_X1 U15935 ( .A1(n14732), .A2(n14379), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9792), .ZN(n13971) );
  AOI21_X1 U15936 ( .B1(n13972), .B2(n14724), .A(n13971), .ZN(n13980) );
  OAI211_X1 U15937 ( .C1(n13974), .C2(n13973), .A(n14728), .B(n13990), .ZN(
        n13979) );
  OAI211_X1 U15938 ( .C1(n13977), .C2(n13976), .A(n14727), .B(n13975), .ZN(
        n13978) );
  NAND4_X1 U15939 ( .A1(n13981), .A2(n13980), .A3(n13979), .A4(n13978), .ZN(
        P1_U3245) );
  NOR2_X1 U15940 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14734), .ZN(n13984) );
  NOR2_X1 U15941 ( .A1(n14020), .A2(n13982), .ZN(n13983) );
  AOI211_X1 U15942 ( .C1(n14715), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13984), .B(
        n13983), .ZN(n13996) );
  OAI211_X1 U15943 ( .C1(n13987), .C2(n13986), .A(n14727), .B(n13985), .ZN(
        n13995) );
  MUX2_X1 U15944 ( .A(n9022), .B(P1_REG2_REG_3__SCAN_IN), .S(n13988), .Z(
        n13991) );
  NAND3_X1 U15945 ( .A1(n13991), .A2(n13990), .A3(n13989), .ZN(n13992) );
  NAND3_X1 U15946 ( .A1(n14728), .A2(n13993), .A3(n13992), .ZN(n13994) );
  NAND3_X1 U15947 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(P1_U3246) );
  OAI21_X1 U15948 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14000) );
  NAND2_X1 U15949 ( .A1(n14000), .A2(n14727), .ZN(n14010) );
  AOI21_X1 U15950 ( .B1(n14715), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14001), 
        .ZN(n14009) );
  OAI21_X1 U15951 ( .B1(n14004), .B2(n14003), .A(n14002), .ZN(n14005) );
  NAND2_X1 U15952 ( .A1(n14005), .A2(n14728), .ZN(n14008) );
  NAND2_X1 U15953 ( .A1(n14724), .A2(n14006), .ZN(n14007) );
  NAND4_X1 U15954 ( .A1(n14010), .A2(n14009), .A3(n14008), .A4(n14007), .ZN(
        P1_U3255) );
  NAND2_X1 U15955 ( .A1(n14012), .A2(n14011), .ZN(n14016) );
  INV_X1 U15956 ( .A(n14013), .ZN(n14014) );
  NAND2_X1 U15957 ( .A1(n14014), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14015) );
  NAND2_X1 U15958 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  XOR2_X1 U15959 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14017), .Z(n14023) );
  XNOR2_X1 U15960 ( .A(n14019), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U15961 ( .A1(n14023), .A2(n14728), .B1(n14727), .B2(n14022), .ZN(
        n14024) );
  MUX2_X1 U15962 ( .A(n14025), .B(n14024), .S(n14635), .Z(n14027) );
  OAI211_X1 U15963 ( .C1(n7728), .C2(n14732), .A(n14027), .B(n14026), .ZN(
        P1_U3262) );
  NAND2_X1 U15964 ( .A1(n14028), .A2(n8808), .ZN(n14266) );
  INV_X1 U15965 ( .A(P1_B_REG_SCAN_IN), .ZN(n14029) );
  NOR2_X1 U15966 ( .A1(n6526), .A2(n14029), .ZN(n14030) );
  NOR2_X1 U15967 ( .A1(n14633), .A2(n14030), .ZN(n14048) );
  NAND2_X1 U15968 ( .A1(n14031), .A2(n14048), .ZN(n14268) );
  NOR2_X1 U15969 ( .A1(n14747), .A2(n14268), .ZN(n14038) );
  INV_X1 U15970 ( .A(n14032), .ZN(n14267) );
  NOR2_X1 U15971 ( .A1(n14267), .A2(n14738), .ZN(n14033) );
  AOI211_X1 U15972 ( .C1(n14747), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14038), 
        .B(n14033), .ZN(n14034) );
  OAI21_X1 U15973 ( .B1(n14266), .B2(n14489), .A(n14034), .ZN(P1_U3263) );
  OAI211_X1 U15974 ( .C1(n14270), .C2(n6820), .A(n14036), .B(n8808), .ZN(
        n14269) );
  AND2_X1 U15975 ( .A1(n14747), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14037) );
  NOR2_X1 U15976 ( .A1(n14038), .A2(n14037), .ZN(n14041) );
  NAND2_X1 U15977 ( .A1(n14039), .A2(n14259), .ZN(n14040) );
  OAI211_X1 U15978 ( .C1(n14269), .C2(n14489), .A(n14041), .B(n14040), .ZN(
        P1_U3264) );
  NAND2_X1 U15979 ( .A1(n14074), .A2(n14043), .ZN(n14044) );
  XNOR2_X1 U15980 ( .A(n14044), .B(n14060), .ZN(n14274) );
  AOI21_X1 U15981 ( .B1(n14273), .B2(n6584), .A(n14674), .ZN(n14046) );
  NAND2_X1 U15982 ( .A1(n14046), .A2(n14045), .ZN(n14275) );
  AND2_X1 U15983 ( .A1(n14048), .A2(n14047), .ZN(n14271) );
  INV_X1 U15984 ( .A(n14271), .ZN(n14050) );
  OAI22_X1 U15985 ( .A1(n14051), .A2(n14050), .B1(n14049), .B2(n14642), .ZN(
        n14052) );
  AOI21_X1 U15986 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14747), .A(n14052), 
        .ZN(n14054) );
  NAND2_X1 U15987 ( .A1(n14273), .A2(n14259), .ZN(n14053) );
  OAI211_X1 U15988 ( .C1(n14275), .C2(n14489), .A(n14054), .B(n14053), .ZN(
        n14065) );
  XOR2_X1 U15989 ( .A(n14060), .B(n14059), .Z(n14061) );
  NAND2_X1 U15990 ( .A1(n14061), .A2(n14494), .ZN(n14278) );
  NOR2_X1 U15991 ( .A1(n14062), .A2(n14631), .ZN(n14272) );
  INV_X1 U15992 ( .A(n14272), .ZN(n14063) );
  AOI21_X1 U15993 ( .B1(n14278), .B2(n14063), .A(n14747), .ZN(n14064) );
  INV_X1 U15994 ( .A(n14066), .ZN(P1_U3356) );
  NAND2_X1 U15995 ( .A1(n14068), .A2(n14221), .ZN(n14071) );
  NAND2_X1 U15996 ( .A1(n14069), .A2(n14222), .ZN(n14070) );
  OAI21_X1 U15997 ( .B1(n14076), .B2(n14075), .A(n14074), .ZN(n14283) );
  NAND2_X1 U15998 ( .A1(n14747), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14077) );
  OAI21_X1 U15999 ( .B1(n14642), .B2(n14078), .A(n14077), .ZN(n14079) );
  AOI21_X1 U16000 ( .B1(n14280), .B2(n14259), .A(n14079), .ZN(n14083) );
  AOI21_X1 U16001 ( .B1(n14280), .B2(n14080), .A(n14674), .ZN(n14081) );
  NAND2_X1 U16002 ( .A1(n14279), .A2(n14743), .ZN(n14082) );
  OAI211_X1 U16003 ( .C1(n14283), .C2(n14247), .A(n14083), .B(n14082), .ZN(
        n14084) );
  INV_X1 U16004 ( .A(n14084), .ZN(n14085) );
  OAI21_X1 U16005 ( .B1(n14282), .B2(n14747), .A(n14085), .ZN(P1_U3265) );
  OAI21_X1 U16006 ( .B1(n7419), .B2(n14087), .A(n14086), .ZN(n14292) );
  XNOR2_X1 U16007 ( .A(n14089), .B(n14088), .ZN(n14092) );
  INV_X1 U16008 ( .A(n14090), .ZN(n14091) );
  AOI21_X1 U16009 ( .B1(n14092), .B2(n14494), .A(n14091), .ZN(n14291) );
  OAI21_X1 U16010 ( .B1(n14093), .B2(n14642), .A(n14291), .ZN(n14094) );
  NAND2_X1 U16011 ( .A1(n14094), .A2(n14639), .ZN(n14100) );
  AOI211_X1 U16012 ( .C1(n14289), .C2(n14106), .A(n14674), .B(n14095), .ZN(
        n14288) );
  OAI22_X1 U16013 ( .A1(n14097), .A2(n14738), .B1(n14096), .B2(n14639), .ZN(
        n14098) );
  AOI21_X1 U16014 ( .B1(n14288), .B2(n14743), .A(n14098), .ZN(n14099) );
  OAI211_X1 U16015 ( .C1(n14292), .C2(n14247), .A(n14100), .B(n14099), .ZN(
        P1_U3267) );
  OAI21_X1 U16016 ( .B1(n14103), .B2(n14102), .A(n14101), .ZN(n14105) );
  AOI21_X1 U16017 ( .B1(n14105), .B2(n14494), .A(n14104), .ZN(n14299) );
  OAI211_X1 U16018 ( .C1(n14107), .C2(n14128), .A(n8808), .B(n14106), .ZN(
        n14296) );
  OR2_X1 U16019 ( .A1(n14109), .A2(n14108), .ZN(n14295) );
  NAND3_X1 U16020 ( .A1(n14295), .A2(n14262), .A3(n14294), .ZN(n14114) );
  NAND2_X1 U16021 ( .A1(n14747), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U16022 ( .B1(n14642), .B2(n14111), .A(n14110), .ZN(n14112) );
  AOI21_X1 U16023 ( .B1(n14293), .B2(n14259), .A(n14112), .ZN(n14113) );
  OAI211_X1 U16024 ( .C1(n14296), .C2(n14489), .A(n14114), .B(n14113), .ZN(
        n14115) );
  INV_X1 U16025 ( .A(n14115), .ZN(n14116) );
  OAI21_X1 U16026 ( .B1(n14299), .B2(n14747), .A(n14116), .ZN(P1_U3268) );
  AOI211_X1 U16027 ( .C1(n11714), .C2(n14118), .A(n14629), .B(n14117), .ZN(
        n14121) );
  INV_X1 U16028 ( .A(n14119), .ZN(n14120) );
  NOR2_X1 U16029 ( .A1(n14121), .A2(n14120), .ZN(n14303) );
  INV_X1 U16030 ( .A(n14122), .ZN(n14123) );
  AOI21_X1 U16031 ( .B1(n14125), .B2(n14124), .A(n14123), .ZN(n14304) );
  INV_X1 U16032 ( .A(n14304), .ZN(n14134) );
  NAND2_X1 U16033 ( .A1(n14301), .A2(n6588), .ZN(n14126) );
  NAND2_X1 U16034 ( .A1(n14126), .A2(n8808), .ZN(n14127) );
  NOR2_X1 U16035 ( .A1(n14128), .A2(n14127), .ZN(n14300) );
  NAND2_X1 U16036 ( .A1(n14300), .A2(n14743), .ZN(n14131) );
  AOI22_X1 U16037 ( .A1(n14747), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14129), 
        .B2(n14735), .ZN(n14130) );
  OAI211_X1 U16038 ( .C1(n14132), .C2(n14738), .A(n14131), .B(n14130), .ZN(
        n14133) );
  AOI21_X1 U16039 ( .B1(n14134), .B2(n14262), .A(n14133), .ZN(n14135) );
  OAI21_X1 U16040 ( .B1(n14303), .B2(n14747), .A(n14135), .ZN(P1_U3269) );
  INV_X1 U16041 ( .A(n14136), .ZN(n14141) );
  XNOR2_X1 U16042 ( .A(n14138), .B(n14137), .ZN(n14139) );
  NAND2_X1 U16043 ( .A1(n14139), .A2(n14494), .ZN(n14312) );
  INV_X1 U16044 ( .A(n14312), .ZN(n14140) );
  AOI211_X1 U16045 ( .C1(n14735), .C2(n14141), .A(n14306), .B(n14140), .ZN(
        n14148) );
  INV_X1 U16046 ( .A(n6588), .ZN(n14142) );
  AOI211_X1 U16047 ( .C1(n14307), .C2(n6681), .A(n14674), .B(n14142), .ZN(
        n14305) );
  OAI22_X1 U16048 ( .A1(n7499), .A2(n14738), .B1(n15417), .B2(n14639), .ZN(
        n14143) );
  AOI21_X1 U16049 ( .B1(n14305), .B2(n14743), .A(n14143), .ZN(n14147) );
  NAND2_X1 U16050 ( .A1(n14145), .A2(n14144), .ZN(n14308) );
  NAND3_X1 U16051 ( .A1(n14309), .A2(n14308), .A3(n14262), .ZN(n14146) );
  OAI211_X1 U16052 ( .C1(n14148), .C2(n14747), .A(n14147), .B(n14146), .ZN(
        P1_U3270) );
  XOR2_X1 U16053 ( .A(n14149), .B(n14150), .Z(n14317) );
  OAI21_X1 U16054 ( .B1(n14166), .B2(n14151), .A(n14150), .ZN(n14152) );
  AOI21_X1 U16055 ( .B1(n6617), .B2(n14152), .A(n14629), .ZN(n14154) );
  NOR2_X1 U16056 ( .A1(n14154), .A2(n14153), .ZN(n14316) );
  NAND2_X1 U16057 ( .A1(n14747), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n14155) );
  OAI21_X1 U16058 ( .B1(n14642), .B2(n14156), .A(n14155), .ZN(n14157) );
  AOI21_X1 U16059 ( .B1(n14314), .B2(n14259), .A(n14157), .ZN(n14160) );
  AOI21_X1 U16060 ( .B1(n14314), .B2(n14169), .A(n14674), .ZN(n14158) );
  AND2_X1 U16061 ( .A1(n14158), .A2(n6681), .ZN(n14313) );
  NAND2_X1 U16062 ( .A1(n14313), .A2(n14743), .ZN(n14159) );
  OAI211_X1 U16063 ( .C1(n14316), .C2(n14747), .A(n14160), .B(n14159), .ZN(
        n14161) );
  INV_X1 U16064 ( .A(n14161), .ZN(n14162) );
  OAI21_X1 U16065 ( .B1(n14317), .B2(n14247), .A(n14162), .ZN(P1_U3271) );
  AND3_X1 U16066 ( .A1(n14180), .A2(n14164), .A3(n14163), .ZN(n14165) );
  NOR3_X1 U16067 ( .A1(n14166), .A2(n14165), .A3(n14629), .ZN(n14168) );
  NOR2_X1 U16068 ( .A1(n14168), .A2(n14167), .ZN(n14321) );
  INV_X1 U16069 ( .A(n14169), .ZN(n14170) );
  AOI211_X1 U16070 ( .C1(n14319), .C2(n14188), .A(n14674), .B(n14170), .ZN(
        n14318) );
  INV_X1 U16071 ( .A(n14319), .ZN(n14173) );
  AOI22_X1 U16072 ( .A1(n14171), .A2(n14735), .B1(n14747), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14172) );
  OAI21_X1 U16073 ( .B1(n14173), .B2(n14738), .A(n14172), .ZN(n14178) );
  INV_X1 U16074 ( .A(n14174), .ZN(n14175) );
  AOI21_X1 U16075 ( .B1(n7398), .B2(n14176), .A(n14175), .ZN(n14322) );
  NOR2_X1 U16076 ( .A1(n14322), .A2(n14247), .ZN(n14177) );
  AOI211_X1 U16077 ( .C1(n14318), .C2(n14743), .A(n14178), .B(n14177), .ZN(
        n14179) );
  OAI21_X1 U16078 ( .B1(n14747), .B2(n14321), .A(n14179), .ZN(P1_U3272) );
  OAI211_X1 U16079 ( .C1(n14182), .C2(n14181), .A(n14180), .B(n14494), .ZN(
        n14185) );
  AOI22_X1 U16080 ( .A1(n14183), .A2(n14222), .B1(n14223), .B2(n14221), .ZN(
        n14184) );
  NAND2_X1 U16081 ( .A1(n14185), .A2(n14184), .ZN(n14329) );
  AOI21_X1 U16082 ( .B1(n14186), .B2(n14735), .A(n14329), .ZN(n14198) );
  OR2_X1 U16083 ( .A1(n14209), .A2(n14325), .ZN(n14187) );
  NAND2_X1 U16084 ( .A1(n14188), .A2(n14187), .ZN(n14326) );
  INV_X1 U16085 ( .A(n14326), .ZN(n14196) );
  INV_X1 U16086 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U16087 ( .A1(n14325), .A2(n14738), .B1(n14639), .B2(n14189), .ZN(
        n14194) );
  NOR2_X1 U16088 ( .A1(n14191), .A2(n14190), .ZN(n14324) );
  INV_X1 U16089 ( .A(n14192), .ZN(n14323) );
  NOR3_X1 U16090 ( .A1(n14324), .A2(n14323), .A3(n14247), .ZN(n14193) );
  AOI211_X1 U16091 ( .C1(n14196), .C2(n14195), .A(n14194), .B(n14193), .ZN(
        n14197) );
  OAI21_X1 U16092 ( .B1(n14198), .B2(n14747), .A(n14197), .ZN(P1_U3273) );
  XNOR2_X1 U16093 ( .A(n14200), .B(n14199), .ZN(n14334) );
  AOI21_X1 U16094 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14204) );
  OAI222_X1 U16095 ( .A1(n14631), .A2(n14206), .B1(n14633), .B2(n14205), .C1(
        n14629), .C2(n14204), .ZN(n14330) );
  NAND2_X1 U16096 ( .A1(n14332), .A2(n14226), .ZN(n14207) );
  NAND2_X1 U16097 ( .A1(n14207), .A2(n8808), .ZN(n14208) );
  NOR2_X1 U16098 ( .A1(n14209), .A2(n14208), .ZN(n14331) );
  NAND2_X1 U16099 ( .A1(n14331), .A2(n14743), .ZN(n14212) );
  AOI22_X1 U16100 ( .A1(n14747), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14210), 
        .B2(n14735), .ZN(n14211) );
  OAI211_X1 U16101 ( .C1(n14213), .C2(n14738), .A(n14212), .B(n14211), .ZN(
        n14214) );
  AOI21_X1 U16102 ( .B1(n14330), .B2(n14639), .A(n14214), .ZN(n14215) );
  OAI21_X1 U16103 ( .B1(n14334), .B2(n14247), .A(n14215), .ZN(P1_U3274) );
  XOR2_X1 U16104 ( .A(n14216), .B(n14218), .Z(n14339) );
  OAI211_X1 U16105 ( .C1(n14219), .C2(n14218), .A(n14217), .B(n14494), .ZN(
        n14225) );
  AOI22_X1 U16106 ( .A1(n14223), .A2(n14222), .B1(n14221), .B2(n14220), .ZN(
        n14224) );
  NAND2_X1 U16107 ( .A1(n14225), .A2(n14224), .ZN(n14335) );
  AOI211_X1 U16108 ( .C1(n14337), .C2(n14235), .A(n14674), .B(n6813), .ZN(
        n14336) );
  NAND2_X1 U16109 ( .A1(n14336), .A2(n14743), .ZN(n14230) );
  INV_X1 U16110 ( .A(n14227), .ZN(n14228) );
  AOI22_X1 U16111 ( .A1(n14747), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14228), 
        .B2(n14735), .ZN(n14229) );
  OAI211_X1 U16112 ( .C1(n14231), .C2(n14738), .A(n14230), .B(n14229), .ZN(
        n14232) );
  AOI21_X1 U16113 ( .B1(n14335), .B2(n14639), .A(n14232), .ZN(n14233) );
  OAI21_X1 U16114 ( .B1(n14247), .B2(n14339), .A(n14233), .ZN(P1_U3275) );
  XNOR2_X1 U16115 ( .A(n14234), .B(n14241), .ZN(n14346) );
  INV_X1 U16116 ( .A(n14622), .ZN(n14237) );
  INV_X1 U16117 ( .A(n14235), .ZN(n14236) );
  AOI211_X1 U16118 ( .C1(n14343), .C2(n14237), .A(n14674), .B(n14236), .ZN(
        n14341) );
  AOI22_X1 U16119 ( .A1(n14747), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14238), 
        .B2(n14735), .ZN(n14239) );
  OAI21_X1 U16120 ( .B1(n14240), .B2(n14738), .A(n14239), .ZN(n14245) );
  XNOR2_X1 U16121 ( .A(n14242), .B(n14241), .ZN(n14243) );
  NAND2_X1 U16122 ( .A1(n14243), .A2(n14494), .ZN(n14344) );
  AOI21_X1 U16123 ( .B1(n14344), .B2(n14340), .A(n14747), .ZN(n14244) );
  AOI211_X1 U16124 ( .C1(n14341), .C2(n14743), .A(n14245), .B(n14244), .ZN(
        n14246) );
  OAI21_X1 U16125 ( .B1(n14247), .B2(n14346), .A(n14246), .ZN(P1_U3276) );
  XNOR2_X1 U16126 ( .A(n14248), .B(n14260), .ZN(n14250) );
  OAI22_X1 U16127 ( .A1(n14250), .A2(n14629), .B1(n14249), .B2(n14631), .ZN(
        n14662) );
  INV_X1 U16128 ( .A(n14657), .ZN(n14251) );
  OAI21_X1 U16129 ( .B1(n14662), .B2(n14251), .A(n14639), .ZN(n14265) );
  OAI22_X1 U16130 ( .A1(n14639), .A2(n9693), .B1(n14252), .B2(n14642), .ZN(
        n14257) );
  INV_X1 U16131 ( .A(n14253), .ZN(n14255) );
  OAI211_X1 U16132 ( .C1(n14659), .C2(n14255), .A(n8808), .B(n14254), .ZN(
        n14658) );
  NOR2_X1 U16133 ( .A1(n14658), .A2(n14489), .ZN(n14256) );
  AOI211_X1 U16134 ( .C1(n14259), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14264) );
  NAND2_X1 U16135 ( .A1(n14261), .A2(n14260), .ZN(n14655) );
  NAND3_X1 U16136 ( .A1(n6959), .A2(n14655), .A3(n14262), .ZN(n14263) );
  NAND3_X1 U16137 ( .A1(n14265), .A2(n14264), .A3(n14263), .ZN(P1_U3279) );
  OAI211_X1 U16138 ( .C1(n14267), .C2(n14793), .A(n14266), .B(n14268), .ZN(
        n14348) );
  MUX2_X1 U16139 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14348), .S(n14808), .Z(
        P1_U3559) );
  MUX2_X1 U16140 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14349), .S(n14808), .Z(
        P1_U3558) );
  AOI211_X1 U16141 ( .C1(n14273), .C2(n14759), .A(n14272), .B(n14271), .ZN(
        n14277) );
  NAND2_X1 U16142 ( .A1(n14274), .A2(n14796), .ZN(n14276) );
  NAND4_X1 U16143 ( .A1(n14276), .A2(n14277), .A3(n14278), .A4(n14275), .ZN(
        n14350) );
  MUX2_X1 U16144 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14350), .S(n14808), .Z(
        P1_U3557) );
  AOI21_X1 U16145 ( .B1(n14759), .B2(n14280), .A(n14279), .ZN(n14281) );
  MUX2_X1 U16146 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14351), .S(n14808), .Z(
        P1_U3556) );
  AOI22_X1 U16147 ( .A1(n14285), .A2(n8808), .B1(n14759), .B2(n14284), .ZN(
        n14286) );
  MUX2_X1 U16148 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14352), .S(n14808), .Z(
        P1_U3555) );
  AOI21_X1 U16149 ( .B1(n14759), .B2(n14289), .A(n14288), .ZN(n14290) );
  OAI211_X1 U16150 ( .C1(n14663), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14353) );
  MUX2_X1 U16151 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14353), .S(n14808), .Z(
        P1_U3554) );
  NAND2_X1 U16152 ( .A1(n14293), .A2(n14759), .ZN(n14298) );
  NAND3_X1 U16153 ( .A1(n14295), .A2(n14796), .A3(n14294), .ZN(n14297) );
  NAND4_X1 U16154 ( .A1(n14299), .A2(n14298), .A3(n14297), .A4(n14296), .ZN(
        n14354) );
  MUX2_X1 U16155 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14354), .S(n14808), .Z(
        P1_U3553) );
  AOI21_X1 U16156 ( .B1(n14759), .B2(n14301), .A(n14300), .ZN(n14302) );
  OAI211_X1 U16157 ( .C1(n14663), .C2(n14304), .A(n14303), .B(n14302), .ZN(
        n14355) );
  MUX2_X1 U16158 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14355), .S(n14808), .Z(
        P1_U3552) );
  AOI211_X1 U16159 ( .C1(n14759), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        n14311) );
  NAND3_X1 U16160 ( .A1(n14309), .A2(n14308), .A3(n14796), .ZN(n14310) );
  NAND3_X1 U16161 ( .A1(n14312), .A2(n14311), .A3(n14310), .ZN(n14356) );
  MUX2_X1 U16162 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14356), .S(n14808), .Z(
        P1_U3551) );
  AOI21_X1 U16163 ( .B1(n14759), .B2(n14314), .A(n14313), .ZN(n14315) );
  OAI211_X1 U16164 ( .C1(n14663), .C2(n14317), .A(n14316), .B(n14315), .ZN(
        n14357) );
  MUX2_X1 U16165 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14357), .S(n14808), .Z(
        P1_U3550) );
  AOI21_X1 U16166 ( .B1(n14759), .B2(n14319), .A(n14318), .ZN(n14320) );
  OAI211_X1 U16167 ( .C1(n14663), .C2(n14322), .A(n14321), .B(n14320), .ZN(
        n14358) );
  MUX2_X1 U16168 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14358), .S(n14808), .Z(
        P1_U3549) );
  NOR3_X1 U16169 ( .A1(n14324), .A2(n14323), .A3(n14663), .ZN(n14328) );
  OAI22_X1 U16170 ( .A1(n14326), .A2(n14674), .B1(n14325), .B2(n14793), .ZN(
        n14327) );
  MUX2_X1 U16171 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14359), .S(n14808), .Z(
        P1_U3548) );
  AOI211_X1 U16172 ( .C1(n14759), .C2(n14332), .A(n14331), .B(n14330), .ZN(
        n14333) );
  OAI21_X1 U16173 ( .B1(n14663), .B2(n14334), .A(n14333), .ZN(n14360) );
  MUX2_X1 U16174 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14360), .S(n14808), .Z(
        P1_U3547) );
  AOI211_X1 U16175 ( .C1(n14759), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        n14338) );
  OAI21_X1 U16176 ( .B1(n14663), .B2(n14339), .A(n14338), .ZN(n14361) );
  MUX2_X1 U16177 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14361), .S(n14808), .Z(
        P1_U3546) );
  INV_X1 U16178 ( .A(n14340), .ZN(n14342) );
  AOI211_X1 U16179 ( .C1(n14759), .C2(n14343), .A(n14342), .B(n14341), .ZN(
        n14345) );
  OAI211_X1 U16180 ( .C1(n14663), .C2(n14346), .A(n14345), .B(n14344), .ZN(
        n14362) );
  MUX2_X1 U16181 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14362), .S(n14808), .Z(
        P1_U3545) );
  MUX2_X1 U16182 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14347), .S(n14808), .Z(
        P1_U3528) );
  MUX2_X1 U16183 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14348), .S(n6528), .Z(
        P1_U3527) );
  MUX2_X1 U16184 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14350), .S(n6528), .Z(
        P1_U3525) );
  MUX2_X1 U16185 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14351), .S(n6528), .Z(
        P1_U3524) );
  MUX2_X1 U16186 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14353), .S(n6528), .Z(
        P1_U3522) );
  MUX2_X1 U16187 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14354), .S(n6528), .Z(
        P1_U3521) );
  MUX2_X1 U16188 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14355), .S(n6528), .Z(
        P1_U3520) );
  MUX2_X1 U16189 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14356), .S(n6528), .Z(
        P1_U3519) );
  MUX2_X1 U16190 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14357), .S(n6528), .Z(
        P1_U3518) );
  MUX2_X1 U16191 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14358), .S(n6528), .Z(
        P1_U3517) );
  MUX2_X1 U16192 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14359), .S(n6528), .Z(
        P1_U3516) );
  MUX2_X1 U16193 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14360), .S(n6528), .Z(
        P1_U3515) );
  MUX2_X1 U16194 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14361), .S(n6528), .Z(
        P1_U3513) );
  MUX2_X1 U16195 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14362), .S(n6528), .Z(
        P1_U3510) );
  OAI222_X1 U16196 ( .A1(n14370), .A2(n14365), .B1(P1_U3086), .B2(n14364), 
        .C1(n14363), .C2(n14372), .ZN(P1_U3326) );
  OAI222_X1 U16197 ( .A1(n14372), .A2(n14367), .B1(n14370), .B2(n14366), .C1(
        P1_U3086), .C2(n6526), .ZN(P1_U3328) );
  OAI222_X1 U16198 ( .A1(n14372), .A2(n14371), .B1(n14370), .B2(n14369), .C1(
        n14368), .C2(P1_U3086), .ZN(P1_U3329) );
  MUX2_X1 U16199 ( .A(n14374), .B(n14373), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16200 ( .A(n14375), .ZN(n14376) );
  MUX2_X1 U16201 ( .A(n14376), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16202 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14412) );
  NOR2_X1 U16203 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14377), .ZN(n14411) );
  INV_X1 U16204 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14733) );
  NOR2_X1 U16205 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14733), .ZN(n14410) );
  INV_X1 U16206 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15157) );
  XNOR2_X1 U16207 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .ZN(n14420) );
  INV_X1 U16208 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14407) );
  INV_X1 U16209 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14404) );
  XNOR2_X1 U16210 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14462) );
  INV_X1 U16211 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14402) );
  INV_X1 U16212 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14424) );
  INV_X1 U16213 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14397) );
  XNOR2_X1 U16214 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14455) );
  INV_X1 U16215 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14395) );
  NOR2_X1 U16216 ( .A1(n14384), .A2(n14385), .ZN(n14387) );
  AND2_X1 U16217 ( .A1(n14388), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14389) );
  NOR2_X1 U16218 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14390), .ZN(n14393) );
  XNOR2_X1 U16219 ( .A(n14390), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14449) );
  INV_X1 U16220 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14391) );
  XOR2_X1 U16221 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14426) );
  NAND2_X1 U16222 ( .A1(n14455), .A2(n14454), .ZN(n14396) );
  NOR2_X1 U16223 ( .A1(n14424), .A2(n14423), .ZN(n14400) );
  INV_X1 U16224 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U16225 ( .A1(n14424), .A2(n14423), .ZN(n14398) );
  XOR2_X1 U16226 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .Z(n14421) );
  NAND2_X1 U16227 ( .A1(n14462), .A2(n14461), .ZN(n14403) );
  INV_X1 U16228 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14405) );
  NAND2_X1 U16229 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14405), .ZN(n14406) );
  NAND2_X1 U16230 ( .A1(n14420), .A2(n14419), .ZN(n14408) );
  OAI22_X1 U16231 ( .A1(n14410), .A2(n14469), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14409), .ZN(n14417) );
  OAI22_X1 U16232 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14412), .B1(n14411), 
        .B2(n14417), .ZN(n14413) );
  NOR2_X1 U16233 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14413), .ZN(n14415) );
  INV_X1 U16234 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14533) );
  XNOR2_X1 U16235 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14413), .ZN(n14473) );
  NOR2_X1 U16236 ( .A1(n14533), .A2(n14473), .ZN(n14414) );
  NOR2_X1 U16237 ( .A1(n14415), .A2(n14414), .ZN(n14519) );
  XOR2_X1 U16238 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14416) );
  XNOR2_X1 U16239 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .ZN(n14418) );
  XNOR2_X1 U16240 ( .A(n14418), .B(n14417), .ZN(n14704) );
  XOR2_X1 U16241 ( .A(n14420), .B(n14419), .Z(n14698) );
  INV_X1 U16242 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14694) );
  XOR2_X1 U16243 ( .A(n14422), .B(n14421), .Z(n14688) );
  XOR2_X1 U16244 ( .A(n14424), .B(n14423), .Z(n14425) );
  XNOR2_X1 U16245 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14425), .ZN(n14460) );
  XOR2_X1 U16246 ( .A(n14427), .B(n14426), .Z(n14453) );
  NAND2_X1 U16247 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14429), .ZN(n14441) );
  INV_X1 U16248 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14839) );
  XNOR2_X1 U16249 ( .A(n14431), .B(n14430), .ZN(n14477) );
  XOR2_X1 U16250 ( .A(n14432), .B(n14433), .Z(n14435) );
  NAND2_X1 U16251 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14435), .ZN(n14437) );
  AOI21_X1 U16252 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14434), .A(n14433), .ZN(
        n15442) );
  NOR2_X1 U16253 ( .A1(n15442), .A2(n15441), .ZN(n15450) );
  NAND2_X1 U16254 ( .A1(n14477), .A2(n14478), .ZN(n14438) );
  NOR2_X1 U16255 ( .A1(n14477), .A2(n14478), .ZN(n14476) );
  XNOR2_X1 U16256 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14439), .ZN(n15446) );
  NAND2_X1 U16257 ( .A1(n15447), .A2(n15446), .ZN(n14440) );
  NOR2_X1 U16258 ( .A1(n15447), .A2(n15446), .ZN(n15445) );
  NAND2_X1 U16259 ( .A1(n14445), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14448) );
  XNOR2_X1 U16260 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14447) );
  XOR2_X1 U16261 ( .A(n14447), .B(n14446), .Z(n14480) );
  NAND2_X1 U16262 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14450), .ZN(n14451) );
  XNOR2_X1 U16263 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14449), .ZN(n15444) );
  XNOR2_X1 U16264 ( .A(n14455), .B(n14454), .ZN(n14457) );
  NAND2_X1 U16265 ( .A1(n14456), .A2(n14457), .ZN(n14458) );
  XNOR2_X1 U16266 ( .A(n14462), .B(n14461), .ZN(n14692) );
  XOR2_X1 U16267 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14464) );
  XOR2_X1 U16268 ( .A(n14465), .B(n14464), .Z(n14466) );
  XOR2_X1 U16269 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14468) );
  XOR2_X1 U16270 ( .A(n14469), .B(n14468), .Z(n14471) );
  AND2_X1 U16271 ( .A1(n14470), .A2(n14471), .ZN(n14702) );
  XNOR2_X1 U16272 ( .A(n14533), .B(n14473), .ZN(n14513) );
  XOR2_X1 U16273 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14474), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16274 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14475) );
  OAI21_X1 U16275 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14475), 
        .ZN(U28) );
  AOI21_X1 U16276 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14479) );
  XNOR2_X1 U16277 ( .A(n14479), .B(n14839), .ZN(SUB_1596_U61) );
  XOR2_X1 U16278 ( .A(n14481), .B(n14480), .Z(SUB_1596_U57) );
  XNOR2_X1 U16279 ( .A(n14482), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16280 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14483), .Z(SUB_1596_U54) );
  XNOR2_X1 U16281 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14484), .ZN(SUB_1596_U70)
         );
  XNOR2_X1 U16282 ( .A(n14486), .B(n14485), .ZN(n14503) );
  OAI211_X1 U16283 ( .C1(n14488), .C2(n14506), .A(n8808), .B(n14487), .ZN(
        n14504) );
  OAI22_X1 U16284 ( .A1(n14503), .A2(n14739), .B1(n14489), .B2(n14504), .ZN(
        n14490) );
  INV_X1 U16285 ( .A(n14490), .ZN(n14502) );
  XNOR2_X1 U16286 ( .A(n14492), .B(n14491), .ZN(n14495) );
  AOI21_X1 U16287 ( .B1(n14495), .B2(n14494), .A(n14493), .ZN(n14505) );
  OAI21_X1 U16288 ( .B1(n14496), .B2(n14503), .A(n14505), .ZN(n14500) );
  NOR2_X1 U16289 ( .A1(n14506), .A2(n14738), .ZN(n14499) );
  OAI22_X1 U16290 ( .A1(n14639), .A2(n9592), .B1(n14497), .B2(n14642), .ZN(
        n14498) );
  AOI211_X1 U16291 ( .C1(n14500), .C2(n14639), .A(n14499), .B(n14498), .ZN(
        n14501) );
  NAND2_X1 U16292 ( .A1(n14502), .A2(n14501), .ZN(P1_U3281) );
  INV_X1 U16293 ( .A(n14503), .ZN(n14508) );
  OAI211_X1 U16294 ( .C1(n14506), .C2(n14793), .A(n14505), .B(n14504), .ZN(
        n14507) );
  AOI21_X1 U16295 ( .B1(n14508), .B2(n14796), .A(n14507), .ZN(n14510) );
  INV_X1 U16296 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U16297 ( .A1(n6528), .A2(n14510), .B1(n14509), .B2(n14797), .ZN(
        P1_U3495) );
  AOI22_X1 U16298 ( .A1(n14808), .A2(n14510), .B1(n10351), .B2(n14806), .ZN(
        P1_U3540) );
  OAI21_X1 U16299 ( .B1(n14513), .B2(n14512), .A(n14511), .ZN(n14514) );
  XNOR2_X1 U16300 ( .A(n14514), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U16301 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14517) );
  OR2_X1 U16302 ( .A1(n14517), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U16303 ( .A1(n14519), .A2(n14518), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n14517), .ZN(n14521) );
  XNOR2_X1 U16304 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14520) );
  XNOR2_X1 U16305 ( .A(n14521), .B(n14520), .ZN(n14522) );
  AOI21_X1 U16306 ( .B1(n14526), .B2(n14525), .A(n14524), .ZN(n14541) );
  OAI21_X1 U16307 ( .B1(n14528), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14527), 
        .ZN(n14539) );
  NAND2_X1 U16308 ( .A1(n14543), .A2(n14529), .ZN(n14531) );
  OAI211_X1 U16309 ( .C1(n14533), .C2(n14532), .A(n14531), .B(n14530), .ZN(
        n14538) );
  AOI211_X1 U16310 ( .C1(n14536), .C2(n14535), .A(n14983), .B(n14534), .ZN(
        n14537) );
  AOI211_X1 U16311 ( .C1(n14990), .C2(n14539), .A(n14538), .B(n14537), .ZN(
        n14540) );
  OAI21_X1 U16312 ( .B1(n14541), .B2(n14994), .A(n14540), .ZN(P3_U3199) );
  AOI22_X1 U16313 ( .A1(n14543), .A2(n14542), .B1(n14987), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14561) );
  OAI21_X1 U16314 ( .B1(n14546), .B2(n14545), .A(n14544), .ZN(n14552) );
  AOI21_X1 U16315 ( .B1(n14549), .B2(n14548), .A(n14547), .ZN(n14550) );
  NOR2_X1 U16316 ( .A1(n14550), .A2(n14983), .ZN(n14551) );
  AOI21_X1 U16317 ( .B1(n14990), .B2(n14552), .A(n14551), .ZN(n14560) );
  INV_X1 U16318 ( .A(n14553), .ZN(n14559) );
  OAI221_X1 U16319 ( .B1(n14557), .B2(n14556), .C1(n14557), .C2(n14555), .A(
        n14554), .ZN(n14558) );
  NAND4_X1 U16320 ( .A1(n14561), .A2(n14560), .A3(n14559), .A4(n14558), .ZN(
        P3_U3200) );
  XNOR2_X1 U16321 ( .A(n14562), .B(n14566), .ZN(n14565) );
  AOI222_X1 U16322 ( .A1(n15068), .A2(n14565), .B1(n14564), .B2(n15065), .C1(
        n14563), .C2(n15062), .ZN(n14588) );
  AOI22_X1 U16323 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n15083), .B1(n15075), 
        .B2(n7692), .ZN(n14572) );
  XNOR2_X1 U16324 ( .A(n14567), .B(n14566), .ZN(n14591) );
  INV_X1 U16325 ( .A(n14568), .ZN(n14569) );
  NOR2_X1 U16326 ( .A1(n14569), .A2(n15054), .ZN(n14590) );
  AOI22_X1 U16327 ( .A1(n14591), .A2(n14570), .B1(n15028), .B2(n14590), .ZN(
        n14571) );
  OAI211_X1 U16328 ( .C1(n15083), .C2(n14588), .A(n14572), .B(n14571), .ZN(
        P3_U3220) );
  INV_X1 U16329 ( .A(n15034), .ZN(n14582) );
  OAI21_X1 U16330 ( .B1(n10909), .B2(n10908), .A(n14573), .ZN(n14600) );
  NAND2_X1 U16331 ( .A1(n14575), .A2(n14574), .ZN(n15004) );
  NAND2_X1 U16332 ( .A1(n15004), .A2(n14996), .ZN(n14577) );
  NAND2_X1 U16333 ( .A1(n14577), .A2(n14576), .ZN(n14579) );
  XNOR2_X1 U16334 ( .A(n14579), .B(n14578), .ZN(n14580) );
  OAI222_X1 U16335 ( .A1(n15046), .A2(n14581), .B1(n15048), .B2(n15019), .C1(
        n14580), .C2(n15053), .ZN(n14598) );
  AOI21_X1 U16336 ( .B1(n14582), .B2(n14600), .A(n14598), .ZN(n14587) );
  NOR2_X1 U16337 ( .A1(n14583), .A2(n15054), .ZN(n14599) );
  AOI22_X1 U16338 ( .A1(n14599), .A2(n15028), .B1(n15075), .B2(n14584), .ZN(
        n14585) );
  OAI221_X1 U16339 ( .B1(n15083), .B2(n14587), .C1(n15080), .C2(n14586), .A(
        n14585), .ZN(P3_U3222) );
  INV_X1 U16340 ( .A(n14588), .ZN(n14589) );
  AOI211_X1 U16341 ( .C1(n14591), .C2(n14601), .A(n14590), .B(n14589), .ZN(
        n14604) );
  INV_X1 U16342 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16343 ( .A1(n15142), .A2(n14604), .B1(n14592), .B2(n15140), .ZN(
        P3_U3472) );
  AND2_X1 U16344 ( .A1(n14593), .A2(n14601), .ZN(n14595) );
  NOR3_X1 U16345 ( .A1(n14596), .A2(n14595), .A3(n14594), .ZN(n14606) );
  AOI22_X1 U16346 ( .A1(n15142), .A2(n14606), .B1(n14597), .B2(n15140), .ZN(
        P3_U3471) );
  AOI211_X1 U16347 ( .C1(n14601), .C2(n14600), .A(n14599), .B(n14598), .ZN(
        n14608) );
  INV_X1 U16348 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U16349 ( .A1(n15142), .A2(n14608), .B1(n14602), .B2(n15140), .ZN(
        P3_U3470) );
  INV_X1 U16350 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14603) );
  AOI22_X1 U16351 ( .A1(n15127), .A2(n14604), .B1(n14603), .B2(n15125), .ZN(
        P3_U3429) );
  INV_X1 U16352 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14605) );
  AOI22_X1 U16353 ( .A1(n15127), .A2(n14606), .B1(n14605), .B2(n15125), .ZN(
        P3_U3426) );
  INV_X1 U16354 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U16355 ( .A1(n15127), .A2(n14608), .B1(n14607), .B2(n15125), .ZN(
        P3_U3423) );
  OAI21_X1 U16356 ( .B1(n14611), .B2(n14610), .A(n14609), .ZN(n14613) );
  AOI222_X1 U16357 ( .A1(n14616), .A2(n14672), .B1(n14615), .B2(n14614), .C1(
        n14613), .C2(n14612), .ZN(n14618) );
  OAI211_X1 U16358 ( .C1(n14620), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        P1_U3236) );
  XOR2_X1 U16359 ( .A(n14621), .B(n14627), .Z(n14647) );
  AOI211_X1 U16360 ( .C1(n14645), .C2(n14623), .A(n14674), .B(n14622), .ZN(
        n14644) );
  INV_X1 U16361 ( .A(n14645), .ZN(n14625) );
  OAI21_X1 U16362 ( .B1(n14625), .B2(n14624), .A(n14639), .ZN(n14634) );
  AOI21_X1 U16363 ( .B1(n14627), .B2(n14626), .A(n6679), .ZN(n14628) );
  OAI222_X1 U16364 ( .A1(n14633), .A2(n14632), .B1(n14631), .B2(n14630), .C1(
        n14629), .C2(n14628), .ZN(n14643) );
  AOI211_X1 U16365 ( .C1(n14644), .C2(n14635), .A(n14634), .B(n14643), .ZN(
        n14636) );
  OAI21_X1 U16366 ( .B1(n14647), .B2(n14637), .A(n14636), .ZN(n14638) );
  OAI21_X1 U16367 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14639), .A(n14638), 
        .ZN(n14640) );
  OAI21_X1 U16368 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(P1_U3277) );
  AOI211_X1 U16369 ( .C1(n14759), .C2(n14645), .A(n14644), .B(n14643), .ZN(
        n14646) );
  OAI21_X1 U16370 ( .B1(n14663), .B2(n14647), .A(n14646), .ZN(n14648) );
  INV_X1 U16371 ( .A(n14648), .ZN(n14682) );
  AOI22_X1 U16372 ( .A1(n14808), .A2(n14682), .B1(n14649), .B2(n14806), .ZN(
        P1_U3544) );
  OAI21_X1 U16373 ( .B1(n7497), .B2(n14793), .A(n14650), .ZN(n14651) );
  AOI21_X1 U16374 ( .B1(n14652), .B2(n14796), .A(n14651), .ZN(n14653) );
  AND2_X1 U16375 ( .A1(n14654), .A2(n14653), .ZN(n14683) );
  AOI22_X1 U16376 ( .A1(n14808), .A2(n14683), .B1(n15326), .B2(n14806), .ZN(
        P1_U3543) );
  AND3_X1 U16377 ( .A1(n6959), .A2(n14796), .A3(n14655), .ZN(n14661) );
  OAI211_X1 U16378 ( .C1(n14659), .C2(n14793), .A(n14658), .B(n14657), .ZN(
        n14660) );
  NOR3_X1 U16379 ( .A1(n14662), .A2(n14661), .A3(n14660), .ZN(n14684) );
  AOI22_X1 U16380 ( .A1(n14808), .A2(n14684), .B1(n10621), .B2(n14806), .ZN(
        P1_U3542) );
  NOR2_X1 U16381 ( .A1(n14664), .A2(n14663), .ZN(n14670) );
  AOI21_X1 U16382 ( .B1(n14666), .B2(n14759), .A(n14665), .ZN(n14667) );
  NAND2_X1 U16383 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  NOR3_X1 U16384 ( .A1(n14671), .A2(n14670), .A3(n14669), .ZN(n14685) );
  AOI22_X1 U16385 ( .A1(n14808), .A2(n14685), .B1(n10606), .B2(n14806), .ZN(
        P1_U3541) );
  INV_X1 U16386 ( .A(n14672), .ZN(n14673) );
  OAI22_X1 U16387 ( .A1(n14675), .A2(n14674), .B1(n14673), .B2(n14793), .ZN(
        n14676) );
  INV_X1 U16388 ( .A(n14676), .ZN(n14679) );
  NAND2_X1 U16389 ( .A1(n14677), .A2(n14796), .ZN(n14678) );
  AOI22_X1 U16390 ( .A1(n14808), .A2(n14687), .B1(n10227), .B2(n14806), .ZN(
        P1_U3539) );
  INV_X1 U16391 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16392 ( .A1(n6528), .A2(n14682), .B1(n14681), .B2(n14797), .ZN(
        P1_U3507) );
  INV_X1 U16393 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15211) );
  AOI22_X1 U16394 ( .A1(n6528), .A2(n14683), .B1(n15211), .B2(n14797), .ZN(
        P1_U3504) );
  AOI22_X1 U16395 ( .A1(n6528), .A2(n14684), .B1(n10620), .B2(n14797), .ZN(
        P1_U3501) );
  AOI22_X1 U16396 ( .A1(n6528), .A2(n14685), .B1(n10605), .B2(n14797), .ZN(
        P1_U3498) );
  INV_X1 U16397 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U16398 ( .A1(n6528), .A2(n14687), .B1(n14686), .B2(n14797), .ZN(
        P1_U3492) );
  AOI21_X1 U16399 ( .B1(n14689), .B2(n14688), .A(n6680), .ZN(n14690) );
  XNOR2_X1 U16400 ( .A(n14690), .B(n9845), .ZN(SUB_1596_U69) );
  AOI21_X1 U16401 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14695) );
  XNOR2_X1 U16402 ( .A(n14695), .B(n14694), .ZN(SUB_1596_U68) );
  XNOR2_X1 U16403 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14696), .ZN(SUB_1596_U67)
         );
  AOI21_X1 U16404 ( .B1(n14699), .B2(n14698), .A(n14697), .ZN(n14700) );
  XOR2_X1 U16405 ( .A(n14700), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16406 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  XOR2_X1 U16407 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14703), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16408 ( .B1(n14705), .B2(n14704), .A(n6654), .ZN(n14706) );
  XNOR2_X1 U16409 ( .A(n14706), .B(n11091), .ZN(SUB_1596_U64) );
  AND2_X1 U16410 ( .A1(n6526), .A2(n14707), .ZN(n14711) );
  NOR2_X1 U16411 ( .A1(n14709), .A2(n14711), .ZN(n14710) );
  MUX2_X1 U16412 ( .A(n14711), .B(n14710), .S(P1_IR_REG_0__SCAN_IN), .Z(n14714) );
  INV_X1 U16413 ( .A(n14712), .ZN(n14713) );
  OR2_X1 U16414 ( .A1(n14714), .A2(n14713), .ZN(n14717) );
  AOI22_X1 U16415 ( .A1(n14715), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14716) );
  OAI21_X1 U16416 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(P1_U3243) );
  AOI21_X1 U16417 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14720), .A(n14719), 
        .ZN(n14721) );
  INV_X1 U16418 ( .A(n14721), .ZN(n14729) );
  OAI21_X1 U16419 ( .B1(n14723), .B2(n15326), .A(n14722), .ZN(n14726) );
  AOI222_X1 U16420 ( .A1(n14729), .A2(n14728), .B1(n14727), .B2(n14726), .C1(
        n14725), .C2(n14724), .ZN(n14731) );
  OAI211_X1 U16421 ( .C1(n14733), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        P1_U3258) );
  AOI22_X1 U16422 ( .A1(n14747), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14735), 
        .B2(n14734), .ZN(n14736) );
  OAI21_X1 U16423 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14742) );
  NOR2_X1 U16424 ( .A1(n14740), .A2(n14739), .ZN(n14741) );
  AOI211_X1 U16425 ( .C1(n14744), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14745) );
  OAI21_X1 U16426 ( .B1(n14747), .B2(n14746), .A(n14745), .ZN(P1_U3290) );
  AND2_X1 U16427 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14749), .ZN(P1_U3294) );
  AND2_X1 U16428 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14749), .ZN(P1_U3295) );
  AND2_X1 U16429 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14749), .ZN(P1_U3296) );
  AND2_X1 U16430 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14749), .ZN(P1_U3297) );
  AND2_X1 U16431 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14749), .ZN(P1_U3298) );
  AND2_X1 U16432 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14749), .ZN(P1_U3299) );
  AND2_X1 U16433 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14749), .ZN(P1_U3300) );
  AND2_X1 U16434 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14749), .ZN(P1_U3301) );
  INV_X1 U16435 ( .A(n14749), .ZN(n14748) );
  NOR2_X1 U16436 ( .A1(n14748), .A2(n15182), .ZN(P1_U3302) );
  AND2_X1 U16437 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14749), .ZN(P1_U3303) );
  NOR2_X1 U16438 ( .A1(n14748), .A2(n15239), .ZN(P1_U3304) );
  AND2_X1 U16439 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14749), .ZN(P1_U3305) );
  AND2_X1 U16440 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14749), .ZN(P1_U3306) );
  NOR2_X1 U16441 ( .A1(n14748), .A2(n15199), .ZN(P1_U3307) );
  INV_X1 U16442 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15265) );
  NOR2_X1 U16443 ( .A1(n14748), .A2(n15265), .ZN(P1_U3308) );
  AND2_X1 U16444 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14749), .ZN(P1_U3309) );
  AND2_X1 U16445 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14749), .ZN(P1_U3310) );
  INV_X1 U16446 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15404) );
  NOR2_X1 U16447 ( .A1(n14748), .A2(n15404), .ZN(P1_U3311) );
  AND2_X1 U16448 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14749), .ZN(P1_U3312) );
  AND2_X1 U16449 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14749), .ZN(P1_U3313) );
  AND2_X1 U16450 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14749), .ZN(P1_U3314) );
  AND2_X1 U16451 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14749), .ZN(P1_U3315) );
  AND2_X1 U16452 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14749), .ZN(P1_U3316) );
  AND2_X1 U16453 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14749), .ZN(P1_U3317) );
  AND2_X1 U16454 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14749), .ZN(P1_U3318) );
  NOR2_X1 U16455 ( .A1(n14748), .A2(n15360), .ZN(P1_U3319) );
  AND2_X1 U16456 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14749), .ZN(P1_U3320) );
  AND2_X1 U16457 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14749), .ZN(P1_U3321) );
  AND2_X1 U16458 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14749), .ZN(P1_U3322) );
  AND2_X1 U16459 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14749), .ZN(P1_U3323) );
  INV_X1 U16460 ( .A(n14750), .ZN(n14756) );
  OAI21_X1 U16461 ( .B1(n14752), .B2(n14793), .A(n14751), .ZN(n14755) );
  INV_X1 U16462 ( .A(n14753), .ZN(n14754) );
  AOI211_X1 U16463 ( .C1(n14796), .C2(n14756), .A(n14755), .B(n14754), .ZN(
        n14798) );
  AOI22_X1 U16464 ( .A1(n6528), .A2(n14798), .B1(n8838), .B2(n14797), .ZN(
        P1_U3462) );
  AOI21_X1 U16465 ( .B1(n14759), .B2(n14758), .A(n14757), .ZN(n14760) );
  OAI211_X1 U16466 ( .C1(n14762), .C2(n14764), .A(n14761), .B(n14760), .ZN(
        n14763) );
  INV_X1 U16467 ( .A(n14763), .ZN(n14799) );
  AOI22_X1 U16468 ( .A1(n6528), .A2(n14799), .B1(n9519), .B2(n14797), .ZN(
        P1_U3474) );
  INV_X1 U16469 ( .A(n14764), .ZN(n14788) );
  INV_X1 U16470 ( .A(n14765), .ZN(n14770) );
  OAI21_X1 U16471 ( .B1(n14767), .B2(n14793), .A(n14766), .ZN(n14769) );
  AOI211_X1 U16472 ( .C1(n14788), .C2(n14770), .A(n14769), .B(n14768), .ZN(
        n14801) );
  AOI22_X1 U16473 ( .A1(n6528), .A2(n14801), .B1(n9751), .B2(n14797), .ZN(
        P1_U3477) );
  INV_X1 U16474 ( .A(n14771), .ZN(n14776) );
  OAI21_X1 U16475 ( .B1(n14773), .B2(n14793), .A(n14772), .ZN(n14775) );
  AOI211_X1 U16476 ( .C1(n14788), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14803) );
  AOI22_X1 U16477 ( .A1(n6528), .A2(n14803), .B1(n9773), .B2(n14797), .ZN(
        P1_U3480) );
  OAI211_X1 U16478 ( .C1(n7495), .C2(n14793), .A(n14778), .B(n14777), .ZN(
        n14779) );
  AOI21_X1 U16479 ( .B1(n14780), .B2(n14796), .A(n14779), .ZN(n14804) );
  INV_X1 U16480 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14781) );
  AOI22_X1 U16481 ( .A1(n6528), .A2(n14804), .B1(n14781), .B2(n14797), .ZN(
        P1_U3483) );
  INV_X1 U16482 ( .A(n14782), .ZN(n14787) );
  OAI21_X1 U16483 ( .B1(n14784), .B2(n14793), .A(n14783), .ZN(n14786) );
  AOI211_X1 U16484 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14805) );
  INV_X1 U16485 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14789) );
  AOI22_X1 U16486 ( .A1(n6528), .A2(n14805), .B1(n14789), .B2(n14797), .ZN(
        P1_U3486) );
  OAI211_X1 U16487 ( .C1(n6824), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14794) );
  AOI21_X1 U16488 ( .B1(n14796), .B2(n14795), .A(n14794), .ZN(n14807) );
  AOI22_X1 U16489 ( .A1(n6528), .A2(n14807), .B1(n10040), .B2(n14797), .ZN(
        P1_U3489) );
  AOI22_X1 U16490 ( .A1(n14808), .A2(n14798), .B1(n8678), .B2(n14806), .ZN(
        P1_U3529) );
  AOI22_X1 U16491 ( .A1(n14808), .A2(n14799), .B1(n9518), .B2(n14806), .ZN(
        P1_U3533) );
  INV_X1 U16492 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U16493 ( .A1(n14808), .A2(n14801), .B1(n14800), .B2(n14806), .ZN(
        P1_U3534) );
  INV_X1 U16494 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14802) );
  AOI22_X1 U16495 ( .A1(n14808), .A2(n14803), .B1(n14802), .B2(n14806), .ZN(
        P1_U3535) );
  AOI22_X1 U16496 ( .A1(n14808), .A2(n14804), .B1(n9936), .B2(n14806), .ZN(
        P1_U3536) );
  AOI22_X1 U16497 ( .A1(n14808), .A2(n14805), .B1(n10028), .B2(n14806), .ZN(
        P1_U3537) );
  AOI22_X1 U16498 ( .A1(n14808), .A2(n14807), .B1(n8768), .B2(n14806), .ZN(
        P1_U3538) );
  NOR2_X1 U16499 ( .A1(n14809), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16500 ( .A1(n14811), .A2(n14810), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8023), .ZN(n14817) );
  AOI211_X1 U16501 ( .C1(n14815), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14816) );
  AOI211_X1 U16502 ( .C1(n14819), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        n14820) );
  OAI21_X1 U16503 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(P2_U3206) );
  INV_X1 U16504 ( .A(n14823), .ZN(n14824) );
  OAI21_X1 U16505 ( .B1(n14826), .B2(n14825), .A(n14824), .ZN(n14831) );
  NOR2_X1 U16506 ( .A1(n14827), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14828) );
  AOI21_X1 U16507 ( .B1(n14865), .B2(n14829), .A(n14828), .ZN(n14830) );
  OAI21_X1 U16508 ( .B1(n14858), .B2(n14831), .A(n14830), .ZN(n14832) );
  INV_X1 U16509 ( .A(n14832), .ZN(n14838) );
  NAND2_X1 U16510 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  NAND3_X1 U16511 ( .A1(n14867), .A2(n14836), .A3(n14835), .ZN(n14837) );
  OAI211_X1 U16512 ( .C1(n14873), .C2(n14839), .A(n14838), .B(n14837), .ZN(
        P2_U3216) );
  INV_X1 U16513 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14857) );
  AOI211_X1 U16514 ( .C1(n14842), .C2(n14841), .A(n14858), .B(n14840), .ZN(
        n14849) );
  INV_X1 U16515 ( .A(n14843), .ZN(n14848) );
  NOR3_X1 U16516 ( .A1(n14846), .A2(n14845), .A3(n14844), .ZN(n14847) );
  NOR3_X1 U16517 ( .A1(n14849), .A2(n14848), .A3(n14847), .ZN(n14856) );
  AOI211_X1 U16518 ( .C1(n14853), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14854) );
  INV_X1 U16519 ( .A(n14854), .ZN(n14855) );
  OAI211_X1 U16520 ( .C1(n14873), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        P2_U3222) );
  INV_X1 U16521 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14872) );
  NOR2_X1 U16522 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8023), .ZN(n14863) );
  AOI211_X1 U16523 ( .C1(n14861), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14862) );
  AOI211_X1 U16524 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14871) );
  OAI211_X1 U16525 ( .C1(n14869), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14870) );
  OAI211_X1 U16526 ( .C1(n14873), .C2(n14872), .A(n14871), .B(n14870), .ZN(
        P2_U3227) );
  NAND2_X1 U16527 ( .A1(n14875), .A2(n14874), .ZN(n14878) );
  AOI22_X1 U16528 ( .A1(n13561), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14876), 
        .B2(n14902), .ZN(n14877) );
  OAI211_X1 U16529 ( .C1(n14880), .C2(n14879), .A(n14878), .B(n14877), .ZN(
        n14881) );
  AOI21_X1 U16530 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14884) );
  OAI21_X1 U16531 ( .B1(n13561), .B2(n14885), .A(n14884), .ZN(P2_U3258) );
  XNOR2_X1 U16532 ( .A(n14887), .B(n14886), .ZN(n14928) );
  AND2_X1 U16533 ( .A1(n14928), .A2(n14888), .ZN(n14906) );
  OAI21_X1 U16534 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14893) );
  NAND2_X1 U16535 ( .A1(n14893), .A2(n14892), .ZN(n14895) );
  NAND2_X1 U16536 ( .A1(n14895), .A2(n14894), .ZN(n14932) );
  AOI21_X1 U16537 ( .B1(n14897), .B2(n14901), .A(n14896), .ZN(n14899) );
  NAND2_X1 U16538 ( .A1(n14899), .A2(n14898), .ZN(n14929) );
  AOI22_X1 U16539 ( .A1(n14903), .A2(n14902), .B1(n14901), .B2(n14900), .ZN(
        n14904) );
  OAI21_X1 U16540 ( .B1(n14929), .B2(n6527), .A(n14904), .ZN(n14905) );
  NOR3_X1 U16541 ( .A1(n14906), .A2(n14932), .A3(n14905), .ZN(n14907) );
  AOI22_X1 U16542 ( .A1(n13561), .A2(n8907), .B1(n14907), .B2(n13598), .ZN(
        P2_U3262) );
  INV_X1 U16543 ( .A(n14909), .ZN(n14910) );
  AND2_X1 U16544 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14910), .ZN(P2_U3266) );
  AND2_X1 U16545 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14910), .ZN(P2_U3267) );
  AND2_X1 U16546 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14910), .ZN(P2_U3268) );
  AND2_X1 U16547 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14910), .ZN(P2_U3269) );
  AND2_X1 U16548 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14910), .ZN(P2_U3270) );
  AND2_X1 U16549 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14910), .ZN(P2_U3271) );
  AND2_X1 U16550 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14910), .ZN(P2_U3272) );
  AND2_X1 U16551 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14910), .ZN(P2_U3273) );
  INV_X1 U16552 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16553 ( .A1(n14909), .A2(n15343), .ZN(P2_U3274) );
  AND2_X1 U16554 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14910), .ZN(P2_U3275) );
  AND2_X1 U16555 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14910), .ZN(P2_U3276) );
  AND2_X1 U16556 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14910), .ZN(P2_U3277) );
  INV_X1 U16557 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15366) );
  NOR2_X1 U16558 ( .A1(n14909), .A2(n15366), .ZN(P2_U3278) );
  INV_X1 U16559 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15406) );
  NOR2_X1 U16560 ( .A1(n14909), .A2(n15406), .ZN(P2_U3279) );
  AND2_X1 U16561 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14910), .ZN(P2_U3280) );
  INV_X1 U16562 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15408) );
  NOR2_X1 U16563 ( .A1(n14909), .A2(n15408), .ZN(P2_U3281) );
  AND2_X1 U16564 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14910), .ZN(P2_U3282) );
  AND2_X1 U16565 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14910), .ZN(P2_U3283) );
  AND2_X1 U16566 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14910), .ZN(P2_U3284) );
  AND2_X1 U16567 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14910), .ZN(P2_U3285) );
  AND2_X1 U16568 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14910), .ZN(P2_U3286) );
  AND2_X1 U16569 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14910), .ZN(P2_U3287) );
  INV_X1 U16570 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15214) );
  NOR2_X1 U16571 ( .A1(n14909), .A2(n15214), .ZN(P2_U3288) );
  AND2_X1 U16572 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14910), .ZN(P2_U3289) );
  AND2_X1 U16573 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14910), .ZN(P2_U3290) );
  AND2_X1 U16574 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14910), .ZN(P2_U3291) );
  AND2_X1 U16575 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14910), .ZN(P2_U3292) );
  INV_X1 U16576 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15144) );
  NOR2_X1 U16577 ( .A1(n14909), .A2(n15144), .ZN(P2_U3293) );
  AND2_X1 U16578 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14910), .ZN(P2_U3294) );
  AND2_X1 U16579 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14910), .ZN(P2_U3295) );
  AOI22_X1 U16580 ( .A1(n14916), .A2(n14912), .B1(n14911), .B2(n14913), .ZN(
        P2_U3416) );
  AOI22_X1 U16581 ( .A1(n14916), .A2(n14915), .B1(n14914), .B2(n14913), .ZN(
        P2_U3417) );
  AOI211_X1 U16582 ( .C1(n14943), .C2(n14919), .A(n14918), .B(n14917), .ZN(
        n14963) );
  AOI22_X1 U16583 ( .A1(n14962), .A2(n14963), .B1(n7267), .B2(n14961), .ZN(
        P2_U3430) );
  INV_X1 U16584 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U16585 ( .A1(n14962), .A2(n14920), .B1(n15171), .B2(n14961), .ZN(
        P2_U3433) );
  INV_X1 U16586 ( .A(n14924), .ZN(n14926) );
  AOI21_X1 U16587 ( .B1(n14953), .B2(n7852), .A(n14921), .ZN(n14923) );
  OAI211_X1 U16588 ( .C1(n14924), .C2(n14955), .A(n14923), .B(n14922), .ZN(
        n14925) );
  AOI21_X1 U16589 ( .B1(n14960), .B2(n14926), .A(n14925), .ZN(n14965) );
  AOI22_X1 U16590 ( .A1(n14962), .A2(n14965), .B1(n7839), .B2(n14961), .ZN(
        P2_U3436) );
  AND2_X1 U16591 ( .A1(n14928), .A2(n14927), .ZN(n14933) );
  OAI21_X1 U16592 ( .B1(n14930), .B2(n14946), .A(n14929), .ZN(n14931) );
  NOR3_X1 U16593 ( .A1(n14933), .A2(n14932), .A3(n14931), .ZN(n14966) );
  INV_X1 U16594 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U16595 ( .A1(n14962), .A2(n14966), .B1(n14934), .B2(n14961), .ZN(
        P2_U3439) );
  INV_X1 U16596 ( .A(n14939), .ZN(n14941) );
  AOI21_X1 U16597 ( .B1(n14953), .B2(n14936), .A(n14935), .ZN(n14937) );
  OAI211_X1 U16598 ( .C1(n14955), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        n14940) );
  AOI21_X1 U16599 ( .B1(n14960), .B2(n14941), .A(n14940), .ZN(n14968) );
  INV_X1 U16600 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14942) );
  AOI22_X1 U16601 ( .A1(n14962), .A2(n14968), .B1(n14942), .B2(n14961), .ZN(
        P2_U3442) );
  NAND2_X1 U16602 ( .A1(n14950), .A2(n14943), .ZN(n14945) );
  OAI211_X1 U16603 ( .C1(n14947), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14948) );
  AOI211_X1 U16604 ( .C1(n14960), .C2(n14950), .A(n14949), .B(n14948), .ZN(
        n14969) );
  AOI22_X1 U16605 ( .A1(n14962), .A2(n14969), .B1(n7882), .B2(n14961), .ZN(
        P2_U3445) );
  AOI21_X1 U16606 ( .B1(n14953), .B2(n14952), .A(n14951), .ZN(n14954) );
  OAI21_X1 U16607 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14957) );
  AOI211_X1 U16608 ( .C1(n14960), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14971) );
  AOI22_X1 U16609 ( .A1(n14962), .A2(n14971), .B1(n7936), .B2(n14961), .ZN(
        P2_U3454) );
  AOI22_X1 U16610 ( .A1(n14972), .A2(n14963), .B1(n9040), .B2(n14970), .ZN(
        P2_U3499) );
  INV_X1 U16611 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U16612 ( .A1(n14972), .A2(n14965), .B1(n14964), .B2(n14970), .ZN(
        P2_U3501) );
  AOI22_X1 U16613 ( .A1(n14972), .A2(n14966), .B1(n7856), .B2(n14970), .ZN(
        P2_U3502) );
  INV_X1 U16614 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16615 ( .A1(n14972), .A2(n14968), .B1(n14967), .B2(n14970), .ZN(
        P2_U3503) );
  AOI22_X1 U16616 ( .A1(n14972), .A2(n14969), .B1(n7883), .B2(n14970), .ZN(
        P2_U3504) );
  AOI22_X1 U16617 ( .A1(n14972), .A2(n14971), .B1(n9629), .B2(n14970), .ZN(
        P2_U3507) );
  NOR2_X1 U16618 ( .A1(P3_U3897), .A2(n14987), .ZN(P3_U3150) );
  AOI21_X1 U16619 ( .B1(n15030), .B2(n14974), .A(n14973), .ZN(n14995) );
  INV_X1 U16620 ( .A(n14975), .ZN(n14980) );
  AOI21_X1 U16621 ( .B1(n14977), .B2(n14979), .A(n14976), .ZN(n14978) );
  AOI21_X1 U16622 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14984) );
  OAI22_X1 U16623 ( .A1(n14984), .A2(n14983), .B1(n14982), .B2(n14981), .ZN(
        n14985) );
  AOI211_X1 U16624 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14987), .A(n14986), .B(
        n14985), .ZN(n14993) );
  OAI21_X1 U16625 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14989), .A(n14988), .ZN(
        n14991) );
  NAND2_X1 U16626 ( .A1(n14991), .A2(n14990), .ZN(n14992) );
  OAI211_X1 U16627 ( .C1(n14995), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        P3_U3191) );
  NAND2_X1 U16628 ( .A1(n14997), .A2(n14996), .ZN(n14998) );
  NAND2_X1 U16629 ( .A1(n14999), .A2(n14998), .ZN(n15122) );
  INV_X1 U16630 ( .A(n15122), .ZN(n15008) );
  AOI22_X1 U16631 ( .A1(n15062), .A2(n15001), .B1(n15000), .B2(n15065), .ZN(
        n15002) );
  OAI21_X1 U16632 ( .B1(n15122), .B2(n15072), .A(n15002), .ZN(n15003) );
  INV_X1 U16633 ( .A(n15003), .ZN(n15007) );
  XNOR2_X1 U16634 ( .A(n15004), .B(n6707), .ZN(n15005) );
  NAND2_X1 U16635 ( .A1(n15005), .A2(n15068), .ZN(n15006) );
  NAND2_X1 U16636 ( .A1(n15007), .A2(n15006), .ZN(n15124) );
  AOI21_X1 U16637 ( .B1(n15025), .B2(n15008), .A(n15124), .ZN(n15014) );
  NAND2_X1 U16638 ( .A1(n15009), .A2(n15073), .ZN(n15120) );
  INV_X1 U16639 ( .A(n15120), .ZN(n15011) );
  AOI22_X1 U16640 ( .A1(n15028), .A2(n15011), .B1(n15075), .B2(n15010), .ZN(
        n15012) );
  OAI221_X1 U16641 ( .B1(n15083), .B2(n15014), .C1(n15080), .C2(n15013), .A(
        n15012), .ZN(P3_U3223) );
  XNOR2_X1 U16642 ( .A(n15016), .B(n15015), .ZN(n15024) );
  INV_X1 U16643 ( .A(n15024), .ZN(n15119) );
  XNOR2_X1 U16644 ( .A(n15018), .B(n15017), .ZN(n15022) );
  OAI22_X1 U16645 ( .A1(n15020), .A2(n15048), .B1(n15019), .B2(n15046), .ZN(
        n15021) );
  AOI21_X1 U16646 ( .B1(n15022), .B2(n15068), .A(n15021), .ZN(n15023) );
  OAI21_X1 U16647 ( .B1(n15072), .B2(n15024), .A(n15023), .ZN(n15116) );
  AOI21_X1 U16648 ( .B1(n15025), .B2(n15119), .A(n15116), .ZN(n15031) );
  NOR2_X1 U16649 ( .A1(n15026), .A2(n15054), .ZN(n15117) );
  AOI22_X1 U16650 ( .A1(n15028), .A2(n15117), .B1(n15075), .B2(n15027), .ZN(
        n15029) );
  OAI221_X1 U16651 ( .B1(n15083), .B2(n15031), .C1(n15080), .C2(n15030), .A(
        n15029), .ZN(P3_U3224) );
  OAI21_X1 U16652 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15035) );
  MUX2_X1 U16653 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15035), .S(n15080), .Z(
        n15036) );
  AOI21_X1 U16654 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15039) );
  OAI21_X1 U16655 ( .B1(n15041), .B2(n15040), .A(n15039), .ZN(P3_U3227) );
  INV_X1 U16656 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15060) );
  XNOR2_X1 U16657 ( .A(n15042), .B(n15044), .ZN(n15052) );
  OAI21_X1 U16658 ( .B1(n15045), .B2(n15044), .A(n15043), .ZN(n15091) );
  OAI22_X1 U16659 ( .A1(n9252), .A2(n15048), .B1(n15047), .B2(n15046), .ZN(
        n15049) );
  AOI21_X1 U16660 ( .B1(n15091), .B2(n15050), .A(n15049), .ZN(n15051) );
  OAI21_X1 U16661 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n15089) );
  INV_X1 U16662 ( .A(n15091), .ZN(n15057) );
  NOR2_X1 U16663 ( .A1(n9876), .A2(n15054), .ZN(n15090) );
  INV_X1 U16664 ( .A(n15090), .ZN(n15055) );
  OAI22_X1 U16665 ( .A1(n15057), .A2(n15078), .B1(n15056), .B2(n15055), .ZN(
        n15058) );
  AOI211_X1 U16666 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15075), .A(n15089), .B(
        n15058), .ZN(n15059) );
  AOI22_X1 U16667 ( .A1(n15083), .A2(n15060), .B1(n15059), .B2(n15080), .ZN(
        P3_U3231) );
  XNOR2_X1 U16668 ( .A(n15067), .B(n15061), .ZN(n15084) );
  AOI22_X1 U16669 ( .A1(n15065), .A2(n15064), .B1(n15063), .B2(n15062), .ZN(
        n15071) );
  XNOR2_X1 U16670 ( .A(n15066), .B(n15067), .ZN(n15069) );
  NAND2_X1 U16671 ( .A1(n15069), .A2(n15068), .ZN(n15070) );
  OAI211_X1 U16672 ( .C1(n15084), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15085) );
  AND2_X1 U16673 ( .A1(n15074), .A2(n15073), .ZN(n15086) );
  AOI22_X1 U16674 ( .A1(n15086), .A2(n15076), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15075), .ZN(n15077) );
  OAI21_X1 U16675 ( .B1(n15084), .B2(n15078), .A(n15077), .ZN(n15079) );
  NOR2_X1 U16676 ( .A1(n15085), .A2(n15079), .ZN(n15081) );
  AOI22_X1 U16677 ( .A1(n15083), .A2(n15082), .B1(n15081), .B2(n15080), .ZN(
        P3_U3232) );
  INV_X1 U16678 ( .A(n15084), .ZN(n15087) );
  AOI211_X1 U16679 ( .C1(n15118), .C2(n15087), .A(n15086), .B(n15085), .ZN(
        n15128) );
  INV_X1 U16680 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U16681 ( .A1(n15127), .A2(n15128), .B1(n15088), .B2(n15125), .ZN(
        P3_U3393) );
  AOI211_X1 U16682 ( .C1(n15118), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15130) );
  INV_X1 U16683 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15201) );
  AOI22_X1 U16684 ( .A1(n15127), .A2(n15130), .B1(n15201), .B2(n15125), .ZN(
        P3_U3396) );
  INV_X1 U16685 ( .A(n15092), .ZN(n15093) );
  AOI211_X1 U16686 ( .C1(n15095), .C2(n15118), .A(n15094), .B(n15093), .ZN(
        n15132) );
  INV_X1 U16687 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U16688 ( .A1(n15127), .A2(n15132), .B1(n15418), .B2(n15125), .ZN(
        P3_U3399) );
  INV_X1 U16689 ( .A(n15096), .ZN(n15099) );
  AOI211_X1 U16690 ( .C1(n15099), .C2(n15118), .A(n15098), .B(n15097), .ZN(
        n15133) );
  INV_X1 U16691 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U16692 ( .A1(n15127), .A2(n15133), .B1(n15100), .B2(n15125), .ZN(
        P3_U3402) );
  INV_X1 U16693 ( .A(n15101), .ZN(n15104) );
  AOI211_X1 U16694 ( .C1(n15104), .C2(n15118), .A(n15103), .B(n15102), .ZN(
        n15134) );
  INV_X1 U16695 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U16696 ( .A1(n15127), .A2(n15134), .B1(n15105), .B2(n15125), .ZN(
        P3_U3405) );
  INV_X1 U16697 ( .A(n15106), .ZN(n15109) );
  AOI211_X1 U16698 ( .C1(n15109), .C2(n15118), .A(n15108), .B(n15107), .ZN(
        n15135) );
  INV_X1 U16699 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U16700 ( .A1(n15127), .A2(n15135), .B1(n15110), .B2(n15125), .ZN(
        P3_U3411) );
  INV_X1 U16701 ( .A(n15118), .ZN(n15121) );
  OAI21_X1 U16702 ( .B1(n15112), .B2(n15121), .A(n15111), .ZN(n15113) );
  NOR2_X1 U16703 ( .A1(n15114), .A2(n15113), .ZN(n15137) );
  INV_X1 U16704 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16705 ( .A1(n15127), .A2(n15137), .B1(n15115), .B2(n15125), .ZN(
        P3_U3414) );
  AOI211_X1 U16706 ( .C1(n15119), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15139) );
  INV_X1 U16707 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16708 ( .A1(n15127), .A2(n15139), .B1(n15169), .B2(n15125), .ZN(
        P3_U3417) );
  OAI21_X1 U16709 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15123) );
  NOR2_X1 U16710 ( .A1(n15124), .A2(n15123), .ZN(n15141) );
  INV_X1 U16711 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15126) );
  AOI22_X1 U16712 ( .A1(n15127), .A2(n15141), .B1(n15126), .B2(n15125), .ZN(
        P3_U3420) );
  AOI22_X1 U16713 ( .A1(n15142), .A2(n15128), .B1(n9126), .B2(n15140), .ZN(
        P3_U3460) );
  AOI22_X1 U16714 ( .A1(n15142), .A2(n15130), .B1(n15129), .B2(n15140), .ZN(
        P3_U3461) );
  INV_X1 U16715 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U16716 ( .A1(n15142), .A2(n15132), .B1(n15131), .B2(n15140), .ZN(
        P3_U3462) );
  AOI22_X1 U16717 ( .A1(n15142), .A2(n15133), .B1(n9095), .B2(n15140), .ZN(
        P3_U3463) );
  INV_X1 U16718 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U16719 ( .A1(n15142), .A2(n15134), .B1(n15405), .B2(n15140), .ZN(
        P3_U3464) );
  INV_X1 U16720 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U16721 ( .A1(n15142), .A2(n15135), .B1(n15364), .B2(n15140), .ZN(
        P3_U3466) );
  AOI22_X1 U16722 ( .A1(n15142), .A2(n15137), .B1(n15136), .B2(n15140), .ZN(
        P3_U3467) );
  INV_X1 U16723 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16724 ( .A1(n15142), .A2(n15139), .B1(n15138), .B2(n15140), .ZN(
        P3_U3468) );
  AOI22_X1 U16725 ( .A1(n15142), .A2(n15141), .B1(n9965), .B2(n15140), .ZN(
        P3_U3469) );
  AOI22_X1 U16726 ( .A1(n15145), .A2(keyinput44), .B1(keyinput97), .B2(n15144), 
        .ZN(n15143) );
  OAI221_X1 U16727 ( .B1(n15145), .B2(keyinput44), .C1(n15144), .C2(keyinput97), .A(n15143), .ZN(n15155) );
  AOI22_X1 U16728 ( .A1(n13496), .A2(keyinput22), .B1(n15147), .B2(keyinput121), .ZN(n15146) );
  OAI221_X1 U16729 ( .B1(n13496), .B2(keyinput22), .C1(n15147), .C2(
        keyinput121), .A(n15146), .ZN(n15154) );
  AOI22_X1 U16730 ( .A1(n15149), .A2(keyinput7), .B1(n15398), .B2(keyinput21), 
        .ZN(n15148) );
  OAI221_X1 U16731 ( .B1(n15149), .B2(keyinput7), .C1(n15398), .C2(keyinput21), 
        .A(n15148), .ZN(n15153) );
  XNOR2_X1 U16732 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput58), .ZN(n15151)
         );
  XNOR2_X1 U16733 ( .A(SI_2_), .B(keyinput43), .ZN(n15150) );
  NAND2_X1 U16734 ( .A1(n15151), .A2(n15150), .ZN(n15152) );
  NOR4_X1 U16735 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15197) );
  AOI22_X1 U16736 ( .A1(n7839), .A2(keyinput108), .B1(keyinput72), .B2(n15157), 
        .ZN(n15156) );
  OAI221_X1 U16737 ( .B1(n7839), .B2(keyinput108), .C1(n15157), .C2(keyinput72), .A(n15156), .ZN(n15167) );
  AOI22_X1 U16738 ( .A1(n15397), .A2(keyinput14), .B1(n15159), .B2(keyinput88), 
        .ZN(n15158) );
  OAI221_X1 U16739 ( .B1(n15397), .B2(keyinput14), .C1(n15159), .C2(keyinput88), .A(n15158), .ZN(n15166) );
  AOI22_X1 U16740 ( .A1(n10641), .A2(keyinput31), .B1(n15161), .B2(keyinput33), 
        .ZN(n15160) );
  OAI221_X1 U16741 ( .B1(n10641), .B2(keyinput31), .C1(n15161), .C2(keyinput33), .A(n15160), .ZN(n15165) );
  XNOR2_X1 U16742 ( .A(SI_8_), .B(keyinput66), .ZN(n15163) );
  XNOR2_X1 U16743 ( .A(SI_18_), .B(keyinput102), .ZN(n15162) );
  NAND2_X1 U16744 ( .A1(n15163), .A2(n15162), .ZN(n15164) );
  NOR4_X1 U16745 ( .A1(n15167), .A2(n15166), .A3(n15165), .A4(n15164), .ZN(
        n15196) );
  AOI22_X1 U16746 ( .A1(n15169), .A2(keyinput84), .B1(n15392), .B2(keyinput67), 
        .ZN(n15168) );
  OAI221_X1 U16747 ( .B1(n15169), .B2(keyinput84), .C1(n15392), .C2(keyinput67), .A(n15168), .ZN(n15179) );
  AOI22_X1 U16748 ( .A1(n15171), .A2(keyinput5), .B1(n8694), .B2(keyinput25), 
        .ZN(n15170) );
  OAI221_X1 U16749 ( .B1(n15171), .B2(keyinput5), .C1(n8694), .C2(keyinput25), 
        .A(n15170), .ZN(n15178) );
  INV_X1 U16750 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15173) );
  INV_X1 U16751 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U16752 ( .A1(n15173), .A2(keyinput27), .B1(keyinput85), .B2(n15393), 
        .ZN(n15172) );
  OAI221_X1 U16753 ( .B1(n15173), .B2(keyinput27), .C1(n15393), .C2(keyinput85), .A(n15172), .ZN(n15177) );
  XOR2_X1 U16754 ( .A(n8495), .B(keyinput83), .Z(n15175) );
  XNOR2_X1 U16755 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput32), .ZN(n15174) );
  NAND2_X1 U16756 ( .A1(n15175), .A2(n15174), .ZN(n15176) );
  NOR4_X1 U16757 ( .A1(n15179), .A2(n15178), .A3(n15177), .A4(n15176), .ZN(
        n15195) );
  AOI22_X1 U16758 ( .A1(n15182), .A2(keyinput91), .B1(n15181), .B2(keyinput45), 
        .ZN(n15180) );
  OAI221_X1 U16759 ( .B1(n15182), .B2(keyinput91), .C1(n15181), .C2(keyinput45), .A(n15180), .ZN(n15193) );
  AOI22_X1 U16760 ( .A1(n15185), .A2(keyinput82), .B1(n15184), .B2(keyinput78), 
        .ZN(n15183) );
  OAI221_X1 U16761 ( .B1(n15185), .B2(keyinput82), .C1(n15184), .C2(keyinput78), .A(n15183), .ZN(n15192) );
  XNOR2_X1 U16762 ( .A(n15186), .B(keyinput56), .ZN(n15191) );
  XOR2_X1 U16763 ( .A(n11798), .B(keyinput124), .Z(n15189) );
  XNOR2_X1 U16764 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput109), .ZN(n15188) );
  XNOR2_X1 U16765 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput104), .ZN(n15187)
         );
  NAND3_X1 U16766 ( .A1(n15189), .A2(n15188), .A3(n15187), .ZN(n15190) );
  NOR4_X1 U16767 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15194) );
  NAND4_X1 U16768 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15355) );
  AOI22_X1 U16769 ( .A1(n12858), .A2(keyinput34), .B1(keyinput115), .B2(n15199), .ZN(n15198) );
  OAI221_X1 U16770 ( .B1(n12858), .B2(keyinput34), .C1(n15199), .C2(
        keyinput115), .A(n15198), .ZN(n15209) );
  INV_X1 U16771 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U16772 ( .A1(n15395), .A2(keyinput80), .B1(n15201), .B2(keyinput57), 
        .ZN(n15200) );
  OAI221_X1 U16773 ( .B1(n15395), .B2(keyinput80), .C1(n15201), .C2(keyinput57), .A(n15200), .ZN(n15208) );
  AOI22_X1 U16774 ( .A1(n15377), .A2(keyinput119), .B1(keyinput29), .B2(n13468), .ZN(n15202) );
  OAI221_X1 U16775 ( .B1(n15377), .B2(keyinput119), .C1(n13468), .C2(
        keyinput29), .A(n15202), .ZN(n15207) );
  INV_X1 U16776 ( .A(keyinput9), .ZN(n15204) );
  AOI22_X1 U16777 ( .A1(n15205), .A2(keyinput54), .B1(P2_WR_REG_SCAN_IN), .B2(
        n15204), .ZN(n15203) );
  OAI221_X1 U16778 ( .B1(n15205), .B2(keyinput54), .C1(n15204), .C2(
        P2_WR_REG_SCAN_IN), .A(n15203), .ZN(n15206) );
  NOR4_X1 U16779 ( .A1(n15209), .A2(n15208), .A3(n15207), .A4(n15206), .ZN(
        n15249) );
  AOI22_X1 U16780 ( .A1(n15211), .A2(keyinput99), .B1(n15376), .B2(keyinput126), .ZN(n15210) );
  OAI221_X1 U16781 ( .B1(n15211), .B2(keyinput99), .C1(n15376), .C2(
        keyinput126), .A(n15210), .ZN(n15220) );
  AOI22_X1 U16782 ( .A1(n15375), .A2(keyinput106), .B1(n10620), .B2(keyinput20), .ZN(n15212) );
  OAI221_X1 U16783 ( .B1(n15375), .B2(keyinput106), .C1(n10620), .C2(
        keyinput20), .A(n15212), .ZN(n15219) );
  AOI22_X1 U16784 ( .A1(n15215), .A2(keyinput90), .B1(keyinput17), .B2(n15214), 
        .ZN(n15213) );
  OAI221_X1 U16785 ( .B1(n15215), .B2(keyinput90), .C1(n15214), .C2(keyinput17), .A(n15213), .ZN(n15218) );
  AOI22_X1 U16786 ( .A1(n15380), .A2(keyinput1), .B1(keyinput125), .B2(n15379), 
        .ZN(n15216) );
  OAI221_X1 U16787 ( .B1(n15380), .B2(keyinput1), .C1(n15379), .C2(keyinput125), .A(n15216), .ZN(n15217) );
  NOR4_X1 U16788 ( .A1(n15220), .A2(n15219), .A3(n15218), .A4(n15217), .ZN(
        n15248) );
  AOI22_X1 U16789 ( .A1(n15223), .A2(keyinput37), .B1(keyinput6), .B2(n15222), 
        .ZN(n15221) );
  OAI221_X1 U16790 ( .B1(n15223), .B2(keyinput37), .C1(n15222), .C2(keyinput6), 
        .A(n15221), .ZN(n15231) );
  AOI22_X1 U16791 ( .A1(n7882), .A2(keyinput62), .B1(keyinput52), .B2(n15378), 
        .ZN(n15224) );
  OAI221_X1 U16792 ( .B1(n7882), .B2(keyinput62), .C1(n15378), .C2(keyinput52), 
        .A(n15224), .ZN(n15230) );
  AOI22_X1 U16793 ( .A1(n11629), .A2(keyinput12), .B1(n15226), .B2(keyinput65), 
        .ZN(n15225) );
  OAI221_X1 U16794 ( .B1(n11629), .B2(keyinput12), .C1(n15226), .C2(keyinput65), .A(n15225), .ZN(n15229) );
  AOI22_X1 U16795 ( .A1(n8838), .A2(keyinput123), .B1(n8869), .B2(keyinput36), 
        .ZN(n15227) );
  OAI221_X1 U16796 ( .B1(n8838), .B2(keyinput123), .C1(n8869), .C2(keyinput36), 
        .A(n15227), .ZN(n15228) );
  NOR4_X1 U16797 ( .A1(n15231), .A2(n15230), .A3(n15229), .A4(n15228), .ZN(
        n15247) );
  INV_X1 U16798 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U16799 ( .A1(n15234), .A2(keyinput63), .B1(n15233), .B2(keyinput53), 
        .ZN(n15232) );
  OAI221_X1 U16800 ( .B1(n15234), .B2(keyinput63), .C1(n15233), .C2(keyinput53), .A(n15232), .ZN(n15237) );
  XNOR2_X1 U16801 ( .A(n15362), .B(keyinput112), .ZN(n15236) );
  XOR2_X1 U16802 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput117), .Z(n15235) );
  OR3_X1 U16803 ( .A1(n15237), .A2(n15236), .A3(n15235), .ZN(n15245) );
  INV_X1 U16804 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U16805 ( .A1(n15240), .A2(keyinput93), .B1(keyinput49), .B2(n15239), 
        .ZN(n15238) );
  OAI221_X1 U16806 ( .B1(n15240), .B2(keyinput93), .C1(n15239), .C2(keyinput49), .A(n15238), .ZN(n15244) );
  AOI22_X1 U16807 ( .A1(n15242), .A2(keyinput92), .B1(n15381), .B2(keyinput122), .ZN(n15241) );
  OAI221_X1 U16808 ( .B1(n15242), .B2(keyinput92), .C1(n15381), .C2(
        keyinput122), .A(n15241), .ZN(n15243) );
  NOR3_X1 U16809 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(n15246) );
  NAND4_X1 U16810 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        n15354) );
  AOI22_X1 U16811 ( .A1(n15252), .A2(keyinput127), .B1(keyinput19), .B2(n15251), .ZN(n15250) );
  OAI221_X1 U16812 ( .B1(n15252), .B2(keyinput127), .C1(n15251), .C2(
        keyinput19), .A(n15250), .ZN(n15256) );
  XNOR2_X1 U16813 ( .A(n15253), .B(keyinput111), .ZN(n15255) );
  XNOR2_X1 U16814 ( .A(n15368), .B(keyinput68), .ZN(n15254) );
  OR3_X1 U16815 ( .A1(n15256), .A2(n15255), .A3(n15254), .ZN(n15263) );
  AOI22_X1 U16816 ( .A1(n15360), .A2(keyinput60), .B1(n15361), .B2(keyinput40), 
        .ZN(n15257) );
  OAI221_X1 U16817 ( .B1(n15360), .B2(keyinput60), .C1(n15361), .C2(keyinput40), .A(n15257), .ZN(n15262) );
  AOI22_X1 U16818 ( .A1(n15260), .A2(keyinput113), .B1(n15259), .B2(keyinput74), .ZN(n15258) );
  OAI221_X1 U16819 ( .B1(n15260), .B2(keyinput113), .C1(n15259), .C2(
        keyinput74), .A(n15258), .ZN(n15261) );
  NOR3_X1 U16820 ( .A1(n15263), .A2(n15262), .A3(n15261), .ZN(n15303) );
  INV_X1 U16821 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U16822 ( .A1(n15365), .A2(keyinput26), .B1(n15265), .B2(keyinput15), 
        .ZN(n15264) );
  OAI221_X1 U16823 ( .B1(n15365), .B2(keyinput26), .C1(n15265), .C2(keyinput15), .A(n15264), .ZN(n15276) );
  INV_X1 U16824 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U16825 ( .A1(n15268), .A2(keyinput2), .B1(keyinput110), .B2(n15267), 
        .ZN(n15266) );
  OAI221_X1 U16826 ( .B1(n15268), .B2(keyinput2), .C1(n15267), .C2(keyinput110), .A(n15266), .ZN(n15275) );
  AOI22_X1 U16827 ( .A1(n15366), .A2(keyinput87), .B1(keyinput10), .B2(n15270), 
        .ZN(n15269) );
  OAI221_X1 U16828 ( .B1(n15366), .B2(keyinput87), .C1(n15270), .C2(keyinput10), .A(n15269), .ZN(n15274) );
  XOR2_X1 U16829 ( .A(n7013), .B(keyinput3), .Z(n15272) );
  XNOR2_X1 U16830 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput46), .ZN(n15271) );
  NAND2_X1 U16831 ( .A1(n15272), .A2(n15271), .ZN(n15273) );
  NOR4_X1 U16832 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15302) );
  INV_X1 U16833 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U16834 ( .A1(n8974), .A2(keyinput48), .B1(n15278), .B2(keyinput13), 
        .ZN(n15277) );
  OAI221_X1 U16835 ( .B1(n8974), .B2(keyinput48), .C1(n15278), .C2(keyinput13), 
        .A(n15277), .ZN(n15287) );
  AOI22_X1 U16836 ( .A1(n15364), .A2(keyinput79), .B1(n9675), .B2(keyinput77), 
        .ZN(n15279) );
  OAI221_X1 U16837 ( .B1(n15364), .B2(keyinput79), .C1(n9675), .C2(keyinput77), 
        .A(n15279), .ZN(n15286) );
  AOI22_X1 U16838 ( .A1(n13112), .A2(keyinput55), .B1(keyinput51), .B2(n15281), 
        .ZN(n15280) );
  OAI221_X1 U16839 ( .B1(n13112), .B2(keyinput55), .C1(n15281), .C2(keyinput51), .A(n15280), .ZN(n15285) );
  XOR2_X1 U16840 ( .A(n15363), .B(keyinput41), .Z(n15283) );
  XNOR2_X1 U16841 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput116), .ZN(n15282) );
  NAND2_X1 U16842 ( .A1(n15283), .A2(n15282), .ZN(n15284) );
  NOR4_X1 U16843 ( .A1(n15287), .A2(n15286), .A3(n15285), .A4(n15284), .ZN(
        n15301) );
  AOI22_X1 U16844 ( .A1(n7707), .A2(keyinput64), .B1(keyinput24), .B2(n13575), 
        .ZN(n15288) );
  OAI221_X1 U16845 ( .B1(n7707), .B2(keyinput64), .C1(n13575), .C2(keyinput24), 
        .A(n15288), .ZN(n15299) );
  AOI22_X1 U16846 ( .A1(n15290), .A2(keyinput39), .B1(keyinput76), .B2(n9126), 
        .ZN(n15289) );
  OAI221_X1 U16847 ( .B1(n15290), .B2(keyinput39), .C1(n9126), .C2(keyinput76), 
        .A(n15289), .ZN(n15298) );
  INV_X1 U16848 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U16849 ( .A1(n15293), .A2(keyinput30), .B1(keyinput69), .B2(n15292), 
        .ZN(n15291) );
  OAI221_X1 U16850 ( .B1(n15293), .B2(keyinput30), .C1(n15292), .C2(keyinput69), .A(n15291), .ZN(n15297) );
  XNOR2_X1 U16851 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput81), .ZN(n15295)
         );
  XNOR2_X1 U16852 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput105), .ZN(n15294) );
  NAND2_X1 U16853 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  NOR4_X1 U16854 ( .A1(n15299), .A2(n15298), .A3(n15297), .A4(n15296), .ZN(
        n15300) );
  NAND4_X1 U16855 ( .A1(n15303), .A2(n15302), .A3(n15301), .A4(n15300), .ZN(
        n15353) );
  AOI22_X1 U16856 ( .A1(n13545), .A2(keyinput75), .B1(n15305), .B2(keyinput11), 
        .ZN(n15304) );
  OAI221_X1 U16857 ( .B1(n13545), .B2(keyinput75), .C1(n15305), .C2(keyinput11), .A(n15304), .ZN(n15314) );
  AOI22_X1 U16858 ( .A1(n15307), .A2(keyinput38), .B1(keyinput100), .B2(n15413), .ZN(n15306) );
  OAI221_X1 U16859 ( .B1(n15307), .B2(keyinput38), .C1(n15413), .C2(
        keyinput100), .A(n15306), .ZN(n15313) );
  XOR2_X1 U16860 ( .A(n15418), .B(keyinput8), .Z(n15311) );
  XNOR2_X1 U16861 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput114), .ZN(n15310) );
  XNOR2_X1 U16862 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput42), .ZN(n15309) );
  XNOR2_X1 U16863 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput16), .ZN(n15308)
         );
  NAND4_X1 U16864 ( .A1(n15311), .A2(n15310), .A3(n15309), .A4(n15308), .ZN(
        n15312) );
  NOR3_X1 U16865 ( .A1(n15314), .A2(n15313), .A3(n15312), .ZN(n15351) );
  AOI22_X1 U16866 ( .A1(n15316), .A2(keyinput0), .B1(n13410), .B2(keyinput47), 
        .ZN(n15315) );
  OAI221_X1 U16867 ( .B1(n15316), .B2(keyinput0), .C1(n13410), .C2(keyinput47), 
        .A(n15315), .ZN(n15324) );
  INV_X1 U16868 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U16869 ( .A1(n15417), .A2(keyinput86), .B1(n15419), .B2(keyinput95), 
        .ZN(n15317) );
  OAI221_X1 U16870 ( .B1(n15417), .B2(keyinput86), .C1(n15419), .C2(keyinput95), .A(n15317), .ZN(n15323) );
  AOI22_X1 U16871 ( .A1(n9010), .A2(keyinput28), .B1(n15420), .B2(keyinput71), 
        .ZN(n15318) );
  OAI221_X1 U16872 ( .B1(n9010), .B2(keyinput28), .C1(n15420), .C2(keyinput71), 
        .A(n15318), .ZN(n15322) );
  XNOR2_X1 U16873 ( .A(SI_3_), .B(keyinput59), .ZN(n15320) );
  XNOR2_X1 U16874 ( .A(SI_19_), .B(keyinput89), .ZN(n15319) );
  NAND2_X1 U16875 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  NOR4_X1 U16876 ( .A1(n15324), .A2(n15323), .A3(n15322), .A4(n15321), .ZN(
        n15350) );
  AOI22_X1 U16877 ( .A1(n15405), .A2(keyinput94), .B1(keyinput18), .B2(n15326), 
        .ZN(n15325) );
  OAI221_X1 U16878 ( .B1(n15405), .B2(keyinput94), .C1(n15326), .C2(keyinput18), .A(n15325), .ZN(n15336) );
  AOI22_X1 U16879 ( .A1(n13585), .A2(keyinput4), .B1(n11073), .B2(keyinput120), 
        .ZN(n15327) );
  OAI221_X1 U16880 ( .B1(n13585), .B2(keyinput4), .C1(n11073), .C2(keyinput120), .A(n15327), .ZN(n15335) );
  AOI22_X1 U16881 ( .A1(n15329), .A2(keyinput101), .B1(n15404), .B2(keyinput70), .ZN(n15328) );
  OAI221_X1 U16882 ( .B1(n15329), .B2(keyinput101), .C1(n15404), .C2(
        keyinput70), .A(n15328), .ZN(n15334) );
  AOI22_X1 U16883 ( .A1(n15332), .A2(keyinput50), .B1(n15331), .B2(keyinput73), 
        .ZN(n15330) );
  OAI221_X1 U16884 ( .B1(n15332), .B2(keyinput50), .C1(n15331), .C2(keyinput73), .A(n15330), .ZN(n15333) );
  NOR4_X1 U16885 ( .A1(n15336), .A2(n15335), .A3(n15334), .A4(n15333), .ZN(
        n15349) );
  INV_X1 U16886 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U16887 ( .A1(n8281), .A2(keyinput96), .B1(n15407), .B2(keyinput107), 
        .ZN(n15337) );
  OAI221_X1 U16888 ( .B1(n8281), .B2(keyinput96), .C1(n15407), .C2(keyinput107), .A(n15337), .ZN(n15341) );
  XNOR2_X1 U16889 ( .A(n15408), .B(keyinput23), .ZN(n15340) );
  XNOR2_X1 U16890 ( .A(n15338), .B(keyinput98), .ZN(n15339) );
  OR3_X1 U16891 ( .A1(n15341), .A2(n15340), .A3(n15339), .ZN(n15347) );
  AOI22_X1 U16892 ( .A1(n15343), .A2(keyinput35), .B1(keyinput61), .B2(n15406), 
        .ZN(n15342) );
  OAI221_X1 U16893 ( .B1(n15343), .B2(keyinput35), .C1(n15406), .C2(keyinput61), .A(n15342), .ZN(n15346) );
  AOI22_X1 U16894 ( .A1(n7197), .A2(keyinput103), .B1(n12911), .B2(keyinput118), .ZN(n15344) );
  OAI221_X1 U16895 ( .B1(n7197), .B2(keyinput103), .C1(n12911), .C2(
        keyinput118), .A(n15344), .ZN(n15345) );
  NOR3_X1 U16896 ( .A1(n15347), .A2(n15346), .A3(n15345), .ZN(n15348) );
  NAND4_X1 U16897 ( .A1(n15351), .A2(n15350), .A3(n15349), .A4(n15348), .ZN(
        n15352) );
  NOR4_X1 U16898 ( .A1(n15355), .A2(n15354), .A3(n15353), .A4(n15352), .ZN(
        n15359) );
  INV_X1 U16899 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15357) );
  INV_X1 U16900 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15356) );
  AOI221_X1 U16901 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n15357), .C2(n15356), .A(P3_RD_REG_SCAN_IN), .ZN(n15358) );
  XNOR2_X1 U16902 ( .A(n15359), .B(n15358), .ZN(n15437) );
  NOR4_X1 U16903 ( .A1(P3_REG2_REG_3__SCAN_IN), .A2(P2_DATAO_REG_7__SCAN_IN), 
        .A3(n15361), .A4(n15360), .ZN(n15435) );
  NOR4_X1 U16904 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), .A3(P1_IR_REG_7__SCAN_IN), .A4(n15362), .ZN(n15434) );
  NAND4_X1 U16905 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(P3_REG1_REG_30__SCAN_IN), 
        .A3(P2_REG1_REG_7__SCAN_IN), .A4(n9675), .ZN(n15374) );
  NAND4_X1 U16906 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(n15364), .A4(n15363), .ZN(n15373) );
  NOR4_X1 U16907 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P2_REG0_REG_29__SCAN_IN), 
        .A3(n15366), .A4(n15365), .ZN(n15371) );
  NOR4_X1 U16908 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_REG1_REG_1__SCAN_IN), 
        .A3(P3_REG3_REG_0__SCAN_IN), .A4(P2_IR_REG_13__SCAN_IN), .ZN(n15370)
         );
  NOR4_X1 U16909 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P2_DATAO_REG_19__SCAN_IN), .A3(P2_IR_REG_2__SCAN_IN), .A4(n13575), .ZN(n15367) );
  AND4_X1 U16910 ( .A1(n7013), .A2(n15368), .A3(P1_IR_REG_10__SCAN_IN), .A4(
        n15367), .ZN(n15369) );
  NAND4_X1 U16911 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(
        P3_D_REG_2__SCAN_IN), .ZN(n15372) );
  NOR3_X1 U16912 ( .A1(n15374), .A2(n15373), .A3(n15372), .ZN(n15433) );
  NAND4_X1 U16913 ( .A1(P2_D_REG_9__SCAN_IN), .A2(SI_9_), .A3(
        P1_REG0_REG_14__SCAN_IN), .A4(n15375), .ZN(n15431) );
  NAND4_X1 U16914 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P2_WR_REG_SCAN_IN), .A4(n15376), .ZN(n15430) );
  NOR4_X1 U16915 ( .A1(P3_REG0_REG_2__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(P1_D_REG_18__SCAN_IN), .A4(n15377), .ZN(n15388) );
  NAND4_X1 U16916 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P1_REG2_REG_30__SCAN_IN), 
        .A3(n7882), .A4(n15378), .ZN(n15385) );
  NAND4_X1 U16917 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(P1_REG1_REG_19__SCAN_IN), 
        .A3(n15380), .A4(n15379), .ZN(n15384) );
  NAND4_X1 U16918 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .A3(P3_DATAO_REG_27__SCAN_IN), .A4(n15381), .ZN(n15383) );
  NAND4_X1 U16919 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .A3(P1_D_REG_21__SCAN_IN), .A4(P1_REG0_REG_1__SCAN_IN), .ZN(n15382) );
  NOR4_X1 U16920 ( .A1(n15385), .A2(n15384), .A3(n15383), .A4(n15382), .ZN(
        n15386) );
  NAND3_X1 U16921 ( .A1(n15388), .A2(n15387), .A3(n15386), .ZN(n15429) );
  NAND4_X1 U16922 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P2_REG1_REG_1__SCAN_IN), 
        .A3(P1_D_REG_0__SCAN_IN), .A4(P1_REG1_REG_27__SCAN_IN), .ZN(n15394) );
  NAND4_X1 U16923 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n15390)
         );
  NAND4_X1 U16924 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_REG0_REG_9__SCAN_IN), 
        .A3(SI_15_), .A4(P2_REG0_REG_1__SCAN_IN), .ZN(n15389) );
  OR4_X1 U16925 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(n15390), .A3(n15389), .A4(
        P3_REG2_REG_8__SCAN_IN), .ZN(n15391) );
  NOR4_X1 U16926 ( .A1(n15394), .A2(n15393), .A3(n15392), .A4(n15391), .ZN(
        n15427) );
  NAND4_X1 U16927 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P1_REG0_REG_29__SCAN_IN), 
        .A3(P2_ADDR_REG_5__SCAN_IN), .A4(n15395), .ZN(n15403) );
  NAND4_X1 U16928 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P1_REG2_REG_16__SCAN_IN), 
        .A3(n15397), .A4(n15396), .ZN(n15402) );
  INV_X1 U16929 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15399) );
  NAND4_X1 U16930 ( .A1(SI_2_), .A2(P2_REG2_REG_22__SCAN_IN), .A3(n15399), 
        .A4(n15398), .ZN(n15400) );
  OR4_X1 U16931 ( .A1(SI_8_), .A2(n15145), .A3(P3_REG3_REG_17__SCAN_IN), .A4(
        n15400), .ZN(n15401) );
  NOR4_X1 U16932 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15403), .A3(n15402), .A4(
        n15401), .ZN(n15426) );
  NAND4_X1 U16933 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(P3_REG3_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_26__SCAN_IN), .A4(n15404), .ZN(n15412) );
  NAND4_X1 U16934 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15405), .A3(n11073), 
        .A4(n13585), .ZN(n15411) );
  NAND4_X1 U16935 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), 
        .A3(n15407), .A4(n15406), .ZN(n15410) );
  NAND4_X1 U16936 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .A3(n15408), .A4(n12911), .ZN(n15409) );
  NOR4_X1 U16937 ( .A1(n15412), .A2(n15411), .A3(n15410), .A4(n15409), .ZN(
        n15425) );
  NAND4_X1 U16938 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), .A3(P1_REG0_REG_28__SCAN_IN), .A4(n15413), .ZN(n15414) );
  NOR3_X1 U16939 ( .A1(n15415), .A2(P3_IR_REG_21__SCAN_IN), .A3(n15414), .ZN(
        n15416) );
  NAND3_X1 U16940 ( .A1(n15416), .A2(P1_DATAO_REG_0__SCAN_IN), .A3(
        P3_REG0_REG_29__SCAN_IN), .ZN(n15423) );
  NAND4_X1 U16941 ( .A1(SI_3_), .A2(n15419), .A3(n15418), .A4(n15417), .ZN(
        n15422) );
  NAND4_X1 U16942 ( .A1(SI_19_), .A2(P2_REG2_REG_28__SCAN_IN), .A3(
        P3_DATAO_REG_2__SCAN_IN), .A4(n15420), .ZN(n15421) );
  NOR3_X1 U16943 ( .A1(n15423), .A2(n15422), .A3(n15421), .ZN(n15424) );
  NAND4_X1 U16944 ( .A1(n15427), .A2(n15426), .A3(n15425), .A4(n15424), .ZN(
        n15428) );
  NOR4_X1 U16945 ( .A1(n15431), .A2(n15430), .A3(n15429), .A4(n15428), .ZN(
        n15432) );
  NAND4_X1 U16946 ( .A1(n15435), .A2(n15434), .A3(n15433), .A4(n15432), .ZN(
        n15436) );
  XNOR2_X1 U16947 ( .A(n15437), .B(n15436), .ZN(U29) );
  XNOR2_X1 U16948 ( .A(n15438), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  XOR2_X1 U16949 ( .A(n15440), .B(n15439), .Z(SUB_1596_U59) );
  AOI21_X1 U16950 ( .B1(n15442), .B2(n15441), .A(n15450), .ZN(SUB_1596_U53) );
  XOR2_X1 U16951 ( .A(n15443), .B(n15444), .Z(SUB_1596_U56) );
  AOI21_X1 U16952 ( .B1(n15447), .B2(n15446), .A(n15445), .ZN(n15448) );
  XNOR2_X1 U16953 ( .A(n15448), .B(n8967), .ZN(SUB_1596_U60) );
  XOR2_X1 U16954 ( .A(n15450), .B(n15449), .Z(SUB_1596_U5) );
  INV_X1 U7325 ( .A(n6893), .ZN(n8256) );
  NAND2_X2 U10124 ( .A1(n8899), .A2(n9161), .ZN(n7832) );
  CLKBUF_X1 U7308 ( .A(n7196), .Z(n6923) );
  CLKBUF_X1 U7309 ( .A(n7857), .Z(n6943) );
  INV_X1 U7339 ( .A(n7645), .ZN(n8361) );
  XNOR2_X1 U7375 ( .A(n11113), .B(n11112), .ZN(n12384) );
  CLKBUF_X1 U7601 ( .A(n7855), .Z(n8257) );
  CLKBUF_X1 U9514 ( .A(n8306), .Z(n6527) );
  CLKBUF_X2 U9538 ( .A(n6538), .Z(n6535) );
endmodule

