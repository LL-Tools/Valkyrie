

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339;

  AND2_X1 U11076 ( .A1(n11338), .A2(n11336), .ZN(n13573) );
  NAND2_X1 U11077 ( .A1(n13616), .A2(n11047), .ZN(n19263) );
  AND2_X1 U11078 ( .A1(n11201), .A2(n11028), .ZN(n19294) );
  AND2_X1 U11079 ( .A1(n13630), .A2(n14921), .ZN(n19309) );
  INV_X1 U11080 ( .A(n11028), .ZN(n15128) );
  NOR2_X1 U11081 ( .A1(n13623), .A2(n13622), .ZN(n13632) );
  NOR2_X1 U11082 ( .A1(n13623), .A2(n13620), .ZN(n13630) );
  AND2_X1 U11083 ( .A1(n12406), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12564) );
  AND2_X1 U11084 ( .A1(n11027), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12559) );
  CLKBUF_X1 U11085 ( .A(n12648), .Z(n13023) );
  AND2_X2 U11086 ( .A1(n12533), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12700) );
  CLKBUF_X2 U11087 ( .A(n17618), .Z(n17590) );
  CLKBUF_X2 U11088 ( .A(n11735), .Z(n13306) );
  CLKBUF_X2 U11089 ( .A(n11511), .Z(n12076) );
  CLKBUF_X2 U11090 ( .A(n11623), .Z(n12055) );
  CLKBUF_X2 U11091 ( .A(n12174), .Z(n13307) );
  BUF_X2 U11092 ( .A(n15360), .Z(n17650) );
  CLKBUF_X2 U11093 ( .A(n17456), .Z(n10998) );
  INV_X2 U11094 ( .A(n11386), .ZN(n20172) );
  CLKBUF_X3 U11095 ( .A(n15348), .Z(n10994) );
  BUF_X1 U11096 ( .A(n12464), .Z(n14806) );
  INV_X2 U11097 ( .A(n20142), .ZN(n17681) );
  INV_X1 U11098 ( .A(n13348), .ZN(n11549) );
  AND4_X1 U11099 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11547) );
  INV_X1 U11100 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21232) );
  CLKBUF_X1 U11101 ( .A(n12365), .Z(n19353) );
  AND2_X1 U11102 ( .A1(n11096), .A2(n14238), .ZN(n12174) );
  AND2_X1 U11103 ( .A1(n11335), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11413) );
  INV_X1 U11104 ( .A(n13975), .ZN(n12397) );
  NAND2_X1 U11105 ( .A1(n12381), .A2(n12380), .ZN(n13975) );
  CLKBUF_X1 U11106 ( .A(n12407), .Z(n11024) );
  BUF_X2 U11107 ( .A(n12405), .Z(n10987) );
  INV_X2 U11108 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12373) );
  CLKBUF_X2 U11109 ( .A(n12407), .Z(n11000) );
  CLKBUF_X1 U11110 ( .A(n19106), .Z(n10969) );
  NOR2_X1 U11111 ( .A1(n18721), .A2(n18687), .ZN(n19106) );
  OAI22_X1 U11112 ( .A1(n20023), .A2(n14601), .B1(n16963), .B2(n14600), .ZN(
        n22094) );
  NAND2_X2 U11113 ( .A1(n19979), .A2(n14544), .ZN(n14601) );
  OAI22_X1 U11114 ( .A1(n20021), .A2(n14601), .B1(n16964), .B2(n14600), .ZN(
        n22056) );
  NAND2_X2 U11115 ( .A1(n19979), .A2(n15202), .ZN(n14600) );
  OR2_X1 U11116 ( .A1(n19218), .A2(n13641), .ZN(n13644) );
  AND3_X1 U11117 ( .A1(n11556), .A2(n14316), .A3(n14234), .ZN(n11565) );
  AND2_X1 U11118 ( .A1(n11411), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11418) );
  CLKBUF_X2 U11119 ( .A(n11710), .Z(n13305) );
  AND2_X1 U11120 ( .A1(n15835), .A2(n13551), .ZN(n11347) );
  AND2_X1 U11121 ( .A1(n14233), .A2(n11546), .ZN(n11569) );
  INV_X1 U11122 ( .A(n12404), .ZN(n10973) );
  INV_X1 U11123 ( .A(n12530), .ZN(n15485) );
  AND2_X2 U11124 ( .A1(n11420), .A2(n14460), .ZN(n11029) );
  OR2_X1 U11125 ( .A1(n15861), .A2(n15860), .ZN(n19956) );
  CLKBUF_X2 U11126 ( .A(n12034), .Z(n14448) );
  AND4_X1 U11127 ( .A1(n11435), .A2(n11433), .A3(n11434), .A4(n11432), .ZN(
        n11051) );
  AND2_X1 U11128 ( .A1(n12395), .A2(n13269), .ZN(n12392) );
  NOR2_X2 U11129 ( .A1(n13975), .A2(n12440), .ZN(n12441) );
  AND2_X2 U11130 ( .A1(n13886), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12532) );
  INV_X1 U11131 ( .A(n17663), .ZN(n17469) );
  NOR2_X2 U11132 ( .A1(n14529), .A2(n14708), .ZN(n14854) );
  INV_X1 U11133 ( .A(n12282), .ZN(n14229) );
  NAND2_X1 U11134 ( .A1(n12393), .A2(n12392), .ZN(n12456) );
  CLKBUF_X2 U11135 ( .A(n13142), .Z(n13242) );
  NOR2_X1 U11136 ( .A1(n11046), .A2(n13994), .ZN(n14002) );
  NOR2_X2 U11137 ( .A1(n14537), .A2(n14538), .ZN(n14539) );
  INV_X1 U11138 ( .A(n17369), .ZN(n17662) );
  CLKBUF_X3 U11139 ( .A(n17364), .Z(n10991) );
  NAND2_X1 U11140 ( .A1(n20759), .A2(n20772), .ZN(n20117) );
  INV_X1 U11141 ( .A(n14356), .ZN(n13464) );
  AND2_X1 U11142 ( .A1(n13563), .A2(n15848), .ZN(n11038) );
  BUF_X1 U11143 ( .A(n19935), .Z(n10972) );
  NAND2_X1 U11144 ( .A1(n14229), .A2(n11476), .ZN(n11558) );
  NOR2_X1 U11146 ( .A1(n16133), .A2(n16126), .ZN(n16125) );
  NAND2_X1 U11147 ( .A1(n14614), .A2(n14613), .ZN(n14537) );
  AOI211_X1 U11148 ( .C1(n19115), .C2(n18606), .A(n14029), .B(n15467), .ZN(
        n14030) );
  NAND3_X1 U11149 ( .A1(n12396), .A2(n12395), .A3(n12426), .ZN(n13955) );
  BUF_X1 U11150 ( .A(n20393), .Z(n20528) );
  INV_X1 U11151 ( .A(n20363), .ZN(n20463) );
  INV_X1 U11152 ( .A(n18156), .ZN(n18166) );
  INV_X1 U11153 ( .A(n13364), .ZN(n15446) );
  NOR2_X2 U11154 ( .A1(n15540), .A2(n15542), .ZN(n15527) );
  NAND2_X1 U11155 ( .A1(n14531), .A2(n14530), .ZN(n14529) );
  NAND2_X2 U11156 ( .A1(n11650), .A2(n14548), .ZN(n14973) );
  NAND2_X1 U11157 ( .A1(n12877), .A2(n14822), .ZN(n14096) );
  INV_X2 U11158 ( .A(n18376), .ZN(n18584) );
  INV_X1 U11159 ( .A(n18291), .ZN(n12459) );
  AOI21_X1 U11160 ( .B1(n16271), .B2(n15459), .A(n14032), .ZN(n15462) );
  INV_X1 U11161 ( .A(n21122), .ZN(n21175) );
  NAND2_X1 U11162 ( .A1(n13462), .A2(n12209), .ZN(n15508) );
  AOI211_X1 U11163 ( .C1(n19965), .C2(n15774), .A(n15773), .B(n15772), .ZN(
        n15775) );
  INV_X1 U11164 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22008) );
  AOI21_X1 U11165 ( .B1(n16623), .B2(n16592), .A(n16616), .ZN(n16608) );
  INV_X1 U11166 ( .A(n18015), .ZN(n18153) );
  AND3_X1 U11167 ( .A1(n11031), .A2(n11552), .A3(n14715), .ZN(n10970) );
  AND4_X1 U11168 ( .A1(n11431), .A2(n11429), .A3(n11430), .A4(n11428), .ZN(
        n10971) );
  INV_X1 U11169 ( .A(n13550), .ZN(n19935) );
  OAI21_X2 U11170 ( .B1(n11289), .B2(n12515), .A(n11199), .ZN(n11198) );
  OAI21_X4 U11171 ( .B1(n15754), .B2(n15755), .A(n10972), .ZN(n15778) );
  NOR2_X2 U11172 ( .A1(n18117), .A2(n20180), .ZN(n18103) );
  OAI21_X1 U11173 ( .B1(n13482), .B2(n13481), .A(n13480), .ZN(n14285) );
  AND2_X1 U11174 ( .A1(n16180), .A2(n16181), .ZN(n16183) );
  NOR2_X2 U11175 ( .A1(n16200), .A2(n16189), .ZN(n16180) );
  NOR2_X4 U11176 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14463) );
  AND2_X4 U11177 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13886) );
  XNOR2_X2 U11178 ( .A(n13501), .B(n21346), .ZN(n14749) );
  NAND2_X2 U11179 ( .A1(n14622), .A2(n13494), .ZN(n13501) );
  INV_X1 U11180 ( .A(n12404), .ZN(n10974) );
  INV_X1 U11181 ( .A(n12404), .ZN(n10975) );
  INV_X1 U11182 ( .A(n10973), .ZN(n10976) );
  INV_X1 U11185 ( .A(n10974), .ZN(n10979) );
  INV_X1 U11186 ( .A(n10974), .ZN(n10980) );
  INV_X1 U11187 ( .A(n10974), .ZN(n10981) );
  INV_X1 U11188 ( .A(n10975), .ZN(n10982) );
  INV_X1 U11189 ( .A(n10975), .ZN(n10983) );
  INV_X1 U11190 ( .A(n10975), .ZN(n10984) );
  AND2_X2 U11191 ( .A1(n11286), .A2(n12878), .ZN(n12404) );
  XNOR2_X2 U11192 ( .A(n13849), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16350) );
  AND2_X2 U11195 ( .A1(n14768), .A2(n14798), .ZN(n10985) );
  INV_X1 U11196 ( .A(n10985), .ZN(n10986) );
  NOR4_X2 U11197 ( .A1(n17239), .A2(n15394), .A3(n15389), .A4(n20797), .ZN(
        n17732) );
  BUF_X4 U11198 ( .A(n12405), .Z(n10988) );
  BUF_X4 U11199 ( .A(n12405), .Z(n10989) );
  NOR2_X2 U11200 ( .A1(n16310), .A2(n16438), .ZN(n16303) );
  NAND2_X1 U11201 ( .A1(n11205), .A2(n11206), .ZN(n14073) );
  XNOR2_X1 U11202 ( .A(n13461), .B(n13330), .ZN(n13591) );
  NAND2_X1 U11203 ( .A1(n11331), .A2(n11330), .ZN(n15776) );
  OAI21_X1 U11204 ( .B1(n11007), .B2(n11348), .A(n11082), .ZN(n16131) );
  AND2_X1 U11205 ( .A1(n19950), .A2(n13559), .ZN(n15860) );
  NAND2_X1 U11206 ( .A1(n14854), .A2(n11807), .ZN(n14910) );
  NOR2_X1 U11207 ( .A1(n13626), .A2(n14803), .ZN(n11201) );
  AND2_X1 U11208 ( .A1(n14936), .A2(n11085), .ZN(n16066) );
  NOR2_X1 U11209 ( .A1(n11797), .A2(n11796), .ZN(n11810) );
  INV_X1 U11210 ( .A(n18006), .ZN(n17894) );
  OAI21_X1 U11211 ( .B1(n15161), .B2(n14848), .A(n12504), .ZN(n14373) );
  INV_X1 U11212 ( .A(n15161), .ZN(n17132) );
  OR2_X1 U11213 ( .A1(n14483), .A2(n11277), .ZN(n16642) );
  NAND2_X1 U11214 ( .A1(n12474), .A2(n12493), .ZN(n12518) );
  NAND2_X1 U11215 ( .A1(n14481), .A2(n14480), .ZN(n14483) );
  NAND2_X1 U11216 ( .A1(n11267), .A2(n11264), .ZN(n14481) );
  NAND2_X1 U11217 ( .A1(n20782), .A2(n20744), .ZN(n21206) );
  NOR2_X1 U11218 ( .A1(n12983), .A2(n12982), .ZN(n14860) );
  INV_X2 U11219 ( .A(n17976), .ZN(n18051) );
  CLKBUF_X1 U11220 ( .A(n12432), .Z(n14011) );
  INV_X4 U11221 ( .A(n20796), .ZN(n20800) );
  INV_X4 U11222 ( .A(n13989), .ZN(n13820) );
  CLKBUF_X2 U11223 ( .A(n12459), .Z(n19574) );
  NAND3_X1 U11224 ( .A1(n15376), .A2(n15375), .A3(n15374), .ZN(n20796) );
  INV_X2 U11225 ( .A(n12394), .ZN(n13269) );
  NOR2_X2 U11227 ( .A1(n13348), .A2(n11553), .ZN(n14715) );
  AND4_X1 U11228 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11493) );
  INV_X2 U11229 ( .A(n21199), .ZN(n10990) );
  CLKBUF_X3 U11230 ( .A(n17652), .Z(n10997) );
  CLKBUF_X2 U11231 ( .A(n11602), .Z(n11584) );
  CLKBUF_X2 U11232 ( .A(n11663), .Z(n11582) );
  CLKBUF_X3 U11233 ( .A(n17341), .Z(n10996) );
  CLKBUF_X2 U11234 ( .A(n11669), .Z(n11589) );
  CLKBUF_X2 U11235 ( .A(n11601), .Z(n11670) );
  CLKBUF_X2 U11236 ( .A(n11664), .Z(n11711) );
  CLKBUF_X2 U11237 ( .A(n11671), .Z(n13313) );
  INV_X2 U11238 ( .A(n15481), .ZN(n12533) );
  CLKBUF_X2 U11239 ( .A(n11022), .Z(n11023) );
  BUF_X2 U11240 ( .A(n11022), .Z(n11001) );
  INV_X1 U11241 ( .A(n22337), .ZN(n22339) );
  INV_X1 U11242 ( .A(n10999), .ZN(n10992) );
  CLKBUF_X2 U11243 ( .A(n19811), .Z(n21288) );
  CLKBUF_X2 U11244 ( .A(n11622), .Z(n11838) );
  BUF_X2 U11245 ( .A(n11583), .Z(n11899) );
  AND2_X1 U11246 ( .A1(n11410), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11096) );
  NOR2_X2 U11247 ( .A1(n20759), .A2(n20772), .ZN(n20775) );
  NAND2_X1 U11248 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20773) );
  AOI21_X1 U11249 ( .B1(n16445), .B2(n18612), .A(n16444), .ZN(n16446) );
  AOI21_X1 U11250 ( .B1(n15462), .B2(n18612), .A(n15461), .ZN(n15463) );
  NAND2_X1 U11251 ( .A1(n11211), .A2(n11212), .ZN(n16310) );
  NAND2_X1 U11252 ( .A1(n11211), .A2(n11209), .ZN(n11213) );
  INV_X1 U11253 ( .A(n16331), .ZN(n11211) );
  AOI21_X1 U11254 ( .B1(n15475), .B2(n15474), .A(n15473), .ZN(n15497) );
  NAND2_X1 U11255 ( .A1(n16335), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16331) );
  NAND2_X1 U11256 ( .A1(n16359), .A2(n16358), .ZN(n16409) );
  INV_X1 U11257 ( .A(n14073), .ZN(n11149) );
  NOR2_X1 U11258 ( .A1(n15445), .A2(n15659), .ZN(n11243) );
  INV_X1 U11259 ( .A(n15620), .ZN(n15767) );
  OR2_X1 U11260 ( .A1(n13573), .A2(n13572), .ZN(n13578) );
  NOR2_X1 U11261 ( .A1(n16117), .A2(n11392), .ZN(n12828) );
  OR2_X1 U11262 ( .A1(n14051), .A2(n12207), .ZN(n15620) );
  NOR2_X1 U11263 ( .A1(n15760), .A2(n15759), .ZN(n15762) );
  AOI211_X1 U11264 ( .C1(n19976), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21416), .B(n19944), .ZN(n19945) );
  AOI211_X1 U11265 ( .C1(n18552), .C2(n18611), .A(n16453), .B(n16452), .ZN(
        n16454) );
  XNOR2_X1 U11266 ( .A(n14002), .B(n14001), .ZN(n18579) );
  NAND2_X1 U11267 ( .A1(n16718), .A2(n11037), .ZN(n16653) );
  NAND2_X1 U11268 ( .A1(n16715), .A2(n16716), .ZN(n16718) );
  XNOR2_X1 U11269 ( .A(n11046), .B(n13247), .ZN(n15504) );
  NAND2_X1 U11270 ( .A1(n16093), .A2(n11046), .ZN(n18564) );
  OR2_X1 U11271 ( .A1(n16101), .A2(n16112), .ZN(n18535) );
  INV_X1 U11272 ( .A(n11007), .ZN(n16138) );
  NAND2_X1 U11273 ( .A1(n15206), .A2(n15212), .ZN(n15210) );
  AND2_X1 U11274 ( .A1(n13687), .A2(n13686), .ZN(n15068) );
  NAND2_X1 U11275 ( .A1(n15869), .A2(n13551), .ZN(n11346) );
  CLKBUF_X1 U11276 ( .A(n15869), .Z(n15870) );
  AND2_X2 U11277 ( .A1(n15593), .A2(n15592), .ZN(n15595) );
  NAND2_X1 U11278 ( .A1(n15872), .A2(n15871), .ZN(n15869) );
  AND2_X1 U11279 ( .A1(n17934), .A2(n21029), .ZN(n17974) );
  OR2_X1 U11280 ( .A1(n15289), .A2(n15292), .ZN(n15293) );
  OR2_X1 U11281 ( .A1(n11347), .A2(n11345), .ZN(n11344) );
  NAND2_X2 U11282 ( .A1(n14903), .A2(n14941), .ZN(n14940) );
  NAND2_X1 U11283 ( .A1(n19929), .A2(n11055), .ZN(n15244) );
  AND2_X1 U11284 ( .A1(n16183), .A2(n13251), .ZN(n13255) );
  XNOR2_X1 U11285 ( .A(n16183), .B(n13251), .ZN(n18563) );
  NAND2_X1 U11286 ( .A1(n13508), .A2(n19912), .ZN(n11342) );
  INV_X1 U11287 ( .A(n14910), .ZN(n11364) );
  OAI211_X1 U11288 ( .C1(n13652), .C2(n13651), .A(n13644), .B(n13643), .ZN(
        n11193) );
  INV_X1 U11289 ( .A(n14911), .ZN(n11818) );
  OR2_X1 U11290 ( .A1(n13550), .A2(n13552), .ZN(n19960) );
  NAND2_X1 U11291 ( .A1(n11176), .A2(n13535), .ZN(n13537) );
  AOI21_X1 U11292 ( .B1(n13530), .B2(n11942), .A(n11817), .ZN(n14911) );
  OR2_X1 U11293 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  AOI22_X1 U11294 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19309), .B1(
        n13699), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U11295 ( .A1(n13616), .A2(n13607), .ZN(n19231) );
  NAND2_X1 U11296 ( .A1(n13616), .A2(n13597), .ZN(n19248) );
  OAI211_X1 U11297 ( .C1(n13516), .C2(n11897), .A(n11805), .B(n11804), .ZN(
        n14855) );
  NAND2_X1 U11298 ( .A1(n13615), .A2(n11047), .ZN(n19170) );
  NAND2_X1 U11299 ( .A1(n13616), .A2(n11050), .ZN(n17047) );
  NAND2_X1 U11300 ( .A1(n13615), .A2(n13607), .ZN(n19135) );
  NAND2_X1 U11301 ( .A1(n13615), .A2(n13597), .ZN(n19155) );
  NOR2_X1 U11302 ( .A1(n15631), .A2(n15556), .ZN(n15557) );
  NAND2_X1 U11303 ( .A1(n11787), .A2(n11808), .ZN(n13520) );
  NAND2_X1 U11304 ( .A1(n11810), .A2(n11809), .ZN(n13542) );
  OR2_X1 U11305 ( .A1(n11797), .A2(n11796), .ZN(n11787) );
  OAI21_X1 U11306 ( .B1(n13621), .B2(n14848), .A(n12522), .ZN(n12524) );
  NAND2_X1 U11307 ( .A1(n11173), .A2(n11760), .ZN(n11797) );
  OAI21_X1 U11308 ( .B1(n18090), .B2(n11317), .A(n11315), .ZN(n18053) );
  INV_X1 U11309 ( .A(n13621), .ZN(n14803) );
  NAND2_X1 U11310 ( .A1(n12497), .A2(n12496), .ZN(n14405) );
  NAND2_X1 U11311 ( .A1(n14355), .A2(n13492), .ZN(n13493) );
  INV_X1 U11312 ( .A(n18171), .ZN(n18161) );
  NAND2_X2 U11313 ( .A1(n15260), .A2(n14510), .ZN(n15725) );
  CLKBUF_X2 U11314 ( .A(n13610), .Z(n11028) );
  NAND2_X1 U11315 ( .A1(n11723), .A2(n11722), .ZN(n14522) );
  XNOR2_X1 U11316 ( .A(n13606), .B(n12495), .ZN(n13610) );
  NAND2_X1 U11317 ( .A1(n16115), .A2(n16103), .ZN(n11232) );
  NAND2_X1 U11318 ( .A1(n14285), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14284) );
  NAND2_X1 U11319 ( .A1(n12501), .A2(n12494), .ZN(n12517) );
  NAND2_X1 U11320 ( .A1(n12501), .A2(n12500), .ZN(n15161) );
  XNOR2_X1 U11321 ( .A(n12493), .B(n12494), .ZN(n13606) );
  XNOR2_X1 U11322 ( .A(n14295), .B(n21960), .ZN(n14445) );
  AND2_X1 U11323 ( .A1(n14295), .A2(n11660), .ZN(n21961) );
  XNOR2_X1 U11324 ( .A(n17722), .B(n17721), .ZN(n18114) );
  AOI21_X2 U11325 ( .B1(n13142), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12473), .ZN(n12493) );
  OR2_X1 U11326 ( .A1(n14861), .A2(n11268), .ZN(n11267) );
  INV_X1 U11327 ( .A(n12469), .ZN(n12494) );
  NOR2_X2 U11328 ( .A1(n21224), .A2(n21206), .ZN(n21122) );
  INV_X1 U11329 ( .A(n13152), .ZN(n11288) );
  NAND2_X1 U11330 ( .A1(n12511), .A2(n12510), .ZN(n13153) );
  OAI21_X1 U11331 ( .B1(n12507), .B2(n14159), .A(n12477), .ZN(n12481) );
  XNOR2_X1 U11332 ( .A(n17965), .B(n17964), .ZN(n20393) );
  OR2_X1 U11333 ( .A1(n12983), .A2(n12979), .ZN(n14339) );
  INV_X2 U11334 ( .A(n13143), .ZN(n13243) );
  AND2_X1 U11335 ( .A1(n12431), .A2(n12430), .ZN(n12454) );
  INV_X2 U11336 ( .A(n20063), .ZN(n20112) );
  OR2_X1 U11337 ( .A1(n14017), .A2(n18286), .ZN(n12453) );
  AOI21_X1 U11338 ( .B1(n14435), .B2(n12978), .A(n12977), .ZN(n12983) );
  NAND2_X1 U11339 ( .A1(n14437), .A2(n14436), .ZN(n14435) );
  NOR2_X2 U11340 ( .A1(n20811), .A2(n21090), .ZN(n17976) );
  AND2_X1 U11341 ( .A1(n11566), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11647) );
  AND2_X1 U11342 ( .A1(n11570), .A2(n11560), .ZN(n11561) );
  AND2_X1 U11343 ( .A1(n14377), .A2(n14378), .ZN(n14376) );
  NAND3_X1 U11344 ( .A1(n15393), .A2(n15418), .A3(n18802), .ZN(n15397) );
  OAI21_X1 U11345 ( .B1(n15425), .B2(n18883), .A(n15389), .ZN(n11093) );
  NAND2_X1 U11346 ( .A1(n12210), .A2(n14715), .ZN(n14234) );
  AND2_X1 U11347 ( .A1(n11614), .A2(n11613), .ZN(n11642) );
  NOR2_X1 U11348 ( .A1(n11575), .A2(n19986), .ZN(n11576) );
  NAND2_X1 U11349 ( .A1(n12427), .A2(n12426), .ZN(n14018) );
  OR2_X1 U11350 ( .A1(n11609), .A2(n11662), .ZN(n11596) );
  AND2_X1 U11351 ( .A1(n11523), .A2(n14578), .ZN(n13581) );
  NAND2_X1 U11352 ( .A1(n12459), .A2(n19628), .ZN(n12877) );
  CLKBUF_X2 U11353 ( .A(n14449), .Z(n11031) );
  BUF_X2 U11354 ( .A(n13269), .Z(n13989) );
  INV_X2 U11355 ( .A(n11407), .ZN(n13252) );
  AND2_X1 U11356 ( .A1(n12273), .A2(n14578), .ZN(n11548) );
  OR2_X1 U11357 ( .A1(n11629), .A2(n11628), .ZN(n13483) );
  AND2_X2 U11358 ( .A1(n11549), .A2(n11553), .ZN(n14214) );
  OR2_X1 U11359 ( .A1(n11595), .A2(n11594), .ZN(n13484) );
  INV_X1 U11360 ( .A(n12419), .ZN(n12415) );
  OR2_X1 U11361 ( .A1(n11608), .A2(n11607), .ZN(n13543) );
  OR2_X1 U11362 ( .A1(n12974), .A2(n12973), .ZN(n13668) );
  AND2_X2 U11363 ( .A1(n11571), .A2(n13348), .ZN(n13364) );
  AND2_X1 U11364 ( .A1(n14307), .A2(n11571), .ZN(n12273) );
  INV_X1 U11365 ( .A(n11574), .ZN(n11522) );
  NAND4_X2 U11366 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n14578) );
  NAND2_X2 U11367 ( .A1(n11172), .A2(n11171), .ZN(n12394) );
  INV_X2 U11368 ( .A(U212), .ZN(n10993) );
  NAND2_X1 U11369 ( .A1(n12327), .A2(n12373), .ZN(n12328) );
  NAND2_X1 U11370 ( .A1(n12335), .A2(n12334), .ZN(n12342) );
  NAND2_X1 U11371 ( .A1(n12322), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12329) );
  NAND2_X2 U11372 ( .A1(U214), .A2(n19989), .ZN(n20050) );
  AND2_X2 U11373 ( .A1(n11035), .A2(n11057), .ZN(n14307) );
  OR2_X2 U11374 ( .A1(n11506), .A2(n11505), .ZN(n11571) );
  AND4_X1 U11375 ( .A1(n11417), .A2(n11416), .A3(n11415), .A4(n11414), .ZN(
        n11427) );
  AND4_X1 U11376 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  AND4_X1 U11377 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11472) );
  AND4_X1 U11378 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11541) );
  AND3_X1 U11379 ( .A1(n11539), .A2(n11538), .A3(n11409), .ZN(n11540) );
  AND4_X1 U11380 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(
        n11496) );
  AND4_X1 U11381 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11453) );
  AND4_X1 U11382 ( .A1(n11484), .A2(n11483), .A3(n11482), .A4(n11481), .ZN(
        n11495) );
  AND4_X1 U11383 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11542) );
  AND4_X1 U11384 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11454) );
  AND4_X1 U11385 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11452) );
  AND4_X1 U11386 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11494) );
  AND4_X1 U11387 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11455) );
  AND4_X1 U11388 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11543) );
  AND4_X1 U11389 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11475) );
  AND4_X1 U11390 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11057) );
  BUF_X2 U11391 ( .A(n17618), .Z(n20777) );
  AND4_X1 U11392 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11474) );
  CLKBUF_X3 U11393 ( .A(n17661), .Z(n17702) );
  NOR2_X1 U11394 ( .A1(n21232), .A2(n20764), .ZN(n17618) );
  AND2_X2 U11395 ( .A1(n13584), .A2(n21935), .ZN(n19979) );
  INV_X2 U11396 ( .A(n21739), .ZN(n17226) );
  INV_X2 U11397 ( .A(n18964), .ZN(U215) );
  NAND2_X2 U11398 ( .A1(n17765), .A2(n21277), .ZN(n21199) );
  AND3_X1 U11399 ( .A1(n12311), .A2(n12310), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12315) );
  INV_X2 U11400 ( .A(n11281), .ZN(n14812) );
  INV_X2 U11401 ( .A(n19737), .ZN(n19797) );
  INV_X2 U11402 ( .A(n21736), .ZN(n17237) );
  AND2_X2 U11403 ( .A1(n11413), .A2(n14238), .ZN(n12034) );
  AND2_X2 U11404 ( .A1(n11096), .A2(n14463), .ZN(n11602) );
  AND2_X2 U11405 ( .A1(n11418), .A2(n11096), .ZN(n11664) );
  INV_X1 U11406 ( .A(n18627), .ZN(n18362) );
  AND2_X2 U11407 ( .A1(n13886), .A2(n12878), .ZN(n12530) );
  AND2_X2 U11408 ( .A1(n14463), .A2(n11419), .ZN(n11583) );
  INV_X2 U11409 ( .A(n12368), .ZN(n10999) );
  NAND2_X1 U11410 ( .A1(n21240), .A2(n21232), .ZN(n20774) );
  NAND2_X1 U11411 ( .A1(n20759), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15309) );
  OR3_X1 U11412 ( .A1(n20759), .A2(n20772), .A3(n20773), .ZN(n11386) );
  NOR2_X1 U11413 ( .A1(n21240), .A2(n20759), .ZN(n20758) );
  INV_X1 U11414 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21683) );
  INV_X2 U11415 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11335) );
  INV_X2 U11416 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20759) );
  NOR2_X1 U11417 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11421) );
  AND2_X1 U11418 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14450) );
  INV_X1 U11419 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14798) );
  INV_X1 U11420 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12878) );
  XNOR2_X1 U11421 ( .A(n13542), .B(n11813), .ZN(n13530) );
  NAND2_X1 U11422 ( .A1(n13542), .A2(n13541), .ZN(n13550) );
  CLKBUF_X1 U11423 ( .A(n13964), .Z(n11002) );
  BUF_X1 U11424 ( .A(n16373), .Z(n11003) );
  NOR2_X2 U11425 ( .A1(n18074), .A2(n21162), .ZN(n18014) );
  NOR2_X2 U11426 ( .A1(n21254), .A2(n21279), .ZN(n21282) );
  CLKBUF_X1 U11427 ( .A(n13938), .Z(n11004) );
  CLKBUF_X1 U11428 ( .A(n14919), .Z(n11005) );
  OAI22_X1 U11429 ( .A1(n19170), .A2(n13618), .B1(n19263), .B2(n13617), .ZN(
        n13619) );
  CLKBUF_X1 U11430 ( .A(n15206), .Z(n11006) );
  NOR2_X2 U11431 ( .A1(n15149), .A2(n15207), .ZN(n15206) );
  NOR2_X2 U11432 ( .A1(n20706), .A2(n20717), .ZN(n20702) );
  AND2_X1 U11433 ( .A1(n11286), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11022) );
  AND2_X1 U11434 ( .A1(n11286), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12407) );
  NOR2_X2 U11435 ( .A1(n19937), .A2(n19936), .ZN(n19943) );
  NOR2_X2 U11436 ( .A1(n13679), .A2(n13680), .ZN(n13674) );
  AND4_X1 U11437 ( .A1(n13673), .A2(n13688), .A3(n13674), .A4(n11162), .ZN(
        n13757) );
  NAND2_X1 U11438 ( .A1(n13796), .A2(n11169), .ZN(n13800) );
  NOR3_X2 U11439 ( .A1(n13880), .A2(n13596), .A3(n16443), .ZN(n16267) );
  INV_X1 U11440 ( .A(n16651), .ZN(n11147) );
  NAND2_X1 U11441 ( .A1(n11205), .A2(n11202), .ZN(n16347) );
  NAND2_X1 U11442 ( .A1(n18291), .A2(n14009), .ZN(n14822) );
  INV_X1 U11443 ( .A(n14009), .ZN(n19628) );
  NAND2_X1 U11444 ( .A1(n14009), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18290) );
  AND2_X1 U11445 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12538) );
  AND2_X2 U11446 ( .A1(n12878), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14768) );
  NOR2_X1 U11447 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12539) );
  AND2_X2 U11448 ( .A1(n16144), .A2(n16145), .ZN(n11007) );
  NAND2_X1 U11449 ( .A1(n11004), .A2(n13937), .ZN(n11008) );
  NAND2_X1 U11450 ( .A1(n13938), .A2(n13937), .ZN(n16429) );
  OAI21_X2 U11451 ( .B1(n13489), .B2(n13481), .A(n13488), .ZN(n13490) );
  NAND3_X1 U11452 ( .A1(n11342), .A2(n13517), .A3(n11341), .ZN(n19918) );
  NAND2_X2 U11453 ( .A1(n13615), .A2(n11050), .ZN(n19144) );
  OR2_X1 U11454 ( .A1(n16705), .A2(n16602), .ZN(n11009) );
  NAND2_X1 U11455 ( .A1(n16601), .A2(n11009), .ZN(n16605) );
  OAI21_X2 U11456 ( .B1(n15809), .B2(n13566), .A(n10972), .ZN(n15966) );
  NAND2_X4 U11457 ( .A1(n11175), .A2(n11038), .ZN(n15809) );
  NAND2_X2 U11458 ( .A1(n11758), .A2(n11683), .ZN(n14519) );
  NAND2_X2 U11459 ( .A1(n13567), .A2(n15966), .ZN(n15754) );
  OR2_X1 U11460 ( .A1(n16598), .A2(n16730), .ZN(n11010) );
  NAND2_X1 U11461 ( .A1(n11010), .A2(n16597), .ZN(P2_U3029) );
  BUF_X4 U11462 ( .A(n13623), .Z(n15096) );
  OR4_X1 U11463 ( .A1(n14084), .A2(n16599), .A3(n14083), .A4(n14082), .ZN(
        P2_U2998) );
  NOR2_X2 U11464 ( .A1(n14883), .A2(n14884), .ZN(n14695) );
  NAND2_X1 U11465 ( .A1(n15249), .A2(n15288), .ZN(n11011) );
  NOR2_X2 U11466 ( .A1(n11011), .A2(n11012), .ZN(n15593) );
  OR2_X1 U11467 ( .A1(n15652), .A2(n15292), .ZN(n11012) );
  NAND2_X1 U11468 ( .A1(n15527), .A2(n15528), .ZN(n11013) );
  XNOR2_X1 U11469 ( .A(n11567), .B(n11647), .ZN(n11014) );
  INV_X1 U11470 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11015) );
  NAND2_X2 U11471 ( .A1(n11562), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11651) );
  XNOR2_X1 U11472 ( .A(n11567), .B(n11647), .ZN(n14628) );
  AND2_X2 U11473 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14460) );
  NAND2_X2 U11474 ( .A1(n15831), .A2(n11403), .ZN(n11175) );
  AND2_X2 U11475 ( .A1(n11096), .A2(n11420), .ZN(n11671) );
  AND2_X2 U11476 ( .A1(n12925), .A2(n13820), .ZN(n12964) );
  AOI21_X1 U11477 ( .B1(n15831), .B2(n19957), .A(n15858), .ZN(n19948) );
  NOR2_X4 U11478 ( .A1(n15133), .A2(n15152), .ZN(n14079) );
  NAND2_X2 U11479 ( .A1(n15244), .A2(n13549), .ZN(n15872) );
  AND2_X1 U11480 ( .A1(n11096), .A2(n11420), .ZN(n11016) );
  OR2_X1 U11481 ( .A1(n14048), .A2(n11380), .ZN(n13462) );
  NAND2_X2 U11482 ( .A1(n14750), .A2(n13502), .ZN(n19914) );
  NAND2_X2 U11483 ( .A1(n14749), .A2(n14751), .ZN(n14750) );
  NOR2_X2 U11484 ( .A1(n14696), .A2(n12571), .ZN(n14903) );
  INV_X1 U11485 ( .A(n11553), .ZN(n11017) );
  INV_X1 U11486 ( .A(n11553), .ZN(n11018) );
  XNOR2_X2 U11487 ( .A(n15736), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15908) );
  XNOR2_X1 U11489 ( .A(n11696), .B(n11695), .ZN(n13482) );
  NAND2_X2 U11490 ( .A1(n11733), .A2(n11732), .ZN(n14530) );
  AND2_X2 U11491 ( .A1(n11420), .A2(n14460), .ZN(n11824) );
  AND2_X1 U11492 ( .A1(n11420), .A2(n14460), .ZN(n11030) );
  AND2_X1 U11493 ( .A1(n11096), .A2(n14238), .ZN(n11021) );
  NAND2_X2 U11494 ( .A1(n11748), .A2(n11725), .ZN(n14521) );
  NAND2_X2 U11495 ( .A1(n11099), .A2(n11098), .ZN(n11758) );
  NOR2_X2 U11496 ( .A1(n15210), .A2(n11359), .ZN(n16144) );
  NOR2_X2 U11497 ( .A1(n12276), .A2(n14570), .ZN(n14122) );
  INV_X1 U11498 ( .A(n14448), .ZN(n11025) );
  INV_X2 U11499 ( .A(n12368), .ZN(n11026) );
  INV_X2 U11500 ( .A(n12368), .ZN(n11027) );
  NAND2_X2 U11501 ( .A1(n12538), .A2(n14798), .ZN(n12368) );
  NAND2_X4 U11502 ( .A1(n12364), .A2(n12363), .ZN(n12425) );
  NOR2_X2 U11503 ( .A1(n11097), .A2(n11555), .ZN(n12210) );
  XNOR2_X2 U11504 ( .A(n11617), .B(n11616), .ZN(n11698) );
  OAI211_X2 U11505 ( .C1(n16097), .C2(n16109), .A(n16099), .B(n16106), .ZN(
        n15475) );
  AND2_X2 U11506 ( .A1(n15229), .A2(n15250), .ZN(n15249) );
  NOR2_X2 U11507 ( .A1(n15196), .A2(n11382), .ZN(n15229) );
  NOR2_X2 U11508 ( .A1(n15569), .A2(n15627), .ZN(n15554) );
  XNOR2_X2 U11509 ( .A(n13489), .B(n11642), .ZN(n11688) );
  OAI21_X4 U11510 ( .B1(n14973), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11596), 
        .ZN(n13489) );
  OAI222_X1 U11511 ( .A1(n15659), .A2(n15771), .B1(n15621), .B2(n19911), .C1(
        n15929), .C2(n15657), .ZN(P1_U2845) );
  AOI21_X2 U11512 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n15740) );
  OAI21_X1 U11513 ( .B1(n15527), .B2(n15528), .A(n11013), .ZN(n15771) );
  AND2_X4 U11514 ( .A1(n11413), .A2(n14463), .ZN(n11710) );
  NOR2_X1 U11515 ( .A1(n13636), .A2(n13635), .ZN(n13637) );
  NAND2_X1 U11516 ( .A1(n18124), .A2(n17719), .ZN(n17722) );
  INV_X1 U11517 ( .A(n11758), .ZN(n11173) );
  NAND2_X1 U11518 ( .A1(n11017), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11661) );
  INV_X1 U11519 ( .A(n13275), .ZN(n13714) );
  AOI21_X1 U11520 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19175), .A(
        n12872), .ZN(n12890) );
  OAI22_X1 U11521 ( .A1(n21244), .A2(n21241), .B1(n21242), .B2(n21243), .ZN(
        n11113) );
  AND2_X1 U11522 ( .A1(n11372), .A2(n15571), .ZN(n11371) );
  INV_X1 U11523 ( .A(n15118), .ZN(n11864) );
  AOI21_X1 U11524 ( .B1(n15872), .B2(n11052), .A(n11343), .ZN(n13557) );
  NAND2_X1 U11525 ( .A1(n11344), .A2(n10972), .ZN(n11343) );
  INV_X1 U11526 ( .A(n14321), .ZN(n13439) );
  NAND2_X1 U11527 ( .A1(n13530), .A2(n13521), .ZN(n11176) );
  NAND2_X1 U11528 ( .A1(n11635), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11662) );
  NOR2_X1 U11529 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12711) );
  NOR2_X1 U11530 ( .A1(n18291), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U11531 ( .A1(n11294), .A2(n11295), .ZN(n11292) );
  NOR2_X1 U11532 ( .A1(n11279), .A2(n15036), .ZN(n11278) );
  NAND2_X1 U11533 ( .A1(n11270), .A2(n11269), .ZN(n11268) );
  INV_X1 U11534 ( .A(n14482), .ZN(n11269) );
  INV_X1 U11535 ( .A(n11271), .ZN(n11270) );
  NOR2_X1 U11536 ( .A1(n14482), .A2(n13015), .ZN(n11266) );
  NOR2_X1 U11537 ( .A1(n11194), .A2(n11193), .ZN(n11192) );
  INV_X1 U11538 ( .A(n13605), .ZN(n11140) );
  NOR2_X1 U11539 ( .A1(n13614), .A2(n13613), .ZN(n11142) );
  NOR2_X1 U11540 ( .A1(n13619), .A2(n13604), .ZN(n11141) );
  NOR2_X1 U11541 ( .A1(n20774), .A2(n15308), .ZN(n17467) );
  NOR2_X1 U11542 ( .A1(n15310), .A2(n20117), .ZN(n17456) );
  NAND2_X1 U11543 ( .A1(n17773), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11325) );
  INV_X1 U11544 ( .A(n18053), .ZN(n17772) );
  AOI21_X1 U11545 ( .B1(n16779), .B2(n21257), .A(n21250), .ZN(n16778) );
  INV_X1 U11546 ( .A(n20799), .ZN(n15387) );
  INV_X1 U11547 ( .A(n18883), .ZN(n15394) );
  AND2_X1 U11548 ( .A1(n13425), .A2(n13350), .ZN(n13351) );
  MUX2_X1 U11549 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13352) );
  AOI21_X1 U11550 ( .B1(n11758), .B2(n11370), .A(n11368), .ZN(n14506) );
  NOR2_X1 U11551 ( .A1(n11687), .A2(n11369), .ZN(n11368) );
  AND2_X1 U11552 ( .A1(n11683), .A2(n11075), .ZN(n11370) );
  INV_X1 U11553 ( .A(n11704), .ZN(n11369) );
  AND2_X1 U11554 ( .A1(n14315), .A2(n14314), .ZN(n14334) );
  INV_X1 U11555 ( .A(n21692), .ZN(n14314) );
  NOR2_X1 U11556 ( .A1(n11353), .A2(n11352), .ZN(n11351) );
  INV_X1 U11557 ( .A(n15151), .ZN(n11352) );
  NAND2_X1 U11558 ( .A1(n14407), .A2(n14825), .ZN(n14777) );
  NAND2_X1 U11559 ( .A1(n13255), .A2(n13254), .ZN(n14005) );
  AND2_X1 U11560 ( .A1(n13269), .A2(n12425), .ZN(n13094) );
  INV_X1 U11561 ( .A(n14018), .ZN(n12909) );
  AND4_X1 U11562 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n13036) );
  AND4_X1 U11563 ( .A1(n13021), .A2(n13020), .A3(n13019), .A4(n13018), .ZN(
        n13037) );
  AOI22_X1 U11564 ( .A1(n21225), .A2(n21223), .B1(n21229), .B2(n21087), .ZN(
        n21254) );
  OAI21_X1 U11565 ( .B1(n18114), .B2(n11126), .A(n11125), .ZN(n18104) );
  AOI21_X1 U11566 ( .B1(n17724), .B2(n20888), .A(n11127), .ZN(n11125) );
  INV_X1 U11567 ( .A(n18106), .ZN(n11127) );
  NAND2_X1 U11568 ( .A1(n11305), .A2(n11304), .ZN(n17954) );
  AND2_X1 U11569 ( .A1(n17931), .A2(n11306), .ZN(n11305) );
  NOR2_X1 U11570 ( .A1(n11307), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11306) );
  INV_X1 U11571 ( .A(n17930), .ZN(n11307) );
  NAND2_X1 U11572 ( .A1(n17932), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U11573 ( .A1(n17902), .A2(n17901), .ZN(n17909) );
  NAND2_X1 U11574 ( .A1(n14839), .A2(n18634), .ZN(n18647) );
  AOI21_X1 U11575 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21241), .A(
        n15401), .ZN(n15402) );
  AND2_X1 U11576 ( .A1(n11786), .A2(n11785), .ZN(n11808) );
  INV_X1 U11577 ( .A(n13483), .ZN(n11637) );
  NAND2_X1 U11578 ( .A1(n14445), .A2(n21683), .ZN(n11723) );
  NAND2_X1 U11579 ( .A1(n12241), .A2(n13521), .ZN(n12263) );
  AND2_X1 U11580 ( .A1(n13716), .A2(n13715), .ZN(n13723) );
  NAND2_X1 U11581 ( .A1(n12944), .A2(n11406), .ZN(n14377) );
  NAND2_X1 U11582 ( .A1(n11143), .A2(n12434), .ZN(n12452) );
  NAND2_X1 U11583 ( .A1(n13600), .A2(n15161), .ZN(n13626) );
  AND2_X1 U11584 ( .A1(n12870), .A2(n12869), .ZN(n12872) );
  AND2_X1 U11585 ( .A1(n12397), .A2(n12440), .ZN(n12395) );
  INV_X1 U11586 ( .A(n13326), .ZN(n12201) );
  NAND2_X1 U11587 ( .A1(n11041), .A2(n11068), .ZN(n11384) );
  AND2_X1 U11588 ( .A1(n11367), .A2(n15015), .ZN(n11366) );
  AND3_X1 U11589 ( .A1(n14227), .A2(n12273), .A3(n13582), .ZN(n14251) );
  AOI21_X1 U11590 ( .B1(n19950), .B2(n11334), .A(n13418), .ZN(n11333) );
  INV_X1 U11591 ( .A(n13564), .ZN(n11334) );
  INV_X1 U11592 ( .A(n15636), .ZN(n11252) );
  NOR2_X1 U11593 ( .A1(n15296), .A2(n11253), .ZN(n11257) );
  OR2_X1 U11594 ( .A1(n11254), .A2(n11255), .ZN(n11253) );
  INV_X1 U11595 ( .A(n15600), .ZN(n11254) );
  NAND2_X1 U11596 ( .A1(n13364), .A2(n14356), .ZN(n13436) );
  NAND2_X1 U11597 ( .A1(n13349), .A2(n13464), .ZN(n13425) );
  AOI21_X1 U11598 ( .B1(n21961), .B2(n21683), .A(n11680), .ZN(n11681) );
  INV_X1 U11599 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21922) );
  NOR2_X1 U11600 ( .A1(n11393), .A2(n11467), .ZN(n11473) );
  NAND2_X1 U11601 ( .A1(n12235), .A2(n12234), .ZN(n12239) );
  OR2_X1 U11602 ( .A1(n12263), .A2(n12239), .ZN(n12270) );
  NAND2_X1 U11603 ( .A1(n11662), .A2(n11661), .ZN(n12248) );
  NOR2_X1 U11604 ( .A1(n13862), .A2(n13860), .ZN(n13864) );
  AND2_X1 U11605 ( .A1(n13823), .A2(n13821), .ZN(n13806) );
  NOR2_X2 U11606 ( .A1(n13800), .A2(n13798), .ZN(n13823) );
  OR2_X1 U11607 ( .A1(n11362), .A2(n16155), .ZN(n11361) );
  NAND2_X1 U11608 ( .A1(n11363), .A2(n16159), .ZN(n11362) );
  INV_X1 U11609 ( .A(n16168), .ZN(n11363) );
  AND2_X1 U11610 ( .A1(n14881), .A2(n11248), .ZN(n11247) );
  INV_X1 U11611 ( .A(n14699), .ZN(n11248) );
  NOR2_X1 U11612 ( .A1(n17069), .A2(n11224), .ZN(n11223) );
  INV_X1 U11613 ( .A(n13148), .ZN(n11287) );
  AND4_X1 U11614 ( .A1(n13032), .A2(n13031), .A3(n13030), .A4(n13029), .ZN(
        n13035) );
  AND2_X1 U11615 ( .A1(n11206), .A2(n11204), .ZN(n11203) );
  INV_X1 U11616 ( .A(n14040), .ZN(n11204) );
  AND2_X1 U11617 ( .A1(n11275), .A2(n11274), .ZN(n11273) );
  INV_X1 U11618 ( .A(n16259), .ZN(n11274) );
  OR2_X1 U11619 ( .A1(n11280), .A2(n14484), .ZN(n11279) );
  INV_X1 U11620 ( .A(n14487), .ZN(n11280) );
  NAND2_X1 U11621 ( .A1(n11207), .A2(n11049), .ZN(n11206) );
  INV_X1 U11622 ( .A(n17072), .ZN(n11207) );
  AND2_X1 U11623 ( .A1(n13942), .A2(n11049), .ZN(n11208) );
  NAND2_X1 U11624 ( .A1(n11272), .A2(n15176), .ZN(n11271) );
  INV_X1 U11625 ( .A(n14952), .ZN(n11272) );
  OR2_X1 U11626 ( .A1(n12858), .A2(n12857), .ZN(n13919) );
  AND2_X1 U11627 ( .A1(n13669), .A2(n13640), .ZN(n11296) );
  OAI21_X1 U11628 ( .B1(n13089), .B2(n17170), .A(n12948), .ZN(n14378) );
  NAND2_X1 U11629 ( .A1(n12491), .A2(n12492), .ZN(n12506) );
  AND3_X1 U11630 ( .A1(n12304), .A2(n12303), .A3(n12373), .ZN(n12309) );
  AOI21_X1 U11631 ( .B1(n17409), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n11122), .ZN(n11121) );
  NOR2_X1 U11632 ( .A1(n15309), .A2(n20773), .ZN(n15306) );
  NOR2_X1 U11633 ( .A1(n17862), .A2(n11157), .ZN(n11156) );
  NOR2_X1 U11634 ( .A1(n18040), .A2(n11167), .ZN(n11166) );
  NOR2_X1 U11635 ( .A1(n20596), .A2(n17720), .ZN(n17692) );
  NOR2_X1 U11636 ( .A1(n21162), .A2(n17772), .ZN(n17774) );
  NAND2_X1 U11637 ( .A1(n11185), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17762) );
  NAND2_X1 U11638 ( .A1(n18136), .A2(n17752), .ZN(n17754) );
  AND2_X1 U11639 ( .A1(n17713), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11132) );
  INV_X1 U11640 ( .A(n17713), .ZN(n11131) );
  NOR2_X1 U11641 ( .A1(n17716), .A2(n17711), .ZN(n17712) );
  NAND2_X1 U11642 ( .A1(n15418), .A2(n20756), .ZN(n17730) );
  NOR2_X1 U11643 ( .A1(n15395), .A2(n15394), .ZN(n20755) );
  INV_X1 U11644 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21234) );
  NAND2_X1 U11645 ( .A1(n11114), .A2(n11113), .ZN(n11112) );
  OR2_X1 U11646 ( .A1(n21245), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11114) );
  INV_X1 U11647 ( .A(n21254), .ZN(n11105) );
  NAND2_X1 U11648 ( .A1(n21253), .A2(n21252), .ZN(n11104) );
  NAND2_X1 U11649 ( .A1(n11107), .A2(n21247), .ZN(n11106) );
  NAND2_X1 U11650 ( .A1(n11108), .A2(n21245), .ZN(n11107) );
  NAND2_X1 U11651 ( .A1(n11110), .A2(n11109), .ZN(n11108) );
  NOR2_X1 U11652 ( .A1(n15646), .A2(n15584), .ZN(n15637) );
  NAND2_X1 U11653 ( .A1(n11257), .A2(n11256), .ZN(n15646) );
  INV_X1 U11654 ( .A(n15643), .ZN(n11256) );
  AND2_X1 U11655 ( .A1(n13391), .A2(n13390), .ZN(n15267) );
  OR2_X1 U11656 ( .A1(n14323), .A2(n13464), .ZN(n11259) );
  NOR2_X1 U11657 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  INV_X1 U11658 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11959) );
  NOR2_X1 U11659 ( .A1(n11916), .A2(n15278), .ZN(n11930) );
  INV_X1 U11660 ( .A(n15028), .ZN(n11367) );
  CLKBUF_X1 U11661 ( .A(n15013), .Z(n15014) );
  INV_X1 U11662 ( .A(n15241), .ZN(n13547) );
  NAND2_X1 U11663 ( .A1(n13510), .A2(n13509), .ZN(n11341) );
  INV_X1 U11664 ( .A(n14505), .ZN(n11702) );
  OR2_X1 U11665 ( .A1(n14310), .A2(n21692), .ZN(n14271) );
  AND2_X1 U11666 ( .A1(n13568), .A2(n11043), .ZN(n11174) );
  AND2_X1 U11667 ( .A1(n15269), .A2(n15232), .ZN(n15253) );
  NOR2_X1 U11668 ( .A1(n13540), .A2(n13481), .ZN(n13541) );
  NAND2_X1 U11669 ( .A1(n21683), .A2(n14557), .ZN(n21871) );
  NAND2_X1 U11670 ( .A1(n14521), .A2(n14519), .ZN(n21894) );
  AND2_X1 U11671 ( .A1(n21961), .A2(n14547), .ZN(n21910) );
  INV_X1 U11672 ( .A(n11020), .ZN(n21865) );
  NOR2_X1 U11673 ( .A1(n21945), .A2(n21871), .ZN(n21998) );
  OR2_X1 U11674 ( .A1(n14519), .A2(n11724), .ZN(n21984) );
  INV_X1 U11675 ( .A(n21984), .ZN(n21989) );
  AND2_X1 U11676 ( .A1(n12894), .A2(n12895), .ZN(n14819) );
  NOR2_X1 U11677 ( .A1(n13869), .A2(n13868), .ZN(n13878) );
  OR2_X1 U11678 ( .A1(n13858), .A2(n13857), .ZN(n13869) );
  NAND2_X1 U11679 ( .A1(n13844), .A2(n11163), .ZN(n13855) );
  NOR2_X1 U11680 ( .A1(n13852), .A2(n11164), .ZN(n11163) );
  INV_X1 U11681 ( .A(n13286), .ZN(n11164) );
  INV_X1 U11682 ( .A(n18483), .ZN(n11217) );
  NAND2_X1 U11683 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11227) );
  NOR2_X2 U11684 ( .A1(n13810), .A2(n13809), .ZN(n13811) );
  OAI21_X1 U11685 ( .B1(n15465), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13997), 
        .ZN(n15113) );
  INV_X1 U11686 ( .A(n14822), .ZN(n13268) );
  AND2_X1 U11687 ( .A1(n14495), .A2(n11084), .ZN(n11358) );
  INV_X1 U11688 ( .A(n12735), .ZN(n11348) );
  NAND2_X1 U11689 ( .A1(n14835), .A2(n12441), .ZN(n12908) );
  NAND2_X1 U11690 ( .A1(n14079), .A2(n11070), .ZN(n16165) );
  INV_X1 U11691 ( .A(n16167), .ZN(n11236) );
  AND2_X1 U11692 ( .A1(n13180), .A2(n13179), .ZN(n14943) );
  XNOR2_X1 U11693 ( .A(n13944), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17072) );
  OR2_X1 U11694 ( .A1(n13939), .A2(n13596), .ZN(n13944) );
  OR2_X1 U11695 ( .A1(n13984), .A2(n16267), .ZN(n13985) );
  OR2_X1 U11696 ( .A1(n13255), .A2(n13254), .ZN(n13256) );
  NAND2_X1 U11697 ( .A1(n16197), .A2(n13084), .ZN(n16200) );
  NAND2_X1 U11698 ( .A1(n18540), .A2(n13276), .ZN(n16296) );
  INV_X1 U11699 ( .A(n16339), .ZN(n11290) );
  AND2_X1 U11700 ( .A1(n13827), .A2(n13826), .ZN(n13843) );
  NAND2_X1 U11701 ( .A1(n16351), .A2(n16350), .ZN(n16349) );
  AND2_X1 U11702 ( .A1(n16078), .A2(n15213), .ZN(n11275) );
  AND2_X1 U11703 ( .A1(n14936), .A2(n16078), .ZN(n16080) );
  AND3_X1 U11704 ( .A1(n13045), .A2(n13044), .A3(n13043), .ZN(n15036) );
  NOR2_X1 U11705 ( .A1(n11266), .A2(n11265), .ZN(n11264) );
  NOR2_X1 U11706 ( .A1(n13596), .A2(n13038), .ZN(n11265) );
  XNOR2_X1 U11707 ( .A(n14373), .B(n12505), .ZN(n14404) );
  NAND2_X1 U11708 ( .A1(n13959), .A2(n12893), .ZN(n15112) );
  OAI21_X1 U11709 ( .B1(n12524), .B2(n12523), .A(n12527), .ZN(n12525) );
  AND2_X1 U11710 ( .A1(n19255), .A2(n19254), .ZN(n19287) );
  AND2_X1 U11711 ( .A1(n19255), .A2(n17161), .ZN(n19242) );
  OR2_X1 U11712 ( .A1(n19625), .A2(n19307), .ZN(n19325) );
  NOR2_X1 U11713 ( .A1(n19255), .A2(n19254), .ZN(n19140) );
  OR2_X1 U11715 ( .A1(n13899), .A2(n12903), .ZN(n14833) );
  BUF_X1 U11716 ( .A(n12456), .Z(n14765) );
  OR2_X1 U11717 ( .A1(n20394), .A2(n11019), .ZN(n11153) );
  NAND2_X1 U11718 ( .A1(n20116), .A2(n20113), .ZN(n20118) );
  NAND2_X1 U11719 ( .A1(n20777), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11180) );
  AND2_X1 U11720 ( .A1(n17664), .A2(n17665), .ZN(n11312) );
  NOR2_X1 U11721 ( .A1(n11134), .A2(n11133), .ZN(n11311) );
  INV_X1 U11722 ( .A(n17666), .ZN(n11133) );
  NAND2_X1 U11723 ( .A1(n20799), .A2(n20615), .ZN(n20746) );
  NOR2_X2 U11724 ( .A1(n17882), .A2(n20429), .ZN(n17892) );
  INV_X1 U11725 ( .A(n20925), .ZN(n18039) );
  INV_X1 U11726 ( .A(n17723), .ZN(n17721) );
  NAND2_X1 U11727 ( .A1(n18114), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18113) );
  NAND2_X1 U11728 ( .A1(n17692), .A2(n17738), .ZN(n21090) );
  NAND2_X1 U11729 ( .A1(n21089), .A2(n21088), .ZN(n21094) );
  NAND2_X1 U11730 ( .A1(n20978), .A2(n11191), .ZN(n21013) );
  INV_X1 U11731 ( .A(n21051), .ZN(n11191) );
  NAND2_X1 U11732 ( .A1(n11308), .A2(n11309), .ZN(n17932) );
  NAND2_X1 U11733 ( .A1(n11309), .A2(n18051), .ZN(n17931) );
  OAI21_X1 U11734 ( .B1(n17827), .B2(n11087), .A(n18051), .ZN(n11326) );
  NAND2_X1 U11735 ( .A1(n11325), .A2(n11320), .ZN(n18012) );
  INV_X1 U11736 ( .A(n11322), .ZN(n11321) );
  AOI21_X1 U11737 ( .B1(n18051), .B2(n11087), .A(n11323), .ZN(n11322) );
  NAND2_X1 U11738 ( .A1(n17976), .A2(n21177), .ZN(n11324) );
  INV_X1 U11739 ( .A(n11325), .ZN(n11319) );
  AOI22_X1 U11740 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U11741 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15376) );
  AOI211_X1 U11742 ( .C1(n10991), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n15373), .B(n15372), .ZN(n15374) );
  AND2_X1 U11743 ( .A1(n11033), .A2(n11124), .ZN(n21227) );
  INV_X1 U11744 ( .A(n16778), .ZN(n11124) );
  NOR2_X1 U11745 ( .A1(n21230), .A2(n21086), .ZN(n21153) );
  NAND2_X1 U11746 ( .A1(n18090), .A2(n17729), .ZN(n18077) );
  NAND2_X1 U11747 ( .A1(n17759), .A2(n18107), .ZN(n18097) );
  OR2_X1 U11748 ( .A1(n18097), .A2(n18098), .ZN(n11185) );
  NAND2_X1 U11749 ( .A1(n18091), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18090) );
  INV_X1 U11750 ( .A(n20726), .ZN(n17694) );
  XNOR2_X1 U11751 ( .A(n20726), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18159) );
  NAND2_X1 U11752 ( .A1(n11093), .A2(n11092), .ZN(n15390) );
  NAND2_X1 U11753 ( .A1(n15392), .A2(n15394), .ZN(n11092) );
  INV_X1 U11754 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U11755 ( .A1(n14111), .A2(n14212), .ZN(n21286) );
  OR2_X1 U11756 ( .A1(n11659), .A2(n11658), .ZN(n11660) );
  XNOR2_X1 U11757 ( .A(n13442), .B(n13441), .ZN(n15879) );
  AND2_X2 U11758 ( .A1(n13467), .A2(n14314), .ZN(n19911) );
  NAND2_X1 U11759 ( .A1(n14257), .A2(n13466), .ZN(n13467) );
  OR2_X1 U11760 ( .A1(n13465), .A2(n13464), .ZN(n13466) );
  NOR2_X1 U11761 ( .A1(n14050), .A2(n11381), .ZN(n14051) );
  INV_X1 U11762 ( .A(n11013), .ZN(n14050) );
  AND2_X1 U11763 ( .A1(n12281), .A2(n14314), .ZN(n15260) );
  OR2_X1 U11764 ( .A1(n14260), .A2(n12280), .ZN(n12281) );
  OR2_X1 U11765 ( .A1(n12207), .A2(n12208), .ZN(n12209) );
  OR2_X1 U11766 ( .A1(n16817), .A2(n14271), .ZN(n21667) );
  XNOR2_X1 U11767 ( .A(n13469), .B(n11245), .ZN(n15906) );
  INV_X1 U11768 ( .A(n13470), .ZN(n11245) );
  NAND2_X1 U11769 ( .A1(n14334), .A2(n14324), .ZN(n21429) );
  INV_X1 U11770 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21975) );
  NAND2_X1 U11771 ( .A1(n16060), .A2(n18584), .ZN(n18482) );
  NAND2_X1 U11772 ( .A1(n16061), .A2(n16377), .ZN(n16060) );
  NAND2_X1 U11773 ( .A1(n15113), .A2(n18423), .ZN(n16077) );
  INV_X1 U11774 ( .A(n18562), .ZN(n18580) );
  NAND2_X1 U11775 ( .A1(n17055), .A2(n14850), .ZN(n18562) );
  INV_X1 U11776 ( .A(n14905), .ZN(n12571) );
  OR2_X1 U11777 ( .A1(n12581), .A2(n12580), .ZN(n14941) );
  INV_X1 U11778 ( .A(n16178), .ZN(n16169) );
  INV_X1 U11779 ( .A(n17144), .ZN(n17043) );
  XNOR2_X1 U11780 ( .A(n11213), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15470) );
  NAND2_X1 U11781 ( .A1(n15504), .A2(n17133), .ZN(n13952) );
  INV_X1 U11782 ( .A(n17119), .ZN(n17131) );
  AND2_X1 U11783 ( .A1(n17117), .A2(n17127), .ZN(n17105) );
  INV_X1 U11784 ( .A(n17105), .ZN(n17125) );
  NAND2_X1 U11785 ( .A1(n18647), .A2(n13949), .ZN(n17117) );
  NAND2_X1 U11786 ( .A1(n15470), .A2(n18612), .ZN(n14044) );
  INV_X1 U11787 ( .A(n11213), .ZN(n14032) );
  XNOR2_X1 U11788 ( .A(n13885), .B(n13884), .ZN(n15464) );
  OAI211_X1 U11789 ( .C1(n18564), .C2(n16705), .A(n11263), .B(n11262), .ZN(
        n11261) );
  INV_X1 U11790 ( .A(n16441), .ZN(n11262) );
  INV_X1 U11791 ( .A(n19321), .ZN(n19307) );
  INV_X1 U11792 ( .A(n16761), .ZN(n18637) );
  NOR2_X1 U11793 ( .A1(n19153), .A2(n19160), .ZN(n19727) );
  NOR2_X1 U11794 ( .A1(n21227), .A2(n20062), .ZN(n20116) );
  NAND2_X1 U11795 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21274), .ZN(n21279) );
  INV_X1 U11796 ( .A(n20523), .ZN(n20479) );
  NOR2_X2 U11797 ( .A1(n20340), .A2(n21264), .ZN(n20523) );
  INV_X1 U11798 ( .A(n20522), .ZN(n20544) );
  INV_X1 U11799 ( .A(n11189), .ZN(n11188) );
  AOI21_X1 U11800 ( .B1(n21066), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11189) );
  INV_X1 U11801 ( .A(n21213), .ZN(n21188) );
  INV_X1 U11802 ( .A(n21186), .ZN(n21113) );
  AND4_X1 U11803 ( .A1(n13737), .A2(n13736), .A3(n13735), .A4(n13734), .ZN(
        n13745) );
  AND4_X1 U11804 ( .A1(n13703), .A2(n13702), .A3(n13701), .A4(n13700), .ZN(
        n13711) );
  NAND2_X1 U11805 ( .A1(n19309), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13625) );
  NAND2_X1 U11806 ( .A1(n12422), .A2(n13269), .ZN(n13964) );
  AOI22_X1 U11807 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U11808 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10981), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12389) );
  INV_X1 U11809 ( .A(n13556), .ZN(n11345) );
  OR2_X1 U11810 ( .A1(n11771), .A2(n11770), .ZN(n13523) );
  OR2_X1 U11811 ( .A1(n11784), .A2(n11783), .ZN(n13532) );
  OR2_X1 U11812 ( .A1(n11721), .A2(n11720), .ZN(n13503) );
  NAND2_X1 U11813 ( .A1(n11573), .A2(n15446), .ZN(n11577) );
  AOI22_X1 U11814 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U11815 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11447) );
  INV_X1 U11816 ( .A(n12258), .ZN(n12241) );
  INV_X1 U11817 ( .A(n12240), .ZN(n12264) );
  AOI21_X1 U11818 ( .B1(n19178), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n19574), .ZN(n13643) );
  AOI21_X1 U11819 ( .B1(n13668), .B2(n13268), .A(n13267), .ZN(n13893) );
  NAND2_X1 U11820 ( .A1(n12466), .A2(n12467), .ZN(n12469) );
  NAND2_X1 U11821 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U11822 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12311) );
  NAND2_X1 U11823 ( .A1(n12532), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12310) );
  XNOR2_X1 U11824 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12869) );
  AND2_X1 U11825 ( .A1(n13963), .A2(n12425), .ZN(n12367) );
  AOI21_X1 U11826 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21234), .A(
        n15400), .ZN(n15406) );
  NOR2_X1 U11827 ( .A1(n17369), .A2(n18841), .ZN(n11122) );
  NAND2_X1 U11828 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21232), .ZN(
        n15307) );
  NOR2_X1 U11829 ( .A1(n20117), .A2(n15307), .ZN(n17661) );
  NOR2_X1 U11830 ( .A1(n20605), .A2(n17710), .ZN(n17693) );
  NAND2_X1 U11831 ( .A1(n11113), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11110) );
  INV_X1 U11832 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11109) );
  INV_X1 U11833 ( .A(n15196), .ZN(n11385) );
  NAND2_X1 U11834 ( .A1(n12208), .A2(n11381), .ZN(n11380) );
  AND2_X1 U11835 ( .A1(n11374), .A2(n11373), .ZN(n11372) );
  INV_X1 U11836 ( .A(n15634), .ZN(n11373) );
  NOR2_X1 U11837 ( .A1(n15583), .A2(n11375), .ZN(n11374) );
  INV_X1 U11838 ( .A(n15647), .ZN(n11375) );
  NAND2_X1 U11839 ( .A1(n11930), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11960) );
  AND3_X1 U11840 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n11799), .ZN(n11789) );
  NOR2_X1 U11841 ( .A1(n14578), .A2(n22008), .ZN(n11788) );
  NOR2_X1 U11842 ( .A1(n15530), .A2(n11241), .ZN(n11240) );
  INV_X1 U11843 ( .A(n15544), .ZN(n11241) );
  OR2_X1 U11844 ( .A1(n11258), .A2(n15297), .ZN(n11255) );
  OR2_X1 U11845 ( .A1(n11745), .A2(n11744), .ZN(n13511) );
  NOR2_X1 U11846 ( .A1(n11662), .A2(n11641), .ZN(n13539) );
  NAND2_X1 U11847 ( .A1(n11519), .A2(n14578), .ZN(n11097) );
  NAND2_X1 U11848 ( .A1(n13486), .A2(n11522), .ZN(n11518) );
  AOI22_X1 U11849 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U11850 ( .B1(n21687), .B2(n14474), .A(n21671), .ZN(n14557) );
  INV_X1 U11851 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21965) );
  MUX2_X1 U11852 ( .A(n12437), .B(n12428), .S(n12440), .Z(n12438) );
  AND2_X1 U11853 ( .A1(n16052), .A2(n16227), .ZN(n11285) );
  OR2_X1 U11854 ( .A1(n13816), .A2(n13814), .ZN(n13810) );
  NAND2_X1 U11855 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U11856 ( .A1(n13806), .A2(n13804), .ZN(n13816) );
  NOR2_X1 U11857 ( .A1(n11155), .A2(n13763), .ZN(n11154) );
  INV_X1 U11858 ( .A(n13717), .ZN(n11162) );
  NAND2_X1 U11859 ( .A1(n11072), .A2(n13673), .ZN(n13718) );
  OAI21_X1 U11860 ( .B1(n13228), .B2(n14411), .A(n11402), .ZN(n12449) );
  NAND2_X1 U11861 ( .A1(n12735), .A2(n16139), .ZN(n11349) );
  NAND3_X1 U11862 ( .A1(n19353), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n18291), 
        .ZN(n12750) );
  NAND2_X1 U11863 ( .A1(n11234), .A2(n16111), .ZN(n11233) );
  INV_X1 U11864 ( .A(n16126), .ZN(n11234) );
  NOR2_X1 U11865 ( .A1(n18382), .A2(n11226), .ZN(n11225) );
  NAND2_X1 U11866 ( .A1(n11223), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11221) );
  INV_X1 U11867 ( .A(n12517), .ZN(n11289) );
  NOR2_X1 U11868 ( .A1(n11200), .A2(n13150), .ZN(n11199) );
  INV_X1 U11869 ( .A(n12481), .ZN(n12482) );
  NAND2_X1 U11870 ( .A1(n12516), .A2(n13148), .ZN(n12485) );
  OR2_X1 U11871 ( .A1(n12940), .A2(n12939), .ZN(n13906) );
  AND2_X1 U11872 ( .A1(n16327), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11302) );
  NOR2_X1 U11873 ( .A1(n13867), .A2(n16307), .ZN(n13870) );
  NOR2_X1 U11874 ( .A1(n18547), .A2(n13596), .ZN(n13872) );
  NOR2_X1 U11875 ( .A1(n16489), .A2(n14026), .ZN(n11212) );
  AND2_X1 U11876 ( .A1(n11285), .A2(n16218), .ZN(n11284) );
  AND2_X1 U11877 ( .A1(n16237), .A2(n11282), .ZN(n16197) );
  AND2_X1 U11878 ( .A1(n11284), .A2(n11283), .ZN(n11282) );
  INV_X1 U11879 ( .A(n16207), .ZN(n11283) );
  AND2_X1 U11880 ( .A1(n13839), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13840) );
  INV_X1 U11881 ( .A(n16172), .ZN(n11237) );
  OR2_X1 U11882 ( .A1(n13014), .A2(n13013), .ZN(n13748) );
  OR2_X1 U11883 ( .A1(n13002), .A2(n13001), .ZN(n13275) );
  OR2_X1 U11884 ( .A1(n12868), .A2(n12867), .ZN(n13638) );
  AND2_X1 U11885 ( .A1(n12456), .A2(n12398), .ZN(n14006) );
  OAI21_X1 U11886 ( .B1(n12456), .B2(n19628), .A(n13249), .ZN(n12904) );
  INV_X1 U11887 ( .A(n13906), .ZN(n16746) );
  NAND2_X1 U11888 ( .A1(n12488), .A2(n19293), .ZN(n12521) );
  NOR2_X1 U11889 ( .A1(n12750), .A2(n13651), .ZN(n12505) );
  MUX2_X1 U11890 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12892), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13959) );
  AND2_X1 U11891 ( .A1(n17142), .A2(n18295), .ZN(n17045) );
  AND3_X1 U11893 ( .A1(n12331), .A2(n12373), .A3(n12330), .ZN(n12335) );
  AOI22_X1 U11894 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12358) );
  AOI221_X1 U11895 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12890), 
        .C1(n16769), .C2(n12890), .A(n12889), .ZN(n13899) );
  NOR2_X1 U11896 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16788), .ZN(
        n12889) );
  AND2_X1 U11897 ( .A1(n18286), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12502) );
  NOR2_X1 U11898 ( .A1(n15392), .A2(n17733), .ZN(n15418) );
  NAND2_X1 U11899 ( .A1(n20772), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15308) );
  NAND2_X1 U11900 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21240), .ZN(
        n15310) );
  OR2_X1 U11901 ( .A1(n20774), .A2(n20117), .ZN(n17369) );
  OR2_X1 U11902 ( .A1(n20773), .A2(n15308), .ZN(n11387) );
  NOR2_X1 U11903 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20764), .ZN(
        n15348) );
  INV_X1 U11904 ( .A(n11182), .ZN(n11181) );
  OAI21_X1 U11905 ( .B1(n17369), .B2(n11184), .A(n11183), .ZN(n11182) );
  INV_X1 U11906 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U11907 ( .A1(n15306), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11183) );
  AOI21_X1 U11908 ( .B1(n15360), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n11136), .ZN(n11135) );
  NOR2_X1 U11909 ( .A1(n15367), .A2(n11137), .ZN(n11136) );
  INV_X1 U11910 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U11911 ( .A1(n17954), .A2(n18051), .B1(n11139), .B2(n17933), .ZN(
        n17934) );
  INV_X1 U11912 ( .A(n17932), .ZN(n11139) );
  NAND2_X1 U11913 ( .A1(n11324), .A2(n21170), .ZN(n11323) );
  NOR2_X1 U11914 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11328) );
  INV_X1 U11915 ( .A(n18078), .ZN(n11317) );
  NOR2_X1 U11916 ( .A1(n17976), .A2(n18077), .ZN(n18045) );
  NAND2_X1 U11917 ( .A1(n18118), .A2(n17756), .ZN(n17757) );
  NAND2_X1 U11918 ( .A1(n17726), .A2(n18104), .ZN(n17792) );
  INV_X1 U11919 ( .A(n20807), .ZN(n15395) );
  NOR2_X1 U11920 ( .A1(n15395), .A2(n17239), .ZN(n15426) );
  NOR2_X1 U11921 ( .A1(n20554), .A2(n16780), .ZN(n15425) );
  NOR2_X1 U11922 ( .A1(n20810), .A2(n15387), .ZN(n20756) );
  INV_X1 U11923 ( .A(n15306), .ZN(n15367) );
  INV_X1 U11924 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15603) );
  AND2_X1 U11925 ( .A1(n11942), .A2(n11883), .ZN(n15220) );
  NAND2_X1 U11926 ( .A1(n11657), .A2(n11656), .ZN(n11658) );
  OR2_X1 U11927 ( .A1(n11651), .A2(n11015), .ZN(n11657) );
  INV_X1 U11928 ( .A(n15559), .ZN(n21553) );
  AND2_X1 U11929 ( .A1(n13438), .A2(n13437), .ZN(n15518) );
  AND3_X1 U11930 ( .A1(n13414), .A2(n13425), .A3(n13413), .ZN(n15643) );
  NOR2_X1 U11931 ( .A1(n19907), .A2(n13374), .ZN(n19899) );
  OR2_X1 U11932 ( .A1(n14329), .A2(n14305), .ZN(n14257) );
  AND2_X1 U11933 ( .A1(n15260), .A2(n12293), .ZN(n15722) );
  AND2_X1 U11934 ( .A1(n14273), .A2(n14272), .ZN(n19801) );
  NOR2_X1 U11935 ( .A1(n14271), .A2(n21726), .ZN(n14272) );
  AND2_X1 U11936 ( .A1(n22008), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13329) );
  AND2_X1 U11937 ( .A1(n13304), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13343) );
  NOR2_X1 U11938 ( .A1(n11013), .A2(n11377), .ZN(n13461) );
  NAND2_X1 U11939 ( .A1(n11379), .A2(n11378), .ZN(n11377) );
  INV_X1 U11940 ( .A(n11380), .ZN(n11379) );
  INV_X1 U11941 ( .A(n13463), .ZN(n11378) );
  NOR2_X1 U11942 ( .A1(n12143), .A2(n15788), .ZN(n12144) );
  NAND2_X1 U11943 ( .A1(n12093), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12143) );
  AND2_X1 U11944 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12092), .ZN(
        n12093) );
  INV_X1 U11945 ( .A(n12091), .ZN(n12092) );
  NOR2_X1 U11946 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  AND2_X1 U11947 ( .A1(n12011), .A2(n12010), .ZN(n15592) );
  NOR2_X1 U11948 ( .A1(n11979), .A2(n15612), .ZN(n11980) );
  NAND2_X1 U11949 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12012) );
  CLKBUF_X1 U11950 ( .A(n15593), .Z(n15594) );
  AND2_X1 U11951 ( .A1(n11978), .A2(n11977), .ZN(n15292) );
  AND2_X1 U11952 ( .A1(n11963), .A2(n11962), .ZN(n15288) );
  NAND2_X1 U11953 ( .A1(n11383), .A2(n15227), .ZN(n11382) );
  INV_X1 U11954 ( .A(n11384), .ZN(n11383) );
  INV_X1 U11955 ( .A(n11911), .ZN(n11894) );
  NOR2_X1 U11956 ( .A1(n11867), .A2(n11866), .ZN(n11868) );
  NAND2_X1 U11957 ( .A1(n11868), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U11958 ( .A1(n11848), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11867) );
  NOR2_X1 U11959 ( .A1(n11833), .A2(n15245), .ZN(n11848) );
  NAND2_X1 U11960 ( .A1(n11814), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11833) );
  AND2_X1 U11961 ( .A1(n11789), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U11962 ( .A1(n14503), .A2(n11704), .ZN(n14531) );
  NOR2_X1 U11963 ( .A1(n15742), .A2(n11337), .ZN(n11336) );
  INV_X1 U11964 ( .A(n11339), .ZN(n11337) );
  AND2_X1 U11965 ( .A1(n15557), .A2(n11238), .ZN(n15519) );
  NOR2_X1 U11966 ( .A1(n11239), .A2(n15518), .ZN(n11238) );
  INV_X1 U11967 ( .A(n11240), .ZN(n11239) );
  NAND2_X1 U11968 ( .A1(n19950), .A2(n11340), .ZN(n11339) );
  INV_X1 U11969 ( .A(n15909), .ZN(n11340) );
  NAND2_X1 U11970 ( .A1(n15557), .A2(n11240), .ZN(n15531) );
  NAND2_X1 U11971 ( .A1(n15557), .A2(n15544), .ZN(n15546) );
  AOI21_X1 U11972 ( .B1(n11333), .B2(n10972), .A(n10972), .ZN(n11330) );
  NOR2_X1 U11973 ( .A1(n11251), .A2(n15628), .ZN(n11249) );
  OAI21_X1 U11974 ( .B1(n15809), .B2(n10972), .A(n11333), .ZN(n13567) );
  NAND2_X1 U11975 ( .A1(n15637), .A2(n15636), .ZN(n15635) );
  NAND2_X1 U11976 ( .A1(n15637), .A2(n11250), .ZN(n15629) );
  AND2_X1 U11977 ( .A1(n13412), .A2(n13411), .ZN(n15600) );
  NOR2_X1 U11978 ( .A1(n15296), .A2(n11255), .ZN(n15656) );
  INV_X1 U11979 ( .A(n11257), .ZN(n15644) );
  NOR2_X1 U11980 ( .A1(n15296), .A2(n15297), .ZN(n15654) );
  AND3_X1 U11981 ( .A1(n13403), .A2(n13425), .A3(n13402), .ZN(n15285) );
  OR2_X1 U11982 ( .A1(n15286), .A2(n15285), .ZN(n15296) );
  AND2_X1 U11983 ( .A1(n13401), .A2(n13400), .ZN(n15252) );
  NAND2_X1 U11984 ( .A1(n15253), .A2(n15252), .ZN(n15286) );
  NAND2_X1 U11985 ( .A1(n15869), .A2(n11347), .ZN(n15847) );
  NOR2_X1 U11986 ( .A1(n19891), .A2(n13395), .ZN(n15269) );
  NAND2_X1 U11987 ( .A1(n11230), .A2(n11229), .ZN(n19891) );
  NOR2_X1 U11988 ( .A1(n15199), .A2(n19894), .ZN(n11229) );
  INV_X1 U11989 ( .A(n19893), .ZN(n11230) );
  OR2_X1 U11990 ( .A1(n13548), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13549) );
  OR2_X1 U11991 ( .A1(n19905), .A2(n19904), .ZN(n19907) );
  NAND2_X1 U11992 ( .A1(n11260), .A2(n13358), .ZN(n14533) );
  INV_X1 U11993 ( .A(n14508), .ZN(n11260) );
  NOR2_X1 U11994 ( .A1(n14533), .A2(n14532), .ZN(n14706) );
  NOR2_X1 U11995 ( .A1(n15881), .A2(n15880), .ZN(n21348) );
  AND2_X1 U11996 ( .A1(n21297), .A2(n21296), .ZN(n21349) );
  NAND2_X1 U11997 ( .A1(n14334), .A2(n14330), .ZN(n21334) );
  AND2_X1 U11998 ( .A1(n13354), .A2(n13353), .ZN(n14323) );
  NAND2_X1 U11999 ( .A1(n15446), .A2(n13360), .ZN(n14321) );
  NAND2_X1 U12000 ( .A1(n14334), .A2(n14455), .ZN(n21296) );
  AND2_X2 U12001 ( .A1(n13348), .A2(n11553), .ZN(n14356) );
  NAND2_X1 U12002 ( .A1(n11640), .A2(n11639), .ZN(n11695) );
  OR2_X1 U12003 ( .A1(n12258), .A2(n11634), .ZN(n11640) );
  INV_X1 U12004 ( .A(n11615), .ZN(n11616) );
  AOI21_X1 U12005 ( .B1(n11696), .B2(n11695), .A(n13539), .ZN(n11689) );
  INV_X1 U12006 ( .A(n11681), .ZN(n11098) );
  OR2_X1 U12007 ( .A1(n11651), .A2(n11335), .ZN(n11709) );
  INV_X1 U12008 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14281) );
  AND2_X1 U12009 ( .A1(n14564), .A2(n14578), .ZN(n11476) );
  INV_X1 U12010 ( .A(n11558), .ZN(n16033) );
  NOR2_X1 U12011 ( .A1(n11571), .A2(n11551), .ZN(n14449) );
  AND2_X1 U12012 ( .A1(n12210), .A2(n14717), .ZN(n14455) );
  NAND2_X1 U12013 ( .A1(n11659), .A2(n11658), .ZN(n14295) );
  OR2_X1 U12014 ( .A1(n21894), .A2(n21920), .ZN(n21876) );
  INV_X1 U12015 ( .A(n11574), .ZN(n14570) );
  NAND2_X1 U12016 ( .A1(n12248), .A2(n12237), .ZN(n12272) );
  INV_X1 U12017 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21722) );
  XNOR2_X1 U12018 ( .A(n13869), .B(n13868), .ZN(n18547) );
  OR2_X1 U12019 ( .A1(n13855), .A2(n13594), .ZN(n13862) );
  NOR2_X1 U12020 ( .A1(n13118), .A2(n16398), .ZN(n13119) );
  NOR2_X1 U12021 ( .A1(n13791), .A2(n11170), .ZN(n11169) );
  NAND2_X1 U12022 ( .A1(n13796), .A2(n13795), .ZN(n13793) );
  NOR2_X1 U12023 ( .A1(n11356), .A2(n13049), .ZN(n11355) );
  INV_X1 U12024 ( .A(n15049), .ZN(n11356) );
  XNOR2_X1 U12025 ( .A(n12789), .B(n11401), .ZN(n16119) );
  XNOR2_X1 U12026 ( .A(n16131), .B(n12770), .ZN(n16124) );
  NAND2_X1 U12027 ( .A1(n16124), .A2(n16123), .ZN(n16122) );
  NAND2_X1 U12028 ( .A1(n12734), .A2(n19574), .ZN(n12735) );
  OR2_X1 U12029 ( .A1(n11361), .A2(n11360), .ZN(n11359) );
  INV_X1 U12030 ( .A(n16150), .ZN(n11360) );
  CLKBUF_X1 U12031 ( .A(n15210), .Z(n15211) );
  AND3_X1 U12032 ( .A1(n13052), .A2(n13051), .A3(n13050), .ZN(n16641) );
  NAND2_X1 U12033 ( .A1(n11278), .A2(n14596), .ZN(n11277) );
  AND2_X1 U12034 ( .A1(n14147), .A2(n18292), .ZN(n17180) );
  INV_X1 U12035 ( .A(n14182), .ZN(n17039) );
  XNOR2_X1 U12036 ( .A(n13101), .B(n13100), .ZN(n15465) );
  INV_X1 U12037 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U12038 ( .A1(n13125), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13131) );
  AND2_X1 U12039 ( .A1(n16049), .A2(n16151), .ZN(n13219) );
  NAND2_X1 U12040 ( .A1(n13123), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13127) );
  NOR2_X2 U12041 ( .A1(n16165), .A2(n16160), .ZN(n16161) );
  NOR2_X1 U12042 ( .A1(n13115), .A2(n16084), .ZN(n13117) );
  NAND2_X1 U12043 ( .A1(n13117), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13118) );
  NAND2_X1 U12044 ( .A1(n13112), .A2(n11034), .ZN(n13113) );
  AND2_X1 U12045 ( .A1(n13112), .A2(n11225), .ZN(n13114) );
  NAND2_X1 U12046 ( .A1(n14539), .A2(n11048), .ZN(n14942) );
  NOR2_X1 U12047 ( .A1(n13110), .A2(n17094), .ZN(n13112) );
  NAND2_X1 U12048 ( .A1(n11220), .A2(n11218), .ZN(n13110) );
  INV_X1 U12049 ( .A(n11221), .ZN(n11220) );
  NOR2_X1 U12050 ( .A1(n13105), .A2(n11219), .ZN(n11218) );
  INV_X1 U12051 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11219) );
  NOR2_X1 U12052 ( .A1(n11221), .A2(n13105), .ZN(n13111) );
  INV_X1 U12053 ( .A(n16430), .ZN(n11145) );
  INV_X1 U12054 ( .A(n18620), .ZN(n13261) );
  INV_X1 U12055 ( .A(n13105), .ZN(n11222) );
  NOR2_X2 U12056 ( .A1(n14501), .A2(n14490), .ZN(n14614) );
  NOR2_X1 U12057 ( .A1(n11210), .A2(n14043), .ZN(n11209) );
  INV_X1 U12058 ( .A(n11212), .ZN(n11210) );
  NOR2_X1 U12059 ( .A1(n16269), .A2(n16268), .ZN(n13987) );
  NAND2_X1 U12060 ( .A1(n16296), .A2(n16438), .ZN(n16288) );
  INV_X1 U12061 ( .A(n16197), .ZN(n16209) );
  NOR2_X1 U12062 ( .A1(n16331), .A2(n16489), .ZN(n16319) );
  AND2_X1 U12063 ( .A1(n16237), .A2(n16052), .ZN(n16228) );
  AND2_X2 U12064 ( .A1(n16064), .A2(n16236), .ZN(n16237) );
  AND2_X1 U12065 ( .A1(n11203), .A2(n11089), .ZN(n11202) );
  NAND2_X1 U12066 ( .A1(n14079), .A2(n11066), .ZN(n16174) );
  AND2_X1 U12067 ( .A1(n13193), .A2(n13192), .ZN(n15152) );
  AND3_X1 U12068 ( .A1(n13059), .A2(n13058), .A3(n13057), .ZN(n18416) );
  AND2_X1 U12069 ( .A1(n18401), .A2(n13832), .ZN(n16420) );
  AND2_X1 U12070 ( .A1(n11301), .A2(n13784), .ZN(n11300) );
  NAND2_X1 U12071 ( .A1(n13777), .A2(n13778), .ZN(n11301) );
  INV_X1 U12072 ( .A(n14943), .ZN(n11246) );
  OR2_X1 U12073 ( .A1(n16686), .A2(n13775), .ZN(n16673) );
  INV_X1 U12074 ( .A(n14483), .ZN(n11276) );
  OR2_X1 U12075 ( .A1(n14483), .A2(n11279), .ZN(n15035) );
  CLKBUF_X1 U12076 ( .A(n13995), .Z(n13996) );
  NOR2_X1 U12077 ( .A1(n14483), .A2(n14484), .ZN(n14486) );
  AND2_X1 U12078 ( .A1(n13017), .A2(n13016), .ZN(n14482) );
  NAND2_X1 U12079 ( .A1(n13934), .A2(n13933), .ZN(n16714) );
  NAND2_X1 U12080 ( .A1(n13929), .A2(n13935), .ZN(n13934) );
  AOI21_X1 U12081 ( .B1(n13932), .B2(n13928), .A(n11396), .ZN(n13933) );
  OR2_X1 U12082 ( .A1(n14861), .A2(n11271), .ZN(n15175) );
  AND3_X1 U12083 ( .A1(n12992), .A2(n12991), .A3(n12990), .ZN(n14952) );
  NAND2_X1 U12084 ( .A1(n11298), .A2(n13640), .ZN(n13671) );
  INV_X1 U12085 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U12086 ( .A1(n14036), .A2(n14819), .ZN(n16586) );
  CLKBUF_X1 U12087 ( .A(n12904), .Z(n12905) );
  XNOR2_X1 U12088 ( .A(n12949), .B(n14376), .ZN(n14437) );
  AND2_X1 U12089 ( .A1(n14021), .A2(n14020), .ZN(n14785) );
  INV_X1 U12090 ( .A(n19160), .ZN(n19256) );
  AND2_X1 U12091 ( .A1(n19152), .A2(n17043), .ZN(n19286) );
  OR2_X1 U12092 ( .A1(n19152), .A2(n17043), .ZN(n19282) );
  INV_X1 U12093 ( .A(n19140), .ZN(n19153) );
  NAND2_X1 U12094 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19313), .ZN(n19627) );
  AOI21_X1 U12095 ( .B1(n21765), .B2(n21762), .A(n18269), .ZN(n20801) );
  OR2_X1 U12096 ( .A1(n20505), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n20518) );
  AOI21_X1 U12097 ( .B1(n20452), .B2(n20451), .A(n20528), .ZN(n20467) );
  NOR2_X1 U12098 ( .A1(n20467), .A2(n20468), .ZN(n20476) );
  OR2_X1 U12099 ( .A1(n20452), .A2(n20528), .ZN(n11168) );
  NOR2_X1 U12100 ( .A1(n20407), .A2(n20528), .ZN(n20408) );
  NOR2_X1 U12101 ( .A1(n20385), .A2(n20386), .ZN(n20394) );
  INV_X1 U12102 ( .A(n20428), .ZN(n20438) );
  AND2_X1 U12103 ( .A1(n18103), .A2(n11166), .ZN(n18041) );
  OAI21_X1 U12104 ( .B1(n17241), .B2(n17240), .A(n21272), .ZN(n20551) );
  NAND2_X1 U12105 ( .A1(n11119), .A2(n15354), .ZN(n20615) );
  NOR2_X1 U12106 ( .A1(n15353), .A2(n11120), .ZN(n11119) );
  NOR2_X1 U12107 ( .A1(n20062), .A2(n16777), .ZN(n18217) );
  NOR2_X1 U12108 ( .A1(n21257), .A2(n20062), .ZN(n20063) );
  NOR2_X1 U12109 ( .A1(n17968), .A2(n20130), .ZN(n18003) );
  NOR2_X1 U12110 ( .A1(n17952), .A2(n20473), .ZN(n17939) );
  INV_X1 U12111 ( .A(n21013), .ZN(n17989) );
  NAND3_X1 U12112 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17952) );
  NAND2_X1 U12113 ( .A1(n17782), .A2(n11040), .ZN(n17882) );
  NAND2_X1 U12114 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17863) );
  INV_X1 U12115 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17862) );
  NOR2_X1 U12116 ( .A1(n17767), .A2(n17766), .ZN(n17782) );
  INV_X1 U12117 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17766) );
  OAI21_X1 U12118 ( .B1(n20130), .B2(n17967), .A(n18751), .ZN(n17923) );
  NAND2_X1 U12119 ( .A1(n18027), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17790) );
  NOR2_X1 U12120 ( .A1(n18039), .A2(n20947), .ZN(n18025) );
  NOR2_X1 U12121 ( .A1(n17811), .A2(n17833), .ZN(n18027) );
  INV_X1 U12122 ( .A(n17923), .ZN(n17966) );
  NAND2_X1 U12123 ( .A1(n18103), .A2(n11165), .ZN(n17811) );
  AND2_X1 U12124 ( .A1(n11166), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11165) );
  NOR2_X1 U12125 ( .A1(n18045), .A2(n21208), .ZN(n20812) );
  NAND2_X1 U12126 ( .A1(n18103), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18080) );
  XNOR2_X1 U12127 ( .A(n17757), .B(n11177), .ZN(n18108) );
  INV_X1 U12128 ( .A(n17758), .ZN(n11177) );
  NAND2_X1 U12129 ( .A1(n18131), .A2(n17755), .ZN(n18119) );
  NAND2_X1 U12130 ( .A1(n18119), .A2(n18120), .ZN(n18118) );
  NOR2_X1 U12131 ( .A1(n17909), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17908) );
  NAND2_X1 U12132 ( .A1(n18012), .A2(n18051), .ZN(n17902) );
  INV_X1 U12133 ( .A(n20978), .ZN(n21151) );
  INV_X1 U12134 ( .A(n20994), .ZN(n21162) );
  INV_X1 U12135 ( .A(n11326), .ZN(n17775) );
  NOR2_X1 U12136 ( .A1(n18024), .A2(n17794), .ZN(n20978) );
  NAND2_X1 U12137 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17796), .ZN(
        n20976) );
  NOR2_X1 U12138 ( .A1(n21152), .A2(n20947), .ZN(n18033) );
  INV_X1 U12139 ( .A(n11316), .ZN(n11315) );
  OAI21_X1 U12140 ( .B1(n17729), .B2(n11317), .A(n17769), .ZN(n11316) );
  OR2_X1 U12141 ( .A1(n17976), .A2(n21208), .ZN(n17769) );
  NAND2_X1 U12142 ( .A1(n17764), .A2(n18075), .ZN(n20925) );
  NAND2_X1 U12143 ( .A1(n17761), .A2(n11186), .ZN(n18076) );
  AOI21_X1 U12144 ( .B1(n11185), .B2(n11039), .A(n11053), .ZN(n11186) );
  XNOR2_X1 U12145 ( .A(n17792), .B(n17727), .ZN(n18091) );
  INV_X1 U12146 ( .A(n17728), .ZN(n17727) );
  XNOR2_X1 U12147 ( .A(n17754), .B(n11178), .ZN(n18132) );
  INV_X1 U12148 ( .A(n17753), .ZN(n11178) );
  NAND2_X1 U12149 ( .A1(n18147), .A2(n17713), .ZN(n17715) );
  NAND2_X1 U12150 ( .A1(n11131), .A2(n17714), .ZN(n11130) );
  NAND2_X1 U12151 ( .A1(n18142), .A2(n18141), .ZN(n18140) );
  NAND2_X1 U12152 ( .A1(n18150), .A2(n17751), .ZN(n18137) );
  NAND2_X1 U12153 ( .A1(n18137), .A2(n18138), .ZN(n18136) );
  NOR2_X1 U12154 ( .A1(n18802), .A2(n15395), .ZN(n20803) );
  OAI21_X1 U12155 ( .B1(n15412), .B2(n15415), .A(n15416), .ZN(n21249) );
  NAND2_X1 U12156 ( .A1(n15387), .A2(n20615), .ZN(n20797) );
  NOR2_X2 U12157 ( .A1(n20054), .A2(n17730), .ZN(n21224) );
  NOR2_X1 U12158 ( .A1(n15336), .A2(n15335), .ZN(n19016) );
  NOR2_X1 U12159 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18678), .ZN(n18966) );
  NOR2_X1 U12160 ( .A1(n15326), .A2(n15325), .ZN(n18883) );
  INV_X1 U12161 ( .A(n20615), .ZN(n18802) );
  NOR2_X1 U12162 ( .A1(n11123), .A2(n11091), .ZN(n11090) );
  INV_X1 U12163 ( .A(n15359), .ZN(n11091) );
  NOR2_X1 U12164 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21144), .ZN(n17877) );
  NOR2_X1 U12165 ( .A1(n11105), .A2(n11104), .ZN(n11103) );
  NAND2_X1 U12166 ( .A1(n11112), .A2(n21246), .ZN(n11111) );
  NOR2_X1 U12167 ( .A1(n21561), .A2(n21539), .ZN(n21625) );
  AND2_X1 U12168 ( .A1(n13453), .A2(n13452), .ZN(n21651) );
  NAND2_X1 U12169 ( .A1(n13453), .A2(n13451), .ZN(n21539) );
  AND2_X1 U12170 ( .A1(n13453), .A2(n13444), .ZN(n21628) );
  XNOR2_X1 U12171 ( .A(n13355), .B(n14323), .ZN(n21477) );
  AND2_X1 U12172 ( .A1(n15559), .A2(n14722), .ZN(n21659) );
  INV_X1 U12173 ( .A(n21539), .ZN(n21562) );
  INV_X1 U12174 ( .A(n21628), .ZN(n21665) );
  INV_X1 U12175 ( .A(n21594), .ZN(n21601) );
  NOR2_X1 U12176 ( .A1(n15720), .A2(n14510), .ZN(n15264) );
  INV_X1 U12177 ( .A(n15264), .ZN(n15259) );
  OR2_X1 U12178 ( .A1(n14212), .A2(n14208), .ZN(n21857) );
  OR2_X2 U12179 ( .A1(n16832), .A2(n14271), .ZN(n21863) );
  INV_X1 U12180 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U12181 ( .A1(n11818), .A2(n11367), .ZN(n11365) );
  NAND2_X1 U12182 ( .A1(n19929), .A2(n13538), .ZN(n15242) );
  INV_X1 U12183 ( .A(n15874), .ZN(n19976) );
  INV_X1 U12184 ( .A(n21667), .ZN(n19978) );
  NAND2_X1 U12185 ( .A1(n11332), .A2(n19950), .ZN(n15965) );
  NAND2_X1 U12186 ( .A1(n15809), .A2(n13564), .ZN(n11332) );
  XNOR2_X1 U12187 ( .A(n11100), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n21422) );
  OAI21_X1 U12188 ( .B1(n19943), .B2(n11102), .A(n11101), .ZN(n11100) );
  OR2_X1 U12189 ( .A1(n15870), .A2(n19950), .ZN(n11102) );
  NAND2_X1 U12190 ( .A1(n19943), .A2(n19950), .ZN(n11101) );
  NAND2_X1 U12191 ( .A1(n19926), .A2(n13529), .ZN(n19931) );
  INV_X1 U12192 ( .A(n21430), .ZN(n21462) );
  INV_X1 U12193 ( .A(n21429), .ZN(n21461) );
  AND2_X1 U12194 ( .A1(n14264), .A2(n14263), .ZN(n21675) );
  INV_X1 U12195 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14465) );
  NOR2_X1 U12196 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U12197 ( .A1(n21989), .A2(n21867), .ZN(n22247) );
  INV_X1 U12198 ( .A(n21906), .ZN(n22272) );
  OAI21_X1 U12199 ( .B1(n14978), .B2(n14983), .A(n21998), .ZN(n15005) );
  OR2_X1 U12200 ( .A1(n14551), .A2(n11020), .ZN(n22277) );
  AND2_X1 U12201 ( .A1(n14633), .A2(n11020), .ZN(n22279) );
  OAI211_X1 U12202 ( .C1(n22284), .C2(n21930), .A(n21929), .B(n21952), .ZN(
        n22287) );
  NOR2_X2 U12203 ( .A1(n21939), .A2(n21983), .ZN(n22298) );
  NAND2_X1 U12204 ( .A1(n14602), .A2(n15721), .ZN(n21974) );
  NAND2_X1 U12205 ( .A1(n14602), .A2(n15715), .ZN(n22047) );
  NAND2_X1 U12206 ( .A1(n14602), .A2(n15703), .ZN(n22122) );
  NAND2_X1 U12207 ( .A1(n14602), .A2(n15697), .ZN(n22159) );
  NAND2_X1 U12208 ( .A1(n14602), .A2(n21805), .ZN(n22196) );
  NAND2_X1 U12209 ( .A1(n14602), .A2(n15686), .ZN(n22233) );
  NOR2_X1 U12210 ( .A1(n21939), .A2(n21866), .ZN(n22306) );
  AOI22_X1 U12211 ( .A1(n21964), .A2(n21970), .B1(n21991), .B2(n21963), .ZN(
        n22311) );
  OAI211_X1 U12212 ( .C1(n22319), .C2(n21999), .A(n21998), .B(n21997), .ZN(
        n22322) );
  NOR2_X2 U12213 ( .A1(n21984), .A2(n21983), .ZN(n22321) );
  INV_X1 U12214 ( .A(n21966), .ZN(n22010) );
  INV_X1 U12215 ( .A(n22043), .ZN(n22054) );
  INV_X1 U12216 ( .A(n22118), .ZN(n22129) );
  INV_X1 U12217 ( .A(n22155), .ZN(n22166) );
  INV_X1 U12218 ( .A(n22229), .ZN(n22240) );
  INV_X1 U12219 ( .A(n22304), .ZN(n22327) );
  INV_X1 U12220 ( .A(n22247), .ZN(n22331) );
  NAND2_X1 U12221 ( .A1(n21677), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21692) );
  AND2_X1 U12222 ( .A1(n16826), .A2(n16825), .ZN(n21693) );
  NOR2_X1 U12223 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21687) );
  INV_X1 U12224 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16839) );
  AND2_X1 U12225 ( .A1(n16839), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21677) );
  INV_X1 U12226 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21930) );
  NAND2_X1 U12227 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21716) );
  NAND2_X1 U12228 ( .A1(n13962), .A2(n13248), .ZN(n14100) );
  NAND2_X1 U12229 ( .A1(n18554), .A2(n18555), .ZN(n18553) );
  AND2_X1 U12230 ( .A1(n13869), .A2(n13859), .ZN(n18540) );
  NAND2_X1 U12231 ( .A1(n18504), .A2(n18505), .ZN(n18503) );
  NAND2_X1 U12232 ( .A1(n13844), .A2(n13286), .ZN(n13853) );
  NAND2_X1 U12233 ( .A1(n11216), .A2(n11215), .ZN(n16047) );
  AOI21_X1 U12234 ( .B1(n18584), .B2(n11217), .A(n13124), .ZN(n11215) );
  NAND2_X1 U12235 ( .A1(n18446), .A2(n18447), .ZN(n18445) );
  INV_X1 U12236 ( .A(n18561), .ZN(n18537) );
  OR3_X1 U12237 ( .A1(n17055), .A2(n13263), .A3(n13262), .ZN(n18520) );
  NAND2_X1 U12238 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n18520), .ZN(n18488) );
  INV_X1 U12239 ( .A(n18488), .ZN(n18577) );
  AND2_X1 U12240 ( .A1(n17055), .A2(n13250), .ZN(n18551) );
  INV_X1 U12241 ( .A(n18551), .ZN(n18578) );
  OR2_X1 U12242 ( .A1(n12622), .A2(n12621), .ZN(n15151) );
  CLKBUF_X1 U12243 ( .A(n15149), .Z(n15150) );
  OR2_X1 U12244 ( .A1(n12570), .A2(n12569), .ZN(n14905) );
  OR2_X1 U12245 ( .A1(n12558), .A2(n12557), .ZN(n14697) );
  AND2_X1 U12246 ( .A1(n11358), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11357) );
  OR2_X1 U12247 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  NAND2_X1 U12248 ( .A1(n16127), .A2(n12425), .ZN(n16178) );
  XNOR2_X1 U12249 ( .A(n15475), .B(n12844), .ZN(n16096) );
  INV_X1 U12250 ( .A(n16251), .ZN(n19615) );
  INV_X1 U12251 ( .A(n19619), .ZN(n16201) );
  XNOR2_X1 U12252 ( .A(n14413), .B(n14414), .ZN(n19254) );
  NAND2_X1 U12253 ( .A1(n12912), .A2(n18634), .ZN(n19613) );
  NOR2_X2 U12254 ( .A1(n19613), .A2(n12425), .ZN(n19619) );
  INV_X1 U12255 ( .A(n19398), .ZN(n19620) );
  NAND2_X1 U12256 ( .A1(n16250), .A2(n14372), .ZN(n14958) );
  BUF_X1 U12257 ( .A(n17200), .Z(n17211) );
  INV_X1 U12258 ( .A(n14131), .ZN(n14166) );
  OR3_X1 U12259 ( .A1(n14100), .A2(n12459), .A3(n18630), .ZN(n14268) );
  INV_X1 U12260 ( .A(n14166), .ZN(n14270) );
  OAI21_X1 U12261 ( .B1(n16101), .B2(n16103), .A(n16102), .ZN(n16450) );
  NAND2_X1 U12262 ( .A1(n13943), .A2(n13942), .ZN(n17071) );
  INV_X1 U12263 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17069) );
  INV_X1 U12264 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17064) );
  INV_X1 U12265 ( .A(n17133), .ZN(n17113) );
  OR2_X1 U12266 ( .A1(n18647), .A2(n18291), .ZN(n17119) );
  AND2_X1 U12267 ( .A1(n17117), .A2(n16785), .ZN(n17133) );
  OAI211_X1 U12268 ( .C1(n16733), .C2(n15498), .A(n15455), .B(n11405), .ZN(
        n15456) );
  OR2_X1 U12269 ( .A1(n16183), .A2(n16182), .ZN(n18549) );
  NAND2_X1 U12270 ( .A1(n16349), .A2(n13851), .ZN(n16340) );
  NAND2_X1 U12271 ( .A1(n14936), .A2(n11275), .ZN(n16260) );
  NAND2_X1 U12272 ( .A1(n16590), .A2(n16586), .ZN(n16740) );
  INV_X1 U12273 ( .A(n16730), .ZN(n18609) );
  INV_X1 U12274 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17147) );
  NAND2_X1 U12275 ( .A1(n15114), .A2(n14375), .ZN(n17144) );
  NAND2_X1 U12276 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17142) );
  INV_X1 U12277 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17156) );
  INV_X1 U12278 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19175) );
  NOR2_X2 U12279 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19321) );
  INV_X1 U12280 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16788) );
  INV_X1 U12281 ( .A(n19254), .ZN(n17161) );
  NAND2_X1 U12282 ( .A1(n15112), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16761) );
  OR2_X1 U12283 ( .A1(n14419), .A2(n14418), .ZN(n14420) );
  AOI21_X1 U12284 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n18631), .A(n15111), .ZN(
        n16762) );
  AOI21_X1 U12285 ( .B1(n19333), .B2(n19336), .A(n19330), .ZN(n19735) );
  INV_X1 U12286 ( .A(n19703), .ZN(n19705) );
  AND2_X1 U12287 ( .A1(n19242), .A2(n19239), .ZN(n19698) );
  AND2_X1 U12288 ( .A1(n19224), .A2(n19223), .ZN(n19675) );
  INV_X1 U12289 ( .A(n19367), .ZN(n19669) );
  AND2_X1 U12290 ( .A1(n19206), .A2(n19239), .ZN(n19674) );
  INV_X1 U12291 ( .A(n19724), .ZN(n19731) );
  INV_X1 U12292 ( .A(n19606), .ZN(n19610) );
  INV_X1 U12293 ( .A(n19565), .ZN(n19569) );
  INV_X1 U12294 ( .A(n19524), .ZN(n19528) );
  INV_X1 U12295 ( .A(n19435), .ZN(n19440) );
  INV_X1 U12296 ( .A(n18644), .ZN(n18634) );
  INV_X1 U12297 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18286) );
  OR2_X1 U12298 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21746), .ZN(n21736) );
  NOR2_X1 U12299 ( .A1(n20507), .A2(n20508), .ZN(n20513) );
  OAI21_X1 U12300 ( .B1(n20512), .B2(P3_REIP_REG_29__SCAN_IN), .A(n20511), 
        .ZN(n11159) );
  AND2_X1 U12301 ( .A1(n11153), .A2(n11152), .ZN(n20407) );
  INV_X1 U12302 ( .A(n20396), .ZN(n11152) );
  INV_X1 U12303 ( .A(n11153), .ZN(n20395) );
  NOR2_X1 U12304 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20359), .ZN(n20377) );
  NOR2_X1 U12305 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20194), .ZN(n20210) );
  NOR2_X1 U12306 ( .A1(n21258), .A2(n20118), .ZN(n20363) );
  AOI211_X2 U12307 ( .C1(n21274), .C2(n21273), .A(n20116), .B(n20115), .ZN(
        n20340) );
  INV_X1 U12308 ( .A(n20504), .ZN(n20543) );
  NOR2_X1 U12309 ( .A1(n20457), .A2(n17517), .ZN(n17522) );
  NOR2_X1 U12310 ( .A1(n20435), .A2(n17527), .ZN(n17533) );
  NOR2_X1 U12311 ( .A1(n20404), .A2(n17497), .ZN(n17534) );
  INV_X1 U12312 ( .A(n17587), .ZN(n17559) );
  NOR2_X1 U12313 ( .A1(n20364), .A2(n17601), .ZN(n17588) );
  NOR2_X1 U12314 ( .A1(n17572), .A2(n17379), .ZN(n17602) );
  NAND2_X1 U12315 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17602), .ZN(n17601) );
  NOR2_X1 U12316 ( .A1(n17571), .A2(n17348), .ZN(n17294) );
  NOR3_X2 U12317 ( .A1(n20800), .A2(n19016), .A3(n20551), .ZN(n17611) );
  NAND2_X1 U12318 ( .A1(n20671), .A2(n20707), .ZN(n20668) );
  INV_X1 U12319 ( .A(n20671), .ZN(n20664) );
  OR2_X1 U12320 ( .A1(n20675), .A2(n20669), .ZN(n20671) );
  NOR2_X1 U12321 ( .A1(n20680), .A2(n20681), .ZN(n20679) );
  NAND2_X1 U12322 ( .A1(n20679), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20675) );
  NOR2_X1 U12323 ( .A1(n20687), .A2(n20650), .ZN(n20656) );
  NAND2_X1 U12324 ( .A1(n20656), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20680) );
  NOR2_X1 U12325 ( .A1(n20693), .A2(n20649), .ZN(n20688) );
  NAND2_X1 U12326 ( .A1(n20688), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20687) );
  INV_X1 U12327 ( .A(n20620), .ZN(n20625) );
  INV_X1 U12328 ( .A(n20641), .ZN(n20637) );
  NAND2_X1 U12329 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20637), .ZN(n20636) );
  NOR2_X1 U12330 ( .A1(n17638), .A2(n17637), .ZN(n20596) );
  NOR2_X1 U12331 ( .A1(n17656), .A2(n11179), .ZN(n17657) );
  AND2_X1 U12332 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20609), .ZN(n20613) );
  INV_X2 U12333 ( .A(n20720), .ZN(n20707) );
  INV_X1 U12334 ( .A(n17660), .ZN(n11138) );
  NAND2_X1 U12335 ( .A1(n17618), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n17669) );
  NOR2_X1 U12336 ( .A1(n20734), .A2(n20746), .ZN(n20727) );
  NOR2_X1 U12337 ( .A1(n17708), .A2(n17707), .ZN(n20740) );
  INV_X1 U12338 ( .A(n20727), .ZN(n20739) );
  CLKBUF_X1 U12339 ( .A(n20098), .Z(n20110) );
  CLKBUF_X1 U12340 ( .A(n20080), .Z(n20109) );
  INV_X1 U12341 ( .A(n20393), .ZN(n20354) );
  NOR2_X1 U12342 ( .A1(n17927), .A2(n17922), .ZN(n18002) );
  NAND2_X1 U12343 ( .A1(n11314), .A2(n21102), .ZN(n17935) );
  NAND2_X1 U12344 ( .A1(n17935), .A2(n21101), .ZN(n21089) );
  NOR2_X1 U12345 ( .A1(n17790), .A2(n17804), .ZN(n18011) );
  INV_X1 U12346 ( .A(n18014), .ZN(n17958) );
  INV_X1 U12347 ( .A(n20964), .ZN(n17796) );
  NOR2_X2 U12348 ( .A1(n20811), .A2(n18170), .ZN(n18086) );
  NAND2_X1 U12349 ( .A1(n18113), .A2(n17724), .ZN(n18105) );
  INV_X1 U12350 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20180) );
  AND2_X1 U12351 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18129) );
  INV_X1 U12352 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18155) );
  INV_X1 U12353 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20130) );
  INV_X1 U12354 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20750) );
  OAI21_X1 U12355 ( .B1(n21045), .B2(n21128), .A(n21044), .ZN(n21066) );
  AND2_X1 U12356 ( .A1(n11303), .A2(n11304), .ZN(n17956) );
  AND2_X1 U12357 ( .A1(n17931), .A2(n17930), .ZN(n11303) );
  AND2_X1 U12358 ( .A1(n11326), .A2(n11327), .ZN(n18013) );
  NOR2_X1 U12359 ( .A1(n11319), .A2(n11318), .ZN(n11327) );
  INV_X1 U12360 ( .A(n11324), .ZN(n11318) );
  NAND2_X1 U12361 ( .A1(n18077), .A2(n18078), .ZN(n17815) );
  NAND2_X1 U12362 ( .A1(n21227), .A2(n20742), .ZN(n21213) );
  INV_X1 U12363 ( .A(n11185), .ZN(n18096) );
  NAND2_X1 U12364 ( .A1(n21216), .A2(n21087), .ZN(n20910) );
  INV_X1 U12365 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18721) );
  INV_X2 U12366 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21240) );
  NAND2_X1 U12367 ( .A1(n20775), .A2(n21240), .ZN(n20764) );
  INV_X1 U12368 ( .A(n11095), .ZN(n15399) );
  AOI211_X2 U12369 ( .C1(n21272), .C2(n21238), .A(n18680), .B(n15430), .ZN(
        n20795) );
  INV_X1 U12370 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19008) );
  INV_X1 U12371 ( .A(n21279), .ZN(n21272) );
  NAND2_X1 U12372 ( .A1(n21263), .A2(n11118), .ZN(n21268) );
  NAND2_X1 U12373 ( .A1(n21710), .A2(n21144), .ZN(n11118) );
  NOR2_X1 U12374 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21277), .ZN(n21274) );
  NOR2_X1 U12375 ( .A1(n21767), .A2(n21765), .ZN(n18269) );
  INV_X1 U12377 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19738) );
  NAND2_X1 U12378 ( .A1(n11244), .A2(n11242), .ZN(P1_U2842) );
  NAND2_X1 U12379 ( .A1(n15906), .A2(n13472), .ZN(n11244) );
  NOR2_X1 U12380 ( .A1(n11243), .A2(n13473), .ZN(n11242) );
  OR2_X1 U12381 ( .A1(n12302), .A2(n12301), .ZN(P1_U2875) );
  OR2_X1 U12382 ( .A1(n14058), .A2(n14057), .ZN(P1_U2876) );
  AOI21_X1 U12383 ( .B1(n15752), .B2(n19979), .A(n15751), .ZN(n15753) );
  INV_X1 U12384 ( .A(n15508), .ZN(n15752) );
  NOR4_X1 U12385 ( .A1(n15896), .A2(n15895), .A3(n15894), .A4(n15893), .ZN(
        n15897) );
  NAND2_X1 U12386 ( .A1(n13141), .A2(n18362), .ZN(n13302) );
  NAND2_X1 U12387 ( .A1(n18482), .A2(n18483), .ZN(n18481) );
  NAND2_X1 U12388 ( .A1(n16077), .A2(n16076), .ZN(n16075) );
  OAI21_X1 U12389 ( .B1(n15464), .B2(n17120), .A(n13954), .ZN(P2_U2984) );
  NAND2_X1 U12390 ( .A1(n14044), .A2(n11388), .ZN(n14045) );
  INV_X1 U12391 ( .A(n11261), .ZN(n16442) );
  OAI21_X1 U12392 ( .B1(n20513), .B2(n11160), .A(n11158), .ZN(P3_U2642) );
  INV_X1 U12393 ( .A(n11161), .ZN(n11160) );
  AOI211_X1 U12394 ( .C1(n20510), .C2(P3_REIP_REG_29__SCAN_IN), .A(n20509), 
        .B(n11159), .ZN(n11158) );
  AOI21_X1 U12395 ( .B1(n20507), .B2(n20508), .A(n20525), .ZN(n11161) );
  INV_X1 U12396 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20157) );
  AOI21_X1 U12397 ( .B1(n11190), .B2(n11188), .A(n11187), .ZN(n21070) );
  AND2_X1 U12398 ( .A1(n21113), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11187) );
  AOI21_X1 U12399 ( .B1(n21067), .B2(n21068), .A(n21154), .ZN(n11190) );
  AOI211_X1 U12400 ( .C1(n21100), .C2(n21099), .A(n21098), .B(n21097), .ZN(
        n21105) );
  OAI21_X1 U12401 ( .B1(n21268), .B2(n11117), .A(n11115), .ZN(P3_U2997) );
  NAND2_X1 U12402 ( .A1(n21259), .A2(n21274), .ZN(n11117) );
  NOR2_X1 U12403 ( .A1(n11088), .A2(n11116), .ZN(n11115) );
  NAND2_X1 U12404 ( .A1(n21260), .A2(n21261), .ZN(n11116) );
  OR2_X1 U12405 ( .A1(n19989), .A2(n20038), .ZN(U212) );
  CLKBUF_X3 U12406 ( .A(n15365), .Z(n17701) );
  OR2_X1 U12407 ( .A1(n15210), .A2(n11362), .ZN(n11032) );
  AND2_X1 U12408 ( .A1(n15595), .A2(n11372), .ZN(n15568) );
  NAND2_X1 U12409 ( .A1(n14079), .A2(n14081), .ZN(n14080) );
  AND2_X1 U12410 ( .A1(n11095), .A2(n11094), .ZN(n11033) );
  AND2_X1 U12411 ( .A1(n11225), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11034) );
  AND2_X2 U12412 ( .A1(n14238), .A2(n14460), .ZN(n11623) );
  AND4_X1 U12413 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11035) );
  NAND2_X1 U12414 ( .A1(n11385), .A2(n11872), .ZN(n15195) );
  OR2_X1 U12415 ( .A1(n18423), .A2(n13116), .ZN(n11036) );
  AND2_X1 U12416 ( .A1(n13759), .A2(n11145), .ZN(n11037) );
  INV_X2 U12417 ( .A(n16127), .ZN(n16176) );
  NAND2_X1 U12418 ( .A1(n14496), .A2(n14495), .ZN(n14489) );
  NAND2_X1 U12419 ( .A1(n11222), .A2(n11223), .ZN(n13104) );
  NAND2_X1 U12420 ( .A1(n11354), .A2(n11355), .ZN(n15048) );
  NAND2_X1 U12421 ( .A1(n11355), .A2(n15138), .ZN(n11353) );
  NOR2_X1 U12422 ( .A1(n17763), .A2(n20903), .ZN(n11039) );
  AND2_X1 U12423 ( .A1(n11156), .A2(n11071), .ZN(n11040) );
  AND2_X1 U12424 ( .A1(n15261), .A2(n15223), .ZN(n11041) );
  AND2_X1 U12425 ( .A1(n11168), .A2(n20451), .ZN(n11042) );
  OR2_X1 U12426 ( .A1(n19950), .A2(n15732), .ZN(n11043) );
  AND2_X1 U12427 ( .A1(n13132), .A2(n11081), .ZN(n13136) );
  AND2_X1 U12428 ( .A1(n11081), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11044) );
  AND2_X2 U12429 ( .A1(n14769), .A2(n12711), .ZN(n12551) );
  OR3_X1 U12430 ( .A1(n13118), .A2(n11228), .A3(n11227), .ZN(n11045) );
  AND2_X1 U12431 ( .A1(n11024), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12592) );
  AND2_X1 U12432 ( .A1(n11205), .A2(n11203), .ZN(n16344) );
  OR2_X1 U12433 ( .A1(n16102), .A2(n16092), .ZN(n11046) );
  INV_X1 U12434 ( .A(n12509), .ZN(n13143) );
  NOR2_X1 U12435 ( .A1(n11028), .A2(n17132), .ZN(n11047) );
  AND2_X1 U12436 ( .A1(n11247), .A2(n14901), .ZN(n11048) );
  NAND2_X1 U12437 ( .A1(n15595), .A2(n15647), .ZN(n15581) );
  AND2_X1 U12438 ( .A1(n11150), .A2(n13877), .ZN(n16269) );
  OR2_X1 U12439 ( .A1(n13939), .A2(n13945), .ZN(n11049) );
  NAND2_X1 U12440 ( .A1(n11299), .A2(n11300), .ZN(n16644) );
  AND2_X1 U12441 ( .A1(n11028), .A2(n15161), .ZN(n11050) );
  NOR3_X1 U12442 ( .A1(n16133), .A2(n11233), .A3(n11235), .ZN(n16101) );
  AND2_X1 U12443 ( .A1(n15871), .A2(n13556), .ZN(n11052) );
  OAI21_X1 U12444 ( .B1(n14414), .B2(n14413), .A(n12506), .ZN(n14418) );
  AND2_X1 U12445 ( .A1(n18098), .A2(n18097), .ZN(n11053) );
  NOR2_X1 U12446 ( .A1(n16119), .A2(n16118), .ZN(n16117) );
  AND2_X1 U12447 ( .A1(n14450), .A2(n11421), .ZN(n11622) );
  INV_X1 U12448 ( .A(n12238), .ZN(n11552) );
  NAND2_X1 U12449 ( .A1(n15595), .A2(n11374), .ZN(n11376) );
  AND2_X1 U12450 ( .A1(n11154), .A2(n13768), .ZN(n11054) );
  INV_X1 U12451 ( .A(n14307), .ZN(n11551) );
  AND2_X1 U12452 ( .A1(n13538), .A2(n13547), .ZN(n11055) );
  NAND2_X1 U12453 ( .A1(n11633), .A2(n11632), .ZN(n11696) );
  INV_X4 U12454 ( .A(n19935), .ZN(n19950) );
  AND4_X1 U12455 ( .A1(n15364), .A2(n15363), .A3(n15362), .A4(n15361), .ZN(
        n11056) );
  INV_X1 U12456 ( .A(n13851), .ZN(n11295) );
  OR2_X1 U12457 ( .A1(n13850), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13851) );
  OR2_X1 U12458 ( .A1(n13856), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11058) );
  AND2_X1 U12459 ( .A1(n13536), .A2(n13529), .ZN(n11059) );
  OR2_X1 U12460 ( .A1(n12908), .A2(n12457), .ZN(n11060) );
  AND2_X1 U12461 ( .A1(n15832), .A2(n15833), .ZN(n15848) );
  OR2_X1 U12462 ( .A1(n16283), .A2(n11302), .ZN(n11061) );
  INV_X1 U12463 ( .A(n11346), .ZN(n15831) );
  AND3_X1 U12464 ( .A1(n17654), .A2(n17655), .A3(n11181), .ZN(n11062) );
  NAND2_X1 U12465 ( .A1(n16122), .A2(n11408), .ZN(n12789) );
  AND2_X1 U12466 ( .A1(n11048), .A2(n11246), .ZN(n11063) );
  OR2_X1 U12467 ( .A1(n11386), .A2(n19008), .ZN(n11064) );
  AND2_X1 U12468 ( .A1(n12418), .A2(n12417), .ZN(n12421) );
  OR2_X1 U12469 ( .A1(n12425), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11407) );
  NAND4_X4 U12470 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13276) );
  AND3_X1 U12471 ( .A1(n11548), .A2(n11553), .A3(n14122), .ZN(n12278) );
  NAND2_X1 U12472 ( .A1(n14417), .A2(n12528), .ZN(n14496) );
  NAND2_X1 U12473 ( .A1(n13112), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13103) );
  AND2_X1 U12474 ( .A1(n14934), .A2(n14935), .ZN(n14936) );
  NOR2_X1 U12475 ( .A1(n15196), .A2(n11384), .ZN(n15228) );
  NAND2_X1 U12476 ( .A1(n13761), .A2(n13760), .ZN(n13762) );
  NOR2_X1 U12477 ( .A1(n15210), .A2(n11361), .ZN(n16148) );
  NOR2_X1 U12478 ( .A1(n15210), .A2(n16168), .ZN(n16158) );
  NOR2_X1 U12479 ( .A1(n14940), .A2(n13049), .ZN(n15022) );
  NOR2_X1 U12480 ( .A1(n14940), .A2(n11353), .ZN(n15136) );
  NAND2_X1 U12481 ( .A1(n11364), .A2(n11818), .ZN(n14909) );
  INV_X1 U12482 ( .A(n14049), .ZN(n11381) );
  AND4_X1 U12483 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13108) );
  NAND2_X1 U12484 ( .A1(n13761), .A2(n11054), .ZN(n13767) );
  AND2_X1 U12485 ( .A1(n14936), .A2(n11273), .ZN(n11065) );
  AND2_X1 U12486 ( .A1(n14081), .A2(n11237), .ZN(n11066) );
  NOR2_X1 U12487 ( .A1(n15050), .A2(n15051), .ZN(n15052) );
  AND2_X1 U12488 ( .A1(n14539), .A2(n11247), .ZN(n14700) );
  NOR2_X1 U12489 ( .A1(n18415), .A2(n18416), .ZN(n14934) );
  AND2_X1 U12490 ( .A1(n11276), .A2(n11278), .ZN(n11067) );
  NAND2_X1 U12491 ( .A1(n16237), .A2(n11284), .ZN(n16206) );
  NAND2_X1 U12492 ( .A1(n16718), .A2(n13759), .ZN(n16432) );
  INV_X1 U12493 ( .A(n13760), .ZN(n11155) );
  AND2_X1 U12494 ( .A1(n16237), .A2(n11285), .ZN(n16217) );
  NAND2_X1 U12495 ( .A1(n14834), .A2(n19628), .ZN(n13249) );
  NOR2_X1 U12496 ( .A1(n13105), .A2(n17069), .ZN(n13106) );
  NAND2_X1 U12497 ( .A1(n11342), .A2(n11341), .ZN(n19917) );
  OAI21_X1 U12498 ( .B1(n16138), .B2(n16139), .A(n12735), .ZN(n16130) );
  NOR2_X1 U12499 ( .A1(n20800), .A2(n15397), .ZN(n20061) );
  INV_X1 U12500 ( .A(n20061), .ZN(n11094) );
  NOR2_X1 U12501 ( .A1(n14910), .A2(n11365), .ZN(n15012) );
  AND2_X1 U12502 ( .A1(n16066), .A2(n16065), .ZN(n16064) );
  NAND2_X1 U12503 ( .A1(n11574), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11897) );
  INV_X1 U12504 ( .A(n11897), .ZN(n11942) );
  OR2_X1 U12505 ( .A1(n11872), .A2(n15220), .ZN(n11068) );
  AND2_X1 U12506 ( .A1(n11300), .A2(n11404), .ZN(n11069) );
  AND2_X1 U12507 ( .A1(n11066), .A2(n11236), .ZN(n11070) );
  INV_X1 U12508 ( .A(n14940), .ZN(n11354) );
  AND2_X1 U12509 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U12510 ( .A1(n13108), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13105) );
  AND2_X1 U12511 ( .A1(n18345), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16430) );
  AND2_X1 U12512 ( .A1(n13688), .A2(n13674), .ZN(n11072) );
  AND2_X1 U12513 ( .A1(n16152), .A2(n13219), .ZN(n16050) );
  AND2_X1 U12514 ( .A1(n17782), .A2(n11156), .ZN(n11073) );
  NAND2_X1 U12515 ( .A1(n17772), .A2(n17770), .ZN(n17827) );
  INV_X1 U12516 ( .A(n17827), .ZN(n11329) );
  AND2_X1 U12517 ( .A1(n13673), .A2(n13674), .ZN(n11074) );
  AND2_X1 U12518 ( .A1(n11942), .A2(n11704), .ZN(n11075) );
  AND2_X1 U12519 ( .A1(n11329), .A2(n11328), .ZN(n11076) );
  AND2_X1 U12520 ( .A1(n11034), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11077) );
  AND2_X1 U12521 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11078) );
  AND2_X1 U12522 ( .A1(n13761), .A2(n11154), .ZN(n11079) );
  INV_X1 U12523 ( .A(n12532), .ZN(n15481) );
  INV_X2 U12524 ( .A(n15485), .ZN(n12531) );
  INV_X1 U12525 ( .A(n18606), .ZN(n16733) );
  AND2_X1 U12526 ( .A1(n14496), .A2(n11358), .ZN(n14536) );
  NOR3_X1 U12527 ( .A1(n13118), .A2(n11228), .A3(n13098), .ZN(n13120) );
  AND2_X1 U12528 ( .A1(n11548), .A2(n14122), .ZN(n14235) );
  NOR2_X1 U12529 ( .A1(n14861), .A2(n14952), .ZN(n11080) );
  NOR2_X1 U12530 ( .A1(n11045), .A2(n16054), .ZN(n13123) );
  AND2_X1 U12531 ( .A1(n13112), .A2(n11077), .ZN(n13102) );
  NOR2_X1 U12532 ( .A1(n13127), .A2(n13126), .ZN(n13125) );
  INV_X1 U12533 ( .A(n16705), .ZN(n18611) );
  NOR2_X1 U12534 ( .A1(n13131), .A2(n13226), .ZN(n13132) );
  INV_X1 U12535 ( .A(n13795), .ZN(n11170) );
  NAND2_X1 U12536 ( .A1(n14539), .A2(n14881), .ZN(n14698) );
  AND2_X1 U12537 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11081) );
  AND2_X1 U12538 ( .A1(n13132), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13134) );
  AND2_X1 U12539 ( .A1(n16132), .A2(n11349), .ZN(n11082) );
  AND2_X1 U12540 ( .A1(n10983), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12675) );
  INV_X1 U12541 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11226) );
  OR2_X1 U12542 ( .A1(n12612), .A2(n12611), .ZN(n15138) );
  INV_X1 U12543 ( .A(n11251), .ZN(n11250) );
  OR2_X1 U12544 ( .A1(n11252), .A2(n15577), .ZN(n11251) );
  INV_X1 U12545 ( .A(n16115), .ZN(n11235) );
  AND2_X1 U12546 ( .A1(n15175), .A2(n13015), .ZN(n11083) );
  AND2_X1 U12547 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11084) );
  AND2_X1 U12548 ( .A1(n11273), .A2(n16246), .ZN(n11085) );
  OR2_X1 U12549 ( .A1(n13118), .A2(n11228), .ZN(n11086) );
  INV_X1 U12550 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U12551 ( .A1(n11328), .A2(n17771), .ZN(n11087) );
  NAND2_X1 U12552 ( .A1(n12532), .A2(n12373), .ZN(n11281) );
  INV_X1 U12553 ( .A(n12877), .ZN(n14835) );
  INV_X1 U12554 ( .A(n18592), .ZN(n11148) );
  AND2_X1 U12555 ( .A1(n21710), .A2(n18233), .ZN(n11088) );
  AND2_X1 U12556 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11089) );
  INV_X1 U12557 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11167) );
  INV_X1 U12558 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11157) );
  INV_X1 U12559 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11224) );
  NOR2_X1 U12560 ( .A1(n20810), .A2(n19015), .ZN(n18877) );
  NOR2_X1 U12561 ( .A1(n15316), .A2(n15315), .ZN(n20810) );
  NOR2_X4 U12563 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21765), .ZN(n18272) );
  AND2_X2 U12564 ( .A1(n11090), .A2(n11056), .ZN(n20799) );
  NAND3_X1 U12565 ( .A1(n20743), .A2(n17732), .A3(n20779), .ZN(n11095) );
  INV_X1 U12566 ( .A(n17731), .ZN(n20754) );
  NAND2_X1 U12567 ( .A1(n20743), .A2(n20779), .ZN(n17731) );
  INV_X2 U12568 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20772) );
  AND2_X2 U12569 ( .A1(n14463), .A2(n14460), .ZN(n11511) );
  AND2_X2 U12570 ( .A1(n11418), .A2(n14460), .ZN(n11669) );
  NAND2_X1 U12571 ( .A1(n11688), .A2(n11689), .ZN(n11645) );
  NAND2_X1 U12572 ( .A1(n11097), .A2(n11017), .ZN(n11520) );
  OAI21_X2 U12573 ( .B1(n14519), .B2(n13481), .A(n13476), .ZN(n14620) );
  INV_X1 U12574 ( .A(n11682), .ZN(n11099) );
  NAND2_X1 U12575 ( .A1(n14307), .A2(n12238), .ZN(n13486) );
  NAND2_X2 U12576 ( .A1(n10971), .A2(n11051), .ZN(n12238) );
  NAND2_X2 U12577 ( .A1(n19926), .A2(n11059), .ZN(n19929) );
  OR2_X2 U12578 ( .A1(n19924), .A2(n19923), .ZN(n19926) );
  NAND3_X1 U12579 ( .A1(n11111), .A2(n11106), .A3(n11103), .ZN(n21255) );
  NAND3_X1 U12580 ( .A1(n15347), .A2(n15355), .A3(n11121), .ZN(n11120) );
  NAND3_X1 U12581 ( .A1(n15358), .A2(n15356), .A3(n15357), .ZN(n11123) );
  INV_X1 U12582 ( .A(n17724), .ZN(n11126) );
  NAND3_X1 U12583 ( .A1(n11129), .A2(n11130), .A3(n11128), .ZN(n18142) );
  NAND3_X1 U12584 ( .A1(n18148), .A2(n18149), .A3(n17714), .ZN(n11128) );
  NAND2_X1 U12585 ( .A1(n18147), .A2(n11132), .ZN(n11129) );
  NAND2_X1 U12586 ( .A1(n18148), .A2(n18149), .ZN(n18147) );
  NAND3_X1 U12587 ( .A1(n17667), .A2(n11064), .A3(n11135), .ZN(n11134) );
  OR2_X2 U12588 ( .A1(n11138), .A2(n11310), .ZN(n20726) );
  NAND4_X1 U12589 ( .A1(n13637), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11298) );
  NAND2_X1 U12590 ( .A1(n12452), .A2(n12451), .ZN(n14017) );
  NAND2_X1 U12591 ( .A1(n14011), .A2(n12440), .ZN(n11143) );
  INV_X1 U12592 ( .A(n11144), .ZN(n12484) );
  NAND2_X1 U12593 ( .A1(n12517), .A2(n12518), .ZN(n11144) );
  NAND2_X1 U12594 ( .A1(n11144), .A2(n12486), .ZN(n13149) );
  AND2_X2 U12595 ( .A1(n14803), .A2(n15096), .ZN(n13615) );
  NAND2_X2 U12596 ( .A1(n13601), .A2(n15128), .ZN(n19218) );
  NOR2_X2 U12597 ( .A1(n13626), .A2(n13621), .ZN(n13601) );
  OR2_X2 U12598 ( .A1(n17111), .A2(n16626), .ZN(n16623) );
  NAND2_X2 U12599 ( .A1(n11147), .A2(n11146), .ZN(n17111) );
  INV_X1 U12600 ( .A(n14074), .ZN(n11146) );
  NAND2_X2 U12601 ( .A1(n11149), .A2(n11148), .ZN(n16651) );
  OAI21_X2 U12602 ( .B1(n16610), .B2(n14075), .A(n14076), .ZN(n14078) );
  OAI21_X2 U12603 ( .B1(n16418), .B2(n16420), .A(n16645), .ZN(n16610) );
  NAND2_X2 U12604 ( .A1(n11299), .A2(n11069), .ZN(n16418) );
  AOI21_X2 U12605 ( .B1(n16394), .B2(n16361), .A(n16360), .ZN(n16364) );
  OAI21_X2 U12606 ( .B1(n16409), .B2(n16406), .A(n16405), .ZN(n16394) );
  XNOR2_X1 U12607 ( .A(n13872), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16289) );
  NAND3_X1 U12608 ( .A1(n11061), .A2(n13870), .A3(n11151), .ZN(n11150) );
  INV_X1 U12609 ( .A(n16289), .ZN(n11151) );
  OR2_X2 U12610 ( .A1(n13767), .A2(n13772), .ZN(n13774) );
  INV_X1 U12611 ( .A(n11168), .ZN(n20453) );
  NAND2_X1 U12612 ( .A1(n12352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U12613 ( .A1(n12347), .A2(n12373), .ZN(n11172) );
  NAND2_X1 U12614 ( .A1(n15778), .A2(n13568), .ZN(n15731) );
  NAND2_X1 U12615 ( .A1(n15778), .A2(n11174), .ZN(n11338) );
  NAND3_X1 U12616 ( .A1(n17653), .A2(n11062), .A3(n11180), .ZN(n11179) );
  INV_X1 U12617 ( .A(n17762), .ZN(n17760) );
  NAND2_X1 U12618 ( .A1(n11297), .A2(n13669), .ZN(n13670) );
  NAND3_X1 U12619 ( .A1(n11192), .A2(n13665), .A3(n13666), .ZN(n11297) );
  NAND4_X1 U12620 ( .A1(n13650), .A2(n13645), .A3(n13649), .A4(n13642), .ZN(
        n11194) );
  NAND3_X2 U12621 ( .A1(n11198), .A2(n11196), .A3(n11195), .ZN(n13621) );
  NAND4_X1 U12622 ( .A1(n12517), .A2(n13148), .A3(n12518), .A4(n13150), .ZN(
        n11195) );
  OAI21_X1 U12623 ( .B1(n11287), .B2(n13150), .A(n11197), .ZN(n11196) );
  NAND2_X1 U12624 ( .A1(n13150), .A2(n12516), .ZN(n11197) );
  XNOR2_X2 U12625 ( .A(n11288), .B(n13153), .ZN(n13150) );
  INV_X1 U12626 ( .A(n12516), .ZN(n11200) );
  NAND2_X2 U12628 ( .A1(n13943), .A2(n11208), .ZN(n11205) );
  NAND2_X1 U12629 ( .A1(n11214), .A2(n18584), .ZN(n16048) );
  OR2_X1 U12630 ( .A1(n16060), .A2(n11217), .ZN(n11214) );
  NAND2_X1 U12631 ( .A1(n16060), .A2(n18584), .ZN(n11216) );
  NAND2_X1 U12632 ( .A1(n13132), .A2(n11044), .ZN(n13138) );
  INV_X1 U12633 ( .A(n13138), .ZN(n13099) );
  NAND2_X1 U12634 ( .A1(n15113), .A2(n11036), .ZN(n18446) );
  NAND3_X1 U12635 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13107) );
  INV_X1 U12636 ( .A(n11231), .ZN(n16102) );
  NOR3_X2 U12637 ( .A1(n16133), .A2(n11233), .A3(n11232), .ZN(n11231) );
  NOR3_X1 U12638 ( .A1(n16133), .A2(n16126), .A3(n11235), .ZN(n16110) );
  AND2_X2 U12639 ( .A1(n14539), .A2(n11063), .ZN(n15019) );
  NAND2_X1 U12640 ( .A1(n15637), .A2(n11249), .ZN(n15631) );
  INV_X1 U12641 ( .A(n15653), .ZN(n11258) );
  NAND2_X1 U12642 ( .A1(n13355), .A2(n11259), .ZN(n14508) );
  OR2_X1 U12643 ( .A1(n18563), .A2(n16733), .ZN(n11263) );
  NOR2_X4 U12644 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11286) );
  NOR2_X1 U12645 ( .A1(n13886), .A2(n11286), .ZN(n14791) );
  NAND2_X2 U12646 ( .A1(n12482), .A2(n12483), .ZN(n13148) );
  NAND2_X1 U12647 ( .A1(n16351), .A2(n11294), .ZN(n11293) );
  AOI21_X2 U12648 ( .B1(n11291), .B2(n13851), .A(n11290), .ZN(n11294) );
  INV_X1 U12649 ( .A(n16350), .ZN(n11291) );
  NAND3_X1 U12650 ( .A1(n11293), .A2(n11058), .A3(n11292), .ZN(n16280) );
  OAI21_X1 U12651 ( .B1(n16351), .B2(n11295), .A(n11294), .ZN(n16338) );
  NAND3_X1 U12652 ( .A1(n11297), .A2(n11298), .A3(n11296), .ZN(n13918) );
  NAND2_X1 U12653 ( .A1(n16653), .A2(n13777), .ZN(n11299) );
  NAND2_X1 U12654 ( .A1(n13995), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12507) );
  NAND2_X2 U12655 ( .A1(n12461), .A2(n12460), .ZN(n13995) );
  NAND2_X1 U12656 ( .A1(n13995), .A2(n11078), .ZN(n12511) );
  OAI211_X1 U12657 ( .C1(n21105), .C2(n21106), .A(n21104), .B(n21103), .ZN(
        P3_U2834) );
  NOR2_X1 U12658 ( .A1(n17903), .A2(n17915), .ZN(n11308) );
  INV_X1 U12659 ( .A(n17908), .ZN(n11309) );
  NAND4_X1 U12660 ( .A1(n17669), .A2(n11312), .A3(n17668), .A4(n11311), .ZN(
        n11310) );
  OAI21_X1 U12661 ( .B1(n17942), .B2(n17976), .A(n11314), .ZN(n21034) );
  NAND2_X1 U12662 ( .A1(n17942), .A2(n17976), .ZN(n11314) );
  AOI21_X1 U12663 ( .B1(n17827), .B2(n18051), .A(n11321), .ZN(n11320) );
  NAND2_X1 U12664 ( .A1(n15809), .A2(n11333), .ZN(n11331) );
  AND2_X2 U12665 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U12666 ( .A1(n11338), .A2(n11339), .ZN(n15744) );
  INV_X1 U12667 ( .A(n14940), .ZN(n11350) );
  NAND2_X1 U12668 ( .A1(n11350), .A2(n11351), .ZN(n15149) );
  NAND2_X1 U12669 ( .A1(n14496), .A2(n11357), .ZN(n14883) );
  NAND3_X1 U12670 ( .A1(n11364), .A2(n11366), .A3(n11818), .ZN(n15013) );
  NAND2_X1 U12671 ( .A1(n15595), .A2(n11371), .ZN(n15569) );
  INV_X1 U12672 ( .A(n11376), .ZN(n15582) );
  NOR2_X1 U12673 ( .A1(n11013), .A2(n14049), .ZN(n12207) );
  NOR2_X2 U12676 ( .A1(n14921), .A2(n13633), .ZN(n19178) );
  AND2_X1 U12677 ( .A1(n17147), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12882) );
  AND2_X2 U12678 ( .A1(n14768), .A2(n12711), .ZN(n13022) );
  AND2_X1 U12679 ( .A1(n15021), .A2(n15050), .ZN(n18389) );
  OR2_X2 U12681 ( .A1(n11758), .A2(n11724), .ZN(n11748) );
  NAND2_X1 U12682 ( .A1(n11650), .A2(n11649), .ZN(n11659) );
  AOI21_X1 U12683 ( .B1(n13987), .B2(n13986), .A(n13985), .ZN(n13993) );
  AOI211_X1 U12684 ( .C1(n16457), .C2(n18612), .A(n16456), .B(n16455), .ZN(
        n16458) );
  XNOR2_X1 U12685 ( .A(n14406), .B(n14405), .ZN(n19152) );
  AOI22_X1 U12686 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12343) );
  OAI21_X1 U12687 ( .B1(n12492), .B2(n12491), .A(n12506), .ZN(n14414) );
  NAND2_X1 U12688 ( .A1(n11698), .A2(n21683), .ZN(n11633) );
  NAND2_X1 U12689 ( .A1(n15554), .A2(n15555), .ZN(n15540) );
  NAND2_X1 U12690 ( .A1(n15527), .A2(n15528), .ZN(n14048) );
  AOI21_X2 U12691 ( .B1(n16418), .B2(n13843), .A(n13842), .ZN(n16351) );
  NOR2_X1 U12692 ( .A1(n15309), .A2(n15310), .ZN(n17341) );
  OR2_X1 U12693 ( .A1(n15460), .A2(n14031), .ZN(n11388) );
  OR2_X1 U12694 ( .A1(n20536), .A2(n20535), .ZN(n11389) );
  OR2_X1 U12695 ( .A1(n19950), .A2(n15757), .ZN(n11390) );
  NOR2_X1 U12696 ( .A1(n21924), .A2(n21944), .ZN(n11391) );
  AND2_X1 U12697 ( .A1(n12789), .A2(n11401), .ZN(n11392) );
  NOR2_X1 U12698 ( .A1(n15309), .A2(n15307), .ZN(n17364) );
  AND2_X1 U12699 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11393) );
  AND2_X1 U12700 ( .A1(n13680), .A2(n13675), .ZN(n11394) );
  AND2_X1 U12701 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21709), .ZN(n21713) );
  INV_X1 U12702 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12217) );
  NOR2_X1 U12703 ( .A1(n18583), .A2(n18585), .ZN(n11395) );
  NOR2_X1 U12704 ( .A1(n15166), .A2(n13753), .ZN(n11396) );
  NOR2_X1 U12705 ( .A1(n18286), .A2(n13904), .ZN(n11397) );
  INV_X1 U12706 ( .A(n12941), .ZN(n13039) );
  NAND2_X1 U12707 ( .A1(n12452), .A2(n12445), .ZN(n11398) );
  INV_X1 U12708 ( .A(n12751), .ZN(n12734) );
  AND2_X1 U12709 ( .A1(n12292), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14544)
         );
  INV_X1 U12710 ( .A(n14303), .ZN(n11554) );
  NAND2_X1 U12711 ( .A1(n17877), .A2(n18166), .ZN(n17967) );
  INV_X1 U12712 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13651) );
  INV_X1 U12713 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17964) );
  INV_X1 U12714 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16054) );
  AND2_X1 U12715 ( .A1(n10972), .A2(n15732), .ZN(n11399) );
  OR2_X1 U12716 ( .A1(n15761), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11400) );
  AND2_X1 U12717 ( .A1(n12788), .A2(n12809), .ZN(n11401) );
  INV_X1 U12718 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17978) );
  INV_X1 U12719 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16769) );
  OR2_X1 U12720 ( .A1(n18647), .A2(n19574), .ZN(n17120) );
  AND2_X1 U12721 ( .A1(n18620), .A2(n12448), .ZN(n11402) );
  INV_X1 U12722 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16320) );
  INV_X1 U12723 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14031) );
  INV_X1 U12724 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17094) );
  AND2_X1 U12725 ( .A1(n15835), .A2(n21427), .ZN(n11403) );
  INV_X1 U12726 ( .A(n18522), .ZN(n13297) );
  OR2_X1 U12727 ( .A1(n18383), .A2(n13788), .ZN(n11404) );
  OR4_X1 U12728 ( .A1(n15454), .A2(n16437), .A3(n16443), .A4(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11405) );
  NOR2_X1 U12729 ( .A1(n15308), .A2(n15307), .ZN(n17652) );
  INV_X1 U12730 ( .A(n21935), .ZN(n22015) );
  INV_X1 U12731 ( .A(n22015), .ZN(n21982) );
  INV_X2 U12732 ( .A(n18751), .ZN(n19011) );
  NAND2_X1 U12733 ( .A1(n13751), .A2(n13750), .ZN(n13931) );
  AND2_X1 U12734 ( .A1(n12975), .A2(n12943), .ZN(n11406) );
  OR2_X1 U12735 ( .A1(n16131), .A2(n12773), .ZN(n11408) );
  AND2_X1 U12736 ( .A1(n11537), .A2(n11536), .ZN(n11409) );
  INV_X1 U12737 ( .A(n14331), .ZN(n11575) );
  OR2_X1 U12738 ( .A1(n12228), .A2(n12242), .ZN(n12213) );
  NAND2_X1 U12739 ( .A1(n13698), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13624) );
  AND2_X1 U12740 ( .A1(n12215), .A2(n12214), .ZN(n12226) );
  OR2_X1 U12741 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12217), .ZN(
        n12220) );
  NAND2_X1 U12742 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  INV_X1 U12743 ( .A(n12440), .ZN(n12433) );
  AOI22_X1 U12744 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12350) );
  OR2_X1 U12745 ( .A1(n11677), .A2(n11676), .ZN(n13474) );
  NAND2_X1 U12746 ( .A1(n14018), .A2(n12433), .ZN(n12434) );
  NAND2_X1 U12747 ( .A1(n12415), .A2(n12428), .ZN(n13963) );
  AOI22_X1 U12748 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12370) );
  INV_X1 U12749 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11412) );
  BUF_X1 U12750 ( .A(n11964), .Z(n13312) );
  AND2_X1 U12751 ( .A1(n11759), .A2(n14522), .ZN(n11760) );
  AND2_X1 U12752 ( .A1(n19950), .A2(n13554), .ZN(n13555) );
  INV_X1 U12753 ( .A(n13484), .ZN(n11609) );
  NOR2_X1 U12754 ( .A1(n11635), .A2(n21683), .ZN(n11611) );
  NAND2_X1 U12755 ( .A1(n12445), .A2(n18291), .ZN(n12446) );
  NAND2_X1 U12756 ( .A1(n12532), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12303) );
  AND2_X1 U12757 ( .A1(n11773), .A2(n11772), .ZN(n11796) );
  INV_X1 U12758 ( .A(n11808), .ZN(n11809) );
  NAND2_X1 U12759 ( .A1(n15446), .A2(n14356), .ZN(n13422) );
  NAND2_X1 U12760 ( .A1(n11611), .A2(n11553), .ZN(n12258) );
  INV_X1 U12761 ( .A(n13931), .ZN(n13753) );
  NAND2_X1 U12762 ( .A1(n13915), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13916) );
  INV_X1 U12763 ( .A(n13630), .ZN(n13631) );
  AND2_X1 U12764 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  NAND2_X1 U12765 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11539) );
  INV_X1 U12766 ( .A(n15197), .ZN(n11872) );
  AND2_X1 U12767 ( .A1(n12168), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12169) );
  NAND2_X1 U12768 ( .A1(n16033), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13326) );
  INV_X1 U12769 ( .A(n13329), .ZN(n11975) );
  INV_X1 U12770 ( .A(n13422), .ZN(n13432) );
  INV_X1 U12771 ( .A(n19932), .ZN(n13536) );
  INV_X1 U12772 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U12773 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12324) );
  INV_X1 U12774 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13904) );
  NOR2_X1 U12775 ( .A1(n13876), .A2(n13875), .ZN(n13877) );
  AND2_X1 U12776 ( .A1(n13069), .A2(n13068), .ZN(n16259) );
  AND2_X1 U12777 ( .A1(n15078), .A2(n13276), .ZN(n16654) );
  NAND2_X1 U12779 ( .A1(n17976), .A2(n21012), .ZN(n17930) );
  INV_X1 U12780 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17714) );
  NAND2_X1 U12781 ( .A1(n20610), .A2(n20726), .ZN(n17710) );
  AOI21_X1 U12782 ( .B1(n15426), .B2(n15423), .A(n20803), .ZN(n15392) );
  INV_X1 U12783 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11866) );
  OR2_X1 U12784 ( .A1(n14254), .A2(n14120), .ZN(n14117) );
  NAND2_X1 U12785 ( .A1(n12169), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13303) );
  INV_X1 U12786 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U12787 ( .A1(n11894), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11916) );
  INV_X1 U12788 ( .A(n12163), .ZN(n12204) );
  NAND2_X1 U12789 ( .A1(n11390), .A2(n15758), .ZN(n15759) );
  AND2_X1 U12790 ( .A1(n15847), .A2(n15848), .ZN(n15999) );
  AND2_X1 U12791 ( .A1(n12238), .A2(n13348), .ZN(n13521) );
  NAND2_X1 U12792 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  NAND2_X1 U12793 ( .A1(n11709), .A2(n11708), .ZN(n21960) );
  AND3_X1 U12794 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21683), .A3(n14557), 
        .ZN(n14603) );
  OR2_X1 U12795 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11753) );
  INV_X1 U12796 ( .A(n16198), .ZN(n13084) );
  AND2_X1 U12797 ( .A1(n12787), .A2(n12786), .ZN(n12805) );
  AND2_X1 U12798 ( .A1(n18291), .A2(n19293), .ZN(n12941) );
  OR2_X1 U12799 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  OR2_X1 U12800 ( .A1(n19674), .A2(n19213), .ZN(n19214) );
  AND2_X1 U12801 ( .A1(n20383), .A2(n20382), .ZN(n20384) );
  INV_X1 U12802 ( .A(n20810), .ZN(n17239) );
  INV_X1 U12803 ( .A(n17967), .ZN(n17879) );
  INV_X1 U12804 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15612) );
  INV_X1 U12805 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15278) );
  INV_X1 U12806 ( .A(n21652), .ZN(n21570) );
  OR2_X1 U12807 ( .A1(n21286), .A2(n13342), .ZN(n15559) );
  AND3_X1 U12808 ( .A1(n13426), .A2(n13425), .A3(n13424), .ZN(n15628) );
  INV_X1 U12809 ( .A(n14507), .ZN(n13358) );
  NAND2_X1 U12810 ( .A1(n12298), .A2(n15202), .ZN(n15724) );
  INV_X1 U12811 ( .A(n11788), .ZN(n12163) );
  NAND2_X1 U12812 ( .A1(n12144), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12167) );
  NOR2_X1 U12813 ( .A1(n12012), .A2(n15603), .ZN(n12013) );
  INV_X1 U12814 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U12815 ( .A1(n21667), .A2(n13586), .ZN(n15874) );
  OAI21_X1 U12816 ( .B1(n13571), .B2(n19950), .A(n13570), .ZN(n13572) );
  AND2_X1 U12817 ( .A1(n13386), .A2(n13385), .ZN(n19894) );
  AND2_X1 U12818 ( .A1(n21349), .A2(n21334), .ZN(n21426) );
  NAND2_X1 U12819 ( .A1(n12272), .A2(n12271), .ZN(n14310) );
  OR2_X1 U12820 ( .A1(n21894), .A2(n21987), .ZN(n22261) );
  AND2_X1 U12821 ( .A1(n16028), .A2(n14445), .ZN(n21943) );
  NOR2_X1 U12822 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21935) );
  OR2_X1 U12823 ( .A1(n14521), .A2(n14677), .ZN(n21939) );
  OR2_X1 U12824 ( .A1(n14520), .A2(n21865), .ZN(n21920) );
  AOI21_X1 U12825 ( .B1(n21975), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21871), 
        .ZN(n22017) );
  INV_X1 U12826 ( .A(n11753), .ZN(n13339) );
  AND2_X1 U12827 ( .A1(n18584), .A2(n15094), .ZN(n15122) );
  INV_X1 U12828 ( .A(n13994), .ZN(n13247) );
  NOR2_X1 U12829 ( .A1(n12545), .A2(n12544), .ZN(n14884) );
  INV_X1 U12830 ( .A(n12525), .ZN(n14419) );
  INV_X1 U12831 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16398) );
  AND2_X1 U12832 ( .A1(n13203), .A2(n13202), .ZN(n16167) );
  INV_X1 U12833 ( .A(n16281), .ZN(n16327) );
  AND2_X1 U12834 ( .A1(n18437), .A2(n13830), .ZN(n16406) );
  INV_X1 U12835 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15062) );
  INV_X1 U12836 ( .A(n16396), .ZN(n18381) );
  AOI21_X1 U12837 ( .B1(n18637), .B2(n18286), .A(n17045), .ZN(n19327) );
  INV_X1 U12838 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19293) );
  INV_X1 U12839 ( .A(n19287), .ZN(n19315) );
  INV_X1 U12840 ( .A(n19242), .ZN(n17160) );
  AND2_X1 U12841 ( .A1(n19214), .A2(n19322), .ZN(n19221) );
  NAND2_X1 U12842 ( .A1(n19152), .A2(n17144), .ZN(n19316) );
  OR2_X1 U12843 ( .A1(n19152), .A2(n17144), .ZN(n19160) );
  INV_X1 U12844 ( .A(n12502), .ZN(n14848) );
  NOR2_X1 U12845 ( .A1(n20393), .A2(n20384), .ZN(n20385) );
  NAND2_X1 U12846 ( .A1(n20363), .A2(n20362), .ZN(n20428) );
  NOR2_X1 U12847 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20267), .ZN(n20283) );
  NOR2_X1 U12848 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20241), .ZN(n20260) );
  INV_X1 U12849 ( .A(n20368), .ZN(n20525) );
  NOR2_X1 U12850 ( .A1(n20808), .A2(n17730), .ZN(n17241) );
  NOR2_X1 U12851 ( .A1(n20722), .A2(n20721), .ZN(n20719) );
  AOI211_X1 U12852 ( .C1(n17701), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15343), .B(n15342), .ZN(n15344) );
  AND2_X1 U12853 ( .A1(n20649), .A2(n20584), .ZN(n20720) );
  OR2_X1 U12854 ( .A1(n20062), .A2(n21710), .ZN(n20553) );
  NOR2_X1 U12855 ( .A1(n20976), .A2(n21051), .ZN(n21046) );
  INV_X1 U12856 ( .A(n18088), .ZN(n18034) );
  INV_X1 U12857 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21208) );
  NAND2_X1 U12858 ( .A1(n17974), .A2(n17973), .ZN(n17995) );
  INV_X1 U12859 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17794) );
  INV_X1 U12860 ( .A(n21153), .ZN(n21130) );
  NOR2_X1 U12861 ( .A1(n20755), .A2(n20753), .ZN(n20744) );
  INV_X1 U12862 ( .A(n21223), .ZN(n21128) );
  AOI21_X1 U12863 ( .B1(n21267), .B2(n17614), .A(n20792), .ZN(n18678) );
  INV_X1 U12864 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21241) );
  NOR2_X1 U12865 ( .A1(n15386), .A2(n15385), .ZN(n20807) );
  AOI211_X1 U12866 ( .C1(n15429), .C2(n21764), .A(n17241), .B(n20804), .ZN(
        n21256) );
  INV_X1 U12867 ( .A(n14271), .ZN(n13338) );
  OAI21_X1 U12868 ( .B1(n15879), .B2(n21665), .A(n13457), .ZN(n13458) );
  INV_X1 U12869 ( .A(n21625), .ZN(n21638) );
  AND2_X1 U12870 ( .A1(n15559), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21652) );
  AND2_X1 U12871 ( .A1(n15559), .A2(n13346), .ZN(n21661) );
  AND2_X1 U12872 ( .A1(n12298), .A2(n14544), .ZN(n15729) );
  INV_X1 U12873 ( .A(n15260), .ZN(n15720) );
  INV_X1 U12874 ( .A(n21801), .ZN(n21858) );
  NAND2_X1 U12875 ( .A1(n15750), .A2(n15749), .ZN(n15751) );
  NAND2_X1 U12876 ( .A1(n12049), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12091) );
  NAND2_X1 U12877 ( .A1(n12013), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U12878 ( .A1(n11961), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11979) );
  AND2_X1 U12879 ( .A1(n11832), .A2(n11831), .ZN(n15028) );
  NOR2_X1 U12880 ( .A1(n11726), .A2(n14893), .ZN(n11799) );
  AND2_X1 U12881 ( .A1(n15874), .A2(n13588), .ZN(n19965) );
  INV_X1 U12882 ( .A(n21334), .ZN(n21407) );
  NAND2_X1 U12883 ( .A1(n16038), .A2(n21683), .ZN(n13585) );
  OAI22_X1 U12884 ( .A1(n21334), .A2(n21351), .B1(n16003), .B2(n21319), .ZN(
        n21396) );
  INV_X1 U12885 ( .A(n21349), .ZN(n21330) );
  NOR2_X1 U12886 ( .A1(n21930), .A2(n14310), .ZN(n21686) );
  INV_X1 U12887 ( .A(n21686), .ZN(n21671) );
  INV_X1 U12888 ( .A(n21876), .ZN(n22255) );
  INV_X1 U12889 ( .A(n22259), .ZN(n22263) );
  INV_X1 U12890 ( .A(n22261), .ZN(n22271) );
  INV_X1 U12891 ( .A(n14979), .ZN(n15009) );
  INV_X1 U12892 ( .A(n22277), .ZN(n14607) );
  OAI211_X1 U12893 ( .C1(n21982), .C2(n14550), .A(n14549), .B(n22017), .ZN(
        n14599) );
  AND2_X1 U12894 ( .A1(n21910), .A2(n21962), .ZN(n21916) );
  OAI211_X1 U12895 ( .C1(n21982), .C2(n14635), .A(n14632), .B(n22017), .ZN(
        n14661) );
  AND2_X1 U12896 ( .A1(n14633), .A2(n21865), .ZN(n22286) );
  INV_X1 U12897 ( .A(n21939), .ZN(n21921) );
  AND2_X1 U12898 ( .A1(n21943), .A2(n21962), .ZN(n21953) );
  NOR2_X2 U12899 ( .A1(n21939), .A2(n21987), .ZN(n22297) );
  AND2_X1 U12900 ( .A1(n14518), .A2(n14517), .ZN(n15709) );
  INV_X1 U12901 ( .A(n21871), .ZN(n14602) );
  INV_X1 U12902 ( .A(n21920), .ZN(n21957) );
  INV_X1 U12903 ( .A(n22081), .ZN(n22092) );
  INV_X1 U12904 ( .A(n22192), .ZN(n22203) );
  INV_X1 U12905 ( .A(n22310), .ZN(n22329) );
  NOR2_X1 U12906 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21722), .ZN(n21724) );
  INV_X1 U12907 ( .A(n21720), .ZN(n19858) );
  NOR2_X1 U12908 ( .A1(n14833), .A2(n14765), .ZN(n13962) );
  NAND3_X1 U12909 ( .A1(n14093), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18644) );
  NAND2_X1 U12910 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  INV_X1 U12911 ( .A(n16237), .ZN(n16238) );
  NAND2_X1 U12912 ( .A1(n18458), .A2(n18459), .ZN(n18457) );
  INV_X1 U12913 ( .A(n18520), .ZN(n18576) );
  NAND2_X1 U12914 ( .A1(n18573), .A2(n13260), .ZN(n18561) );
  OR2_X1 U12915 ( .A1(n12699), .A2(n12698), .ZN(n16145) );
  OR2_X1 U12916 ( .A1(n12602), .A2(n12601), .ZN(n15049) );
  INV_X1 U12917 ( .A(n14404), .ZN(n14406) );
  INV_X1 U12918 ( .A(n14267), .ZN(n14220) );
  INV_X1 U12919 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16084) );
  AND2_X1 U12920 ( .A1(n14945), .A2(n14944), .ZN(n18367) );
  INV_X1 U12921 ( .A(n17120), .ZN(n17135) );
  INV_X1 U12922 ( .A(n17117), .ZN(n17126) );
  NOR2_X1 U12923 ( .A1(n16723), .A2(n16702), .ZN(n18615) );
  AND2_X1 U12924 ( .A1(n13982), .A2(n18634), .ZN(n14036) );
  INV_X1 U12925 ( .A(n18604), .ZN(n18612) );
  AND2_X1 U12926 ( .A1(n14036), .A2(n14008), .ZN(n18606) );
  INV_X1 U12927 ( .A(n19327), .ZN(n19313) );
  AOI22_X1 U12928 ( .A1(n19338), .A2(n19337), .B1(n19336), .B2(n19335), .ZN(
        n19730) );
  NOR2_X2 U12929 ( .A1(n19316), .A2(n19315), .ZN(n19732) );
  OAI21_X1 U12930 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(n19699) );
  OAI21_X1 U12931 ( .B1(n19246), .B2(n19257), .A(n19245), .ZN(n19693) );
  OAI211_X1 U12932 ( .C1(n19221), .C2(n19216), .A(n19313), .B(n19215), .ZN(
        n19676) );
  AND2_X1 U12933 ( .A1(n19206), .A2(n19286), .ZN(n19462) );
  NOR2_X1 U12934 ( .A1(n19255), .A2(n17161), .ZN(n19206) );
  INV_X1 U12935 ( .A(n19319), .ZN(n19339) );
  INV_X1 U12936 ( .A(n19483), .ZN(n19488) );
  INV_X1 U12937 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21746) );
  NAND2_X1 U12938 ( .A1(n21272), .A2(n21228), .ZN(n20062) );
  INV_X1 U12939 ( .A(n21249), .ZN(n21228) );
  NOR2_X1 U12940 ( .A1(n20475), .A2(n20474), .ZN(n20514) );
  NOR2_X1 U12941 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20405), .ZN(n20432) );
  NOR2_X1 U12942 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20380), .ZN(n20401) );
  NOR2_X1 U12943 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20323), .ZN(n20348) );
  NOR2_X1 U12944 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20294), .ZN(n20317) );
  NOR2_X1 U12945 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20214), .ZN(n20240) );
  INV_X1 U12946 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20153) );
  INV_X1 U12947 ( .A(n20340), .ZN(n20547) );
  AND2_X1 U12948 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17559), .ZN(n17484) );
  NAND2_X1 U12949 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17294), .ZN(n17379) );
  INV_X1 U12950 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20181) );
  INV_X1 U12951 ( .A(n20649), .ZN(n20585) );
  NOR2_X1 U12952 ( .A1(n20631), .A2(n20636), .ZN(n20630) );
  NAND2_X1 U12953 ( .A1(n20702), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20701) );
  NAND3_X1 U12954 ( .A1(n17628), .A2(n17627), .A3(n17626), .ZN(n21086) );
  INV_X1 U12955 ( .A(n19016), .ZN(n20113) );
  NOR2_X1 U12956 ( .A1(n20110), .A2(n20063), .ZN(n20080) );
  NOR2_X1 U12957 ( .A1(n11094), .A2(n20553), .ZN(n20098) );
  NOR3_X2 U12958 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18156), .A3(n20750), 
        .ZN(n18006) );
  INV_X1 U12959 ( .A(n20812), .ZN(n21152) );
  AOI21_X2 U12960 ( .B1(n20058), .B2(n21277), .A(n21282), .ZN(n18156) );
  AND2_X1 U12961 ( .A1(n21080), .A2(n21216), .ZN(n21081) );
  NOR2_X1 U12962 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21267), .ZN(n17765) );
  NOR2_X2 U12963 ( .A1(n20796), .A2(n21175), .ZN(n21223) );
  NOR2_X2 U12964 ( .A1(n20811), .A2(n20910), .ZN(n21220) );
  NOR2_X1 U12965 ( .A1(n21154), .A2(n21128), .ZN(n21014) );
  NOR2_X1 U12966 ( .A1(n20800), .A2(n21175), .ZN(n21087) );
  NOR2_X1 U12967 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21264), .ZN(
        n20792) );
  NAND2_X1 U12968 ( .A1(n18173), .A2(n18966), .ZN(n18751) );
  INV_X1 U12969 ( .A(n18951), .ZN(n19109) );
  INV_X1 U12970 ( .A(n18993), .ZN(n19091) );
  INV_X1 U12971 ( .A(n19066), .ZN(n19079) );
  INV_X1 U12972 ( .A(n19060), .ZN(n19073) );
  INV_X1 U12973 ( .A(n19048), .ZN(n19062) );
  INV_X1 U12974 ( .A(n18980), .ZN(n19056) );
  INV_X1 U12975 ( .A(n19042), .ZN(n19050) );
  INV_X1 U12976 ( .A(n19036), .ZN(n19044) );
  INV_X1 U12977 ( .A(n18834), .ZN(n18838) );
  INV_X1 U12978 ( .A(n18748), .ZN(n18755) );
  INV_X1 U12979 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21144) );
  INV_X1 U12980 ( .A(n21764), .ZN(n21710) );
  INV_X1 U12981 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21709) );
  NAND2_X1 U12982 ( .A1(n12278), .A2(n13338), .ZN(n14212) );
  INV_X1 U12983 ( .A(n21286), .ZN(n15450) );
  INV_X1 U12984 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21936) );
  INV_X1 U12985 ( .A(n13458), .ZN(n13459) );
  INV_X1 U12986 ( .A(n21661), .ZN(n21591) );
  INV_X1 U12987 ( .A(n21651), .ZN(n21649) );
  INV_X1 U12988 ( .A(n21659), .ZN(n21642) );
  NAND2_X1 U12989 ( .A1(n19911), .A2(n13471), .ZN(n15657) );
  OR2_X1 U12990 ( .A1(n14056), .A2(n14055), .ZN(n14057) );
  NAND2_X1 U12991 ( .A1(n19801), .A2(n11553), .ZN(n14434) );
  INV_X1 U12992 ( .A(n19801), .ZN(n19820) );
  INV_X1 U12993 ( .A(n21843), .ZN(n21801) );
  OR2_X1 U12994 ( .A1(n15249), .A2(n15251), .ZN(n21592) );
  INV_X1 U12995 ( .A(n19965), .ZN(n19982) );
  NAND2_X1 U12996 ( .A1(n14334), .A2(n14320), .ZN(n21430) );
  INV_X1 U12997 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U12998 ( .A1(n21874), .A2(n21872), .B1(n11391), .B2(n21945), .ZN(
        n22252) );
  OR2_X1 U12999 ( .A1(n21894), .A2(n21983), .ZN(n22259) );
  AOI22_X1 U13000 ( .A1(n21887), .A2(n21890), .B1(n21911), .B2(n21945), .ZN(
        n22267) );
  OR2_X1 U13001 ( .A1(n21894), .A2(n21866), .ZN(n22269) );
  OR2_X1 U13002 ( .A1(n14551), .A2(n21865), .ZN(n14979) );
  AOI22_X1 U13003 ( .A1(n21912), .A2(n21916), .B1(n21991), .B2(n21911), .ZN(
        n22283) );
  INV_X1 U13004 ( .A(n22279), .ZN(n14660) );
  NAND2_X1 U13005 ( .A1(n21921), .A2(n21957), .ZN(n22295) );
  AOI22_X1 U13006 ( .A1(n21946), .A2(n21953), .B1(n21945), .B2(n21992), .ZN(
        n22302) );
  INV_X1 U13007 ( .A(n14682), .ZN(n14764) );
  NAND2_X1 U13008 ( .A1(n14602), .A2(n15709), .ZN(n22085) );
  NAND2_X1 U13009 ( .A1(n14602), .A2(n15681), .ZN(n22310) );
  NAND2_X1 U13010 ( .A1(n21989), .A2(n21957), .ZN(n22317) );
  INV_X1 U13011 ( .A(n22000), .ZN(n22022) );
  NAND2_X1 U13012 ( .A1(n21989), .A2(n21988), .ZN(n22335) );
  INV_X1 U13013 ( .A(n21696), .ZN(n16802) );
  OR2_X1 U13014 ( .A1(n13447), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21726) );
  NAND2_X1 U13015 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22339), .ZN(n21720) );
  INV_X1 U13016 ( .A(n19855), .ZN(n19860) );
  NAND2_X1 U13017 ( .A1(n14100), .A2(n18307), .ZN(n17055) );
  INV_X1 U13018 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21698) );
  AND2_X1 U13019 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  NAND2_X1 U13020 ( .A1(n17055), .A2(n13296), .ZN(n18522) );
  OR2_X1 U13021 ( .A1(n14833), .A2(n14146), .ZN(n18307) );
  NAND2_X1 U13022 ( .A1(n14417), .A2(n14420), .ZN(n19255) );
  AND2_X1 U13023 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  INV_X1 U13024 ( .A(n19613), .ZN(n16250) );
  AND2_X1 U13025 ( .A1(n16201), .A2(n19398), .ZN(n19404) );
  NAND2_X1 U13026 ( .A1(n16250), .A2(n12942), .ZN(n19398) );
  NAND2_X1 U13027 ( .A1(n17180), .A2(n12445), .ZN(n14402) );
  INV_X1 U13028 ( .A(n17180), .ZN(n17213) );
  OAI21_X1 U13029 ( .B1(n14100), .B2(n18630), .A(n14267), .ZN(n14131) );
  OR2_X1 U13030 ( .A1(n14100), .A2(n18291), .ZN(n14267) );
  INV_X1 U13031 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18413) );
  INV_X1 U13032 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18382) );
  INV_X1 U13033 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17079) );
  NOR2_X1 U13034 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  NAND2_X1 U13035 ( .A1(n14036), .A2(n14033), .ZN(n18604) );
  NAND2_X1 U13036 ( .A1(n14036), .A2(n13983), .ZN(n16730) );
  INV_X1 U13037 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19302) );
  INV_X1 U13038 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19531) );
  NAND2_X1 U13039 ( .A1(n19287), .A2(n19286), .ZN(n19723) );
  AOI21_X1 U13040 ( .B1(n19278), .B2(n19277), .A(n19276), .ZN(n19710) );
  NAND2_X1 U13041 ( .A1(n19287), .A2(n19256), .ZN(n19703) );
  NAND2_X1 U13042 ( .A1(n19242), .A2(n19286), .ZN(n19696) );
  NAND2_X1 U13043 ( .A1(n19256), .A2(n19242), .ZN(n19684) );
  AND2_X1 U13044 ( .A1(n19205), .A2(n19204), .ZN(n19367) );
  INV_X1 U13045 ( .A(n19462), .ZN(n19672) );
  NAND2_X1 U13046 ( .A1(n19256), .A2(n19206), .ZN(n19660) );
  NAND2_X1 U13047 ( .A1(n19140), .A2(n19286), .ZN(n19648) );
  INV_X1 U13048 ( .A(n19727), .ZN(n19636) );
  INV_X1 U13049 ( .A(n21701), .ZN(n17178) );
  INV_X1 U13050 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21752) );
  INV_X1 U13051 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21703) );
  AOI21_X1 U13052 ( .B1(n20538), .B2(n20537), .A(n11389), .ZN(n20539) );
  INV_X1 U13053 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20473) );
  INV_X1 U13054 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20239) );
  AND2_X1 U13055 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17522), .ZN(n17516) );
  AND2_X1 U13056 ( .A1(n17611), .A2(n20649), .ZN(n17609) );
  INV_X2 U13057 ( .A(n17609), .ZN(n17606) );
  INV_X1 U13058 ( .A(n21086), .ZN(n20811) );
  NOR2_X1 U13059 ( .A1(n17649), .A2(n17648), .ZN(n20605) );
  NAND2_X1 U13060 ( .A1(n18217), .A2(n20113), .ZN(n18235) );
  INV_X1 U13061 ( .A(n18217), .ZN(n18216) );
  OR4_X1 U13062 ( .A1(n17959), .A2(n17958), .A3(n21016), .A4(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17960) );
  INV_X1 U13063 ( .A(n18086), .ZN(n18035) );
  INV_X1 U13064 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21195) );
  NAND2_X1 U13065 ( .A1(n21282), .A2(n20796), .ZN(n18170) );
  INV_X1 U13066 ( .A(n21220), .ZN(n21139) );
  INV_X1 U13067 ( .A(n21216), .ZN(n21154) );
  NAND2_X1 U13068 ( .A1(n21199), .A2(n21154), .ZN(n21186) );
  INV_X1 U13069 ( .A(n21014), .ZN(n21008) );
  INV_X1 U13070 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18683) );
  INV_X1 U13071 ( .A(n20795), .ZN(n20793) );
  INV_X1 U13072 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18841) );
  INV_X1 U13073 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18760) );
  INV_X1 U13074 ( .A(n19069), .ZN(n19054) );
  INV_X1 U13075 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21277) );
  INV_X1 U13076 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21264) );
  INV_X1 U13077 ( .A(n16773), .ZN(n21706) );
  NAND2_X1 U13078 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21764) );
  INV_X1 U13079 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20898) );
  INV_X1 U13080 ( .A(n18272), .ZN(n18271) );
  NOR2_X1 U13081 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14072), .ZN(n19010)
         );
  INV_X1 U13082 ( .A(n19797), .ZN(n19786) );
  OAI211_X1 U13083 ( .C1(n14067), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        P1_U2874) );
  OAI21_X1 U13084 ( .B1(n13302), .B2(n11395), .A(n13301), .ZN(P2_U2825) );
  INV_X1 U13085 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U13086 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12174), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11417) );
  INV_X1 U13087 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11411) );
  AND2_X2 U13088 ( .A1(n11413), .A2(n11418), .ZN(n11663) );
  NOR2_X2 U13089 ( .A1(n11412), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11420) );
  NOR2_X4 U13090 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11419) );
  AND2_X2 U13091 ( .A1(n11420), .A2(n11419), .ZN(n11735) );
  AOI22_X1 U13092 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U13093 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U13094 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11414) );
  AND2_X2 U13095 ( .A1(n11418), .A2(n11419), .ZN(n11601) );
  AOI22_X1 U13096 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11425) );
  AND2_X2 U13097 ( .A1(n11419), .A2(n14238), .ZN(n11964) );
  AOI22_X1 U13098 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U13099 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U13100 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11422) );
  AND2_X4 U13101 ( .A1(n11427), .A2(n11426), .ZN(n11574) );
  AOI22_X1 U13102 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U13103 ( .A1(n12174), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U13104 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11710), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U13105 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11669), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U13106 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11583), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U13107 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11511), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U13108 ( .A1(n11016), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U13109 ( .A1(n11574), .A2(n12238), .ZN(n12282) );
  NAND2_X1 U13110 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11439) );
  NAND2_X1 U13111 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11438) );
  NAND2_X1 U13112 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11437) );
  NAND2_X1 U13113 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11436) );
  NAND2_X1 U13114 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11443) );
  NAND2_X1 U13115 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U13116 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U13117 ( .A1(n11622), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11440) );
  NAND2_X1 U13118 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11446) );
  NAND2_X1 U13119 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11445) );
  NAND2_X1 U13120 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11444) );
  NAND2_X1 U13121 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11451) );
  NAND2_X1 U13122 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11450) );
  NAND2_X1 U13123 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U13124 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11448) );
  INV_X2 U13125 ( .A(n11547), .ZN(n14564) );
  NAND2_X1 U13126 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11459) );
  NAND2_X1 U13127 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U13128 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11457) );
  NAND2_X1 U13129 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U13130 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U13131 ( .A1(n12174), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U13132 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11461) );
  NAND2_X1 U13133 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11460) );
  NAND2_X1 U13134 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U13135 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U13136 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11464) );
  NAND3_X1 U13137 ( .A1(n11466), .A2(n11465), .A3(n11464), .ZN(n11467) );
  NAND2_X1 U13138 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11471) );
  NAND2_X1 U13139 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11470) );
  NAND2_X1 U13140 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U13141 ( .A1(n11622), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11468) );
  NAND2_X1 U13142 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U13143 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11479) );
  NAND2_X1 U13144 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11478) );
  NAND2_X1 U13145 ( .A1(n11622), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U13146 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11484) );
  NAND2_X1 U13147 ( .A1(n12174), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11483) );
  NAND2_X1 U13148 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11482) );
  NAND2_X1 U13149 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11481) );
  NAND2_X1 U13150 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U13151 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11487) );
  NAND2_X1 U13152 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11486) );
  NAND2_X1 U13153 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11485) );
  NAND2_X1 U13154 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U13155 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U13156 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11490) );
  NAND2_X1 U13157 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11489) );
  NAND4_X4 U13158 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(
        n11553) );
  AOI22_X1 U13159 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U13160 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U13161 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U13162 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11497) );
  NAND4_X1 U13163 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11506) );
  AOI22_X1 U13164 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U13165 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U13166 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U13167 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U13168 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  AND2_X1 U13169 ( .A1(n11017), .A2(n11571), .ZN(n13477) );
  AOI22_X1 U13170 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11021), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U13171 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11664), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U13172 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U13173 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11583), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U13174 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11601), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U13175 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11622), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U13176 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11512) );
  AND2_X2 U13177 ( .A1(n11547), .A2(n12238), .ZN(n13583) );
  NAND2_X1 U13178 ( .A1(n13583), .A2(n11018), .ZN(n11516) );
  AOI22_X1 U13179 ( .A1(n11558), .A2(n13477), .B1(n11551), .B2(n11516), .ZN(
        n11521) );
  NAND2_X1 U13180 ( .A1(n14564), .A2(n11574), .ZN(n11517) );
  NAND2_X1 U13181 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  AND2_X1 U13182 ( .A1(n11521), .A2(n11520), .ZN(n14233) );
  NAND2_X1 U13183 ( .A1(n11552), .A2(n11522), .ZN(n11523) );
  NAND2_X1 U13184 ( .A1(n13581), .A2(n11635), .ZN(n14230) );
  NAND2_X1 U13185 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U13186 ( .A1(n11671), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U13187 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U13188 ( .A1(n11511), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11524) );
  NAND2_X1 U13189 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U13190 ( .A1(n11663), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U13191 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U13192 ( .A1(n11601), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U13193 ( .A1(n12174), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U13194 ( .A1(n11664), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U13195 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11533) );
  NAND2_X1 U13196 ( .A1(n11583), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U13197 ( .A1(n11669), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U13198 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U13199 ( .A1(n11622), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11536) );
  NAND4_X4 U13200 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n13348) );
  NAND2_X1 U13201 ( .A1(n13583), .A2(n13364), .ZN(n11544) );
  NAND2_X1 U13202 ( .A1(n11017), .A2(n13348), .ZN(n14255) );
  NAND2_X1 U13203 ( .A1(n11544), .A2(n14255), .ZN(n11545) );
  AOI21_X1 U13204 ( .B1(n14230), .B2(n14214), .A(n11545), .ZN(n11546) );
  NAND2_X1 U13205 ( .A1(n11552), .A2(n11547), .ZN(n12276) );
  AOI21_X1 U13206 ( .B1(n21722), .B2(P1_STATE_REG_2__SCAN_IN), .A(n21724), 
        .ZN(n13447) );
  NAND2_X1 U13207 ( .A1(n11549), .A2(n13447), .ZN(n11550) );
  NAND2_X1 U13208 ( .A1(n12278), .A2(n11550), .ZN(n11556) );
  NAND2_X1 U13209 ( .A1(n14570), .A2(n14578), .ZN(n14303) );
  NAND2_X1 U13210 ( .A1(n10970), .A2(n11554), .ZN(n14316) );
  INV_X1 U13211 ( .A(n11571), .ZN(n13347) );
  NAND2_X1 U13212 ( .A1(n13583), .A2(n13347), .ZN(n11555) );
  INV_X1 U13213 ( .A(n14230), .ZN(n11557) );
  NAND2_X1 U13214 ( .A1(n11557), .A2(n12282), .ZN(n11559) );
  NAND2_X1 U13215 ( .A1(n11559), .A2(n11558), .ZN(n11570) );
  INV_X1 U13216 ( .A(n11031), .ZN(n11560) );
  NAND3_X1 U13217 ( .A1(n11569), .A2(n11565), .A3(n11561), .ZN(n11562) );
  XNOR2_X1 U13218 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21923) );
  OR2_X1 U13219 ( .A1(n21677), .A2(n21965), .ZN(n11646) );
  OAI21_X1 U13220 ( .B1(n13585), .B2(n21923), .A(n11646), .ZN(n11563) );
  INV_X1 U13221 ( .A(n11563), .ZN(n11564) );
  OAI21_X2 U13222 ( .B1(n11651), .B2(n11412), .A(n11564), .ZN(n11567) );
  INV_X1 U13223 ( .A(n11565), .ZN(n11566) );
  MUX2_X1 U13224 ( .A(n13585), .B(n21677), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11568) );
  OAI21_X2 U13225 ( .B1(n11651), .B2(n14281), .A(n11568), .ZN(n11617) );
  INV_X1 U13226 ( .A(n11570), .ZN(n11579) );
  INV_X1 U13227 ( .A(n14715), .ZN(n15447) );
  NAND2_X1 U13228 ( .A1(n12282), .A2(n11571), .ZN(n11572) );
  AND2_X1 U13229 ( .A1(n15447), .A2(n11572), .ZN(n11573) );
  NAND2_X1 U13230 ( .A1(n11031), .A2(n11574), .ZN(n14331) );
  NAND2_X1 U13231 ( .A1(n16038), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19986) );
  AOI21_X1 U13232 ( .B1(n11579), .B2(n13348), .A(n11578), .ZN(n11580) );
  NAND2_X1 U13233 ( .A1(n11569), .A2(n11580), .ZN(n11615) );
  NAND2_X1 U13234 ( .A1(n11617), .A2(n11615), .ZN(n11581) );
  OR2_X2 U13235 ( .A1(n14628), .A2(n11581), .ZN(n11650) );
  NAND2_X1 U13236 ( .A1(n11014), .A2(n11581), .ZN(n14548) );
  AOI22_X1 U13237 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U13238 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U13239 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13240 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U13241 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11595) );
  AOI22_X1 U13242 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U13243 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U13244 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U13245 ( .A1(n11711), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U13246 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11594) );
  AOI22_X1 U13247 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14448), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13248 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U13249 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U13250 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U13251 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11608) );
  AOI22_X1 U13252 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13253 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U13254 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13255 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U13256 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  OAI22_X1 U13257 ( .A1(n11662), .A2(n13543), .B1(n11661), .B2(n11609), .ZN(
        n11610) );
  INV_X1 U13258 ( .A(n11610), .ZN(n11614) );
  INV_X1 U13259 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11612) );
  OR2_X1 U13260 ( .A1(n12258), .A2(n11612), .ZN(n11613) );
  INV_X1 U13261 ( .A(n11662), .ZN(n11631) );
  AOI22_X1 U13262 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U13263 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U13264 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U13265 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U13266 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n11629) );
  AOI22_X1 U13267 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U13268 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U13269 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U13270 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11624) );
  NAND4_X1 U13271 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11628) );
  XNOR2_X1 U13272 ( .A(n11637), .B(n13543), .ZN(n11630) );
  NAND2_X1 U13273 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  INV_X1 U13274 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U13275 ( .A1(n11635), .A2(n13543), .ZN(n11636) );
  OAI211_X1 U13276 ( .C1(n11637), .C2(n11553), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n11636), .ZN(n11638) );
  INV_X1 U13277 ( .A(n11638), .ZN(n11639) );
  INV_X1 U13278 ( .A(n13543), .ZN(n11641) );
  INV_X1 U13279 ( .A(n13489), .ZN(n11643) );
  NAND2_X1 U13280 ( .A1(n11643), .A2(n11642), .ZN(n11644) );
  NAND2_X1 U13281 ( .A1(n11645), .A2(n11644), .ZN(n11682) );
  INV_X1 U13282 ( .A(n11646), .ZN(n11648) );
  OAI21_X1 U13283 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11648), .A(
        n11647), .ZN(n11649) );
  NAND2_X1 U13284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U13285 ( .A1(n21922), .A2(n11652), .ZN(n11654) );
  NAND2_X1 U13286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22007) );
  INV_X1 U13287 ( .A(n22007), .ZN(n11653) );
  NAND2_X1 U13288 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11653), .ZN(
        n22004) );
  NAND2_X1 U13289 ( .A1(n11654), .A2(n22004), .ZN(n14980) );
  OAI22_X1 U13290 ( .A1(n13585), .A2(n14980), .B1(n21677), .B2(n21922), .ZN(
        n11655) );
  INV_X1 U13291 ( .A(n11655), .ZN(n11656) );
  INV_X1 U13292 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U13293 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U13294 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U13295 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U13296 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U13297 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11677) );
  AOI22_X1 U13298 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U13299 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U13300 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U13301 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11672) );
  NAND4_X1 U13302 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n11676) );
  NAND2_X1 U13303 ( .A1(n12248), .A2(n13474), .ZN(n11678) );
  OAI21_X1 U13304 ( .B1(n12258), .B2(n11679), .A(n11678), .ZN(n11680) );
  NAND2_X1 U13305 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  NAND2_X1 U13306 ( .A1(n11554), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11749) );
  XNOR2_X1 U13307 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14723) );
  AOI21_X1 U13308 ( .B1(n13339), .B2(n14723), .A(n13329), .ZN(n11685) );
  NAND2_X1 U13309 ( .A1(n12204), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11684) );
  OAI211_X1 U13310 ( .C1(n11749), .C2(n11015), .A(n11685), .B(n11684), .ZN(
        n11686) );
  INV_X1 U13311 ( .A(n11686), .ZN(n11687) );
  NAND2_X1 U13312 ( .A1(n13329), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11704) );
  INV_X1 U13313 ( .A(n14506), .ZN(n11703) );
  XNOR2_X2 U13314 ( .A(n11688), .B(n11689), .ZN(n14520) );
  NAND2_X1 U13315 ( .A1(n14520), .A2(n11942), .ZN(n11694) );
  INV_X1 U13316 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21474) );
  NOR2_X1 U13317 ( .A1(n21474), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11690) );
  AOI21_X1 U13318 ( .B1(n12204), .B2(P1_EAX_REG_1__SCAN_IN), .A(n11690), .ZN(
        n11691) );
  OAI21_X1 U13319 ( .B1(n11749), .B2(n11412), .A(n11691), .ZN(n11692) );
  INV_X1 U13320 ( .A(n11692), .ZN(n11693) );
  NAND2_X1 U13321 ( .A1(n11694), .A2(n11693), .ZN(n14366) );
  NAND2_X1 U13322 ( .A1(n11020), .A2(n11574), .ZN(n11697) );
  NAND2_X1 U13323 ( .A1(n11697), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U13324 ( .A1(n11788), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n22008), .ZN(n11699) );
  OAI21_X1 U13325 ( .B1(n14281), .B2(n11749), .A(n11699), .ZN(n11700) );
  AOI21_X1 U13326 ( .B1(n11698), .B2(n11942), .A(n11700), .ZN(n14289) );
  OR2_X1 U13327 ( .A1(n14288), .A2(n14289), .ZN(n14286) );
  NAND2_X1 U13328 ( .A1(n14289), .A2(n13339), .ZN(n11701) );
  NAND2_X1 U13329 ( .A1(n14286), .A2(n11701), .ZN(n14365) );
  NAND2_X1 U13330 ( .A1(n14366), .A2(n14365), .ZN(n14505) );
  NAND2_X1 U13331 ( .A1(n11703), .A2(n11702), .ZN(n14503) );
  INV_X1 U13332 ( .A(n13585), .ZN(n11707) );
  INV_X1 U13333 ( .A(n22004), .ZN(n11705) );
  NAND2_X1 U13334 ( .A1(n11705), .A2(n12217), .ZN(n14662) );
  NAND2_X1 U13335 ( .A1(n22004), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U13336 ( .A1(n14662), .A2(n11706), .ZN(n21924) );
  INV_X1 U13337 ( .A(n21677), .ZN(n16828) );
  AOI22_X1 U13338 ( .A1(n11707), .A2(n21924), .B1(n16828), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U13339 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U13340 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U13341 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U13342 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11712) );
  NAND4_X1 U13343 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11721) );
  AOI22_X1 U13344 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U13345 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U13346 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U13347 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U13348 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11720) );
  AOI22_X1 U13349 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12248), .B2(n13503), .ZN(n11722) );
  INV_X1 U13350 ( .A(n14522), .ZN(n11724) );
  NAND2_X1 U13351 ( .A1(n11758), .A2(n11724), .ZN(n11725) );
  OR2_X2 U13352 ( .A1(n14521), .A2(n11897), .ZN(n11733) );
  NAND2_X1 U13353 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11726) );
  INV_X1 U13354 ( .A(n11726), .ZN(n11728) );
  INV_X1 U13355 ( .A(n11799), .ZN(n11727) );
  OAI21_X1 U13356 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11728), .A(
        n11727), .ZN(n14888) );
  AOI22_X1 U13357 ( .A1(n13339), .A2(n14888), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U13358 ( .A1(n12204), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11729) );
  OAI211_X1 U13359 ( .C1(n11749), .C2(n11335), .A(n11730), .B(n11729), .ZN(
        n11731) );
  INV_X1 U13360 ( .A(n11731), .ZN(n11732) );
  INV_X1 U13361 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11734) );
  OR2_X1 U13362 ( .A1(n12258), .A2(n11734), .ZN(n11747) );
  AOI22_X1 U13363 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14448), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U13364 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11582), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U13365 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13305), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U13366 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U13367 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11745) );
  AOI22_X1 U13368 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11589), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U13369 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U13370 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U13371 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U13372 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11744) );
  NAND2_X1 U13373 ( .A1(n12248), .A2(n13511), .ZN(n11746) );
  NAND2_X1 U13374 ( .A1(n11747), .A2(n11746), .ZN(n11759) );
  XNOR2_X1 U13375 ( .A(n11748), .B(n11759), .ZN(n13507) );
  INV_X1 U13376 ( .A(n11749), .ZN(n11750) );
  NAND2_X1 U13377 ( .A1(n11750), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11756) );
  INV_X1 U13378 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11751) );
  AOI21_X1 U13379 ( .B1(n11751), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11752) );
  AOI21_X1 U13380 ( .B1(n12204), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11752), .ZN(
        n11755) );
  XNOR2_X1 U13381 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n11799), .ZN(
        n21493) );
  NOR2_X1 U13382 ( .A1(n21493), .A2(n11753), .ZN(n11754) );
  AOI21_X1 U13383 ( .B1(n11756), .B2(n11755), .A(n11754), .ZN(n11757) );
  AOI21_X1 U13384 ( .B1(n13507), .B2(n11942), .A(n11757), .ZN(n14708) );
  INV_X1 U13385 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11761) );
  OR2_X1 U13386 ( .A1(n12258), .A2(n11761), .ZN(n11773) );
  AOI22_X1 U13387 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U13388 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U13389 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U13390 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11762) );
  NAND4_X1 U13391 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n11771) );
  AOI22_X1 U13392 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U13393 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U13394 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U13395 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U13396 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11770) );
  NAND2_X1 U13397 ( .A1(n12248), .A2(n13523), .ZN(n11772) );
  INV_X1 U13398 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11774) );
  OR2_X1 U13399 ( .A1(n12258), .A2(n11774), .ZN(n11786) );
  AOI22_X1 U13400 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U13401 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U13402 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13403 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11775) );
  NAND4_X1 U13404 ( .A1(n11778), .A2(n11777), .A3(n11776), .A4(n11775), .ZN(
        n11784) );
  AOI22_X1 U13405 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U13406 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U13407 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U13408 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U13409 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  NAND2_X1 U13410 ( .A1(n12248), .A2(n13532), .ZN(n11785) );
  INV_X1 U13411 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11794) );
  INV_X1 U13412 ( .A(n11814), .ZN(n11791) );
  INV_X1 U13413 ( .A(n11789), .ZN(n11803) );
  INV_X1 U13414 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21510) );
  NAND2_X1 U13415 ( .A1(n11803), .A2(n21510), .ZN(n11790) );
  NAND2_X1 U13416 ( .A1(n11791), .A2(n11790), .ZN(n21512) );
  NOR2_X1 U13417 ( .A1(n11975), .A2(n21510), .ZN(n11792) );
  AOI21_X1 U13418 ( .B1(n21512), .B2(n13339), .A(n11792), .ZN(n11793) );
  OAI21_X1 U13419 ( .B1(n12163), .B2(n11794), .A(n11793), .ZN(n11795) );
  AOI21_X1 U13420 ( .B1(n13520), .B2(n11942), .A(n11795), .ZN(n14950) );
  INV_X1 U13421 ( .A(n14950), .ZN(n11806) );
  NAND2_X1 U13422 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  NAND2_X1 U13423 ( .A1(n11787), .A2(n11798), .ZN(n13516) );
  INV_X1 U13424 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U13425 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11799), .ZN(
        n11800) );
  NAND2_X1 U13426 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  NAND2_X1 U13427 ( .A1(n11803), .A2(n11802), .ZN(n21499) );
  AOI22_X1 U13428 ( .A1(n21499), .A2(n13339), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U13429 ( .A1(n12204), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11804) );
  AND2_X1 U13430 ( .A1(n11806), .A2(n14855), .ZN(n11807) );
  INV_X1 U13431 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U13432 ( .A1(n12248), .A2(n13543), .ZN(n11811) );
  OAI21_X1 U13433 ( .B1(n12258), .B2(n11812), .A(n11811), .ZN(n11813) );
  INV_X1 U13434 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11816) );
  OAI21_X1 U13435 ( .B1(n11814), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11833), .ZN(n21524) );
  AOI22_X1 U13436 ( .A1(n21524), .A2(n13339), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11815) );
  OAI21_X1 U13437 ( .B1(n12163), .B2(n11816), .A(n11815), .ZN(n11817) );
  XNOR2_X1 U13438 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11833), .ZN(
        n21534) );
  INV_X1 U13439 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15245) );
  OAI22_X1 U13440 ( .A1(n11753), .A2(n21534), .B1(n11975), .B2(n15245), .ZN(
        n11819) );
  AOI21_X1 U13441 ( .B1(n12204), .B2(P1_EAX_REG_8__SCAN_IN), .A(n11819), .ZN(
        n11832) );
  AOI22_X1 U13442 ( .A1(n11711), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U13443 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U13444 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U13445 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11820) );
  NAND4_X1 U13446 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11830) );
  AOI22_X1 U13447 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14448), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U13448 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U13449 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U13450 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U13451 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11829) );
  OAI21_X1 U13452 ( .B1(n11830), .B2(n11829), .A(n11942), .ZN(n11831) );
  XOR2_X1 U13453 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11848), .Z(n21549) );
  AOI22_X1 U13454 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U13455 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U13456 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U13457 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U13458 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11844) );
  AOI22_X1 U13459 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U13460 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U13461 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U13462 ( .A1(n11711), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U13463 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11843) );
  OR2_X1 U13464 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  AOI22_X1 U13465 ( .A1(n11942), .A2(n11845), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U13466 ( .A1(n11788), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11846) );
  OAI211_X1 U13467 ( .C1(n21549), .C2(n11753), .A(n11847), .B(n11846), .ZN(
        n15015) );
  INV_X1 U13468 ( .A(n15013), .ZN(n11865) );
  XNOR2_X1 U13469 ( .A(n11867), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n21560) );
  INV_X1 U13470 ( .A(n21560), .ZN(n11863) );
  AOI22_X1 U13471 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11582), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U13472 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U13473 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U13474 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11849) );
  NAND4_X1 U13475 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11858) );
  AOI22_X1 U13476 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U13477 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U13478 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U13479 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U13480 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  NOR2_X1 U13481 ( .A1(n11858), .A2(n11857), .ZN(n11861) );
  NAND2_X1 U13482 ( .A1(n13329), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11860) );
  NAND2_X1 U13483 ( .A1(n11788), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U13484 ( .C1(n11897), .C2(n11861), .A(n11860), .B(n11859), .ZN(
        n11862) );
  AOI21_X1 U13485 ( .B1(n11863), .B2(n13339), .A(n11862), .ZN(n15118) );
  NAND2_X1 U13486 ( .A1(n11865), .A2(n11864), .ZN(n15196) );
  OR2_X1 U13487 ( .A1(n11868), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U13488 ( .A1(n11869), .A2(n11911), .ZN(n21575) );
  INV_X1 U13489 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15205) );
  INV_X1 U13490 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11870) );
  OAI22_X1 U13491 ( .A1(n12163), .A2(n15205), .B1(n11975), .B2(n11870), .ZN(
        n11871) );
  AOI21_X1 U13492 ( .B1(n21575), .B2(n13339), .A(n11871), .ZN(n15197) );
  AOI22_X1 U13493 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U13494 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U13495 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U13496 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U13497 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11882) );
  AOI22_X1 U13498 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U13499 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U13500 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U13501 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U13502 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11881) );
  OR2_X1 U13503 ( .A1(n11882), .A2(n11881), .ZN(n11883) );
  AOI22_X1 U13504 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U13505 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U13506 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U13507 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11884) );
  NAND4_X1 U13508 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n11893) );
  AOI22_X1 U13509 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U13510 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U13511 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U13512 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U13513 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11892) );
  NOR2_X1 U13514 ( .A1(n11893), .A2(n11892), .ZN(n11898) );
  XNOR2_X1 U13515 ( .A(n11916), .B(n15278), .ZN(n15864) );
  NAND2_X1 U13516 ( .A1(n15864), .A2(n13339), .ZN(n11896) );
  AOI22_X1 U13517 ( .A1(n11788), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n13329), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11895) );
  OAI211_X1 U13518 ( .C1(n11898), .C2(n11897), .A(n11896), .B(n11895), .ZN(
        n15261) );
  INV_X1 U13519 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U13520 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13305), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U13521 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14448), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U13522 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U13523 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11900) );
  NAND4_X1 U13524 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11909) );
  AOI22_X1 U13525 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U13526 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11670), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U13527 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U13528 ( .A1(n11711), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U13529 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11908) );
  OR2_X1 U13530 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  NAND2_X1 U13531 ( .A1(n11942), .A2(n11910), .ZN(n11915) );
  XNOR2_X1 U13532 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11911), .ZN(
        n21584) );
  INV_X1 U13533 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11912) );
  OAI22_X1 U13534 ( .A1(n21584), .A2(n11753), .B1(n11975), .B2(n11912), .ZN(
        n11913) );
  INV_X1 U13535 ( .A(n11913), .ZN(n11914) );
  OAI211_X1 U13536 ( .C1(n12163), .C2(n15226), .A(n11915), .B(n11914), .ZN(
        n15223) );
  INV_X1 U13537 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15236) );
  XNOR2_X1 U13538 ( .A(n15236), .B(n11930), .ZN(n19964) );
  AOI22_X1 U13539 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U13540 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U13541 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U13542 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U13543 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11926) );
  AOI22_X1 U13544 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U13545 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U13546 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U13547 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U13548 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11925) );
  OR2_X1 U13549 ( .A1(n11926), .A2(n11925), .ZN(n11927) );
  AOI22_X1 U13550 ( .A1(n11942), .A2(n11927), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11929) );
  NAND2_X1 U13551 ( .A1(n11788), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11928) );
  OAI211_X1 U13552 ( .C1(n19964), .C2(n11753), .A(n11929), .B(n11928), .ZN(
        n15227) );
  XNOR2_X1 U13553 ( .A(n11960), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21588) );
  AOI22_X1 U13554 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U13555 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13556 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U13557 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U13558 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11940) );
  AOI22_X1 U13559 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U13560 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U13561 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U13562 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U13563 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  OR2_X1 U13564 ( .A1(n11940), .A2(n11939), .ZN(n11941) );
  AOI22_X1 U13565 ( .A1(n11942), .A2(n11941), .B1(n13329), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11944) );
  NAND2_X1 U13566 ( .A1(n11788), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11943) );
  OAI211_X1 U13567 ( .C1(n21588), .C2(n11753), .A(n11944), .B(n11943), .ZN(
        n15250) );
  AOI22_X1 U13568 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U13569 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U13570 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U13571 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11945) );
  NAND4_X1 U13572 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11954) );
  AOI22_X1 U13573 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U13574 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U13575 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U13576 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11949) );
  NAND4_X1 U13577 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11953) );
  NOR2_X1 U13578 ( .A1(n11954), .A2(n11953), .ZN(n11958) );
  NAND2_X1 U13579 ( .A1(n22008), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U13580 ( .A1(n11753), .A2(n11955), .ZN(n11956) );
  AOI21_X1 U13581 ( .B1(n12204), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11956), .ZN(
        n11957) );
  OAI21_X1 U13582 ( .B1(n13326), .B2(n11958), .A(n11957), .ZN(n11963) );
  OAI21_X1 U13583 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11961), .A(
        n11979), .ZN(n21605) );
  OR2_X1 U13584 ( .A1(n11753), .A2(n21605), .ZN(n11962) );
  NAND2_X1 U13585 ( .A1(n15249), .A2(n15288), .ZN(n15289) );
  AOI22_X1 U13586 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13587 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13588 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U13589 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11965) );
  NAND4_X1 U13590 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(
        n11974) );
  AOI22_X1 U13591 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13592 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U13593 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U13594 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U13595 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  OAI21_X1 U13596 ( .B1(n11974), .B2(n11973), .A(n12201), .ZN(n11978) );
  XNOR2_X1 U13597 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11979), .ZN(
        n15843) );
  OAI22_X1 U13598 ( .A1(n15843), .A2(n11753), .B1(n11975), .B2(n15612), .ZN(
        n11976) );
  AOI21_X1 U13599 ( .B1(n12204), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11976), .ZN(
        n11977) );
  OR2_X1 U13600 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U13601 ( .A1(n11981), .A2(n12012), .ZN(n21617) );
  AOI22_X1 U13602 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13603 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U13604 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U13605 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11982) );
  NAND4_X1 U13606 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11991) );
  AOI22_X1 U13607 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U13608 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U13609 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U13610 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U13611 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11990) );
  NOR2_X1 U13612 ( .A1(n11991), .A2(n11990), .ZN(n11994) );
  OAI21_X1 U13613 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21936), .A(
        n22008), .ZN(n11993) );
  NAND2_X1 U13614 ( .A1(n11788), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n11992) );
  OAI211_X1 U13615 ( .C1(n13326), .C2(n11994), .A(n11993), .B(n11992), .ZN(
        n11995) );
  OAI21_X1 U13616 ( .B1(n21617), .B2(n11753), .A(n11995), .ZN(n15652) );
  AOI22_X1 U13617 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U13618 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14448), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U13619 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U13620 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U13621 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12005) );
  AOI22_X1 U13622 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U13623 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U13624 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U13625 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U13626 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NOR2_X1 U13627 ( .A1(n12005), .A2(n12004), .ZN(n12009) );
  NAND2_X1 U13628 ( .A1(n22008), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U13629 ( .A1(n11753), .A2(n12006), .ZN(n12007) );
  AOI21_X1 U13630 ( .B1(n12204), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12007), .ZN(
        n12008) );
  OAI21_X1 U13631 ( .B1(n13326), .B2(n12009), .A(n12008), .ZN(n12011) );
  XNOR2_X1 U13632 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12012), .ZN(
        n15820) );
  NAND2_X1 U13633 ( .A1(n15820), .A2(n13339), .ZN(n12010) );
  OR2_X1 U13634 ( .A1(n12013), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U13635 ( .A1(n12014), .A2(n12048), .ZN(n19975) );
  INV_X1 U13636 ( .A(n19975), .ZN(n21630) );
  AOI22_X1 U13637 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U13638 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U13639 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U13640 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U13641 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12024) );
  AOI22_X1 U13642 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11582), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U13643 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13306), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U13644 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14448), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U13645 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11670), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U13646 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12023) );
  OR2_X1 U13647 ( .A1(n12024), .A2(n12023), .ZN(n12028) );
  INV_X1 U13648 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U13649 ( .A1(n22008), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12025) );
  OAI211_X1 U13650 ( .C1(n12163), .C2(n12026), .A(n11753), .B(n12025), .ZN(
        n12027) );
  AOI21_X1 U13651 ( .B1(n12201), .B2(n12028), .A(n12027), .ZN(n12029) );
  AOI21_X1 U13652 ( .B1(n21630), .B2(n13339), .A(n12029), .ZN(n15647) );
  AOI22_X1 U13653 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U13654 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U13655 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U13656 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12030) );
  NAND4_X1 U13657 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12040) );
  AOI22_X1 U13658 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U13659 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U13660 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13661 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U13662 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  NOR2_X1 U13663 ( .A1(n12040), .A2(n12039), .ZN(n12044) );
  NAND2_X1 U13664 ( .A1(n22008), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U13665 ( .A1(n11753), .A2(n12041), .ZN(n12042) );
  AOI21_X1 U13666 ( .B1(n12204), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12042), .ZN(
        n12043) );
  OAI21_X1 U13667 ( .B1(n13326), .B2(n12044), .A(n12043), .ZN(n12046) );
  XNOR2_X1 U13668 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12048), .ZN(
        n15586) );
  NAND2_X1 U13669 ( .A1(n13339), .A2(n15586), .ZN(n12045) );
  NAND2_X1 U13670 ( .A1(n12046), .A2(n12045), .ZN(n15583) );
  OR2_X1 U13671 ( .A1(n12049), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12050) );
  NAND2_X1 U13672 ( .A1(n12050), .A2(n12091), .ZN(n21643) );
  INV_X1 U13673 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13674 ( .A1(n11711), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U13675 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U13676 ( .A1(n13312), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13677 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12051) );
  NAND4_X1 U13678 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12061) );
  AOI22_X1 U13679 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U13680 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U13681 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U13682 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12056) );
  NAND4_X1 U13683 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n12060) );
  OAI21_X1 U13684 ( .B1(n12061), .B2(n12060), .A(n12201), .ZN(n12063) );
  AOI21_X1 U13685 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22008), .A(
        n13339), .ZN(n12062) );
  OAI211_X1 U13686 ( .C1(n12163), .C2(n12064), .A(n12063), .B(n12062), .ZN(
        n12065) );
  OAI21_X1 U13687 ( .B1(n21643), .B2(n11753), .A(n12065), .ZN(n15634) );
  AOI22_X1 U13688 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14448), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U13689 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U13690 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U13691 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U13692 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12075) );
  AOI22_X1 U13693 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U13694 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U13695 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13696 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U13697 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12074) );
  NOR2_X1 U13698 ( .A1(n12075), .A2(n12074), .ZN(n12097) );
  AOI22_X1 U13699 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13700 ( .A1(n11964), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U13701 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U13702 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U13703 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U13704 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U13705 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U13706 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13707 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U13708 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NOR2_X1 U13709 ( .A1(n12086), .A2(n12085), .ZN(n12098) );
  XOR2_X1 U13710 ( .A(n12097), .B(n12098), .Z(n12087) );
  NAND2_X1 U13711 ( .A1(n12201), .A2(n12087), .ZN(n12090) );
  INV_X1 U13712 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15803) );
  NOR2_X1 U13713 ( .A1(n15803), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12088) );
  AOI211_X1 U13714 ( .C1(n12204), .C2(P1_EAX_REG_23__SCAN_IN), .A(n13339), .B(
        n12088), .ZN(n12089) );
  XNOR2_X1 U13715 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12091), .ZN(
        n15807) );
  AOI22_X1 U13716 ( .A1(n12090), .A2(n12089), .B1(n13339), .B2(n15807), .ZN(
        n15571) );
  INV_X1 U13717 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12095) );
  INV_X1 U13718 ( .A(n12093), .ZN(n12094) );
  NAND2_X1 U13719 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  NAND2_X1 U13720 ( .A1(n12143), .A2(n12096), .ZN(n21658) );
  NOR2_X1 U13721 ( .A1(n12098), .A2(n12097), .ZN(n12124) );
  AOI22_X1 U13722 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13723 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13724 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13725 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U13726 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12108) );
  AOI22_X1 U13727 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U13728 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13729 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U13730 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U13731 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12107) );
  OR2_X1 U13732 ( .A1(n12108), .A2(n12107), .ZN(n12123) );
  XNOR2_X1 U13733 ( .A(n12124), .B(n12123), .ZN(n12111) );
  AOI21_X1 U13734 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n22008), .A(
        n13339), .ZN(n12110) );
  NAND2_X1 U13735 ( .A1(n11788), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12109) );
  OAI211_X1 U13736 ( .C1(n12111), .C2(n13326), .A(n12110), .B(n12109), .ZN(
        n12112) );
  OAI21_X1 U13737 ( .B1(n11753), .B2(n21658), .A(n12112), .ZN(n15627) );
  AOI22_X1 U13738 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13739 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U13740 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U13741 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U13742 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12122) );
  AOI22_X1 U13743 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U13744 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U13745 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U13746 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U13747 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12121) );
  NOR2_X1 U13748 ( .A1(n12122), .A2(n12121), .ZN(n12130) );
  NAND2_X1 U13749 ( .A1(n12124), .A2(n12123), .ZN(n12129) );
  XOR2_X1 U13750 ( .A(n12130), .B(n12129), .Z(n12125) );
  NAND2_X1 U13751 ( .A1(n12125), .A2(n12201), .ZN(n12128) );
  NOR2_X1 U13752 ( .A1(n15788), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12126) );
  AOI211_X1 U13753 ( .C1(n12204), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13339), .B(
        n12126), .ZN(n12127) );
  XNOR2_X1 U13754 ( .A(n12143), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15792) );
  AOI22_X1 U13755 ( .A1(n12128), .A2(n12127), .B1(n13339), .B2(n15792), .ZN(
        n15555) );
  NOR2_X1 U13756 ( .A1(n12130), .A2(n12129), .ZN(n12160) );
  AOI22_X1 U13757 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13758 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U13759 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U13760 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12131) );
  NAND4_X1 U13761 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12140) );
  AOI22_X1 U13762 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U13763 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U13764 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U13765 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U13766 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12139) );
  OR2_X1 U13767 ( .A1(n12140), .A2(n12139), .ZN(n12159) );
  XNOR2_X1 U13768 ( .A(n12160), .B(n12159), .ZN(n12141) );
  NOR2_X1 U13769 ( .A1(n12141), .A2(n13326), .ZN(n12148) );
  INV_X1 U13770 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21834) );
  NOR2_X1 U13771 ( .A1(n21936), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12142) );
  OAI22_X1 U13772 ( .A1(n12163), .A2(n21834), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12142), .ZN(n12147) );
  INV_X1 U13773 ( .A(n12144), .ZN(n12145) );
  INV_X1 U13774 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15547) );
  NAND2_X1 U13775 ( .A1(n12145), .A2(n15547), .ZN(n12146) );
  NAND2_X1 U13776 ( .A1(n12167), .A2(n12146), .ZN(n15782) );
  OAI22_X1 U13777 ( .A1(n12148), .A2(n12147), .B1(n11753), .B2(n15782), .ZN(
        n15542) );
  XNOR2_X1 U13778 ( .A(n12167), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15774) );
  AOI22_X1 U13779 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13306), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13780 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11670), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U13781 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U13782 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12055), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12149) );
  NAND4_X1 U13783 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12158) );
  AOI22_X1 U13784 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13313), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U13785 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13305), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U13786 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13787 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U13788 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NOR2_X1 U13789 ( .A1(n12158), .A2(n12157), .ZN(n12173) );
  NAND2_X1 U13790 ( .A1(n12160), .A2(n12159), .ZN(n12172) );
  XOR2_X1 U13791 ( .A(n12173), .B(n12172), .Z(n12165) );
  INV_X1 U13792 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U13793 ( .A1(n22008), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12161) );
  OAI211_X1 U13794 ( .C1(n12163), .C2(n12162), .A(n11753), .B(n12161), .ZN(
        n12164) );
  AOI21_X1 U13795 ( .B1(n12165), .B2(n12201), .A(n12164), .ZN(n12166) );
  AOI21_X1 U13796 ( .B1(n13339), .B2(n15774), .A(n12166), .ZN(n15528) );
  INV_X1 U13797 ( .A(n12167), .ZN(n12168) );
  INV_X1 U13798 ( .A(n12169), .ZN(n12170) );
  INV_X1 U13799 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15517) );
  NAND2_X1 U13800 ( .A1(n12170), .A2(n15517), .ZN(n12171) );
  NAND2_X1 U13801 ( .A1(n13303), .A2(n12171), .ZN(n15765) );
  NOR2_X1 U13802 ( .A1(n12173), .A2(n12172), .ZN(n12200) );
  AOI22_X1 U13803 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13307), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U13804 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U13805 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U13806 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U13807 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U13808 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U13809 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U13810 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U13811 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U13812 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  OR2_X1 U13813 ( .A1(n12184), .A2(n12183), .ZN(n12199) );
  XNOR2_X1 U13814 ( .A(n12200), .B(n12199), .ZN(n12187) );
  AOI21_X1 U13815 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n22008), .A(
        n13339), .ZN(n12186) );
  NAND2_X1 U13816 ( .A1(n11788), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12185) );
  OAI211_X1 U13817 ( .C1(n12187), .C2(n13326), .A(n12186), .B(n12185), .ZN(
        n12188) );
  OAI21_X1 U13818 ( .B1(n11753), .B2(n15765), .A(n12188), .ZN(n14049) );
  AOI22_X1 U13819 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11589), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U13820 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13306), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U13821 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U13822 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12189) );
  NAND4_X1 U13823 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12198) );
  AOI22_X1 U13824 ( .A1(n13305), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U13825 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U13826 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11964), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U13827 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U13828 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12197) );
  NOR2_X1 U13829 ( .A1(n12198), .A2(n12197), .ZN(n13321) );
  NAND2_X1 U13830 ( .A1(n12200), .A2(n12199), .ZN(n13320) );
  XOR2_X1 U13831 ( .A(n13321), .B(n13320), .Z(n12202) );
  NAND2_X1 U13832 ( .A1(n12202), .A2(n12201), .ZN(n12206) );
  INV_X1 U13833 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15747) );
  NOR2_X1 U13834 ( .A1(n15747), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12203) );
  AOI211_X1 U13835 ( .C1(n12204), .C2(P1_EAX_REG_29__SCAN_IN), .A(n13339), .B(
        n12203), .ZN(n12205) );
  XNOR2_X1 U13836 ( .A(n13303), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15746) );
  AOI22_X1 U13837 ( .A1(n12206), .A2(n12205), .B1(n13339), .B2(n15746), .ZN(
        n12208) );
  NAND2_X1 U13838 ( .A1(n12210), .A2(n11017), .ZN(n14254) );
  NAND2_X1 U13839 ( .A1(n21965), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12212) );
  NAND2_X1 U13840 ( .A1(n11411), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U13841 ( .A1(n12212), .A2(n12211), .ZN(n12228) );
  NAND2_X1 U13842 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21975), .ZN(
        n12242) );
  NAND2_X1 U13843 ( .A1(n12213), .A2(n12212), .ZN(n12225) );
  NAND2_X1 U13844 ( .A1(n21922), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12215) );
  NAND2_X1 U13845 ( .A1(n11015), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12214) );
  NAND2_X1 U13846 ( .A1(n12225), .A2(n12226), .ZN(n12216) );
  NAND2_X1 U13847 ( .A1(n12216), .A2(n12215), .ZN(n12219) );
  NAND2_X1 U13848 ( .A1(n12219), .A2(n12220), .ZN(n12233) );
  NAND2_X1 U13849 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14465), .ZN(
        n12234) );
  NAND2_X1 U13850 ( .A1(n12233), .A2(n12234), .ZN(n12218) );
  NAND2_X1 U13851 ( .A1(n12217), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12230) );
  NAND2_X1 U13852 ( .A1(n12218), .A2(n12230), .ZN(n12224) );
  INV_X1 U13853 ( .A(n12219), .ZN(n12222) );
  NAND2_X1 U13854 ( .A1(n12230), .A2(n12220), .ZN(n12221) );
  NAND2_X1 U13855 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  NAND2_X1 U13856 ( .A1(n12224), .A2(n12223), .ZN(n12240) );
  XOR2_X1 U13857 ( .A(n12226), .B(n12225), .Z(n12257) );
  INV_X1 U13858 ( .A(n12242), .ZN(n12227) );
  XNOR2_X1 U13859 ( .A(n12228), .B(n12227), .ZN(n12249) );
  NAND2_X1 U13860 ( .A1(n12257), .A2(n12249), .ZN(n12229) );
  OR2_X1 U13861 ( .A1(n12240), .A2(n12229), .ZN(n12236) );
  NAND2_X1 U13862 ( .A1(n16841), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12231) );
  AND2_X1 U13863 ( .A1(n12231), .A2(n12230), .ZN(n12232) );
  NAND2_X1 U13864 ( .A1(n12233), .A2(n12232), .ZN(n12235) );
  NAND2_X1 U13865 ( .A1(n12236), .A2(n12239), .ZN(n14120) );
  NAND2_X1 U13866 ( .A1(n11549), .A2(n21716), .ZN(n12275) );
  INV_X1 U13867 ( .A(n12239), .ZN(n12237) );
  NOR2_X1 U13868 ( .A1(n12241), .A2(n12264), .ZN(n12266) );
  NAND2_X1 U13869 ( .A1(n12248), .A2(n12257), .ZN(n12255) );
  INV_X1 U13870 ( .A(n12255), .ZN(n12262) );
  AOI21_X1 U13871 ( .B1(n11549), .B2(n12238), .A(n14715), .ZN(n12256) );
  INV_X1 U13872 ( .A(n12256), .ZN(n12261) );
  OAI22_X1 U13873 ( .A1(n21683), .A2(n12238), .B1(n12258), .B2(n12249), .ZN(
        n12247) );
  NOR3_X1 U13874 ( .A1(n13348), .A2(n12249), .A3(n12247), .ZN(n12254) );
  INV_X1 U13875 ( .A(n13583), .ZN(n14224) );
  OAI21_X1 U13876 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21975), .A(
        n12242), .ZN(n12244) );
  INV_X1 U13877 ( .A(n12244), .ZN(n12243) );
  OAI211_X1 U13878 ( .C1(n11018), .C2(n14224), .A(n12256), .B(n12243), .ZN(
        n12246) );
  INV_X1 U13879 ( .A(n12248), .ZN(n12250) );
  OAI21_X1 U13880 ( .B1(n12250), .B2(n12244), .A(n12263), .ZN(n12245) );
  NAND2_X1 U13881 ( .A1(n12246), .A2(n12245), .ZN(n12253) );
  AOI21_X1 U13882 ( .B1(n12248), .B2(n13348), .A(n12247), .ZN(n12252) );
  AOI21_X1 U13883 ( .B1(n12250), .B2(n13521), .A(n12249), .ZN(n12251) );
  OAI22_X1 U13884 ( .A1(n12254), .A2(n12253), .B1(n12252), .B2(n12251), .ZN(
        n12260) );
  OAI211_X1 U13885 ( .C1(n12258), .C2(n12257), .A(n12256), .B(n12255), .ZN(
        n12259) );
  AOI22_X1 U13886 ( .A1(n12262), .A2(n12261), .B1(n12260), .B2(n12259), .ZN(
        n12265) );
  OAI22_X1 U13887 ( .A1(n12266), .A2(n12265), .B1(n12264), .B2(n12263), .ZN(
        n12267) );
  AOI21_X1 U13888 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21683), .A(
        n12267), .ZN(n12268) );
  INV_X1 U13889 ( .A(n12268), .ZN(n12269) );
  AND2_X1 U13890 ( .A1(n12273), .A2(n14715), .ZN(n12274) );
  NAND2_X1 U13891 ( .A1(n16033), .A2(n12274), .ZN(n14121) );
  OAI22_X1 U13892 ( .A1(n14117), .A2(n12275), .B1(n14310), .B2(n14121), .ZN(
        n14260) );
  INV_X1 U13893 ( .A(n12276), .ZN(n12277) );
  INV_X1 U13894 ( .A(n14578), .ZN(n13471) );
  NAND4_X1 U13895 ( .A1(n12277), .A2(n13471), .A3(n11031), .A4(n14570), .ZN(
        n13465) );
  NAND2_X1 U13896 ( .A1(n13348), .A2(n21716), .ZN(n14208) );
  NOR2_X1 U13897 ( .A1(n14310), .A2(n14208), .ZN(n12279) );
  NAND2_X1 U13898 ( .A1(n12278), .A2(n12279), .ZN(n14249) );
  OAI21_X1 U13899 ( .B1(n13465), .B2(n15447), .A(n14249), .ZN(n12280) );
  NAND2_X1 U13900 ( .A1(n12282), .A2(n14578), .ZN(n14510) );
  NOR2_X1 U13901 ( .A1(n15508), .A2(n15725), .ZN(n12302) );
  NOR2_X1 U13902 ( .A1(n15720), .A2(n14303), .ZN(n12298) );
  NOR4_X1 U13903 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12286) );
  NOR4_X1 U13904 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12285) );
  NOR4_X1 U13905 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12284) );
  NOR4_X1 U13906 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12283) );
  AND4_X1 U13907 ( .A1(n12286), .A2(n12285), .A3(n12284), .A4(n12283), .ZN(
        n12291) );
  NOR4_X1 U13908 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12289) );
  NOR4_X1 U13909 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12288) );
  NOR4_X1 U13910 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12287) );
  INV_X1 U13911 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19821) );
  AND4_X1 U13912 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n19821), .ZN(
        n12290) );
  NAND2_X1 U13913 ( .A1(n12291), .A2(n12290), .ZN(n12292) );
  INV_X1 U13914 ( .A(DATAI_29_), .ZN(n12297) );
  NOR2_X1 U13915 ( .A1(n13471), .A2(n12238), .ZN(n12293) );
  INV_X2 U13916 ( .A(n14544), .ZN(n15202) );
  INV_X1 U13917 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20014) );
  OR2_X1 U13918 ( .A1(n15202), .A2(n20014), .ZN(n12295) );
  NAND2_X1 U13919 ( .A1(n15202), .A2(DATAI_13_), .ZN(n12294) );
  NAND2_X1 U13920 ( .A1(n12295), .A2(n12294), .ZN(n21848) );
  AOI22_X1 U13921 ( .A1(n15722), .A2(n21848), .B1(n15720), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n12296) );
  OAI21_X1 U13922 ( .B1(n15724), .B2(n12297), .A(n12296), .ZN(n12300) );
  AND2_X1 U13923 ( .A1(n15729), .A2(BUF1_REG_29__SCAN_IN), .ZN(n12299) );
  OR2_X1 U13924 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  INV_X1 U13925 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12305) );
  AND2_X2 U13926 ( .A1(n12305), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14769) );
  AND2_X4 U13927 ( .A1(n14769), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12405) );
  AOI22_X1 U13928 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10981), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12308) );
  AND2_X4 U13929 ( .A1(n12539), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12406) );
  AOI22_X1 U13930 ( .A1(n11000), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12307) );
  AND2_X4 U13931 ( .A1(n14768), .A2(n14798), .ZN(n12529) );
  AOI22_X1 U13932 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12306) );
  NAND4_X1 U13933 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12317) );
  AOI22_X1 U13934 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U13935 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10979), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U13936 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12312) );
  NAND4_X1 U13937 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12316) );
  NAND2_X1 U13938 ( .A1(n12317), .A2(n12316), .ZN(n12365) );
  AOI22_X1 U13939 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U13940 ( .A1(n11023), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U13941 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U13942 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10979), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12318) );
  NAND4_X1 U13943 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n12322) );
  AOI22_X1 U13944 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U13945 ( .A1(n11000), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U13946 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12323) );
  NAND4_X1 U13947 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        n12327) );
  NAND2_X4 U13948 ( .A1(n12329), .A2(n12328), .ZN(n18291) );
  INV_X1 U13949 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19572) );
  NOR2_X1 U13950 ( .A1(n12750), .A2(n19572), .ZN(n12492) );
  AOI22_X1 U13951 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U13952 ( .A1(n11023), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U13953 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U13954 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U13955 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12336) );
  AND2_X1 U13956 ( .A1(n12336), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12340) );
  AOI22_X1 U13957 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10980), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U13958 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U13959 ( .A1(n11024), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U13960 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12341) );
  NAND2_X2 U13961 ( .A1(n12342), .A2(n12341), .ZN(n12419) );
  AOI22_X1 U13962 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U13963 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U13964 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U13965 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  AOI22_X1 U13966 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U13967 ( .A1(n12405), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U13968 ( .A1(n11000), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U13969 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  NAND2_X2 U13970 ( .A1(n12365), .A2(n12394), .ZN(n12428) );
  AOI22_X1 U13971 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U13972 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10987), .B1(
        n10980), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U13974 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12532), .B1(
        n12530), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12353) );
  NAND4_X1 U13975 ( .A1(n12356), .A2(n12355), .A3(n12354), .A4(n12353), .ZN(
        n12357) );
  NAND2_X1 U13976 ( .A1(n12357), .A2(n12373), .ZN(n12364) );
  AOI22_X1 U13977 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U13978 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U13979 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12359) );
  NAND4_X1 U13980 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  NAND2_X1 U13981 ( .A1(n12362), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12363) );
  INV_X2 U13982 ( .A(n12365), .ZN(n12422) );
  NAND2_X1 U13983 ( .A1(n13964), .A2(n12428), .ZN(n12366) );
  NAND2_X1 U13984 ( .A1(n12366), .A2(n12419), .ZN(n13970) );
  NAND2_X1 U13985 ( .A1(n12367), .A2(n13970), .ZN(n12432) );
  INV_X1 U13986 ( .A(n12432), .ZN(n12393) );
  AOI22_X1 U13987 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10980), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U13988 ( .A1(n11000), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U13989 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U13990 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12374) );
  NAND2_X1 U13991 ( .A1(n12374), .A2(n12373), .ZN(n12381) );
  AOI22_X1 U13992 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U13993 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U13994 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U13995 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U13996 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12379) );
  NAND2_X1 U13997 ( .A1(n12379), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12380) );
  AOI22_X1 U13998 ( .A1(n11023), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U13999 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U14000 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12382) );
  NAND4_X1 U14001 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12391) );
  AOI22_X1 U14002 ( .A1(n11000), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U14003 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U14004 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12386) );
  NAND4_X1 U14005 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12390) );
  MUX2_X2 U14006 ( .A(n12391), .B(n12390), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12440) );
  AND2_X1 U14007 ( .A1(n12394), .A2(n12425), .ZN(n12396) );
  NAND2_X1 U14008 ( .A1(n12419), .A2(n12422), .ZN(n12416) );
  INV_X1 U14009 ( .A(n12416), .ZN(n12426) );
  NAND3_X1 U14010 ( .A1(n13955), .A2(n12397), .A3(n18291), .ZN(n12398) );
  AOI22_X1 U14011 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U14012 ( .A1(n11001), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U14013 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U14014 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U14015 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12403) );
  NAND2_X1 U14016 ( .A1(n12403), .A2(n12373), .ZN(n12414) );
  AOI22_X1 U14017 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U14018 ( .A1(n11024), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12406), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U14019 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U14020 ( .A1(n12530), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12532), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U14021 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12412) );
  NAND2_X1 U14022 ( .A1(n12412), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12413) );
  NAND2_X2 U14023 ( .A1(n12414), .A2(n12413), .ZN(n14009) );
  INV_X1 U14024 ( .A(n18290), .ZN(n12445) );
  NAND2_X1 U14025 ( .A1(n14006), .A2(n12445), .ZN(n12431) );
  NAND2_X1 U14026 ( .A1(n12415), .A2(n12425), .ZN(n12435) );
  NAND2_X1 U14027 ( .A1(n12435), .A2(n12416), .ZN(n12418) );
  NAND2_X1 U14028 ( .A1(n12428), .A2(n12440), .ZN(n12417) );
  AND4_X1 U14029 ( .A1(n13975), .A2(n12419), .A3(n12394), .A4(n12425), .ZN(
        n12420) );
  AND2_X2 U14030 ( .A1(n12421), .A2(n12420), .ZN(n14834) );
  INV_X1 U14031 ( .A(n14834), .ZN(n16764) );
  AOI21_X1 U14032 ( .B1(n12422), .B2(n12394), .A(n13975), .ZN(n12423) );
  NAND2_X1 U14033 ( .A1(n12421), .A2(n12423), .ZN(n12424) );
  NAND2_X1 U14034 ( .A1(n16764), .A2(n12424), .ZN(n14010) );
  NOR2_X1 U14035 ( .A1(n12394), .A2(n12425), .ZN(n12427) );
  AND2_X1 U14036 ( .A1(n12428), .A2(n19574), .ZN(n12450) );
  NAND3_X1 U14037 ( .A1(n14010), .A2(n14018), .A3(n12450), .ZN(n12429) );
  NOR2_X1 U14038 ( .A1(n14009), .A2(n18286), .ZN(n18293) );
  NAND2_X1 U14039 ( .A1(n12429), .A2(n18293), .ZN(n12430) );
  NAND2_X2 U14040 ( .A1(n12454), .A2(n11398), .ZN(n12512) );
  NAND2_X1 U14041 ( .A1(n12512), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12444) );
  INV_X1 U14042 ( .A(n12435), .ZN(n12436) );
  NAND2_X1 U14043 ( .A1(n14096), .A2(n12436), .ZN(n12439) );
  NAND3_X1 U14044 ( .A1(n12459), .A2(n19353), .A3(n13269), .ZN(n12437) );
  NOR2_X2 U14045 ( .A1(n12439), .A2(n12438), .ZN(n12894) );
  NAND2_X1 U14046 ( .A1(n12894), .A2(n12441), .ZN(n12460) );
  INV_X1 U14047 ( .A(n12441), .ZN(n13969) );
  NOR2_X1 U14048 ( .A1(n13969), .A2(n14822), .ZN(n12442) );
  NAND2_X1 U14049 ( .A1(n12909), .A2(n12442), .ZN(n14408) );
  NAND2_X1 U14050 ( .A1(n12460), .A2(n14408), .ZN(n14789) );
  INV_X2 U14051 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U14052 ( .A1(n18286), .A2(n14093), .ZN(n18620) );
  AOI22_X1 U14053 ( .A1(n14789), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n13261), .ZN(n12443) );
  NAND2_X1 U14054 ( .A1(n12444), .A2(n12443), .ZN(n12498) );
  NOR2_X2 U14055 ( .A1(n14765), .A2(n12446), .ZN(n12509) );
  NOR2_X2 U14056 ( .A1(n12446), .A2(n13969), .ZN(n12447) );
  NAND2_X4 U14057 ( .A1(n12447), .A2(n12909), .ZN(n13228) );
  INV_X1 U14058 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14411) );
  NAND2_X1 U14059 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12448) );
  AOI21_X1 U14060 ( .B1(n12509), .B2(P2_REIP_REG_0__SCAN_IN), .A(n12449), .ZN(
        n12455) );
  INV_X1 U14061 ( .A(n12450), .ZN(n12451) );
  AND3_X1 U14062 ( .A1(n12455), .A2(n12454), .A3(n12453), .ZN(n12463) );
  INV_X1 U14063 ( .A(n12904), .ZN(n12458) );
  NAND2_X1 U14064 ( .A1(n12422), .A2(n12425), .ZN(n13093) );
  INV_X1 U14065 ( .A(n13093), .ZN(n12922) );
  NAND2_X1 U14066 ( .A1(n12922), .A2(n13269), .ZN(n12457) );
  NAND2_X1 U14067 ( .A1(n12458), .A2(n11060), .ZN(n12464) );
  NAND2_X1 U14068 ( .A1(n12464), .A2(n19574), .ZN(n12461) );
  NAND2_X1 U14069 ( .A1(n13995), .A2(n11397), .ZN(n12462) );
  NAND2_X1 U14070 ( .A1(n12463), .A2(n12462), .ZN(n12499) );
  NAND2_X1 U14071 ( .A1(n12498), .A2(n12499), .ZN(n12468) );
  BUF_X2 U14072 ( .A(n12468), .Z(n12501) );
  NAND2_X1 U14073 ( .A1(n12512), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12467) );
  AND2_X1 U14074 ( .A1(n13261), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12465) );
  AOI21_X1 U14075 ( .B1(n14806), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12465), 
        .ZN(n12466) );
  INV_X1 U14076 ( .A(n12468), .ZN(n12470) );
  NAND2_X1 U14077 ( .A1(n12470), .A2(n12469), .ZN(n12474) );
  INV_X1 U14078 ( .A(n12507), .ZN(n13142) );
  INV_X1 U14079 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12472) );
  INV_X2 U14080 ( .A(n13228), .ZN(n13159) );
  AOI22_X1 U14081 ( .A1(n13159), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12471) );
  OAI21_X1 U14082 ( .B1(n13143), .B2(n12472), .A(n12471), .ZN(n12473) );
  INV_X1 U14083 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12475) );
  INV_X1 U14084 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14161) );
  OAI22_X1 U14085 ( .A1(n13228), .A2(n12475), .B1(n14093), .B2(n14161), .ZN(
        n12476) );
  AOI21_X1 U14086 ( .B1(n12509), .B2(P2_REIP_REG_2__SCAN_IN), .A(n12476), .ZN(
        n12477) );
  NAND2_X1 U14087 ( .A1(n12512), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12479) );
  AOI21_X1 U14088 ( .B1(n18286), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12478) );
  NAND2_X1 U14089 ( .A1(n12479), .A2(n12478), .ZN(n12480) );
  NAND2_X1 U14090 ( .A1(n12481), .A2(n12480), .ZN(n12516) );
  INV_X1 U14091 ( .A(n12480), .ZN(n12483) );
  NAND2_X1 U14092 ( .A1(n12484), .A2(n12485), .ZN(n12487) );
  INV_X1 U14093 ( .A(n12485), .ZN(n12486) );
  NAND2_X2 U14094 ( .A1(n12487), .A2(n13149), .ZN(n13623) );
  NAND2_X1 U14095 ( .A1(n13623), .A2(n12502), .ZN(n12490) );
  NAND2_X1 U14096 ( .A1(n12422), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12488) );
  NAND2_X1 U14097 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19272) );
  XNOR2_X1 U14098 ( .A(n19272), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19163) );
  AOI22_X1 U14099 ( .A1(n12521), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19321), .B2(n19163), .ZN(n12489) );
  NAND2_X1 U14100 ( .A1(n12490), .A2(n12489), .ZN(n12491) );
  INV_X1 U14101 ( .A(n12501), .ZN(n12495) );
  NAND2_X1 U14102 ( .A1(n13610), .A2(n12502), .ZN(n12497) );
  NAND2_X1 U14103 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17147), .ZN(
        n19288) );
  NAND2_X1 U14104 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19302), .ZN(
        n19305) );
  NAND2_X1 U14105 ( .A1(n19288), .A2(n19305), .ZN(n17044) );
  AND2_X1 U14106 ( .A1(n19321), .A2(n17044), .ZN(n19289) );
  AOI21_X1 U14107 ( .B1(n12521), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19289), .ZN(n12496) );
  NOR2_X1 U14108 ( .A1(n19307), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12503) );
  AOI21_X1 U14109 ( .B1(n12521), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12503), .ZN(n12504) );
  OAI22_X1 U14110 ( .A1(n14405), .A2(n14404), .B1(n12505), .B2(n14373), .ZN(
        n14413) );
  INV_X1 U14111 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13271) );
  INV_X1 U14112 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14920) );
  OAI22_X1 U14113 ( .A1(n13228), .A2(n13271), .B1(n14093), .B2(n14920), .ZN(
        n12508) );
  AOI21_X1 U14114 ( .B1(n12509), .B2(P2_REIP_REG_3__SCAN_IN), .A(n12508), .ZN(
        n12510) );
  NAND2_X1 U14115 ( .A1(n12512), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12514) );
  NAND2_X1 U14116 ( .A1(n13261), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12513) );
  NAND2_X1 U14117 ( .A1(n12514), .A2(n12513), .ZN(n13152) );
  INV_X1 U14118 ( .A(n12518), .ZN(n12515) );
  OAI21_X1 U14119 ( .B1(n19272), .B2(n17156), .A(n19175), .ZN(n12520) );
  INV_X1 U14120 ( .A(n19272), .ZN(n12519) );
  NOR2_X1 U14121 ( .A1(n17156), .A2(n19175), .ZN(n19149) );
  NAND2_X1 U14122 ( .A1(n12519), .A2(n19149), .ZN(n19134) );
  AND3_X1 U14123 ( .A1(n12520), .A2(n19134), .A3(n19321), .ZN(n19161) );
  AOI21_X1 U14124 ( .B1(n12521), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19161), .ZN(n12522) );
  NOR2_X1 U14125 ( .A1(n12750), .A2(n19531), .ZN(n12523) );
  NAND2_X1 U14126 ( .A1(n12524), .A2(n12523), .ZN(n12527) );
  NAND2_X1 U14127 ( .A1(n14418), .A2(n14419), .ZN(n14417) );
  NAND2_X1 U14128 ( .A1(n12422), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12526) );
  AND2_X1 U14129 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  INV_X1 U14130 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19493) );
  NOR2_X1 U14131 ( .A1(n12750), .A2(n19493), .ZN(n14495) );
  INV_X1 U14132 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19395) );
  INV_X1 U14133 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14610) );
  AND2_X2 U14134 ( .A1(n10989), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12848) );
  AND2_X2 U14135 ( .A1(n10985), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12930) );
  AOI22_X1 U14136 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12930), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U14137 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12536) );
  AND2_X2 U14138 ( .A1(n10987), .A2(n12373), .ZN(n13028) );
  AOI22_X1 U14139 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12535) );
  AND2_X2 U14140 ( .A1(n12531), .A2(n12373), .ZN(n13033) );
  AOI22_X1 U14141 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12534) );
  NAND4_X1 U14142 ( .A1(n12537), .A2(n12536), .A3(n12535), .A4(n12534), .ZN(
        n12545) );
  AND2_X1 U14143 ( .A1(n12406), .A2(n12373), .ZN(n12648) );
  AOI22_X1 U14144 ( .A1(n12648), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12543) );
  AND2_X2 U14145 ( .A1(n12531), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12637) );
  AOI22_X1 U14146 ( .A1(n12637), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12542) );
  AND2_X1 U14147 ( .A1(n12711), .A2(n12538), .ZN(n12550) );
  AOI22_X1 U14148 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12541) );
  AND2_X1 U14149 ( .A1(n12539), .A2(n12711), .ZN(n12552) );
  AOI22_X1 U14150 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12540) );
  NAND4_X1 U14151 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12544) );
  AOI22_X1 U14152 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U14153 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U14154 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U14155 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U14156 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12558) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U14158 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U14159 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U14160 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12553) );
  NAND4_X1 U14161 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12557) );
  NAND2_X1 U14162 ( .A1(n14695), .A2(n14697), .ZN(n14696) );
  AOI22_X1 U14163 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U14164 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12562) );
  AOI22_X1 U14165 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U14166 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12700), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12560) );
  NAND4_X1 U14167 ( .A1(n12563), .A2(n12562), .A3(n12561), .A4(n12560), .ZN(
        n12570) );
  AOI22_X1 U14168 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U14169 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n14812), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U14170 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U14171 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12565) );
  NAND4_X1 U14172 ( .A1(n12568), .A2(n12567), .A3(n12566), .A4(n12565), .ZN(
        n12569) );
  AOI22_X1 U14173 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U14174 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U14175 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12572) );
  NAND4_X1 U14177 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12581) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U14179 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U14180 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U14181 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12576) );
  NAND4_X1 U14182 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12580) );
  AOI22_X1 U14183 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12930), .B1(
        n12848), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U14184 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13028), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U14185 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U14186 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U14187 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12591) );
  AOI22_X1 U14188 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U14189 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U14190 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U14191 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U14192 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12590) );
  NOR2_X1 U14193 ( .A1(n12591), .A2(n12590), .ZN(n13049) );
  AOI22_X1 U14194 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U14195 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U14196 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U14197 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U14198 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12602) );
  AOI22_X1 U14199 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U14200 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U14201 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U14202 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12597) );
  NAND4_X1 U14203 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12601) );
  AOI22_X1 U14204 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U14205 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U14206 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U14207 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12603) );
  NAND4_X1 U14208 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12612) );
  AOI22_X1 U14209 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U14210 ( .A1(n12637), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U14211 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U14212 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12607) );
  NAND4_X1 U14213 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n12611) );
  AOI22_X1 U14214 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U14215 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U14216 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14217 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12613) );
  NAND4_X1 U14218 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12622) );
  AOI22_X1 U14219 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U14220 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U14221 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U14222 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U14223 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  AOI22_X1 U14224 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U14225 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U14226 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U14227 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12623) );
  NAND4_X1 U14228 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n12632) );
  AOI22_X1 U14229 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14230 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U14231 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U14232 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12627) );
  NAND4_X1 U14233 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12631) );
  NOR2_X1 U14234 ( .A1(n12632), .A2(n12631), .ZN(n15207) );
  AOI22_X1 U14235 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U14236 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U14237 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U14238 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12633) );
  NAND4_X1 U14239 ( .A1(n12636), .A2(n12635), .A3(n12634), .A4(n12633), .ZN(
        n12643) );
  AOI22_X1 U14240 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U14241 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U14242 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U14243 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12638) );
  NAND4_X1 U14244 ( .A1(n12641), .A2(n12640), .A3(n12639), .A4(n12638), .ZN(
        n12642) );
  OR2_X1 U14245 ( .A1(n12643), .A2(n12642), .ZN(n15212) );
  AOI22_X1 U14246 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14247 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14248 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U14249 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12644) );
  NAND4_X1 U14250 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12654) );
  AOI22_X1 U14251 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U14252 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U14253 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U14254 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12649) );
  NAND4_X1 U14255 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n12653) );
  NOR2_X1 U14256 ( .A1(n12654), .A2(n12653), .ZN(n16168) );
  AOI22_X1 U14257 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n12675), .ZN(n12658) );
  AOI22_X1 U14258 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U14259 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U14260 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n12592), .ZN(n12655) );
  NAND4_X1 U14261 ( .A1(n12658), .A2(n12657), .A3(n12656), .A4(n12655), .ZN(
        n12664) );
  AOI22_X1 U14262 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U14263 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U14264 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U14265 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n12552), .ZN(n12659) );
  NAND4_X1 U14266 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n12659), .ZN(
        n12663) );
  OR2_X1 U14267 ( .A1(n12664), .A2(n12663), .ZN(n16159) );
  AOI22_X1 U14268 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U14269 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U14270 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U14271 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n12592), .ZN(n12665) );
  NAND4_X1 U14272 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12674) );
  AOI22_X1 U14273 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U14274 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U14275 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U14276 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n12552), .ZN(n12669) );
  NAND4_X1 U14277 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  NOR2_X1 U14278 ( .A1(n12674), .A2(n12673), .ZN(n16155) );
  AOI22_X1 U14279 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12683) );
  INV_X1 U14280 ( .A(n12848), .ZN(n12678) );
  INV_X1 U14281 ( .A(n12675), .ZN(n12677) );
  INV_X1 U14282 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12676) );
  OAI22_X1 U14283 ( .A1(n12678), .A2(n14610), .B1(n12677), .B2(n12676), .ZN(
        n12679) );
  INV_X1 U14284 ( .A(n12679), .ZN(n12682) );
  AOI22_X1 U14285 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U14286 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U14287 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12689) );
  AOI22_X1 U14288 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U14289 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U14290 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U14291 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12684) );
  NAND4_X1 U14292 ( .A1(n12687), .A2(n12686), .A3(n12685), .A4(n12684), .ZN(
        n12688) );
  OR2_X1 U14293 ( .A1(n12689), .A2(n12688), .ZN(n16150) );
  AOI22_X1 U14294 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U14295 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U14296 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U14297 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U14298 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12699) );
  AOI22_X1 U14299 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U14300 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U14301 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U14302 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12694) );
  NAND4_X1 U14303 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12698) );
  AOI22_X1 U14304 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U14305 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U14306 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U14307 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12701) );
  NAND4_X1 U14308 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12710) );
  AOI22_X1 U14309 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U14310 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12637), .B1(
        n13033), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U14311 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U14312 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12705) );
  NAND4_X1 U14313 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n12705), .ZN(
        n12709) );
  NOR2_X1 U14314 ( .A1(n12710), .A2(n12709), .ZN(n12730) );
  AOI22_X1 U14315 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11023), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U14316 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U14317 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12718) );
  INV_X1 U14318 ( .A(n12406), .ZN(n15483) );
  INV_X1 U14319 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U14320 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12714) );
  INV_X1 U14321 ( .A(n12711), .ZN(n12713) );
  NAND2_X1 U14322 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12712) );
  NAND2_X1 U14323 ( .A1(n12713), .A2(n12712), .ZN(n15482) );
  OAI211_X1 U14324 ( .C1(n15483), .C2(n12715), .A(n12714), .B(n15482), .ZN(
        n12716) );
  INV_X1 U14325 ( .A(n12716), .ZN(n12717) );
  NAND4_X1 U14326 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        n12729) );
  AOI22_X1 U14327 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11000), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U14328 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U14329 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12725) );
  INV_X1 U14330 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U14331 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12721) );
  INV_X1 U14332 ( .A(n15482), .ZN(n12819) );
  OAI211_X1 U14333 ( .C1(n15483), .C2(n12722), .A(n12721), .B(n12819), .ZN(
        n12723) );
  INV_X1 U14334 ( .A(n12723), .ZN(n12724) );
  NAND4_X1 U14335 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12728) );
  NAND2_X1 U14336 ( .A1(n12729), .A2(n12728), .ZN(n12731) );
  XNOR2_X1 U14337 ( .A(n12730), .B(n12731), .ZN(n16139) );
  INV_X1 U14338 ( .A(n12730), .ZN(n12733) );
  INV_X1 U14339 ( .A(n12731), .ZN(n12732) );
  NAND2_X1 U14340 ( .A1(n12733), .A2(n12732), .ZN(n12751) );
  AOI22_X1 U14341 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U14342 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14343 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U14344 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12736) );
  OAI211_X1 U14345 ( .C1(n15483), .C2(n13651), .A(n12736), .B(n15482), .ZN(
        n12737) );
  INV_X1 U14346 ( .A(n12737), .ZN(n12738) );
  NAND4_X1 U14347 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12749) );
  AOI22_X1 U14348 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U14349 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U14350 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12745) );
  INV_X1 U14351 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U14352 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12742) );
  OAI211_X1 U14353 ( .C1(n15483), .C2(n13641), .A(n12742), .B(n12819), .ZN(
        n12743) );
  INV_X1 U14354 ( .A(n12743), .ZN(n12744) );
  NAND4_X1 U14355 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n12748) );
  NAND2_X1 U14356 ( .A1(n12749), .A2(n12748), .ZN(n12752) );
  NOR2_X1 U14357 ( .A1(n12751), .A2(n12752), .ZN(n12769) );
  INV_X1 U14358 ( .A(n12750), .ZN(n12809) );
  NAND2_X1 U14359 ( .A1(n12809), .A2(n12734), .ZN(n12753) );
  AOI22_X1 U14360 ( .A1(n12769), .A2(n18291), .B1(n12753), .B2(n12752), .ZN(
        n16132) );
  AOI22_X1 U14361 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11024), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U14362 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10980), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U14363 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U14364 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12754) );
  OAI211_X1 U14365 ( .C1(n15483), .C2(n19572), .A(n12754), .B(n15482), .ZN(
        n12755) );
  INV_X1 U14366 ( .A(n12755), .ZN(n12756) );
  NAND4_X1 U14367 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12768) );
  AOI22_X1 U14368 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11000), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U14369 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10979), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U14370 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12764) );
  INV_X1 U14371 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U14372 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12760) );
  OAI211_X1 U14373 ( .C1(n15483), .C2(n12761), .A(n12760), .B(n12819), .ZN(
        n12762) );
  INV_X1 U14374 ( .A(n12762), .ZN(n12763) );
  NAND4_X1 U14375 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12767) );
  AND2_X1 U14376 ( .A1(n12768), .A2(n12767), .ZN(n12771) );
  NAND2_X1 U14377 ( .A1(n12769), .A2(n12771), .ZN(n12807) );
  OAI211_X1 U14378 ( .C1(n12769), .C2(n12771), .A(n12809), .B(n12807), .ZN(
        n12773) );
  INV_X1 U14379 ( .A(n12773), .ZN(n12770) );
  INV_X1 U14380 ( .A(n12771), .ZN(n12772) );
  NOR2_X1 U14381 ( .A1(n18291), .A2(n12772), .ZN(n16123) );
  AOI22_X1 U14382 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11023), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U14383 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U14384 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12777) );
  NAND2_X1 U14385 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12774) );
  OAI211_X1 U14386 ( .C1(n15483), .C2(n19531), .A(n12774), .B(n15482), .ZN(
        n12775) );
  INV_X1 U14387 ( .A(n12775), .ZN(n12776) );
  NAND4_X1 U14388 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12787) );
  AOI22_X1 U14389 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11000), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U14390 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10981), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U14391 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11026), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12783) );
  INV_X1 U14392 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13602) );
  NAND2_X1 U14393 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12780) );
  OAI211_X1 U14394 ( .C1(n15483), .C2(n13602), .A(n12780), .B(n12819), .ZN(
        n12781) );
  INV_X1 U14395 ( .A(n12781), .ZN(n12782) );
  NAND4_X1 U14396 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12782), .ZN(
        n12786) );
  XNOR2_X1 U14397 ( .A(n12807), .B(n12805), .ZN(n12788) );
  NAND2_X1 U14398 ( .A1(n19574), .A2(n12805), .ZN(n16118) );
  AOI22_X1 U14399 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U14400 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10984), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U14401 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12793) );
  NAND2_X1 U14402 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12790) );
  OAI211_X1 U14403 ( .C1(n15483), .C2(n19493), .A(n12790), .B(n15482), .ZN(
        n12791) );
  INV_X1 U14404 ( .A(n12791), .ZN(n12792) );
  NAND4_X1 U14405 ( .A1(n12795), .A2(n12794), .A3(n12793), .A4(n12792), .ZN(
        n12804) );
  AOI22_X1 U14406 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U14407 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10983), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U14408 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11027), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12800) );
  INV_X1 U14409 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12797) );
  NAND2_X1 U14410 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12796) );
  OAI211_X1 U14411 ( .C1(n15483), .C2(n12797), .A(n12796), .B(n12819), .ZN(
        n12798) );
  INV_X1 U14412 ( .A(n12798), .ZN(n12799) );
  NAND4_X1 U14413 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12803) );
  NAND2_X1 U14414 ( .A1(n12804), .A2(n12803), .ZN(n12812) );
  INV_X1 U14415 ( .A(n12812), .ZN(n12811) );
  INV_X1 U14416 ( .A(n12805), .ZN(n12806) );
  OR2_X1 U14417 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  INV_X1 U14418 ( .A(n12808), .ZN(n12810) );
  OR2_X1 U14419 ( .A1(n12808), .A2(n12812), .ZN(n16098) );
  OAI211_X1 U14420 ( .C1(n12811), .C2(n12810), .A(n16098), .B(n12809), .ZN(
        n12827) );
  NOR2_X2 U14421 ( .A1(n12828), .A2(n12827), .ZN(n16097) );
  NOR2_X1 U14422 ( .A1(n18291), .A2(n12812), .ZN(n16109) );
  OAI21_X1 U14423 ( .B1(n15483), .B2(n14610), .A(n15482), .ZN(n12815) );
  INV_X1 U14424 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12813) );
  INV_X1 U14425 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13694) );
  OAI22_X1 U14426 ( .A1(n15485), .A2(n12813), .B1(n10992), .B2(n13694), .ZN(
        n12814) );
  AOI211_X1 U14427 ( .C1(n12533), .C2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12815), .B(n12814), .ZN(n12818) );
  AOI22_X1 U14428 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11024), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U14429 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10981), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12816) );
  NAND3_X1 U14430 ( .A1(n12818), .A2(n12817), .A3(n12816), .ZN(n12826) );
  INV_X1 U14431 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U14432 ( .B1(n15483), .B2(n13692), .A(n12819), .ZN(n12821) );
  INV_X1 U14433 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13693) );
  INV_X1 U14434 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13695) );
  OAI22_X1 U14435 ( .A1(n15485), .A2(n13693), .B1(n10992), .B2(n13695), .ZN(
        n12820) );
  AOI211_X1 U14436 ( .C1(n12533), .C2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n12821), .B(n12820), .ZN(n12824) );
  AOI22_X1 U14437 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11000), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U14438 ( .A1(n10985), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10976), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12822) );
  NAND3_X1 U14439 ( .A1(n12824), .A2(n12823), .A3(n12822), .ZN(n12825) );
  AND2_X1 U14440 ( .A1(n12826), .A2(n12825), .ZN(n16099) );
  NAND2_X1 U14441 ( .A1(n12828), .A2(n12827), .ZN(n16106) );
  INV_X1 U14442 ( .A(n16098), .ZN(n12829) );
  NAND3_X1 U14443 ( .A1(n12829), .A2(n16099), .A3(n18291), .ZN(n15474) );
  AOI22_X1 U14444 ( .A1(n10989), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11000), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U14445 ( .A1(n10979), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U14446 ( .A1(n12831), .A2(n12830), .ZN(n12843) );
  INV_X1 U14447 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U14448 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12531), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12833) );
  AOI21_X1 U14449 ( .B1(n12406), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n15482), .ZN(n12832) );
  OAI211_X1 U14450 ( .C1(n15481), .C2(n12834), .A(n12833), .B(n12832), .ZN(
        n12842) );
  OAI21_X1 U14451 ( .B1(n15483), .B2(n19395), .A(n15482), .ZN(n12837) );
  INV_X1 U14452 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12835) );
  INV_X1 U14453 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13727) );
  OAI22_X1 U14454 ( .A1(n15485), .A2(n12835), .B1(n10992), .B2(n13727), .ZN(
        n12836) );
  AOI211_X1 U14455 ( .C1(n12533), .C2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12837), .B(n12836), .ZN(n12840) );
  AOI22_X1 U14456 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11023), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U14457 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10982), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12838) );
  NAND3_X1 U14458 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(n12841) );
  OAI21_X1 U14459 ( .B1(n12843), .B2(n12842), .A(n12841), .ZN(n15473) );
  XNOR2_X1 U14460 ( .A(n15474), .B(n15473), .ZN(n12844) );
  MUX2_X1 U14461 ( .A(n19302), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12881) );
  NAND2_X1 U14462 ( .A1(n12881), .A2(n12882), .ZN(n12846) );
  NAND2_X1 U14463 ( .A1(n19302), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12845) );
  NAND2_X1 U14464 ( .A1(n12846), .A2(n12845), .ZN(n12875) );
  XNOR2_X1 U14465 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U14466 ( .A1(n12875), .A2(n12874), .ZN(n12873) );
  NAND2_X1 U14467 ( .A1(n17156), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12847) );
  NAND2_X1 U14468 ( .A1(n12873), .A2(n12847), .ZN(n12870) );
  NAND3_X1 U14469 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12890), .A3(
        n16769), .ZN(n12900) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U14471 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U14472 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12849) );
  NAND4_X1 U14474 ( .A1(n12852), .A2(n12851), .A3(n12850), .A4(n12849), .ZN(
        n12858) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U14476 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13033), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U14478 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12853) );
  NAND4_X1 U14479 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12857) );
  MUX2_X1 U14480 ( .A(n12900), .B(n13919), .S(n13268), .Z(n13274) );
  AOI22_X1 U14481 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U14483 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U14484 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12859) );
  NAND4_X1 U14485 ( .A1(n12862), .A2(n12861), .A3(n12860), .A4(n12859), .ZN(
        n12868) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13023), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13033), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U14489 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12863) );
  NAND4_X1 U14490 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  NOR2_X1 U14491 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  NOR2_X1 U14492 ( .A1(n12872), .A2(n12871), .ZN(n12896) );
  MUX2_X1 U14493 ( .A(n13638), .B(n12896), .S(n14822), .Z(n13272) );
  NAND2_X1 U14494 ( .A1(n13274), .A2(n13272), .ZN(n13898) );
  OAI21_X1 U14495 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12897) );
  INV_X1 U14496 ( .A(n12897), .ZN(n12876) );
  AND2_X1 U14497 ( .A1(n14822), .A2(n12876), .ZN(n13267) );
  AOI21_X1 U14498 ( .B1(n18290), .B2(n18291), .A(n12876), .ZN(n12886) );
  AND2_X1 U14499 ( .A1(n12878), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12879) );
  NOR2_X1 U14500 ( .A1(n12882), .A2(n12879), .ZN(n13676) );
  NAND2_X1 U14501 ( .A1(n13676), .A2(n12881), .ZN(n12880) );
  NAND2_X1 U14502 ( .A1(n13268), .A2(n12880), .ZN(n12884) );
  INV_X1 U14503 ( .A(n12881), .ZN(n13894) );
  XNOR2_X1 U14504 ( .A(n13894), .B(n12882), .ZN(n12901) );
  OAI211_X1 U14505 ( .C1(n18291), .C2(n13676), .A(n19628), .B(n12901), .ZN(
        n12883) );
  OAI211_X1 U14506 ( .C1(n12877), .C2(n12897), .A(n12884), .B(n12883), .ZN(
        n12885) );
  OAI21_X1 U14507 ( .B1(n13267), .B2(n12886), .A(n12885), .ZN(n12887) );
  AND3_X1 U14508 ( .A1(n12900), .A2(n12896), .A3(n12887), .ZN(n12888) );
  AOI21_X1 U14509 ( .B1(n13898), .B2(n14822), .A(n12888), .ZN(n12891) );
  OR2_X1 U14510 ( .A1(n12891), .A2(n13899), .ZN(n12892) );
  NAND2_X1 U14511 ( .A1(n13899), .A2(n12445), .ZN(n12893) );
  AND3_X1 U14512 ( .A1(n12397), .A2(n19574), .A3(n13820), .ZN(n12895) );
  INV_X1 U14513 ( .A(n12896), .ZN(n12898) );
  NOR2_X1 U14514 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  NAND2_X1 U14515 ( .A1(n12900), .A2(n12899), .ZN(n13890) );
  INV_X1 U14516 ( .A(n12901), .ZN(n12902) );
  NOR2_X1 U14517 ( .A1(n13890), .A2(n12902), .ZN(n12903) );
  NAND2_X1 U14518 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21735) );
  AND2_X1 U14519 ( .A1(n14096), .A2(n21735), .ZN(n14829) );
  NAND2_X1 U14520 ( .A1(n12905), .A2(n14829), .ZN(n12906) );
  NOR2_X1 U14521 ( .A1(n14833), .A2(n12906), .ZN(n12907) );
  AOI21_X1 U14522 ( .B1(n15112), .B2(n14819), .A(n12907), .ZN(n14779) );
  INV_X1 U14523 ( .A(n12908), .ZN(n12910) );
  NAND2_X1 U14524 ( .A1(n12910), .A2(n12909), .ZN(n12911) );
  NAND2_X1 U14525 ( .A1(n14779), .A2(n12911), .ZN(n12912) );
  INV_X1 U14526 ( .A(n12428), .ZN(n12942) );
  NOR4_X1 U14527 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12916) );
  NOR4_X1 U14528 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12915) );
  NOR4_X1 U14529 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12914) );
  NOR4_X1 U14530 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U14531 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12921) );
  NOR4_X1 U14532 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12919) );
  NOR4_X1 U14533 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12918) );
  NOR4_X1 U14534 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12917) );
  NAND4_X1 U14535 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n19738), .ZN(
        n12920) );
  OAI21_X4 U14536 ( .B1(n12921), .B2(n12920), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14182) );
  NAND2_X1 U14537 ( .A1(n12922), .A2(n14182), .ZN(n12923) );
  NOR2_X2 U14538 ( .A1(n19613), .A2(n12923), .ZN(n19617) );
  NAND2_X2 U14539 ( .A1(n13094), .A2(n12925), .ZN(n13089) );
  INV_X1 U14540 ( .A(n13089), .ZN(n13085) );
  INV_X1 U14541 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n12924) );
  INV_X1 U14542 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14025) );
  OAI22_X1 U14543 ( .A1(n11407), .A2(n12924), .B1(n13039), .B2(n14025), .ZN(
        n12927) );
  INV_X1 U14544 ( .A(n12964), .ZN(n13038) );
  NOR2_X1 U14545 ( .A1(n13038), .A2(n14884), .ZN(n12926) );
  AOI211_X1 U14546 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n13085), .A(n12927), .B(
        n12926), .ZN(n14484) );
  OR2_X1 U14547 ( .A1(n13089), .A2(n12472), .ZN(n12929) );
  AOI22_X1 U14548 ( .A1(n13252), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12941), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12928) );
  NAND2_X1 U14549 ( .A1(n12929), .A2(n12928), .ZN(n12963) );
  INV_X1 U14550 ( .A(n12963), .ZN(n12949) );
  AOI22_X1 U14551 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U14552 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U14553 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U14554 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12931) );
  NAND4_X1 U14555 ( .A1(n12934), .A2(n12933), .A3(n12932), .A4(n12931), .ZN(
        n12940) );
  AOI22_X1 U14556 ( .A1(n12648), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U14557 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U14558 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U14559 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12935) );
  NAND4_X1 U14560 ( .A1(n12938), .A2(n12937), .A3(n12936), .A4(n12935), .ZN(
        n12939) );
  NAND2_X1 U14561 ( .A1(n12964), .A2(n13906), .ZN(n12944) );
  NAND2_X1 U14562 ( .A1(n12942), .A2(n12941), .ZN(n12975) );
  MUX2_X1 U14563 ( .A(n12425), .B(n17147), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12943) );
  INV_X1 U14564 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n17170) );
  INV_X1 U14565 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U14566 ( .A1(n18291), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12945) );
  OAI211_X1 U14567 ( .C1(n12425), .C2(n12946), .A(n12945), .B(n19293), .ZN(
        n12947) );
  INV_X1 U14568 ( .A(n12947), .ZN(n12948) );
  AOI22_X1 U14569 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13023), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U14570 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U14571 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12675), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U14572 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13033), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12950) );
  NAND4_X1 U14573 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n12959) );
  AOI22_X1 U14574 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U14575 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U14576 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12637), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U14577 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12954) );
  NAND4_X1 U14578 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12958) );
  NOR2_X1 U14579 ( .A1(n12959), .A2(n12958), .ZN(n13908) );
  OR2_X1 U14580 ( .A1(n13908), .A2(n13038), .ZN(n12962) );
  AND2_X1 U14581 ( .A1(n12428), .A2(n12425), .ZN(n14372) );
  INV_X1 U14582 ( .A(n14372), .ZN(n12960) );
  MUX2_X1 U14583 ( .A(n12960), .B(n19302), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12961) );
  AND2_X1 U14584 ( .A1(n12962), .A2(n12961), .ZN(n14436) );
  OR2_X1 U14585 ( .A1(n14376), .A2(n12963), .ZN(n12978) );
  AOI22_X1 U14586 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13028), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U14587 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n12848), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U14588 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U14589 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12700), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U14590 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n12974) );
  AOI22_X1 U14591 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12648), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U14592 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13033), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U14593 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U14594 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12969) );
  NAND4_X1 U14595 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12973) );
  NAND2_X1 U14596 ( .A1(n12964), .A2(n13668), .ZN(n12976) );
  OAI211_X1 U14597 ( .C1(n19293), .C2(n17156), .A(n12976), .B(n12975), .ZN(
        n12977) );
  AND3_X1 U14598 ( .A1(n14435), .A2(n12978), .A3(n12977), .ZN(n12979) );
  INV_X1 U14599 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17217) );
  OR2_X1 U14600 ( .A1(n13089), .A2(n17217), .ZN(n12981) );
  INV_X2 U14601 ( .A(n13039), .ZN(n13090) );
  AOI22_X1 U14602 ( .A1(n13252), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13090), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U14603 ( .A1(n12981), .A2(n12980), .ZN(n14340) );
  NOR2_X1 U14604 ( .A1(n14339), .A2(n14340), .ZN(n12982) );
  INV_X1 U14605 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17218) );
  NAND2_X1 U14606 ( .A1(n13252), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U14607 ( .A1(n13090), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12984) );
  OAI211_X1 U14608 ( .C1(n19293), .C2(n19175), .A(n12985), .B(n12984), .ZN(
        n12986) );
  INV_X1 U14609 ( .A(n12986), .ZN(n12988) );
  NAND2_X1 U14610 ( .A1(n12964), .A2(n13638), .ZN(n12987) );
  OAI211_X1 U14611 ( .C1(n13089), .C2(n17218), .A(n12988), .B(n12987), .ZN(
        n14859) );
  NAND2_X1 U14612 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  INV_X1 U14613 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12989) );
  OR2_X1 U14614 ( .A1(n13089), .A2(n12989), .ZN(n12992) );
  AOI22_X1 U14615 ( .A1(n13252), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13090), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U14616 ( .A1(n12964), .A2(n13919), .ZN(n12990) );
  AOI22_X1 U14617 ( .A1(n13085), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n13252), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U14618 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14619 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U14620 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U14621 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12993) );
  NAND4_X1 U14622 ( .A1(n12996), .A2(n12995), .A3(n12994), .A4(n12993), .ZN(
        n13002) );
  AOI22_X1 U14623 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U14624 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12637), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U14625 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14626 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12997) );
  NAND4_X1 U14627 ( .A1(n13000), .A2(n12999), .A3(n12998), .A4(n12997), .ZN(
        n13001) );
  AOI22_X1 U14628 ( .A1(n12964), .A2(n13275), .B1(n13090), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U14629 ( .A1(n13004), .A2(n13003), .ZN(n15176) );
  AOI22_X1 U14630 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U14631 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12592), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14632 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12559), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U14633 ( .A1(n13033), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U14634 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13014) );
  AOI22_X1 U14635 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12564), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U14636 ( .A1(n12637), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12700), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U14637 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U14638 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13009) );
  NAND4_X1 U14639 ( .A1(n13012), .A2(n13011), .A3(n13010), .A4(n13009), .ZN(
        n13013) );
  NAND2_X1 U14640 ( .A1(n13748), .A2(n12964), .ZN(n13015) );
  INV_X1 U14641 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n18334) );
  OR2_X1 U14642 ( .A1(n13089), .A2(n18334), .ZN(n13017) );
  AOI22_X1 U14643 ( .A1(n13252), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13090), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U14644 ( .A1(n12848), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13021) );
  NAND2_X1 U14645 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13020) );
  NAND2_X1 U14646 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13019) );
  NAND2_X1 U14647 ( .A1(n12559), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13018) );
  AOI22_X1 U14648 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13022), .B1(
        n12550), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U14649 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U14650 ( .A1(n13023), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13025) );
  NAND2_X1 U14651 ( .A1(n12564), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13024) );
  NAND2_X1 U14652 ( .A1(n13028), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13032) );
  NAND2_X1 U14653 ( .A1(n12592), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13031) );
  NAND2_X1 U14654 ( .A1(n12700), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13030) );
  NAND2_X1 U14655 ( .A1(n12637), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13029) );
  AOI22_X1 U14656 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13033), .B1(
        n14812), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13034) );
  INV_X1 U14657 ( .A(n13276), .ZN(n13596) );
  INV_X1 U14658 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16707) );
  INV_X1 U14659 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18347) );
  INV_X1 U14660 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17196) );
  OAI222_X1 U14661 ( .A1(n16707), .A2(n13039), .B1(n13089), .B2(n18347), .C1(
        n11407), .C2(n17196), .ZN(n14480) );
  INV_X1 U14662 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U14663 ( .A1(n13252), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13090), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U14664 ( .A1(n12964), .A2(n14697), .ZN(n13040) );
  OAI211_X1 U14665 ( .C1(n13089), .C2(n13042), .A(n13041), .B(n13040), .ZN(
        n14487) );
  INV_X1 U14666 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n15038) );
  OR2_X1 U14667 ( .A1(n13089), .A2(n15038), .ZN(n13045) );
  AOI22_X1 U14668 ( .A1(n13252), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U14669 ( .A1(n12964), .A2(n14905), .ZN(n13043) );
  INV_X1 U14670 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16663) );
  AOI22_X1 U14671 ( .A1(n13252), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U14672 ( .A1(n12964), .A2(n14941), .ZN(n13046) );
  OAI211_X1 U14673 ( .C1(n13089), .C2(n16663), .A(n13047), .B(n13046), .ZN(
        n14596) );
  INV_X1 U14674 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13048) );
  OR2_X1 U14675 ( .A1(n13089), .A2(n13048), .ZN(n13052) );
  AOI22_X1 U14676 ( .A1(n13252), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13051) );
  INV_X1 U14677 ( .A(n13049), .ZN(n15024) );
  NAND2_X1 U14678 ( .A1(n12964), .A2(n15024), .ZN(n13050) );
  NOR2_X2 U14679 ( .A1(n16642), .A2(n16641), .ZN(n14675) );
  INV_X1 U14680 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U14681 ( .A1(n13252), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U14682 ( .A1(n12964), .A2(n15049), .ZN(n13053) );
  OAI211_X1 U14683 ( .C1(n13089), .C2(n13055), .A(n13054), .B(n13053), .ZN(
        n14674) );
  NAND2_X1 U14684 ( .A1(n14675), .A2(n14674), .ZN(n18415) );
  INV_X1 U14685 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13056) );
  OR2_X1 U14686 ( .A1(n13089), .A2(n13056), .ZN(n13059) );
  AOI22_X1 U14687 ( .A1(n13252), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13058) );
  NAND2_X1 U14688 ( .A1(n12964), .A2(n15138), .ZN(n13057) );
  INV_X1 U14689 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U14690 ( .A1(n13252), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13061) );
  NAND2_X1 U14691 ( .A1(n12964), .A2(n15151), .ZN(n13060) );
  OAI211_X1 U14692 ( .C1(n13089), .C2(n13062), .A(n13061), .B(n13060), .ZN(
        n14935) );
  INV_X1 U14693 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n13063) );
  OR2_X1 U14694 ( .A1(n13089), .A2(n13063), .ZN(n13065) );
  AOI22_X1 U14695 ( .A1(n13252), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13064) );
  NAND2_X1 U14696 ( .A1(n13065), .A2(n13064), .ZN(n16078) );
  INV_X1 U14697 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18439) );
  OR2_X1 U14698 ( .A1(n13089), .A2(n18439), .ZN(n13067) );
  AOI22_X1 U14699 ( .A1(n13252), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13066) );
  NAND2_X1 U14700 ( .A1(n13067), .A2(n13066), .ZN(n15213) );
  INV_X1 U14701 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n18452) );
  OR2_X1 U14702 ( .A1(n13089), .A2(n18452), .ZN(n13069) );
  AOI22_X1 U14703 ( .A1(n13252), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13068) );
  INV_X1 U14704 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17220) );
  OR2_X1 U14705 ( .A1(n13089), .A2(n17220), .ZN(n13071) );
  AOI22_X1 U14706 ( .A1(n13252), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U14707 ( .A1(n13071), .A2(n13070), .ZN(n16246) );
  INV_X1 U14708 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17221) );
  OR2_X1 U14709 ( .A1(n13089), .A2(n17221), .ZN(n13073) );
  AOI22_X1 U14710 ( .A1(n13252), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13072) );
  NAND2_X1 U14711 ( .A1(n13073), .A2(n13072), .ZN(n16065) );
  INV_X1 U14712 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18474) );
  OR2_X1 U14713 ( .A1(n13089), .A2(n18474), .ZN(n13075) );
  AOI22_X1 U14714 ( .A1(n13252), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U14715 ( .A1(n13075), .A2(n13074), .ZN(n16236) );
  INV_X1 U14716 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U14717 ( .A1(n13252), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13076) );
  OAI21_X1 U14718 ( .B1(n13089), .B2(n13077), .A(n13076), .ZN(n16052) );
  INV_X1 U14719 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U14720 ( .A1(n13252), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13078) );
  OAI21_X1 U14721 ( .B1(n13089), .B2(n17222), .A(n13078), .ZN(n16227) );
  INV_X1 U14722 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U14723 ( .A1(n13252), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13079) );
  OAI21_X1 U14724 ( .B1(n13089), .B2(n17223), .A(n13079), .ZN(n16218) );
  NAND2_X1 U14725 ( .A1(n13085), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U14726 ( .A1(n13252), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13080) );
  AND2_X1 U14727 ( .A1(n13081), .A2(n13080), .ZN(n16207) );
  NAND2_X1 U14728 ( .A1(n13085), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U14729 ( .A1(n13252), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13082) );
  AND2_X1 U14730 ( .A1(n13083), .A2(n13082), .ZN(n16198) );
  NAND2_X1 U14731 ( .A1(n13085), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U14732 ( .A1(n13252), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13086) );
  AND2_X1 U14733 ( .A1(n13087), .A2(n13086), .ZN(n16189) );
  INV_X1 U14734 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16291) );
  AOI22_X1 U14735 ( .A1(n13252), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13088) );
  OAI21_X1 U14736 ( .B1(n13089), .B2(n16291), .A(n13088), .ZN(n16181) );
  INV_X1 U14737 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U14738 ( .A1(n13252), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13091) );
  OAI21_X1 U14739 ( .B1(n13089), .B2(n17227), .A(n13091), .ZN(n13251) );
  INV_X1 U14740 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14392) );
  OAI22_X1 U14741 ( .A1(n16201), .A2(n18563), .B1(n16250), .B2(n14392), .ZN(
        n13092) );
  AOI21_X1 U14742 ( .B1(n19617), .B2(BUF2_REG_29__SCAN_IN), .A(n13092), .ZN(
        n13096) );
  NOR3_X2 U14743 ( .A1(n19613), .A2(n14182), .A3(n13093), .ZN(n19616) );
  NAND2_X1 U14744 ( .A1(n16250), .A2(n13094), .ZN(n16251) );
  AOI22_X1 U14745 ( .A1(n17039), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n14182), .ZN(n14676) );
  INV_X1 U14746 ( .A(n14676), .ZN(n14138) );
  AOI22_X1 U14747 ( .A1(n19616), .A2(BUF1_REG_29__SCAN_IN), .B1(n19615), .B2(
        n14138), .ZN(n13095) );
  OAI21_X1 U14748 ( .B1(n16096), .B2(n19398), .A(n13097), .ZN(P2_U2890) );
  NAND2_X1 U14749 ( .A1(n13102), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13115) );
  INV_X1 U14750 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U14751 ( .A1(n13099), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13101) );
  INV_X1 U14752 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U14753 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13997) );
  AOI21_X1 U14754 ( .B1(n18413), .B2(n13113), .A(n13102), .ZN(n18410) );
  AOI21_X1 U14755 ( .B1(n18382), .B2(n13103), .A(n13114), .ZN(n18388) );
  AOI21_X1 U14756 ( .B1(n17094), .B2(n13110), .A(n13112), .ZN(n17086) );
  AOI21_X1 U14757 ( .B1(n17079), .B2(n13104), .A(n13111), .ZN(n17070) );
  AOI21_X1 U14758 ( .B1(n17069), .B2(n13105), .A(n13106), .ZN(n18329) );
  AOI21_X1 U14759 ( .B1(n17064), .B2(n13107), .A(n13108), .ZN(n18312) );
  INV_X1 U14760 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U14761 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n14161), .B2(n14089), .ZN(
        n15095) );
  AOI22_X1 U14762 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18286), .ZN(n15124) );
  AOI22_X1 U14763 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14089), .B2(n18286), .ZN(
        n15123) );
  NAND2_X1 U14764 ( .A1(n15124), .A2(n15123), .ZN(n15094) );
  NOR2_X1 U14765 ( .A1(n15095), .A2(n15094), .ZN(n14960) );
  NOR2_X1 U14766 ( .A1(n14089), .A2(n14161), .ZN(n13109) );
  OAI21_X1 U14767 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13109), .A(
        n13107), .ZN(n14961) );
  NAND2_X1 U14768 ( .A1(n14960), .A2(n14961), .ZN(n18309) );
  NOR2_X1 U14769 ( .A1(n18312), .A2(n18309), .ZN(n18317) );
  OAI21_X1 U14770 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13108), .A(
        n13105), .ZN(n18319) );
  NAND2_X1 U14771 ( .A1(n18317), .A2(n18319), .ZN(n18328) );
  NOR2_X1 U14772 ( .A1(n18329), .A2(n18328), .ZN(n18342) );
  OAI21_X1 U14773 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13106), .A(
        n13104), .ZN(n18344) );
  NAND2_X1 U14774 ( .A1(n18342), .A2(n18344), .ZN(n15076) );
  NOR2_X1 U14775 ( .A1(n17070), .A2(n15076), .ZN(n18358) );
  OAI21_X1 U14776 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n13111), .A(
        n13110), .ZN(n18359) );
  NAND2_X1 U14777 ( .A1(n18358), .A2(n18359), .ZN(n15033) );
  NOR2_X1 U14778 ( .A1(n17086), .A2(n15033), .ZN(n18377) );
  OAI21_X1 U14779 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13112), .A(
        n13103), .ZN(n18380) );
  NAND2_X1 U14780 ( .A1(n18377), .A2(n18380), .ZN(n18386) );
  NOR2_X1 U14781 ( .A1(n18388), .A2(n18386), .ZN(n18397) );
  OAI21_X1 U14782 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n13114), .A(
        n13113), .ZN(n18408) );
  NAND2_X1 U14783 ( .A1(n18397), .A2(n18408), .ZN(n18396) );
  NOR2_X1 U14784 ( .A1(n18410), .A2(n18396), .ZN(n18425) );
  OAI21_X1 U14785 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n13102), .A(
        n13115), .ZN(n18430) );
  NAND2_X1 U14786 ( .A1(n18425), .A2(n18430), .ZN(n18423) );
  AOI21_X1 U14787 ( .B1(n16084), .B2(n13115), .A(n13117), .ZN(n13116) );
  INV_X1 U14788 ( .A(n13116), .ZN(n16076) );
  OAI21_X1 U14789 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13117), .A(
        n13118), .ZN(n18447) );
  NAND2_X1 U14790 ( .A1(n15113), .A2(n18445), .ZN(n18458) );
  AOI21_X1 U14791 ( .B1(n13118), .B2(n16398), .A(n13119), .ZN(n16395) );
  INV_X1 U14792 ( .A(n16395), .ZN(n18459) );
  NAND2_X1 U14793 ( .A1(n18584), .A2(n18457), .ZN(n18469) );
  OAI21_X1 U14794 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n13119), .A(
        n11086), .ZN(n18470) );
  NAND2_X1 U14795 ( .A1(n18469), .A2(n18470), .ZN(n18468) );
  NAND2_X1 U14796 ( .A1(n18584), .A2(n18468), .ZN(n16061) );
  INV_X1 U14797 ( .A(n13120), .ZN(n13122) );
  NAND2_X1 U14798 ( .A1(n13098), .A2(n11086), .ZN(n13121) );
  NAND2_X1 U14799 ( .A1(n13122), .A2(n13121), .ZN(n16377) );
  OAI21_X1 U14800 ( .B1(n13120), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11045), .ZN(n18483) );
  AOI21_X1 U14801 ( .B1(n11045), .B2(n16054), .A(n13123), .ZN(n13124) );
  INV_X1 U14802 ( .A(n13124), .ZN(n16353) );
  NAND2_X1 U14803 ( .A1(n16047), .A2(n18584), .ZN(n18495) );
  OAI21_X1 U14804 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n13123), .A(
        n13127), .ZN(n18496) );
  NAND2_X1 U14805 ( .A1(n18495), .A2(n18496), .ZN(n18494) );
  NAND2_X1 U14806 ( .A1(n18584), .A2(n18494), .ZN(n18504) );
  INV_X1 U14807 ( .A(n13125), .ZN(n13130) );
  NAND2_X1 U14808 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  NAND2_X1 U14809 ( .A1(n13130), .A2(n13128), .ZN(n18505) );
  NAND2_X1 U14810 ( .A1(n18503), .A2(n18584), .ZN(n18514) );
  INV_X1 U14811 ( .A(n13131), .ZN(n13129) );
  AOI21_X1 U14812 ( .B1(n16320), .B2(n13130), .A(n13129), .ZN(n16322) );
  INV_X1 U14813 ( .A(n16322), .ZN(n18515) );
  NAND2_X1 U14814 ( .A1(n18514), .A2(n18515), .ZN(n18513) );
  NAND2_X1 U14815 ( .A1(n18513), .A2(n18584), .ZN(n18529) );
  AND2_X1 U14816 ( .A1(n13131), .A2(n13226), .ZN(n13133) );
  OR2_X1 U14817 ( .A1(n13133), .A2(n13132), .ZN(n18530) );
  NAND2_X1 U14818 ( .A1(n18529), .A2(n18530), .ZN(n18528) );
  NAND2_X1 U14819 ( .A1(n18528), .A2(n18584), .ZN(n18542) );
  INV_X1 U14820 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16299) );
  INV_X1 U14821 ( .A(n13132), .ZN(n13135) );
  AOI21_X1 U14822 ( .B1(n16299), .B2(n13135), .A(n13134), .ZN(n16302) );
  INV_X1 U14823 ( .A(n16302), .ZN(n18543) );
  NAND2_X1 U14824 ( .A1(n18542), .A2(n18543), .ZN(n18541) );
  NAND2_X1 U14825 ( .A1(n18541), .A2(n18584), .ZN(n18554) );
  NOR2_X1 U14826 ( .A1(n13134), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13137) );
  OR2_X1 U14827 ( .A1(n13136), .A2(n13137), .ZN(n18555) );
  NAND2_X1 U14828 ( .A1(n18553), .A2(n18584), .ZN(n18567) );
  OR2_X1 U14829 ( .A1(n13136), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13139) );
  AND2_X1 U14830 ( .A1(n13139), .A2(n13138), .ZN(n16276) );
  INV_X1 U14831 ( .A(n16276), .ZN(n18568) );
  NAND2_X1 U14832 ( .A1(n18567), .A2(n18568), .ZN(n18566) );
  NAND2_X1 U14833 ( .A1(n18566), .A2(n18584), .ZN(n18583) );
  INV_X1 U14834 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13140) );
  XNOR2_X1 U14835 ( .A(n13138), .B(n13140), .ZN(n18585) );
  NAND2_X1 U14836 ( .A1(n18583), .A2(n18585), .ZN(n13141) );
  INV_X1 U14837 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19335) );
  NAND4_X1 U14838 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18286), .A3(n19335), 
        .A4(n21698), .ZN(n18627) );
  NAND2_X1 U14839 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13147) );
  INV_X1 U14840 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n13287) );
  INV_X1 U14841 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13144) );
  OAI22_X1 U14842 ( .A1(n13228), .A2(n13287), .B1(n14093), .B2(n13144), .ZN(
        n13145) );
  AOI21_X1 U14843 ( .B1(n13243), .B2(P2_REIP_REG_23__SCAN_IN), .A(n13145), 
        .ZN(n13146) );
  NAND2_X1 U14844 ( .A1(n13147), .A2(n13146), .ZN(n16141) );
  NAND2_X1 U14845 ( .A1(n13149), .A2(n13148), .ZN(n13151) );
  NAND2_X1 U14846 ( .A1(n13151), .A2(n13150), .ZN(n13155) );
  OR2_X1 U14847 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  NAND2_X1 U14848 ( .A1(n13155), .A2(n13154), .ZN(n14499) );
  INV_X1 U14849 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U14850 ( .A1(n13243), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U14851 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13156) );
  OAI211_X1 U14852 ( .C1(n13273), .C2(n13228), .A(n13157), .B(n13156), .ZN(
        n13158) );
  AOI21_X1 U14853 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13158), .ZN(n14498) );
  OR2_X2 U14854 ( .A1(n14499), .A2(n14498), .ZN(n14501) );
  NAND2_X1 U14855 ( .A1(n13243), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U14856 ( .A1(n13159), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13160) );
  NAND2_X1 U14857 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  AOI21_X1 U14858 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13162), .ZN(n14490) );
  NAND2_X1 U14859 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13165) );
  INV_X1 U14860 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14618) );
  OAI22_X1 U14861 ( .A1(n13228), .A2(n14618), .B1(n14093), .B2(n17069), .ZN(
        n13163) );
  AOI21_X1 U14862 ( .B1(n13243), .B2(P2_REIP_REG_6__SCAN_IN), .A(n13163), .ZN(
        n13164) );
  NAND2_X1 U14863 ( .A1(n13165), .A2(n13164), .ZN(n14613) );
  NAND2_X1 U14864 ( .A1(n13243), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U14865 ( .A1(n13159), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13166) );
  NAND2_X1 U14866 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  AOI21_X1 U14867 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13168), .ZN(n14538) );
  NAND2_X1 U14868 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13171) );
  INV_X1 U14869 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13278) );
  OAI22_X1 U14870 ( .A1(n13228), .A2(n13278), .B1(n14093), .B2(n17079), .ZN(
        n13169) );
  AOI21_X1 U14871 ( .B1(n13243), .B2(P2_REIP_REG_8__SCAN_IN), .A(n13169), .ZN(
        n13170) );
  NAND2_X1 U14872 ( .A1(n13171), .A2(n13170), .ZN(n14881) );
  NAND2_X1 U14873 ( .A1(n13243), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U14874 ( .A1(n13159), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13172) );
  NAND2_X1 U14875 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  AOI21_X1 U14876 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13174), .ZN(n14699) );
  NAND2_X1 U14877 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13177) );
  INV_X1 U14878 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13279) );
  OAI22_X1 U14879 ( .A1(n13228), .A2(n13279), .B1(n14093), .B2(n17094), .ZN(
        n13175) );
  AOI21_X1 U14880 ( .B1(n13243), .B2(P2_REIP_REG_10__SCAN_IN), .A(n13175), 
        .ZN(n13176) );
  NAND2_X1 U14881 ( .A1(n13177), .A2(n13176), .ZN(n14901) );
  NAND2_X1 U14882 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13180) );
  INV_X1 U14883 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13280) );
  OAI22_X1 U14884 ( .A1(n13228), .A2(n13280), .B1(n14093), .B2(n11226), .ZN(
        n13178) );
  AOI21_X1 U14885 ( .B1(n13243), .B2(P2_REIP_REG_11__SCAN_IN), .A(n13178), 
        .ZN(n13179) );
  NAND2_X1 U14886 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13183) );
  INV_X1 U14887 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13281) );
  OAI22_X1 U14888 ( .A1(n13228), .A2(n13281), .B1(n14093), .B2(n18382), .ZN(
        n13181) );
  AOI21_X1 U14889 ( .B1(n13243), .B2(P2_REIP_REG_12__SCAN_IN), .A(n13181), 
        .ZN(n13182) );
  NAND2_X1 U14890 ( .A1(n13183), .A2(n13182), .ZN(n15020) );
  NAND2_X1 U14891 ( .A1(n15019), .A2(n15020), .ZN(n15050) );
  NAND2_X1 U14892 ( .A1(n13243), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U14893 ( .A1(n13159), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n13184) );
  NAND2_X1 U14894 ( .A1(n13185), .A2(n13184), .ZN(n13186) );
  AOI21_X1 U14895 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n13186), .ZN(n15051) );
  NAND2_X1 U14896 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13189) );
  INV_X1 U14897 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13282) );
  OAI22_X1 U14898 ( .A1(n13228), .A2(n13282), .B1(n14093), .B2(n18413), .ZN(
        n13187) );
  AOI21_X1 U14899 ( .B1(n13243), .B2(P2_REIP_REG_14__SCAN_IN), .A(n13187), 
        .ZN(n13188) );
  NAND2_X1 U14900 ( .A1(n13189), .A2(n13188), .ZN(n15134) );
  NAND2_X1 U14901 ( .A1(n15052), .A2(n15134), .ZN(n15133) );
  NAND2_X1 U14902 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13193) );
  INV_X1 U14903 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13283) );
  INV_X1 U14904 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13190) );
  OAI22_X1 U14905 ( .A1(n13228), .A2(n13283), .B1(n14093), .B2(n13190), .ZN(
        n13191) );
  AOI21_X1 U14906 ( .B1(n13243), .B2(P2_REIP_REG_15__SCAN_IN), .A(n13191), 
        .ZN(n13192) );
  NAND2_X1 U14907 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13197) );
  INV_X1 U14908 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13194) );
  OAI22_X1 U14909 ( .A1(n13228), .A2(n13194), .B1(n14093), .B2(n16084), .ZN(
        n13195) );
  AOI21_X1 U14910 ( .B1(n13243), .B2(P2_REIP_REG_16__SCAN_IN), .A(n13195), 
        .ZN(n13196) );
  NAND2_X1 U14911 ( .A1(n13197), .A2(n13196), .ZN(n14081) );
  NAND2_X1 U14912 ( .A1(n13243), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U14913 ( .A1(n13159), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n13198) );
  NAND2_X1 U14914 ( .A1(n13199), .A2(n13198), .ZN(n13200) );
  AOI21_X1 U14915 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13200), .ZN(n16172) );
  NAND2_X1 U14916 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13203) );
  INV_X1 U14917 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n13284) );
  OAI22_X1 U14918 ( .A1(n13228), .A2(n13284), .B1(n14093), .B2(n16398), .ZN(
        n13201) );
  AOI21_X1 U14919 ( .B1(n13243), .B2(P2_REIP_REG_18__SCAN_IN), .A(n13201), 
        .ZN(n13202) );
  INV_X1 U14920 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n13285) );
  NAND2_X1 U14921 ( .A1(n13243), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U14922 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13204) );
  OAI211_X1 U14923 ( .C1(n13285), .C2(n13228), .A(n13205), .B(n13204), .ZN(
        n13206) );
  AOI21_X1 U14924 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n13206), .ZN(n16160) );
  NAND2_X1 U14925 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13210) );
  INV_X1 U14926 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n13207) );
  OAI22_X1 U14927 ( .A1(n13228), .A2(n13207), .B1(n14093), .B2(n13098), .ZN(
        n13208) );
  AOI21_X1 U14928 ( .B1(n13243), .B2(P2_REIP_REG_20__SCAN_IN), .A(n13208), 
        .ZN(n13209) );
  NAND2_X1 U14929 ( .A1(n13210), .A2(n13209), .ZN(n16062) );
  AND2_X2 U14930 ( .A1(n16161), .A2(n16062), .ZN(n16152) );
  NAND2_X1 U14931 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13214) );
  INV_X1 U14932 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n13211) );
  OAI22_X1 U14933 ( .A1(n13228), .A2(n13211), .B1(n14093), .B2(n16054), .ZN(
        n13212) );
  AOI21_X1 U14934 ( .B1(n13243), .B2(P2_REIP_REG_22__SCAN_IN), .A(n13212), 
        .ZN(n13213) );
  NAND2_X1 U14935 ( .A1(n13214), .A2(n13213), .ZN(n16049) );
  NAND2_X1 U14936 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13218) );
  INV_X1 U14937 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n13819) );
  INV_X1 U14938 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13215) );
  OAI22_X1 U14939 ( .A1(n13228), .A2(n13819), .B1(n14093), .B2(n13215), .ZN(
        n13216) );
  AOI21_X1 U14940 ( .B1(n13243), .B2(P2_REIP_REG_21__SCAN_IN), .A(n13216), 
        .ZN(n13217) );
  NAND2_X1 U14941 ( .A1(n13218), .A2(n13217), .ZN(n16151) );
  NAND2_X1 U14942 ( .A1(n16141), .A2(n16050), .ZN(n16140) );
  NAND2_X1 U14943 ( .A1(n13243), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U14944 ( .A1(n13159), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n13220) );
  NAND2_X1 U14945 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  AOI21_X1 U14946 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n13222), .ZN(n16135) );
  OR2_X2 U14947 ( .A1(n16140), .A2(n16135), .ZN(n16133) );
  NAND2_X1 U14948 ( .A1(n13243), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U14949 ( .A1(n13159), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n13223) );
  NAND2_X1 U14950 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  AOI21_X1 U14951 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n13225), .ZN(n16126) );
  NAND2_X1 U14952 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13231) );
  INV_X1 U14953 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n13227) );
  OAI22_X1 U14954 ( .A1(n13228), .A2(n13227), .B1(n14093), .B2(n13226), .ZN(
        n13229) );
  AOI21_X1 U14955 ( .B1(n13243), .B2(P2_REIP_REG_26__SCAN_IN), .A(n13229), 
        .ZN(n13230) );
  NAND2_X1 U14956 ( .A1(n13231), .A2(n13230), .ZN(n16115) );
  NAND2_X1 U14957 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13234) );
  INV_X1 U14958 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13290) );
  OAI22_X1 U14959 ( .A1(n13228), .A2(n13290), .B1(n14093), .B2(n16299), .ZN(
        n13232) );
  AOI21_X1 U14960 ( .B1(n13243), .B2(P2_REIP_REG_27__SCAN_IN), .A(n13232), 
        .ZN(n13233) );
  NAND2_X1 U14961 ( .A1(n13234), .A2(n13233), .ZN(n16111) );
  NAND2_X1 U14962 ( .A1(n13242), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13238) );
  INV_X1 U14963 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n13291) );
  INV_X1 U14964 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13235) );
  OAI22_X1 U14965 ( .A1(n13228), .A2(n13291), .B1(n14093), .B2(n13235), .ZN(
        n13236) );
  AOI21_X1 U14966 ( .B1(n13243), .B2(P2_REIP_REG_28__SCAN_IN), .A(n13236), 
        .ZN(n13237) );
  NAND2_X1 U14967 ( .A1(n13238), .A2(n13237), .ZN(n16103) );
  NAND2_X1 U14968 ( .A1(n13243), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U14969 ( .A1(n13159), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n13239) );
  NAND2_X1 U14970 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  AOI21_X1 U14971 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13241), .ZN(n16092) );
  NAND2_X1 U14972 ( .A1(n13243), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U14973 ( .A1(n13159), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13244) );
  NAND2_X1 U14974 ( .A1(n13245), .A2(n13244), .ZN(n13246) );
  AOI21_X1 U14975 ( .B1(n13242), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13246), .ZN(n13994) );
  AND2_X1 U14976 ( .A1(n14009), .A2(n18634), .ZN(n13248) );
  OR2_X1 U14977 ( .A1(n13249), .A2(n18644), .ZN(n14146) );
  INV_X1 U14978 ( .A(n21735), .ZN(n18630) );
  NOR2_X1 U14979 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n18630), .ZN(n13294) );
  AND2_X1 U14980 ( .A1(n13268), .A2(n13294), .ZN(n13250) );
  INV_X1 U14981 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U14982 ( .A1(n13252), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U14983 ( .B1(n13089), .B2(n17228), .A(n13253), .ZN(n13254) );
  NAND2_X1 U14984 ( .A1(n14005), .A2(n13256), .ZN(n15498) );
  NAND2_X1 U14985 ( .A1(n19574), .A2(n14009), .ZN(n14820) );
  NAND2_X2 U14986 ( .A1(n17237), .A2(n21752), .ZN(n17230) );
  NOR2_X1 U14987 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n21749) );
  NAND2_X1 U14988 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21749), .ZN(n17215) );
  NAND2_X1 U14989 ( .A1(n17230), .A2(n17215), .ZN(n18292) );
  NAND2_X1 U14990 ( .A1(n21735), .A2(n18292), .ZN(n14831) );
  NOR2_X1 U14991 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14831), .ZN(n13258) );
  INV_X1 U14992 ( .A(n13258), .ZN(n13257) );
  NOR2_X1 U14993 ( .A1(n14820), .A2(n13257), .ZN(n14850) );
  OR2_X1 U14994 ( .A1(n14267), .A2(n13258), .ZN(n18573) );
  OR2_X1 U14995 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13294), .ZN(n13259) );
  OR2_X1 U14996 ( .A1(n14100), .A2(n13259), .ZN(n13260) );
  NOR2_X1 U14997 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18286), .ZN(n18629) );
  NAND3_X1 U14998 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n18629), .A3(n14093), 
        .ZN(n18641) );
  INV_X1 U14999 ( .A(n18641), .ZN(n13263) );
  NAND2_X1 U15000 ( .A1(n13261), .A2(n19321), .ZN(n14035) );
  NAND2_X1 U15001 ( .A1(n18381), .A2(n18627), .ZN(n13262) );
  AOI22_X1 U15002 ( .A1(n18561), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18577), .ZN(n13265) );
  NAND2_X1 U15003 ( .A1(n18576), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13264) );
  OAI211_X1 U15004 ( .C1(n15498), .C2(n18562), .A(n13265), .B(n13264), .ZN(
        n13266) );
  AOI21_X1 U15005 ( .B1(n15504), .B2(n18551), .A(n13266), .ZN(n13300) );
  MUX2_X1 U15006 ( .A(n13893), .B(P2_EBX_REG_2__SCAN_IN), .S(n13989), .Z(
        n13679) );
  INV_X1 U15007 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U15008 ( .A1(n14411), .A2(n14409), .ZN(n13270) );
  MUX2_X1 U15009 ( .A(n13908), .B(n13270), .S(n13989), .Z(n13680) );
  MUX2_X1 U15010 ( .A(n13272), .B(n13271), .S(n13989), .Z(n13673) );
  MUX2_X1 U15011 ( .A(n13274), .B(n13273), .S(n13989), .Z(n13688) );
  MUX2_X1 U15012 ( .A(n13714), .B(P2_EBX_REG_5__SCAN_IN), .S(n13989), .Z(
        n13717) );
  MUX2_X1 U15013 ( .A(n13748), .B(n14618), .S(n13989), .Z(n13756) );
  AND2_X2 U15014 ( .A1(n13757), .A2(n13756), .ZN(n13761) );
  INV_X1 U15015 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13277) );
  MUX2_X1 U15016 ( .A(n13277), .B(n13276), .S(n13820), .Z(n13760) );
  NOR2_X1 U15017 ( .A1(n13820), .A2(n13278), .ZN(n13763) );
  NAND2_X1 U15018 ( .A1(n13989), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13768) );
  NOR2_X1 U15019 ( .A1(n13820), .A2(n13279), .ZN(n13772) );
  NOR2_X1 U15020 ( .A1(n13820), .A2(n13280), .ZN(n13765) );
  OR2_X2 U15021 ( .A1(n13774), .A2(n13765), .ZN(n13786) );
  NOR2_X1 U15022 ( .A1(n13820), .A2(n13281), .ZN(n13785) );
  NOR2_X4 U15023 ( .A1(n13786), .A2(n13785), .ZN(n13796) );
  NAND2_X1 U15024 ( .A1(n13989), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13795) );
  NOR2_X1 U15025 ( .A1(n13820), .A2(n13282), .ZN(n13791) );
  NOR2_X1 U15026 ( .A1(n13820), .A2(n13283), .ZN(n13798) );
  NAND2_X1 U15027 ( .A1(n13989), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U15028 ( .A1(n13989), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13804) );
  NOR2_X1 U15029 ( .A1(n13820), .A2(n13284), .ZN(n13814) );
  NOR2_X1 U15030 ( .A1(n13820), .A2(n13285), .ZN(n13809) );
  NAND2_X1 U15031 ( .A1(n13989), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13789) );
  AND2_X2 U15032 ( .A1(n13811), .A2(n13789), .ZN(n13844) );
  OAI21_X1 U15033 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(P2_EBX_REG_22__SCAN_IN), 
        .A(n13989), .ZN(n13286) );
  NOR2_X1 U15034 ( .A1(n13820), .A2(n13287), .ZN(n13852) );
  INV_X1 U15035 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n13288) );
  NOR2_X1 U15036 ( .A1(n13820), .A2(n13288), .ZN(n13594) );
  INV_X1 U15037 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n13289) );
  NOR2_X1 U15038 ( .A1(n13820), .A2(n13289), .ZN(n13860) );
  NAND2_X1 U15039 ( .A1(n13989), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n13863) );
  NAND2_X1 U15040 ( .A1(n13864), .A2(n13863), .ZN(n13858) );
  NOR2_X1 U15041 ( .A1(n13820), .A2(n13290), .ZN(n13857) );
  NOR2_X1 U15042 ( .A1(n13820), .A2(n13291), .ZN(n13868) );
  NAND2_X1 U15043 ( .A1(n13989), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U15044 ( .A1(n13878), .A2(n13879), .ZN(n13988) );
  INV_X1 U15045 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13292) );
  NOR2_X1 U15046 ( .A1(n13820), .A2(n13292), .ZN(n13293) );
  XNOR2_X1 U15047 ( .A(n13988), .B(n13293), .ZN(n13882) );
  INV_X1 U15048 ( .A(n13882), .ZN(n13298) );
  INV_X1 U15049 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16091) );
  NOR2_X1 U15050 ( .A1(n13294), .A2(n16091), .ZN(n13295) );
  AND2_X1 U15051 ( .A1(n13268), .A2(n13295), .ZN(n13296) );
  INV_X1 U15052 ( .A(n13303), .ZN(n13304) );
  XNOR2_X1 U15053 ( .A(n13343), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15738) );
  AOI22_X1 U15054 ( .A1(n13306), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13305), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13311) );
  AOI22_X1 U15055 ( .A1(n13307), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U15056 ( .A1(n14448), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U15057 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13308) );
  NAND4_X1 U15058 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13319) );
  AOI22_X1 U15059 ( .A1(n11582), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11711), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U15060 ( .A1(n13313), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13312), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U15061 ( .A1(n11589), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U15062 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13314) );
  NAND4_X1 U15063 ( .A1(n13317), .A2(n13316), .A3(n13315), .A4(n13314), .ZN(
        n13318) );
  NOR2_X1 U15064 ( .A1(n13319), .A2(n13318), .ZN(n13323) );
  NOR2_X1 U15065 ( .A1(n13321), .A2(n13320), .ZN(n13322) );
  XOR2_X1 U15066 ( .A(n13323), .B(n13322), .Z(n13327) );
  AOI21_X1 U15067 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n22008), .A(
        n13339), .ZN(n13325) );
  NAND2_X1 U15068 ( .A1(n12204), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13324) );
  OAI211_X1 U15069 ( .C1(n13327), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        n13328) );
  OAI21_X1 U15070 ( .B1(n11753), .B2(n15738), .A(n13328), .ZN(n13463) );
  AOI22_X1 U15071 ( .A1(n12204), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13329), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13330) );
  AND2_X1 U15072 ( .A1(n15260), .A2(n13471), .ZN(n13331) );
  NAND2_X1 U15073 ( .A1(n13591), .A2(n13331), .ZN(n13336) );
  AOI22_X1 U15074 ( .A1(n15729), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15720), .ZN(n13332) );
  INV_X1 U15075 ( .A(n13332), .ZN(n13334) );
  INV_X1 U15076 ( .A(DATAI_31_), .ZN(n14574) );
  NOR2_X1 U15077 ( .A1(n15724), .A2(n14574), .ZN(n13333) );
  NOR2_X1 U15078 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  NAND2_X1 U15079 ( .A1(n13336), .A2(n13335), .ZN(P1_U2873) );
  INV_X1 U15080 ( .A(n14117), .ZN(n13337) );
  NAND2_X1 U15081 ( .A1(n13337), .A2(n14314), .ZN(n14111) );
  NAND2_X1 U15082 ( .A1(n13339), .A2(n21683), .ZN(n16837) );
  NAND2_X1 U15083 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21687), .ZN(n16834) );
  INV_X1 U15084 ( .A(n16834), .ZN(n13340) );
  NAND2_X1 U15085 ( .A1(n13340), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13341) );
  OR2_X2 U15086 ( .A1(n13585), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21616) );
  OAI211_X1 U15087 ( .C1(n16839), .C2(n16837), .A(n13341), .B(n21616), .ZN(
        n13342) );
  NAND2_X1 U15088 ( .A1(n13343), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13345) );
  INV_X1 U15089 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13344) );
  XNOR2_X1 U15090 ( .A(n13345), .B(n13344), .ZN(n14721) );
  NOR2_X1 U15091 ( .A1(n14721), .A2(n16839), .ZN(n13346) );
  NAND2_X1 U15092 ( .A1(n13591), .A2(n21661), .ZN(n13460) );
  NAND2_X1 U15093 ( .A1(n13347), .A2(n11553), .ZN(n13360) );
  OAI22_X1 U15094 ( .A1(n14321), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n13464), .ZN(n13470) );
  INV_X1 U15095 ( .A(n13360), .ZN(n13349) );
  NAND2_X1 U15096 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13350) );
  NAND2_X1 U15097 ( .A1(n13352), .A2(n13351), .ZN(n13355) );
  INV_X1 U15098 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14876) );
  NAND2_X1 U15099 ( .A1(n15446), .A2(n14876), .ZN(n13354) );
  NAND2_X1 U15100 ( .A1(n13360), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13353) );
  MUX2_X1 U15101 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13357) );
  NAND3_X1 U15102 ( .A1(n15446), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n13464), .ZN(n13356) );
  AND3_X1 U15103 ( .A1(n13357), .A2(n13425), .A3(n13356), .ZN(n14507) );
  MUX2_X1 U15104 ( .A(n13422), .B(n15446), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13359) );
  OAI21_X1 U15105 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14321), .A(
        n13359), .ZN(n14532) );
  MUX2_X1 U15106 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13363) );
  NAND2_X1 U15107 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13361) );
  AND2_X1 U15108 ( .A1(n13425), .A2(n13361), .ZN(n13362) );
  NAND2_X1 U15109 ( .A1(n13363), .A2(n13362), .ZN(n14705) );
  NAND2_X1 U15110 ( .A1(n14706), .A2(n14705), .ZN(n19905) );
  INV_X1 U15111 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U15112 ( .A1(n13432), .A2(n19910), .ZN(n13367) );
  INV_X1 U15113 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21365) );
  NAND2_X1 U15114 ( .A1(n14356), .A2(n19910), .ZN(n13365) );
  OAI211_X1 U15115 ( .C1(n13364), .C2(n21365), .A(n13365), .B(n13360), .ZN(
        n13366) );
  NAND2_X1 U15116 ( .A1(n13367), .A2(n13366), .ZN(n19904) );
  INV_X1 U15117 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19903) );
  NAND2_X1 U15118 ( .A1(n13432), .A2(n19903), .ZN(n13370) );
  INV_X1 U15119 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21377) );
  NAND2_X1 U15120 ( .A1(n14356), .A2(n19903), .ZN(n13368) );
  OAI211_X1 U15121 ( .C1(n13364), .C2(n21377), .A(n13368), .B(n13360), .ZN(
        n13369) );
  AND2_X1 U15122 ( .A1(n13370), .A2(n13369), .ZN(n19896) );
  MUX2_X1 U15123 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13373) );
  NAND2_X1 U15124 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13371) );
  AND2_X1 U15125 ( .A1(n13425), .A2(n13371), .ZN(n13372) );
  NAND2_X1 U15126 ( .A1(n13373), .A2(n13372), .ZN(n19897) );
  NAND2_X1 U15127 ( .A1(n19896), .A2(n19897), .ZN(n13374) );
  MUX2_X1 U15128 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13377) );
  NAND2_X1 U15129 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13375) );
  AND2_X1 U15130 ( .A1(n13425), .A2(n13375), .ZN(n13376) );
  NAND2_X1 U15131 ( .A1(n13377), .A2(n13376), .ZN(n15086) );
  INV_X1 U15132 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15091) );
  NAND2_X1 U15133 ( .A1(n13432), .A2(n15091), .ZN(n13380) );
  INV_X1 U15134 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21398) );
  NAND2_X1 U15135 ( .A1(n14356), .A2(n15091), .ZN(n13378) );
  OAI211_X1 U15136 ( .C1(n13364), .C2(n21398), .A(n13378), .B(n13360), .ZN(
        n13379) );
  AND2_X1 U15137 ( .A1(n13380), .A2(n13379), .ZN(n15087) );
  AND2_X1 U15138 ( .A1(n15086), .A2(n15087), .ZN(n13381) );
  NAND2_X1 U15139 ( .A1(n19899), .A2(n13381), .ZN(n19893) );
  INV_X1 U15140 ( .A(n13436), .ZN(n13382) );
  INV_X1 U15141 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21566) );
  NAND2_X1 U15142 ( .A1(n13382), .A2(n21566), .ZN(n13386) );
  INV_X1 U15143 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19936) );
  NAND2_X1 U15144 ( .A1(n13360), .A2(n19936), .ZN(n13384) );
  NAND2_X1 U15145 ( .A1(n14356), .A2(n21566), .ZN(n13383) );
  NAND3_X1 U15146 ( .A1(n13384), .A2(n15446), .A3(n13383), .ZN(n13385) );
  INV_X1 U15147 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21417) );
  NAND2_X1 U15148 ( .A1(n21417), .A2(n13439), .ZN(n13388) );
  MUX2_X1 U15149 ( .A(n13422), .B(n15446), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13387) );
  NAND2_X1 U15150 ( .A1(n13388), .A2(n13387), .ZN(n15199) );
  INV_X1 U15151 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U15152 ( .A1(n13432), .A2(n15271), .ZN(n13391) );
  NAND2_X1 U15153 ( .A1(n14356), .A2(n15271), .ZN(n13389) );
  OAI211_X1 U15154 ( .C1(n13364), .C2(n13552), .A(n13389), .B(n13360), .ZN(
        n13390) );
  INV_X1 U15155 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U15156 ( .A1(n13360), .A2(n13559), .ZN(n13393) );
  INV_X1 U15157 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21581) );
  NAND2_X1 U15158 ( .A1(n14356), .A2(n21581), .ZN(n13392) );
  NAND3_X1 U15159 ( .A1(n13393), .A2(n15446), .A3(n13392), .ZN(n13394) );
  OAI21_X1 U15160 ( .B1(n13436), .B2(P1_EBX_REG_12__SCAN_IN), .A(n13394), .ZN(
        n19890) );
  NAND2_X1 U15161 ( .A1(n15267), .A2(n19890), .ZN(n13395) );
  MUX2_X1 U15162 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13398) );
  NAND2_X1 U15163 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13396) );
  AND2_X1 U15164 ( .A1(n13425), .A2(n13396), .ZN(n13397) );
  NAND2_X1 U15165 ( .A1(n13398), .A2(n13397), .ZN(n15232) );
  INV_X1 U15166 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15255) );
  NAND2_X1 U15167 ( .A1(n13432), .A2(n15255), .ZN(n13401) );
  INV_X1 U15168 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16005) );
  NAND2_X1 U15169 ( .A1(n14356), .A2(n15255), .ZN(n13399) );
  OAI211_X1 U15170 ( .C1(n13364), .C2(n16005), .A(n13399), .B(n13360), .ZN(
        n13400) );
  MUX2_X1 U15171 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13403) );
  NAND2_X1 U15172 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13402) );
  INV_X1 U15173 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U15174 ( .A1(n13432), .A2(n13404), .ZN(n13407) );
  INV_X1 U15175 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U15176 ( .A1(n14356), .A2(n13404), .ZN(n13405) );
  OAI211_X1 U15177 ( .C1(n13364), .C2(n13558), .A(n13405), .B(n13360), .ZN(
        n13406) );
  NAND2_X1 U15178 ( .A1(n13407), .A2(n13406), .ZN(n15297) );
  MUX2_X1 U15179 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13410) );
  NAND2_X1 U15180 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13408) );
  AND2_X1 U15181 ( .A1(n13425), .A2(n13408), .ZN(n13409) );
  NAND2_X1 U15182 ( .A1(n13410), .A2(n13409), .ZN(n15653) );
  MUX2_X1 U15183 ( .A(n13422), .B(n15446), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13412) );
  INV_X1 U15184 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U15185 ( .A1(n13439), .A2(n15985), .ZN(n13411) );
  MUX2_X1 U15186 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13414) );
  NAND2_X1 U15187 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13413) );
  INV_X1 U15188 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15639) );
  NAND2_X1 U15189 ( .A1(n13432), .A2(n15639), .ZN(n13417) );
  INV_X1 U15190 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21456) );
  NAND2_X1 U15191 ( .A1(n14356), .A2(n15639), .ZN(n13415) );
  OAI211_X1 U15192 ( .C1(n13364), .C2(n21456), .A(n13415), .B(n13360), .ZN(
        n13416) );
  NAND2_X1 U15193 ( .A1(n13417), .A2(n13416), .ZN(n15584) );
  INV_X1 U15194 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U15195 ( .A1(n13360), .A2(n13418), .ZN(n13420) );
  INV_X1 U15196 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21650) );
  NAND2_X1 U15197 ( .A1(n14356), .A2(n21650), .ZN(n13419) );
  NAND3_X1 U15198 ( .A1(n13420), .A2(n15446), .A3(n13419), .ZN(n13421) );
  OAI21_X1 U15199 ( .B1(n13436), .B2(P1_EBX_REG_22__SCAN_IN), .A(n13421), .ZN(
        n15636) );
  MUX2_X1 U15200 ( .A(n13422), .B(n15446), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13423) );
  OAI21_X1 U15201 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14321), .A(
        n13423), .ZN(n15577) );
  MUX2_X1 U15202 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13426) );
  NAND2_X1 U15203 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13424) );
  INV_X1 U15204 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15623) );
  NAND2_X1 U15205 ( .A1(n13432), .A2(n15623), .ZN(n13429) );
  INV_X1 U15206 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15947) );
  NAND2_X1 U15207 ( .A1(n14356), .A2(n15623), .ZN(n13427) );
  OAI211_X1 U15208 ( .C1(n13364), .C2(n15947), .A(n13427), .B(n13360), .ZN(
        n13428) );
  NAND2_X1 U15209 ( .A1(n13429), .A2(n13428), .ZN(n15556) );
  INV_X1 U15210 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15779) );
  NAND2_X1 U15211 ( .A1(n13360), .A2(n15779), .ZN(n13430) );
  OAI211_X1 U15212 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n13464), .A(n13430), .B(
        n15446), .ZN(n13431) );
  OAI21_X1 U15213 ( .B1(n13436), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13431), .ZN(
        n15544) );
  INV_X1 U15214 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U15215 ( .A1(n13432), .A2(n15621), .ZN(n13435) );
  INV_X1 U15216 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U15217 ( .A1(n14356), .A2(n15621), .ZN(n13433) );
  OAI211_X1 U15218 ( .C1(n13364), .C2(n15757), .A(n13433), .B(n13360), .ZN(
        n13434) );
  NAND2_X1 U15219 ( .A1(n13435), .A2(n13434), .ZN(n15530) );
  MUX2_X1 U15220 ( .A(n13436), .B(n13360), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13438) );
  NAND2_X1 U15221 ( .A1(n13464), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13437) );
  INV_X1 U15222 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15618) );
  AND2_X1 U15223 ( .A1(n14356), .A2(n15618), .ZN(n13440) );
  INV_X1 U15224 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15913) );
  AOI21_X1 U15225 ( .B1(n13439), .B2(n15913), .A(n13440), .ZN(n13468) );
  MUX2_X1 U15226 ( .A(n13440), .B(n13468), .S(n15446), .Z(n15510) );
  NAND2_X1 U15227 ( .A1(n15519), .A2(n15510), .ZN(n15509) );
  MUX2_X1 U15228 ( .A(n13470), .B(n15446), .S(n15509), .Z(n13442) );
  OAI22_X1 U15229 ( .A1(n14321), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n13464), .ZN(n13441) );
  NOR2_X1 U15230 ( .A1(n15450), .A2(n11018), .ZN(n13453) );
  INV_X1 U15231 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15616) );
  AOI21_X1 U15232 ( .B1(n21716), .B2(n21936), .A(n15616), .ZN(n13443) );
  AND2_X1 U15233 ( .A1(n13348), .A2(n13443), .ZN(n13444) );
  INV_X1 U15234 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n19838) );
  INV_X1 U15235 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21576) );
  NAND4_X1 U15236 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_14__SCAN_IN), .A4(P1_REIP_REG_17__SCAN_IN), .ZN(n13445) );
  NOR3_X1 U15237 ( .A1(n19838), .A2(n21576), .A3(n13445), .ZN(n13446) );
  AND4_X1 U15238 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(n13446), .ZN(n21626) );
  NAND2_X1 U15239 ( .A1(n21626), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15590) );
  INV_X1 U15240 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n19842) );
  OR2_X1 U15241 ( .A1(n15590), .A2(n19842), .ZN(n21639) );
  INV_X1 U15242 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21635) );
  NOR2_X1 U15243 ( .A1(n21639), .A2(n21635), .ZN(n15560) );
  NAND4_X1 U15244 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n21494)
         );
  INV_X1 U15245 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21506) );
  NOR2_X1 U15246 ( .A1(n21494), .A2(n21506), .ZN(n21508) );
  NAND2_X1 U15247 ( .A1(n21508), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21518) );
  INV_X1 U15248 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21529) );
  NOR2_X1 U15249 ( .A1(n21518), .A2(n21529), .ZN(n21530) );
  NAND2_X1 U15250 ( .A1(n21530), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21540) );
  INV_X1 U15251 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21552) );
  NOR2_X1 U15252 ( .A1(n21540), .A2(n21552), .ZN(n21563) );
  NAND2_X1 U15253 ( .A1(n21563), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n21561) );
  INV_X1 U15254 ( .A(n21726), .ZN(n14118) );
  OAI21_X1 U15255 ( .B1(n13348), .B2(n14118), .A(n21716), .ZN(n14301) );
  NOR2_X1 U15256 ( .A1(n14301), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13451) );
  NAND2_X1 U15257 ( .A1(n15560), .A2(n21625), .ZN(n15573) );
  INV_X1 U15258 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n19846) );
  NOR2_X1 U15259 ( .A1(n15573), .A2(n19846), .ZN(n21656) );
  NAND2_X1 U15260 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n21656), .ZN(n15561) );
  INV_X1 U15261 ( .A(n15561), .ZN(n13448) );
  NAND3_X1 U15262 ( .A1(n13448), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_26__SCAN_IN), .ZN(n15552) );
  INV_X1 U15263 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n19851) );
  NOR2_X1 U15264 ( .A1(n15552), .A2(n19851), .ZN(n15529) );
  NAND2_X1 U15265 ( .A1(n15529), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15516) );
  INV_X1 U15266 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n19857) );
  NOR2_X1 U15267 ( .A1(n15516), .A2(n19857), .ZN(n15438) );
  AND2_X1 U15268 ( .A1(n15438), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U15269 ( .A1(n21539), .A2(n15559), .ZN(n21594) );
  NOR2_X1 U15270 ( .A1(n13449), .A2(n21601), .ZN(n15437) );
  INV_X1 U15271 ( .A(n13449), .ZN(n13455) );
  AND2_X1 U15272 ( .A1(n13348), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13450) );
  NOR2_X1 U15273 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  AOI22_X1 U15274 ( .A1(n21651), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21652), .ZN(n13454) );
  OAI21_X1 U15275 ( .B1(n13455), .B2(P1_REIP_REG_31__SCAN_IN), .A(n13454), 
        .ZN(n13456) );
  AOI21_X1 U15276 ( .B1(n15437), .B2(P1_REIP_REG_31__SCAN_IN), .A(n13456), 
        .ZN(n13457) );
  NAND2_X1 U15277 ( .A1(n13460), .A2(n13459), .ZN(P1_U2809) );
  INV_X1 U15278 ( .A(n15740), .ZN(n15445) );
  INV_X1 U15279 ( .A(n12273), .ZN(n14225) );
  NOR2_X1 U15280 ( .A1(n14225), .A2(n11558), .ZN(n14240) );
  NAND2_X1 U15281 ( .A1(n14240), .A2(n14356), .ZN(n14329) );
  INV_X1 U15282 ( .A(n14310), .ZN(n14305) );
  NAND2_X2 U15283 ( .A1(n14578), .A2(n19911), .ZN(n15659) );
  INV_X1 U15284 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15442) );
  NOR2_X1 U15285 ( .A1(n19911), .A2(n15442), .ZN(n13473) );
  AOI22_X1 U15286 ( .A1(n15509), .A2(n13364), .B1(n13468), .B2(n15519), .ZN(
        n13469) );
  INV_X1 U15287 ( .A(n15657), .ZN(n13472) );
  NAND2_X1 U15288 ( .A1(n13484), .A2(n13483), .ZN(n13496) );
  INV_X1 U15289 ( .A(n13474), .ZN(n13495) );
  XNOR2_X1 U15290 ( .A(n13496), .B(n13495), .ZN(n13475) );
  AOI21_X1 U15291 ( .B1(n13475), .B2(n14214), .A(n13477), .ZN(n13476) );
  INV_X1 U15292 ( .A(n13521), .ZN(n13481) );
  INV_X1 U15293 ( .A(n14214), .ZN(n21291) );
  INV_X1 U15294 ( .A(n13477), .ZN(n13478) );
  OAI21_X1 U15295 ( .B1(n21291), .B2(n13483), .A(n13478), .ZN(n13479) );
  INV_X1 U15296 ( .A(n13479), .ZN(n13480) );
  OAI211_X1 U15297 ( .C1(n13484), .C2(n13483), .A(n14214), .B(n13496), .ZN(
        n13485) );
  INV_X1 U15298 ( .A(n13485), .ZN(n13487) );
  NOR2_X1 U15299 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  XNOR2_X1 U15300 ( .A(n14284), .B(n13490), .ZN(n14354) );
  NAND2_X1 U15301 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14355) );
  INV_X1 U15302 ( .A(n13490), .ZN(n13491) );
  OR2_X1 U15303 ( .A1(n14284), .A2(n13491), .ZN(n13492) );
  INV_X1 U15304 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21336) );
  XNOR2_X1 U15305 ( .A(n13493), .B(n21336), .ZN(n14621) );
  NAND2_X1 U15306 ( .A1(n14620), .A2(n14621), .ZN(n14622) );
  NAND2_X1 U15307 ( .A1(n13493), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13494) );
  INV_X1 U15308 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21346) );
  OR2_X1 U15309 ( .A1(n14521), .A2(n13481), .ZN(n13500) );
  NAND2_X1 U15310 ( .A1(n13496), .A2(n13495), .ZN(n13504) );
  INV_X1 U15311 ( .A(n13503), .ZN(n13497) );
  XNOR2_X1 U15312 ( .A(n13504), .B(n13497), .ZN(n13498) );
  NAND2_X1 U15313 ( .A1(n13498), .A2(n14214), .ZN(n13499) );
  NAND2_X1 U15314 ( .A1(n13500), .A2(n13499), .ZN(n14751) );
  NAND2_X1 U15315 ( .A1(n13501), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13502) );
  NAND2_X1 U15316 ( .A1(n19914), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13508) );
  NAND2_X1 U15317 ( .A1(n13504), .A2(n13503), .ZN(n13513) );
  XNOR2_X1 U15318 ( .A(n13513), .B(n13511), .ZN(n13505) );
  AND2_X1 U15319 ( .A1(n13505), .A2(n14214), .ZN(n13506) );
  AOI21_X1 U15320 ( .B1(n13507), .B2(n13521), .A(n13506), .ZN(n19912) );
  INV_X1 U15321 ( .A(n19914), .ZN(n13510) );
  INV_X1 U15322 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13509) );
  INV_X1 U15323 ( .A(n13511), .ZN(n13512) );
  OR2_X1 U15324 ( .A1(n13513), .A2(n13512), .ZN(n13522) );
  XNOR2_X1 U15325 ( .A(n13522), .B(n13523), .ZN(n13514) );
  NAND2_X1 U15326 ( .A1(n13514), .A2(n14214), .ZN(n13515) );
  OAI21_X1 U15327 ( .B1(n13516), .B2(n13481), .A(n13515), .ZN(n13518) );
  XNOR2_X1 U15328 ( .A(n13518), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19920) );
  INV_X1 U15329 ( .A(n19920), .ZN(n13517) );
  NAND2_X1 U15330 ( .A1(n13518), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13519) );
  NAND2_X1 U15331 ( .A1(n19918), .A2(n13519), .ZN(n19924) );
  NAND3_X1 U15332 ( .A1(n13542), .A2(n13521), .A3(n13520), .ZN(n13527) );
  INV_X1 U15333 ( .A(n13522), .ZN(n13524) );
  NAND2_X1 U15334 ( .A1(n13524), .A2(n13523), .ZN(n13531) );
  XNOR2_X1 U15335 ( .A(n13531), .B(n13532), .ZN(n13525) );
  NAND2_X1 U15336 ( .A1(n13525), .A2(n14214), .ZN(n13526) );
  NAND2_X1 U15337 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  XNOR2_X1 U15338 ( .A(n13528), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19923) );
  OR2_X1 U15339 ( .A1(n13528), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13529) );
  INV_X1 U15340 ( .A(n13531), .ZN(n13533) );
  NAND2_X1 U15341 ( .A1(n13533), .A2(n13532), .ZN(n13545) );
  XNOR2_X1 U15342 ( .A(n13545), .B(n13543), .ZN(n13534) );
  NAND2_X1 U15343 ( .A1(n13534), .A2(n14214), .ZN(n13535) );
  XNOR2_X1 U15344 ( .A(n13537), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19932) );
  NAND2_X1 U15345 ( .A1(n13537), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13538) );
  INV_X1 U15346 ( .A(n13539), .ZN(n13540) );
  NAND2_X1 U15347 ( .A1(n14214), .A2(n13543), .ZN(n13544) );
  OR2_X1 U15348 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  NAND2_X1 U15349 ( .A1(n19950), .A2(n13546), .ZN(n13548) );
  XNOR2_X1 U15350 ( .A(n13548), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15241) );
  XNOR2_X1 U15351 ( .A(n19950), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15871) );
  NAND2_X1 U15352 ( .A1(n19950), .A2(n21398), .ZN(n13551) );
  INV_X1 U15353 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U15354 ( .A1(n19950), .A2(n13552), .ZN(n13553) );
  NAND2_X1 U15355 ( .A1(n19960), .A2(n13553), .ZN(n15861) );
  NAND3_X1 U15356 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13554) );
  NOR2_X2 U15357 ( .A1(n19956), .A2(n13555), .ZN(n15835) );
  INV_X1 U15358 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16000) );
  AND3_X1 U15359 ( .A1(n16005), .A2(n13558), .A3(n16000), .ZN(n13556) );
  INV_X1 U15360 ( .A(n13557), .ZN(n13563) );
  NAND2_X1 U15361 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21424) );
  NOR2_X1 U15362 ( .A1(n21424), .A2(n13558), .ZN(n21427) );
  OR2_X1 U15363 ( .A1(n19950), .A2(n13559), .ZN(n15859) );
  NOR2_X1 U15364 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13560) );
  OR2_X1 U15365 ( .A1(n19950), .A2(n13560), .ZN(n15857) );
  AND2_X1 U15366 ( .A1(n15859), .A2(n15857), .ZN(n15832) );
  INV_X1 U15367 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13561) );
  OR2_X1 U15368 ( .A1(n19950), .A2(n13561), .ZN(n13562) );
  AND2_X1 U15369 ( .A1(n19960), .A2(n13562), .ZN(n15833) );
  NAND3_X1 U15370 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15977) );
  INV_X1 U15371 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15810) );
  NOR2_X1 U15372 ( .A1(n15977), .A2(n15810), .ZN(n13564) );
  INV_X1 U15373 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13565) );
  NAND4_X1 U15374 ( .A1(n21456), .A2(n13565), .A3(n15985), .A4(n15810), .ZN(
        n13566) );
  INV_X1 U15375 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15953) );
  INV_X1 U15376 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15959) );
  NAND3_X1 U15377 ( .A1(n15953), .A2(n15947), .A3(n15959), .ZN(n15755) );
  AND2_X1 U15378 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15944) );
  NAND2_X1 U15379 ( .A1(n15944), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15886) );
  NAND2_X1 U15380 ( .A1(n19950), .A2(n15886), .ZN(n15777) );
  NAND3_X1 U15381 ( .A1(n15776), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15777), .ZN(n13568) );
  AND2_X1 U15382 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15909) );
  NOR2_X1 U15383 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15732) );
  AND2_X1 U15384 ( .A1(n19950), .A2(n15913), .ZN(n15742) );
  XNOR2_X1 U15385 ( .A(n19950), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13569) );
  INV_X1 U15386 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15903) );
  NAND2_X1 U15387 ( .A1(n19950), .A2(n15903), .ZN(n13574) );
  NAND3_X1 U15388 ( .A1(n13573), .A2(n13569), .A3(n13574), .ZN(n13579) );
  NOR2_X1 U15389 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13571) );
  INV_X1 U15390 ( .A(n13569), .ZN(n13570) );
  NOR2_X1 U15391 ( .A1(n19950), .A2(n15913), .ZN(n15743) );
  INV_X1 U15392 ( .A(n13574), .ZN(n13575) );
  AOI211_X1 U15393 ( .C1(n10972), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15743), .B(n13575), .ZN(n13576) );
  OR2_X1 U15394 ( .A1(n13576), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13577) );
  NAND3_X1 U15395 ( .A1(n13579), .A2(n13578), .A3(n13577), .ZN(n15898) );
  NAND2_X1 U15396 ( .A1(n13583), .A2(n11574), .ZN(n13580) );
  AND2_X1 U15397 ( .A1(n13581), .A2(n13580), .ZN(n14227) );
  NAND2_X1 U15398 ( .A1(n11558), .A2(n11018), .ZN(n13582) );
  NAND2_X1 U15399 ( .A1(n14251), .A2(n13583), .ZN(n16817) );
  OR2_X2 U15400 ( .A1(n15898), .A2(n21667), .ZN(n13593) );
  NAND3_X1 U15401 ( .A1(n21683), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21680) );
  INV_X1 U15402 ( .A(n21680), .ZN(n13584) );
  NAND2_X1 U15403 ( .A1(n22015), .A2(n13585), .ZN(n21287) );
  NAND2_X1 U15404 ( .A1(n21287), .A2(n21683), .ZN(n13586) );
  NAND2_X1 U15405 ( .A1(n21683), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16829) );
  NAND2_X1 U15406 ( .A1(n21936), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13587) );
  AND2_X1 U15407 ( .A1(n16829), .A2(n13587), .ZN(n14290) );
  INV_X1 U15408 ( .A(n14290), .ZN(n13588) );
  INV_X1 U15409 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n19861) );
  NOR2_X1 U15410 ( .A1(n21616), .A2(n19861), .ZN(n15894) );
  AOI21_X1 U15411 ( .B1(n19976), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15894), .ZN(n13589) );
  OAI21_X1 U15412 ( .B1(n19982), .B2(n14721), .A(n13589), .ZN(n13590) );
  AOI21_X1 U15413 ( .B1(n13591), .B2(n19979), .A(n13590), .ZN(n13592) );
  NAND2_X1 U15414 ( .A1(n13593), .A2(n13592), .ZN(P1_U2968) );
  INV_X1 U15415 ( .A(n13594), .ZN(n13595) );
  XNOR2_X1 U15416 ( .A(n13855), .B(n13595), .ZN(n18500) );
  NAND2_X1 U15417 ( .A1(n18500), .A2(n13276), .ZN(n16281) );
  NAND2_X1 U15418 ( .A1(n17132), .A2(n13606), .ZN(n13620) );
  INV_X1 U15419 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13599) );
  INV_X1 U15420 ( .A(n13620), .ZN(n13597) );
  INV_X1 U15421 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13598) );
  OAI22_X1 U15422 ( .A1(n19155), .A2(n13599), .B1(n19248), .B2(n13598), .ZN(
        n13605) );
  INV_X1 U15423 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13603) );
  INV_X1 U15424 ( .A(n13623), .ZN(n13600) );
  NAND2_X1 U15425 ( .A1(n13601), .A2(n11028), .ZN(n19192) );
  OAI22_X1 U15426 ( .A1(n13603), .A2(n19192), .B1(n19218), .B2(n13602), .ZN(
        n13604) );
  OR2_X1 U15427 ( .A1(n15161), .A2(n13606), .ZN(n13622) );
  INV_X1 U15428 ( .A(n13622), .ZN(n13607) );
  INV_X1 U15429 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13609) );
  INV_X1 U15430 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13608) );
  OAI22_X1 U15431 ( .A1(n19135), .A2(n13609), .B1(n19231), .B2(n13608), .ZN(
        n13614) );
  INV_X1 U15432 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13612) );
  INV_X1 U15433 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13611) );
  OAI22_X1 U15434 ( .A1(n19144), .A2(n13612), .B1(n17047), .B2(n13611), .ZN(
        n13613) );
  INV_X1 U15435 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13618) );
  INV_X1 U15436 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13617) );
  BUF_X2 U15437 ( .A(n13621), .Z(n14921) );
  AND2_X2 U15438 ( .A1(n13632), .A2(n14921), .ZN(n13698) );
  AND2_X1 U15439 ( .A1(n13625), .A2(n13624), .ZN(n13629) );
  NAND2_X1 U15440 ( .A1(n19334), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13628) );
  NAND2_X1 U15441 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13627) );
  NAND3_X1 U15442 ( .A1(n13629), .A2(n13628), .A3(n13627), .ZN(n13636) );
  NOR2_X2 U15443 ( .A1(n13631), .A2(n14921), .ZN(n13699) );
  INV_X1 U15444 ( .A(n13632), .ZN(n13633) );
  AOI22_X1 U15445 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13699), .B1(
        n19178), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13634) );
  INV_X1 U15446 ( .A(n13634), .ZN(n13635) );
  INV_X1 U15447 ( .A(n13638), .ZN(n13639) );
  NAND2_X1 U15448 ( .A1(n13639), .A2(n19574), .ZN(n13640) );
  NAND2_X1 U15449 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13642) );
  INV_X1 U15450 ( .A(n19334), .ZN(n13652) );
  INV_X1 U15451 ( .A(n19144), .ZN(n13646) );
  NAND2_X1 U15452 ( .A1(n13646), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13650) );
  INV_X1 U15453 ( .A(n13698), .ZN(n13648) );
  INV_X1 U15454 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13647) );
  INV_X1 U15455 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13654) );
  INV_X1 U15456 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13653) );
  OAI22_X1 U15457 ( .A1(n19170), .A2(n13654), .B1(n19263), .B2(n13653), .ZN(
        n13658) );
  INV_X1 U15458 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13656) );
  INV_X1 U15459 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13655) );
  OAI22_X1 U15460 ( .A1(n13656), .A2(n19248), .B1(n17047), .B2(n13655), .ZN(
        n13657) );
  NOR2_X1 U15461 ( .A1(n13658), .A2(n13657), .ZN(n13666) );
  INV_X1 U15462 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13660) );
  INV_X1 U15463 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13659) );
  OAI22_X1 U15464 ( .A1(n19192), .A2(n13660), .B1(n19135), .B2(n13659), .ZN(
        n13664) );
  INV_X1 U15465 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13662) );
  INV_X1 U15466 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13661) );
  OAI22_X1 U15467 ( .A1(n19155), .A2(n13662), .B1(n19231), .B2(n13661), .ZN(
        n13663) );
  NOR2_X1 U15468 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  NOR2_X1 U15469 ( .A1(n16746), .A2(n13908), .ZN(n13667) );
  NAND2_X1 U15470 ( .A1(n19574), .A2(n13667), .ZN(n13903) );
  INV_X1 U15471 ( .A(n13668), .ZN(n13902) );
  NAND2_X1 U15472 ( .A1(n13903), .A2(n13902), .ZN(n13669) );
  NAND2_X1 U15473 ( .A1(n13671), .A2(n13670), .ZN(n13672) );
  XNOR2_X1 U15475 ( .A(n13674), .B(n13673), .ZN(n14964) );
  OAI21_X2 U15476 ( .B1(n14919), .B2(n13276), .A(n14964), .ZN(n14916) );
  NAND2_X1 U15477 ( .A1(n14916), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13684) );
  NAND3_X1 U15478 ( .A1(n13989), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n13675) );
  INV_X1 U15479 ( .A(n13676), .ZN(n13889) );
  MUX2_X1 U15480 ( .A(n13889), .B(n16746), .S(n13268), .Z(n13895) );
  MUX2_X1 U15481 ( .A(n13895), .B(n14411), .S(n13989), .Z(n16749) );
  NOR2_X1 U15482 ( .A1(n16749), .A2(n13904), .ZN(n13677) );
  NAND2_X1 U15483 ( .A1(n11394), .A2(n13677), .ZN(n13678) );
  XOR2_X1 U15484 ( .A(n11394), .B(n13677), .Z(n14086) );
  NAND2_X1 U15485 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14086), .ZN(
        n14085) );
  NAND2_X1 U15486 ( .A1(n13678), .A2(n14085), .ZN(n14155) );
  INV_X1 U15487 ( .A(n13679), .ZN(n13681) );
  XNOR2_X1 U15488 ( .A(n13681), .B(n13680), .ZN(n15097) );
  NOR2_X1 U15489 ( .A1(n14155), .A2(n15097), .ZN(n14154) );
  OR2_X1 U15490 ( .A1(n14154), .A2(n14159), .ZN(n13683) );
  NAND2_X1 U15491 ( .A1(n14155), .A2(n15097), .ZN(n13682) );
  AND2_X1 U15492 ( .A1(n13683), .A2(n13682), .ZN(n14914) );
  NAND2_X1 U15493 ( .A1(n13684), .A2(n14914), .ZN(n13687) );
  INV_X1 U15494 ( .A(n14916), .ZN(n13685) );
  NAND2_X1 U15495 ( .A1(n13685), .A2(n15062), .ZN(n13686) );
  OAI21_X1 U15496 ( .B1(n11074), .B2(n13688), .A(n13718), .ZN(n18303) );
  XNOR2_X1 U15497 ( .A(n18303), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15069) );
  NAND2_X1 U15498 ( .A1(n15068), .A2(n15069), .ZN(n15072) );
  INV_X1 U15499 ( .A(n18303), .ZN(n13689) );
  NAND2_X1 U15500 ( .A1(n13689), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13690) );
  NAND2_X1 U15501 ( .A1(n15072), .A2(n13690), .ZN(n15171) );
  INV_X1 U15502 ( .A(n13918), .ZN(n13691) );
  OAI22_X1 U15503 ( .A1(n13693), .A2(n19192), .B1(n19218), .B2(n13692), .ZN(
        n13697) );
  OAI22_X1 U15504 ( .A1(n19135), .A2(n13695), .B1(n19231), .B2(n13694), .ZN(
        n13696) );
  NOR2_X1 U15505 ( .A1(n13697), .A2(n13696), .ZN(n13713) );
  INV_X1 U15506 ( .A(n19263), .ZN(n19266) );
  INV_X1 U15507 ( .A(n17047), .ZN(n17040) );
  AOI22_X1 U15508 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19266), .B1(
        n17040), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U15509 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13698), .B1(
        n19178), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19309), .B1(
        n13699), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13702) );
  NAND2_X1 U15511 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13701) );
  NAND2_X1 U15512 ( .A1(n19334), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13700) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13705) );
  INV_X1 U15514 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13704) );
  OAI22_X1 U15515 ( .A1(n13705), .A2(n19170), .B1(n19144), .B2(n13704), .ZN(
        n13709) );
  INV_X1 U15516 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13707) );
  INV_X1 U15517 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13706) );
  OAI22_X1 U15518 ( .A1(n19155), .A2(n13707), .B1(n19248), .B2(n13706), .ZN(
        n13708) );
  NOR2_X1 U15519 ( .A1(n13709), .A2(n13708), .ZN(n13710) );
  NAND4_X1 U15520 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        n13716) );
  NAND2_X1 U15521 ( .A1(n13714), .A2(n19574), .ZN(n13715) );
  NAND2_X1 U15522 ( .A1(n13926), .A2(n13596), .ZN(n13719) );
  XNOR2_X1 U15523 ( .A(n13718), .B(n13717), .ZN(n18320) );
  NAND2_X1 U15524 ( .A1(n13719), .A2(n18320), .ZN(n13720) );
  INV_X1 U15525 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15178) );
  XNOR2_X1 U15526 ( .A(n13720), .B(n15178), .ZN(n15172) );
  NAND2_X1 U15527 ( .A1(n15171), .A2(n15172), .ZN(n15170) );
  NAND2_X1 U15528 ( .A1(n13720), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13721) );
  NAND2_X1 U15529 ( .A1(n15170), .A2(n13721), .ZN(n16715) );
  INV_X1 U15530 ( .A(n13722), .ZN(n13724) );
  NAND2_X1 U15531 ( .A1(n13724), .A2(n13723), .ZN(n13752) );
  INV_X1 U15532 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13726) );
  INV_X1 U15533 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13725) );
  OAI22_X1 U15534 ( .A1(n13726), .A2(n19218), .B1(n19192), .B2(n13725), .ZN(
        n13730) );
  INV_X1 U15535 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13728) );
  OAI22_X1 U15536 ( .A1(n19135), .A2(n13728), .B1(n19231), .B2(n13727), .ZN(
        n13729) );
  NOR2_X1 U15537 ( .A1(n13730), .A2(n13729), .ZN(n13747) );
  INV_X1 U15538 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13732) );
  INV_X1 U15539 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13731) );
  OAI22_X1 U15540 ( .A1(n19144), .A2(n13732), .B1(n19263), .B2(n13731), .ZN(
        n13733) );
  INV_X1 U15541 ( .A(n13733), .ZN(n13746) );
  AOI22_X1 U15542 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19309), .B1(
        n19178), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U15543 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13698), .B1(
        n13699), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U15544 ( .A1(n19334), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13735) );
  NAND2_X1 U15545 ( .A1(n19294), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13734) );
  INV_X1 U15546 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13739) );
  INV_X1 U15547 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13738) );
  OAI22_X1 U15548 ( .A1(n19155), .A2(n13739), .B1(n19248), .B2(n13738), .ZN(
        n13743) );
  INV_X1 U15549 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13741) );
  INV_X1 U15550 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13740) );
  OAI22_X1 U15551 ( .A1(n19170), .A2(n13741), .B1(n17047), .B2(n13740), .ZN(
        n13742) );
  NOR2_X1 U15552 ( .A1(n13743), .A2(n13742), .ZN(n13744) );
  NAND4_X1 U15553 ( .A1(n13747), .A2(n13746), .A3(n13745), .A4(n13744), .ZN(
        n13751) );
  INV_X1 U15554 ( .A(n13748), .ZN(n13749) );
  NAND2_X1 U15555 ( .A1(n13749), .A2(n19574), .ZN(n13750) );
  NAND2_X1 U15556 ( .A1(n13752), .A2(n13931), .ZN(n13755) );
  INV_X1 U15557 ( .A(n13752), .ZN(n13754) );
  NAND2_X1 U15558 ( .A1(n13754), .A2(n13753), .ZN(n13939) );
  NAND2_X1 U15559 ( .A1(n13755), .A2(n13939), .ZN(n13928) );
  XNOR2_X1 U15560 ( .A(n13757), .B(n13756), .ZN(n18331) );
  OAI21_X2 U15561 ( .B1(n13928), .B2(n13276), .A(n18331), .ZN(n13758) );
  INV_X1 U15562 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16719) );
  XNOR2_X1 U15563 ( .A(n13758), .B(n16719), .ZN(n16716) );
  NAND2_X1 U15564 ( .A1(n13758), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13759) );
  XNOR2_X1 U15565 ( .A(n13761), .B(n11155), .ZN(n18345) );
  INV_X1 U15566 ( .A(n13763), .ZN(n13764) );
  XNOR2_X1 U15567 ( .A(n13762), .B(n13764), .ZN(n15078) );
  INV_X1 U15568 ( .A(n16654), .ZN(n17074) );
  NOR2_X1 U15569 ( .A1(n17074), .A2(n14025), .ZN(n13778) );
  NAND2_X1 U15570 ( .A1(n13774), .A2(n13765), .ZN(n13766) );
  NAND2_X1 U15571 ( .A1(n13786), .A2(n13766), .ZN(n18374) );
  INV_X1 U15572 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16665) );
  OAI21_X1 U15573 ( .B1(n18374), .B2(n13596), .A(n16665), .ZN(n16658) );
  OR2_X1 U15574 ( .A1(n11079), .A2(n13768), .ZN(n13769) );
  NAND2_X1 U15575 ( .A1(n13767), .A2(n13769), .ZN(n18355) );
  OR2_X1 U15576 ( .A1(n18355), .A2(n13596), .ZN(n13781) );
  INV_X1 U15577 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U15578 ( .A1(n13781), .A2(n16698), .ZN(n16689) );
  INV_X1 U15579 ( .A(n18345), .ZN(n13770) );
  NAND2_X1 U15580 ( .A1(n13770), .A2(n16707), .ZN(n17073) );
  OAI211_X1 U15581 ( .C1(n16654), .C2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n16689), .B(n17073), .ZN(n13771) );
  INV_X1 U15582 ( .A(n13771), .ZN(n13776) );
  NAND2_X1 U15583 ( .A1(n13767), .A2(n13772), .ZN(n13773) );
  NAND2_X1 U15584 ( .A1(n13774), .A2(n13773), .ZN(n15044) );
  OR2_X1 U15585 ( .A1(n15044), .A2(n13596), .ZN(n13779) );
  INV_X1 U15586 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U15587 ( .A1(n13779), .A2(n13775), .ZN(n16675) );
  AND3_X1 U15588 ( .A1(n16658), .A2(n13776), .A3(n16675), .ZN(n13777) );
  INV_X1 U15589 ( .A(n13779), .ZN(n13780) );
  NAND2_X1 U15590 ( .A1(n13780), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16676) );
  INV_X1 U15591 ( .A(n13781), .ZN(n13782) );
  NAND2_X1 U15592 ( .A1(n13782), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16691) );
  NAND2_X1 U15593 ( .A1(n16676), .A2(n16691), .ZN(n16657) );
  NAND2_X1 U15594 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13783) );
  NOR2_X1 U15595 ( .A1(n18374), .A2(n13783), .ZN(n16659) );
  NOR2_X1 U15596 ( .A1(n16657), .A2(n16659), .ZN(n13784) );
  AND2_X1 U15597 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  OR2_X1 U15598 ( .A1(n13787), .A2(n13796), .ZN(n18383) );
  NAND2_X1 U15599 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13788) );
  NOR2_X1 U15600 ( .A1(n13811), .A2(n13789), .ZN(n13790) );
  OR2_X1 U15601 ( .A1(n13844), .A2(n13790), .ZN(n16074) );
  NOR2_X1 U15602 ( .A1(n16074), .A2(n13596), .ZN(n16363) );
  INV_X1 U15603 ( .A(n13791), .ZN(n13792) );
  XNOR2_X1 U15604 ( .A(n13793), .B(n13792), .ZN(n18411) );
  NAND2_X1 U15605 ( .A1(n18411), .A2(n13276), .ZN(n13794) );
  INV_X1 U15606 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18596) );
  NAND2_X1 U15607 ( .A1(n13794), .A2(n18596), .ZN(n17107) );
  XNOR2_X1 U15608 ( .A(n13796), .B(n11170), .ZN(n18401) );
  NAND2_X1 U15609 ( .A1(n18401), .A2(n13276), .ZN(n13797) );
  INV_X1 U15610 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16631) );
  NAND2_X1 U15611 ( .A1(n13797), .A2(n16631), .ZN(n16419) );
  AND2_X1 U15612 ( .A1(n17107), .A2(n16419), .ZN(n13802) );
  INV_X1 U15613 ( .A(n13798), .ZN(n13799) );
  XNOR2_X1 U15614 ( .A(n13800), .B(n13799), .ZN(n18429) );
  NAND2_X1 U15615 ( .A1(n18429), .A2(n13276), .ZN(n13801) );
  INV_X1 U15616 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16626) );
  NAND2_X1 U15617 ( .A1(n13801), .A2(n16626), .ZN(n16613) );
  NAND2_X1 U15618 ( .A1(n13802), .A2(n16613), .ZN(n14075) );
  OAI21_X1 U15619 ( .B1(n18383), .B2(n13596), .A(n16630), .ZN(n16645) );
  INV_X1 U15620 ( .A(n16645), .ZN(n13803) );
  NOR2_X1 U15621 ( .A1(n14075), .A2(n13803), .ZN(n13808) );
  INV_X1 U15622 ( .A(n13804), .ZN(n13805) );
  XNOR2_X1 U15623 ( .A(n13806), .B(n13805), .ZN(n18437) );
  NAND2_X1 U15624 ( .A1(n18437), .A2(n13276), .ZN(n13807) );
  INV_X1 U15625 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16593) );
  NAND2_X1 U15626 ( .A1(n13807), .A2(n16593), .ZN(n16405) );
  OAI211_X1 U15627 ( .C1(n16363), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n13808), .B(n16405), .ZN(n13818) );
  AND2_X1 U15628 ( .A1(n13810), .A2(n13809), .ZN(n13812) );
  OR2_X1 U15629 ( .A1(n13812), .A2(n13811), .ZN(n18463) );
  NOR2_X1 U15630 ( .A1(n18463), .A2(n13596), .ZN(n13828) );
  INV_X1 U15631 ( .A(n13828), .ZN(n13813) );
  INV_X1 U15632 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16565) );
  NAND2_X1 U15633 ( .A1(n13813), .A2(n16565), .ZN(n16382) );
  INV_X1 U15634 ( .A(n13814), .ZN(n13815) );
  XNOR2_X1 U15635 ( .A(n13816), .B(n13815), .ZN(n18450) );
  NAND2_X1 U15636 ( .A1(n18450), .A2(n13276), .ZN(n13817) );
  INV_X1 U15637 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16402) );
  NAND2_X1 U15638 ( .A1(n13817), .A2(n16402), .ZN(n16392) );
  NAND2_X1 U15639 ( .A1(n16382), .A2(n16392), .ZN(n16360) );
  NOR2_X1 U15640 ( .A1(n13818), .A2(n16360), .ZN(n13827) );
  NOR2_X1 U15641 ( .A1(n13820), .A2(n13819), .ZN(n13845) );
  XNOR2_X1 U15642 ( .A(n13844), .B(n13845), .ZN(n18480) );
  NAND2_X1 U15643 ( .A1(n18480), .A2(n13276), .ZN(n16366) );
  INV_X1 U15644 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U15645 ( .A1(n16366), .A2(n16345), .ZN(n13825) );
  INV_X1 U15646 ( .A(n13821), .ZN(n13822) );
  XNOR2_X1 U15647 ( .A(n13823), .B(n13822), .ZN(n16081) );
  NAND2_X1 U15648 ( .A1(n16081), .A2(n13276), .ZN(n13824) );
  XNOR2_X1 U15649 ( .A(n13824), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14077) );
  AND2_X1 U15650 ( .A1(n13825), .A2(n14077), .ZN(n13826) );
  NAND2_X1 U15651 ( .A1(n13828), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16383) );
  AND2_X1 U15652 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13829) );
  NAND2_X1 U15653 ( .A1(n18450), .A2(n13829), .ZN(n16391) );
  AND2_X1 U15654 ( .A1(n16383), .A2(n16391), .ZN(n16361) );
  NAND2_X1 U15655 ( .A1(n16363), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13838) );
  AND2_X1 U15656 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13830) );
  AND2_X1 U15657 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13831) );
  NAND2_X1 U15658 ( .A1(n16081), .A2(n13831), .ZN(n16358) );
  AND2_X1 U15659 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13832) );
  INV_X1 U15660 ( .A(n16420), .ZN(n13835) );
  AND2_X1 U15661 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13833) );
  NAND2_X1 U15662 ( .A1(n18429), .A2(n13833), .ZN(n16612) );
  AND2_X1 U15663 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13834) );
  NAND2_X1 U15664 ( .A1(n18411), .A2(n13834), .ZN(n17106) );
  NAND4_X1 U15665 ( .A1(n16358), .A2(n13835), .A3(n16612), .A4(n17106), .ZN(
        n13836) );
  NOR2_X1 U15666 ( .A1(n16406), .A2(n13836), .ZN(n13837) );
  NAND3_X1 U15667 ( .A1(n16361), .A2(n13838), .A3(n13837), .ZN(n13841) );
  INV_X1 U15668 ( .A(n16366), .ZN(n13839) );
  NAND2_X1 U15669 ( .A1(n13989), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n13848) );
  INV_X1 U15670 ( .A(n13844), .ZN(n13846) );
  NOR2_X1 U15671 ( .A1(n13846), .A2(n13845), .ZN(n13847) );
  XOR2_X1 U15672 ( .A(n13848), .B(n13847), .Z(n16046) );
  NAND2_X1 U15673 ( .A1(n16046), .A2(n13276), .ZN(n13849) );
  INV_X1 U15674 ( .A(n13849), .ZN(n13850) );
  NAND2_X1 U15675 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  NAND2_X1 U15676 ( .A1(n13855), .A2(n13854), .ZN(n18487) );
  NOR2_X1 U15677 ( .A1(n18487), .A2(n13596), .ZN(n13856) );
  XOR2_X1 U15678 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n13856), .Z(
        n16339) );
  INV_X1 U15679 ( .A(n16280), .ZN(n16283) );
  NAND2_X1 U15680 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  INV_X1 U15681 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16438) );
  INV_X1 U15682 ( .A(n13860), .ZN(n13861) );
  XNOR2_X1 U15683 ( .A(n13862), .B(n13861), .ZN(n18510) );
  NAND2_X1 U15684 ( .A1(n18510), .A2(n13276), .ZN(n13873) );
  INV_X1 U15685 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16489) );
  NAND2_X1 U15686 ( .A1(n13873), .A2(n16489), .ZN(n16314) );
  OAI211_X1 U15687 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16327), .A(
        n16288), .B(n16314), .ZN(n13867) );
  XNOR2_X1 U15688 ( .A(n13864), .B(n13863), .ZN(n18523) );
  INV_X1 U15689 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14026) );
  NOR3_X1 U15690 ( .A1(n18523), .A2(n13596), .A3(n14026), .ZN(n13874) );
  INV_X1 U15691 ( .A(n18523), .ZN(n13865) );
  AOI21_X1 U15692 ( .B1(n13865), .B2(n13276), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13866) );
  NOR2_X1 U15693 ( .A1(n13874), .A2(n13866), .ZN(n16284) );
  INV_X1 U15694 ( .A(n16284), .ZN(n16307) );
  INV_X1 U15695 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16448) );
  NAND2_X1 U15696 ( .A1(n16448), .A2(n16438), .ZN(n13871) );
  AND2_X1 U15697 ( .A1(n13872), .A2(n13871), .ZN(n13876) );
  NOR2_X1 U15698 ( .A1(n13873), .A2(n16489), .ZN(n16316) );
  NOR2_X1 U15699 ( .A1(n13874), .A2(n16316), .ZN(n16285) );
  INV_X1 U15700 ( .A(n16285), .ZN(n13875) );
  XOR2_X1 U15701 ( .A(n13879), .B(n13878), .Z(n18560) );
  AOI21_X1 U15702 ( .B1(n18560), .B2(n13276), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16268) );
  INV_X1 U15703 ( .A(n18560), .ZN(n13880) );
  INV_X1 U15704 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16443) );
  NOR2_X1 U15705 ( .A1(n13987), .A2(n16267), .ZN(n13885) );
  NAND2_X1 U15706 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13881) );
  NOR2_X1 U15707 ( .A1(n13882), .A2(n13881), .ZN(n13984) );
  INV_X1 U15708 ( .A(n13984), .ZN(n13883) );
  INV_X1 U15709 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15459) );
  OAI21_X1 U15710 ( .B1(n13882), .B2(n13596), .A(n15459), .ZN(n13986) );
  NAND2_X1 U15711 ( .A1(n13883), .A2(n13986), .ZN(n13884) );
  NAND2_X1 U15712 ( .A1(n13886), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13887) );
  NAND2_X1 U15713 ( .A1(n13887), .A2(n16769), .ZN(n16765) );
  INV_X1 U15714 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13888) );
  OAI21_X1 U15715 ( .B1(n12848), .B2(n16765), .A(n13888), .ZN(n17141) );
  NOR2_X1 U15716 ( .A1(n13890), .A2(n13889), .ZN(n13891) );
  NOR2_X1 U15717 ( .A1(n14833), .A2(n13891), .ZN(n13892) );
  MUX2_X1 U15718 ( .A(n17141), .B(n13892), .S(n14093), .Z(n18632) );
  NOR2_X1 U15719 ( .A1(n13955), .A2(n14822), .ZN(n13983) );
  NAND2_X1 U15720 ( .A1(n18632), .A2(n13983), .ZN(n13901) );
  OAI21_X1 U15721 ( .B1(n13895), .B2(n13894), .A(n13893), .ZN(n13896) );
  INV_X1 U15722 ( .A(n13896), .ZN(n13897) );
  NOR2_X1 U15723 ( .A1(n13898), .A2(n13897), .ZN(n13900) );
  NOR2_X1 U15724 ( .A1(n13900), .A2(n13899), .ZN(n14821) );
  NOR2_X1 U15725 ( .A1(n13955), .A2(n14820), .ZN(n14033) );
  NAND2_X1 U15726 ( .A1(n14821), .A2(n14033), .ZN(n13976) );
  NAND2_X1 U15727 ( .A1(n13901), .A2(n13976), .ZN(n14839) );
  NAND2_X1 U15728 ( .A1(n14919), .A2(n15062), .ZN(n13914) );
  XNOR2_X1 U15729 ( .A(n13903), .B(n13902), .ZN(n13910) );
  NOR2_X1 U15730 ( .A1(n13904), .A2(n13906), .ZN(n16744) );
  INV_X1 U15731 ( .A(n13908), .ZN(n13905) );
  NAND2_X1 U15732 ( .A1(n16744), .A2(n13905), .ZN(n13909) );
  NOR2_X1 U15733 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13906), .ZN(
        n13907) );
  XOR2_X1 U15734 ( .A(n13908), .B(n13907), .Z(n14088) );
  NAND2_X1 U15735 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14088), .ZN(
        n14087) );
  NAND2_X1 U15736 ( .A1(n13909), .A2(n14087), .ZN(n13911) );
  AND2_X1 U15737 ( .A1(n13910), .A2(n13911), .ZN(n14158) );
  NOR2_X1 U15738 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14158), .ZN(
        n13912) );
  NOR2_X1 U15739 ( .A1(n13911), .A2(n13910), .ZN(n14157) );
  OR2_X1 U15740 ( .A1(n13912), .A2(n14157), .ZN(n14917) );
  INV_X1 U15741 ( .A(n14917), .ZN(n13913) );
  NAND2_X1 U15742 ( .A1(n13914), .A2(n13913), .ZN(n13917) );
  INV_X1 U15743 ( .A(n14919), .ZN(n13915) );
  NAND2_X1 U15744 ( .A1(n13917), .A2(n13916), .ZN(n13922) );
  INV_X1 U15745 ( .A(n13919), .ZN(n13920) );
  XNOR2_X1 U15746 ( .A(n13922), .B(n13923), .ZN(n15057) );
  INV_X1 U15747 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U15748 ( .A1(n15057), .A2(n15174), .ZN(n15059) );
  INV_X1 U15749 ( .A(n13922), .ZN(n13924) );
  NAND2_X1 U15750 ( .A1(n13924), .A2(n13923), .ZN(n13925) );
  NAND2_X2 U15751 ( .A1(n15059), .A2(n13925), .ZN(n15169) );
  NAND2_X1 U15752 ( .A1(n13926), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15166) );
  NAND2_X1 U15753 ( .A1(n15169), .A2(n15166), .ZN(n13936) );
  INV_X1 U15754 ( .A(n13926), .ZN(n13927) );
  NAND2_X1 U15755 ( .A1(n13927), .A2(n15178), .ZN(n15167) );
  NAND2_X1 U15756 ( .A1(n13936), .A2(n15167), .ZN(n13929) );
  INV_X1 U15757 ( .A(n13928), .ZN(n13935) );
  INV_X1 U15758 ( .A(n15167), .ZN(n13930) );
  NOR2_X1 U15759 ( .A1(n15169), .A2(n13930), .ZN(n13932) );
  NAND2_X1 U15760 ( .A1(n16714), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13938) );
  NAND3_X1 U15761 ( .A1(n13936), .A2(n13935), .A3(n15167), .ZN(n13937) );
  XNOR2_X1 U15762 ( .A(n13939), .B(n13596), .ZN(n13940) );
  XNOR2_X1 U15763 ( .A(n13940), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16428) );
  NAND2_X1 U15764 ( .A1(n16429), .A2(n16428), .ZN(n13943) );
  INV_X1 U15765 ( .A(n13940), .ZN(n13941) );
  NAND2_X1 U15766 ( .A1(n13941), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13942) );
  NAND2_X1 U15767 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13945) );
  NAND3_X1 U15768 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18592) );
  NAND3_X1 U15769 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14074) );
  NOR2_X1 U15770 ( .A1(n18592), .A2(n14074), .ZN(n16540) );
  NAND3_X1 U15771 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16539) );
  NOR2_X1 U15772 ( .A1(n16402), .A2(n16539), .ZN(n16374) );
  AND2_X1 U15773 ( .A1(n16540), .A2(n16374), .ZN(n16545) );
  NAND2_X1 U15774 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16529) );
  INV_X1 U15775 ( .A(n16529), .ZN(n13946) );
  NAND2_X1 U15776 ( .A1(n16545), .A2(n13946), .ZN(n14040) );
  INV_X1 U15777 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16512) );
  NOR2_X2 U15778 ( .A1(n16347), .A2(n16512), .ZN(n16335) );
  NAND3_X1 U15779 ( .A1(n16303), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16271) );
  AND2_X1 U15780 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15453) );
  AND2_X1 U15781 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U15782 ( .A1(n15453), .A2(n13947), .ZN(n14043) );
  INV_X1 U15783 ( .A(n17142), .ZN(n13948) );
  NOR2_X1 U15784 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13948), .ZN(n17149) );
  NAND2_X1 U15785 ( .A1(n17149), .A2(n18286), .ZN(n13949) );
  NAND2_X1 U15786 ( .A1(n21698), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U15787 ( .A1(n14848), .A2(n13950), .ZN(n17127) );
  AND2_X1 U15788 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16785) );
  NOR2_X1 U15789 ( .A1(n14035), .A2(n17228), .ZN(n15452) );
  AOI21_X1 U15790 ( .B1(n17126), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15452), .ZN(n13951) );
  OAI211_X1 U15791 ( .C1(n18585), .C2(n17125), .A(n13952), .B(n13951), .ZN(
        n13953) );
  AOI21_X1 U15792 ( .B1(n15462), .B2(n17131), .A(n13953), .ZN(n13954) );
  INV_X1 U15793 ( .A(n13955), .ZN(n14823) );
  NAND2_X1 U15794 ( .A1(n18632), .A2(n14823), .ZN(n13957) );
  NAND2_X1 U15795 ( .A1(n13962), .A2(n21735), .ZN(n13956) );
  NAND2_X1 U15796 ( .A1(n13957), .A2(n13956), .ZN(n13958) );
  NAND2_X1 U15797 ( .A1(n13958), .A2(n18291), .ZN(n13981) );
  NAND2_X1 U15798 ( .A1(n15112), .A2(n18291), .ZN(n14773) );
  AOI21_X1 U15799 ( .B1(n13959), .B2(n19628), .A(n12419), .ZN(n13960) );
  NAND2_X1 U15800 ( .A1(n14773), .A2(n13960), .ZN(n13980) );
  INV_X1 U15801 ( .A(n14831), .ZN(n13961) );
  NAND2_X1 U15802 ( .A1(n13962), .A2(n13961), .ZN(n13974) );
  NAND2_X1 U15803 ( .A1(n13963), .A2(n12397), .ZN(n13972) );
  NAND2_X1 U15804 ( .A1(n14372), .A2(n11002), .ZN(n13966) );
  INV_X1 U15805 ( .A(n14820), .ZN(n13965) );
  NAND2_X1 U15806 ( .A1(n13966), .A2(n13965), .ZN(n14012) );
  NAND2_X1 U15807 ( .A1(n12425), .A2(n14009), .ZN(n13967) );
  OAI211_X1 U15808 ( .C1(n12435), .C2(n18291), .A(n12397), .B(n13967), .ZN(
        n13968) );
  NAND4_X1 U15809 ( .A1(n13970), .A2(n13969), .A3(n14012), .A4(n13968), .ZN(
        n13971) );
  AOI21_X1 U15810 ( .B1(n13249), .B2(n13972), .A(n13971), .ZN(n13973) );
  NAND2_X1 U15811 ( .A1(n13974), .A2(n13973), .ZN(n14776) );
  INV_X1 U15812 ( .A(n18292), .ZN(n21744) );
  NAND2_X1 U15813 ( .A1(n18291), .A2(n21744), .ZN(n18296) );
  NAND3_X1 U15814 ( .A1(n18296), .A2(n21735), .A3(n13975), .ZN(n13977) );
  OAI21_X1 U15815 ( .B1(n14833), .B2(n13977), .A(n13976), .ZN(n13978) );
  NOR2_X1 U15816 ( .A1(n14776), .A2(n13978), .ZN(n13979) );
  NAND3_X1 U15817 ( .A1(n13981), .A2(n13980), .A3(n13979), .ZN(n13982) );
  NOR2_X1 U15818 ( .A1(n13988), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13990) );
  MUX2_X1 U15819 ( .A(n13762), .B(n13990), .S(n13989), .Z(n18575) );
  NAND2_X1 U15820 ( .A1(n18575), .A2(n13276), .ZN(n13991) );
  XOR2_X1 U15821 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13991), .Z(
        n13992) );
  XNOR2_X1 U15822 ( .A(n13993), .B(n13992), .ZN(n15472) );
  INV_X1 U15823 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n17229) );
  INV_X1 U15824 ( .A(n13997), .ZN(n13998) );
  NAND2_X1 U15825 ( .A1(n13996), .A2(n13998), .ZN(n14000) );
  AOI22_X1 U15826 ( .A1(n13159), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13999) );
  OAI211_X1 U15827 ( .C1(n13143), .C2(n17229), .A(n14000), .B(n13999), .ZN(
        n14001) );
  NAND2_X1 U15828 ( .A1(n14036), .A2(n13996), .ZN(n16705) );
  AOI22_X1 U15829 ( .A1(n13252), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n13090), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U15830 ( .B1(n13089), .B2(n17229), .A(n14003), .ZN(n14004) );
  XNOR2_X1 U15831 ( .A(n14005), .B(n14004), .ZN(n19115) );
  AND2_X1 U15832 ( .A1(n12905), .A2(n18291), .ZN(n14007) );
  INV_X1 U15833 ( .A(n12894), .ZN(n14767) );
  NOR2_X1 U15834 ( .A1(n14006), .A2(n14767), .ZN(n14825) );
  OR2_X1 U15835 ( .A1(n14007), .A2(n14825), .ZN(n14008) );
  INV_X1 U15836 ( .A(n16540), .ZN(n16588) );
  MUX2_X1 U15837 ( .A(n14010), .B(n12397), .S(n14009), .Z(n14016) );
  NAND2_X1 U15838 ( .A1(n14011), .A2(n18291), .ZN(n14766) );
  NAND2_X1 U15839 ( .A1(n14766), .A2(n14012), .ZN(n14014) );
  NOR2_X1 U15840 ( .A1(n14096), .A2(n12419), .ZN(n14013) );
  AOI21_X1 U15841 ( .B1(n14014), .B2(n12440), .A(n14013), .ZN(n14015) );
  AND2_X1 U15842 ( .A1(n14016), .A2(n14015), .ZN(n14021) );
  OAI211_X1 U15843 ( .C1(n12877), .C2(n14018), .A(n14017), .B(n14096), .ZN(
        n14019) );
  NAND2_X1 U15844 ( .A1(n14019), .A2(n12441), .ZN(n14020) );
  NAND2_X1 U15845 ( .A1(n14785), .A2(n14408), .ZN(n14022) );
  NAND2_X1 U15846 ( .A1(n14036), .A2(n14022), .ZN(n16590) );
  NAND2_X1 U15847 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16739) );
  NOR2_X1 U15848 ( .A1(n14159), .A2(n16739), .ZN(n14343) );
  INV_X1 U15849 ( .A(n14343), .ZN(n14023) );
  NAND2_X1 U15850 ( .A1(n16586), .A2(n14023), .ZN(n14024) );
  NAND2_X1 U15851 ( .A1(n16740), .A2(n14024), .ZN(n16723) );
  INV_X1 U15852 ( .A(n16739), .ZN(n14338) );
  NOR2_X1 U15853 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14338), .ZN(
        n14927) );
  NOR4_X1 U15854 ( .A1(n14927), .A2(n15178), .A3(n15062), .A4(n15174), .ZN(
        n16720) );
  NAND2_X1 U15855 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16720), .ZN(
        n16702) );
  NOR2_X1 U15856 ( .A1(n14025), .A2(n16707), .ZN(n14034) );
  NAND2_X1 U15857 ( .A1(n18615), .A2(n14034), .ZN(n18590) );
  NOR2_X1 U15858 ( .A1(n16588), .A2(n18590), .ZN(n16627) );
  NAND2_X1 U15859 ( .A1(n16374), .A2(n16627), .ZN(n16549) );
  NOR3_X1 U15860 ( .A1(n16345), .A2(n16529), .A3(n16549), .ZN(n16517) );
  NAND3_X1 U15861 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n16517), .ZN(n16483) );
  INV_X1 U15862 ( .A(n16483), .ZN(n14027) );
  NOR2_X1 U15863 ( .A1(n14026), .A2(n16489), .ZN(n16471) );
  AND2_X1 U15864 ( .A1(n14027), .A2(n16471), .ZN(n14028) );
  NAND2_X1 U15865 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14028), .ZN(
        n16437) );
  NOR3_X1 U15866 ( .A1(n14043), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16437), .ZN(n14029) );
  NOR2_X1 U15867 ( .A1(n14035), .A2(n17229), .ZN(n15467) );
  OAI21_X1 U15868 ( .B1(n18579), .B2(n16705), .A(n14030), .ZN(n14046) );
  INV_X1 U15869 ( .A(n16740), .ZN(n16751) );
  INV_X1 U15870 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16520) );
  NOR2_X1 U15871 ( .A1(n16512), .A2(n16520), .ZN(n16505) );
  INV_X1 U15872 ( .A(n14034), .ZN(n18614) );
  NOR2_X1 U15873 ( .A1(n16702), .A2(n18614), .ZN(n14038) );
  NOR2_X1 U15874 ( .A1(n16586), .A2(n14038), .ZN(n14037) );
  INV_X1 U15875 ( .A(n14035), .ZN(n16396) );
  NOR2_X1 U15876 ( .A1(n14036), .A2(n16396), .ZN(n16738) );
  OR2_X1 U15877 ( .A1(n14037), .A2(n16738), .ZN(n16542) );
  NAND2_X1 U15878 ( .A1(n14343), .A2(n14038), .ZN(n16587) );
  INV_X1 U15879 ( .A(n16587), .ZN(n16544) );
  NOR2_X1 U15880 ( .A1(n16590), .A2(n16544), .ZN(n14039) );
  NOR2_X1 U15881 ( .A1(n16542), .A2(n14039), .ZN(n16699) );
  NAND2_X1 U15882 ( .A1(n16740), .A2(n14040), .ZN(n14041) );
  NAND2_X1 U15883 ( .A1(n16699), .A2(n14041), .ZN(n16528) );
  AND2_X1 U15884 ( .A1(n16740), .A2(n16345), .ZN(n14042) );
  NOR2_X1 U15885 ( .A1(n16528), .A2(n14042), .ZN(n16519) );
  OAI21_X1 U15886 ( .B1(n16751), .B2(n16505), .A(n16519), .ZN(n16502) );
  NOR2_X1 U15887 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16483), .ZN(
        n16496) );
  NOR2_X1 U15888 ( .A1(n16502), .A2(n16496), .ZN(n16490) );
  OAI21_X1 U15889 ( .B1(n16751), .B2(n16471), .A(n16490), .ZN(n16465) );
  AOI21_X1 U15890 ( .B1(n16740), .B2(n14043), .A(n16465), .ZN(n15460) );
  OAI21_X1 U15891 ( .B1(n16730), .B2(n15472), .A(n14047), .ZN(P2_U3015) );
  NOR2_X1 U15892 ( .A1(n15620), .A2(n15725), .ZN(n14058) );
  INV_X1 U15893 ( .A(DATAI_28_), .ZN(n16951) );
  INV_X1 U15894 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20012) );
  OR2_X1 U15895 ( .A1(n15202), .A2(n20012), .ZN(n14053) );
  NAND2_X1 U15896 ( .A1(n15202), .A2(DATAI_12_), .ZN(n14052) );
  NAND2_X1 U15897 ( .A1(n14053), .A2(n14052), .ZN(n15225) );
  AOI22_X1 U15898 ( .A1(n15722), .A2(n15225), .B1(n15720), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14054) );
  OAI21_X1 U15899 ( .B1(n15724), .B2(n16951), .A(n14054), .ZN(n14056) );
  AND2_X1 U15900 ( .A1(n15729), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14055) );
  INV_X1 U15901 ( .A(n15729), .ZN(n14067) );
  INV_X1 U15902 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14066) );
  INV_X1 U15903 ( .A(DATAI_30_), .ZN(n16949) );
  INV_X1 U15904 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20016) );
  OR2_X1 U15905 ( .A1(n15202), .A2(n20016), .ZN(n14060) );
  NAND2_X1 U15906 ( .A1(n15202), .A2(DATAI_14_), .ZN(n14059) );
  NAND2_X1 U15907 ( .A1(n14060), .A2(n14059), .ZN(n21855) );
  AOI22_X1 U15908 ( .A1(n15722), .A2(n21855), .B1(n15720), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14061) );
  OAI21_X1 U15909 ( .B1(n15724), .B2(n16949), .A(n14061), .ZN(n14062) );
  INV_X1 U15910 ( .A(n14062), .ZN(n14065) );
  INV_X1 U15911 ( .A(n15725), .ZN(n14063) );
  NAND2_X1 U15912 ( .A1(n15740), .A2(n14063), .ZN(n14064) );
  INV_X1 U15913 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20052) );
  INV_X1 U15914 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22338) );
  NOR4_X1 U15915 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20052), .A4(n22338), .ZN(n14069) );
  NOR4_X1 U15916 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14068) );
  NAND3_X1 U15917 ( .A1(n14544), .A2(n14069), .A3(n14068), .ZN(U214) );
  NOR2_X1 U15918 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14071) );
  NOR4_X1 U15919 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14070) );
  NAND4_X1 U15920 ( .A1(n14071), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14070), .ZN(n14072) );
  OR2_X1 U15921 ( .A1(n14182), .A2(n14072), .ZN(n19989) );
  INV_X2 U15922 ( .A(U214), .ZN(n20038) );
  INV_X1 U15923 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16607) );
  NOR2_X1 U15924 ( .A1(n16607), .A2(n16623), .ZN(n16414) );
  AOI211_X1 U15925 ( .C1(n16623), .C2(n16607), .A(n16414), .B(n17119), .ZN(
        n14084) );
  NOR2_X1 U15926 ( .A1(n14035), .A2(n13063), .ZN(n16599) );
  OAI22_X1 U15927 ( .A1(n16084), .A2(n17117), .B1(n17125), .B2(n16076), .ZN(
        n14083) );
  AND2_X1 U15928 ( .A1(n16612), .A2(n17106), .ZN(n14076) );
  NAND2_X1 U15929 ( .A1(n14078), .A2(n14077), .ZN(n16359) );
  OAI21_X1 U15930 ( .B1(n14078), .B2(n14077), .A(n16359), .ZN(n16603) );
  OAI21_X1 U15931 ( .B1(n14079), .B2(n14081), .A(n14080), .ZN(n16602) );
  OAI22_X1 U15932 ( .A1(n16603), .A2(n17120), .B1(n17113), .B2(n16602), .ZN(
        n14082) );
  OAI21_X1 U15933 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14086), .A(
        n14085), .ZN(n16731) );
  NOR2_X1 U15934 ( .A1(n16731), .A2(n17120), .ZN(n14092) );
  OAI21_X1 U15935 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14088), .A(
        n14087), .ZN(n16736) );
  OAI22_X1 U15936 ( .A1(n16736), .A2(n17119), .B1(n17117), .B2(n14089), .ZN(
        n14091) );
  OAI22_X1 U15937 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17125), .B1(
        n17113), .B2(n15128), .ZN(n14090) );
  NOR2_X1 U15938 ( .A1(n14035), .A2(n12472), .ZN(n16735) );
  OR4_X1 U15939 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n16735), .ZN(
        P2_U3013) );
  NAND2_X1 U15940 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17614) );
  NOR2_X1 U15941 ( .A1(n21277), .A2(n17614), .ZN(n16775) );
  OAI211_X1 U15942 ( .C1(n20773), .C2(n20759), .A(n15367), .B(n15410), .ZN(
        n17615) );
  NAND2_X1 U15943 ( .A1(n20750), .A2(n21144), .ZN(n21267) );
  INV_X1 U15944 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21284) );
  INV_X1 U15945 ( .A(n16775), .ZN(n21262) );
  NOR2_X1 U15946 ( .A1(n21284), .A2(n21262), .ZN(n15430) );
  AOI211_X2 U15947 ( .C1(n16775), .C2(n17615), .A(n18966), .B(n15430), .ZN(
        n18178) );
  AND2_X1 U15948 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18178), .ZN(
        P3_U2867) );
  INV_X1 U15949 ( .A(n18307), .ZN(n14095) );
  INV_X1 U15950 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14094) );
  NAND2_X1 U15951 ( .A1(n19321), .A2(n14093), .ZN(n17056) );
  OAI211_X1 U15952 ( .C1(n14095), .C2(n14094), .A(n14100), .B(n17056), .ZN(
        P2_U2814) );
  INV_X1 U15953 ( .A(n14096), .ZN(n14099) );
  INV_X1 U15954 ( .A(n17055), .ZN(n18288) );
  INV_X1 U15955 ( .A(n17056), .ZN(n14097) );
  OAI21_X1 U15956 ( .B1(n14097), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18288), 
        .ZN(n14098) );
  OAI21_X1 U15957 ( .B1(n14099), .B2(n18288), .A(n14098), .ZN(P2_U3612) );
  INV_X1 U15958 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U15959 ( .A1(n17039), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14182), .ZN(n19405) );
  NOR2_X1 U15960 ( .A1(n14268), .A2(n19405), .ZN(n14169) );
  AOI21_X1 U15961 ( .B1(n14220), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14169), .ZN(
        n14101) );
  OAI21_X1 U15962 ( .B1(n14131), .B2(n14102), .A(n14101), .ZN(P2_U2957) );
  INV_X1 U15963 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14104) );
  INV_X1 U15964 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20001) );
  INV_X1 U15965 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20595) );
  AOI22_X1 U15966 ( .A1(n17039), .A2(n20001), .B1(n20595), .B2(n14182), .ZN(
        n19344) );
  INV_X1 U15967 ( .A(n19344), .ZN(n19352) );
  NOR2_X1 U15968 ( .A1(n14268), .A2(n19352), .ZN(n14205) );
  AOI21_X1 U15969 ( .B1(n14220), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14205), .ZN(
        n14103) );
  OAI21_X1 U15970 ( .B1(n14131), .B2(n14104), .A(n14103), .ZN(P2_U2958) );
  INV_X1 U15971 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U15972 ( .A1(n17039), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14182), .ZN(n19131) );
  NOR2_X1 U15973 ( .A1(n14268), .A2(n19131), .ZN(n14190) );
  AOI21_X1 U15974 ( .B1(n14220), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14190), .ZN(
        n14105) );
  OAI21_X1 U15975 ( .B1(n14131), .B2(n14106), .A(n14105), .ZN(P2_U2959) );
  INV_X1 U15976 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U15977 ( .A1(n17039), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14182), .ZN(n16222) );
  NOR2_X1 U15978 ( .A1(n14268), .A2(n16222), .ZN(n14199) );
  AOI21_X1 U15979 ( .B1(n14220), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14199), .ZN(
        n14107) );
  OAI21_X1 U15980 ( .B1(n14131), .B2(n14108), .A(n14107), .ZN(P2_U2960) );
  INV_X1 U15981 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14110) );
  INV_X1 U15982 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n19997) );
  INV_X1 U15983 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20604) );
  AOI22_X1 U15984 ( .A1(n17039), .A2(n19997), .B1(n20604), .B2(n14182), .ZN(
        n19445) );
  INV_X1 U15985 ( .A(n19445), .ZN(n19451) );
  NOR2_X1 U15986 ( .A1(n14268), .A2(n19451), .ZN(n14202) );
  AOI21_X1 U15987 ( .B1(n14220), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14202), .ZN(
        n14109) );
  OAI21_X1 U15988 ( .B1(n14131), .B2(n14110), .A(n14109), .ZN(P2_U2956) );
  INV_X1 U15989 ( .A(n14111), .ZN(n14114) );
  INV_X1 U15990 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14113) );
  AND2_X1 U15991 ( .A1(n21935), .A2(n16839), .ZN(n15448) );
  INV_X1 U15992 ( .A(n15448), .ZN(n14112) );
  OAI211_X1 U15993 ( .C1(n14114), .C2(n14113), .A(n14212), .B(n14112), .ZN(
        P1_U2801) );
  INV_X1 U15994 ( .A(n12278), .ZN(n14116) );
  AND2_X1 U15995 ( .A1(n14310), .A2(n15447), .ZN(n14115) );
  AOI21_X1 U15996 ( .B1(n14117), .B2(n14116), .A(n14115), .ZN(n19983) );
  INV_X1 U15997 ( .A(n14255), .ZN(n14717) );
  NOR2_X1 U15998 ( .A1(n14717), .A2(n14214), .ZN(n14239) );
  OR2_X1 U15999 ( .A1(n14239), .A2(n14118), .ZN(n14119) );
  NAND2_X1 U16000 ( .A1(n14119), .A2(n21716), .ZN(n21289) );
  NAND2_X1 U16001 ( .A1(n19983), .A2(n21289), .ZN(n16820) );
  AND2_X1 U16002 ( .A1(n16820), .A2(n14314), .ZN(n21669) );
  INV_X1 U16003 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n14130) );
  INV_X1 U16004 ( .A(n14120), .ZN(n14300) );
  AND2_X1 U16005 ( .A1(n16817), .A2(n14121), .ZN(n14319) );
  NAND3_X1 U16006 ( .A1(n14122), .A2(n12273), .A3(n11553), .ZN(n14123) );
  NAND2_X1 U16007 ( .A1(n14319), .A2(n14123), .ZN(n14124) );
  NAND2_X1 U16008 ( .A1(n14124), .A2(n14310), .ZN(n14126) );
  OR2_X1 U16009 ( .A1(n14329), .A2(n14310), .ZN(n14125) );
  OAI211_X1 U16010 ( .C1(n14300), .C2(n14254), .A(n14126), .B(n14125), .ZN(
        n14127) );
  NAND2_X1 U16011 ( .A1(n14127), .A2(n14578), .ZN(n16818) );
  INV_X1 U16012 ( .A(n16818), .ZN(n14128) );
  NAND2_X1 U16013 ( .A1(n21669), .A2(n14128), .ZN(n14129) );
  OAI21_X1 U16014 ( .B1(n21669), .B2(n14130), .A(n14129), .ZN(P1_U3484) );
  INV_X1 U16015 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17206) );
  NAND2_X1 U16016 ( .A1(n14166), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14132) );
  INV_X1 U16017 ( .A(n14268), .ZN(n14142) );
  MUX2_X1 U16018 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14182), .Z(n19122) );
  NAND2_X1 U16019 ( .A1(n14142), .A2(n19122), .ZN(n14136) );
  OAI211_X1 U16020 ( .C1(n17206), .C2(n14267), .A(n14132), .B(n14136), .ZN(
        P2_U2979) );
  INV_X1 U16021 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U16022 ( .A1(n14166), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14134) );
  NOR2_X1 U16023 ( .A1(n14182), .A2(n20016), .ZN(n14133) );
  AOI21_X1 U16024 ( .B1(n14182), .B2(BUF2_REG_14__SCAN_IN), .A(n14133), .ZN(
        n15500) );
  INV_X1 U16025 ( .A(n15500), .ZN(n19119) );
  NAND2_X1 U16026 ( .A1(n14142), .A2(n19119), .ZN(n14144) );
  OAI211_X1 U16027 ( .C1(n14403), .C2(n14267), .A(n14134), .B(n14144), .ZN(
        P2_U2966) );
  INV_X1 U16028 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17202) );
  NAND2_X1 U16029 ( .A1(n14166), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14135) );
  MUX2_X1 U16030 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14182), .Z(n19125) );
  NAND2_X1 U16031 ( .A1(n14142), .A2(n19125), .ZN(n14140) );
  OAI211_X1 U16032 ( .C1(n17202), .C2(n14267), .A(n14135), .B(n14140), .ZN(
        P2_U2977) );
  INV_X1 U16033 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U16034 ( .A1(n14166), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14137) );
  OAI211_X1 U16035 ( .C1(n14396), .C2(n14267), .A(n14137), .B(n14136), .ZN(
        P2_U2964) );
  NAND2_X1 U16036 ( .A1(n14166), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U16037 ( .A1(n14142), .A2(n14138), .ZN(n14218) );
  OAI211_X1 U16038 ( .C1(n14267), .C2(n14392), .A(n14139), .B(n14218), .ZN(
        P2_U2965) );
  INV_X1 U16039 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U16040 ( .A1(n14166), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14141) );
  OAI211_X1 U16041 ( .C1(n14390), .C2(n14267), .A(n14141), .B(n14140), .ZN(
        P2_U2962) );
  INV_X1 U16042 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16191) );
  NAND2_X1 U16043 ( .A1(n14166), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U16044 ( .A1(n17039), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n14182), .ZN(n14598) );
  INV_X1 U16045 ( .A(n14598), .ZN(n16188) );
  NAND2_X1 U16046 ( .A1(n14142), .A2(n16188), .ZN(n14222) );
  OAI211_X1 U16047 ( .C1(n14267), .C2(n16191), .A(n14143), .B(n14222), .ZN(
        P2_U2963) );
  INV_X1 U16048 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17210) );
  NAND2_X1 U16049 ( .A1(n14166), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14145) );
  OAI211_X1 U16050 ( .C1(n17210), .C2(n14267), .A(n14145), .B(n14144), .ZN(
        P2_U2981) );
  INV_X1 U16051 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16221) );
  OAI21_X1 U16052 ( .B1(n14773), .B2(n14146), .A(n14267), .ZN(n14147) );
  NOR2_X1 U16053 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17142), .ZN(n17200) );
  NOR2_X4 U16054 ( .A1(n17180), .A2(n17211), .ZN(n17192) );
  AOI22_X1 U16055 ( .A1(n17211), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14148) );
  OAI21_X1 U16056 ( .B1(n16221), .B2(n14402), .A(n14148), .ZN(P2_U2927) );
  INV_X1 U16057 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16211) );
  AOI22_X1 U16058 ( .A1(n17211), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U16059 ( .B1(n16211), .B2(n14402), .A(n14149), .ZN(P2_U2926) );
  INV_X1 U16060 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16231) );
  AOI22_X1 U16061 ( .A1(n17211), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14150) );
  OAI21_X1 U16062 ( .B1(n16231), .B2(n14402), .A(n14150), .ZN(P2_U2928) );
  INV_X1 U16063 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16241) );
  AOI22_X1 U16064 ( .A1(n17211), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U16065 ( .B1(n16241), .B2(n14402), .A(n14151), .ZN(P2_U2930) );
  INV_X1 U16066 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U16067 ( .A1(n17211), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14152) );
  OAI21_X1 U16068 ( .B1(n14153), .B2(n14402), .A(n14152), .ZN(P2_U2929) );
  AOI21_X1 U16069 ( .B1(n15097), .B2(n14155), .A(n14154), .ZN(n14156) );
  XNOR2_X1 U16070 ( .A(n14156), .B(n14159), .ZN(n14350) );
  INV_X1 U16071 ( .A(n14350), .ZN(n14165) );
  NOR2_X1 U16072 ( .A1(n14158), .A2(n14157), .ZN(n14160) );
  XNOR2_X1 U16073 ( .A(n14160), .B(n14159), .ZN(n14349) );
  NOR2_X1 U16074 ( .A1(n14035), .A2(n17217), .ZN(n14341) );
  NOR2_X1 U16075 ( .A1(n17117), .A2(n14161), .ZN(n14162) );
  AOI211_X1 U16076 ( .C1(n14349), .C2(n17131), .A(n14341), .B(n14162), .ZN(
        n14164) );
  AOI22_X1 U16077 ( .A1(n15095), .A2(n17105), .B1(n17133), .B2(n15096), .ZN(
        n14163) );
  OAI211_X1 U16078 ( .C1(n14165), .C2(n17120), .A(n14164), .B(n14163), .ZN(
        P2_U3012) );
  INV_X1 U16079 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U16080 ( .A1(n17039), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14182), .ZN(n19532) );
  NOR2_X1 U16081 ( .A1(n14268), .A2(n19532), .ZN(n14172) );
  AOI21_X1 U16082 ( .B1(n14220), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14172), .ZN(
        n14167) );
  OAI21_X1 U16083 ( .B1(n14270), .B2(n14168), .A(n14167), .ZN(P2_U2954) );
  INV_X1 U16084 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14171) );
  AOI21_X1 U16085 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n14220), .A(n14169), .ZN(
        n14170) );
  OAI21_X1 U16086 ( .B1(n14270), .B2(n14171), .A(n14170), .ZN(P2_U2972) );
  INV_X1 U16087 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14174) );
  AOI21_X1 U16088 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n14220), .A(n14172), .ZN(
        n14173) );
  OAI21_X1 U16089 ( .B1(n14270), .B2(n14174), .A(n14173), .ZN(P2_U2969) );
  INV_X1 U16090 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14176) );
  INV_X1 U16091 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n19991) );
  INV_X1 U16092 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19012) );
  AOI22_X1 U16093 ( .A1(n17039), .A2(n19991), .B1(n19012), .B2(n14182), .ZN(
        n19614) );
  INV_X1 U16094 ( .A(n19614), .ZN(n19626) );
  NOR2_X1 U16095 ( .A1(n14268), .A2(n19626), .ZN(n14179) );
  AOI21_X1 U16096 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n14220), .A(n14179), .ZN(
        n14175) );
  OAI21_X1 U16097 ( .B1(n14270), .B2(n14176), .A(n14175), .ZN(P2_U2967) );
  INV_X1 U16098 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U16099 ( .A1(n17039), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14182), .ZN(n17042) );
  NOR2_X1 U16100 ( .A1(n14268), .A2(n17042), .ZN(n14193) );
  AOI21_X1 U16101 ( .B1(n14220), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14193), .ZN(
        n14177) );
  OAI21_X1 U16102 ( .B1(n14270), .B2(n14178), .A(n14177), .ZN(P2_U2955) );
  INV_X1 U16103 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14181) );
  AOI21_X1 U16104 ( .B1(n14220), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14179), .ZN(
        n14180) );
  OAI21_X1 U16105 ( .B1(n14270), .B2(n14181), .A(n14180), .ZN(P2_U2952) );
  INV_X1 U16106 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U16107 ( .A1(n17039), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14182), .ZN(n19573) );
  NOR2_X1 U16108 ( .A1(n14268), .A2(n19573), .ZN(n14185) );
  AOI21_X1 U16109 ( .B1(n14220), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14185), .ZN(
        n14183) );
  OAI21_X1 U16110 ( .B1(n14270), .B2(n14184), .A(n14183), .ZN(P2_U2953) );
  INV_X1 U16111 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14187) );
  AOI21_X1 U16112 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14220), .A(n14185), .ZN(
        n14186) );
  OAI21_X1 U16113 ( .B1(n14270), .B2(n14187), .A(n14186), .ZN(P2_U2968) );
  INV_X1 U16114 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U16115 ( .A1(n17039), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n14182), .ZN(n16212) );
  NOR2_X1 U16116 ( .A1(n14268), .A2(n16212), .ZN(n14196) );
  AOI21_X1 U16117 ( .B1(n14220), .B2(P2_EAX_REG_25__SCAN_IN), .A(n14196), .ZN(
        n14188) );
  OAI21_X1 U16118 ( .B1(n14270), .B2(n14189), .A(n14188), .ZN(P2_U2961) );
  INV_X1 U16119 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14192) );
  AOI21_X1 U16120 ( .B1(n14220), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14190), .ZN(
        n14191) );
  OAI21_X1 U16121 ( .B1(n14270), .B2(n14192), .A(n14191), .ZN(P2_U2974) );
  INV_X1 U16122 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14195) );
  AOI21_X1 U16123 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n14220), .A(n14193), .ZN(
        n14194) );
  OAI21_X1 U16124 ( .B1(n14270), .B2(n14195), .A(n14194), .ZN(P2_U2970) );
  INV_X1 U16125 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14198) );
  AOI21_X1 U16126 ( .B1(n14220), .B2(P2_EAX_REG_9__SCAN_IN), .A(n14196), .ZN(
        n14197) );
  OAI21_X1 U16127 ( .B1(n14270), .B2(n14198), .A(n14197), .ZN(P2_U2976) );
  INV_X1 U16128 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14201) );
  AOI21_X1 U16129 ( .B1(P2_EAX_REG_8__SCAN_IN), .B2(n14220), .A(n14199), .ZN(
        n14200) );
  OAI21_X1 U16130 ( .B1(n14270), .B2(n14201), .A(n14200), .ZN(P2_U2975) );
  INV_X1 U16131 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14204) );
  AOI21_X1 U16132 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n14220), .A(n14202), .ZN(
        n14203) );
  OAI21_X1 U16133 ( .B1(n14270), .B2(n14204), .A(n14203), .ZN(P2_U2971) );
  INV_X1 U16134 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14207) );
  AOI21_X1 U16135 ( .B1(n14220), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14205), .ZN(
        n14206) );
  OAI21_X1 U16136 ( .B1(n14270), .B2(n14207), .A(n14206), .ZN(P2_U2973) );
  NAND2_X1 U16137 ( .A1(n12278), .A2(n11549), .ZN(n16832) );
  INV_X1 U16138 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14216) );
  INV_X1 U16139 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14209) );
  OR2_X1 U16140 ( .A1(n15202), .A2(n14209), .ZN(n14211) );
  NAND2_X1 U16141 ( .A1(n15202), .A2(DATAI_15_), .ZN(n14210) );
  AND2_X1 U16142 ( .A1(n14211), .A2(n14210), .ZN(n15258) );
  INV_X1 U16143 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14215) );
  INV_X1 U16144 ( .A(n14212), .ZN(n14213) );
  OAI21_X2 U16145 ( .B1(n14214), .B2(n21716), .A(n14213), .ZN(n21843) );
  OAI222_X1 U16146 ( .A1(n21863), .A2(n14216), .B1(n21857), .B2(n15258), .C1(
        n14215), .C2(n21801), .ZN(P1_U2967) );
  INV_X1 U16147 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14219) );
  NAND2_X1 U16148 ( .A1(n14220), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14217) );
  OAI211_X1 U16149 ( .C1(n14270), .C2(n14219), .A(n14218), .B(n14217), .ZN(
        P2_U2980) );
  INV_X1 U16150 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14223) );
  NAND2_X1 U16151 ( .A1(n14220), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14221) );
  OAI211_X1 U16152 ( .C1(n14270), .C2(n14223), .A(n14222), .B(n14221), .ZN(
        P2_U2978) );
  AOI22_X1 U16153 ( .A1(n14321), .A2(n14225), .B1(n14224), .B2(n14717), .ZN(
        n14226) );
  OAI21_X1 U16154 ( .B1(n14227), .B2(n15446), .A(n14226), .ZN(n14228) );
  INV_X1 U16155 ( .A(n14228), .ZN(n14232) );
  MUX2_X1 U16156 ( .A(n14230), .B(n11549), .S(n14229), .Z(n14231) );
  NAND2_X1 U16157 ( .A1(n14231), .A2(n11553), .ZN(n14252) );
  AND3_X1 U16158 ( .A1(n14233), .A2(n14232), .A3(n14252), .ZN(n14332) );
  NOR2_X1 U16159 ( .A1(n14235), .A2(n10970), .ZN(n14236) );
  AND2_X1 U16160 ( .A1(n14234), .A2(n14236), .ZN(n14237) );
  NAND2_X1 U16161 ( .A1(n14332), .A2(n14237), .ZN(n16037) );
  NAND2_X1 U16162 ( .A1(n21961), .A2(n16037), .ZN(n14247) );
  INV_X1 U16163 ( .A(n14238), .ZN(n16032) );
  NAND2_X1 U16164 ( .A1(n16032), .A2(n11015), .ZN(n14451) );
  NAND2_X1 U16165 ( .A1(n14238), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14446) );
  NAND2_X1 U16166 ( .A1(n14451), .A2(n14446), .ZN(n14241) );
  INV_X1 U16167 ( .A(n14241), .ZN(n14248) );
  NAND2_X1 U16168 ( .A1(n11031), .A2(n14248), .ZN(n14244) );
  XNOR2_X1 U16169 ( .A(n11015), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14242) );
  AND2_X1 U16170 ( .A1(n14240), .A2(n14239), .ZN(n14453) );
  AOI22_X1 U16171 ( .A1(n14455), .A2(n14242), .B1(n14453), .B2(n14241), .ZN(
        n14243) );
  OAI21_X1 U16172 ( .B1(n16037), .B2(n14244), .A(n14243), .ZN(n14245) );
  INV_X1 U16173 ( .A(n14245), .ZN(n14246) );
  NAND2_X1 U16174 ( .A1(n14247), .A2(n14246), .ZN(n14444) );
  INV_X1 U16175 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14359) );
  NOR2_X1 U16176 ( .A1(n16839), .A2(n14359), .ZN(n16041) );
  INV_X1 U16177 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15888) );
  INV_X1 U16178 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U16179 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n15888), .B2(n15882), .ZN(
        n16039) );
  AOI222_X1 U16180 ( .A1(n14444), .A2(n16038), .B1(n16041), .B2(n16039), .C1(
        n14248), .C2(n21686), .ZN(n14266) );
  INV_X1 U16181 ( .A(n21716), .ZN(n16835) );
  OR3_X1 U16182 ( .A1(n14310), .A2(n16835), .A3(n21726), .ZN(n16827) );
  NAND2_X1 U16183 ( .A1(n14249), .A2(n16827), .ZN(n14250) );
  OAI21_X1 U16184 ( .B1(n14455), .B2(n14235), .A(n14250), .ZN(n14258) );
  NAND2_X1 U16185 ( .A1(n14252), .A2(n14251), .ZN(n14253) );
  NAND2_X1 U16186 ( .A1(n14254), .A2(n14253), .ZN(n14312) );
  OR2_X1 U16187 ( .A1(n14255), .A2(n11551), .ZN(n14256) );
  NAND4_X1 U16188 ( .A1(n14258), .A2(n14312), .A3(n14257), .A4(n14256), .ZN(
        n14259) );
  OR2_X1 U16189 ( .A1(n14260), .A2(n14259), .ZN(n14464) );
  NAND2_X1 U16190 ( .A1(n14464), .A2(n14314), .ZN(n14264) );
  INV_X1 U16191 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21668) );
  NAND2_X1 U16192 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21682) );
  NOR3_X1 U16193 ( .A1(n21683), .A2(n21668), .A3(n21682), .ZN(n14262) );
  NOR2_X1 U16194 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21930), .ZN(n14261) );
  NOR2_X1 U16195 ( .A1(n14262), .A2(n14261), .ZN(n14263) );
  NAND2_X1 U16196 ( .A1(n21675), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14265) );
  OAI21_X1 U16197 ( .B1(n14266), .B2(n21675), .A(n14265), .ZN(P1_U3472) );
  INV_X1 U16198 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14269) );
  AOI22_X1 U16199 ( .A1(n17039), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14182), .ZN(n14939) );
  INV_X1 U16200 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17214) );
  OAI222_X1 U16201 ( .A1(n14270), .A2(n14269), .B1(n14268), .B2(n14939), .C1(
        n14267), .C2(n17214), .ZN(P2_U2982) );
  INV_X1 U16202 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21818) );
  INV_X1 U16203 ( .A(n14455), .ZN(n16035) );
  NAND2_X1 U16204 ( .A1(n16035), .A2(n16832), .ZN(n14273) );
  NOR2_X1 U16205 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21682), .ZN(n19811) );
  NOR2_X4 U16206 ( .A1(n19801), .A2(n21288), .ZN(n19808) );
  AOI22_X1 U16207 ( .A1(n19811), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U16208 ( .B1(n21818), .B2(n14434), .A(n14274), .ZN(P1_U2913) );
  INV_X1 U16209 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21808) );
  AOI22_X1 U16210 ( .A1(n21288), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14275) );
  OAI21_X1 U16211 ( .B1(n21808), .B2(n14434), .A(n14275), .ZN(P1_U2915) );
  INV_X1 U16212 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21828) );
  AOI22_X1 U16213 ( .A1(n21288), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14276) );
  OAI21_X1 U16214 ( .B1(n21828), .B2(n14434), .A(n14276), .ZN(P1_U2911) );
  INV_X1 U16215 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21823) );
  AOI22_X1 U16216 ( .A1(n21288), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14277) );
  OAI21_X1 U16217 ( .B1(n21823), .B2(n14434), .A(n14277), .ZN(P1_U2912) );
  AOI22_X1 U16218 ( .A1(n21288), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14278) );
  OAI21_X1 U16219 ( .B1(n12064), .B2(n14434), .A(n14278), .ZN(P1_U2914) );
  INV_X1 U16220 ( .A(n11698), .ZN(n14477) );
  INV_X1 U16221 ( .A(n16037), .ZN(n14279) );
  OAI22_X1 U16222 ( .A1(n14477), .A2(n14279), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11558), .ZN(n16804) );
  OAI22_X1 U16223 ( .A1(n16839), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21671), .ZN(n14280) );
  AOI21_X1 U16224 ( .B1(n16804), .B2(n16038), .A(n14280), .ZN(n14283) );
  NOR2_X1 U16225 ( .A1(n16035), .A2(n14281), .ZN(n16803) );
  AOI22_X1 U16226 ( .A1(n21675), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n16038), .B2(n16803), .ZN(n14282) );
  OAI21_X1 U16227 ( .B1(n14283), .B2(n21675), .A(n14282), .ZN(P1_U3474) );
  OAI21_X1 U16228 ( .B1(n14285), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14284), .ZN(n14337) );
  INV_X1 U16229 ( .A(n14286), .ZN(n14287) );
  AOI21_X1 U16230 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n14879) );
  NAND2_X1 U16231 ( .A1(n14879), .A2(n19979), .ZN(n14294) );
  NAND2_X1 U16232 ( .A1(n14290), .A2(n15874), .ZN(n14292) );
  INV_X1 U16233 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14291) );
  NOR2_X1 U16234 ( .A1(n21616), .A2(n14291), .ZN(n14327) );
  AOI21_X1 U16235 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14292), .A(
        n14327), .ZN(n14293) );
  OAI211_X1 U16236 ( .C1(n21667), .C2(n14337), .A(n14294), .B(n14293), .ZN(
        P1_U2999) );
  INV_X1 U16237 ( .A(n21960), .ZN(n14547) );
  OR2_X1 U16238 ( .A1(n14295), .A2(n14547), .ZN(n14296) );
  XNOR2_X1 U16239 ( .A(n14296), .B(n14465), .ZN(n21484) );
  INV_X1 U16240 ( .A(n21675), .ZN(n16044) );
  INV_X1 U16241 ( .A(n14234), .ZN(n14297) );
  NAND3_X1 U16242 ( .A1(n16044), .A2(n16038), .A3(n14297), .ZN(n14298) );
  OAI22_X1 U16243 ( .A1(n21484), .A2(n14298), .B1(n14465), .B2(n16044), .ZN(
        P1_U3468) );
  AOI21_X1 U16244 ( .B1(n13348), .B2(n21726), .A(n16835), .ZN(n14299) );
  NAND2_X1 U16245 ( .A1(n14300), .A2(n14299), .ZN(n14309) );
  INV_X1 U16246 ( .A(n14301), .ZN(n14302) );
  NAND2_X1 U16247 ( .A1(n14235), .A2(n14302), .ZN(n14304) );
  NAND3_X1 U16248 ( .A1(n14304), .A2(n11553), .A3(n14303), .ZN(n14306) );
  NAND2_X1 U16249 ( .A1(n14306), .A2(n14305), .ZN(n14308) );
  MUX2_X1 U16250 ( .A(n14309), .B(n14308), .S(n14307), .Z(n14313) );
  NAND3_X1 U16251 ( .A1(n14310), .A2(n16033), .A3(n13348), .ZN(n14311) );
  NAND3_X1 U16252 ( .A1(n14313), .A2(n14312), .A3(n14311), .ZN(n14315) );
  INV_X1 U16253 ( .A(n14316), .ZN(n14317) );
  AOI22_X1 U16254 ( .A1(n14317), .A2(n14564), .B1(n14235), .B2(n14356), .ZN(
        n14318) );
  NAND3_X1 U16255 ( .A1(n14319), .A2(n14318), .A3(n14234), .ZN(n14320) );
  NOR2_X1 U16256 ( .A1(n14321), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14322) );
  OR2_X1 U16257 ( .A1(n14323), .A2(n14322), .ZN(n14875) );
  INV_X1 U16258 ( .A(n14875), .ZN(n14328) );
  OAI21_X1 U16259 ( .B1(n14316), .B2(n14564), .A(n16832), .ZN(n14324) );
  INV_X2 U16260 ( .A(n21616), .ZN(n21457) );
  NOR2_X1 U16261 ( .A1(n21457), .A2(n14334), .ZN(n15881) );
  INV_X1 U16262 ( .A(n15881), .ZN(n14325) );
  AOI21_X1 U16263 ( .B1(n21296), .B2(n14325), .A(n14359), .ZN(n14326) );
  AOI211_X1 U16264 ( .C1(n14328), .C2(n21461), .A(n14327), .B(n14326), .ZN(
        n14336) );
  INV_X1 U16265 ( .A(n14329), .ZN(n14330) );
  NAND2_X1 U16266 ( .A1(n14332), .A2(n14331), .ZN(n14333) );
  NAND2_X1 U16267 ( .A1(n14334), .A2(n14333), .ZN(n21297) );
  AOI21_X1 U16268 ( .B1(n21334), .B2(n21297), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14357) );
  INV_X1 U16269 ( .A(n14357), .ZN(n14335) );
  OAI211_X1 U16270 ( .C1(n14337), .C2(n21430), .A(n14336), .B(n14335), .ZN(
        P1_U3031) );
  NOR2_X1 U16271 ( .A1(n16590), .A2(n14343), .ZN(n14925) );
  INV_X1 U16272 ( .A(n14925), .ZN(n14353) );
  INV_X1 U16273 ( .A(n16738), .ZN(n16750) );
  OAI21_X1 U16274 ( .B1(n14338), .B2(n16590), .A(n16750), .ZN(n14348) );
  XNOR2_X1 U16275 ( .A(n14339), .B(n14340), .ZN(n17151) );
  AOI21_X1 U16276 ( .B1(n18606), .B2(n17151), .A(n14341), .ZN(n14346) );
  INV_X1 U16277 ( .A(n16586), .ZN(n14342) );
  OAI21_X1 U16278 ( .B1(n14343), .B2(n14927), .A(n14342), .ZN(n14345) );
  NAND2_X1 U16279 ( .A1(n18611), .A2(n15096), .ZN(n14344) );
  NAND3_X1 U16280 ( .A1(n14346), .A2(n14345), .A3(n14344), .ZN(n14347) );
  AOI21_X1 U16281 ( .B1(n14348), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14347), .ZN(n14352) );
  AOI22_X1 U16282 ( .A1(n14350), .A2(n18609), .B1(n18612), .B2(n14349), .ZN(
        n14351) );
  OAI211_X1 U16283 ( .C1(n14353), .C2(n16739), .A(n14352), .B(n14351), .ZN(
        P2_U3044) );
  OR2_X1 U16284 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14369) );
  NAND3_X1 U16285 ( .A1(n14369), .A2(n14355), .A3(n21462), .ZN(n14364) );
  XNOR2_X1 U16286 ( .A(n21477), .B(n14356), .ZN(n14424) );
  OAI21_X1 U16287 ( .B1(n14357), .B2(n15881), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14358) );
  OAI21_X1 U16288 ( .B1(n14424), .B2(n21429), .A(n14358), .ZN(n14362) );
  NAND2_X1 U16289 ( .A1(n14359), .A2(n21296), .ZN(n15890) );
  INV_X1 U16290 ( .A(n15890), .ZN(n14360) );
  NOR3_X1 U16291 ( .A1(n21426), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14360), .ZN(n14361) );
  AOI211_X1 U16292 ( .C1(n21457), .C2(P1_REIP_REG_1__SCAN_IN), .A(n14362), .B(
        n14361), .ZN(n14363) );
  NAND2_X1 U16293 ( .A1(n14364), .A2(n14363), .ZN(P1_U3030) );
  OAI21_X1 U16294 ( .B1(n14366), .B2(n14365), .A(n14505), .ZN(n21472) );
  INV_X1 U16295 ( .A(n19979), .ZN(n19947) );
  INV_X1 U16296 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14367) );
  OAI22_X1 U16297 ( .A1(n15874), .A2(n21474), .B1(n21616), .B2(n14367), .ZN(
        n14368) );
  AOI21_X1 U16298 ( .B1(n19965), .B2(n21474), .A(n14368), .ZN(n14371) );
  NAND3_X1 U16299 ( .A1(n14369), .A2(n14355), .A3(n19978), .ZN(n14370) );
  OAI211_X1 U16300 ( .C1(n21472), .C2(n19947), .A(n14371), .B(n14370), .ZN(
        P1_U2998) );
  INV_X1 U16301 ( .A(n14373), .ZN(n15114) );
  NAND2_X1 U16302 ( .A1(n18291), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14374) );
  NAND4_X1 U16303 ( .A1(n14374), .A2(n19353), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19293), .ZN(n14375) );
  INV_X1 U16304 ( .A(n14376), .ZN(n14382) );
  INV_X1 U16305 ( .A(n14377), .ZN(n14380) );
  INV_X1 U16306 ( .A(n14378), .ZN(n14379) );
  NAND2_X1 U16307 ( .A1(n14380), .A2(n14379), .ZN(n14381) );
  NAND2_X1 U16308 ( .A1(n14382), .A2(n14381), .ZN(n15157) );
  INV_X1 U16309 ( .A(n15157), .ZN(n16748) );
  NOR2_X1 U16310 ( .A1(n17144), .A2(n15157), .ZN(n14439) );
  INV_X1 U16311 ( .A(n14439), .ZN(n14383) );
  OAI211_X1 U16312 ( .C1(n17043), .C2(n16748), .A(n14383), .B(n19620), .ZN(
        n14385) );
  AOI22_X1 U16313 ( .A1(n19619), .A2(n16748), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19613), .ZN(n14384) );
  OAI211_X1 U16314 ( .C1(n14958), .C2(n19626), .A(n14385), .B(n14384), .ZN(
        P2_U2919) );
  INV_X1 U16315 ( .A(n14879), .ZN(n14516) );
  OAI222_X1 U16316 ( .A1(n14875), .A2(n15657), .B1(n14876), .B2(n19911), .C1(
        n14516), .C2(n15659), .ZN(P1_U2872) );
  INV_X1 U16317 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U16318 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17192), .B1(n17211), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14386) );
  OAI21_X1 U16319 ( .B1(n14387), .B2(n14402), .A(n14386), .ZN(P2_U2935) );
  AOI22_X1 U16320 ( .A1(n17211), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14388) );
  OAI21_X1 U16321 ( .B1(n16191), .B2(n14402), .A(n14388), .ZN(P2_U2924) );
  AOI22_X1 U16322 ( .A1(n17211), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14389) );
  OAI21_X1 U16323 ( .B1(n14390), .B2(n14402), .A(n14389), .ZN(P2_U2925) );
  AOI22_X1 U16324 ( .A1(n17211), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14391) );
  OAI21_X1 U16325 ( .B1(n14392), .B2(n14402), .A(n14391), .ZN(P2_U2922) );
  INV_X1 U16326 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14394) );
  AOI22_X1 U16327 ( .A1(n17211), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14393) );
  OAI21_X1 U16328 ( .B1(n14394), .B2(n14402), .A(n14393), .ZN(P2_U2931) );
  AOI22_X1 U16329 ( .A1(n17211), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14395) );
  OAI21_X1 U16330 ( .B1(n14396), .B2(n14402), .A(n14395), .ZN(P2_U2923) );
  INV_X1 U16331 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U16332 ( .A1(n17200), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14397) );
  OAI21_X1 U16333 ( .B1(n14398), .B2(n14402), .A(n14397), .ZN(P2_U2933) );
  INV_X1 U16334 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U16335 ( .A1(n17200), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14399) );
  OAI21_X1 U16336 ( .B1(n16249), .B2(n14402), .A(n14399), .ZN(P2_U2932) );
  INV_X1 U16337 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U16338 ( .A1(n17200), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14400) );
  OAI21_X1 U16339 ( .B1(n15216), .B2(n14402), .A(n14400), .ZN(P2_U2934) );
  AOI22_X1 U16340 ( .A1(n17200), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14401) );
  OAI21_X1 U16341 ( .B1(n14403), .B2(n14402), .A(n14401), .ZN(P2_U2921) );
  INV_X1 U16342 ( .A(n15112), .ZN(n14407) );
  AOI21_X4 U16343 ( .B1(n14777), .B2(n14408), .A(n18644), .ZN(n16127) );
  MUX2_X1 U16344 ( .A(n14409), .B(n15128), .S(n16127), .Z(n14410) );
  OAI21_X1 U16345 ( .B1(n19152), .B2(n16178), .A(n14410), .ZN(P2_U2886) );
  MUX2_X1 U16346 ( .A(n14411), .B(n15161), .S(n16127), .Z(n14412) );
  OAI21_X1 U16347 ( .B1(n17144), .B2(n16178), .A(n14412), .ZN(P2_U2887) );
  NOR2_X1 U16348 ( .A1(n16127), .A2(n12475), .ZN(n14415) );
  AOI21_X1 U16349 ( .B1(n16127), .B2(n15096), .A(n14415), .ZN(n14416) );
  OAI21_X1 U16350 ( .B1(n19254), .B2(n16178), .A(n14416), .ZN(P2_U2885) );
  MUX2_X1 U16351 ( .A(n14921), .B(n13271), .S(n16176), .Z(n14421) );
  OAI21_X1 U16352 ( .B1(n19255), .B2(n16178), .A(n14421), .ZN(P2_U2884) );
  INV_X1 U16353 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n21777) );
  AOI22_X1 U16354 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19808), .B1(n19811), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14422) );
  OAI21_X1 U16355 ( .B1(n21777), .B2(n14434), .A(n14422), .ZN(P1_U2920) );
  INV_X1 U16356 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14423) );
  OAI222_X1 U16357 ( .A1(n14424), .A2(n15657), .B1(n19911), .B2(n14423), .C1(
        n21472), .C2(n15659), .ZN(P1_U2871) );
  INV_X1 U16358 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n21783) );
  AOI22_X1 U16359 ( .A1(n19811), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14425) );
  OAI21_X1 U16360 ( .B1(n21783), .B2(n14434), .A(n14425), .ZN(P1_U2919) );
  INV_X1 U16361 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n21789) );
  AOI22_X1 U16362 ( .A1(n21288), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14426) );
  OAI21_X1 U16363 ( .B1(n21789), .B2(n14434), .A(n14426), .ZN(P1_U2918) );
  INV_X1 U16364 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21845) );
  AOI22_X1 U16365 ( .A1(n21288), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14427) );
  OAI21_X1 U16366 ( .B1(n21845), .B2(n14434), .A(n14427), .ZN(P1_U2908) );
  AOI22_X1 U16367 ( .A1(n21288), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14428) );
  OAI21_X1 U16368 ( .B1(n12162), .B2(n14434), .A(n14428), .ZN(P1_U2909) );
  AOI22_X1 U16369 ( .A1(n21288), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14429) );
  OAI21_X1 U16370 ( .B1(n21834), .B2(n14434), .A(n14429), .ZN(P1_U2910) );
  AOI22_X1 U16371 ( .A1(n21288), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14430) );
  OAI21_X1 U16372 ( .B1(n12026), .B2(n14434), .A(n14430), .ZN(P1_U2916) );
  INV_X1 U16373 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n21795) );
  AOI22_X1 U16374 ( .A1(n21288), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14431) );
  OAI21_X1 U16375 ( .B1(n21795), .B2(n14434), .A(n14431), .ZN(P1_U2917) );
  INV_X1 U16376 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21851) );
  AOI22_X1 U16377 ( .A1(n21288), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14432) );
  OAI21_X1 U16378 ( .B1(n21851), .B2(n14434), .A(n14432), .ZN(P1_U2907) );
  INV_X1 U16379 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21860) );
  AOI22_X1 U16380 ( .A1(n21288), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U16381 ( .B1(n21860), .B2(n14434), .A(n14433), .ZN(P1_U2906) );
  OAI21_X1 U16382 ( .B1(n14437), .B2(n14436), .A(n14435), .ZN(n17158) );
  INV_X1 U16383 ( .A(n17158), .ZN(n16732) );
  NAND2_X1 U16384 ( .A1(n19152), .A2(n16732), .ZN(n14668) );
  OAI21_X1 U16385 ( .B1(n19152), .B2(n16732), .A(n14668), .ZN(n14438) );
  NOR2_X1 U16386 ( .A1(n14438), .A2(n14439), .ZN(n14670) );
  AOI21_X1 U16387 ( .B1(n14439), .B2(n14438), .A(n14670), .ZN(n14443) );
  AOI22_X1 U16388 ( .A1(n19619), .A2(n17158), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19613), .ZN(n14442) );
  INV_X1 U16389 ( .A(n14958), .ZN(n19397) );
  INV_X1 U16390 ( .A(n19573), .ZN(n14440) );
  NAND2_X1 U16391 ( .A1(n19397), .A2(n14440), .ZN(n14441) );
  OAI211_X1 U16392 ( .C1(n14443), .C2(n19398), .A(n14442), .B(n14441), .ZN(
        P2_U2918) );
  MUX2_X1 U16393 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14444), .S(
        n14464), .Z(n16810) );
  NAND2_X1 U16394 ( .A1(n14446), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14447) );
  NAND2_X1 U16395 ( .A1(n11025), .A2(n14447), .ZN(n21670) );
  NAND2_X1 U16396 ( .A1(n11031), .A2(n21670), .ZN(n14457) );
  XNOR2_X1 U16397 ( .A(n14450), .B(n11335), .ZN(n14454) );
  XNOR2_X1 U16398 ( .A(n14451), .B(n11335), .ZN(n14452) );
  AOI22_X1 U16399 ( .A1(n14455), .A2(n14454), .B1(n14453), .B2(n14452), .ZN(
        n14456) );
  OAI21_X1 U16400 ( .B1(n16037), .B2(n14457), .A(n14456), .ZN(n14458) );
  AOI21_X1 U16401 ( .B1(n14445), .B2(n16037), .A(n14458), .ZN(n21674) );
  MUX2_X1 U16402 ( .A(n11335), .B(n21674), .S(n14464), .Z(n16812) );
  INV_X1 U16403 ( .A(n16812), .ZN(n14459) );
  NAND3_X1 U16404 ( .A1(n16810), .A2(n14459), .A3(n16839), .ZN(n14462) );
  AND2_X1 U16405 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21668), .ZN(n14468) );
  NAND2_X1 U16406 ( .A1(n14468), .A2(n14460), .ZN(n14461) );
  NAND2_X1 U16407 ( .A1(n14462), .A2(n14461), .ZN(n16824) );
  INV_X1 U16408 ( .A(n14463), .ZN(n16031) );
  NAND2_X1 U16409 ( .A1(n16824), .A2(n16031), .ZN(n14472) );
  OAI21_X1 U16410 ( .B1(n21484), .B2(n14234), .A(n14464), .ZN(n14467) );
  INV_X1 U16411 ( .A(n14464), .ZN(n16806) );
  AOI21_X1 U16412 ( .B1(n16806), .B2(n14465), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n14466) );
  NAND2_X1 U16413 ( .A1(n14467), .A2(n14466), .ZN(n14470) );
  NAND2_X1 U16414 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14468), .ZN(
        n14469) );
  NAND2_X1 U16415 ( .A1(n14470), .A2(n14469), .ZN(n16822) );
  INV_X1 U16416 ( .A(n16822), .ZN(n14471) );
  NAND2_X1 U16417 ( .A1(n14472), .A2(n14471), .ZN(n14476) );
  NOR2_X1 U16418 ( .A1(n21683), .A2(n21682), .ZN(n14473) );
  OAI21_X1 U16419 ( .B1(n14476), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14473), .ZN(
        n14475) );
  INV_X1 U16420 ( .A(n21682), .ZN(n14474) );
  NAND2_X1 U16421 ( .A1(n14475), .A2(n21871), .ZN(n16840) );
  NOR2_X1 U16422 ( .A1(n14476), .A2(n21682), .ZN(n21690) );
  NAND2_X1 U16423 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21930), .ZN(n14524) );
  INV_X1 U16424 ( .A(n14524), .ZN(n16029) );
  OAI22_X1 U16425 ( .A1(n11020), .A2(n22015), .B1(n14477), .B2(n16029), .ZN(
        n14478) );
  OAI21_X1 U16426 ( .B1(n21690), .B2(n14478), .A(n16840), .ZN(n14479) );
  OAI21_X1 U16427 ( .B1(n16840), .B2(n21975), .A(n14479), .ZN(P1_U3478) );
  OAI21_X1 U16428 ( .B1(n14481), .B2(n14480), .A(n14483), .ZN(n18349) );
  OAI222_X1 U16429 ( .A1(n14958), .A2(n19131), .B1(n18349), .B2(n19404), .C1(
        n17196), .C2(n16250), .ZN(P2_U2912) );
  XNOR2_X1 U16430 ( .A(n11083), .B(n14482), .ZN(n18337) );
  INV_X1 U16431 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17194) );
  OAI222_X1 U16432 ( .A1(n14958), .A2(n19352), .B1(n18337), .B2(n19404), .C1(
        n17194), .C2(n16250), .ZN(P2_U2913) );
  AOI21_X1 U16433 ( .B1(n14484), .B2(n14483), .A(n14486), .ZN(n18605) );
  INV_X1 U16434 ( .A(n18605), .ZN(n14485) );
  OAI222_X1 U16435 ( .A1(n14958), .A2(n16222), .B1(n14485), .B2(n19404), .C1(
        n12924), .C2(n16250), .ZN(P2_U2911) );
  OR2_X1 U16436 ( .A1(n14487), .A2(n14486), .ZN(n14488) );
  NAND2_X1 U16437 ( .A1(n14488), .A2(n15035), .ZN(n18366) );
  INV_X1 U16438 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17199) );
  OAI222_X1 U16439 ( .A1(n14958), .A2(n16212), .B1(n18366), .B2(n19404), .C1(
        n17199), .C2(n16250), .ZN(P2_U2910) );
  XOR2_X1 U16440 ( .A(n14489), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14494)
         );
  AND2_X1 U16441 ( .A1(n14501), .A2(n14490), .ZN(n14491) );
  OR2_X1 U16442 ( .A1(n14491), .A2(n14614), .ZN(n18323) );
  NOR2_X1 U16443 ( .A1(n18323), .A2(n16176), .ZN(n14492) );
  AOI21_X1 U16444 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n16176), .A(n14492), .ZN(
        n14493) );
  OAI21_X1 U16445 ( .B1(n14494), .B2(n16178), .A(n14493), .ZN(P2_U2882) );
  OR2_X1 U16446 ( .A1(n14496), .A2(n14495), .ZN(n14497) );
  NAND2_X1 U16447 ( .A1(n14489), .A2(n14497), .ZN(n19399) );
  NAND2_X1 U16448 ( .A1(n14499), .A2(n14498), .ZN(n14500) );
  NAND2_X1 U16449 ( .A1(n14501), .A2(n14500), .ZN(n18306) );
  MUX2_X1 U16450 ( .A(n18306), .B(n13273), .S(n16176), .Z(n14502) );
  OAI21_X1 U16451 ( .B1(n19399), .B2(n16178), .A(n14502), .ZN(P2_U2883) );
  INV_X1 U16452 ( .A(n14503), .ZN(n14504) );
  AOI21_X1 U16453 ( .B1(n14506), .B2(n14505), .A(n14504), .ZN(n14626) );
  INV_X1 U16454 ( .A(n14626), .ZN(n14731) );
  INV_X1 U16455 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U16456 ( .A1(n14508), .A2(n14507), .ZN(n14509) );
  NAND2_X1 U16457 ( .A1(n14533), .A2(n14509), .ZN(n21323) );
  OAI222_X1 U16458 ( .A1(n14731), .A2(n15659), .B1(n19911), .B2(n14719), .C1(
        n21323), .C2(n15657), .ZN(P1_U2870) );
  INV_X1 U16459 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21786) );
  INV_X1 U16460 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n14511) );
  OR2_X1 U16461 ( .A1(n15202), .A2(n14511), .ZN(n14513) );
  NAND2_X1 U16462 ( .A1(n15202), .A2(DATAI_1_), .ZN(n14512) );
  NAND2_X1 U16463 ( .A1(n14513), .A2(n14512), .ZN(n15715) );
  INV_X1 U16464 ( .A(n15715), .ZN(n21781) );
  OAI222_X1 U16465 ( .A1(n15725), .A2(n21472), .B1(n15260), .B2(n21786), .C1(
        n15259), .C2(n21781), .ZN(P1_U2903) );
  INV_X1 U16466 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21780) );
  OR2_X1 U16467 ( .A1(n15202), .A2(n19991), .ZN(n14515) );
  NAND2_X1 U16468 ( .A1(n15202), .A2(DATAI_0_), .ZN(n14514) );
  NAND2_X1 U16469 ( .A1(n14515), .A2(n14514), .ZN(n15721) );
  INV_X1 U16470 ( .A(n15721), .ZN(n21775) );
  OAI222_X1 U16471 ( .A1(n15725), .A2(n14516), .B1(n15260), .B2(n21780), .C1(
        n15259), .C2(n21775), .ZN(P1_U2904) );
  INV_X1 U16472 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21792) );
  OR2_X1 U16473 ( .A1(n15202), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14518) );
  INV_X1 U16474 ( .A(DATAI_2_), .ZN(n16854) );
  NAND2_X1 U16475 ( .A1(n15202), .A2(n16854), .ZN(n14517) );
  INV_X1 U16476 ( .A(n15709), .ZN(n21787) );
  OAI222_X1 U16477 ( .A1(n14731), .A2(n15725), .B1(n15260), .B2(n21792), .C1(
        n15259), .C2(n21787), .ZN(P1_U2902) );
  NAND2_X1 U16478 ( .A1(n14520), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16022) );
  INV_X1 U16479 ( .A(n16022), .ZN(n16025) );
  NAND2_X1 U16480 ( .A1(n21989), .A2(n16025), .ZN(n22013) );
  INV_X1 U16481 ( .A(n22013), .ZN(n14523) );
  NOR2_X1 U16482 ( .A1(n14519), .A2(n14522), .ZN(n14546) );
  AND2_X1 U16483 ( .A1(n14546), .A2(n14520), .ZN(n14633) );
  NAND2_X1 U16484 ( .A1(n14633), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14631) );
  OAI21_X1 U16485 ( .B1(n14523), .B2(n14521), .A(n14631), .ZN(n14525) );
  AOI22_X1 U16486 ( .A1(n14525), .A2(n21982), .B1(n14524), .B2(n14445), .ZN(
        n14528) );
  INV_X1 U16487 ( .A(n16840), .ZN(n14527) );
  NAND2_X1 U16488 ( .A1(n14527), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14526) );
  OAI21_X1 U16489 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(P1_U3475) );
  OAI21_X1 U16490 ( .B1(n14531), .B2(n14530), .A(n14529), .ZN(n14900) );
  AND2_X1 U16491 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  NOR2_X1 U16492 ( .A1(n14706), .A2(n14534), .ZN(n21341) );
  INV_X1 U16493 ( .A(n19911), .ZN(n15650) );
  AOI22_X1 U16494 ( .A1(n21341), .A2(n13472), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15650), .ZN(n14535) );
  OAI21_X1 U16495 ( .B1(n14900), .B2(n15659), .A(n14535), .ZN(P1_U2869) );
  XNOR2_X1 U16496 ( .A(n14536), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U16497 ( .A1(n14538), .A2(n14537), .ZN(n14541) );
  INV_X1 U16498 ( .A(n14539), .ZN(n14540) );
  NAND2_X1 U16499 ( .A1(n14541), .A2(n14540), .ZN(n18348) );
  MUX2_X1 U16500 ( .A(n13277), .B(n18348), .S(n16127), .Z(n14542) );
  OAI21_X1 U16501 ( .B1(n14543), .B2(n16178), .A(n14542), .ZN(P2_U2880) );
  INV_X1 U16502 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20046) );
  OAI22_X1 U16503 ( .A1(n20046), .A2(n14601), .B1(n12297), .B2(n14600), .ZN(
        n22199) );
  INV_X1 U16504 ( .A(n22199), .ZN(n22208) );
  INV_X1 U16505 ( .A(n14520), .ZN(n14545) );
  NAND2_X1 U16506 ( .A1(n14546), .A2(n14545), .ZN(n14551) );
  NAND3_X1 U16507 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21965), .A3(
        n12217), .ZN(n14976) );
  INV_X1 U16508 ( .A(n14976), .ZN(n14550) );
  INV_X1 U16509 ( .A(n14548), .ZN(n21976) );
  NOR2_X1 U16510 ( .A1(n21975), .A2(n14976), .ZN(n14558) );
  AOI21_X1 U16511 ( .B1(n21910), .B2(n21976), .A(n14558), .ZN(n14553) );
  OAI211_X1 U16512 ( .C1(n14551), .C2(n21936), .A(n21982), .B(n14553), .ZN(
        n14549) );
  NAND2_X1 U16513 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14561) );
  INV_X1 U16514 ( .A(DATAI_21_), .ZN(n14552) );
  INV_X1 U16515 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20029) );
  OAI22_X1 U16516 ( .A1(n14552), .A2(n14600), .B1(n20029), .B2(n14601), .ZN(
        n22205) );
  OAI22_X1 U16517 ( .A1(n14553), .A2(n22015), .B1(n14976), .B2(n22008), .ZN(
        n14554) );
  INV_X1 U16518 ( .A(n14554), .ZN(n14605) );
  OR2_X1 U16519 ( .A1(n15202), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14556) );
  INV_X1 U16520 ( .A(DATAI_5_), .ZN(n16990) );
  NAND2_X1 U16521 ( .A1(n15202), .A2(n16990), .ZN(n14555) );
  AND2_X1 U16522 ( .A1(n14556), .A2(n14555), .ZN(n21805) );
  NAND2_X1 U16523 ( .A1(n14603), .A2(n12238), .ZN(n22192) );
  INV_X1 U16524 ( .A(n14558), .ZN(n14604) );
  OAI22_X1 U16525 ( .A1(n14605), .A2(n22196), .B1(n22192), .B2(n14604), .ZN(
        n14559) );
  AOI21_X1 U16526 ( .B1(n14607), .B2(n22205), .A(n14559), .ZN(n14560) );
  OAI211_X1 U16527 ( .C1(n22208), .C2(n14979), .A(n14561), .B(n14560), .ZN(
        P1_U3078) );
  INV_X1 U16528 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20044) );
  OAI22_X1 U16529 ( .A1(n20044), .A2(n14601), .B1(n16951), .B2(n14600), .ZN(
        n22162) );
  INV_X1 U16530 ( .A(n22162), .ZN(n22171) );
  NAND2_X1 U16531 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14567) );
  INV_X1 U16532 ( .A(DATAI_20_), .ZN(n16880) );
  INV_X1 U16533 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20027) );
  OAI22_X1 U16534 ( .A1(n16880), .A2(n14600), .B1(n20027), .B2(n14601), .ZN(
        n22168) );
  OR2_X1 U16535 ( .A1(n15202), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14563) );
  INV_X1 U16536 ( .A(DATAI_4_), .ZN(n16992) );
  NAND2_X1 U16537 ( .A1(n15202), .A2(n16992), .ZN(n14562) );
  AND2_X1 U16538 ( .A1(n14563), .A2(n14562), .ZN(n15697) );
  NAND2_X1 U16539 ( .A1(n14603), .A2(n14564), .ZN(n22155) );
  OAI22_X1 U16540 ( .A1(n14605), .A2(n22159), .B1(n22155), .B2(n14604), .ZN(
        n14565) );
  AOI21_X1 U16541 ( .B1(n14607), .B2(n22168), .A(n14565), .ZN(n14566) );
  OAI211_X1 U16542 ( .C1(n22171), .C2(n14979), .A(n14567), .B(n14566), .ZN(
        P1_U3077) );
  OAI22_X1 U16543 ( .A1(n14066), .A2(n14601), .B1(n16949), .B2(n14600), .ZN(
        n22236) );
  INV_X1 U16544 ( .A(n22236), .ZN(n22245) );
  NAND2_X1 U16545 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14573) );
  INV_X1 U16546 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20031) );
  INV_X1 U16547 ( .A(DATAI_22_), .ZN(n16961) );
  OAI22_X1 U16548 ( .A1(n20031), .A2(n14601), .B1(n16961), .B2(n14600), .ZN(
        n22242) );
  OR2_X1 U16549 ( .A1(n15202), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14569) );
  INV_X1 U16550 ( .A(DATAI_6_), .ZN(n16856) );
  NAND2_X1 U16551 ( .A1(n15202), .A2(n16856), .ZN(n14568) );
  AND2_X1 U16552 ( .A1(n14569), .A2(n14568), .ZN(n15686) );
  NAND2_X1 U16553 ( .A1(n14603), .A2(n14570), .ZN(n22229) );
  OAI22_X1 U16554 ( .A1(n14605), .A2(n22233), .B1(n22229), .B2(n14604), .ZN(
        n14571) );
  AOI21_X1 U16555 ( .B1(n14607), .B2(n22242), .A(n14571), .ZN(n14572) );
  OAI211_X1 U16556 ( .C1(n22245), .C2(n14979), .A(n14573), .B(n14572), .ZN(
        P1_U3079) );
  INV_X1 U16557 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20049) );
  OAI22_X1 U16558 ( .A1(n14574), .A2(n14600), .B1(n20049), .B2(n14601), .ZN(
        n22320) );
  INV_X1 U16559 ( .A(n22320), .ZN(n22336) );
  NAND2_X1 U16560 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14581) );
  INV_X1 U16561 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20033) );
  INV_X1 U16562 ( .A(DATAI_23_), .ZN(n16960) );
  OAI22_X1 U16563 ( .A1(n20033), .A2(n14601), .B1(n16960), .B2(n14600), .ZN(
        n22332) );
  INV_X1 U16564 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n14575) );
  OR2_X1 U16565 ( .A1(n15202), .A2(n14575), .ZN(n14577) );
  NAND2_X1 U16566 ( .A1(n15202), .A2(DATAI_7_), .ZN(n14576) );
  NAND2_X1 U16567 ( .A1(n14577), .A2(n14576), .ZN(n15681) );
  NAND2_X1 U16568 ( .A1(n14603), .A2(n14578), .ZN(n22304) );
  OAI22_X1 U16569 ( .A1(n14605), .A2(n22310), .B1(n22304), .B2(n14604), .ZN(
        n14579) );
  AOI21_X1 U16570 ( .B1(n14607), .B2(n22332), .A(n14579), .ZN(n14580) );
  OAI211_X1 U16571 ( .C1(n22336), .C2(n14979), .A(n14581), .B(n14580), .ZN(
        P1_U3080) );
  INV_X1 U16572 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20042) );
  INV_X1 U16573 ( .A(DATAI_27_), .ZN(n14582) );
  OAI22_X1 U16574 ( .A1(n20042), .A2(n14601), .B1(n14582), .B2(n14600), .ZN(
        n22125) );
  INV_X1 U16575 ( .A(n22125), .ZN(n22134) );
  NAND2_X1 U16576 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14588) );
  INV_X1 U16577 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20025) );
  INV_X1 U16578 ( .A(DATAI_19_), .ZN(n16944) );
  OAI22_X1 U16579 ( .A1(n20025), .A2(n14601), .B1(n16944), .B2(n14600), .ZN(
        n22131) );
  INV_X1 U16580 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n14583) );
  OR2_X1 U16581 ( .A1(n15202), .A2(n14583), .ZN(n14585) );
  NAND2_X1 U16582 ( .A1(n15202), .A2(DATAI_3_), .ZN(n14584) );
  NAND2_X1 U16583 ( .A1(n14585), .A2(n14584), .ZN(n15703) );
  NAND2_X1 U16584 ( .A1(n14603), .A2(n11571), .ZN(n22118) );
  OAI22_X1 U16585 ( .A1(n14605), .A2(n22122), .B1(n22118), .B2(n14604), .ZN(
        n14586) );
  AOI21_X1 U16586 ( .B1(n14607), .B2(n22131), .A(n14586), .ZN(n14587) );
  OAI211_X1 U16587 ( .C1(n22134), .C2(n14979), .A(n14588), .B(n14587), .ZN(
        P1_U3076) );
  INV_X1 U16588 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20040) );
  INV_X1 U16589 ( .A(DATAI_26_), .ZN(n14589) );
  OAI22_X1 U16590 ( .A1(n20040), .A2(n14601), .B1(n14589), .B2(n14600), .ZN(
        n22088) );
  INV_X1 U16591 ( .A(n22088), .ZN(n22097) );
  NAND2_X1 U16592 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14592) );
  INV_X1 U16593 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20023) );
  INV_X1 U16594 ( .A(DATAI_18_), .ZN(n16963) );
  NAND2_X1 U16595 ( .A1(n14603), .A2(n11551), .ZN(n22081) );
  OAI22_X1 U16596 ( .A1(n14605), .A2(n22085), .B1(n22081), .B2(n14604), .ZN(
        n14590) );
  AOI21_X1 U16597 ( .B1(n14607), .B2(n22094), .A(n14590), .ZN(n14591) );
  OAI211_X1 U16598 ( .C1(n22097), .C2(n14979), .A(n14592), .B(n14591), .ZN(
        P1_U3075) );
  INV_X1 U16599 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20037) );
  INV_X1 U16600 ( .A(DATAI_25_), .ZN(n16868) );
  OAI22_X1 U16601 ( .A1(n20037), .A2(n14601), .B1(n16868), .B2(n14600), .ZN(
        n22050) );
  INV_X1 U16602 ( .A(n22050), .ZN(n22059) );
  NAND2_X1 U16603 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14595) );
  INV_X1 U16604 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20021) );
  INV_X1 U16605 ( .A(DATAI_17_), .ZN(n16964) );
  NAND2_X1 U16606 ( .A1(n14603), .A2(n13348), .ZN(n22043) );
  OAI22_X1 U16607 ( .A1(n14605), .A2(n22047), .B1(n22043), .B2(n14604), .ZN(
        n14593) );
  AOI21_X1 U16608 ( .B1(n14607), .B2(n22056), .A(n14593), .ZN(n14594) );
  OAI211_X1 U16609 ( .C1(n22059), .C2(n14979), .A(n14595), .B(n14594), .ZN(
        P1_U3074) );
  OR2_X1 U16610 ( .A1(n14596), .A2(n11067), .ZN(n14597) );
  NAND2_X1 U16611 ( .A1(n14597), .A2(n16642), .ZN(n18370) );
  INV_X1 U16612 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17204) );
  OAI222_X1 U16613 ( .A1(n14958), .A2(n14598), .B1(n18370), .B2(n19404), .C1(
        n17204), .C2(n16250), .ZN(P2_U2908) );
  INV_X1 U16614 ( .A(DATAI_24_), .ZN(n16946) );
  INV_X1 U16615 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20035) );
  OAI22_X1 U16616 ( .A1(n16946), .A2(n14600), .B1(n20035), .B2(n14601), .ZN(
        n22000) );
  NAND2_X1 U16617 ( .A1(n14599), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14609) );
  INV_X1 U16618 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20019) );
  INV_X1 U16619 ( .A(DATAI_16_), .ZN(n16943) );
  OAI22_X1 U16620 ( .A1(n20019), .A2(n14601), .B1(n16943), .B2(n14600), .ZN(
        n22019) );
  NAND2_X1 U16621 ( .A1(n14603), .A2(n11553), .ZN(n21966) );
  OAI22_X1 U16622 ( .A1(n14605), .A2(n21974), .B1(n21966), .B2(n14604), .ZN(
        n14606) );
  AOI21_X1 U16623 ( .B1(n14607), .B2(n22019), .A(n14606), .ZN(n14608) );
  OAI211_X1 U16624 ( .C1(n22022), .C2(n14979), .A(n14609), .B(n14608), .ZN(
        P1_U3073) );
  NOR2_X1 U16625 ( .A1(n14489), .A2(n14610), .ZN(n14612) );
  INV_X1 U16626 ( .A(n14536), .ZN(n14611) );
  OAI211_X1 U16627 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14612), .A(
        n14611), .B(n16169), .ZN(n14617) );
  OR2_X1 U16628 ( .A1(n14614), .A2(n14613), .ZN(n14615) );
  AND2_X1 U16629 ( .A1(n14615), .A2(n14537), .ZN(n18335) );
  NAND2_X1 U16630 ( .A1(n18335), .A2(n16127), .ZN(n14616) );
  OAI211_X1 U16631 ( .C1(n16127), .C2(n14618), .A(n14617), .B(n14616), .ZN(
        P2_U2881) );
  INV_X1 U16632 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n21798) );
  INV_X1 U16633 ( .A(n15703), .ZN(n21793) );
  OAI222_X1 U16634 ( .A1(n15725), .A2(n14900), .B1(n15260), .B2(n21798), .C1(
        n15259), .C2(n21793), .ZN(P1_U2901) );
  AOI22_X1 U16635 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21457), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14619) );
  OAI21_X1 U16636 ( .B1(n19982), .B2(n14723), .A(n14619), .ZN(n14625) );
  NOR2_X1 U16637 ( .A1(n14621), .A2(n14620), .ZN(n21321) );
  INV_X1 U16638 ( .A(n14622), .ZN(n14623) );
  NOR3_X1 U16639 ( .A1(n21321), .A2(n14623), .A3(n21667), .ZN(n14624) );
  AOI211_X1 U16640 ( .C1(n19979), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n14627) );
  INV_X1 U16641 ( .A(n14627), .ZN(P1_U2997) );
  NOR2_X1 U16642 ( .A1(n22007), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14635) );
  INV_X1 U16643 ( .A(n11014), .ZN(n14629) );
  NAND2_X1 U16644 ( .A1(n14629), .A2(n11698), .ZN(n21898) );
  INV_X1 U16645 ( .A(n21898), .ZN(n22005) );
  INV_X1 U16646 ( .A(n14662), .ZN(n14630) );
  AOI21_X1 U16647 ( .B1(n21910), .B2(n22005), .A(n14630), .ZN(n14634) );
  NAND3_X1 U16648 ( .A1(n14631), .A2(n21982), .A3(n14634), .ZN(n14632) );
  NAND2_X1 U16649 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14641) );
  INV_X1 U16650 ( .A(n14634), .ZN(n14638) );
  INV_X1 U16651 ( .A(n14635), .ZN(n14636) );
  NOR2_X1 U16652 ( .A1(n22008), .A2(n14636), .ZN(n14637) );
  AOI21_X1 U16653 ( .B1(n14638), .B2(n21935), .A(n14637), .ZN(n14663) );
  OAI22_X1 U16654 ( .A1(n14663), .A2(n22122), .B1(n14662), .B2(n22118), .ZN(
        n14639) );
  AOI21_X1 U16655 ( .B1(n22286), .B2(n22131), .A(n14639), .ZN(n14640) );
  OAI211_X1 U16656 ( .C1(n14660), .C2(n22134), .A(n14641), .B(n14640), .ZN(
        P1_U3092) );
  NAND2_X1 U16657 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14644) );
  OAI22_X1 U16658 ( .A1(n14663), .A2(n22047), .B1(n14662), .B2(n22043), .ZN(
        n14642) );
  AOI21_X1 U16659 ( .B1(n22286), .B2(n22056), .A(n14642), .ZN(n14643) );
  OAI211_X1 U16660 ( .C1(n14660), .C2(n22059), .A(n14644), .B(n14643), .ZN(
        P1_U3090) );
  NAND2_X1 U16661 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14647) );
  OAI22_X1 U16662 ( .A1(n14663), .A2(n22159), .B1(n14662), .B2(n22155), .ZN(
        n14645) );
  AOI21_X1 U16663 ( .B1(n22286), .B2(n22168), .A(n14645), .ZN(n14646) );
  OAI211_X1 U16664 ( .C1(n14660), .C2(n22171), .A(n14647), .B(n14646), .ZN(
        P1_U3093) );
  NAND2_X1 U16665 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14650) );
  OAI22_X1 U16666 ( .A1(n14663), .A2(n22233), .B1(n14662), .B2(n22229), .ZN(
        n14648) );
  AOI21_X1 U16667 ( .B1(n22286), .B2(n22242), .A(n14648), .ZN(n14649) );
  OAI211_X1 U16668 ( .C1(n14660), .C2(n22245), .A(n14650), .B(n14649), .ZN(
        P1_U3095) );
  NAND2_X1 U16669 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14653) );
  OAI22_X1 U16670 ( .A1(n14663), .A2(n22196), .B1(n14662), .B2(n22192), .ZN(
        n14651) );
  AOI21_X1 U16671 ( .B1(n22286), .B2(n22205), .A(n14651), .ZN(n14652) );
  OAI211_X1 U16672 ( .C1(n14660), .C2(n22208), .A(n14653), .B(n14652), .ZN(
        P1_U3094) );
  NAND2_X1 U16673 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14656) );
  OAI22_X1 U16674 ( .A1(n14663), .A2(n22085), .B1(n14662), .B2(n22081), .ZN(
        n14654) );
  AOI21_X1 U16675 ( .B1(n22286), .B2(n22094), .A(n14654), .ZN(n14655) );
  OAI211_X1 U16676 ( .C1(n14660), .C2(n22097), .A(n14656), .B(n14655), .ZN(
        P1_U3091) );
  NAND2_X1 U16677 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14659) );
  OAI22_X1 U16678 ( .A1(n14663), .A2(n22310), .B1(n14662), .B2(n22304), .ZN(
        n14657) );
  AOI21_X1 U16679 ( .B1(n22286), .B2(n22332), .A(n14657), .ZN(n14658) );
  OAI211_X1 U16680 ( .C1(n14660), .C2(n22336), .A(n14659), .B(n14658), .ZN(
        P1_U3096) );
  INV_X1 U16681 ( .A(n22286), .ZN(n14667) );
  INV_X1 U16682 ( .A(n22019), .ZN(n22003) );
  NAND2_X1 U16683 ( .A1(n14661), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14666) );
  OAI22_X1 U16684 ( .A1(n14663), .A2(n21974), .B1(n14662), .B2(n21966), .ZN(
        n14664) );
  AOI21_X1 U16685 ( .B1(n22279), .B2(n22000), .A(n14664), .ZN(n14665) );
  OAI211_X1 U16686 ( .C1(n14667), .C2(n22003), .A(n14666), .B(n14665), .ZN(
        P1_U3089) );
  INV_X1 U16687 ( .A(n14668), .ZN(n14669) );
  NOR2_X1 U16688 ( .A1(n14670), .A2(n14669), .ZN(n14864) );
  INV_X1 U16689 ( .A(n17151), .ZN(n15104) );
  XNOR2_X1 U16690 ( .A(n14864), .B(n15104), .ZN(n14863) );
  XNOR2_X1 U16691 ( .A(n14863), .B(n19254), .ZN(n14671) );
  NAND2_X1 U16692 ( .A1(n14671), .A2(n19620), .ZN(n14673) );
  AOI22_X1 U16693 ( .A1(n19619), .A2(n17151), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19613), .ZN(n14672) );
  OAI211_X1 U16694 ( .C1(n19532), .C2(n14958), .A(n14673), .B(n14672), .ZN(
        P2_U2917) );
  INV_X1 U16695 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17208) );
  XNOR2_X1 U16696 ( .A(n14675), .B(n14674), .ZN(n18402) );
  OAI222_X1 U16697 ( .A1(n14958), .A2(n14676), .B1(n16250), .B2(n17208), .C1(
        n19404), .C2(n18402), .ZN(P2_U2906) );
  NAND3_X1 U16698 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21922), .ZN(n21947) );
  INV_X1 U16699 ( .A(n21947), .ZN(n14684) );
  INV_X1 U16700 ( .A(n14519), .ZN(n14677) );
  INV_X1 U16701 ( .A(n21961), .ZN(n16028) );
  NAND2_X1 U16702 ( .A1(n21943), .A2(n22005), .ZN(n14679) );
  NOR2_X1 U16703 ( .A1(n21975), .A2(n21947), .ZN(n14758) );
  INV_X1 U16704 ( .A(n14758), .ZN(n14678) );
  NAND2_X1 U16705 ( .A1(n14679), .A2(n14678), .ZN(n14683) );
  INV_X1 U16706 ( .A(n14683), .ZN(n14680) );
  OAI211_X1 U16707 ( .C1(n21939), .C2(n16022), .A(n21982), .B(n14680), .ZN(
        n14681) );
  OAI211_X1 U16708 ( .C1(n21935), .C2(n14684), .A(n14681), .B(n22017), .ZN(
        n14682) );
  INV_X1 U16709 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U16710 ( .A1(n14520), .A2(n11020), .ZN(n21987) );
  NAND2_X1 U16711 ( .A1(n14520), .A2(n21865), .ZN(n21866) );
  INV_X1 U16712 ( .A(n22306), .ZN(n14745) );
  INV_X1 U16713 ( .A(n22242), .ZN(n22239) );
  INV_X1 U16714 ( .A(n22233), .ZN(n22241) );
  NAND2_X1 U16715 ( .A1(n14683), .A2(n21982), .ZN(n14686) );
  NAND2_X1 U16716 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14684), .ZN(n14685) );
  NAND2_X1 U16717 ( .A1(n14686), .A2(n14685), .ZN(n14757) );
  AOI22_X1 U16718 ( .A1(n22240), .A2(n14758), .B1(n22241), .B2(n14757), .ZN(
        n14687) );
  OAI21_X1 U16719 ( .B1(n14745), .B2(n22239), .A(n14687), .ZN(n14688) );
  AOI21_X1 U16720 ( .B1(n22236), .B2(n22297), .A(n14688), .ZN(n14689) );
  OAI21_X1 U16721 ( .B1(n14764), .B2(n14690), .A(n14689), .ZN(P1_U3127) );
  INV_X1 U16722 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14694) );
  INV_X1 U16723 ( .A(n22332), .ZN(n22325) );
  AOI22_X1 U16724 ( .A1(n22327), .A2(n14758), .B1(n22329), .B2(n14757), .ZN(
        n14691) );
  OAI21_X1 U16725 ( .B1(n14745), .B2(n22325), .A(n14691), .ZN(n14692) );
  AOI21_X1 U16726 ( .B1(n22320), .B2(n22297), .A(n14692), .ZN(n14693) );
  OAI21_X1 U16727 ( .B1(n14764), .B2(n14694), .A(n14693), .ZN(P1_U3128) );
  INV_X1 U16728 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n18354) );
  OAI211_X1 U16729 ( .C1(n14695), .C2(n14697), .A(n14696), .B(n16169), .ZN(
        n14704) );
  NAND2_X1 U16730 ( .A1(n14699), .A2(n14698), .ZN(n14702) );
  INV_X1 U16731 ( .A(n14700), .ZN(n14701) );
  AND2_X1 U16732 ( .A1(n14702), .A2(n14701), .ZN(n18361) );
  NAND2_X1 U16733 ( .A1(n16127), .A2(n18361), .ZN(n14703) );
  OAI211_X1 U16734 ( .C1(n16127), .C2(n18354), .A(n14704), .B(n14703), .ZN(
        P2_U2878) );
  OR2_X1 U16735 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  AND2_X1 U16736 ( .A1(n19905), .A2(n14707), .ZN(n21332) );
  INV_X1 U16737 ( .A(n21332), .ZN(n21482) );
  XOR2_X1 U16738 ( .A(n14529), .B(n14708), .Z(n21490) );
  INV_X1 U16739 ( .A(n21490), .ZN(n14710) );
  INV_X1 U16740 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14709) );
  OAI222_X1 U16741 ( .A1(n21482), .A2(n15657), .B1(n15659), .B2(n14710), .C1(
        n14709), .C2(n19911), .ZN(P1_U2868) );
  INV_X1 U16742 ( .A(n15697), .ZN(n21799) );
  INV_X1 U16743 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21804) );
  OAI222_X1 U16744 ( .A1(n15259), .A2(n21799), .B1(n15725), .B2(n14710), .C1(
        n21804), .C2(n15260), .ZN(P1_U2900) );
  INV_X1 U16745 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14714) );
  INV_X1 U16746 ( .A(n22205), .ZN(n22202) );
  INV_X1 U16747 ( .A(n22196), .ZN(n22204) );
  AOI22_X1 U16748 ( .A1(n22203), .A2(n14758), .B1(n22204), .B2(n14757), .ZN(
        n14711) );
  OAI21_X1 U16749 ( .B1(n14745), .B2(n22202), .A(n14711), .ZN(n14712) );
  AOI21_X1 U16750 ( .B1(n22199), .B2(n22297), .A(n14712), .ZN(n14713) );
  OAI21_X1 U16751 ( .B1(n14764), .B2(n14714), .A(n14713), .ZN(P1_U3126) );
  NAND2_X1 U16752 ( .A1(n21286), .A2(n14715), .ZN(n14716) );
  NAND2_X1 U16753 ( .A1(n21591), .A2(n14716), .ZN(n21497) );
  INV_X1 U16754 ( .A(n21497), .ZN(n21471) );
  NAND2_X1 U16755 ( .A1(n21286), .A2(n14717), .ZN(n21483) );
  INV_X1 U16756 ( .A(n21483), .ZN(n14897) );
  INV_X1 U16757 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14718) );
  NAND3_X1 U16758 ( .A1(n21562), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n14718), 
        .ZN(n14728) );
  OAI21_X1 U16759 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21539), .A(n15559), .ZN(
        n14889) );
  OAI22_X1 U16760 ( .A1(n14719), .A2(n21649), .B1(n21665), .B2(n21323), .ZN(
        n14720) );
  AOI21_X1 U16761 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n14889), .A(n14720), .ZN(
        n14727) );
  AND2_X1 U16762 ( .A1(n14721), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14722) );
  INV_X1 U16763 ( .A(n14723), .ZN(n14724) );
  NAND2_X1 U16764 ( .A1(n21659), .A2(n14724), .ZN(n14726) );
  NAND2_X1 U16765 ( .A1(n21652), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14725) );
  NAND4_X1 U16766 ( .A1(n14728), .A2(n14727), .A3(n14726), .A4(n14725), .ZN(
        n14729) );
  AOI21_X1 U16767 ( .B1(n21961), .B2(n14897), .A(n14729), .ZN(n14730) );
  OAI21_X1 U16768 ( .B1(n14731), .B2(n21471), .A(n14730), .ZN(P1_U2838) );
  INV_X1 U16769 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14735) );
  INV_X1 U16770 ( .A(n22056), .ZN(n22053) );
  INV_X1 U16771 ( .A(n22047), .ZN(n22055) );
  AOI22_X1 U16772 ( .A1(n22054), .A2(n14758), .B1(n22055), .B2(n14757), .ZN(
        n14732) );
  OAI21_X1 U16773 ( .B1(n14745), .B2(n22053), .A(n14732), .ZN(n14733) );
  AOI21_X1 U16774 ( .B1(n22050), .B2(n22297), .A(n14733), .ZN(n14734) );
  OAI21_X1 U16775 ( .B1(n14764), .B2(n14735), .A(n14734), .ZN(P1_U3122) );
  INV_X1 U16776 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14739) );
  INV_X1 U16777 ( .A(n22094), .ZN(n22091) );
  INV_X1 U16778 ( .A(n22085), .ZN(n22093) );
  AOI22_X1 U16779 ( .A1(n22092), .A2(n14758), .B1(n22093), .B2(n14757), .ZN(
        n14736) );
  OAI21_X1 U16780 ( .B1(n14745), .B2(n22091), .A(n14736), .ZN(n14737) );
  AOI21_X1 U16781 ( .B1(n22088), .B2(n22297), .A(n14737), .ZN(n14738) );
  OAI21_X1 U16782 ( .B1(n14764), .B2(n14739), .A(n14738), .ZN(P1_U3123) );
  INV_X1 U16783 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14743) );
  INV_X1 U16784 ( .A(n22168), .ZN(n22165) );
  INV_X1 U16785 ( .A(n22159), .ZN(n22167) );
  AOI22_X1 U16786 ( .A1(n22166), .A2(n14758), .B1(n22167), .B2(n14757), .ZN(
        n14740) );
  OAI21_X1 U16787 ( .B1(n14745), .B2(n22165), .A(n14740), .ZN(n14741) );
  AOI21_X1 U16788 ( .B1(n22162), .B2(n22297), .A(n14741), .ZN(n14742) );
  OAI21_X1 U16789 ( .B1(n14764), .B2(n14743), .A(n14742), .ZN(P1_U3125) );
  INV_X1 U16790 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14748) );
  INV_X1 U16791 ( .A(n22131), .ZN(n22128) );
  INV_X1 U16792 ( .A(n22122), .ZN(n22130) );
  AOI22_X1 U16793 ( .A1(n22129), .A2(n14758), .B1(n22130), .B2(n14757), .ZN(
        n14744) );
  OAI21_X1 U16794 ( .B1(n14745), .B2(n22128), .A(n14744), .ZN(n14746) );
  AOI21_X1 U16795 ( .B1(n22125), .B2(n22297), .A(n14746), .ZN(n14747) );
  OAI21_X1 U16796 ( .B1(n14764), .B2(n14748), .A(n14747), .ZN(P1_U3124) );
  OAI21_X1 U16797 ( .B1(n14749), .B2(n14751), .A(n14750), .ZN(n14752) );
  INV_X1 U16798 ( .A(n14752), .ZN(n21343) );
  NAND2_X1 U16799 ( .A1(n21343), .A2(n19978), .ZN(n14756) );
  INV_X1 U16800 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14753) );
  NOR2_X1 U16801 ( .A1(n21616), .A2(n14753), .ZN(n21340) );
  NOR2_X1 U16802 ( .A1(n19982), .A2(n14888), .ZN(n14754) );
  AOI211_X1 U16803 ( .C1(n19976), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n21340), .B(n14754), .ZN(n14755) );
  OAI211_X1 U16804 ( .C1(n19947), .C2(n14900), .A(n14756), .B(n14755), .ZN(
        P1_U2996) );
  INV_X1 U16805 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14763) );
  INV_X1 U16806 ( .A(n22297), .ZN(n14760) );
  INV_X1 U16807 ( .A(n21974), .ZN(n22011) );
  AOI22_X1 U16808 ( .A1(n22010), .A2(n14758), .B1(n22011), .B2(n14757), .ZN(
        n14759) );
  OAI21_X1 U16809 ( .B1(n14760), .B2(n22022), .A(n14759), .ZN(n14761) );
  AOI21_X1 U16810 ( .B1(n22019), .B2(n22306), .A(n14761), .ZN(n14762) );
  OAI21_X1 U16811 ( .B1(n14764), .B2(n14763), .A(n14762), .ZN(P1_U3121) );
  INV_X1 U16812 ( .A(n14765), .ZN(n14851) );
  INV_X1 U16813 ( .A(n14785), .ZN(n14815) );
  NAND2_X1 U16814 ( .A1(n14806), .A2(n12305), .ZN(n14771) );
  NAND2_X1 U16815 ( .A1(n14767), .A2(n14766), .ZN(n14781) );
  OAI21_X1 U16816 ( .B1(n14769), .B2(n14768), .A(n14781), .ZN(n14770) );
  NAND2_X1 U16817 ( .A1(n14771), .A2(n14770), .ZN(n14772) );
  AOI21_X1 U16818 ( .B1(n11028), .B2(n14815), .A(n14772), .ZN(n16758) );
  INV_X1 U16819 ( .A(n14773), .ZN(n14775) );
  NOR2_X1 U16820 ( .A1(n13249), .A2(n14831), .ZN(n14774) );
  NAND2_X1 U16821 ( .A1(n14775), .A2(n14774), .ZN(n14780) );
  INV_X1 U16822 ( .A(n14776), .ZN(n14778) );
  AND4_X1 U16823 ( .A1(n14780), .A2(n14779), .A3(n14778), .A4(n14777), .ZN(
        n15110) );
  INV_X1 U16824 ( .A(n16758), .ZN(n14786) );
  INV_X1 U16825 ( .A(n14781), .ZN(n14783) );
  INV_X1 U16826 ( .A(n14806), .ZN(n14782) );
  MUX2_X1 U16827 ( .A(n14783), .B(n14782), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14784) );
  OAI21_X1 U16828 ( .B1(n15161), .B2(n14785), .A(n14784), .ZN(n15115) );
  AOI211_X1 U16829 ( .C1(n14786), .C2(n19302), .A(n17147), .B(n15115), .ZN(
        n14787) );
  AOI211_X1 U16830 ( .C1(n16758), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15110), .B(n14787), .ZN(n14802) );
  NAND2_X1 U16831 ( .A1(n15096), .A2(n14815), .ZN(n14797) );
  INV_X1 U16832 ( .A(n12538), .ZN(n14788) );
  NAND2_X1 U16833 ( .A1(n14788), .A2(n14798), .ZN(n14808) );
  INV_X1 U16834 ( .A(n14808), .ZN(n14794) );
  NAND2_X1 U16835 ( .A1(n14789), .A2(n15481), .ZN(n14807) );
  OR2_X1 U16836 ( .A1(n14825), .A2(n14819), .ZN(n14804) );
  NAND2_X1 U16837 ( .A1(n15481), .A2(n14808), .ZN(n14790) );
  NAND2_X1 U16838 ( .A1(n14804), .A2(n14790), .ZN(n14793) );
  NAND2_X1 U16839 ( .A1(n14806), .A2(n14791), .ZN(n14792) );
  OAI211_X1 U16840 ( .C1(n14794), .C2(n14807), .A(n14793), .B(n14792), .ZN(
        n14795) );
  INV_X1 U16841 ( .A(n14795), .ZN(n14796) );
  NAND2_X1 U16842 ( .A1(n14797), .A2(n14796), .ZN(n15146) );
  OR2_X1 U16843 ( .A1(n15146), .A2(n15110), .ZN(n14800) );
  NAND2_X1 U16844 ( .A1(n15110), .A2(n14798), .ZN(n14799) );
  NAND2_X1 U16845 ( .A1(n14800), .A2(n14799), .ZN(n14843) );
  NOR2_X1 U16846 ( .A1(n14843), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14801) );
  OAI22_X1 U16847 ( .A1(n14802), .A2(n14801), .B1(n17156), .B2(n15146), .ZN(
        n14818) );
  AOI22_X1 U16848 ( .A1(n14804), .A2(n14808), .B1(n13886), .B2(n14806), .ZN(
        n14811) );
  INV_X1 U16849 ( .A(n13886), .ZN(n14805) );
  NAND2_X1 U16850 ( .A1(n14806), .A2(n14805), .ZN(n14809) );
  AND3_X1 U16851 ( .A1(n14809), .A2(n14808), .A3(n14807), .ZN(n14810) );
  MUX2_X1 U16852 ( .A(n14811), .B(n14810), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14813) );
  NAND2_X1 U16853 ( .A1(n14813), .A2(n11281), .ZN(n14814) );
  AOI21_X1 U16854 ( .B1(n14803), .B2(n14815), .A(n14814), .ZN(n16760) );
  INV_X1 U16855 ( .A(n15110), .ZN(n14816) );
  MUX2_X1 U16856 ( .A(n12373), .B(n16760), .S(n14816), .Z(n14844) );
  OR2_X1 U16857 ( .A1(n14844), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14817) );
  AOI221_X1 U16858 ( .B1(n14818), .B2(n14817), .C1(n14844), .C2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14846) );
  INV_X1 U16859 ( .A(n14819), .ZN(n14828) );
  OAI22_X1 U16860 ( .A1(n18632), .A2(n14822), .B1(n14821), .B2(n14820), .ZN(
        n14824) );
  NAND2_X1 U16861 ( .A1(n14824), .A2(n14823), .ZN(n14827) );
  AOI22_X1 U16862 ( .A1(n15112), .A2(n14825), .B1(n12905), .B2(n14833), .ZN(
        n14826) );
  OAI211_X1 U16863 ( .C1(n14828), .C2(n15112), .A(n14827), .B(n14826), .ZN(
        n18646) );
  INV_X1 U16864 ( .A(n14829), .ZN(n14830) );
  NAND3_X1 U16865 ( .A1(n12905), .A2(n14831), .A3(n14830), .ZN(n14832) );
  NOR2_X1 U16866 ( .A1(n14833), .A2(n14832), .ZN(n18645) );
  OAI21_X1 U16867 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18645), .ZN(n14837) );
  NAND3_X1 U16868 ( .A1(n14834), .A2(n14835), .A3(n16765), .ZN(n14836) );
  NAND2_X1 U16869 ( .A1(n14837), .A2(n14836), .ZN(n14838) );
  OR2_X1 U16870 ( .A1(n14839), .A2(n14838), .ZN(n14840) );
  NOR2_X1 U16871 ( .A1(n18646), .A2(n14840), .ZN(n14842) );
  NAND2_X1 U16872 ( .A1(n15110), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14841) );
  OAI211_X1 U16873 ( .C1(n14844), .C2(n14843), .A(n14842), .B(n14841), .ZN(
        n14845) );
  OR2_X1 U16874 ( .A1(n14846), .A2(n14845), .ZN(n18635) );
  INV_X1 U16875 ( .A(n18635), .ZN(n14847) );
  NAND3_X1 U16876 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n14847), .A3(n14093), 
        .ZN(n14849) );
  AOI22_X1 U16877 ( .A1(n14851), .A2(n14850), .B1(n14849), .B2(n14848), .ZN(
        n18633) );
  OAI21_X1 U16878 ( .B1(n18633), .B2(n18286), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14853) );
  NOR2_X1 U16879 ( .A1(n18286), .A2(n17142), .ZN(n18631) );
  INV_X1 U16880 ( .A(n18631), .ZN(n14852) );
  NAND2_X1 U16881 ( .A1(n14853), .A2(n14852), .ZN(P2_U3593) );
  NAND2_X1 U16882 ( .A1(n14854), .A2(n14855), .ZN(n14949) );
  OR2_X1 U16883 ( .A1(n14854), .A2(n14855), .ZN(n14856) );
  AND2_X1 U16884 ( .A1(n14949), .A2(n14856), .ZN(n21498) );
  INV_X1 U16885 ( .A(n21498), .ZN(n14858) );
  AOI22_X1 U16886 ( .A1(n15264), .A2(n21805), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n15720), .ZN(n14857) );
  OAI21_X1 U16887 ( .B1(n14858), .B2(n15725), .A(n14857), .ZN(P1_U2899) );
  OR2_X1 U16888 ( .A1(n14860), .A2(n14859), .ZN(n14862) );
  NAND2_X1 U16889 ( .A1(n14862), .A2(n14861), .ZN(n14967) );
  NAND2_X1 U16890 ( .A1(n14863), .A2(n17161), .ZN(n14867) );
  INV_X1 U16891 ( .A(n14967), .ZN(n17164) );
  XNOR2_X1 U16892 ( .A(n19255), .B(n17164), .ZN(n14865) );
  NAND2_X1 U16893 ( .A1(n14864), .A2(n17151), .ZN(n14866) );
  NAND3_X1 U16894 ( .A1(n14867), .A2(n14865), .A3(n14866), .ZN(n14954) );
  INV_X1 U16895 ( .A(n14954), .ZN(n14869) );
  AOI21_X1 U16896 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n14868) );
  OAI21_X1 U16897 ( .B1(n14869), .B2(n14868), .A(n19620), .ZN(n14872) );
  INV_X1 U16898 ( .A(n17042), .ZN(n14870) );
  AOI22_X1 U16899 ( .A1(n19397), .A2(n14870), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19613), .ZN(n14871) );
  OAI211_X1 U16900 ( .C1(n14967), .C2(n16201), .A(n14872), .B(n14871), .ZN(
        P2_U2916) );
  OAI21_X1 U16901 ( .B1(n21652), .B2(n21659), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U16902 ( .A1(n14897), .A2(n11698), .ZN(n14873) );
  OAI211_X1 U16903 ( .C1(n21665), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        n14878) );
  OAI22_X1 U16904 ( .A1(n21601), .A2(n14291), .B1(n14876), .B2(n21649), .ZN(
        n14877) );
  AOI211_X1 U16905 ( .C1(n14879), .C2(n21497), .A(n14878), .B(n14877), .ZN(
        n14880) );
  INV_X1 U16906 ( .A(n14880), .ZN(P1_U2840) );
  OR2_X1 U16907 ( .A1(n14881), .A2(n14539), .ZN(n14882) );
  AND2_X1 U16908 ( .A1(n14698), .A2(n14882), .ZN(n18610) );
  INV_X1 U16909 ( .A(n18610), .ZN(n15081) );
  NOR2_X1 U16910 ( .A1(n16176), .A2(n15081), .ZN(n14886) );
  AOI211_X1 U16911 ( .C1(n14884), .C2(n14883), .A(n16178), .B(n14695), .ZN(
        n14885) );
  AOI211_X1 U16912 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n16176), .A(n14886), .B(
        n14885), .ZN(n14887) );
  INV_X1 U16913 ( .A(n14887), .ZN(P2_U2879) );
  NAND2_X1 U16914 ( .A1(n21651), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14892) );
  INV_X1 U16915 ( .A(n14888), .ZN(n14890) );
  AOI22_X1 U16916 ( .A1(n21659), .A2(n14890), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n14889), .ZN(n14891) );
  OAI211_X1 U16917 ( .C1(n21570), .C2(n14893), .A(n14892), .B(n14891), .ZN(
        n14896) );
  AOI21_X1 U16918 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14894) );
  AOI211_X1 U16919 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n14894), .B(n21539), .ZN(n14895) );
  AOI211_X1 U16920 ( .C1(n21341), .C2(n21628), .A(n14896), .B(n14895), .ZN(
        n14899) );
  NAND2_X1 U16921 ( .A1(n14445), .A2(n14897), .ZN(n14898) );
  OAI211_X1 U16922 ( .C1(n14900), .C2(n21471), .A(n14899), .B(n14898), .ZN(
        P1_U2837) );
  OR2_X1 U16923 ( .A1(n14901), .A2(n14700), .ZN(n14902) );
  AND2_X1 U16924 ( .A1(n14902), .A2(n14942), .ZN(n17087) );
  INV_X1 U16925 ( .A(n17087), .ZN(n16682) );
  INV_X1 U16926 ( .A(n14696), .ZN(n14906) );
  INV_X1 U16927 ( .A(n14903), .ZN(n14904) );
  OAI211_X1 U16928 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n16169), .ZN(
        n14908) );
  NAND2_X1 U16929 ( .A1(n16176), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14907) );
  OAI211_X1 U16930 ( .C1(n16682), .C2(n16176), .A(n14908), .B(n14907), .ZN(
        P2_U2877) );
  NAND2_X1 U16931 ( .A1(n14910), .A2(n14911), .ZN(n14912) );
  AND2_X1 U16932 ( .A1(n14909), .A2(n14912), .ZN(n21526) );
  INV_X1 U16933 ( .A(n21526), .ZN(n14913) );
  INV_X1 U16934 ( .A(n15681), .ZN(n21816) );
  OAI222_X1 U16935 ( .A1(n15725), .A2(n14913), .B1(n15260), .B2(n11816), .C1(
        n15259), .C2(n21816), .ZN(P1_U2897) );
  XNOR2_X1 U16936 ( .A(n14914), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14915) );
  XNOR2_X1 U16937 ( .A(n14916), .B(n14915), .ZN(n14933) );
  XNOR2_X1 U16938 ( .A(n14917), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14918) );
  XNOR2_X1 U16939 ( .A(n11005), .B(n14918), .ZN(n14931) );
  OAI22_X1 U16940 ( .A1(n17218), .A2(n18381), .B1(n17125), .B2(n14961), .ZN(
        n14923) );
  OAI22_X1 U16941 ( .A1(n17113), .A2(n14921), .B1(n14920), .B2(n17117), .ZN(
        n14922) );
  AOI211_X1 U16942 ( .C1(n14931), .C2(n17131), .A(n14923), .B(n14922), .ZN(
        n14924) );
  OAI21_X1 U16943 ( .B1(n14933), .B2(n17120), .A(n14924), .ZN(P2_U3011) );
  INV_X1 U16944 ( .A(n14927), .ZN(n14926) );
  NOR2_X1 U16945 ( .A1(n16738), .A2(n14925), .ZN(n16703) );
  OAI21_X1 U16946 ( .B1(n16586), .B2(n14926), .A(n16703), .ZN(n15061) );
  NOR2_X1 U16947 ( .A1(n16723), .A2(n14927), .ZN(n15060) );
  MUX2_X1 U16948 ( .A(n15061), .B(n15060), .S(n15062), .Z(n14930) );
  AOI22_X1 U16949 ( .A1(n18611), .A2(n14803), .B1(n16396), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n14928) );
  OAI21_X1 U16950 ( .B1(n14967), .B2(n16733), .A(n14928), .ZN(n14929) );
  AOI211_X1 U16951 ( .C1(n14931), .C2(n18612), .A(n14930), .B(n14929), .ZN(
        n14932) );
  OAI21_X1 U16952 ( .B1(n14933), .B2(n16730), .A(n14932), .ZN(P2_U3043) );
  OR2_X1 U16953 ( .A1(n14935), .A2(n14934), .ZN(n14938) );
  INV_X1 U16954 ( .A(n14936), .ZN(n14937) );
  NAND2_X1 U16955 ( .A1(n14938), .A2(n14937), .ZN(n18436) );
  OAI222_X1 U16956 ( .A1(n14958), .A2(n14939), .B1(n18436), .B2(n19404), .C1(
        n17214), .C2(n16250), .ZN(P2_U2904) );
  OAI211_X1 U16957 ( .C1(n14903), .C2(n14941), .A(n14940), .B(n16169), .ZN(
        n14947) );
  NAND2_X1 U16958 ( .A1(n14943), .A2(n14942), .ZN(n14945) );
  INV_X1 U16959 ( .A(n15019), .ZN(n14944) );
  NAND2_X1 U16960 ( .A1(n16127), .A2(n18367), .ZN(n14946) );
  OAI211_X1 U16961 ( .C1(n16127), .C2(n13280), .A(n14947), .B(n14946), .ZN(
        P2_U2876) );
  INV_X1 U16962 ( .A(n19897), .ZN(n14948) );
  XNOR2_X1 U16963 ( .A(n19907), .B(n14948), .ZN(n21509) );
  XOR2_X1 U16964 ( .A(n14950), .B(n14949), .Z(n21514) );
  INV_X1 U16965 ( .A(n21514), .ZN(n14959) );
  INV_X1 U16966 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14951) );
  OAI222_X1 U16967 ( .A1(n15657), .A2(n21509), .B1(n15659), .B2(n14959), .C1(
        n14951), .C2(n19911), .ZN(P1_U2866) );
  NAND2_X1 U16968 ( .A1(n19255), .A2(n14967), .ZN(n14953) );
  AOI21_X1 U16969 ( .B1(n14952), .B2(n14861), .A(n11080), .ZN(n18302) );
  AOI21_X1 U16970 ( .B1(n14954), .B2(n14953), .A(n18302), .ZN(n19400) );
  XOR2_X1 U16971 ( .A(n19399), .B(n19400), .Z(n14955) );
  NAND2_X1 U16972 ( .A1(n14955), .A2(n19620), .ZN(n14957) );
  AOI22_X1 U16973 ( .A1(n19619), .A2(n18302), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19613), .ZN(n14956) );
  OAI211_X1 U16974 ( .C1(n19451), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        P2_U2915) );
  INV_X1 U16975 ( .A(n15686), .ZN(n21812) );
  OAI222_X1 U16976 ( .A1(n15259), .A2(n21812), .B1(n15260), .B2(n11794), .C1(
        n15725), .C2(n14959), .ZN(P1_U2898) );
  NOR2_X1 U16977 ( .A1(n18376), .A2(n14960), .ZN(n14962) );
  XNOR2_X1 U16978 ( .A(n14962), .B(n14961), .ZN(n14963) );
  NAND2_X1 U16979 ( .A1(n14963), .A2(n18362), .ZN(n14972) );
  OAI22_X1 U16980 ( .A1(n18522), .A2(n14964), .B1(n18488), .B2(n14920), .ZN(
        n14965) );
  AOI21_X1 U16981 ( .B1(n18576), .B2(P2_REIP_REG_3__SCAN_IN), .A(n14965), .ZN(
        n14966) );
  OAI21_X1 U16982 ( .B1(n18537), .B2(n13271), .A(n14966), .ZN(n14969) );
  NOR2_X1 U16983 ( .A1(n14967), .A2(n18562), .ZN(n14968) );
  AOI211_X1 U16984 ( .C1(n18551), .C2(n14803), .A(n14969), .B(n14968), .ZN(
        n14971) );
  OAI211_X1 U16985 ( .C1(n19255), .C2(n18307), .A(n14972), .B(n14971), .ZN(
        P2_U2852) );
  AOI21_X1 U16986 ( .B1(n14979), .B2(n22269), .A(n21936), .ZN(n14974) );
  AOI21_X1 U16987 ( .B1(n21910), .B2(n14973), .A(n14974), .ZN(n14975) );
  NOR2_X1 U16988 ( .A1(n14975), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14978) );
  NOR2_X1 U16989 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14976), .ZN(
        n14983) );
  INV_X1 U16990 ( .A(n14980), .ZN(n14977) );
  NOR2_X1 U16991 ( .A1(n14977), .A2(n22008), .ZN(n21945) );
  NAND2_X1 U16992 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14986) );
  INV_X1 U16993 ( .A(n21923), .ZN(n21944) );
  NOR2_X1 U16994 ( .A1(n14980), .A2(n22008), .ZN(n21991) );
  INV_X1 U16995 ( .A(n21910), .ZN(n14981) );
  INV_X1 U16996 ( .A(n14973), .ZN(n21962) );
  NOR3_X1 U16997 ( .A1(n14981), .A2(n21962), .A3(n22015), .ZN(n14982) );
  AOI21_X1 U16998 ( .B1(n11391), .B2(n21991), .A(n14982), .ZN(n15007) );
  INV_X1 U16999 ( .A(n14983), .ZN(n15006) );
  OAI22_X1 U17000 ( .A1(n15007), .A2(n22196), .B1(n22192), .B2(n15006), .ZN(
        n14984) );
  AOI21_X1 U17001 ( .B1(n15009), .B2(n22205), .A(n14984), .ZN(n14985) );
  OAI211_X1 U17002 ( .C1(n22269), .C2(n22208), .A(n14986), .B(n14985), .ZN(
        P1_U3070) );
  NAND2_X1 U17003 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14989) );
  OAI22_X1 U17004 ( .A1(n15007), .A2(n22233), .B1(n22229), .B2(n15006), .ZN(
        n14987) );
  AOI21_X1 U17005 ( .B1(n15009), .B2(n22242), .A(n14987), .ZN(n14988) );
  OAI211_X1 U17006 ( .C1(n22269), .C2(n22245), .A(n14989), .B(n14988), .ZN(
        P1_U3071) );
  NAND2_X1 U17007 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14992) );
  OAI22_X1 U17008 ( .A1(n15007), .A2(n22047), .B1(n22043), .B2(n15006), .ZN(
        n14990) );
  AOI21_X1 U17009 ( .B1(n15009), .B2(n22056), .A(n14990), .ZN(n14991) );
  OAI211_X1 U17010 ( .C1(n22269), .C2(n22059), .A(n14992), .B(n14991), .ZN(
        P1_U3066) );
  NAND2_X1 U17011 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14995) );
  OAI22_X1 U17012 ( .A1(n15007), .A2(n21974), .B1(n21966), .B2(n15006), .ZN(
        n14993) );
  AOI21_X1 U17013 ( .B1(n15009), .B2(n22019), .A(n14993), .ZN(n14994) );
  OAI211_X1 U17014 ( .C1(n22269), .C2(n22022), .A(n14995), .B(n14994), .ZN(
        P1_U3065) );
  NAND2_X1 U17015 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14998) );
  OAI22_X1 U17016 ( .A1(n15007), .A2(n22159), .B1(n22155), .B2(n15006), .ZN(
        n14996) );
  AOI21_X1 U17017 ( .B1(n15009), .B2(n22168), .A(n14996), .ZN(n14997) );
  OAI211_X1 U17018 ( .C1(n22269), .C2(n22171), .A(n14998), .B(n14997), .ZN(
        P1_U3069) );
  NAND2_X1 U17019 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15001) );
  OAI22_X1 U17020 ( .A1(n15007), .A2(n22310), .B1(n22304), .B2(n15006), .ZN(
        n14999) );
  AOI21_X1 U17021 ( .B1(n15009), .B2(n22332), .A(n14999), .ZN(n15000) );
  OAI211_X1 U17022 ( .C1(n22269), .C2(n22336), .A(n15001), .B(n15000), .ZN(
        P1_U3072) );
  NAND2_X1 U17023 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n15004) );
  OAI22_X1 U17024 ( .A1(n15007), .A2(n22122), .B1(n22118), .B2(n15006), .ZN(
        n15002) );
  AOI21_X1 U17025 ( .B1(n15009), .B2(n22131), .A(n15002), .ZN(n15003) );
  OAI211_X1 U17026 ( .C1(n22269), .C2(n22134), .A(n15004), .B(n15003), .ZN(
        P1_U3068) );
  NAND2_X1 U17027 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15011) );
  OAI22_X1 U17028 ( .A1(n15007), .A2(n22085), .B1(n22081), .B2(n15006), .ZN(
        n15008) );
  AOI21_X1 U17029 ( .B1(n15009), .B2(n22094), .A(n15008), .ZN(n15010) );
  OAI211_X1 U17030 ( .C1(n22269), .C2(n22097), .A(n15011), .B(n15010), .ZN(
        P1_U3067) );
  OAI21_X1 U17031 ( .B1(n15012), .B2(n15015), .A(n15014), .ZN(n15878) );
  INV_X1 U17032 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15018) );
  OR2_X1 U17033 ( .A1(n15202), .A2(BUF1_REG_9__SCAN_IN), .ZN(n15017) );
  INV_X1 U17034 ( .A(DATAI_9_), .ZN(n16858) );
  NAND2_X1 U17035 ( .A1(n15202), .A2(n16858), .ZN(n15016) );
  NAND2_X1 U17036 ( .A1(n15017), .A2(n15016), .ZN(n21826) );
  OAI222_X1 U17037 ( .A1(n15878), .A2(n15725), .B1(n15018), .B2(n15260), .C1(
        n21826), .C2(n15259), .ZN(P1_U2895) );
  OR2_X1 U17038 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  INV_X1 U17039 ( .A(n18389), .ZN(n15027) );
  INV_X1 U17040 ( .A(n15022), .ZN(n15023) );
  OAI211_X1 U17041 ( .C1(n11354), .C2(n15024), .A(n15023), .B(n16169), .ZN(
        n15026) );
  NAND2_X1 U17042 ( .A1(n16176), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15025) );
  OAI211_X1 U17043 ( .C1(n15027), .C2(n16176), .A(n15026), .B(n15025), .ZN(
        P2_U2875) );
  XNOR2_X1 U17044 ( .A(n19899), .B(n15086), .ZN(n21531) );
  XNOR2_X1 U17045 ( .A(n14909), .B(n15028), .ZN(n21533) );
  INV_X1 U17046 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15029) );
  OAI222_X1 U17047 ( .A1(n15657), .A2(n21531), .B1(n15659), .B2(n21533), .C1(
        n15029), .C2(n19911), .ZN(P1_U2864) );
  OR2_X1 U17048 ( .A1(n15202), .A2(BUF1_REG_8__SCAN_IN), .ZN(n15031) );
  INV_X1 U17049 ( .A(DATAI_8_), .ZN(n16978) );
  NAND2_X1 U17050 ( .A1(n15202), .A2(n16978), .ZN(n15030) );
  NAND2_X1 U17051 ( .A1(n15031), .A2(n15030), .ZN(n21821) );
  INV_X1 U17052 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15032) );
  OAI222_X1 U17053 ( .A1(n15259), .A2(n21821), .B1(n15725), .B2(n21533), .C1(
        n15032), .C2(n15260), .ZN(P1_U2896) );
  NAND2_X1 U17054 ( .A1(n18584), .A2(n15033), .ZN(n15034) );
  XNOR2_X1 U17055 ( .A(n17086), .B(n15034), .ZN(n15046) );
  AOI21_X1 U17056 ( .B1(n15036), .B2(n15035), .A(n11067), .ZN(n15037) );
  INV_X1 U17057 ( .A(n15037), .ZN(n19127) );
  OAI22_X1 U17058 ( .A1(n18562), .A2(n19127), .B1(n18520), .B2(n15038), .ZN(
        n15041) );
  NAND2_X1 U17059 ( .A1(n18551), .A2(n17087), .ZN(n15039) );
  OAI211_X1 U17060 ( .C1(n18488), .C2(n17094), .A(n15039), .B(n14035), .ZN(
        n15040) );
  NOR2_X1 U17061 ( .A1(n15041), .A2(n15040), .ZN(n15043) );
  NAND2_X1 U17062 ( .A1(n18561), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15042) );
  OAI211_X1 U17063 ( .C1(n15044), .C2(n18522), .A(n15043), .B(n15042), .ZN(
        n15045) );
  AOI21_X1 U17064 ( .B1(n15046), .B2(n18362), .A(n15045), .ZN(n15047) );
  INV_X1 U17065 ( .A(n15047), .ZN(P2_U2845) );
  INV_X1 U17066 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18395) );
  OAI211_X1 U17067 ( .C1(n15022), .C2(n15049), .A(n15048), .B(n16169), .ZN(
        n15056) );
  NAND2_X1 U17068 ( .A1(n15051), .A2(n15050), .ZN(n15054) );
  INV_X1 U17069 ( .A(n15052), .ZN(n15053) );
  NAND2_X1 U17070 ( .A1(n15054), .A2(n15053), .ZN(n16424) );
  INV_X1 U17071 ( .A(n16424), .ZN(n18403) );
  NAND2_X1 U17072 ( .A1(n16127), .A2(n18403), .ZN(n15055) );
  OAI211_X1 U17073 ( .C1(n16127), .C2(n18395), .A(n15056), .B(n15055), .ZN(
        P2_U2874) );
  OR2_X1 U17074 ( .A1(n15057), .A2(n15174), .ZN(n15058) );
  NAND2_X1 U17075 ( .A1(n15059), .A2(n15058), .ZN(n17058) );
  INV_X1 U17076 ( .A(n17058), .ZN(n15075) );
  NOR2_X1 U17077 ( .A1(n18306), .A2(n16705), .ZN(n15067) );
  NAND2_X1 U17078 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15060), .ZN(
        n15173) );
  INV_X1 U17079 ( .A(n15061), .ZN(n15064) );
  NAND2_X1 U17080 ( .A1(n16740), .A2(n15062), .ZN(n15063) );
  AND2_X1 U17081 ( .A1(n15064), .A2(n15063), .ZN(n15179) );
  NAND2_X1 U17082 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16396), .ZN(n15065) );
  OAI221_X1 U17083 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15173), .C1(
        n15174), .C2(n15179), .A(n15065), .ZN(n15066) );
  AOI211_X1 U17084 ( .C1(n18302), .C2(n18606), .A(n15067), .B(n15066), .ZN(
        n15074) );
  INV_X1 U17085 ( .A(n15068), .ZN(n15071) );
  INV_X1 U17086 ( .A(n15069), .ZN(n15070) );
  NAND2_X1 U17087 ( .A1(n15071), .A2(n15070), .ZN(n17057) );
  NAND3_X1 U17088 ( .A1(n17057), .A2(n18609), .A3(n15072), .ZN(n15073) );
  OAI211_X1 U17089 ( .C1(n15075), .C2(n18604), .A(n15074), .B(n15073), .ZN(
        P2_U3042) );
  NAND2_X1 U17090 ( .A1(n18584), .A2(n15076), .ZN(n15077) );
  XNOR2_X1 U17091 ( .A(n17070), .B(n15077), .ZN(n15084) );
  AOI22_X1 U17092 ( .A1(n13297), .A2(n15078), .B1(n18561), .B2(
        P2_EBX_REG_8__SCAN_IN), .ZN(n15079) );
  OAI21_X1 U17093 ( .B1(n17079), .B2(n18488), .A(n15079), .ZN(n15083) );
  AOI22_X1 U17094 ( .A1(n18580), .A2(n18605), .B1(n18576), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n15080) );
  OAI211_X1 U17095 ( .C1(n18578), .C2(n15081), .A(n15080), .B(n14035), .ZN(
        n15082) );
  AOI211_X1 U17096 ( .C1(n15084), .C2(n18362), .A(n15083), .B(n15082), .ZN(
        n15085) );
  INV_X1 U17097 ( .A(n15085), .ZN(P2_U2847) );
  INV_X1 U17098 ( .A(n15878), .ZN(n21546) );
  INV_X1 U17099 ( .A(n15659), .ZN(n19908) );
  NAND2_X1 U17100 ( .A1(n19899), .A2(n15086), .ZN(n15089) );
  INV_X1 U17101 ( .A(n15087), .ZN(n15088) );
  NAND2_X1 U17102 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  NAND2_X1 U17103 ( .A1(n15090), .A2(n19893), .ZN(n21543) );
  OAI22_X1 U17104 ( .A1(n21543), .A2(n15657), .B1(n15091), .B2(n19911), .ZN(
        n15092) );
  AOI21_X1 U17105 ( .B1(n21546), .B2(n19908), .A(n15092), .ZN(n15093) );
  INV_X1 U17106 ( .A(n15093), .ZN(P1_U2863) );
  XOR2_X1 U17107 ( .A(n15095), .B(n15122), .Z(n15108) );
  NAND2_X1 U17108 ( .A1(n15096), .A2(n18551), .ZN(n15102) );
  INV_X1 U17109 ( .A(n15097), .ZN(n15098) );
  OAI22_X1 U17110 ( .A1(n18522), .A2(n15098), .B1(n18488), .B2(n14161), .ZN(
        n15100) );
  NOR2_X1 U17111 ( .A1(n18520), .A2(n17217), .ZN(n15099) );
  NOR2_X1 U17112 ( .A1(n15100), .A2(n15099), .ZN(n15101) );
  OAI211_X1 U17113 ( .C1(n18537), .C2(n12475), .A(n15102), .B(n15101), .ZN(
        n15103) );
  INV_X1 U17114 ( .A(n15103), .ZN(n15106) );
  OR2_X1 U17115 ( .A1(n15104), .A2(n18562), .ZN(n15105) );
  OAI211_X1 U17116 ( .C1(n19254), .C2(n18307), .A(n15106), .B(n15105), .ZN(
        n15107) );
  AOI21_X1 U17117 ( .B1(n15108), .B2(n18362), .A(n15107), .ZN(n15109) );
  INV_X1 U17118 ( .A(n15109), .ZN(P2_U2853) );
  OAI22_X1 U17119 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19293), .B1(n15110), 
        .B2(n18644), .ZN(n15111) );
  NAND2_X1 U17120 ( .A1(n14093), .A2(n19293), .ZN(n18621) );
  INV_X1 U17121 ( .A(n18621), .ZN(n15145) );
  INV_X1 U17122 ( .A(n15113), .ZN(n18376) );
  NOR2_X1 U17123 ( .A1(n18376), .A2(n15124), .ZN(n15156) );
  AOI21_X1 U17124 ( .B1(n18376), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15156), .ZN(n15144) );
  AOI222_X1 U17125 ( .A1(n15115), .A2(n15145), .B1(n15114), .B2(n18637), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15144), .ZN(n15117) );
  NAND2_X1 U17126 ( .A1(n16762), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15116) );
  OAI21_X1 U17127 ( .B1(n16762), .B2(n15117), .A(n15116), .ZN(P2_U3601) );
  XOR2_X1 U17128 ( .A(n15118), .B(n15014), .Z(n19940) );
  INV_X1 U17129 ( .A(n19940), .ZN(n21558) );
  INV_X1 U17130 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20008) );
  OR2_X1 U17131 ( .A1(n15202), .A2(n20008), .ZN(n15120) );
  NAND2_X1 U17132 ( .A1(n15202), .A2(DATAI_10_), .ZN(n15119) );
  NAND2_X1 U17133 ( .A1(n15120), .A2(n15119), .ZN(n21831) );
  AOI22_X1 U17134 ( .A1(n15264), .A2(n21831), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15720), .ZN(n15121) );
  OAI21_X1 U17135 ( .B1(n21558), .B2(n15725), .A(n15121), .ZN(P1_U2894) );
  OAI21_X1 U17136 ( .B1(n15124), .B2(n15123), .A(n15122), .ZN(n15142) );
  NOR2_X1 U17137 ( .A1(n18627), .A2(n18584), .ZN(n18431) );
  INV_X1 U17138 ( .A(n18431), .ZN(n18407) );
  OAI22_X1 U17139 ( .A1(n15142), .A2(n18627), .B1(n18407), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15125) );
  INV_X1 U17140 ( .A(n15125), .ZN(n15132) );
  AOI22_X1 U17141 ( .A1(n13297), .A2(n11394), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18577), .ZN(n15127) );
  NAND2_X1 U17142 ( .A1(n18576), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15126) );
  OAI211_X1 U17143 ( .C1(n16732), .C2(n18562), .A(n15127), .B(n15126), .ZN(
        n15130) );
  NOR2_X1 U17144 ( .A1(n15128), .A2(n18578), .ZN(n15129) );
  AOI211_X1 U17145 ( .C1(P2_EBX_REG_1__SCAN_IN), .C2(n18561), .A(n15130), .B(
        n15129), .ZN(n15131) );
  OAI211_X1 U17146 ( .C1(n18307), .C2(n19152), .A(n15132), .B(n15131), .ZN(
        P2_U2854) );
  OR2_X1 U17147 ( .A1(n15134), .A2(n15052), .ZN(n15135) );
  NAND2_X1 U17148 ( .A1(n15133), .A2(n15135), .ZN(n18417) );
  INV_X1 U17149 ( .A(n15048), .ZN(n15139) );
  INV_X1 U17150 ( .A(n15136), .ZN(n15137) );
  OAI211_X1 U17151 ( .C1(n15139), .C2(n15138), .A(n15137), .B(n16169), .ZN(
        n15141) );
  NAND2_X1 U17152 ( .A1(n16176), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15140) );
  OAI211_X1 U17153 ( .C1(n18417), .C2(n16176), .A(n15141), .B(n15140), .ZN(
        P2_U2873) );
  INV_X1 U17154 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15143) );
  OAI21_X1 U17155 ( .B1(n18584), .B2(n15143), .A(n15142), .ZN(n16756) );
  NOR2_X1 U17156 ( .A1(n15144), .A2(n14093), .ZN(n16755) );
  AOI222_X1 U17157 ( .A1(n15146), .A2(n15145), .B1(n16756), .B2(n16755), .C1(
        n17161), .C2(n18637), .ZN(n15148) );
  NAND2_X1 U17158 ( .A1(n16762), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15147) );
  OAI21_X1 U17159 ( .B1(n15148), .B2(n16762), .A(n15147), .ZN(P2_U3599) );
  OAI211_X1 U17160 ( .C1(n15136), .C2(n15151), .A(n15150), .B(n16169), .ZN(
        n15155) );
  AND2_X1 U17161 ( .A1(n15133), .A2(n15152), .ZN(n15153) );
  OR2_X1 U17162 ( .A1(n14079), .A2(n15153), .ZN(n16621) );
  INV_X1 U17163 ( .A(n16621), .ZN(n18433) );
  NAND2_X1 U17164 ( .A1(n18433), .A2(n16127), .ZN(n15154) );
  OAI211_X1 U17165 ( .C1(n16127), .C2(n13283), .A(n15155), .B(n15154), .ZN(
        P2_U2872) );
  NAND2_X1 U17166 ( .A1(n15156), .A2(n18362), .ZN(n15165) );
  OAI21_X1 U17167 ( .B1(n18577), .B2(n18431), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15160) );
  OAI22_X1 U17168 ( .A1(n17170), .A2(n18520), .B1(n18562), .B2(n15157), .ZN(
        n15158) );
  INV_X1 U17169 ( .A(n15158), .ZN(n15159) );
  OAI211_X1 U17170 ( .C1(n18522), .C2(n16749), .A(n15160), .B(n15159), .ZN(
        n15163) );
  NOR2_X1 U17171 ( .A1(n18578), .A2(n15161), .ZN(n15162) );
  AOI211_X1 U17172 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n18561), .A(n15163), .B(
        n15162), .ZN(n15164) );
  OAI211_X1 U17173 ( .C1(n17144), .C2(n18307), .A(n15165), .B(n15164), .ZN(
        P2_U2855) );
  NAND2_X1 U17174 ( .A1(n15167), .A2(n15166), .ZN(n15168) );
  XNOR2_X1 U17175 ( .A(n15169), .B(n15168), .ZN(n15194) );
  OAI21_X1 U17176 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n15187) );
  INV_X1 U17177 ( .A(n15187), .ZN(n15185) );
  AOI221_X1 U17178 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n15178), .C2(n15174), .A(
        n15173), .ZN(n15184) );
  OAI21_X1 U17179 ( .B1(n11080), .B2(n15176), .A(n15175), .ZN(n19403) );
  INV_X1 U17180 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15177) );
  OAI22_X1 U17181 ( .A1(n18323), .A2(n16705), .B1(n18381), .B2(n15177), .ZN(
        n15181) );
  NOR2_X1 U17182 ( .A1(n15179), .A2(n15178), .ZN(n15180) );
  NOR2_X1 U17183 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  OAI21_X1 U17184 ( .B1(n19403), .B2(n16733), .A(n15182), .ZN(n15183) );
  AOI211_X1 U17185 ( .C1(n15185), .C2(n18609), .A(n15184), .B(n15183), .ZN(
        n15186) );
  OAI21_X1 U17186 ( .B1(n18604), .B2(n15194), .A(n15186), .ZN(P2_U3041) );
  NOR2_X1 U17187 ( .A1(n15187), .A2(n17120), .ZN(n15192) );
  NOR2_X1 U17188 ( .A1(n18323), .A2(n17113), .ZN(n15191) );
  OAI22_X1 U17189 ( .A1(n15177), .A2(n18381), .B1(n17125), .B2(n18319), .ZN(
        n15190) );
  INV_X1 U17190 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15188) );
  NOR2_X1 U17191 ( .A1(n17117), .A2(n15188), .ZN(n15189) );
  NOR4_X1 U17192 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15193) );
  OAI21_X1 U17193 ( .B1(n17119), .B2(n15194), .A(n15193), .ZN(P2_U3009) );
  NAND2_X1 U17194 ( .A1(n15196), .A2(n15197), .ZN(n15198) );
  NAND2_X1 U17195 ( .A1(n15195), .A2(n15198), .ZN(n15222) );
  XNOR2_X1 U17196 ( .A(n15222), .B(n15220), .ZN(n21573) );
  INV_X1 U17197 ( .A(n21573), .ZN(n19946) );
  OAI21_X1 U17198 ( .B1(n19893), .B2(n19894), .A(n15199), .ZN(n15200) );
  AND2_X1 U17199 ( .A1(n15200), .A2(n19891), .ZN(n21568) );
  AOI22_X1 U17200 ( .A1(n21568), .A2(n13472), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15650), .ZN(n15201) );
  OAI21_X1 U17201 ( .B1(n19946), .B2(n15659), .A(n15201), .ZN(P1_U2861) );
  INV_X1 U17202 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20010) );
  OR2_X1 U17203 ( .A1(n15202), .A2(n20010), .ZN(n15204) );
  NAND2_X1 U17204 ( .A1(n15202), .A2(DATAI_11_), .ZN(n15203) );
  NAND2_X1 U17205 ( .A1(n15204), .A2(n15203), .ZN(n15660) );
  INV_X1 U17206 ( .A(n15660), .ZN(n21838) );
  OAI222_X1 U17207 ( .A1(n19946), .A2(n15725), .B1(n15205), .B2(n15260), .C1(
        n15259), .C2(n21838), .ZN(P1_U2893) );
  AOI21_X1 U17208 ( .B1(n15207), .B2(n15150), .A(n11006), .ZN(n19621) );
  NAND2_X1 U17209 ( .A1(n19621), .A2(n16169), .ZN(n15209) );
  NAND2_X1 U17210 ( .A1(n16176), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15208) );
  OAI211_X1 U17211 ( .C1(n16602), .C2(n16176), .A(n15209), .B(n15208), .ZN(
        P2_U2871) );
  OAI21_X1 U17212 ( .B1(n11006), .B2(n15212), .A(n15211), .ZN(n16179) );
  INV_X1 U17213 ( .A(n15213), .ZN(n15214) );
  XNOR2_X1 U17214 ( .A(n16080), .B(n15214), .ZN(n18440) );
  NAND2_X1 U17215 ( .A1(n19619), .A2(n18440), .ZN(n15215) );
  OAI21_X1 U17216 ( .B1(n16250), .B2(n15216), .A(n15215), .ZN(n15218) );
  INV_X1 U17217 ( .A(n19616), .ZN(n16252) );
  OAI22_X1 U17218 ( .A1(n16252), .A2(n20021), .B1(n19573), .B2(n16251), .ZN(
        n15217) );
  AOI211_X1 U17219 ( .C1(n19617), .C2(BUF2_REG_17__SCAN_IN), .A(n15218), .B(
        n15217), .ZN(n15219) );
  OAI21_X1 U17220 ( .B1(n16179), .B2(n19398), .A(n15219), .ZN(P2_U2902) );
  INV_X1 U17221 ( .A(n15220), .ZN(n15221) );
  OAI21_X1 U17222 ( .B1(n15222), .B2(n15221), .A(n15195), .ZN(n15224) );
  NAND2_X1 U17223 ( .A1(n15224), .A2(n15223), .ZN(n15263) );
  OAI21_X1 U17224 ( .B1(n15224), .B2(n15223), .A(n15263), .ZN(n19889) );
  INV_X1 U17225 ( .A(n15225), .ZN(n21842) );
  OAI222_X1 U17226 ( .A1(n19889), .A2(n15725), .B1(n15226), .B2(n15260), .C1(
        n15259), .C2(n21842), .ZN(P1_U2892) );
  INV_X1 U17227 ( .A(n15227), .ZN(n15231) );
  INV_X1 U17228 ( .A(n15228), .ZN(n15230) );
  AOI21_X1 U17229 ( .B1(n15231), .B2(n15230), .A(n15229), .ZN(n19966) );
  INV_X1 U17230 ( .A(n19966), .ZN(n15240) );
  XOR2_X1 U17231 ( .A(n15232), .B(n15269), .Z(n21314) );
  AOI22_X1 U17232 ( .A1(n21314), .A2(n13472), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15650), .ZN(n15233) );
  OAI21_X1 U17233 ( .B1(n15240), .B2(n15659), .A(n15233), .ZN(P1_U2858) );
  AOI22_X1 U17234 ( .A1(n15264), .A2(n21855), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15720), .ZN(n15234) );
  OAI21_X1 U17235 ( .B1(n15240), .B2(n15725), .A(n15234), .ZN(P1_U2890) );
  AOI22_X1 U17236 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(n21651), .B1(n21628), 
        .B2(n21314), .ZN(n15235) );
  OAI211_X1 U17237 ( .C1(n21570), .C2(n15236), .A(n15235), .B(n21616), .ZN(
        n15238) );
  INV_X1 U17238 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21310) );
  INV_X1 U17239 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21580) );
  NOR3_X1 U17240 ( .A1(n21576), .A2(n21580), .A3(n21638), .ZN(n15274) );
  NAND2_X1 U17241 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15274), .ZN(n15275) );
  NOR2_X1 U17242 ( .A1(n21310), .A2(n15275), .ZN(n21595) );
  AOI211_X1 U17243 ( .C1(n21310), .C2(n15275), .A(n21595), .B(n21601), .ZN(
        n15237) );
  AOI211_X1 U17244 ( .C1(n19964), .C2(n21659), .A(n15238), .B(n15237), .ZN(
        n15239) );
  OAI21_X1 U17245 ( .B1(n15240), .B2(n21591), .A(n15239), .ZN(P1_U2826) );
  NAND2_X1 U17246 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  NAND2_X1 U17247 ( .A1(n15244), .A2(n15243), .ZN(n21383) );
  NAND2_X1 U17248 ( .A1(n21383), .A2(n19978), .ZN(n15248) );
  NAND2_X1 U17249 ( .A1(n21457), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21379) );
  OAI21_X1 U17250 ( .B1(n15874), .B2(n15245), .A(n21379), .ZN(n15246) );
  AOI21_X1 U17251 ( .B1(n19965), .B2(n21534), .A(n15246), .ZN(n15247) );
  OAI211_X1 U17252 ( .C1(n21533), .C2(n19947), .A(n15248), .B(n15247), .ZN(
        P1_U2991) );
  NOR2_X1 U17253 ( .A1(n15229), .A2(n15250), .ZN(n15251) );
  OR2_X1 U17254 ( .A1(n15253), .A2(n15252), .ZN(n15254) );
  NAND2_X1 U17255 ( .A1(n15286), .A2(n15254), .ZN(n21598) );
  OAI22_X1 U17256 ( .A1(n21598), .A2(n15657), .B1(n15255), .B2(n19911), .ZN(
        n15256) );
  INV_X1 U17257 ( .A(n15256), .ZN(n15257) );
  OAI21_X1 U17258 ( .B1(n21592), .B2(n15659), .A(n15257), .ZN(P1_U2857) );
  OAI222_X1 U17259 ( .A1(n21592), .A2(n15725), .B1(n15260), .B2(n14216), .C1(
        n15259), .C2(n15258), .ZN(P1_U2889) );
  INV_X1 U17260 ( .A(n15261), .ZN(n15262) );
  AOI21_X1 U17261 ( .B1(n15263), .B2(n15262), .A(n15228), .ZN(n15866) );
  INV_X1 U17262 ( .A(n15866), .ZN(n15266) );
  AOI22_X1 U17263 ( .A1(n15264), .A2(n21848), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15720), .ZN(n15265) );
  OAI21_X1 U17264 ( .B1(n15266), .B2(n15725), .A(n15265), .ZN(P1_U2891) );
  INV_X1 U17265 ( .A(n19891), .ZN(n15268) );
  AOI21_X1 U17266 ( .B1(n15268), .B2(n19890), .A(n15267), .ZN(n15270) );
  OR2_X1 U17267 ( .A1(n15270), .A2(n15269), .ZN(n15276) );
  OAI22_X1 U17268 ( .A1(n15276), .A2(n15657), .B1(n15271), .B2(n19911), .ZN(
        n15272) );
  AOI21_X1 U17269 ( .B1(n15866), .B2(n19908), .A(n15272), .ZN(n15273) );
  INV_X1 U17270 ( .A(n15273), .ZN(P1_U2859) );
  AOI21_X1 U17271 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n21594), .A(n15274), 
        .ZN(n15284) );
  INV_X1 U17272 ( .A(n15275), .ZN(n15283) );
  NAND2_X1 U17273 ( .A1(n15866), .A2(n21661), .ZN(n15282) );
  INV_X1 U17274 ( .A(n15864), .ZN(n15280) );
  INV_X1 U17275 ( .A(n15276), .ZN(n21305) );
  AOI22_X1 U17276 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n21651), .B1(n21628), 
        .B2(n21305), .ZN(n15277) );
  OAI211_X1 U17277 ( .C1(n21570), .C2(n15278), .A(n15277), .B(n21616), .ZN(
        n15279) );
  AOI21_X1 U17278 ( .B1(n21659), .B2(n15280), .A(n15279), .ZN(n15281) );
  OAI211_X1 U17279 ( .C1(n15284), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        P1_U2827) );
  NAND2_X1 U17280 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  NAND2_X1 U17281 ( .A1(n15296), .A2(n15287), .ZN(n21614) );
  INV_X1 U17282 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15291) );
  OR2_X1 U17283 ( .A1(n15249), .A2(n15288), .ZN(n15290) );
  AND2_X1 U17284 ( .A1(n15290), .A2(n15289), .ZN(n21612) );
  INV_X1 U17285 ( .A(n21612), .ZN(n15726) );
  OAI222_X1 U17286 ( .A1(n15657), .A2(n21614), .B1(n15291), .B2(n19911), .C1(
        n15726), .C2(n15659), .ZN(P1_U2856) );
  INV_X1 U17287 ( .A(n15289), .ZN(n15295) );
  INV_X1 U17288 ( .A(n15292), .ZN(n15294) );
  OAI21_X1 U17289 ( .B1(n15295), .B2(n15294), .A(n15293), .ZN(n15846) );
  AOI21_X1 U17290 ( .B1(n15297), .B2(n15296), .A(n15654), .ZN(n21436) );
  AOI22_X1 U17291 ( .A1(n21436), .A2(n13472), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15650), .ZN(n15298) );
  OAI21_X1 U17292 ( .B1(n15846), .B2(n15659), .A(n15298), .ZN(P1_U2855) );
  AND2_X1 U17293 ( .A1(n21264), .A2(n17614), .ZN(n20058) );
  NAND2_X1 U17294 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18128) );
  NAND2_X1 U17295 ( .A1(n20058), .A2(n18128), .ZN(n15433) );
  OAI21_X1 U17296 ( .B1(n18721), .B2(n21264), .A(n15433), .ZN(n18175) );
  INV_X1 U17297 ( .A(n18175), .ZN(n15299) );
  NOR2_X1 U17298 ( .A1(n18178), .A2(n15299), .ZN(n15301) );
  NOR3_X1 U17299 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n21703), .ZN(n18173) );
  NOR2_X1 U17300 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21264), .ZN(
        n18676) );
  OR3_X1 U17301 ( .A1(n18173), .A2(n18676), .A3(n18178), .ZN(n15300) );
  MUX2_X1 U17302 ( .A(n15301), .B(n15300), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X4 U17303 ( .A(n11387), .ZN(n17671) );
  AOI22_X1 U17304 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15305) );
  NOR2_X2 U17305 ( .A1(n15308), .A2(n15310), .ZN(n15360) );
  CLKBUF_X3 U17306 ( .A(n17467), .Z(n17643) );
  AOI22_X1 U17307 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15304) );
  NAND3_X1 U17308 ( .A1(n21232), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n20758), .ZN(n20142) );
  AOI22_X1 U17309 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15303) );
  AOI22_X1 U17310 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15302) );
  NAND4_X1 U17311 ( .A1(n15305), .A2(n15304), .A3(n15303), .A4(n15302), .ZN(
        n15316) );
  NOR2_X2 U17312 ( .A1(n20773), .A2(n20117), .ZN(n17663) );
  INV_X4 U17313 ( .A(n17469), .ZN(n17700) );
  INV_X4 U17314 ( .A(n15367), .ZN(n17409) );
  AOI22_X1 U17315 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15314) );
  AOI22_X1 U17316 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15313) );
  AOI22_X1 U17317 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15312) );
  NOR2_X2 U17318 ( .A1(n20774), .A2(n15309), .ZN(n15365) );
  AOI22_X1 U17319 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15311) );
  NAND4_X1 U17320 ( .A1(n15314), .A2(n15313), .A3(n15312), .A4(n15311), .ZN(
        n15315) );
  AOI22_X1 U17321 ( .A1(n10998), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U17322 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U17323 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15318) );
  AOI22_X1 U17324 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15317) );
  NAND4_X1 U17325 ( .A1(n15320), .A2(n15319), .A3(n15318), .A4(n15317), .ZN(
        n15326) );
  AOI22_X1 U17326 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15324) );
  AOI22_X1 U17327 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U17328 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U17329 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15321) );
  NAND4_X1 U17330 ( .A1(n15324), .A2(n15323), .A3(n15322), .A4(n15321), .ZN(
        n15325) );
  AOI22_X1 U17331 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15330) );
  AOI22_X1 U17332 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15329) );
  AOI22_X1 U17333 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U17334 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15327) );
  NAND4_X1 U17335 ( .A1(n15330), .A2(n15329), .A3(n15328), .A4(n15327), .ZN(
        n15336) );
  AOI22_X1 U17336 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15334) );
  AOI22_X1 U17337 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U17338 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U17339 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15331) );
  NAND4_X1 U17340 ( .A1(n15334), .A2(n15333), .A3(n15332), .A4(n15331), .ZN(
        n15335) );
  AOI22_X1 U17341 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U17342 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U17343 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15337) );
  OAI21_X1 U17344 ( .B1(n17369), .B2(n18760), .A(n15337), .ZN(n15343) );
  AOI22_X1 U17345 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U17346 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15340) );
  AOI22_X1 U17347 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U17348 ( .A1(n20777), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15338) );
  NAND4_X1 U17349 ( .A1(n15341), .A2(n15340), .A3(n15339), .A4(n15338), .ZN(
        n15342) );
  NAND3_X2 U17350 ( .A1(n15346), .A2(n15345), .A3(n15344), .ZN(n20649) );
  NAND2_X1 U17351 ( .A1(n19016), .A2(n20649), .ZN(n15389) );
  AOI22_X1 U17352 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U17353 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U17354 ( .A1(n10998), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15347) );
  AOI22_X1 U17355 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U17356 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U17357 ( .A1(n20777), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U17358 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15349) );
  NAND4_X1 U17359 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15353) );
  AOI22_X1 U17360 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15359) );
  INV_X2 U17361 ( .A(n17369), .ZN(n17695) );
  AOI22_X1 U17362 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15358) );
  AOI22_X1 U17363 ( .A1(n20777), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15357) );
  AOI22_X1 U17364 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U17365 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U17366 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15360), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U17367 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15362) );
  AOI22_X1 U17368 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U17369 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15366) );
  OAI21_X1 U17370 ( .B1(n17369), .B2(n19008), .A(n15366), .ZN(n15373) );
  AOI22_X1 U17371 ( .A1(n10998), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15371) );
  AOI22_X1 U17372 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U17373 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U17374 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15368) );
  NAND4_X1 U17375 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(n15368), .ZN(
        n15372) );
  NAND2_X1 U17376 ( .A1(n20796), .A2(n19016), .ZN(n16779) );
  AOI22_X1 U17377 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U17378 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15379) );
  AOI22_X1 U17379 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U17380 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15377) );
  NAND4_X1 U17381 ( .A1(n15380), .A2(n15379), .A3(n15378), .A4(n15377), .ZN(
        n15386) );
  AOI22_X1 U17382 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U17383 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15360), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U17384 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U17385 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15381) );
  NAND4_X1 U17386 ( .A1(n15384), .A2(n15383), .A3(n15382), .A4(n15381), .ZN(
        n15385) );
  NAND2_X1 U17387 ( .A1(n16779), .A2(n20807), .ZN(n15419) );
  NOR2_X1 U17388 ( .A1(n20799), .A2(n20615), .ZN(n15396) );
  INV_X1 U17389 ( .A(n15396), .ZN(n15423) );
  OAI21_X1 U17390 ( .B1(n20113), .B2(n15395), .A(n20746), .ZN(n15427) );
  INV_X1 U17391 ( .A(n20756), .ZN(n15388) );
  NAND3_X1 U17392 ( .A1(n15423), .A2(n15427), .A3(n15388), .ZN(n15393) );
  OAI221_X1 U17393 ( .B1(n20810), .B2(n20649), .C1(n20810), .C2(n20797), .A(
        n15393), .ZN(n15391) );
  NAND2_X1 U17394 ( .A1(n20113), .A2(n20800), .ZN(n16780) );
  AND2_X1 U17395 ( .A1(n20649), .A2(n20746), .ZN(n20554) );
  AOI211_X2 U17396 ( .C1(n20797), .C2(n15419), .A(n15391), .B(n15390), .ZN(
        n20779) );
  NAND2_X1 U17397 ( .A1(n20649), .A2(n15394), .ZN(n17733) );
  OR2_X2 U17398 ( .A1(n20796), .A2(n15397), .ZN(n21257) );
  NAND2_X1 U17399 ( .A1(n17732), .A2(n15395), .ZN(n15420) );
  AND2_X2 U17400 ( .A1(n15420), .A2(n15397), .ZN(n21250) );
  NAND2_X1 U17401 ( .A1(n15396), .A2(n20755), .ZN(n17238) );
  NAND2_X1 U17402 ( .A1(n20800), .A2(n19016), .ZN(n20552) );
  NOR3_X1 U17403 ( .A1(n20585), .A2(n17238), .A3(n20552), .ZN(n20741) );
  NOR3_X1 U17404 ( .A1(n16778), .A2(n20741), .A3(n20061), .ZN(n20743) );
  OAI21_X1 U17405 ( .B1(n20773), .B2(n20759), .A(n15410), .ZN(n15398) );
  NAND2_X1 U17406 ( .A1(n15399), .A2(n15398), .ZN(n21253) );
  NOR2_X1 U17407 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20790) );
  INV_X1 U17408 ( .A(n20790), .ZN(n20767) );
  NOR2_X1 U17409 ( .A1(n21253), .A2(n20767), .ZN(n15431) );
  INV_X2 U17410 ( .A(n21713), .ZN(n21765) );
  NAND2_X1 U17411 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21709), .ZN(n21762) );
  INV_X1 U17412 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21767) );
  NAND2_X1 U17413 ( .A1(n20801), .A2(n16778), .ZN(n16777) );
  AOI22_X1 U17414 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n21234), .B2(n20759), .ZN(
        n15417) );
  NAND2_X1 U17415 ( .A1(n18721), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15414) );
  XNOR2_X1 U17416 ( .A(n15417), .B(n15414), .ZN(n15412) );
  NOR2_X1 U17417 ( .A1(n15417), .A2(n15414), .ZN(n15400) );
  AOI22_X1 U17418 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n21241), .B2(n21240), .ZN(
        n15405) );
  NOR2_X1 U17419 ( .A1(n15406), .A2(n15405), .ZN(n15401) );
  AOI22_X1 U17420 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15410), .B1(
        n15402), .B2(n21232), .ZN(n15407) );
  NOR2_X1 U17421 ( .A1(n15402), .A2(n21232), .ZN(n15408) );
  NAND2_X1 U17422 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15410), .ZN(
        n15403) );
  OAI22_X1 U17423 ( .A1(n15407), .A2(n18683), .B1(n15408), .B2(n15403), .ZN(
        n15404) );
  INV_X1 U17424 ( .A(n15404), .ZN(n15413) );
  XOR2_X1 U17425 ( .A(n15406), .B(n15405), .Z(n17735) );
  NAND2_X1 U17426 ( .A1(n15413), .A2(n17735), .ZN(n15415) );
  OAI21_X1 U17427 ( .B1(n18683), .B2(n15408), .A(n15407), .ZN(n15409) );
  OAI21_X1 U17428 ( .B1(n15410), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15409), .ZN(n15411) );
  INV_X1 U17429 ( .A(n15411), .ZN(n15416) );
  AOI21_X1 U17430 ( .B1(n11033), .B2(n16777), .A(n21249), .ZN(n15429) );
  OAI211_X1 U17431 ( .C1(n18721), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n15414), .B(n15413), .ZN(n17734) );
  OAI211_X1 U17432 ( .C1(n17734), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n20808) );
  AOI211_X1 U17433 ( .C1(n20746), .C2(n17239), .A(n17733), .B(n15419), .ZN(
        n15422) );
  INV_X1 U17434 ( .A(n15420), .ZN(n15421) );
  AOI21_X1 U17435 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(n15424) );
  AOI211_X1 U17436 ( .C1(n15427), .C2(n15426), .A(n15425), .B(n15424), .ZN(
        n15428) );
  INV_X1 U17437 ( .A(n15428), .ZN(n20804) );
  INV_X1 U17438 ( .A(n21256), .ZN(n21238) );
  NOR2_X1 U17439 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21264), .ZN(n18680) );
  MUX2_X1 U17440 ( .A(n15431), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20795), .Z(P3_U3284) );
  AOI21_X1 U17441 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18175), .A(
        n18173), .ZN(n15432) );
  NOR2_X1 U17442 ( .A1(n18178), .A2(n15432), .ZN(n15436) );
  NOR2_X1 U17443 ( .A1(n21234), .A2(n21241), .ZN(n18674) );
  AOI21_X1 U17444 ( .B1(n21264), .B2(n15433), .A(n18674), .ZN(n15434) );
  NOR3_X1 U17445 ( .A1(n18676), .A2(n18178), .A3(n15434), .ZN(n18176) );
  INV_X1 U17446 ( .A(n18176), .ZN(n15435) );
  MUX2_X1 U17447 ( .A(n15436), .B(n15435), .S(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Z(P3_U2865) );
  OAI21_X1 U17448 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n15438), .A(n15437), 
        .ZN(n15441) );
  INV_X1 U17449 ( .A(n15738), .ZN(n15439) );
  AOI22_X1 U17450 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21652), .B1(
        n21659), .B2(n15439), .ZN(n15440) );
  OAI211_X1 U17451 ( .C1(n21649), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        n15443) );
  AOI21_X1 U17452 ( .B1(n21628), .B2(n15906), .A(n15443), .ZN(n15444) );
  OAI21_X1 U17453 ( .B1(n15445), .B2(n21591), .A(n15444), .ZN(P1_U2810) );
  AND2_X1 U17454 ( .A1(n15447), .A2(n15446), .ZN(n15451) );
  OAI21_X1 U17455 ( .B1(n15448), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n15450), 
        .ZN(n15449) );
  OAI21_X1 U17456 ( .B1(n15451), .B2(n15450), .A(n15449), .ZN(P1_U3487) );
  INV_X1 U17457 ( .A(n15452), .ZN(n15455) );
  INV_X1 U17458 ( .A(n15453), .ZN(n15454) );
  INV_X1 U17459 ( .A(n15456), .ZN(n15458) );
  NAND2_X1 U17460 ( .A1(n15504), .A2(n18611), .ZN(n15457) );
  OAI211_X1 U17461 ( .C1(n15460), .C2(n15459), .A(n15458), .B(n15457), .ZN(
        n15461) );
  OAI21_X1 U17462 ( .B1(n15464), .B2(n16730), .A(n15463), .ZN(P2_U3016) );
  NOR2_X1 U17463 ( .A1(n17125), .A2(n15465), .ZN(n15466) );
  AOI211_X1 U17464 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n17126), .A(
        n15467), .B(n15466), .ZN(n15468) );
  OAI21_X1 U17465 ( .B1(n18579), .B2(n17113), .A(n15468), .ZN(n15469) );
  AOI21_X1 U17466 ( .B1(n15470), .B2(n17131), .A(n15469), .ZN(n15471) );
  OAI21_X1 U17467 ( .B1(n15472), .B2(n17120), .A(n15471), .ZN(P2_U2983) );
  AOI22_X1 U17468 ( .A1(n10988), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U17469 ( .A1(n12529), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10980), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U17470 ( .A1(n15477), .A2(n15476), .ZN(n15494) );
  INV_X1 U17471 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U17472 ( .A1(n12531), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15479) );
  AOI21_X1 U17473 ( .B1(n12406), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15482), .ZN(n15478) );
  OAI211_X1 U17474 ( .C1(n15481), .C2(n15480), .A(n15479), .B(n15478), .ZN(
        n15493) );
  INV_X1 U17475 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19343) );
  OAI21_X1 U17476 ( .B1(n15483), .B2(n19343), .A(n15482), .ZN(n15488) );
  INV_X1 U17477 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15486) );
  INV_X1 U17478 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15484) );
  OAI22_X1 U17479 ( .A1(n10986), .A2(n15486), .B1(n15485), .B2(n15484), .ZN(
        n15487) );
  AOI211_X1 U17480 ( .C1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n12533), .A(
        n15488), .B(n15487), .ZN(n15491) );
  AOI22_X1 U17481 ( .A1(n10987), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11001), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U17482 ( .A1(n10981), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10999), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15489) );
  NAND3_X1 U17483 ( .A1(n15491), .A2(n15490), .A3(n15489), .ZN(n15492) );
  OAI21_X1 U17484 ( .B1(n15494), .B2(n15493), .A(n15492), .ZN(n15495) );
  INV_X1 U17485 ( .A(n15495), .ZN(n15496) );
  XNOR2_X1 U17486 ( .A(n15497), .B(n15496), .ZN(n15507) );
  INV_X1 U17487 ( .A(n15498), .ZN(n15499) );
  AOI22_X1 U17488 ( .A1(n19616), .A2(BUF1_REG_30__SCAN_IN), .B1(n15499), .B2(
        n19619), .ZN(n15503) );
  OAI22_X1 U17489 ( .A1(n16251), .A2(n15500), .B1(n16250), .B2(n14403), .ZN(
        n15501) );
  AOI21_X1 U17490 ( .B1(n19617), .B2(BUF2_REG_30__SCAN_IN), .A(n15501), .ZN(
        n15502) );
  OAI211_X1 U17491 ( .C1(n15507), .C2(n19398), .A(n15503), .B(n15502), .ZN(
        P2_U2889) );
  NAND2_X1 U17492 ( .A1(n16176), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15506) );
  NAND2_X1 U17493 ( .A1(n15504), .A2(n16127), .ZN(n15505) );
  OAI211_X1 U17494 ( .C1(n15507), .C2(n16178), .A(n15506), .B(n15505), .ZN(
        P2_U2857) );
  OAI21_X1 U17495 ( .B1(n15519), .B2(n15510), .A(n15509), .ZN(n15617) );
  INV_X1 U17496 ( .A(n15617), .ZN(n15916) );
  AOI22_X1 U17497 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21652), .B1(
        n21659), .B2(n15746), .ZN(n15511) );
  OAI21_X1 U17498 ( .B1(n21649), .B2(n15618), .A(n15511), .ZN(n15514) );
  NAND3_X1 U17499 ( .A1(n15516), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n21594), 
        .ZN(n15512) );
  OAI21_X1 U17500 ( .B1(n15516), .B2(P1_REIP_REG_29__SCAN_IN), .A(n15512), 
        .ZN(n15513) );
  AOI211_X1 U17501 ( .C1(n15916), .C2(n21628), .A(n15514), .B(n15513), .ZN(
        n15515) );
  OAI21_X1 U17502 ( .B1(n15508), .B2(n21591), .A(n15515), .ZN(P1_U2811) );
  INV_X1 U17503 ( .A(n15516), .ZN(n15526) );
  AOI21_X1 U17504 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n21594), .A(n15529), 
        .ZN(n15525) );
  NAND2_X1 U17505 ( .A1(n15767), .A2(n21661), .ZN(n15524) );
  OAI22_X1 U17506 ( .A1(n15517), .A2(n21570), .B1(n21642), .B2(n15765), .ZN(
        n15522) );
  AND2_X1 U17507 ( .A1(n15531), .A2(n15518), .ZN(n15520) );
  OR2_X1 U17508 ( .A1(n15520), .A2(n15519), .ZN(n15922) );
  NOR2_X1 U17509 ( .A1(n15922), .A2(n21665), .ZN(n15521) );
  AOI211_X1 U17510 ( .C1(n21651), .C2(P1_EBX_REG_28__SCAN_IN), .A(n15522), .B(
        n15521), .ZN(n15523) );
  OAI211_X1 U17511 ( .C1(n15526), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        P1_U2812) );
  INV_X1 U17512 ( .A(n15529), .ZN(n15538) );
  OAI21_X1 U17513 ( .B1(n21601), .B2(n19851), .A(n15552), .ZN(n15537) );
  INV_X1 U17514 ( .A(n15546), .ZN(n15533) );
  INV_X1 U17515 ( .A(n15530), .ZN(n15532) );
  OAI21_X1 U17516 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15929) );
  AOI22_X1 U17517 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21652), .B1(
        n21659), .B2(n15774), .ZN(n15535) );
  NAND2_X1 U17518 ( .A1(n21651), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15534) );
  OAI211_X1 U17519 ( .C1(n15929), .C2(n21665), .A(n15535), .B(n15534), .ZN(
        n15536) );
  AOI21_X1 U17520 ( .B1(n15538), .B2(n15537), .A(n15536), .ZN(n15539) );
  OAI21_X1 U17521 ( .B1(n15771), .B2(n21591), .A(n15539), .ZN(P1_U2813) );
  AOI21_X1 U17523 ( .B1(n15542), .B2(n15541), .A(n15527), .ZN(n15784) );
  INV_X1 U17524 ( .A(n15784), .ZN(n15666) );
  INV_X1 U17525 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n19849) );
  INV_X1 U17526 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15543) );
  OAI22_X1 U17527 ( .A1(n15561), .A2(n19849), .B1(n21601), .B2(n15543), .ZN(
        n15551) );
  OR2_X1 U17528 ( .A1(n15557), .A2(n15544), .ZN(n15545) );
  NAND2_X1 U17529 ( .A1(n15546), .A2(n15545), .ZN(n15935) );
  OAI22_X1 U17530 ( .A1(n15547), .A2(n21570), .B1(n21642), .B2(n15782), .ZN(
        n15548) );
  AOI21_X1 U17531 ( .B1(n21651), .B2(P1_EBX_REG_26__SCAN_IN), .A(n15548), .ZN(
        n15549) );
  OAI21_X1 U17532 ( .B1(n15935), .B2(n21665), .A(n15549), .ZN(n15550) );
  AOI21_X1 U17533 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15553) );
  OAI21_X1 U17534 ( .B1(n15666), .B2(n21591), .A(n15553), .ZN(P1_U2814) );
  OAI21_X1 U17535 ( .B1(n15554), .B2(n15555), .A(n15541), .ZN(n15789) );
  AND2_X1 U17536 ( .A1(n15631), .A2(n15556), .ZN(n15558) );
  OR2_X1 U17537 ( .A1(n15558), .A2(n15557), .ZN(n15624) );
  INV_X1 U17538 ( .A(n15624), .ZN(n15950) );
  NOR2_X1 U17539 ( .A1(n21553), .A2(n21561), .ZN(n15587) );
  AND3_X1 U17540 ( .A1(n15560), .A2(P1_REIP_REG_23__SCAN_IN), .A3(n15587), 
        .ZN(n15572) );
  AOI211_X1 U17541 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n15572), .A(n21601), 
        .B(n19849), .ZN(n15566) );
  INV_X1 U17542 ( .A(n15792), .ZN(n15564) );
  OAI22_X1 U17543 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15561), .B1(n15623), 
        .B2(n21649), .ZN(n15562) );
  AOI21_X1 U17544 ( .B1(n21652), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15562), .ZN(n15563) );
  OAI21_X1 U17545 ( .B1(n21642), .B2(n15564), .A(n15563), .ZN(n15565) );
  AOI211_X1 U17546 ( .C1(n15950), .C2(n21628), .A(n15566), .B(n15565), .ZN(
        n15567) );
  OAI21_X1 U17547 ( .B1(n15789), .B2(n21591), .A(n15567), .ZN(P1_U2815) );
  BUF_X1 U17548 ( .A(n15569), .Z(n15570) );
  OAI21_X1 U17549 ( .B1(n15568), .B2(n15571), .A(n15570), .ZN(n15804) );
  NOR2_X1 U17550 ( .A1(n21601), .A2(n15572), .ZN(n21657) );
  NAND2_X1 U17551 ( .A1(n19846), .A2(n15573), .ZN(n15576) );
  INV_X1 U17552 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15574) );
  OAI22_X1 U17553 ( .A1(n15803), .A2(n21570), .B1(n15574), .B2(n21649), .ZN(
        n15575) );
  AOI21_X1 U17554 ( .B1(n21657), .B2(n15576), .A(n15575), .ZN(n15580) );
  NAND2_X1 U17555 ( .A1(n15635), .A2(n15577), .ZN(n15578) );
  AND2_X1 U17556 ( .A1(n15629), .A2(n15578), .ZN(n21460) );
  AOI22_X1 U17557 ( .A1(n21460), .A2(n21628), .B1(n21659), .B2(n15807), .ZN(
        n15579) );
  OAI211_X1 U17558 ( .C1(n15804), .C2(n21591), .A(n15580), .B(n15579), .ZN(
        P1_U2817) );
  AOI21_X1 U17559 ( .B1(n15583), .B2(n15581), .A(n15582), .ZN(n15816) );
  INV_X1 U17560 ( .A(n15816), .ZN(n15693) );
  AND2_X1 U17561 ( .A1(n15646), .A2(n15584), .ZN(n15585) );
  OR2_X1 U17562 ( .A1(n15637), .A2(n15585), .ZN(n15640) );
  INV_X1 U17563 ( .A(n15640), .ZN(n21451) );
  INV_X1 U17564 ( .A(n15586), .ZN(n15814) );
  OAI22_X1 U17565 ( .A1(n15814), .A2(n21642), .B1(n21570), .B2(n12047), .ZN(
        n15589) );
  INV_X1 U17566 ( .A(n15587), .ZN(n21567) );
  OAI21_X1 U17567 ( .B1(n15590), .B2(n21567), .A(n21594), .ZN(n21637) );
  OAI22_X1 U17568 ( .A1(n15639), .A2(n21649), .B1(n19842), .B2(n21637), .ZN(
        n15588) );
  AOI211_X1 U17569 ( .C1(n21628), .C2(n21451), .A(n15589), .B(n15588), .ZN(
        n15591) );
  OR3_X1 U17570 ( .A1(n15590), .A2(n21638), .A3(P1_REIP_REG_21__SCAN_IN), .ZN(
        n21636) );
  OAI211_X1 U17571 ( .C1(n15693), .C2(n21591), .A(n15591), .B(n21636), .ZN(
        P1_U2819) );
  INV_X1 U17572 ( .A(n15592), .ZN(n15597) );
  INV_X1 U17573 ( .A(n15594), .ZN(n15596) );
  AOI21_X1 U17574 ( .B1(n15597), .B2(n15596), .A(n15595), .ZN(n15824) );
  INV_X1 U17575 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21428) );
  INV_X1 U17576 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21600) );
  NAND2_X1 U17577 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21595), .ZN(n21599) );
  NOR2_X1 U17578 ( .A1(n21600), .A2(n21599), .ZN(n21602) );
  NAND2_X1 U17579 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21602), .ZN(n15599) );
  NOR3_X1 U17580 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21428), .A3(n15599), 
        .ZN(n15608) );
  INV_X1 U17581 ( .A(n15599), .ZN(n15598) );
  NOR2_X1 U17582 ( .A1(n21601), .A2(n15598), .ZN(n21620) );
  NOR2_X1 U17583 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15599), .ZN(n21619) );
  OAI21_X1 U17584 ( .B1(n21620), .B2(n21619), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15606) );
  OR2_X1 U17585 ( .A1(n15656), .A2(n15600), .ZN(n15601) );
  AND2_X1 U17586 ( .A1(n15644), .A2(n15601), .ZN(n21444) );
  AOI22_X1 U17587 ( .A1(n15820), .A2(n21659), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n21651), .ZN(n15602) );
  OAI211_X1 U17588 ( .C1(n21570), .C2(n15603), .A(n15602), .B(n21616), .ZN(
        n15604) );
  AOI21_X1 U17589 ( .B1(n21628), .B2(n21444), .A(n15604), .ZN(n15605) );
  NAND2_X1 U17590 ( .A1(n15606), .A2(n15605), .ZN(n15607) );
  AOI211_X1 U17591 ( .C1(n15824), .C2(n21661), .A(n15608), .B(n15607), .ZN(
        n15609) );
  INV_X1 U17592 ( .A(n15609), .ZN(P1_U2821) );
  OAI21_X1 U17593 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21602), .A(n21620), 
        .ZN(n15610) );
  INV_X1 U17594 ( .A(n15610), .ZN(n15614) );
  AOI22_X1 U17595 ( .A1(n15843), .A2(n21659), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n21651), .ZN(n15611) );
  OAI211_X1 U17596 ( .C1(n21570), .C2(n15612), .A(n15611), .B(n21616), .ZN(
        n15613) );
  AOI211_X1 U17597 ( .C1(n21436), .C2(n21628), .A(n15614), .B(n15613), .ZN(
        n15615) );
  OAI21_X1 U17598 ( .B1(n15846), .B2(n21591), .A(n15615), .ZN(P1_U2823) );
  OAI22_X1 U17599 ( .A1(n15879), .A2(n15657), .B1(n19911), .B2(n15616), .ZN(
        P1_U2841) );
  OAI222_X1 U17600 ( .A1(n15659), .A2(n15508), .B1(n15618), .B2(n19911), .C1(
        n15617), .C2(n15657), .ZN(P1_U2843) );
  INV_X1 U17601 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15619) );
  OAI222_X1 U17602 ( .A1(n15659), .A2(n15620), .B1(n15619), .B2(n19911), .C1(
        n15922), .C2(n15657), .ZN(P1_U2844) );
  INV_X1 U17603 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15622) );
  OAI222_X1 U17604 ( .A1(n15659), .A2(n15666), .B1(n15622), .B2(n19911), .C1(
        n15935), .C2(n15657), .ZN(P1_U2846) );
  OAI22_X1 U17605 ( .A1(n15624), .A2(n15657), .B1(n15623), .B2(n19911), .ZN(
        n15625) );
  INV_X1 U17606 ( .A(n15625), .ZN(n15626) );
  OAI21_X1 U17607 ( .B1(n15789), .B2(n15659), .A(n15626), .ZN(P1_U2847) );
  AOI21_X1 U17608 ( .B1(n15627), .B2(n15570), .A(n15554), .ZN(n21662) );
  INV_X1 U17609 ( .A(n21662), .ZN(n15677) );
  INV_X1 U17610 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15632) );
  NAND2_X1 U17611 ( .A1(n15629), .A2(n15628), .ZN(n15630) );
  NAND2_X1 U17612 ( .A1(n15631), .A2(n15630), .ZN(n21666) );
  OAI222_X1 U17613 ( .A1(n15659), .A2(n15677), .B1(n15632), .B2(n19911), .C1(
        n21666), .C2(n15657), .ZN(P1_U2848) );
  AOI22_X1 U17614 ( .A1(n21460), .A2(n13472), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15650), .ZN(n15633) );
  OAI21_X1 U17615 ( .B1(n15804), .B2(n15659), .A(n15633), .ZN(P1_U2849) );
  AOI21_X1 U17616 ( .B1(n15634), .B2(n11376), .A(n15568), .ZN(n21646) );
  INV_X1 U17617 ( .A(n21646), .ZN(n15688) );
  OAI21_X1 U17618 ( .B1(n15637), .B2(n15636), .A(n15635), .ZN(n21644) );
  INV_X1 U17619 ( .A(n21644), .ZN(n15980) );
  AOI22_X1 U17620 ( .A1(n15980), .A2(n13472), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15650), .ZN(n15638) );
  OAI21_X1 U17621 ( .B1(n15688), .B2(n15659), .A(n15638), .ZN(P1_U2850) );
  OAI22_X1 U17622 ( .A1(n15640), .A2(n15657), .B1(n15639), .B2(n19911), .ZN(
        n15641) );
  INV_X1 U17623 ( .A(n15641), .ZN(n15642) );
  OAI21_X1 U17624 ( .B1(n15693), .B2(n15659), .A(n15642), .ZN(P1_U2851) );
  NAND2_X1 U17625 ( .A1(n15644), .A2(n15643), .ZN(n15645) );
  NAND2_X1 U17626 ( .A1(n15646), .A2(n15645), .ZN(n21627) );
  INV_X1 U17627 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15649) );
  OR2_X1 U17628 ( .A1(n15595), .A2(n15647), .ZN(n15648) );
  AND2_X1 U17629 ( .A1(n15581), .A2(n15648), .ZN(n21631) );
  INV_X1 U17630 ( .A(n21631), .ZN(n15699) );
  OAI222_X1 U17631 ( .A1(n15657), .A2(n21627), .B1(n15649), .B2(n19911), .C1(
        n15699), .C2(n15659), .ZN(P1_U2852) );
  INV_X1 U17632 ( .A(n15824), .ZN(n15705) );
  AOI22_X1 U17633 ( .A1(n21444), .A2(n13472), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15650), .ZN(n15651) );
  OAI21_X1 U17634 ( .B1(n15705), .B2(n15659), .A(n15651), .ZN(P1_U2853) );
  AOI21_X1 U17635 ( .B1(n15652), .B2(n15293), .A(n15594), .ZN(n21621) );
  INV_X1 U17636 ( .A(n21621), .ZN(n15711) );
  INV_X1 U17637 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15658) );
  NOR2_X1 U17638 ( .A1(n15654), .A2(n15653), .ZN(n15655) );
  OR2_X1 U17639 ( .A1(n15656), .A2(n15655), .ZN(n21624) );
  OAI222_X1 U17640 ( .A1(n15711), .A2(n15659), .B1(n15658), .B2(n19911), .C1(
        n15657), .C2(n21624), .ZN(P1_U2854) );
  AOI22_X1 U17641 ( .A1(n15722), .A2(n15660), .B1(n15720), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n15661) );
  OAI21_X1 U17642 ( .B1(n15724), .B2(n14582), .A(n15661), .ZN(n15663) );
  NOR2_X1 U17643 ( .A1(n15771), .A2(n15725), .ZN(n15662) );
  AOI211_X1 U17644 ( .C1(n15729), .C2(BUF1_REG_27__SCAN_IN), .A(n15663), .B(
        n15662), .ZN(n15664) );
  INV_X1 U17645 ( .A(n15664), .ZN(P1_U2877) );
  AOI22_X1 U17646 ( .A1(n15722), .A2(n21831), .B1(n15720), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n15665) );
  OAI21_X1 U17647 ( .B1(n15724), .B2(n14589), .A(n15665), .ZN(n15668) );
  NOR2_X1 U17648 ( .A1(n15666), .A2(n15725), .ZN(n15667) );
  AOI211_X1 U17649 ( .C1(BUF1_REG_26__SCAN_IN), .C2(n15729), .A(n15668), .B(
        n15667), .ZN(n15669) );
  INV_X1 U17650 ( .A(n15669), .ZN(P1_U2878) );
  INV_X1 U17651 ( .A(n21826), .ZN(n15670) );
  AOI22_X1 U17652 ( .A1(n15722), .A2(n15670), .B1(n15720), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n15671) );
  OAI21_X1 U17653 ( .B1(n15724), .B2(n16868), .A(n15671), .ZN(n15673) );
  NOR2_X1 U17654 ( .A1(n15789), .A2(n15725), .ZN(n15672) );
  AOI211_X1 U17655 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n15729), .A(n15673), .B(
        n15672), .ZN(n15674) );
  INV_X1 U17656 ( .A(n15674), .ZN(P1_U2879) );
  INV_X1 U17657 ( .A(n21821), .ZN(n15675) );
  AOI22_X1 U17658 ( .A1(n15722), .A2(n15675), .B1(n15720), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n15676) );
  OAI21_X1 U17659 ( .B1(n16946), .B2(n15724), .A(n15676), .ZN(n15679) );
  NOR2_X1 U17660 ( .A1(n15677), .A2(n15725), .ZN(n15678) );
  AOI211_X1 U17661 ( .C1(n15729), .C2(BUF1_REG_24__SCAN_IN), .A(n15679), .B(
        n15678), .ZN(n15680) );
  INV_X1 U17662 ( .A(n15680), .ZN(P1_U2880) );
  AOI22_X1 U17663 ( .A1(n15722), .A2(n15681), .B1(n15720), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n15682) );
  OAI21_X1 U17664 ( .B1(n15724), .B2(n16960), .A(n15682), .ZN(n15684) );
  NOR2_X1 U17665 ( .A1(n15804), .A2(n15725), .ZN(n15683) );
  AOI211_X1 U17666 ( .C1(n15729), .C2(BUF1_REG_23__SCAN_IN), .A(n15684), .B(
        n15683), .ZN(n15685) );
  INV_X1 U17667 ( .A(n15685), .ZN(P1_U2881) );
  AOI22_X1 U17668 ( .A1(n15722), .A2(n15686), .B1(n15720), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n15687) );
  OAI21_X1 U17669 ( .B1(n15724), .B2(n16961), .A(n15687), .ZN(n15690) );
  NOR2_X1 U17670 ( .A1(n15688), .A2(n15725), .ZN(n15689) );
  AOI211_X1 U17671 ( .C1(n15729), .C2(BUF1_REG_22__SCAN_IN), .A(n15690), .B(
        n15689), .ZN(n15691) );
  INV_X1 U17672 ( .A(n15691), .ZN(P1_U2882) );
  AOI22_X1 U17673 ( .A1(n15722), .A2(n21805), .B1(n15720), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U17674 ( .B1(n15724), .B2(n14552), .A(n15692), .ZN(n15695) );
  NOR2_X1 U17675 ( .A1(n15693), .A2(n15725), .ZN(n15694) );
  AOI211_X1 U17676 ( .C1(n15729), .C2(BUF1_REG_21__SCAN_IN), .A(n15695), .B(
        n15694), .ZN(n15696) );
  INV_X1 U17677 ( .A(n15696), .ZN(P1_U2883) );
  AOI22_X1 U17678 ( .A1(n15722), .A2(n15697), .B1(n15720), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n15698) );
  OAI21_X1 U17679 ( .B1(n16880), .B2(n15724), .A(n15698), .ZN(n15701) );
  NOR2_X1 U17680 ( .A1(n15699), .A2(n15725), .ZN(n15700) );
  AOI211_X1 U17681 ( .C1(n15729), .C2(BUF1_REG_20__SCAN_IN), .A(n15701), .B(
        n15700), .ZN(n15702) );
  INV_X1 U17682 ( .A(n15702), .ZN(P1_U2884) );
  AOI22_X1 U17683 ( .A1(n15722), .A2(n15703), .B1(n15720), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n15704) );
  OAI21_X1 U17684 ( .B1(n15724), .B2(n16944), .A(n15704), .ZN(n15707) );
  NOR2_X1 U17685 ( .A1(n15705), .A2(n15725), .ZN(n15706) );
  AOI211_X1 U17686 ( .C1(n15729), .C2(BUF1_REG_19__SCAN_IN), .A(n15707), .B(
        n15706), .ZN(n15708) );
  INV_X1 U17687 ( .A(n15708), .ZN(P1_U2885) );
  AOI22_X1 U17688 ( .A1(n15722), .A2(n15709), .B1(n15720), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n15710) );
  OAI21_X1 U17689 ( .B1(n16963), .B2(n15724), .A(n15710), .ZN(n15713) );
  NOR2_X1 U17690 ( .A1(n15711), .A2(n15725), .ZN(n15712) );
  AOI211_X1 U17691 ( .C1(n15729), .C2(BUF1_REG_18__SCAN_IN), .A(n15713), .B(
        n15712), .ZN(n15714) );
  INV_X1 U17692 ( .A(n15714), .ZN(P1_U2886) );
  AOI22_X1 U17693 ( .A1(n15722), .A2(n15715), .B1(n15720), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n15716) );
  OAI21_X1 U17694 ( .B1(n15724), .B2(n16964), .A(n15716), .ZN(n15718) );
  NOR2_X1 U17695 ( .A1(n15846), .A2(n15725), .ZN(n15717) );
  AOI211_X1 U17696 ( .C1(n15729), .C2(BUF1_REG_17__SCAN_IN), .A(n15718), .B(
        n15717), .ZN(n15719) );
  INV_X1 U17697 ( .A(n15719), .ZN(P1_U2887) );
  AOI22_X1 U17698 ( .A1(n15722), .A2(n15721), .B1(n15720), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n15723) );
  OAI21_X1 U17699 ( .B1(n16943), .B2(n15724), .A(n15723), .ZN(n15728) );
  NOR2_X1 U17700 ( .A1(n15726), .A2(n15725), .ZN(n15727) );
  AOI211_X1 U17701 ( .C1(n15729), .C2(BUF1_REG_16__SCAN_IN), .A(n15728), .B(
        n15727), .ZN(n15730) );
  INV_X1 U17702 ( .A(n15730), .ZN(P1_U2888) );
  OR2_X2 U17703 ( .A1(n15731), .A2(n11399), .ZN(n15735) );
  NAND3_X1 U17704 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15900) );
  NAND2_X1 U17705 ( .A1(n15731), .A2(n15900), .ZN(n15734) );
  INV_X1 U17706 ( .A(n15743), .ZN(n15733) );
  AND3_X2 U17707 ( .A1(n15735), .A2(n15734), .A3(n15733), .ZN(n15736) );
  NAND2_X1 U17708 ( .A1(n21457), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15902) );
  NAND2_X1 U17709 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15737) );
  OAI211_X1 U17710 ( .C1(n19982), .C2(n15738), .A(n15902), .B(n15737), .ZN(
        n15739) );
  AOI21_X1 U17711 ( .B1(n15740), .B2(n19979), .A(n15739), .ZN(n15741) );
  OAI21_X1 U17712 ( .B1(n15908), .B2(n21667), .A(n15741), .ZN(P1_U2969) );
  NOR2_X1 U17713 ( .A1(n15743), .A2(n15742), .ZN(n15745) );
  XOR2_X1 U17714 ( .A(n15745), .B(n15744), .Z(n15918) );
  NAND2_X1 U17715 ( .A1(n15746), .A2(n19965), .ZN(n15750) );
  NAND2_X1 U17716 ( .A1(n21457), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15912) );
  OAI21_X1 U17717 ( .B1(n15874), .B2(n15747), .A(n15912), .ZN(n15748) );
  INV_X1 U17718 ( .A(n15748), .ZN(n15749) );
  OAI21_X1 U17719 ( .B1(n21667), .B2(n15918), .A(n15753), .ZN(P1_U2970) );
  NAND2_X1 U17720 ( .A1(n15754), .A2(n15777), .ZN(n15761) );
  OAI21_X1 U17721 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15755), .A(
        n15761), .ZN(n15756) );
  INV_X1 U17722 ( .A(n15756), .ZN(n15760) );
  NAND2_X1 U17723 ( .A1(n19950), .A2(n15779), .ZN(n15758) );
  NAND2_X1 U17724 ( .A1(n15762), .A2(n11400), .ZN(n15763) );
  XOR2_X1 U17725 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15763), .Z(
        n15926) );
  INV_X1 U17726 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n19854) );
  NOR2_X1 U17727 ( .A1(n21616), .A2(n19854), .ZN(n15921) );
  AOI21_X1 U17728 ( .B1(n19976), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15921), .ZN(n15764) );
  OAI21_X1 U17729 ( .B1(n19982), .B2(n15765), .A(n15764), .ZN(n15766) );
  AOI21_X1 U17730 ( .B1(n15767), .B2(n19979), .A(n15766), .ZN(n15768) );
  OAI21_X1 U17731 ( .B1(n21667), .B2(n15926), .A(n15768), .ZN(P1_U2971) );
  XNOR2_X1 U17732 ( .A(n19950), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15769) );
  XNOR2_X1 U17733 ( .A(n15731), .B(n15769), .ZN(n15934) );
  INV_X1 U17734 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15770) );
  NAND2_X1 U17735 ( .A1(n21457), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15927) );
  OAI21_X1 U17736 ( .B1(n15874), .B2(n15770), .A(n15927), .ZN(n15773) );
  NOR2_X1 U17737 ( .A1(n15771), .A2(n19947), .ZN(n15772) );
  OAI21_X1 U17738 ( .B1(n15934), .B2(n21667), .A(n15775), .ZN(P1_U2972) );
  NAND3_X1 U17739 ( .A1(n15778), .A2(n15776), .A3(n15777), .ZN(n15780) );
  XNOR2_X1 U17740 ( .A(n15780), .B(n15779), .ZN(n15943) );
  NAND2_X1 U17741 ( .A1(n21457), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U17742 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15781) );
  OAI211_X1 U17743 ( .C1(n19982), .C2(n15782), .A(n15937), .B(n15781), .ZN(
        n15783) );
  AOI21_X1 U17744 ( .B1(n15784), .B2(n19979), .A(n15783), .ZN(n15785) );
  OAI21_X1 U17745 ( .B1(n21667), .B2(n15943), .A(n15785), .ZN(P1_U2973) );
  NOR2_X1 U17746 ( .A1(n15754), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15786) );
  NAND2_X1 U17747 ( .A1(n10972), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15800) );
  OAI211_X1 U17748 ( .C1(n15786), .C2(n15944), .A(n15776), .B(n15800), .ZN(
        n15787) );
  XNOR2_X1 U17749 ( .A(n15787), .B(n15947), .ZN(n15952) );
  NAND2_X1 U17750 ( .A1(n21457), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15946) );
  OAI21_X1 U17751 ( .B1(n15874), .B2(n15788), .A(n15946), .ZN(n15791) );
  NOR2_X1 U17752 ( .A1(n15789), .A2(n19947), .ZN(n15790) );
  AOI211_X1 U17753 ( .C1(n19965), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15793) );
  OAI21_X1 U17754 ( .B1(n21667), .B2(n15952), .A(n15793), .ZN(P1_U2974) );
  NAND2_X1 U17755 ( .A1(n15754), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15795) );
  INV_X1 U17756 ( .A(n15754), .ZN(n15802) );
  NAND2_X1 U17757 ( .A1(n15802), .A2(n15953), .ZN(n15794) );
  MUX2_X1 U17758 ( .A(n15795), .B(n15794), .S(n10972), .Z(n15796) );
  XNOR2_X1 U17759 ( .A(n15796), .B(n15959), .ZN(n15964) );
  INV_X1 U17760 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21655) );
  NOR2_X1 U17761 ( .A1(n21616), .A2(n21655), .ZN(n15955) );
  AOI21_X1 U17762 ( .B1(n19976), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15955), .ZN(n15797) );
  OAI21_X1 U17763 ( .B1(n19982), .B2(n21658), .A(n15797), .ZN(n15798) );
  AOI21_X1 U17764 ( .B1(n21662), .B2(n19979), .A(n15798), .ZN(n15799) );
  OAI21_X1 U17765 ( .B1(n21667), .B2(n15964), .A(n15799), .ZN(P1_U2975) );
  OAI21_X1 U17766 ( .B1(n10972), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15800), .ZN(n15801) );
  XNOR2_X1 U17767 ( .A(n15802), .B(n15801), .ZN(n21459) );
  OAI22_X1 U17768 ( .A1(n15874), .A2(n15803), .B1(n21616), .B2(n19846), .ZN(
        n15806) );
  NOR2_X1 U17769 ( .A1(n15804), .A2(n19947), .ZN(n15805) );
  AOI211_X1 U17770 ( .C1(n19965), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15808) );
  OAI21_X1 U17771 ( .B1(n21459), .B2(n21667), .A(n15808), .ZN(P1_U2976) );
  MUX2_X1 U17772 ( .A(n15810), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .S(
        n19950), .Z(n15827) );
  NAND2_X1 U17773 ( .A1(n15809), .A2(n15827), .ZN(n15826) );
  OAI21_X1 U17774 ( .B1(n15810), .B2(n19950), .A(n15826), .ZN(n15819) );
  AOI22_X1 U17775 ( .A1(n15819), .A2(n15985), .B1(n19950), .B2(n15826), .ZN(
        n15984) );
  NOR2_X1 U17776 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15985), .ZN(
        n15989) );
  INV_X1 U17777 ( .A(n15989), .ZN(n15811) );
  OAI211_X1 U17778 ( .C1(n13565), .C2(n19950), .A(n15984), .B(n15811), .ZN(
        n15812) );
  XNOR2_X1 U17779 ( .A(n15812), .B(n21456), .ZN(n21450) );
  AOI22_X1 U17780 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n21457), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15813) );
  OAI21_X1 U17781 ( .B1(n19982), .B2(n15814), .A(n15813), .ZN(n15815) );
  AOI21_X1 U17782 ( .B1(n15816), .B2(n19979), .A(n15815), .ZN(n15817) );
  OAI21_X1 U17783 ( .B1(n21450), .B2(n21667), .A(n15817), .ZN(P1_U2978) );
  MUX2_X1 U17784 ( .A(n15985), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n19950), .Z(n15818) );
  XNOR2_X1 U17785 ( .A(n15819), .B(n15818), .ZN(n21443) );
  INV_X1 U17786 ( .A(n15820), .ZN(n15822) );
  AOI22_X1 U17787 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n21457), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15821) );
  OAI21_X1 U17788 ( .B1(n19982), .B2(n15822), .A(n15821), .ZN(n15823) );
  AOI21_X1 U17789 ( .B1(n15824), .B2(n19979), .A(n15823), .ZN(n15825) );
  OAI21_X1 U17790 ( .B1(n21443), .B2(n21667), .A(n15825), .ZN(P1_U2980) );
  OAI21_X1 U17791 ( .B1(n15809), .B2(n15827), .A(n15826), .ZN(n21431) );
  AOI22_X1 U17792 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n21457), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15828) );
  OAI21_X1 U17793 ( .B1(n21617), .B2(n19982), .A(n15828), .ZN(n15829) );
  AOI21_X1 U17794 ( .B1(n21621), .B2(n19979), .A(n15829), .ZN(n15830) );
  OAI21_X1 U17795 ( .B1(n21667), .B2(n21431), .A(n15830), .ZN(P1_U2981) );
  NAND2_X1 U17796 ( .A1(n11346), .A2(n15832), .ZN(n19959) );
  OAI21_X1 U17797 ( .B1(n19950), .B2(n16005), .A(n15833), .ZN(n15834) );
  AOI21_X1 U17798 ( .B1(n19959), .B2(n15835), .A(n15834), .ZN(n15836) );
  INV_X1 U17799 ( .A(n15836), .ZN(n15839) );
  AOI21_X1 U17800 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19950), .A(
        n15836), .ZN(n15837) );
  AOI21_X1 U17801 ( .B1(n13550), .B2(n16000), .A(n15837), .ZN(n15838) );
  OAI21_X1 U17802 ( .B1(n16000), .B2(n15839), .A(n15838), .ZN(n15840) );
  XNOR2_X1 U17803 ( .A(n15840), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21437) );
  NAND2_X1 U17804 ( .A1(n21437), .A2(n19978), .ZN(n15845) );
  INV_X1 U17805 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15841) );
  OAI22_X1 U17806 ( .A1(n15874), .A2(n15612), .B1(n21616), .B2(n15841), .ZN(
        n15842) );
  AOI21_X1 U17807 ( .B1(n19965), .B2(n15843), .A(n15842), .ZN(n15844) );
  OAI211_X1 U17808 ( .C1(n19947), .C2(n15846), .A(n15845), .B(n15844), .ZN(
        P1_U2982) );
  MUX2_X1 U17809 ( .A(n16005), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n19950), .Z(n15849) );
  NAND2_X1 U17810 ( .A1(n19950), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15998) );
  MUX2_X1 U17811 ( .A(n15849), .B(n15998), .S(n15999), .Z(n15850) );
  NAND3_X1 U17812 ( .A1(n15999), .A2(n10972), .A3(n16005), .ZN(n15997) );
  NAND2_X1 U17813 ( .A1(n15850), .A2(n15997), .ZN(n16016) );
  NAND2_X1 U17814 ( .A1(n16016), .A2(n19978), .ZN(n15855) );
  INV_X1 U17815 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15851) );
  NOR2_X1 U17816 ( .A1(n21616), .A2(n15851), .ZN(n16018) );
  INV_X1 U17817 ( .A(n21588), .ZN(n15852) );
  NOR2_X1 U17818 ( .A1(n19982), .A2(n15852), .ZN(n15853) );
  AOI211_X1 U17819 ( .C1(n19976), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16018), .B(n15853), .ZN(n15854) );
  OAI211_X1 U17820 ( .C1(n19947), .C2(n21592), .A(n15855), .B(n15854), .ZN(
        P1_U2984) );
  NAND2_X1 U17821 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15856) );
  NAND2_X1 U17822 ( .A1(n19950), .A2(n15856), .ZN(n19957) );
  INV_X1 U17823 ( .A(n15857), .ZN(n15858) );
  INV_X1 U17824 ( .A(n15860), .ZN(n19949) );
  AND3_X1 U17825 ( .A1(n19948), .A2(n19949), .A3(n15859), .ZN(n19951) );
  NOR2_X1 U17826 ( .A1(n19951), .A2(n15860), .ZN(n15862) );
  XNOR2_X1 U17827 ( .A(n15862), .B(n15861), .ZN(n21306) );
  INV_X1 U17828 ( .A(n21306), .ZN(n15868) );
  AOI22_X1 U17829 ( .A1(n19976), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21457), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15863) );
  OAI21_X1 U17830 ( .B1(n19982), .B2(n15864), .A(n15863), .ZN(n15865) );
  AOI21_X1 U17831 ( .B1(n15866), .B2(n19979), .A(n15865), .ZN(n15867) );
  OAI21_X1 U17832 ( .B1(n15868), .B2(n21667), .A(n15867), .ZN(P1_U2986) );
  OAI21_X1 U17833 ( .B1(n15872), .B2(n15871), .A(n15870), .ZN(n21392) );
  NAND2_X1 U17834 ( .A1(n21392), .A2(n19978), .ZN(n15877) );
  INV_X1 U17835 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15873) );
  NAND2_X1 U17836 ( .A1(n21457), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n21388) );
  OAI21_X1 U17837 ( .B1(n15874), .B2(n15873), .A(n21388), .ZN(n15875) );
  AOI21_X1 U17838 ( .B1(n21549), .B2(n19965), .A(n15875), .ZN(n15876) );
  OAI211_X1 U17839 ( .C1(n19947), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        P1_U2990) );
  NOR2_X1 U17840 ( .A1(n15879), .A2(n21429), .ZN(n15896) );
  NOR2_X1 U17841 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21297), .ZN(
        n15880) );
  NOR2_X1 U17842 ( .A1(n13418), .A2(n15977), .ZN(n15883) );
  AND4_X1 U17843 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n21427), .ZN(n15973) );
  INV_X1 U17844 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21378) );
  INV_X1 U17845 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21357) );
  NOR3_X1 U17846 ( .A1(n21378), .A2(n21377), .A3(n21357), .ZN(n21397) );
  NAND3_X1 U17847 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n21397), .ZN(n16002) );
  NAND2_X1 U17848 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21337) );
  NOR3_X1 U17849 ( .A1(n21336), .A2(n15882), .A3(n21337), .ZN(n21366) );
  NAND2_X1 U17850 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21366), .ZN(
        n16003) );
  OR2_X1 U17851 ( .A1(n16002), .A2(n16003), .ZN(n16006) );
  NOR3_X1 U17852 ( .A1(n13559), .A2(n21417), .A3(n16006), .ZN(n21304) );
  NAND2_X1 U17853 ( .A1(n15973), .A2(n21304), .ZN(n15974) );
  INV_X1 U17854 ( .A(n15974), .ZN(n15968) );
  NAND2_X1 U17855 ( .A1(n15883), .A2(n15968), .ZN(n15891) );
  AOI21_X1 U17856 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21322) );
  NOR2_X1 U17857 ( .A1(n21322), .A2(n21337), .ZN(n21358) );
  NAND2_X1 U17858 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21358), .ZN(
        n21351) );
  NOR2_X1 U17859 ( .A1(n16002), .A2(n21351), .ZN(n16007) );
  NAND2_X1 U17860 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16007), .ZN(
        n21406) );
  NOR2_X1 U17861 ( .A1(n13559), .A2(n21406), .ZN(n21298) );
  NAND2_X1 U17862 ( .A1(n15973), .A2(n21298), .ZN(n15970) );
  NOR3_X1 U17863 ( .A1(n15970), .A2(n13418), .A3(n15977), .ZN(n15892) );
  AOI21_X1 U17864 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15892), .A(
        n21334), .ZN(n15884) );
  AOI21_X1 U17865 ( .B1(n21330), .B2(n15891), .A(n15884), .ZN(n15885) );
  NAND2_X1 U17866 ( .A1(n21348), .A2(n15885), .ZN(n21458) );
  INV_X1 U17867 ( .A(n15886), .ZN(n15936) );
  NOR2_X1 U17868 ( .A1(n21426), .A2(n15936), .ZN(n15887) );
  NOR2_X1 U17869 ( .A1(n21458), .A2(n15887), .ZN(n15948) );
  AND2_X1 U17870 ( .A1(n15948), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15939) );
  NAND2_X1 U17871 ( .A1(n21348), .A2(n21426), .ZN(n21350) );
  INV_X1 U17872 ( .A(n21350), .ZN(n21372) );
  NOR2_X1 U17873 ( .A1(n15939), .A2(n21372), .ZN(n15932) );
  NOR2_X1 U17874 ( .A1(n15932), .A2(n15903), .ZN(n15899) );
  INV_X1 U17875 ( .A(n15900), .ZN(n15889) );
  AOI211_X1 U17876 ( .C1(n15899), .C2(n15889), .A(n21372), .B(n15888), .ZN(
        n15895) );
  NAND2_X1 U17877 ( .A1(n21330), .A2(n15890), .ZN(n21319) );
  NOR2_X1 U17878 ( .A1(n15891), .A2(n21319), .ZN(n15954) );
  AOI21_X1 U17879 ( .B1(n21407), .B2(n15892), .A(n15954), .ZN(n21466) );
  INV_X1 U17880 ( .A(n21466), .ZN(n15956) );
  NAND3_X1 U17881 ( .A1(n15956), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15936), .ZN(n15928) );
  NOR4_X1 U17882 ( .A1(n15928), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15903), .A4(n15900), .ZN(n15893) );
  OAI21_X1 U17883 ( .B1(n15898), .B2(n21430), .A(n15897), .ZN(P1_U3000) );
  NOR3_X1 U17884 ( .A1(n15899), .A2(n15900), .A3(n15928), .ZN(n15905) );
  INV_X1 U17885 ( .A(n15939), .ZN(n15901) );
  OAI21_X1 U17886 ( .B1(n15901), .B2(n15900), .A(n21350), .ZN(n15914) );
  OAI21_X1 U17887 ( .B1(n15914), .B2(n15903), .A(n15902), .ZN(n15904) );
  AOI211_X1 U17888 ( .C1(n15906), .C2(n21461), .A(n15905), .B(n15904), .ZN(
        n15907) );
  OAI21_X1 U17889 ( .B1(n15908), .B2(n21430), .A(n15907), .ZN(P1_U3001) );
  INV_X1 U17890 ( .A(n15928), .ZN(n15910) );
  NAND3_X1 U17891 ( .A1(n15910), .A2(n15909), .A3(n15913), .ZN(n15911) );
  OAI211_X1 U17892 ( .C1(n15914), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        n15915) );
  AOI21_X1 U17893 ( .B1(n15916), .B2(n21461), .A(n15915), .ZN(n15917) );
  OAI21_X1 U17894 ( .B1(n15918), .B2(n21430), .A(n15917), .ZN(P1_U3002) );
  XNOR2_X1 U17895 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15919) );
  NOR2_X1 U17896 ( .A1(n15928), .A2(n15919), .ZN(n15920) );
  AOI211_X1 U17897 ( .C1(n15932), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15921), .B(n15920), .ZN(n15925) );
  INV_X1 U17898 ( .A(n15922), .ZN(n15923) );
  NAND2_X1 U17899 ( .A1(n15923), .A2(n21461), .ZN(n15924) );
  OAI211_X1 U17900 ( .C1(n15926), .C2(n21430), .A(n15925), .B(n15924), .ZN(
        P1_U3003) );
  OAI21_X1 U17901 ( .B1(n15928), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15927), .ZN(n15931) );
  NOR2_X1 U17902 ( .A1(n15929), .A2(n21429), .ZN(n15930) );
  AOI211_X1 U17903 ( .C1(n15932), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15931), .B(n15930), .ZN(n15933) );
  OAI21_X1 U17904 ( .B1(n15934), .B2(n21430), .A(n15933), .ZN(P1_U3004) );
  INV_X1 U17905 ( .A(n15935), .ZN(n15941) );
  AOI21_X1 U17906 ( .B1(n15956), .B2(n15936), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15938) );
  OAI21_X1 U17907 ( .B1(n15939), .B2(n15938), .A(n15937), .ZN(n15940) );
  AOI21_X1 U17908 ( .B1(n15941), .B2(n21461), .A(n15940), .ZN(n15942) );
  OAI21_X1 U17909 ( .B1(n15943), .B2(n21430), .A(n15942), .ZN(P1_U3005) );
  NAND3_X1 U17910 ( .A1(n15956), .A2(n15944), .A3(n15947), .ZN(n15945) );
  OAI211_X1 U17911 ( .C1(n15948), .C2(n15947), .A(n15946), .B(n15945), .ZN(
        n15949) );
  AOI21_X1 U17912 ( .B1(n15950), .B2(n21461), .A(n15949), .ZN(n15951) );
  OAI21_X1 U17913 ( .B1(n15952), .B2(n21430), .A(n15951), .ZN(P1_U3006) );
  INV_X1 U17914 ( .A(n21666), .ZN(n15962) );
  AOI21_X1 U17915 ( .B1(n15954), .B2(n15953), .A(n21458), .ZN(n15960) );
  INV_X1 U17916 ( .A(n15955), .ZN(n15958) );
  NAND3_X1 U17917 ( .A1(n15956), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15959), .ZN(n15957) );
  OAI211_X1 U17918 ( .C1(n15960), .C2(n15959), .A(n15958), .B(n15957), .ZN(
        n15961) );
  AOI21_X1 U17919 ( .B1(n15962), .B2(n21461), .A(n15961), .ZN(n15963) );
  OAI21_X1 U17920 ( .B1(n15964), .B2(n21430), .A(n15963), .ZN(P1_U3007) );
  NAND2_X1 U17921 ( .A1(n15966), .A2(n15965), .ZN(n15967) );
  XNOR2_X1 U17922 ( .A(n15967), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19977) );
  INV_X1 U17923 ( .A(n19977), .ZN(n15983) );
  NAND2_X1 U17924 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15975) );
  OAI21_X1 U17925 ( .B1(n21349), .B2(n15968), .A(n21348), .ZN(n15969) );
  AOI21_X1 U17926 ( .B1(n21407), .B2(n15970), .A(n15969), .ZN(n15991) );
  INV_X1 U17927 ( .A(n15991), .ZN(n21442) );
  OAI21_X1 U17928 ( .B1(n15975), .B2(n21442), .A(n21350), .ZN(n21455) );
  INV_X1 U17929 ( .A(n21455), .ZN(n15976) );
  INV_X1 U17930 ( .A(n21298), .ZN(n15972) );
  NAND2_X1 U17931 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21304), .ZN(
        n15971) );
  OAI22_X1 U17932 ( .A1(n21334), .A2(n15972), .B1(n21297), .B2(n15971), .ZN(
        n21301) );
  NAND2_X1 U17933 ( .A1(n15973), .A2(n21301), .ZN(n15992) );
  OAI21_X1 U17934 ( .B1(n15974), .B2(n21296), .A(n15992), .ZN(n15990) );
  INV_X1 U17935 ( .A(n15990), .ZN(n21448) );
  NOR3_X1 U17936 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21448), .A3(
        n15975), .ZN(n21449) );
  OAI21_X1 U17937 ( .B1(n15976), .B2(n21449), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15982) );
  NOR2_X1 U17938 ( .A1(n21616), .A2(n21635), .ZN(n15979) );
  NOR3_X1 U17939 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21448), .A3(
        n15977), .ZN(n15978) );
  AOI211_X1 U17940 ( .C1(n15980), .C2(n21461), .A(n15979), .B(n15978), .ZN(
        n15981) );
  OAI211_X1 U17941 ( .C1(n15983), .C2(n21430), .A(n15982), .B(n15981), .ZN(
        P1_U3009) );
  OAI21_X1 U17942 ( .B1(n15985), .B2(n19950), .A(n15984), .ZN(n15986) );
  XNOR2_X1 U17943 ( .A(n15986), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n19972) );
  INV_X1 U17944 ( .A(n19972), .ZN(n15996) );
  INV_X1 U17945 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15987) );
  OAI22_X1 U17946 ( .A1(n21627), .A2(n21429), .B1(n21616), .B2(n15987), .ZN(
        n15988) );
  AOI21_X1 U17947 ( .B1(n15990), .B2(n15989), .A(n15988), .ZN(n15995) );
  OAI221_X1 U17948 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21296), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15992), .A(n15991), .ZN(
        n15993) );
  NAND2_X1 U17949 ( .A1(n15993), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15994) );
  OAI211_X1 U17950 ( .C1(n15996), .C2(n21430), .A(n15995), .B(n15994), .ZN(
        P1_U3011) );
  OAI21_X1 U17951 ( .B1(n15999), .B2(n15998), .A(n15997), .ZN(n16001) );
  XNOR2_X1 U17952 ( .A(n16001), .B(n16000), .ZN(n19969) );
  NAND3_X1 U17953 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16008) );
  INV_X1 U17954 ( .A(n16002), .ZN(n16004) );
  NAND2_X1 U17955 ( .A1(n16004), .A2(n21396), .ZN(n21412) );
  NOR2_X1 U17956 ( .A1(n16008), .A2(n21412), .ZN(n21315) );
  NAND2_X1 U17957 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21315), .ZN(
        n21423) );
  NOR3_X1 U17958 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16005), .A3(
        n21423), .ZN(n16014) );
  NOR2_X1 U17959 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21423), .ZN(
        n16017) );
  INV_X1 U17960 ( .A(n21426), .ZN(n16009) );
  INV_X1 U17961 ( .A(n21348), .ZN(n21300) );
  AOI21_X1 U17962 ( .B1(n21330), .B2(n16006), .A(n21300), .ZN(n21409) );
  OAI21_X1 U17963 ( .B1(n16007), .B2(n21334), .A(n21409), .ZN(n21419) );
  AOI221_X1 U17964 ( .B1(n13561), .B2(n16009), .C1(n16008), .C2(n16009), .A(
        n21419), .ZN(n21425) );
  INV_X1 U17965 ( .A(n21425), .ZN(n16010) );
  OAI21_X1 U17966 ( .B1(n16017), .B2(n16010), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16012) );
  OR2_X1 U17967 ( .A1(n21616), .A2(n21600), .ZN(n16011) );
  OAI211_X1 U17968 ( .C1(n21614), .C2(n21429), .A(n16012), .B(n16011), .ZN(
        n16013) );
  AOI211_X1 U17969 ( .C1(n19969), .C2(n21462), .A(n16014), .B(n16013), .ZN(
        n16015) );
  INV_X1 U17970 ( .A(n16015), .ZN(P1_U3015) );
  NAND2_X1 U17971 ( .A1(n16016), .A2(n21462), .ZN(n16021) );
  INV_X1 U17972 ( .A(n21598), .ZN(n16019) );
  AOI211_X1 U17973 ( .C1(n21461), .C2(n16019), .A(n16018), .B(n16017), .ZN(
        n16020) );
  OAI211_X1 U17974 ( .C1(n21425), .C2(n16005), .A(n16021), .B(n16020), .ZN(
        P1_U3016) );
  NAND2_X1 U17975 ( .A1(n16022), .A2(n21982), .ZN(n21895) );
  NOR2_X1 U17976 ( .A1(n14520), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16023) );
  OAI22_X1 U17977 ( .A1(n21895), .A2(n16023), .B1(n14973), .B2(n16029), .ZN(
        n16024) );
  MUX2_X1 U17978 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16024), .S(
        n16840), .Z(P1_U3477) );
  NAND2_X1 U17979 ( .A1(n16025), .A2(n21982), .ZN(n16026) );
  MUX2_X1 U17980 ( .A(n21895), .B(n16026), .S(n14519), .Z(n16027) );
  OAI21_X1 U17981 ( .B1(n16029), .B2(n16028), .A(n16027), .ZN(n16030) );
  MUX2_X1 U17982 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n16030), .S(
        n16840), .Z(P1_U3476) );
  NAND3_X1 U17983 ( .A1(n16033), .A2(n16032), .A3(n16031), .ZN(n16034) );
  OAI21_X1 U17984 ( .B1(n16035), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n16034), .ZN(n16036) );
  AOI21_X1 U17985 ( .B1(n21962), .B2(n16037), .A(n16036), .ZN(n16805) );
  INV_X1 U17986 ( .A(n16038), .ZN(n21673) );
  INV_X1 U17987 ( .A(n16039), .ZN(n16042) );
  NOR3_X1 U17988 ( .A1(n14463), .A2(n14238), .A3(n21671), .ZN(n16040) );
  AOI21_X1 U17989 ( .B1(n16042), .B2(n16041), .A(n16040), .ZN(n16043) );
  OAI21_X1 U17990 ( .B1(n16805), .B2(n21673), .A(n16043), .ZN(n16045) );
  MUX2_X1 U17991 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16045), .S(
        n16044), .Z(P1_U3473) );
  INV_X1 U17992 ( .A(n16046), .ZN(n16059) );
  OAI211_X1 U17993 ( .C1(n16353), .C2(n16048), .A(n18362), .B(n16047), .ZN(
        n16058) );
  AOI21_X1 U17994 ( .B1(n16152), .B2(n16151), .A(n16049), .ZN(n16051) );
  NOR2_X1 U17995 ( .A1(n16051), .A2(n16050), .ZN(n16352) );
  NOR2_X1 U17996 ( .A1(n16052), .A2(n16237), .ZN(n16053) );
  OR2_X1 U17997 ( .A1(n16228), .A2(n16053), .ZN(n19346) );
  OAI22_X1 U17998 ( .A1(n18537), .A2(n13211), .B1(n18562), .B2(n19346), .ZN(
        n16056) );
  OAI22_X1 U17999 ( .A1(n16054), .A2(n18488), .B1(n13077), .B2(n18520), .ZN(
        n16055) );
  AOI211_X1 U18000 ( .C1(n16352), .C2(n18551), .A(n16056), .B(n16055), .ZN(
        n16057) );
  OAI211_X1 U18001 ( .C1(n16059), .C2(n18522), .A(n16058), .B(n16057), .ZN(
        P2_U2833) );
  OAI211_X1 U18002 ( .C1(n16061), .C2(n16377), .A(n18362), .B(n16060), .ZN(
        n16073) );
  NOR2_X1 U18003 ( .A1(n16161), .A2(n16062), .ZN(n16063) );
  OR2_X1 U18004 ( .A1(n16152), .A2(n16063), .ZN(n16553) );
  INV_X1 U18005 ( .A(n16553), .ZN(n16071) );
  NOR2_X1 U18006 ( .A1(n16066), .A2(n16065), .ZN(n16067) );
  NOR2_X1 U18007 ( .A1(n16064), .A2(n16067), .ZN(n19446) );
  OAI22_X1 U18008 ( .A1(n13098), .A2(n18488), .B1(n17221), .B2(n18520), .ZN(
        n16068) );
  AOI21_X1 U18009 ( .B1(n18580), .B2(n19446), .A(n16068), .ZN(n16069) );
  OAI21_X1 U18010 ( .B1(n18537), .B2(n13207), .A(n16069), .ZN(n16070) );
  AOI21_X1 U18011 ( .B1(n16071), .B2(n18551), .A(n16070), .ZN(n16072) );
  OAI211_X1 U18012 ( .C1(n18522), .C2(n16074), .A(n16073), .B(n16072), .ZN(
        P2_U2835) );
  OAI211_X1 U18013 ( .C1(n16077), .C2(n16076), .A(n18362), .B(n16075), .ZN(
        n16088) );
  NOR2_X1 U18014 ( .A1(n16078), .A2(n14936), .ZN(n16079) );
  NOR2_X1 U18015 ( .A1(n16080), .A2(n16079), .ZN(n19618) );
  NOR2_X1 U18016 ( .A1(n16602), .A2(n18578), .ZN(n16086) );
  AOI21_X1 U18017 ( .B1(P2_REIP_REG_16__SCAN_IN), .B2(n18576), .A(n16396), 
        .ZN(n16083) );
  AOI22_X1 U18018 ( .A1(n16081), .A2(n13297), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18561), .ZN(n16082) );
  OAI211_X1 U18019 ( .C1(n16084), .C2(n18488), .A(n16083), .B(n16082), .ZN(
        n16085) );
  AOI211_X1 U18020 ( .C1(n19618), .C2(n18580), .A(n16086), .B(n16085), .ZN(
        n16087) );
  NAND2_X1 U18021 ( .A1(n16088), .A2(n16087), .ZN(P2_U2839) );
  INV_X1 U18022 ( .A(n18579), .ZN(n16089) );
  NAND2_X1 U18023 ( .A1(n16089), .A2(n16127), .ZN(n16090) );
  OAI21_X1 U18024 ( .B1(n16127), .B2(n16091), .A(n16090), .ZN(P2_U2856) );
  NAND2_X1 U18025 ( .A1(n16102), .A2(n16092), .ZN(n16093) );
  NOR2_X1 U18026 ( .A1(n18564), .A2(n16176), .ZN(n16094) );
  AOI21_X1 U18027 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16176), .A(n16094), .ZN(
        n16095) );
  OAI21_X1 U18028 ( .B1(n16096), .B2(n16178), .A(n16095), .ZN(P2_U2858) );
  INV_X1 U18029 ( .A(n16097), .ZN(n16107) );
  NAND2_X1 U18030 ( .A1(n16107), .A2(n16098), .ZN(n16100) );
  XNOR2_X1 U18031 ( .A(n16100), .B(n16099), .ZN(n16187) );
  NOR2_X1 U18032 ( .A1(n16450), .A2(n16176), .ZN(n16104) );
  AOI21_X1 U18033 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16176), .A(n16104), .ZN(
        n16105) );
  OAI21_X1 U18034 ( .B1(n16187), .B2(n16178), .A(n16105), .ZN(P2_U2859) );
  NAND2_X1 U18035 ( .A1(n16107), .A2(n16106), .ZN(n16108) );
  XOR2_X1 U18036 ( .A(n16109), .B(n16108), .Z(n16195) );
  NOR2_X1 U18037 ( .A1(n16110), .A2(n16111), .ZN(n16112) );
  NOR2_X1 U18038 ( .A1(n18535), .A2(n16176), .ZN(n16113) );
  AOI21_X1 U18039 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16176), .A(n16113), .ZN(
        n16114) );
  OAI21_X1 U18040 ( .B1(n16195), .B2(n16178), .A(n16114), .ZN(P2_U2860) );
  NOR2_X1 U18041 ( .A1(n16125), .A2(n16115), .ZN(n16116) );
  OR2_X1 U18042 ( .A1(n16110), .A2(n16116), .ZN(n18526) );
  AOI21_X1 U18043 ( .B1(n16119), .B2(n16118), .A(n16117), .ZN(n16196) );
  NAND2_X1 U18044 ( .A1(n16196), .A2(n16169), .ZN(n16121) );
  NAND2_X1 U18045 ( .A1(n16176), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16120) );
  OAI211_X1 U18046 ( .C1(n18526), .C2(n16176), .A(n16121), .B(n16120), .ZN(
        P2_U2861) );
  OAI21_X1 U18047 ( .B1(n16124), .B2(n16123), .A(n16122), .ZN(n16216) );
  NAND2_X1 U18048 ( .A1(n16176), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16129) );
  AOI21_X1 U18049 ( .B1(n16126), .B2(n16133), .A(n16125), .ZN(n18512) );
  NAND2_X1 U18050 ( .A1(n18512), .A2(n16127), .ZN(n16128) );
  OAI211_X1 U18051 ( .C1(n16216), .C2(n16178), .A(n16129), .B(n16128), .ZN(
        P2_U2862) );
  OAI21_X1 U18052 ( .B1(n16130), .B2(n16132), .A(n16131), .ZN(n16226) );
  NAND2_X1 U18053 ( .A1(n16176), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16137) );
  INV_X1 U18054 ( .A(n16133), .ZN(n16134) );
  AOI21_X1 U18055 ( .B1(n16135), .B2(n16140), .A(n16134), .ZN(n18502) );
  NAND2_X1 U18056 ( .A1(n18502), .A2(n16127), .ZN(n16136) );
  OAI211_X1 U18057 ( .C1(n16226), .C2(n16178), .A(n16137), .B(n16136), .ZN(
        P2_U2863) );
  XNOR2_X1 U18058 ( .A(n16138), .B(n16139), .ZN(n16235) );
  OAI21_X1 U18059 ( .B1(n16141), .B2(n16050), .A(n16140), .ZN(n18489) );
  NOR2_X1 U18060 ( .A1(n16176), .A2(n18489), .ZN(n16142) );
  AOI21_X1 U18061 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16176), .A(n16142), .ZN(
        n16143) );
  OAI21_X1 U18062 ( .B1(n16235), .B2(n16178), .A(n16143), .ZN(P2_U2864) );
  OAI21_X1 U18063 ( .B1(n16144), .B2(n16145), .A(n16138), .ZN(n19345) );
  NAND2_X1 U18064 ( .A1(n16176), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16147) );
  NAND2_X1 U18065 ( .A1(n16352), .A2(n16127), .ZN(n16146) );
  OAI211_X1 U18066 ( .C1(n19345), .C2(n16178), .A(n16147), .B(n16146), .ZN(
        P2_U2865) );
  INV_X1 U18067 ( .A(n16144), .ZN(n16149) );
  OAI21_X1 U18068 ( .B1(n16148), .B2(n16150), .A(n16149), .ZN(n16245) );
  XNOR2_X1 U18069 ( .A(n16152), .B(n16151), .ZN(n18478) );
  NOR2_X1 U18070 ( .A1(n18478), .A2(n16176), .ZN(n16153) );
  AOI21_X1 U18071 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n16176), .A(n16153), .ZN(
        n16154) );
  OAI21_X1 U18072 ( .B1(n16245), .B2(n16178), .A(n16154), .ZN(P2_U2866) );
  AOI21_X1 U18073 ( .B1(n16155), .B2(n11032), .A(n16148), .ZN(n19447) );
  NAND2_X1 U18074 ( .A1(n19447), .A2(n16169), .ZN(n16157) );
  NAND2_X1 U18075 ( .A1(n16176), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16156) );
  OAI211_X1 U18076 ( .C1(n16553), .C2(n16176), .A(n16157), .B(n16156), .ZN(
        P2_U2867) );
  OAI21_X1 U18077 ( .B1(n16158), .B2(n16159), .A(n11032), .ZN(n16256) );
  AND2_X1 U18078 ( .A1(n16165), .A2(n16160), .ZN(n16162) );
  OR2_X1 U18079 ( .A1(n16162), .A2(n16161), .ZN(n18466) );
  NOR2_X1 U18080 ( .A1(n18466), .A2(n16176), .ZN(n16163) );
  AOI21_X1 U18081 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16176), .A(n16163), .ZN(
        n16164) );
  OAI21_X1 U18082 ( .B1(n16256), .B2(n16178), .A(n16164), .ZN(P2_U2868) );
  INV_X1 U18083 ( .A(n16165), .ZN(n16166) );
  AOI21_X1 U18084 ( .B1(n16167), .B2(n16174), .A(n16166), .ZN(n16572) );
  INV_X1 U18085 ( .A(n16572), .ZN(n18454) );
  AOI21_X1 U18086 ( .B1(n16168), .B2(n15211), .A(n16158), .ZN(n16257) );
  NAND2_X1 U18087 ( .A1(n16257), .A2(n16169), .ZN(n16171) );
  NAND2_X1 U18088 ( .A1(n16176), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16170) );
  OAI211_X1 U18089 ( .C1(n18454), .C2(n16176), .A(n16171), .B(n16170), .ZN(
        P2_U2869) );
  NAND2_X1 U18090 ( .A1(n14080), .A2(n16172), .ZN(n16173) );
  NAND2_X1 U18091 ( .A1(n16174), .A2(n16173), .ZN(n18442) );
  NOR2_X1 U18092 ( .A1(n18442), .A2(n16176), .ZN(n16175) );
  AOI21_X1 U18093 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16176), .A(n16175), .ZN(
        n16177) );
  OAI21_X1 U18094 ( .B1(n16179), .B2(n16178), .A(n16177), .ZN(P2_U2870) );
  AOI22_X1 U18095 ( .A1(n19616), .A2(BUF1_REG_28__SCAN_IN), .B1(n19615), .B2(
        n19122), .ZN(n16186) );
  NOR2_X1 U18096 ( .A1(n16180), .A2(n16181), .ZN(n16182) );
  OAI22_X1 U18097 ( .A1(n16201), .A2(n18549), .B1(n16250), .B2(n14396), .ZN(
        n16184) );
  AOI21_X1 U18098 ( .B1(n19617), .B2(BUF2_REG_28__SCAN_IN), .A(n16184), .ZN(
        n16185) );
  OAI211_X1 U18099 ( .C1(n16187), .C2(n19398), .A(n16186), .B(n16185), .ZN(
        P2_U2891) );
  AOI22_X1 U18100 ( .A1(n19616), .A2(BUF1_REG_27__SCAN_IN), .B1(n19615), .B2(
        n16188), .ZN(n16194) );
  AND2_X1 U18101 ( .A1(n16200), .A2(n16189), .ZN(n16190) );
  OR2_X1 U18102 ( .A1(n16190), .A2(n16180), .ZN(n18546) );
  OAI22_X1 U18103 ( .A1(n16201), .A2(n18546), .B1(n16250), .B2(n16191), .ZN(
        n16192) );
  AOI21_X1 U18104 ( .B1(n19617), .B2(BUF2_REG_27__SCAN_IN), .A(n16192), .ZN(
        n16193) );
  OAI211_X1 U18105 ( .C1(n16195), .C2(n19398), .A(n16194), .B(n16193), .ZN(
        P2_U2892) );
  INV_X1 U18106 ( .A(n16196), .ZN(n16205) );
  AOI22_X1 U18107 ( .A1(n19616), .A2(BUF1_REG_26__SCAN_IN), .B1(n19615), .B2(
        n19125), .ZN(n16204) );
  NAND2_X1 U18108 ( .A1(n16209), .A2(n16198), .ZN(n16199) );
  NAND2_X1 U18109 ( .A1(n16200), .A2(n16199), .ZN(n18525) );
  OAI22_X1 U18110 ( .A1(n16201), .A2(n18525), .B1(n16250), .B2(n14390), .ZN(
        n16202) );
  AOI21_X1 U18111 ( .B1(n19617), .B2(BUF2_REG_26__SCAN_IN), .A(n16202), .ZN(
        n16203) );
  OAI211_X1 U18112 ( .C1(n16205), .C2(n19398), .A(n16204), .B(n16203), .ZN(
        P2_U2893) );
  NAND2_X1 U18113 ( .A1(n16206), .A2(n16207), .ZN(n16208) );
  AND2_X1 U18114 ( .A1(n16209), .A2(n16208), .ZN(n18511) );
  NAND2_X1 U18115 ( .A1(n19619), .A2(n18511), .ZN(n16210) );
  OAI21_X1 U18116 ( .B1(n16250), .B2(n16211), .A(n16210), .ZN(n16214) );
  OAI22_X1 U18117 ( .A1(n16252), .A2(n20037), .B1(n16212), .B2(n16251), .ZN(
        n16213) );
  AOI211_X1 U18118 ( .C1(n19617), .C2(BUF2_REG_25__SCAN_IN), .A(n16214), .B(
        n16213), .ZN(n16215) );
  OAI21_X1 U18119 ( .B1(n16216), .B2(n19398), .A(n16215), .ZN(P2_U2894) );
  OR2_X1 U18120 ( .A1(n16217), .A2(n16218), .ZN(n16219) );
  AND2_X1 U18121 ( .A1(n16206), .A2(n16219), .ZN(n18501) );
  NAND2_X1 U18122 ( .A1(n19619), .A2(n18501), .ZN(n16220) );
  OAI21_X1 U18123 ( .B1(n16250), .B2(n16221), .A(n16220), .ZN(n16224) );
  OAI22_X1 U18124 ( .A1(n16252), .A2(n20035), .B1(n16222), .B2(n16251), .ZN(
        n16223) );
  AOI211_X1 U18125 ( .C1(n19617), .C2(BUF2_REG_24__SCAN_IN), .A(n16224), .B(
        n16223), .ZN(n16225) );
  OAI21_X1 U18126 ( .B1(n16226), .B2(n19398), .A(n16225), .ZN(P2_U2895) );
  NOR2_X1 U18127 ( .A1(n16228), .A2(n16227), .ZN(n16229) );
  OR2_X1 U18128 ( .A1(n16217), .A2(n16229), .ZN(n18499) );
  INV_X1 U18129 ( .A(n18499), .ZN(n16510) );
  NAND2_X1 U18130 ( .A1(n19619), .A2(n16510), .ZN(n16230) );
  OAI21_X1 U18131 ( .B1(n16250), .B2(n16231), .A(n16230), .ZN(n16233) );
  OAI22_X1 U18132 ( .A1(n16252), .A2(n20033), .B1(n19131), .B2(n16251), .ZN(
        n16232) );
  AOI211_X1 U18133 ( .C1(n19617), .C2(BUF2_REG_23__SCAN_IN), .A(n16233), .B(
        n16232), .ZN(n16234) );
  OAI21_X1 U18134 ( .B1(n16235), .B2(n19398), .A(n16234), .ZN(P2_U2896) );
  OR2_X1 U18135 ( .A1(n16064), .A2(n16236), .ZN(n16239) );
  NAND2_X1 U18136 ( .A1(n16239), .A2(n16238), .ZN(n18486) );
  INV_X1 U18137 ( .A(n18486), .ZN(n16532) );
  NAND2_X1 U18138 ( .A1(n19619), .A2(n16532), .ZN(n16240) );
  OAI21_X1 U18139 ( .B1(n16250), .B2(n16241), .A(n16240), .ZN(n16243) );
  OAI22_X1 U18140 ( .A1(n16252), .A2(n20029), .B1(n19405), .B2(n16251), .ZN(
        n16242) );
  AOI211_X1 U18141 ( .C1(n19617), .C2(BUF2_REG_21__SCAN_IN), .A(n16243), .B(
        n16242), .ZN(n16244) );
  OAI21_X1 U18142 ( .B1(n16245), .B2(n19398), .A(n16244), .ZN(P2_U2898) );
  XNOR2_X1 U18143 ( .A(n11065), .B(n16246), .ZN(n18465) );
  INV_X1 U18144 ( .A(n18465), .ZN(n16247) );
  NAND2_X1 U18145 ( .A1(n19619), .A2(n16247), .ZN(n16248) );
  OAI21_X1 U18146 ( .B1(n16250), .B2(n16249), .A(n16248), .ZN(n16254) );
  OAI22_X1 U18147 ( .A1(n16252), .A2(n20025), .B1(n17042), .B2(n16251), .ZN(
        n16253) );
  AOI211_X1 U18148 ( .C1(n19617), .C2(BUF2_REG_19__SCAN_IN), .A(n16254), .B(
        n16253), .ZN(n16255) );
  OAI21_X1 U18149 ( .B1(n16256), .B2(n19398), .A(n16255), .ZN(P2_U2900) );
  NAND2_X1 U18150 ( .A1(n16257), .A2(n19620), .ZN(n16266) );
  INV_X1 U18151 ( .A(n19532), .ZN(n16258) );
  AOI22_X1 U18152 ( .A1(n19616), .A2(BUF1_REG_18__SCAN_IN), .B1(n19615), .B2(
        n16258), .ZN(n16265) );
  AND2_X1 U18153 ( .A1(n16260), .A2(n16259), .ZN(n16261) );
  OR2_X1 U18154 ( .A1(n16261), .A2(n11065), .ZN(n18453) );
  INV_X1 U18155 ( .A(n18453), .ZN(n16262) );
  AOI22_X1 U18156 ( .A1(n19619), .A2(n16262), .B1(n19613), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16264) );
  NAND2_X1 U18157 ( .A1(n19617), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16263) );
  NAND4_X1 U18158 ( .A1(n16266), .A2(n16265), .A3(n16264), .A4(n16263), .ZN(
        P2_U2901) );
  NOR2_X1 U18159 ( .A1(n16268), .A2(n16267), .ZN(n16270) );
  XOR2_X1 U18160 ( .A(n16270), .B(n16269), .Z(n16447) );
  INV_X1 U18161 ( .A(n16271), .ZN(n16273) );
  AOI21_X1 U18162 ( .B1(n16303), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16272) );
  NOR2_X1 U18163 ( .A1(n16273), .A2(n16272), .ZN(n16445) );
  INV_X1 U18164 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16274) );
  OR2_X1 U18165 ( .A1(n18381), .A2(n17227), .ZN(n16439) );
  OAI21_X1 U18166 ( .B1(n17117), .B2(n16274), .A(n16439), .ZN(n16275) );
  AOI21_X1 U18167 ( .B1(n17105), .B2(n16276), .A(n16275), .ZN(n16277) );
  OAI21_X1 U18168 ( .B1(n18564), .B2(n17113), .A(n16277), .ZN(n16278) );
  AOI21_X1 U18169 ( .B1(n16445), .B2(n17131), .A(n16278), .ZN(n16279) );
  OAI21_X1 U18170 ( .B1(n16447), .B2(n17120), .A(n16279), .ZN(P2_U2985) );
  INV_X1 U18171 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16484) );
  OAI21_X1 U18172 ( .B1(n16329), .B2(n16484), .A(n16281), .ZN(n16282) );
  OAI21_X1 U18173 ( .B1(n16283), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16282), .ZN(n16306) );
  NAND2_X1 U18174 ( .A1(n16284), .A2(n16314), .ZN(n16286) );
  OAI21_X1 U18175 ( .B1(n16306), .B2(n16286), .A(n16285), .ZN(n16298) );
  INV_X1 U18176 ( .A(n16296), .ZN(n16287) );
  AOI22_X1 U18177 ( .A1(n16298), .A2(n16288), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16287), .ZN(n16290) );
  XNOR2_X1 U18178 ( .A(n16290), .B(n16289), .ZN(n16459) );
  XOR2_X1 U18179 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n16303), .Z(
        n16457) );
  NOR2_X1 U18180 ( .A1(n14035), .A2(n16291), .ZN(n16453) );
  NOR2_X1 U18181 ( .A1(n17125), .A2(n18555), .ZN(n16292) );
  AOI211_X1 U18182 ( .C1(n17126), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16453), .B(n16292), .ZN(n16293) );
  OAI21_X1 U18183 ( .B1(n16450), .B2(n17113), .A(n16293), .ZN(n16294) );
  AOI21_X1 U18184 ( .B1(n16457), .B2(n17131), .A(n16294), .ZN(n16295) );
  OAI21_X1 U18185 ( .B1(n16459), .B2(n17120), .A(n16295), .ZN(P2_U2986) );
  XNOR2_X1 U18186 ( .A(n16296), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16297) );
  XNOR2_X1 U18187 ( .A(n16298), .B(n16297), .ZN(n16470) );
  NAND2_X1 U18188 ( .A1(n16396), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16461) );
  OAI21_X1 U18189 ( .B1(n17117), .B2(n16299), .A(n16461), .ZN(n16301) );
  NOR2_X1 U18190 ( .A1(n18535), .A2(n17113), .ZN(n16300) );
  AOI211_X1 U18191 ( .C1(n17105), .C2(n16302), .A(n16301), .B(n16300), .ZN(
        n16305) );
  INV_X1 U18192 ( .A(n16303), .ZN(n16467) );
  NAND2_X1 U18193 ( .A1(n16310), .A2(n16438), .ZN(n16466) );
  NAND3_X1 U18194 ( .A1(n16467), .A2(n17131), .A3(n16466), .ZN(n16304) );
  OAI211_X1 U18195 ( .C1(n16470), .C2(n17120), .A(n16305), .B(n16304), .ZN(
        P2_U2987) );
  INV_X1 U18196 ( .A(n16306), .ZN(n16318) );
  OAI21_X1 U18197 ( .B1(n16318), .B2(n16316), .A(n16314), .ZN(n16308) );
  XNOR2_X1 U18198 ( .A(n16308), .B(n16307), .ZN(n16482) );
  INV_X1 U18199 ( .A(n18526), .ZN(n16475) );
  INV_X1 U18200 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18521) );
  NOR2_X1 U18201 ( .A1(n14035), .A2(n18521), .ZN(n16474) );
  AOI21_X1 U18202 ( .B1(n17126), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16474), .ZN(n16309) );
  OAI21_X1 U18203 ( .B1(n17125), .B2(n18530), .A(n16309), .ZN(n16312) );
  OAI21_X1 U18204 ( .B1(n16319), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16310), .ZN(n16477) );
  NOR2_X1 U18205 ( .A1(n16477), .A2(n17119), .ZN(n16311) );
  AOI211_X1 U18206 ( .C1(n17133), .C2(n16475), .A(n16312), .B(n16311), .ZN(
        n16313) );
  OAI21_X1 U18207 ( .B1(n16482), .B2(n17120), .A(n16313), .ZN(P2_U2988) );
  INV_X1 U18208 ( .A(n16314), .ZN(n16315) );
  NOR2_X1 U18209 ( .A1(n16316), .A2(n16315), .ZN(n16317) );
  XNOR2_X1 U18210 ( .A(n16318), .B(n16317), .ZN(n16494) );
  AOI21_X1 U18211 ( .B1(n16489), .B2(n16331), .A(n16319), .ZN(n16492) );
  INV_X1 U18212 ( .A(n18512), .ZN(n16324) );
  INV_X1 U18213 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17224) );
  NOR2_X1 U18214 ( .A1(n14035), .A2(n17224), .ZN(n16486) );
  NOR2_X1 U18215 ( .A1(n17117), .A2(n16320), .ZN(n16321) );
  AOI211_X1 U18216 ( .C1(n16322), .C2(n17105), .A(n16486), .B(n16321), .ZN(
        n16323) );
  OAI21_X1 U18217 ( .B1(n17113), .B2(n16324), .A(n16323), .ZN(n16325) );
  AOI21_X1 U18218 ( .B1(n16492), .B2(n17131), .A(n16325), .ZN(n16326) );
  OAI21_X1 U18219 ( .B1(n16494), .B2(n17120), .A(n16326), .ZN(P2_U2989) );
  XNOR2_X1 U18220 ( .A(n16327), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16328) );
  XNOR2_X1 U18221 ( .A(n16329), .B(n16328), .ZN(n16504) );
  NOR2_X1 U18222 ( .A1(n14035), .A2(n17223), .ZN(n16495) );
  AOI21_X1 U18223 ( .B1(n17126), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16495), .ZN(n16330) );
  OAI21_X1 U18224 ( .B1(n17125), .B2(n18505), .A(n16330), .ZN(n16333) );
  OAI21_X1 U18225 ( .B1(n16335), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16331), .ZN(n16499) );
  NOR2_X1 U18226 ( .A1(n16499), .A2(n17119), .ZN(n16332) );
  AOI211_X1 U18227 ( .C1(n18502), .C2(n17133), .A(n16333), .B(n16332), .ZN(
        n16334) );
  OAI21_X1 U18228 ( .B1(n16504), .B2(n17120), .A(n16334), .ZN(P2_U2990) );
  INV_X1 U18229 ( .A(n16347), .ZN(n16337) );
  INV_X1 U18230 ( .A(n16335), .ZN(n16336) );
  OAI21_X1 U18231 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16337), .A(
        n16336), .ZN(n16516) );
  OAI21_X1 U18232 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(n16514) );
  OAI22_X1 U18233 ( .A1(n17117), .A2(n13144), .B1(n17125), .B2(n18496), .ZN(
        n16342) );
  OAI22_X1 U18234 ( .A1(n17113), .A2(n18489), .B1(n17222), .B2(n14035), .ZN(
        n16341) );
  AOI211_X1 U18235 ( .C1(n16514), .C2(n17135), .A(n16342), .B(n16341), .ZN(
        n16343) );
  OAI21_X1 U18236 ( .B1(n17119), .B2(n16516), .A(n16343), .ZN(P2_U2991) );
  INV_X1 U18237 ( .A(n16344), .ZN(n16346) );
  NOR2_X1 U18238 ( .A1(n16346), .A2(n16345), .ZN(n16348) );
  OAI21_X1 U18239 ( .B1(n16348), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16347), .ZN(n16527) );
  OAI21_X1 U18240 ( .B1(n16351), .B2(n16350), .A(n16349), .ZN(n16525) );
  INV_X1 U18241 ( .A(n16352), .ZN(n16522) );
  OAI22_X1 U18242 ( .A1(n14035), .A2(n13077), .B1(n17125), .B2(n16353), .ZN(
        n16354) );
  AOI21_X1 U18243 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17126), .A(
        n16354), .ZN(n16355) );
  OAI21_X1 U18244 ( .B1(n16522), .B2(n17113), .A(n16355), .ZN(n16356) );
  AOI21_X1 U18245 ( .B1(n16525), .B2(n17135), .A(n16356), .ZN(n16357) );
  OAI21_X1 U18246 ( .B1(n17119), .B2(n16527), .A(n16357), .ZN(P2_U2992) );
  INV_X1 U18247 ( .A(n16363), .ZN(n16362) );
  XNOR2_X1 U18248 ( .A(n16364), .B(n16362), .ZN(n16373) );
  AND2_X1 U18249 ( .A1(n16364), .A2(n16363), .ZN(n16365) );
  AOI21_X1 U18250 ( .B1(n16373), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16365), .ZN(n16368) );
  XOR2_X1 U18251 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n16366), .Z(
        n16367) );
  XNOR2_X1 U18252 ( .A(n16368), .B(n16367), .ZN(n16538) );
  XOR2_X1 U18253 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n16344), .Z(
        n16536) );
  NOR2_X1 U18254 ( .A1(n14035), .A2(n18474), .ZN(n16531) );
  NOR2_X1 U18255 ( .A1(n17125), .A2(n18483), .ZN(n16369) );
  AOI211_X1 U18256 ( .C1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17126), .A(
        n16531), .B(n16369), .ZN(n16370) );
  OAI21_X1 U18257 ( .B1(n18478), .B2(n17113), .A(n16370), .ZN(n16371) );
  AOI21_X1 U18258 ( .B1(n16536), .B2(n17131), .A(n16371), .ZN(n16372) );
  OAI21_X1 U18259 ( .B1(n16538), .B2(n17120), .A(n16372), .ZN(P2_U2993) );
  XNOR2_X1 U18260 ( .A(n11003), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16560) );
  INV_X1 U18261 ( .A(n16374), .ZN(n16375) );
  NOR2_X1 U18262 ( .A1(n17111), .A2(n16375), .ZN(n16401) );
  AOI21_X1 U18263 ( .B1(n16401), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16376) );
  NOR2_X1 U18264 ( .A1(n16376), .A2(n16344), .ZN(n16558) );
  NOR2_X1 U18265 ( .A1(n14035), .A2(n17221), .ZN(n16550) );
  NOR2_X1 U18266 ( .A1(n17125), .A2(n16377), .ZN(n16378) );
  AOI211_X1 U18267 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n17126), .A(
        n16550), .B(n16378), .ZN(n16379) );
  OAI21_X1 U18268 ( .B1(n17113), .B2(n16553), .A(n16379), .ZN(n16380) );
  AOI21_X1 U18269 ( .B1(n16558), .B2(n17131), .A(n16380), .ZN(n16381) );
  OAI21_X1 U18270 ( .B1(n16560), .B2(n17120), .A(n16381), .ZN(P2_U2994) );
  NAND2_X1 U18271 ( .A1(n16383), .A2(n16382), .ZN(n16386) );
  INV_X1 U18272 ( .A(n16392), .ZN(n16384) );
  AOI21_X1 U18273 ( .B1(n16394), .B2(n16391), .A(n16384), .ZN(n16385) );
  XOR2_X1 U18274 ( .A(n16386), .B(n16385), .Z(n16571) );
  XNOR2_X1 U18275 ( .A(n16401), .B(n16565), .ZN(n16569) );
  NOR2_X1 U18276 ( .A1(n14035), .A2(n17220), .ZN(n16563) );
  NOR2_X1 U18277 ( .A1(n17125), .A2(n18470), .ZN(n16387) );
  AOI211_X1 U18278 ( .C1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17126), .A(
        n16563), .B(n16387), .ZN(n16388) );
  OAI21_X1 U18279 ( .B1(n17113), .B2(n18466), .A(n16388), .ZN(n16389) );
  AOI21_X1 U18280 ( .B1(n16569), .B2(n17131), .A(n16389), .ZN(n16390) );
  OAI21_X1 U18281 ( .B1(n16571), .B2(n17120), .A(n16390), .ZN(P2_U2995) );
  NAND2_X1 U18282 ( .A1(n16392), .A2(n16391), .ZN(n16393) );
  XNOR2_X1 U18283 ( .A(n16394), .B(n16393), .ZN(n16581) );
  NAND2_X1 U18284 ( .A1(n17105), .A2(n16395), .ZN(n16397) );
  NAND2_X1 U18285 ( .A1(n16396), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16573) );
  OAI211_X1 U18286 ( .C1(n16398), .C2(n17117), .A(n16397), .B(n16573), .ZN(
        n16399) );
  AOI21_X1 U18287 ( .B1(n16572), .B2(n17133), .A(n16399), .ZN(n16404) );
  INV_X1 U18288 ( .A(n17111), .ZN(n16400) );
  INV_X1 U18289 ( .A(n16539), .ZN(n16543) );
  NAND2_X1 U18290 ( .A1(n16400), .A2(n16543), .ZN(n16413) );
  AOI21_X1 U18291 ( .B1(n16402), .B2(n16413), .A(n16401), .ZN(n16578) );
  NAND2_X1 U18292 ( .A1(n16578), .A2(n17131), .ZN(n16403) );
  OAI211_X1 U18293 ( .C1(n16581), .C2(n17120), .A(n16404), .B(n16403), .ZN(
        P2_U2996) );
  INV_X1 U18294 ( .A(n16405), .ZN(n16407) );
  NOR2_X1 U18295 ( .A1(n16407), .A2(n16406), .ZN(n16408) );
  XNOR2_X1 U18296 ( .A(n16409), .B(n16408), .ZN(n16598) );
  INV_X1 U18297 ( .A(n18442), .ZN(n16412) );
  NOR2_X1 U18298 ( .A1(n18439), .A2(n18381), .ZN(n16583) );
  INV_X1 U18299 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16410) );
  OAI22_X1 U18300 ( .A1(n16410), .A2(n17117), .B1(n17125), .B2(n18447), .ZN(
        n16411) );
  AOI211_X1 U18301 ( .C1(n16412), .C2(n17133), .A(n16583), .B(n16411), .ZN(
        n16416) );
  OAI211_X1 U18302 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16414), .A(
        n16413), .B(n17131), .ZN(n16415) );
  OAI211_X1 U18303 ( .C1(n16598), .C2(n17120), .A(n16416), .B(n16415), .ZN(
        P2_U2997) );
  OAI21_X1 U18304 ( .B1(n16651), .B2(n16630), .A(n16631), .ZN(n16417) );
  NAND2_X1 U18305 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18591) );
  OR2_X1 U18306 ( .A1(n16651), .A2(n18591), .ZN(n17110) );
  NAND2_X1 U18307 ( .A1(n16417), .A2(n17110), .ZN(n16637) );
  NAND2_X1 U18308 ( .A1(n16418), .A2(n16645), .ZN(n16422) );
  INV_X1 U18309 ( .A(n16419), .ZN(n16609) );
  NOR2_X1 U18310 ( .A1(n16609), .A2(n16420), .ZN(n16421) );
  XNOR2_X1 U18311 ( .A(n16422), .B(n16421), .ZN(n16634) );
  OAI22_X1 U18312 ( .A1(n13055), .A2(n18381), .B1(n17125), .B2(n18408), .ZN(
        n16426) );
  INV_X1 U18313 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16423) );
  OAI22_X1 U18314 ( .A1(n17113), .A2(n16424), .B1(n17117), .B2(n16423), .ZN(
        n16425) );
  AOI211_X1 U18315 ( .C1(n16634), .C2(n17135), .A(n16426), .B(n16425), .ZN(
        n16427) );
  OAI21_X1 U18316 ( .B1(n16637), .B2(n17119), .A(n16427), .ZN(P2_U3001) );
  XNOR2_X1 U18317 ( .A(n11008), .B(n16428), .ZN(n16713) );
  INV_X1 U18318 ( .A(n17073), .ZN(n16431) );
  NOR2_X1 U18319 ( .A1(n16431), .A2(n16430), .ZN(n16433) );
  XOR2_X1 U18320 ( .A(n16433), .B(n16432), .Z(n16711) );
  OAI22_X1 U18321 ( .A1(n18347), .A2(n14035), .B1(n17125), .B2(n18344), .ZN(
        n16435) );
  OAI22_X1 U18322 ( .A1(n17113), .A2(n18348), .B1(n17117), .B2(n11224), .ZN(
        n16434) );
  AOI211_X1 U18323 ( .C1(n16711), .C2(n17135), .A(n16435), .B(n16434), .ZN(
        n16436) );
  OAI21_X1 U18324 ( .B1(n17119), .B2(n16713), .A(n16436), .ZN(P2_U3007) );
  NOR2_X1 U18325 ( .A1(n16437), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16460) );
  NOR2_X1 U18326 ( .A1(n16465), .A2(n16460), .ZN(n16449) );
  OR2_X1 U18327 ( .A1(n16438), .A2(n16437), .ZN(n16451) );
  XNOR2_X1 U18328 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16440) );
  OAI21_X1 U18329 ( .B1(n16451), .B2(n16440), .A(n16439), .ZN(n16441) );
  OAI21_X1 U18330 ( .B1(n16449), .B2(n16443), .A(n16442), .ZN(n16444) );
  OAI21_X1 U18331 ( .B1(n16447), .B2(n16730), .A(n16446), .ZN(P2_U3017) );
  NOR2_X1 U18332 ( .A1(n16449), .A2(n16448), .ZN(n16456) );
  INV_X1 U18333 ( .A(n16450), .ZN(n18552) );
  NOR2_X1 U18334 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16451), .ZN(
        n16452) );
  OAI21_X1 U18335 ( .B1(n18549), .B2(n16733), .A(n16454), .ZN(n16455) );
  OAI21_X1 U18336 ( .B1(n16459), .B2(n16730), .A(n16458), .ZN(P2_U3018) );
  NOR2_X1 U18337 ( .A1(n18535), .A2(n16705), .ZN(n16464) );
  INV_X1 U18338 ( .A(n16460), .ZN(n16462) );
  OAI211_X1 U18339 ( .C1(n16733), .C2(n18546), .A(n16462), .B(n16461), .ZN(
        n16463) );
  AOI211_X1 U18340 ( .C1(n16465), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16464), .B(n16463), .ZN(n16469) );
  NAND3_X1 U18341 ( .A1(n16467), .A2(n18612), .A3(n16466), .ZN(n16468) );
  OAI211_X1 U18342 ( .C1(n16470), .C2(n16730), .A(n16469), .B(n16468), .ZN(
        P2_U3019) );
  INV_X1 U18343 ( .A(n16490), .ZN(n16480) );
  AOI21_X1 U18344 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16472) );
  NOR3_X1 U18345 ( .A1(n16472), .A2(n16471), .A3(n16483), .ZN(n16473) );
  AOI211_X1 U18346 ( .C1(n18611), .C2(n16475), .A(n16474), .B(n16473), .ZN(
        n16476) );
  OAI21_X1 U18347 ( .B1(n16733), .B2(n18525), .A(n16476), .ZN(n16479) );
  NOR2_X1 U18348 ( .A1(n16477), .A2(n18604), .ZN(n16478) );
  AOI211_X1 U18349 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16480), .A(
        n16479), .B(n16478), .ZN(n16481) );
  OAI21_X1 U18350 ( .B1(n16482), .B2(n16730), .A(n16481), .ZN(P2_U3020) );
  NOR3_X1 U18351 ( .A1(n16484), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16483), .ZN(n16485) );
  AOI211_X1 U18352 ( .C1(n18606), .C2(n18511), .A(n16486), .B(n16485), .ZN(
        n16488) );
  NAND2_X1 U18353 ( .A1(n18611), .A2(n18512), .ZN(n16487) );
  OAI211_X1 U18354 ( .C1(n16490), .C2(n16489), .A(n16488), .B(n16487), .ZN(
        n16491) );
  AOI21_X1 U18355 ( .B1(n16492), .B2(n18612), .A(n16491), .ZN(n16493) );
  OAI21_X1 U18356 ( .B1(n16494), .B2(n16730), .A(n16493), .ZN(P2_U3021) );
  INV_X1 U18357 ( .A(n18501), .ZN(n16498) );
  AOI211_X1 U18358 ( .C1(n18611), .C2(n18502), .A(n16496), .B(n16495), .ZN(
        n16497) );
  OAI21_X1 U18359 ( .B1(n16733), .B2(n16498), .A(n16497), .ZN(n16501) );
  NOR2_X1 U18360 ( .A1(n16499), .A2(n18604), .ZN(n16500) );
  AOI211_X1 U18361 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16502), .A(
        n16501), .B(n16500), .ZN(n16503) );
  OAI21_X1 U18362 ( .B1(n16504), .B2(n16730), .A(n16503), .ZN(P2_U3022) );
  AOI21_X1 U18363 ( .B1(n16512), .B2(n16520), .A(n16505), .ZN(n16507) );
  NOR2_X1 U18364 ( .A1(n14035), .A2(n17222), .ZN(n16506) );
  AOI21_X1 U18365 ( .B1(n16507), .B2(n16517), .A(n16506), .ZN(n16508) );
  OAI21_X1 U18366 ( .B1(n16705), .B2(n18489), .A(n16508), .ZN(n16509) );
  AOI21_X1 U18367 ( .B1(n18606), .B2(n16510), .A(n16509), .ZN(n16511) );
  OAI21_X1 U18368 ( .B1(n16519), .B2(n16512), .A(n16511), .ZN(n16513) );
  AOI21_X1 U18369 ( .B1(n16514), .B2(n18609), .A(n16513), .ZN(n16515) );
  OAI21_X1 U18370 ( .B1(n18604), .B2(n16516), .A(n16515), .ZN(P2_U3023) );
  INV_X1 U18371 ( .A(n16517), .ZN(n16521) );
  NAND2_X1 U18372 ( .A1(n16396), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16518) );
  OAI221_X1 U18373 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16521), 
        .C1(n16520), .C2(n16519), .A(n16518), .ZN(n16524) );
  OAI22_X1 U18374 ( .A1(n16522), .A2(n16705), .B1(n16733), .B2(n19346), .ZN(
        n16523) );
  AOI211_X1 U18375 ( .C1(n16525), .C2(n18609), .A(n16524), .B(n16523), .ZN(
        n16526) );
  OAI21_X1 U18376 ( .B1(n18604), .B2(n16527), .A(n16526), .ZN(P2_U3024) );
  NAND2_X1 U18377 ( .A1(n16528), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16534) );
  NOR3_X1 U18378 ( .A1(n16529), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16549), .ZN(n16530) );
  AOI211_X1 U18379 ( .C1(n18606), .C2(n16532), .A(n16531), .B(n16530), .ZN(
        n16533) );
  OAI211_X1 U18380 ( .C1(n18478), .C2(n16705), .A(n16534), .B(n16533), .ZN(
        n16535) );
  AOI21_X1 U18381 ( .B1(n16536), .B2(n18612), .A(n16535), .ZN(n16537) );
  OAI21_X1 U18382 ( .B1(n16538), .B2(n16730), .A(n16537), .ZN(P2_U3025) );
  INV_X1 U18383 ( .A(n16627), .ZN(n16582) );
  NOR3_X1 U18384 ( .A1(n16582), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16539), .ZN(n16575) );
  NOR2_X1 U18385 ( .A1(n16586), .A2(n16540), .ZN(n16541) );
  NOR2_X1 U18386 ( .A1(n16542), .A2(n16541), .ZN(n16589) );
  NAND2_X1 U18387 ( .A1(n16590), .A2(n16543), .ZN(n16547) );
  NAND2_X1 U18388 ( .A1(n16545), .A2(n16544), .ZN(n16546) );
  NAND3_X1 U18389 ( .A1(n16740), .A2(n16547), .A3(n16546), .ZN(n16548) );
  NAND2_X1 U18390 ( .A1(n16589), .A2(n16548), .ZN(n16577) );
  NOR2_X1 U18391 ( .A1(n16575), .A2(n16577), .ZN(n16561) );
  INV_X1 U18392 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16556) );
  XNOR2_X1 U18393 ( .A(n16565), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16551) );
  INV_X1 U18394 ( .A(n16549), .ZN(n16564) );
  AOI21_X1 U18395 ( .B1(n16551), .B2(n16564), .A(n16550), .ZN(n16552) );
  OAI21_X1 U18396 ( .B1(n16553), .B2(n16705), .A(n16552), .ZN(n16554) );
  AOI21_X1 U18397 ( .B1(n18606), .B2(n19446), .A(n16554), .ZN(n16555) );
  OAI21_X1 U18398 ( .B1(n16561), .B2(n16556), .A(n16555), .ZN(n16557) );
  AOI21_X1 U18399 ( .B1(n16558), .B2(n18612), .A(n16557), .ZN(n16559) );
  OAI21_X1 U18400 ( .B1(n16560), .B2(n16730), .A(n16559), .ZN(P2_U3026) );
  NOR2_X1 U18401 ( .A1(n16561), .A2(n16565), .ZN(n16568) );
  NOR2_X1 U18402 ( .A1(n18466), .A2(n16705), .ZN(n16562) );
  AOI211_X1 U18403 ( .C1(n16565), .C2(n16564), .A(n16563), .B(n16562), .ZN(
        n16566) );
  OAI21_X1 U18404 ( .B1(n18465), .B2(n16733), .A(n16566), .ZN(n16567) );
  AOI211_X1 U18405 ( .C1(n16569), .C2(n18612), .A(n16568), .B(n16567), .ZN(
        n16570) );
  OAI21_X1 U18406 ( .B1(n16571), .B2(n16730), .A(n16570), .ZN(P2_U3027) );
  NAND2_X1 U18407 ( .A1(n16572), .A2(n18611), .ZN(n16574) );
  OAI211_X1 U18408 ( .C1(n16733), .C2(n18453), .A(n16574), .B(n16573), .ZN(
        n16576) );
  AOI211_X1 U18409 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16577), .A(
        n16576), .B(n16575), .ZN(n16580) );
  NAND2_X1 U18410 ( .A1(n16578), .A2(n18612), .ZN(n16579) );
  OAI211_X1 U18411 ( .C1(n16581), .C2(n16730), .A(n16580), .B(n16579), .ZN(
        P2_U3028) );
  AOI221_X1 U18412 ( .B1(n17111), .B2(n16582), .C1(n18604), .C2(n16582), .A(
        n16626), .ZN(n16600) );
  NAND3_X1 U18413 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16600), .A3(
        n16593), .ZN(n16585) );
  INV_X1 U18414 ( .A(n16583), .ZN(n16584) );
  OAI211_X1 U18415 ( .C1(n16705), .C2(n18442), .A(n16585), .B(n16584), .ZN(
        n16596) );
  NAND2_X1 U18416 ( .A1(n18604), .A2(n16586), .ZN(n16592) );
  NOR3_X1 U18417 ( .A1(n16588), .A2(n16626), .A3(n16587), .ZN(n16591) );
  OAI21_X1 U18418 ( .B1(n16591), .B2(n16590), .A(n16589), .ZN(n16616) );
  OAI21_X1 U18419 ( .B1(n16740), .B2(n18612), .A(n16607), .ZN(n16594) );
  AOI21_X1 U18420 ( .B1(n16608), .B2(n16594), .A(n16593), .ZN(n16595) );
  AOI211_X1 U18421 ( .C1(n18606), .C2(n18440), .A(n16596), .B(n16595), .ZN(
        n16597) );
  AOI21_X1 U18422 ( .B1(n16600), .B2(n16607), .A(n16599), .ZN(n16601) );
  NOR2_X1 U18423 ( .A1(n16603), .A2(n16730), .ZN(n16604) );
  AOI211_X1 U18424 ( .C1(n18606), .C2(n19618), .A(n16605), .B(n16604), .ZN(
        n16606) );
  OAI21_X1 U18425 ( .B1(n16608), .B2(n16607), .A(n16606), .ZN(P2_U3030) );
  NOR2_X1 U18426 ( .A1(n16610), .A2(n16609), .ZN(n17109) );
  INV_X1 U18427 ( .A(n17106), .ZN(n16611) );
  OAI21_X1 U18428 ( .B1(n17109), .B2(n16611), .A(n17107), .ZN(n16615) );
  NAND2_X1 U18429 ( .A1(n16613), .A2(n16612), .ZN(n16614) );
  XNOR2_X1 U18430 ( .A(n16615), .B(n16614), .ZN(n17121) );
  NAND2_X1 U18431 ( .A1(n16616), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16620) );
  INV_X1 U18432 ( .A(n18436), .ZN(n16618) );
  NOR2_X1 U18433 ( .A1(n13062), .A2(n18381), .ZN(n16617) );
  AOI21_X1 U18434 ( .B1(n18606), .B2(n16618), .A(n16617), .ZN(n16619) );
  OAI211_X1 U18435 ( .C1(n16705), .C2(n16621), .A(n16620), .B(n16619), .ZN(
        n16625) );
  NAND2_X1 U18436 ( .A1(n17111), .A2(n16626), .ZN(n16622) );
  NAND2_X1 U18437 ( .A1(n16623), .A2(n16622), .ZN(n17118) );
  NOR2_X1 U18438 ( .A1(n17118), .A2(n18604), .ZN(n16624) );
  AOI211_X1 U18439 ( .C1(n16627), .C2(n16626), .A(n16625), .B(n16624), .ZN(
        n16628) );
  OAI21_X1 U18440 ( .B1(n17121), .B2(n16730), .A(n16628), .ZN(P2_U3031) );
  OAI22_X1 U18441 ( .A1(n16733), .A2(n18402), .B1(n13055), .B2(n18381), .ZN(
        n16633) );
  NOR3_X1 U18442 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18592), .A3(
        n18590), .ZN(n16639) );
  OAI21_X1 U18443 ( .B1(n11148), .B2(n16751), .A(n16699), .ZN(n16640) );
  NOR2_X1 U18444 ( .A1(n16639), .A2(n16640), .ZN(n18595) );
  INV_X1 U18445 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16630) );
  NOR2_X1 U18446 ( .A1(n18592), .A2(n18590), .ZN(n16629) );
  NAND2_X1 U18447 ( .A1(n16629), .A2(n16631), .ZN(n18594) );
  OAI22_X1 U18448 ( .A1(n18595), .A2(n16631), .B1(n16630), .B2(n18594), .ZN(
        n16632) );
  AOI211_X1 U18449 ( .C1(n18403), .C2(n18611), .A(n16633), .B(n16632), .ZN(
        n16636) );
  NAND2_X1 U18450 ( .A1(n16634), .A2(n18609), .ZN(n16635) );
  OAI211_X1 U18451 ( .C1(n16637), .C2(n18604), .A(n16636), .B(n16635), .ZN(
        P2_U3033) );
  XNOR2_X1 U18452 ( .A(n16651), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17101) );
  NAND2_X1 U18453 ( .A1(n17101), .A2(n18612), .ZN(n16650) );
  NOR2_X1 U18454 ( .A1(n13048), .A2(n18381), .ZN(n16638) );
  AOI211_X1 U18455 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16640), .A(
        n16639), .B(n16638), .ZN(n16649) );
  XNOR2_X1 U18456 ( .A(n16642), .B(n16641), .ZN(n19124) );
  INV_X1 U18457 ( .A(n19124), .ZN(n16643) );
  AOI22_X1 U18458 ( .A1(n18611), .A2(n18389), .B1(n18606), .B2(n16643), .ZN(
        n16648) );
  NAND2_X1 U18459 ( .A1(n11404), .A2(n16645), .ZN(n16646) );
  XNOR2_X1 U18460 ( .A(n16644), .B(n16646), .ZN(n17102) );
  NAND2_X1 U18461 ( .A1(n17102), .A2(n18609), .ZN(n16647) );
  NAND4_X1 U18462 ( .A1(n16650), .A2(n16649), .A3(n16648), .A4(n16647), .ZN(
        P2_U3034) );
  OR2_X1 U18463 ( .A1(n14073), .A2(n16698), .ZN(n16686) );
  INV_X1 U18464 ( .A(n16673), .ZN(n16652) );
  OAI21_X1 U18465 ( .B1(n16652), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16651), .ZN(n17097) );
  OAI21_X1 U18466 ( .B1(n16653), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n17073), .ZN(n16656) );
  AOI21_X1 U18467 ( .B1(n16653), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n16654), .ZN(n16655) );
  NOR2_X1 U18468 ( .A1(n16656), .A2(n16655), .ZN(n16688) );
  NAND2_X1 U18469 ( .A1(n16688), .A2(n16689), .ZN(n16674) );
  INV_X1 U18470 ( .A(n16674), .ZN(n16692) );
  AOI21_X1 U18471 ( .B1(n16692), .B2(n16675), .A(n16657), .ZN(n16662) );
  INV_X1 U18472 ( .A(n16658), .ZN(n16660) );
  NOR2_X1 U18473 ( .A1(n16660), .A2(n16659), .ZN(n16661) );
  XNOR2_X1 U18474 ( .A(n16662), .B(n16661), .ZN(n17095) );
  NOR4_X1 U18475 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n13775), .A3(
        n16698), .A4(n18590), .ZN(n16670) );
  OAI22_X1 U18476 ( .A1(n16733), .A2(n18370), .B1(n18381), .B2(n16663), .ZN(
        n16667) );
  INV_X1 U18477 ( .A(n16699), .ZN(n16664) );
  AOI21_X1 U18478 ( .B1(n16698), .B2(n16740), .A(n16664), .ZN(n16681) );
  INV_X1 U18479 ( .A(n18590), .ZN(n16693) );
  NAND3_X1 U18480 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16693), .A3(
        n13775), .ZN(n16680) );
  AOI21_X1 U18481 ( .B1(n16681), .B2(n16680), .A(n16665), .ZN(n16666) );
  AOI211_X1 U18482 ( .C1(n18611), .C2(n18367), .A(n16667), .B(n16666), .ZN(
        n16668) );
  INV_X1 U18483 ( .A(n16668), .ZN(n16669) );
  AOI211_X1 U18484 ( .C1(n17095), .C2(n18609), .A(n16670), .B(n16669), .ZN(
        n16671) );
  OAI21_X1 U18485 ( .B1(n18604), .B2(n17097), .A(n16671), .ZN(P2_U3035) );
  NAND2_X1 U18486 ( .A1(n16686), .A2(n13775), .ZN(n16672) );
  NAND2_X1 U18487 ( .A1(n16673), .A2(n16672), .ZN(n17090) );
  NAND2_X1 U18488 ( .A1(n16674), .A2(n16691), .ZN(n16678) );
  NAND2_X1 U18489 ( .A1(n16676), .A2(n16675), .ZN(n16677) );
  XNOR2_X1 U18490 ( .A(n16678), .B(n16677), .ZN(n17088) );
  NAND2_X1 U18491 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n16396), .ZN(n16679) );
  OAI211_X1 U18492 ( .C1(n16681), .C2(n13775), .A(n16680), .B(n16679), .ZN(
        n16684) );
  OAI22_X1 U18493 ( .A1(n16733), .A2(n19127), .B1(n16705), .B2(n16682), .ZN(
        n16683) );
  AOI211_X1 U18494 ( .C1(n17088), .C2(n18609), .A(n16684), .B(n16683), .ZN(
        n16685) );
  OAI21_X1 U18495 ( .B1(n18604), .B2(n17090), .A(n16685), .ZN(P2_U3036) );
  INV_X1 U18496 ( .A(n14073), .ZN(n16687) );
  OAI21_X1 U18497 ( .B1(n16687), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16686), .ZN(n17081) );
  AOI21_X1 U18498 ( .B1(n16689), .B2(n16691), .A(n16688), .ZN(n16690) );
  AOI21_X1 U18499 ( .B1(n16692), .B2(n16691), .A(n16690), .ZN(n17080) );
  NAND2_X1 U18500 ( .A1(n16693), .A2(n16698), .ZN(n16697) );
  NOR2_X1 U18501 ( .A1(n13042), .A2(n18381), .ZN(n16695) );
  NOR2_X1 U18502 ( .A1(n16733), .A2(n18366), .ZN(n16694) );
  AOI211_X1 U18503 ( .C1(n18361), .C2(n18611), .A(n16695), .B(n16694), .ZN(
        n16696) );
  OAI211_X1 U18504 ( .C1(n16699), .C2(n16698), .A(n16697), .B(n16696), .ZN(
        n16700) );
  AOI21_X1 U18505 ( .B1(n17080), .B2(n18609), .A(n16700), .ZN(n16701) );
  OAI21_X1 U18506 ( .B1(n18604), .B2(n17081), .A(n16701), .ZN(P2_U3037) );
  INV_X1 U18507 ( .A(n16702), .ZN(n16704) );
  OAI21_X1 U18508 ( .B1(n16751), .B2(n16704), .A(n16703), .ZN(n18607) );
  OAI22_X1 U18509 ( .A1(n16705), .A2(n18348), .B1(n18347), .B2(n14035), .ZN(
        n16706) );
  AOI21_X1 U18510 ( .B1(n18607), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16706), .ZN(n16709) );
  NAND2_X1 U18511 ( .A1(n18615), .A2(n16707), .ZN(n16708) );
  OAI211_X1 U18512 ( .C1(n18349), .C2(n16733), .A(n16709), .B(n16708), .ZN(
        n16710) );
  AOI21_X1 U18513 ( .B1(n16711), .B2(n18609), .A(n16710), .ZN(n16712) );
  OAI21_X1 U18514 ( .B1(n16713), .B2(n18604), .A(n16712), .ZN(P2_U3039) );
  XNOR2_X1 U18515 ( .A(n16714), .B(n16719), .ZN(n17066) );
  INV_X1 U18516 ( .A(n17066), .ZN(n16729) );
  OR2_X1 U18517 ( .A1(n16716), .A2(n16715), .ZN(n16717) );
  AND2_X1 U18518 ( .A1(n16718), .A2(n16717), .ZN(n17065) );
  NAND2_X1 U18519 ( .A1(n16720), .A2(n16719), .ZN(n16724) );
  NOR2_X1 U18520 ( .A1(n18334), .A2(n18381), .ZN(n16721) );
  AOI21_X1 U18521 ( .B1(n18335), .B2(n18611), .A(n16721), .ZN(n16722) );
  OAI21_X1 U18522 ( .B1(n16724), .B2(n16723), .A(n16722), .ZN(n16725) );
  AOI21_X1 U18523 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18607), .A(
        n16725), .ZN(n16726) );
  OAI21_X1 U18524 ( .B1(n18337), .B2(n16733), .A(n16726), .ZN(n16727) );
  AOI21_X1 U18525 ( .B1(n17065), .B2(n18609), .A(n16727), .ZN(n16728) );
  OAI21_X1 U18526 ( .B1(n16729), .B2(n18604), .A(n16728), .ZN(P2_U3040) );
  OAI22_X1 U18527 ( .A1(n16733), .A2(n16732), .B1(n16731), .B2(n16730), .ZN(
        n16734) );
  AOI211_X1 U18528 ( .C1(n18611), .C2(n11028), .A(n16735), .B(n16734), .ZN(
        n16743) );
  INV_X1 U18529 ( .A(n16736), .ZN(n16737) );
  AOI22_X1 U18530 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16738), .B1(
        n18612), .B2(n16737), .ZN(n16742) );
  OAI211_X1 U18531 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16740), .B(n16739), .ZN(n16741) );
  NAND3_X1 U18532 ( .A1(n16743), .A2(n16742), .A3(n16741), .ZN(P2_U3045) );
  NOR2_X1 U18533 ( .A1(n18381), .A2(n17170), .ZN(n17129) );
  INV_X1 U18534 ( .A(n16744), .ZN(n16745) );
  OAI21_X1 U18535 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16746), .A(
        n16745), .ZN(n17128) );
  NOR2_X1 U18536 ( .A1(n18604), .A2(n17128), .ZN(n16747) );
  AOI211_X1 U18537 ( .C1(n16748), .C2(n18606), .A(n17129), .B(n16747), .ZN(
        n16754) );
  XNOR2_X1 U18538 ( .A(n16749), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17134) );
  AOI22_X1 U18539 ( .A1(n17132), .A2(n18611), .B1(n18609), .B2(n17134), .ZN(
        n16753) );
  MUX2_X1 U18540 ( .A(n16751), .B(n16750), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16752) );
  NAND3_X1 U18541 ( .A1(n16754), .A2(n16753), .A3(n16752), .ZN(P2_U3046) );
  INV_X1 U18542 ( .A(n16755), .ZN(n16757) );
  OAI222_X1 U18543 ( .A1(n16761), .A2(n19152), .B1(n18621), .B2(n16758), .C1(
        n16757), .C2(n16756), .ZN(n16759) );
  INV_X1 U18544 ( .A(n16762), .ZN(n16770) );
  MUX2_X1 U18545 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16759), .S(
        n16770), .Z(P2_U3600) );
  OAI22_X1 U18546 ( .A1(n19255), .A2(n16761), .B1(n16760), .B2(n18621), .ZN(
        n16763) );
  MUX2_X1 U18547 ( .A(n16763), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16762), .Z(P2_U3596) );
  INV_X1 U18548 ( .A(n16765), .ZN(n16766) );
  NOR4_X1 U18549 ( .A1(n16764), .A2(n16766), .A3(n12877), .A4(n18621), .ZN(
        n16767) );
  NAND2_X1 U18550 ( .A1(n16770), .A2(n16767), .ZN(n16768) );
  OAI21_X1 U18551 ( .B1(n16770), .B2(n16769), .A(n16768), .ZN(P2_U3595) );
  INV_X1 U18552 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16771) );
  INV_X1 U18553 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21756) );
  OAI21_X1 U18554 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21756), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18236) );
  NAND2_X1 U18555 ( .A1(n21765), .A2(n18236), .ZN(n16773) );
  INV_X1 U18556 ( .A(n21706), .ZN(n16772) );
  INV_X1 U18557 ( .A(BS16), .ZN(n17005) );
  NAND2_X1 U18558 ( .A1(n21767), .A2(n21756), .ZN(n21708) );
  AOI21_X1 U18559 ( .B1(n17005), .B2(n21708), .A(n16772), .ZN(n21702) );
  AOI21_X1 U18560 ( .B1(n16771), .B2(n16772), .A(n21702), .ZN(P3_U3280) );
  AND2_X1 U18561 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16772), .ZN(P3_U3028) );
  AND2_X1 U18562 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16772), .ZN(P3_U3027) );
  AND2_X1 U18563 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16772), .ZN(P3_U3026) );
  AND2_X1 U18564 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16772), .ZN(P3_U3025) );
  AND2_X1 U18565 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16772), .ZN(P3_U3024) );
  AND2_X1 U18566 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16772), .ZN(P3_U3023) );
  AND2_X1 U18567 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16772), .ZN(P3_U3022) );
  AND2_X1 U18568 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16772), .ZN(P3_U3021) );
  AND2_X1 U18569 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16772), .ZN(
        P3_U3020) );
  AND2_X1 U18570 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16772), .ZN(
        P3_U3019) );
  AND2_X1 U18571 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16772), .ZN(
        P3_U3018) );
  AND2_X1 U18572 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16772), .ZN(
        P3_U3017) );
  AND2_X1 U18573 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16772), .ZN(
        P3_U3016) );
  AND2_X1 U18574 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16773), .ZN(
        P3_U3015) );
  AND2_X1 U18575 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16773), .ZN(
        P3_U3014) );
  AND2_X1 U18576 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16773), .ZN(
        P3_U3013) );
  AND2_X1 U18577 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16773), .ZN(
        P3_U3012) );
  AND2_X1 U18578 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16773), .ZN(
        P3_U3011) );
  AND2_X1 U18579 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16773), .ZN(
        P3_U3010) );
  AND2_X1 U18580 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16773), .ZN(
        P3_U3009) );
  AND2_X1 U18581 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16773), .ZN(
        P3_U3008) );
  AND2_X1 U18582 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16773), .ZN(
        P3_U3007) );
  AND2_X1 U18583 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16773), .ZN(
        P3_U3006) );
  AND2_X1 U18584 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16773), .ZN(
        P3_U3005) );
  AND2_X1 U18585 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16773), .ZN(
        P3_U3004) );
  AND2_X1 U18586 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16772), .ZN(
        P3_U3003) );
  AND2_X1 U18587 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16772), .ZN(
        P3_U3002) );
  AND2_X1 U18588 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16772), .ZN(
        P3_U3001) );
  AND2_X1 U18589 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16772), .ZN(
        P3_U3000) );
  AND2_X1 U18590 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16773), .ZN(
        P3_U2999) );
  AOI21_X1 U18591 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16776)
         );
  NAND4_X1 U18592 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n21710), .A4(n21144), .ZN(n21260) );
  INV_X1 U18593 ( .A(n21260), .ZN(n16774) );
  AOI211_X1 U18594 ( .C1(n18128), .C2(n16776), .A(n16775), .B(n16774), .ZN(
        P3_U2998) );
  NAND2_X1 U18595 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17877), .ZN(n21265) );
  INV_X2 U18596 ( .A(n21265), .ZN(n18233) );
  NOR2_X4 U18597 ( .A1(n18233), .A2(n18217), .ZN(n18226) );
  AND2_X1 U18598 ( .A1(n18226), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NOR2_X1 U18599 ( .A1(n17765), .A2(n20116), .ZN(n16782) );
  INV_X1 U18600 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n16781) );
  NAND2_X1 U18601 ( .A1(n16780), .A2(n16779), .ZN(n20054) );
  AOI22_X1 U18602 ( .A1(n16782), .A2(n16781), .B1(n20116), .B2(n20054), .ZN(
        P3_U3298) );
  INV_X1 U18603 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18197) );
  NAND2_X1 U18604 ( .A1(n19016), .A2(n20116), .ZN(n20550) );
  INV_X1 U18605 ( .A(n20550), .ZN(n20171) );
  AOI21_X1 U18606 ( .B1(n16782), .B2(n18197), .A(n20171), .ZN(P3_U3299) );
  NOR2_X1 U18607 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21746), .ZN(n21742) );
  AOI21_X1 U18608 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21742), .A(n21749), 
        .ZN(n16784) );
  INV_X1 U18609 ( .A(n16784), .ZN(n21701) );
  INV_X1 U18610 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U18611 ( .A1(n21752), .A2(n21746), .ZN(n16783) );
  AOI21_X1 U18612 ( .B1(n17005), .B2(n16783), .A(n17178), .ZN(n21697) );
  AOI21_X1 U18613 ( .B1(n17178), .B2(n16799), .A(n21697), .ZN(P2_U3591) );
  AND2_X1 U18614 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17178), .ZN(P2_U3208) );
  AND2_X1 U18615 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n16784), .ZN(P2_U3207) );
  AND2_X1 U18616 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17178), .ZN(P2_U3206) );
  AND2_X1 U18617 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17178), .ZN(P2_U3205) );
  AND2_X1 U18618 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17178), .ZN(P2_U3204) );
  AND2_X1 U18619 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17178), .ZN(P2_U3203) );
  AND2_X1 U18620 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n16784), .ZN(P2_U3202) );
  AND2_X1 U18621 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n16784), .ZN(P2_U3201) );
  AND2_X1 U18622 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16784), .ZN(
        P2_U3200) );
  AND2_X1 U18623 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16784), .ZN(
        P2_U3199) );
  AND2_X1 U18624 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16784), .ZN(
        P2_U3198) );
  AND2_X1 U18625 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16784), .ZN(
        P2_U3197) );
  AND2_X1 U18626 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16784), .ZN(
        P2_U3196) );
  AND2_X1 U18627 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16784), .ZN(
        P2_U3195) );
  AND2_X1 U18628 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16784), .ZN(
        P2_U3194) );
  AND2_X1 U18629 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n16784), .ZN(
        P2_U3193) );
  AND2_X1 U18630 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n16784), .ZN(
        P2_U3192) );
  AND2_X1 U18631 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n16784), .ZN(
        P2_U3191) );
  AND2_X1 U18632 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17178), .ZN(
        P2_U3190) );
  AND2_X1 U18633 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17178), .ZN(
        P2_U3189) );
  AND2_X1 U18634 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17178), .ZN(
        P2_U3188) );
  AND2_X1 U18635 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17178), .ZN(
        P2_U3187) );
  AND2_X1 U18636 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n16784), .ZN(
        P2_U3186) );
  AND2_X1 U18637 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17178), .ZN(
        P2_U3185) );
  AND2_X1 U18638 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17178), .ZN(
        P2_U3184) );
  AND2_X1 U18639 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17178), .ZN(
        P2_U3183) );
  AND2_X1 U18640 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17178), .ZN(
        P2_U3182) );
  AND2_X1 U18641 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17178), .ZN(
        P2_U3181) );
  AND2_X1 U18642 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17178), .ZN(
        P2_U3180) );
  AND2_X1 U18643 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17178), .ZN(
        P2_U3179) );
  NAND2_X1 U18644 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n21735), .ZN(n18622) );
  AOI21_X1 U18645 ( .B1(n16785), .B2(n18286), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16786) );
  AOI221_X1 U18646 ( .B1(n18622), .B2(n16786), .C1(n14093), .C2(n16786), .A(
        n18631), .ZN(P2_U3178) );
  INV_X1 U18647 ( .A(n18632), .ZN(n16787) );
  OAI21_X1 U18648 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n18286), .ZN(n18636) );
  INV_X1 U18649 ( .A(n18636), .ZN(n18295) );
  AOI221_X1 U18650 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n18631), .C1(n16787), .C2(
        n18631), .A(n19313), .ZN(n17168) );
  INV_X1 U18651 ( .A(n17168), .ZN(n17166) );
  NOR2_X1 U18652 ( .A1(n16788), .A2(n17166), .ZN(P2_U3047) );
  AND2_X1 U18653 ( .A1(n17192), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18654 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16792) );
  NOR4_X1 U18655 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16791) );
  NOR4_X1 U18656 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16790) );
  NOR4_X1 U18657 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16789) );
  NAND4_X1 U18658 ( .A1(n16792), .A2(n16791), .A3(n16790), .A4(n16789), .ZN(
        n16798) );
  NOR4_X1 U18659 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16796) );
  AOI211_X1 U18660 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16795) );
  NOR4_X1 U18661 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16794) );
  NOR4_X1 U18662 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16793) );
  NAND4_X1 U18663 ( .A1(n16796), .A2(n16795), .A3(n16794), .A4(n16793), .ZN(
        n16797) );
  NOR2_X1 U18664 ( .A1(n16798), .A2(n16797), .ZN(n17176) );
  INV_X1 U18665 ( .A(n17176), .ZN(n17175) );
  NOR2_X1 U18666 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17175), .ZN(n17169) );
  INV_X1 U18667 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21700) );
  NAND3_X1 U18668 ( .A1(n17170), .A2(n21700), .A3(n16799), .ZN(n17174) );
  INV_X1 U18669 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U18670 ( .A1(n17169), .A2(n17174), .B1(n17175), .B2(n17234), .ZN(
        P2_U2821) );
  INV_X1 U18671 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U18672 ( .A1(n17169), .A2(n17170), .B1(n17175), .B2(n17232), .ZN(
        P2_U2820) );
  INV_X1 U18673 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21732) );
  OR2_X2 U18674 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21722), .ZN(n22337) );
  OAI21_X1 U18675 ( .B1(n21724), .B2(n21732), .A(n22337), .ZN(n16801) );
  INV_X1 U18676 ( .A(n16801), .ZN(n21696) );
  NOR2_X1 U18677 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21715) );
  OAI21_X1 U18678 ( .B1(BS16), .B2(n21715), .A(n21696), .ZN(n21694) );
  OAI21_X1 U18679 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21696), .A(n21694), 
        .ZN(n16800) );
  INV_X1 U18680 ( .A(n16800), .ZN(P1_U3464) );
  AND2_X1 U18681 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n16801), .ZN(P1_U3193) );
  AND2_X1 U18682 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n16802), .ZN(P1_U3192) );
  AND2_X1 U18683 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n16801), .ZN(P1_U3191) );
  AND2_X1 U18684 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n16802), .ZN(P1_U3190) );
  AND2_X1 U18685 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n16801), .ZN(P1_U3189) );
  AND2_X1 U18686 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n16802), .ZN(P1_U3188) );
  AND2_X1 U18687 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n16801), .ZN(P1_U3187) );
  AND2_X1 U18688 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n16801), .ZN(P1_U3186) );
  AND2_X1 U18689 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n16801), .ZN(
        P1_U3185) );
  AND2_X1 U18690 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n16801), .ZN(
        P1_U3184) );
  AND2_X1 U18691 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n16801), .ZN(
        P1_U3183) );
  AND2_X1 U18692 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n16802), .ZN(
        P1_U3182) );
  AND2_X1 U18693 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n16802), .ZN(
        P1_U3181) );
  AND2_X1 U18694 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n16802), .ZN(
        P1_U3180) );
  AND2_X1 U18695 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n16802), .ZN(
        P1_U3179) );
  AND2_X1 U18696 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n16802), .ZN(
        P1_U3178) );
  AND2_X1 U18697 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n16801), .ZN(
        P1_U3177) );
  AND2_X1 U18698 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n16801), .ZN(
        P1_U3176) );
  AND2_X1 U18699 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n16801), .ZN(
        P1_U3175) );
  AND2_X1 U18700 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n16801), .ZN(
        P1_U3174) );
  AND2_X1 U18701 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n16801), .ZN(
        P1_U3173) );
  AND2_X1 U18702 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n16801), .ZN(
        P1_U3172) );
  AND2_X1 U18703 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n16802), .ZN(
        P1_U3171) );
  AND2_X1 U18704 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n16802), .ZN(
        P1_U3170) );
  AND2_X1 U18705 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n16802), .ZN(
        P1_U3169) );
  AND2_X1 U18706 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n16802), .ZN(
        P1_U3168) );
  AND2_X1 U18707 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n16802), .ZN(
        P1_U3167) );
  AND2_X1 U18708 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n16802), .ZN(
        P1_U3166) );
  AND2_X1 U18709 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n16802), .ZN(
        P1_U3165) );
  AND2_X1 U18710 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n16802), .ZN(
        P1_U3164) );
  NOR3_X1 U18711 ( .A1(n16804), .A2(n16803), .A3(n21975), .ZN(n16809) );
  AOI211_X1 U18712 ( .C1(n16809), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16806), .B(n16805), .ZN(n16807) );
  INV_X1 U18713 ( .A(n16807), .ZN(n16808) );
  OAI21_X1 U18714 ( .B1(n16809), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16808), .ZN(n16811) );
  AOI222_X1 U18715 ( .A1(n21922), .A2(n16811), .B1(n21922), .B2(n16810), .C1(
        n16811), .C2(n16810), .ZN(n16814) );
  OR2_X1 U18716 ( .A1(n16814), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16813) );
  NAND2_X1 U18717 ( .A1(n16813), .A2(n16812), .ZN(n16816) );
  NAND2_X1 U18718 ( .A1(n16814), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16815) );
  NAND3_X1 U18719 ( .A1(n16816), .A2(n16815), .A3(n16841), .ZN(n16826) );
  NOR2_X1 U18720 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n16819) );
  OAI211_X1 U18721 ( .C1(n16820), .C2(n16819), .A(n16818), .B(n16817), .ZN(
        n16821) );
  OR2_X1 U18722 ( .A1(n16822), .A2(n16821), .ZN(n16823) );
  NOR2_X1 U18723 ( .A1(n16824), .A2(n16823), .ZN(n16825) );
  INV_X1 U18724 ( .A(n21693), .ZN(n16833) );
  OR2_X1 U18725 ( .A1(n16827), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16831) );
  OAI21_X1 U18726 ( .B1(n21716), .B2(n16829), .A(n16828), .ZN(n16830) );
  OAI21_X1 U18727 ( .B1(n16832), .B2(n16831), .A(n16830), .ZN(n16836) );
  AOI221_X1 U18728 ( .B1(n21683), .B2(n16839), .C1(n16833), .C2(n16839), .A(
        n16836), .ZN(n21685) );
  NOR2_X1 U18729 ( .A1(n21685), .A2(n21683), .ZN(n21684) );
  OAI211_X1 U18730 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21716), .A(n21684), 
        .B(n16834), .ZN(n21689) );
  NOR2_X1 U18731 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21683), .ZN(n21679) );
  AOI21_X1 U18732 ( .B1(n16835), .B2(n21679), .A(n16839), .ZN(n21678) );
  AND3_X1 U18733 ( .A1(n21678), .A2(n16837), .A3(n16836), .ZN(n16838) );
  AOI21_X1 U18734 ( .B1(n16839), .B2(n21689), .A(n16838), .ZN(P1_U3162) );
  NOR2_X1 U18735 ( .A1(n16841), .A2(n16840), .ZN(P1_U3032) );
  AND2_X1 U18736 ( .A1(n19808), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18737 ( .A1(n21724), .A2(n21732), .ZN(n16843) );
  INV_X1 U18738 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n16842) );
  AOI21_X1 U18739 ( .B1(n16843), .B2(n16842), .A(n22339), .ZN(P1_U2802) );
  OAI22_X1 U18740 ( .A1(n19842), .A2(keyinput_62), .B1(keyinput_61), .B2(
        P1_REIP_REG_22__SCAN_IN), .ZN(n16844) );
  AOI221_X1 U18741 ( .B1(n19842), .B2(keyinput_62), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_61), .A(n16844), .ZN(n17038) );
  XNOR2_X1 U18742 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n16926)
         );
  OAI22_X1 U18743 ( .A1(n19857), .A2(keyinput_54), .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .ZN(n16845) );
  AOI221_X1 U18744 ( .B1(n19857), .B2(keyinput_54), .C1(keyinput_55), .C2(
        P1_REIP_REG_28__SCAN_IN), .A(n16845), .ZN(n16923) );
  INV_X1 U18745 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19888) );
  INV_X1 U18746 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21723) );
  AOI22_X1 U18747 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_46), .B1(n21723), 
        .B2(keyinput_43), .ZN(n16846) );
  OAI221_X1 U18748 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_46), .C1(n21723), 
        .C2(keyinput_43), .A(n16846), .ZN(n16849) );
  AOI22_X1 U18749 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_45), .B1(n21936), 
        .B2(keyinput_44), .ZN(n16847) );
  OAI221_X1 U18750 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .C1(n21936), 
        .C2(keyinput_44), .A(n16847), .ZN(n16848) );
  AOI211_X1 U18751 ( .C1(keyinput_47), .C2(P1_W_R_N_REG_SCAN_IN), .A(n16849), 
        .B(n16848), .ZN(n16850) );
  OAI21_X1 U18752 ( .B1(keyinput_47), .B2(P1_W_R_N_REG_SCAN_IN), .A(n16850), 
        .ZN(n16914) );
  INV_X1 U18753 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n19988) );
  INV_X1 U18754 ( .A(keyinput_42), .ZN(n16912) );
  INV_X1 U18755 ( .A(keyinput_41), .ZN(n16910) );
  INV_X1 U18756 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n16939) );
  OAI22_X1 U18757 ( .A1(n16939), .A2(keyinput_38), .B1(P1_ADS_N_REG_SCAN_IN), 
        .B2(keyinput_39), .ZN(n16851) );
  AOI221_X1 U18758 ( .B1(n16939), .B2(keyinput_38), .C1(keyinput_39), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n16851), .ZN(n16907) );
  INV_X1 U18759 ( .A(READY1), .ZN(n17001) );
  INV_X1 U18760 ( .A(NA), .ZN(n21768) );
  AOI22_X1 U18761 ( .A1(HOLD), .A2(keyinput_33), .B1(DATAI_0_), .B2(
        keyinput_32), .ZN(n16852) );
  OAI221_X1 U18762 ( .B1(HOLD), .B2(keyinput_33), .C1(DATAI_0_), .C2(
        keyinput_32), .A(n16852), .ZN(n16899) );
  OAI22_X1 U18763 ( .A1(n16854), .A2(keyinput_30), .B1(keyinput_29), .B2(
        DATAI_3_), .ZN(n16853) );
  AOI221_X1 U18764 ( .B1(n16854), .B2(keyinput_30), .C1(DATAI_3_), .C2(
        keyinput_29), .A(n16853), .ZN(n16896) );
  INV_X1 U18765 ( .A(keyinput_28), .ZN(n16894) );
  AOI22_X1 U18766 ( .A1(DATAI_8_), .A2(keyinput_24), .B1(n16856), .B2(
        keyinput_26), .ZN(n16855) );
  OAI221_X1 U18767 ( .B1(DATAI_8_), .B2(keyinput_24), .C1(n16856), .C2(
        keyinput_26), .A(n16855), .ZN(n16863) );
  INV_X1 U18768 ( .A(DATAI_12_), .ZN(n16979) );
  AOI22_X1 U18769 ( .A1(n16858), .A2(keyinput_23), .B1(n16979), .B2(
        keyinput_20), .ZN(n16857) );
  OAI221_X1 U18770 ( .B1(n16858), .B2(keyinput_23), .C1(n16979), .C2(
        keyinput_20), .A(n16857), .ZN(n16862) );
  XNOR2_X1 U18771 ( .A(DATAI_10_), .B(keyinput_22), .ZN(n16861) );
  INV_X1 U18772 ( .A(DATAI_11_), .ZN(n16983) );
  AOI22_X1 U18773 ( .A1(DATAI_7_), .A2(keyinput_25), .B1(n16983), .B2(
        keyinput_21), .ZN(n16859) );
  OAI221_X1 U18774 ( .B1(DATAI_7_), .B2(keyinput_25), .C1(n16983), .C2(
        keyinput_21), .A(n16859), .ZN(n16860) );
  NOR4_X1 U18775 ( .A1(n16863), .A2(n16862), .A3(n16861), .A4(n16860), .ZN(
        n16891) );
  INV_X1 U18776 ( .A(DATAI_15_), .ZN(n16971) );
  OAI22_X1 U18777 ( .A1(n16971), .A2(keyinput_17), .B1(keyinput_18), .B2(
        DATAI_14_), .ZN(n16864) );
  AOI221_X1 U18778 ( .B1(n16971), .B2(keyinput_17), .C1(DATAI_14_), .C2(
        keyinput_18), .A(n16864), .ZN(n16888) );
  OAI22_X1 U18779 ( .A1(n16964), .A2(keyinput_15), .B1(keyinput_13), .B2(
        DATAI_19_), .ZN(n16865) );
  AOI221_X1 U18780 ( .B1(n16964), .B2(keyinput_15), .C1(DATAI_19_), .C2(
        keyinput_13), .A(n16865), .ZN(n16886) );
  OAI22_X1 U18781 ( .A1(DATAI_18_), .A2(keyinput_14), .B1(DATAI_16_), .B2(
        keyinput_16), .ZN(n16866) );
  AOI221_X1 U18782 ( .B1(DATAI_18_), .B2(keyinput_14), .C1(keyinput_16), .C2(
        DATAI_16_), .A(n16866), .ZN(n16885) );
  OAI22_X1 U18783 ( .A1(n16868), .A2(keyinput_7), .B1(DATAI_26_), .B2(
        keyinput_6), .ZN(n16867) );
  AOI221_X1 U18784 ( .B1(n16868), .B2(keyinput_7), .C1(keyinput_6), .C2(
        DATAI_26_), .A(n16867), .ZN(n16876) );
  OAI22_X1 U18785 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .ZN(n16869) );
  AOI221_X1 U18786 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n16869), .ZN(n16874) );
  AOI22_X1 U18787 ( .A1(DATAI_29_), .A2(keyinput_3), .B1(DATAI_30_), .B2(
        keyinput_2), .ZN(n16870) );
  OAI221_X1 U18788 ( .B1(DATAI_29_), .B2(keyinput_3), .C1(DATAI_30_), .C2(
        keyinput_2), .A(n16870), .ZN(n16873) );
  OAI22_X1 U18789 ( .A1(n16951), .A2(keyinput_4), .B1(keyinput_5), .B2(
        DATAI_27_), .ZN(n16871) );
  AOI221_X1 U18790 ( .B1(n16951), .B2(keyinput_4), .C1(DATAI_27_), .C2(
        keyinput_5), .A(n16871), .ZN(n16872) );
  OAI21_X1 U18791 ( .B1(n16874), .B2(n16873), .A(n16872), .ZN(n16875) );
  OAI211_X1 U18792 ( .C1(n16946), .C2(keyinput_8), .A(n16876), .B(n16875), 
        .ZN(n16877) );
  AOI21_X1 U18793 ( .B1(n16946), .B2(keyinput_8), .A(n16877), .ZN(n16883) );
  AOI22_X1 U18794 ( .A1(n16960), .A2(keyinput_9), .B1(keyinput_10), .B2(n16961), .ZN(n16878) );
  OAI221_X1 U18795 ( .B1(n16960), .B2(keyinput_9), .C1(n16961), .C2(
        keyinput_10), .A(n16878), .ZN(n16882) );
  OAI22_X1 U18796 ( .A1(n16880), .A2(keyinput_12), .B1(keyinput_11), .B2(
        DATAI_21_), .ZN(n16879) );
  AOI221_X1 U18797 ( .B1(n16880), .B2(keyinput_12), .C1(DATAI_21_), .C2(
        keyinput_11), .A(n16879), .ZN(n16881) );
  OAI21_X1 U18798 ( .B1(n16883), .B2(n16882), .A(n16881), .ZN(n16884) );
  NAND3_X1 U18799 ( .A1(n16886), .A2(n16885), .A3(n16884), .ZN(n16887) );
  AOI22_X1 U18800 ( .A1(n16888), .A2(n16887), .B1(keyinput_19), .B2(DATAI_13_), 
        .ZN(n16889) );
  OAI21_X1 U18801 ( .B1(keyinput_19), .B2(DATAI_13_), .A(n16889), .ZN(n16890)
         );
  AOI22_X1 U18802 ( .A1(n16891), .A2(n16890), .B1(keyinput_27), .B2(DATAI_5_), 
        .ZN(n16892) );
  OAI21_X1 U18803 ( .B1(keyinput_27), .B2(DATAI_5_), .A(n16892), .ZN(n16893)
         );
  OAI221_X1 U18804 ( .B1(DATAI_4_), .B2(n16894), .C1(n16992), .C2(keyinput_28), 
        .A(n16893), .ZN(n16895) );
  OAI211_X1 U18805 ( .C1(DATAI_1_), .C2(keyinput_31), .A(n16896), .B(n16895), 
        .ZN(n16897) );
  AOI21_X1 U18806 ( .B1(DATAI_1_), .B2(keyinput_31), .A(n16897), .ZN(n16898)
         );
  OAI22_X1 U18807 ( .A1(keyinput_34), .A2(n21768), .B1(n16899), .B2(n16898), 
        .ZN(n16900) );
  AOI21_X1 U18808 ( .B1(keyinput_34), .B2(n21768), .A(n16900), .ZN(n16904) );
  INV_X1 U18809 ( .A(READY2), .ZN(n16902) );
  AOI22_X1 U18810 ( .A1(BS16), .A2(keyinput_35), .B1(n16902), .B2(keyinput_37), 
        .ZN(n16901) );
  OAI221_X1 U18811 ( .B1(BS16), .B2(keyinput_35), .C1(n16902), .C2(keyinput_37), .A(n16901), .ZN(n16903) );
  AOI211_X1 U18812 ( .C1(n17001), .C2(keyinput_36), .A(n16904), .B(n16903), 
        .ZN(n16905) );
  OAI21_X1 U18813 ( .B1(n17001), .B2(keyinput_36), .A(n16905), .ZN(n16906) );
  OAI211_X1 U18814 ( .C1(P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_40), .A(
        n16907), .B(n16906), .ZN(n16908) );
  AOI21_X1 U18815 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_40), .A(n16908), .ZN(n16909) );
  AOI221_X1 U18816 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(n16910), .C1(n22338), 
        .C2(keyinput_41), .A(n16909), .ZN(n16911) );
  AOI221_X1 U18817 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .C1(n19988), 
        .C2(n16912), .A(n16911), .ZN(n16913) );
  OAI22_X1 U18818 ( .A1(keyinput_48), .A2(n19888), .B1(n16914), .B2(n16913), 
        .ZN(n16915) );
  AOI21_X1 U18819 ( .B1(keyinput_48), .B2(n19888), .A(n16915), .ZN(n16921) );
  INV_X1 U18820 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U18821 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_49), .B1(
        n19875), .B2(keyinput_50), .ZN(n16916) );
  OAI221_X1 U18822 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_49), .C1(
        n19875), .C2(keyinput_50), .A(n16916), .ZN(n16920) );
  XOR2_X1 U18823 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .Z(
        n16919) );
  OAI22_X1 U18824 ( .A1(n19861), .A2(keyinput_52), .B1(keyinput_53), .B2(
        P1_REIP_REG_30__SCAN_IN), .ZN(n16917) );
  AOI221_X1 U18825 ( .B1(n19861), .B2(keyinput_52), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_53), .A(n16917), .ZN(n16918) );
  OAI211_X1 U18826 ( .C1(n16921), .C2(n16920), .A(n16919), .B(n16918), .ZN(
        n16922) );
  AOI22_X1 U18827 ( .A1(n16923), .A2(n16922), .B1(keyinput_56), .B2(
        P1_REIP_REG_27__SCAN_IN), .ZN(n16924) );
  OAI21_X1 U18828 ( .B1(keyinput_56), .B2(P1_REIP_REG_27__SCAN_IN), .A(n16924), 
        .ZN(n16925) );
  AOI22_X1 U18829 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_58), .B1(n16926), .B2(n16925), .ZN(n16929) );
  AOI22_X1 U18830 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_60), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .ZN(n16927) );
  OAI221_X1 U18831 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_59), .A(n16927), .ZN(n16928) );
  AOI221_X1 U18832 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n16929), .C1(
        keyinput_58), .C2(n16929), .A(n16928), .ZN(n17037) );
  OAI22_X1 U18833 ( .A1(n21655), .A2(keyinput_123), .B1(n19846), .B2(
        keyinput_124), .ZN(n16930) );
  AOI221_X1 U18834 ( .B1(n21655), .B2(keyinput_123), .C1(keyinput_124), .C2(
        n19846), .A(n16930), .ZN(n17031) );
  OAI22_X1 U18835 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_126), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_125), .ZN(n16931) );
  AOI221_X1 U18836 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_126), .C1(
        keyinput_125), .C2(P1_REIP_REG_22__SCAN_IN), .A(n16931), .ZN(n17030)
         );
  INV_X1 U18837 ( .A(keyinput_122), .ZN(n17028) );
  INV_X1 U18838 ( .A(keyinput_121), .ZN(n17026) );
  OAI22_X1 U18839 ( .A1(n19857), .A2(keyinput_118), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_119), .ZN(n16932) );
  AOI221_X1 U18840 ( .B1(n19857), .B2(keyinput_118), .C1(keyinput_119), .C2(
        P1_REIP_REG_28__SCAN_IN), .A(n16932), .ZN(n17023) );
  AOI22_X1 U18841 ( .A1(keyinput_109), .A2(P1_MORE_REG_SCAN_IN), .B1(n21723), 
        .B2(keyinput_107), .ZN(n16933) );
  OAI221_X1 U18842 ( .B1(keyinput_109), .B2(P1_MORE_REG_SCAN_IN), .C1(n21723), 
        .C2(keyinput_107), .A(n16933), .ZN(n16936) );
  AOI22_X1 U18843 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_110), .B1(n20052), 
        .B2(keyinput_111), .ZN(n16934) );
  OAI221_X1 U18844 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_110), .C1(n20052), 
        .C2(keyinput_111), .A(n16934), .ZN(n16935) );
  AOI211_X1 U18845 ( .C1(keyinput_108), .C2(P1_STATEBS16_REG_SCAN_IN), .A(
        n16936), .B(n16935), .ZN(n16937) );
  OAI21_X1 U18846 ( .B1(keyinput_108), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        n16937), .ZN(n17014) );
  INV_X1 U18847 ( .A(keyinput_106), .ZN(n17012) );
  INV_X1 U18848 ( .A(keyinput_105), .ZN(n17010) );
  OAI22_X1 U18849 ( .A1(n16939), .A2(keyinput_102), .B1(P1_ADS_N_REG_SCAN_IN), 
        .B2(keyinput_103), .ZN(n16938) );
  AOI221_X1 U18850 ( .B1(n16939), .B2(keyinput_102), .C1(keyinput_103), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n16938), .ZN(n17007) );
  AOI22_X1 U18851 ( .A1(HOLD), .A2(keyinput_97), .B1(DATAI_0_), .B2(
        keyinput_96), .ZN(n16940) );
  OAI221_X1 U18852 ( .B1(HOLD), .B2(keyinput_97), .C1(DATAI_0_), .C2(
        keyinput_96), .A(n16940), .ZN(n16998) );
  OAI22_X1 U18853 ( .A1(DATAI_3_), .A2(keyinput_93), .B1(keyinput_95), .B2(
        DATAI_1_), .ZN(n16941) );
  AOI221_X1 U18854 ( .B1(DATAI_3_), .B2(keyinput_93), .C1(DATAI_1_), .C2(
        keyinput_95), .A(n16941), .ZN(n16995) );
  INV_X1 U18855 ( .A(keyinput_92), .ZN(n16993) );
  INV_X1 U18856 ( .A(keyinput_91), .ZN(n16989) );
  XNOR2_X1 U18857 ( .A(DATAI_13_), .B(keyinput_83), .ZN(n16987) );
  OAI22_X1 U18858 ( .A1(n16944), .A2(keyinput_77), .B1(n16943), .B2(
        keyinput_80), .ZN(n16942) );
  AOI221_X1 U18859 ( .B1(n16944), .B2(keyinput_77), .C1(keyinput_80), .C2(
        n16943), .A(n16942), .ZN(n16974) );
  OAI22_X1 U18860 ( .A1(n16946), .A2(keyinput_72), .B1(DATAI_25_), .B2(
        keyinput_71), .ZN(n16945) );
  AOI221_X1 U18861 ( .B1(n16946), .B2(keyinput_72), .C1(keyinput_71), .C2(
        DATAI_25_), .A(n16945), .ZN(n16956) );
  OAI22_X1 U18862 ( .A1(DATAI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n16947) );
  AOI221_X1 U18863 ( .B1(DATAI_31_), .B2(keyinput_65), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_64), .A(n16947), .ZN(n16954)
         );
  AOI22_X1 U18864 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(n16949), .B2(
        keyinput_66), .ZN(n16948) );
  OAI221_X1 U18865 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(n16949), .C2(
        keyinput_66), .A(n16948), .ZN(n16953) );
  OAI22_X1 U18866 ( .A1(n16951), .A2(keyinput_68), .B1(DATAI_27_), .B2(
        keyinput_69), .ZN(n16950) );
  AOI221_X1 U18867 ( .B1(n16951), .B2(keyinput_68), .C1(keyinput_69), .C2(
        DATAI_27_), .A(n16950), .ZN(n16952) );
  OAI21_X1 U18868 ( .B1(n16954), .B2(n16953), .A(n16952), .ZN(n16955) );
  OAI211_X1 U18869 ( .C1(DATAI_26_), .C2(keyinput_70), .A(n16956), .B(n16955), 
        .ZN(n16957) );
  AOI21_X1 U18870 ( .B1(DATAI_26_), .B2(keyinput_70), .A(n16957), .ZN(n16968)
         );
  OAI22_X1 U18871 ( .A1(DATAI_21_), .A2(keyinput_75), .B1(DATAI_20_), .B2(
        keyinput_76), .ZN(n16958) );
  AOI221_X1 U18872 ( .B1(DATAI_21_), .B2(keyinput_75), .C1(keyinput_76), .C2(
        DATAI_20_), .A(n16958), .ZN(n16967) );
  AOI22_X1 U18873 ( .A1(n16961), .A2(keyinput_74), .B1(n16960), .B2(
        keyinput_73), .ZN(n16959) );
  OAI221_X1 U18874 ( .B1(n16961), .B2(keyinput_74), .C1(n16960), .C2(
        keyinput_73), .A(n16959), .ZN(n16966) );
  AOI22_X1 U18875 ( .A1(n16964), .A2(keyinput_79), .B1(n16963), .B2(
        keyinput_78), .ZN(n16962) );
  OAI221_X1 U18876 ( .B1(n16964), .B2(keyinput_79), .C1(n16963), .C2(
        keyinput_78), .A(n16962), .ZN(n16965) );
  AOI221_X1 U18877 ( .B1(n16968), .B2(n16967), .C1(n16966), .C2(n16967), .A(
        n16965), .ZN(n16973) );
  INV_X1 U18878 ( .A(DATAI_14_), .ZN(n16970) );
  AOI22_X1 U18879 ( .A1(n16971), .A2(keyinput_81), .B1(n16970), .B2(
        keyinput_82), .ZN(n16969) );
  OAI221_X1 U18880 ( .B1(n16971), .B2(keyinput_81), .C1(n16970), .C2(
        keyinput_82), .A(n16969), .ZN(n16972) );
  AOI21_X1 U18881 ( .B1(n16974), .B2(n16973), .A(n16972), .ZN(n16986) );
  OAI22_X1 U18882 ( .A1(DATAI_9_), .A2(keyinput_87), .B1(DATAI_6_), .B2(
        keyinput_90), .ZN(n16975) );
  AOI221_X1 U18883 ( .B1(DATAI_9_), .B2(keyinput_87), .C1(keyinput_90), .C2(
        DATAI_6_), .A(n16975), .ZN(n16985) );
  OAI22_X1 U18884 ( .A1(DATAI_10_), .A2(keyinput_86), .B1(DATAI_7_), .B2(
        keyinput_89), .ZN(n16976) );
  AOI221_X1 U18885 ( .B1(DATAI_10_), .B2(keyinput_86), .C1(keyinput_89), .C2(
        DATAI_7_), .A(n16976), .ZN(n16981) );
  OAI22_X1 U18886 ( .A1(n16979), .A2(keyinput_84), .B1(n16978), .B2(
        keyinput_88), .ZN(n16977) );
  AOI221_X1 U18887 ( .B1(n16979), .B2(keyinput_84), .C1(keyinput_88), .C2(
        n16978), .A(n16977), .ZN(n16980) );
  OAI211_X1 U18888 ( .C1(n16983), .C2(keyinput_85), .A(n16981), .B(n16980), 
        .ZN(n16982) );
  AOI21_X1 U18889 ( .B1(n16983), .B2(keyinput_85), .A(n16982), .ZN(n16984) );
  OAI211_X1 U18890 ( .C1(n16987), .C2(n16986), .A(n16985), .B(n16984), .ZN(
        n16988) );
  OAI221_X1 U18891 ( .B1(DATAI_5_), .B2(keyinput_91), .C1(n16990), .C2(n16989), 
        .A(n16988), .ZN(n16991) );
  OAI221_X1 U18892 ( .B1(DATAI_4_), .B2(n16993), .C1(n16992), .C2(keyinput_92), 
        .A(n16991), .ZN(n16994) );
  OAI211_X1 U18893 ( .C1(DATAI_2_), .C2(keyinput_94), .A(n16995), .B(n16994), 
        .ZN(n16996) );
  AOI21_X1 U18894 ( .B1(DATAI_2_), .B2(keyinput_94), .A(n16996), .ZN(n16997)
         );
  OAI22_X1 U18895 ( .A1(keyinput_98), .A2(n21768), .B1(n16998), .B2(n16997), 
        .ZN(n16999) );
  AOI21_X1 U18896 ( .B1(keyinput_98), .B2(n21768), .A(n16999), .ZN(n17003) );
  AOI22_X1 U18897 ( .A1(READY2), .A2(keyinput_101), .B1(n17001), .B2(
        keyinput_100), .ZN(n17000) );
  OAI221_X1 U18898 ( .B1(READY2), .B2(keyinput_101), .C1(n17001), .C2(
        keyinput_100), .A(n17000), .ZN(n17002) );
  AOI211_X1 U18899 ( .C1(n17005), .C2(keyinput_99), .A(n17003), .B(n17002), 
        .ZN(n17004) );
  OAI21_X1 U18900 ( .B1(n17005), .B2(keyinput_99), .A(n17004), .ZN(n17006) );
  OAI211_X1 U18901 ( .C1(P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_104), .A(
        n17007), .B(n17006), .ZN(n17008) );
  AOI21_X1 U18902 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_104), .A(
        n17008), .ZN(n17009) );
  AOI221_X1 U18903 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(n17010), .C1(n22338), 
        .C2(keyinput_105), .A(n17009), .ZN(n17011) );
  AOI221_X1 U18904 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n17012), .C1(n19988), .C2(
        keyinput_106), .A(n17011), .ZN(n17013) );
  OAI22_X1 U18905 ( .A1(keyinput_112), .A2(n19888), .B1(n17014), .B2(n17013), 
        .ZN(n17015) );
  AOI21_X1 U18906 ( .B1(keyinput_112), .B2(n19888), .A(n17015), .ZN(n17021) );
  INV_X1 U18907 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U18908 ( .A1(n19875), .A2(keyinput_114), .B1(keyinput_113), .B2(
        n19883), .ZN(n17016) );
  OAI221_X1 U18909 ( .B1(n19875), .B2(keyinput_114), .C1(n19883), .C2(
        keyinput_113), .A(n17016), .ZN(n17020) );
  OAI22_X1 U18910 ( .A1(n19861), .A2(keyinput_116), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_117), .ZN(n17017) );
  AOI221_X1 U18911 ( .B1(n19861), .B2(keyinput_116), .C1(keyinput_117), .C2(
        P1_REIP_REG_30__SCAN_IN), .A(n17017), .ZN(n17019) );
  XNOR2_X1 U18912 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_115), .ZN(
        n17018) );
  OAI211_X1 U18913 ( .C1(n17021), .C2(n17020), .A(n17019), .B(n17018), .ZN(
        n17022) );
  AOI22_X1 U18914 ( .A1(keyinput_120), .A2(n19851), .B1(n17023), .B2(n17022), 
        .ZN(n17024) );
  OAI21_X1 U18915 ( .B1(n19851), .B2(keyinput_120), .A(n17024), .ZN(n17025) );
  OAI221_X1 U18916 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n17026), .C1(n15543), 
        .C2(keyinput_121), .A(n17025), .ZN(n17027) );
  OAI221_X1 U18917 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n17028), .C1(n19849), 
        .C2(keyinput_122), .A(n17027), .ZN(n17029) );
  NAND3_X1 U18918 ( .A1(n17031), .A2(n17030), .A3(n17029), .ZN(n17033) );
  AOI21_X1 U18919 ( .B1(keyinput_127), .B2(n17033), .A(P1_REIP_REG_20__SCAN_IN), .ZN(n17035) );
  INV_X1 U18920 ( .A(keyinput_127), .ZN(n17032) );
  AOI21_X1 U18921 ( .B1(n17033), .B2(n17032), .A(keyinput_63), .ZN(n17034) );
  AOI22_X1 U18922 ( .A1(keyinput_63), .A2(n17035), .B1(P1_REIP_REG_20__SCAN_IN), .B2(n17034), .ZN(n17036) );
  AOI21_X1 U18923 ( .B1(n17038), .B2(n17037), .A(n17036), .ZN(n17053) );
  NOR3_X4 U18924 ( .A1(n17039), .A2(n21698), .A3(n19325), .ZN(n19631) );
  NOR3_X4 U18925 ( .A1(n21698), .A2(n14182), .A3(n19325), .ZN(n19632) );
  AOI22_X1 U18926 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19632), .ZN(n19521) );
  INV_X1 U18927 ( .A(n19289), .ZN(n19142) );
  NOR2_X1 U18928 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17156), .ZN(
        n19243) );
  INV_X1 U18929 ( .A(n19243), .ZN(n19240) );
  NOR2_X1 U18930 ( .A1(n19288), .A2(n19240), .ZN(n19685) );
  OAI21_X1 U18931 ( .B1(n17040), .B2(n19685), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17041) );
  OAI21_X1 U18932 ( .B1(n19142), .B2(n19240), .A(n17041), .ZN(n19686) );
  NOR2_X2 U18933 ( .A1(n17042), .A2(n19625), .ZN(n19527) );
  NOR2_X2 U18934 ( .A1(n12433), .A2(n19627), .ZN(n19525) );
  AOI22_X1 U18935 ( .A1(n19686), .A2(n19527), .B1(n19525), .B2(n19685), .ZN(
        n17051) );
  AOI22_X1 U18936 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19631), .ZN(n19524) );
  NOR2_X2 U18937 ( .A1(n17160), .A2(n19282), .ZN(n19688) );
  NAND2_X1 U18938 ( .A1(n19160), .A2(n19316), .ZN(n19187) );
  OR2_X1 U18939 ( .A1(n21698), .A2(n19187), .ZN(n19292) );
  INV_X1 U18940 ( .A(n17044), .ZN(n19162) );
  OAI22_X1 U18941 ( .A1(n17160), .A2(n19292), .B1(n19162), .B2(n19240), .ZN(
        n17049) );
  AND2_X1 U18942 ( .A1(n17045), .A2(n19293), .ZN(n19329) );
  INV_X1 U18943 ( .A(n19329), .ZN(n19262) );
  INV_X1 U18944 ( .A(n19685), .ZN(n17046) );
  OAI211_X1 U18945 ( .C1(n17047), .C2(n19262), .A(n17046), .B(n19307), .ZN(
        n17048) );
  NAND3_X1 U18946 ( .A1(n17049), .A2(n17048), .A3(n19313), .ZN(n19687) );
  AOI22_X1 U18947 ( .A1(n19528), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17050) );
  OAI211_X1 U18948 ( .C1(n19521), .C2(n19696), .A(n17051), .B(n17050), .ZN(
        n17052) );
  XOR2_X1 U18949 ( .A(n17053), .B(n17052), .Z(P2_U3099) );
  INV_X1 U18950 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17054) );
  OAI22_X1 U18951 ( .A1(n18286), .A2(n17056), .B1(n17055), .B2(n17054), .ZN(
        P2_U2816) );
  AOI22_X1 U18952 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n18312), .ZN(n17063) );
  NAND3_X1 U18953 ( .A1(n17057), .A2(n17135), .A3(n15072), .ZN(n17060) );
  NAND2_X1 U18954 ( .A1(n17058), .A2(n17131), .ZN(n17059) );
  OAI211_X1 U18955 ( .C1(n17113), .C2(n18306), .A(n17060), .B(n17059), .ZN(
        n17061) );
  INV_X1 U18956 ( .A(n17061), .ZN(n17062) );
  OAI211_X1 U18957 ( .C1(n17064), .C2(n17117), .A(n17063), .B(n17062), .ZN(
        P2_U3010) );
  AOI22_X1 U18958 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n18329), .ZN(n17068) );
  AOI222_X1 U18959 ( .A1(n17066), .A2(n17131), .B1(n17133), .B2(n18335), .C1(
        n17135), .C2(n17065), .ZN(n17067) );
  OAI211_X1 U18960 ( .C1(n17069), .C2(n17117), .A(n17068), .B(n17067), .ZN(
        P2_U3008) );
  AOI22_X1 U18961 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n17070), .ZN(n17078) );
  XOR2_X1 U18962 ( .A(n17072), .B(n17071), .Z(n18613) );
  NAND2_X1 U18963 ( .A1(n16653), .A2(n17073), .ZN(n17076) );
  XNOR2_X1 U18964 ( .A(n17074), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17075) );
  XNOR2_X1 U18965 ( .A(n17076), .B(n17075), .ZN(n18608) );
  AOI222_X1 U18966 ( .A1(n18613), .A2(n17131), .B1(n17133), .B2(n18610), .C1(
        n17135), .C2(n18608), .ZN(n17077) );
  OAI211_X1 U18967 ( .C1(n17079), .C2(n17117), .A(n17078), .B(n17077), .ZN(
        P2_U3006) );
  AOI22_X1 U18968 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17126), .B1(
        P2_REIP_REG_9__SCAN_IN), .B2(n16396), .ZN(n17085) );
  INV_X1 U18969 ( .A(n17080), .ZN(n17082) );
  OAI22_X1 U18970 ( .A1(n17082), .A2(n17120), .B1(n17119), .B2(n17081), .ZN(
        n17083) );
  AOI21_X1 U18971 ( .B1(n17133), .B2(n18361), .A(n17083), .ZN(n17084) );
  OAI211_X1 U18972 ( .C1(n17125), .C2(n18359), .A(n17085), .B(n17084), .ZN(
        P2_U3005) );
  AOI22_X1 U18973 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n17086), .ZN(n17093) );
  AOI22_X1 U18974 ( .A1(n17088), .A2(n17135), .B1(n17133), .B2(n17087), .ZN(
        n17089) );
  OAI21_X1 U18975 ( .B1(n17090), .B2(n17119), .A(n17089), .ZN(n17091) );
  INV_X1 U18976 ( .A(n17091), .ZN(n17092) );
  OAI211_X1 U18977 ( .C1(n17094), .C2(n17117), .A(n17093), .B(n17092), .ZN(
        P2_U3004) );
  AOI22_X1 U18978 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17126), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n16396), .ZN(n17100) );
  INV_X1 U18979 ( .A(n17095), .ZN(n17096) );
  OAI22_X1 U18980 ( .A1(n17097), .A2(n17119), .B1(n17096), .B2(n17120), .ZN(
        n17098) );
  AOI21_X1 U18981 ( .B1(n17133), .B2(n18367), .A(n17098), .ZN(n17099) );
  OAI211_X1 U18982 ( .C1(n17125), .C2(n18380), .A(n17100), .B(n17099), .ZN(
        P2_U3003) );
  AOI22_X1 U18983 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n18388), .ZN(n17104) );
  AOI222_X1 U18984 ( .A1(n17102), .A2(n17135), .B1(n17133), .B2(n18389), .C1(
        n17131), .C2(n17101), .ZN(n17103) );
  OAI211_X1 U18985 ( .C1(n18382), .C2(n17117), .A(n17104), .B(n17103), .ZN(
        P2_U3002) );
  AOI22_X1 U18986 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n16396), .B1(n17105), 
        .B2(n18410), .ZN(n17116) );
  NAND2_X1 U18987 ( .A1(n17107), .A2(n17106), .ZN(n17108) );
  XNOR2_X1 U18988 ( .A(n17109), .B(n17108), .ZN(n18600) );
  NAND2_X1 U18989 ( .A1(n17110), .A2(n18596), .ZN(n17112) );
  NAND2_X1 U18990 ( .A1(n17112), .A2(n17111), .ZN(n18603) );
  OAI22_X1 U18991 ( .A1(n18603), .A2(n17119), .B1(n17113), .B2(n18417), .ZN(
        n17114) );
  AOI21_X1 U18992 ( .B1(n17135), .B2(n18600), .A(n17114), .ZN(n17115) );
  OAI211_X1 U18993 ( .C1(n18413), .C2(n17117), .A(n17116), .B(n17115), .ZN(
        P2_U3000) );
  AOI22_X1 U18994 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17126), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n16396), .ZN(n17124) );
  OAI22_X1 U18995 ( .A1(n17121), .A2(n17120), .B1(n17119), .B2(n17118), .ZN(
        n17122) );
  AOI21_X1 U18996 ( .B1(n17133), .B2(n18433), .A(n17122), .ZN(n17123) );
  OAI211_X1 U18997 ( .C1(n17125), .C2(n18430), .A(n17124), .B(n17123), .ZN(
        P2_U2999) );
  OAI21_X1 U18998 ( .B1(n17127), .B2(n17126), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17140) );
  INV_X1 U18999 ( .A(n17128), .ZN(n17130) );
  AOI21_X1 U19000 ( .B1(n17131), .B2(n17130), .A(n17129), .ZN(n17138) );
  NAND2_X1 U19001 ( .A1(n17133), .A2(n17132), .ZN(n17137) );
  NAND2_X1 U19002 ( .A1(n17135), .A2(n17134), .ZN(n17136) );
  AND3_X1 U19003 ( .A1(n17138), .A2(n17137), .A3(n17136), .ZN(n17139) );
  NAND2_X1 U19004 ( .A1(n17140), .A2(n17139), .ZN(P2_U3014) );
  INV_X1 U19005 ( .A(n17149), .ZN(n18289) );
  INV_X1 U19006 ( .A(n17141), .ZN(n17143) );
  OAI22_X1 U19007 ( .A1(n17144), .A2(n18289), .B1(n17143), .B2(n17142), .ZN(
        n17145) );
  AOI21_X1 U19008 ( .B1(n17147), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17145), 
        .ZN(n17146) );
  OAI22_X1 U19009 ( .A1(n17147), .A2(n17166), .B1(n17168), .B2(n17146), .ZN(
        P2_U3605) );
  OR2_X1 U19010 ( .A1(n19152), .A2(n21698), .ZN(n19133) );
  INV_X1 U19011 ( .A(n19133), .ZN(n17148) );
  NAND2_X1 U19012 ( .A1(n19254), .A2(n17148), .ZN(n19273) );
  NAND2_X1 U19013 ( .A1(n17148), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17150) );
  AND2_X1 U19014 ( .A1(n17150), .A2(n17149), .ZN(n17163) );
  NAND2_X1 U19015 ( .A1(n17163), .A2(n17161), .ZN(n17153) );
  NAND2_X1 U19016 ( .A1(n17151), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17152) );
  OAI211_X1 U19017 ( .C1(n19273), .C2(n19307), .A(n17153), .B(n17152), .ZN(
        n17154) );
  INV_X1 U19018 ( .A(n17154), .ZN(n17155) );
  AOI22_X1 U19019 ( .A1(n17168), .A2(n17156), .B1(n17155), .B2(n17166), .ZN(
        P2_U3603) );
  OAI21_X1 U19020 ( .B1(n21698), .B2(n19307), .A(n19152), .ZN(n17157) );
  AOI22_X1 U19021 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n17158), .B1(n17163), 
        .B2(n17157), .ZN(n17159) );
  AOI22_X1 U19022 ( .A1(n17168), .A2(n19302), .B1(n17159), .B2(n17166), .ZN(
        P2_U3604) );
  NOR2_X1 U19023 ( .A1(n17160), .A2(n19133), .ZN(n19234) );
  INV_X1 U19024 ( .A(n19234), .ZN(n17162) );
  NAND2_X1 U19025 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19206), .ZN(n19188) );
  NAND2_X1 U19026 ( .A1(n17162), .A2(n19188), .ZN(n17165) );
  INV_X1 U19027 ( .A(n19255), .ZN(n19274) );
  AOI222_X1 U19028 ( .A1(n17165), .A2(n19321), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n17164), .C1(n19274), .C2(n17163), .ZN(n17167) );
  AOI22_X1 U19029 ( .A1(n17168), .A2(n19175), .B1(n17167), .B2(n17166), .ZN(
        P2_U3602) );
  NAND2_X1 U19030 ( .A1(n17169), .A2(n21700), .ZN(n17173) );
  OAI21_X1 U19031 ( .B1(n12472), .B2(n17170), .A(n17176), .ZN(n17171) );
  OAI21_X1 U19032 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17176), .A(n17171), 
        .ZN(n17172) );
  OAI221_X1 U19033 ( .B1(n17173), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17173), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17172), .ZN(P2_U2822) );
  INV_X1 U19034 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17236) );
  OAI221_X1 U19035 ( .B1(n17176), .B2(n17236), .C1(n17175), .C2(n17174), .A(
        n17173), .ZN(P2_U2823) );
  MUX2_X1 U19036 ( .A(P2_M_IO_N_REG_SCAN_IN), .B(P2_MEMORYFETCH_REG_SCAN_IN), 
        .S(n17237), .Z(P2_U3611) );
  INV_X1 U19037 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17177) );
  AOI22_X1 U19038 ( .A1(n17237), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17177), 
        .B2(n21736), .ZN(P2_U3608) );
  INV_X1 U19039 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21755) );
  INV_X1 U19040 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17179) );
  OAI21_X1 U19041 ( .B1(n21755), .B2(n17179), .A(n17178), .ZN(P2_U2815) );
  AOI22_X1 U19042 ( .A1(n17211), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17181) );
  OAI21_X1 U19043 ( .B1(n12946), .B2(n17213), .A(n17181), .ZN(P2_U2951) );
  INV_X1 U19044 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U19045 ( .A1(n17211), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17182) );
  OAI21_X1 U19046 ( .B1(n17183), .B2(n17213), .A(n17182), .ZN(P2_U2950) );
  INV_X1 U19047 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U19048 ( .A1(n17211), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U19049 ( .B1(n17185), .B2(n17213), .A(n17184), .ZN(P2_U2949) );
  INV_X1 U19050 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U19051 ( .A1(n17200), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U19052 ( .B1(n17187), .B2(n17213), .A(n17186), .ZN(P2_U2948) );
  INV_X1 U19053 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U19054 ( .A1(n17211), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U19055 ( .B1(n17189), .B2(n17213), .A(n17188), .ZN(P2_U2947) );
  INV_X1 U19056 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U19057 ( .A1(n17200), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17190) );
  OAI21_X1 U19058 ( .B1(n17191), .B2(n17213), .A(n17190), .ZN(P2_U2946) );
  AOI22_X1 U19059 ( .A1(n17200), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17193) );
  OAI21_X1 U19060 ( .B1(n17194), .B2(n17213), .A(n17193), .ZN(P2_U2945) );
  AOI22_X1 U19061 ( .A1(n17200), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U19062 ( .B1(n17196), .B2(n17213), .A(n17195), .ZN(P2_U2944) );
  AOI22_X1 U19063 ( .A1(n17200), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17197) );
  OAI21_X1 U19064 ( .B1(n12924), .B2(n17213), .A(n17197), .ZN(P2_U2943) );
  AOI22_X1 U19065 ( .A1(n17211), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17198) );
  OAI21_X1 U19066 ( .B1(n17199), .B2(n17213), .A(n17198), .ZN(P2_U2942) );
  AOI22_X1 U19067 ( .A1(n17200), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17201) );
  OAI21_X1 U19068 ( .B1(n17202), .B2(n17213), .A(n17201), .ZN(P2_U2941) );
  AOI22_X1 U19069 ( .A1(n17211), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17203) );
  OAI21_X1 U19070 ( .B1(n17204), .B2(n17213), .A(n17203), .ZN(P2_U2940) );
  AOI22_X1 U19071 ( .A1(n17211), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U19072 ( .B1(n17206), .B2(n17213), .A(n17205), .ZN(P2_U2939) );
  AOI22_X1 U19073 ( .A1(n17211), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17207) );
  OAI21_X1 U19074 ( .B1(n17208), .B2(n17213), .A(n17207), .ZN(P2_U2938) );
  AOI22_X1 U19075 ( .A1(n17211), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17209) );
  OAI21_X1 U19076 ( .B1(n17210), .B2(n17213), .A(n17209), .ZN(P2_U2937) );
  AOI22_X1 U19077 ( .A1(n17211), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17192), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17212) );
  OAI21_X1 U19078 ( .B1(n17214), .B2(n17213), .A(n17212), .ZN(P2_U2936) );
  AOI21_X1 U19079 ( .B1(n21755), .B2(n17215), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17216) );
  AOI21_X1 U19080 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17237), .A(n17216), 
        .ZN(P2_U2817) );
  NOR2_X1 U19081 ( .A1(n21752), .A2(n21736), .ZN(n21739) );
  OAI222_X1 U19082 ( .A1(n17230), .A2(n17217), .B1(n19738), .B2(n17237), .C1(
        n12472), .C2(n17226), .ZN(P2_U3212) );
  INV_X1 U19083 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19740) );
  OAI222_X1 U19084 ( .A1(n17230), .A2(n17218), .B1(n19740), .B2(n17237), .C1(
        n17217), .C2(n17226), .ZN(P2_U3213) );
  INV_X1 U19085 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19742) );
  OAI222_X1 U19086 ( .A1(n17230), .A2(n12989), .B1(n19742), .B2(n17237), .C1(
        n17218), .C2(n17226), .ZN(P2_U3214) );
  INV_X1 U19087 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19744) );
  OAI222_X1 U19088 ( .A1(n17230), .A2(n15177), .B1(n19744), .B2(n17237), .C1(
        n12989), .C2(n17226), .ZN(P2_U3215) );
  INV_X1 U19089 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19746) );
  OAI222_X1 U19090 ( .A1(n17230), .A2(n18334), .B1(n19746), .B2(n17237), .C1(
        n15177), .C2(n17226), .ZN(P2_U3216) );
  INV_X1 U19091 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19748) );
  OAI222_X1 U19092 ( .A1(n17230), .A2(n18347), .B1(n19748), .B2(n17237), .C1(
        n18334), .C2(n17226), .ZN(P2_U3217) );
  INV_X1 U19093 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17219) );
  INV_X1 U19094 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19750) );
  OAI222_X1 U19095 ( .A1(n17230), .A2(n17219), .B1(n19750), .B2(n17237), .C1(
        n18347), .C2(n17226), .ZN(P2_U3218) );
  INV_X1 U19096 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19752) );
  OAI222_X1 U19097 ( .A1(n17230), .A2(n13042), .B1(n19752), .B2(n17237), .C1(
        n17219), .C2(n17226), .ZN(P2_U3219) );
  INV_X1 U19098 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19754) );
  OAI222_X1 U19099 ( .A1(n17226), .A2(n13042), .B1(n19754), .B2(n17237), .C1(
        n15038), .C2(n17230), .ZN(P2_U3220) );
  INV_X1 U19100 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19756) );
  OAI222_X1 U19101 ( .A1(n17226), .A2(n15038), .B1(n19756), .B2(n17237), .C1(
        n16663), .C2(n17230), .ZN(P2_U3221) );
  INV_X1 U19102 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19758) );
  OAI222_X1 U19103 ( .A1(n17226), .A2(n16663), .B1(n19758), .B2(n17237), .C1(
        n13048), .C2(n17230), .ZN(P2_U3222) );
  INV_X1 U19104 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U19105 ( .A1(n17226), .A2(n13048), .B1(n19760), .B2(n17237), .C1(
        n13055), .C2(n17230), .ZN(P2_U3223) );
  INV_X1 U19106 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U19107 ( .A1(n17226), .A2(n13055), .B1(n19762), .B2(n17237), .C1(
        n13056), .C2(n17230), .ZN(P2_U3224) );
  INV_X1 U19108 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19764) );
  OAI222_X1 U19109 ( .A1(n17226), .A2(n13056), .B1(n19764), .B2(n17237), .C1(
        n13062), .C2(n17230), .ZN(P2_U3225) );
  INV_X1 U19110 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19766) );
  OAI222_X1 U19111 ( .A1(n17226), .A2(n13062), .B1(n19766), .B2(n17237), .C1(
        n13063), .C2(n17230), .ZN(P2_U3226) );
  INV_X1 U19112 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19768) );
  OAI222_X1 U19113 ( .A1(n17226), .A2(n13063), .B1(n19768), .B2(n17237), .C1(
        n18439), .C2(n17230), .ZN(P2_U3227) );
  INV_X1 U19114 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19770) );
  OAI222_X1 U19115 ( .A1(n17226), .A2(n18439), .B1(n19770), .B2(n17237), .C1(
        n18452), .C2(n17230), .ZN(P2_U3228) );
  INV_X1 U19116 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19772) );
  OAI222_X1 U19117 ( .A1(n17230), .A2(n17220), .B1(n19772), .B2(n17237), .C1(
        n18452), .C2(n17226), .ZN(P2_U3229) );
  INV_X1 U19118 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19774) );
  OAI222_X1 U19119 ( .A1(n17226), .A2(n17220), .B1(n19774), .B2(n17237), .C1(
        n17221), .C2(n17230), .ZN(P2_U3230) );
  INV_X1 U19120 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19776) );
  OAI222_X1 U19121 ( .A1(n17230), .A2(n18474), .B1(n19776), .B2(n17237), .C1(
        n17221), .C2(n17226), .ZN(P2_U3231) );
  INV_X1 U19122 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19778) );
  OAI222_X1 U19123 ( .A1(n17230), .A2(n13077), .B1(n19778), .B2(n17237), .C1(
        n18474), .C2(n17226), .ZN(P2_U3232) );
  INV_X1 U19124 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19780) );
  OAI222_X1 U19125 ( .A1(n17230), .A2(n17222), .B1(n19780), .B2(n17237), .C1(
        n13077), .C2(n17226), .ZN(P2_U3233) );
  INV_X1 U19126 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19782) );
  OAI222_X1 U19127 ( .A1(n17230), .A2(n17223), .B1(n19782), .B2(n17237), .C1(
        n17222), .C2(n17226), .ZN(P2_U3234) );
  INV_X1 U19128 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19784) );
  OAI222_X1 U19129 ( .A1(n17230), .A2(n17224), .B1(n19784), .B2(n17237), .C1(
        n17223), .C2(n17226), .ZN(P2_U3235) );
  INV_X1 U19130 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19787) );
  OAI222_X1 U19131 ( .A1(n17226), .A2(n17224), .B1(n19787), .B2(n17237), .C1(
        n18521), .C2(n17230), .ZN(P2_U3236) );
  INV_X1 U19132 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17225) );
  INV_X1 U19133 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19789) );
  OAI222_X1 U19134 ( .A1(n17230), .A2(n17225), .B1(n19789), .B2(n17237), .C1(
        n18521), .C2(n17226), .ZN(P2_U3237) );
  INV_X1 U19135 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19791) );
  OAI222_X1 U19136 ( .A1(n17226), .A2(n17225), .B1(n19791), .B2(n17237), .C1(
        n16291), .C2(n17230), .ZN(P2_U3238) );
  INV_X1 U19137 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19793) );
  OAI222_X1 U19138 ( .A1(n17226), .A2(n16291), .B1(n19793), .B2(n17237), .C1(
        n17227), .C2(n17230), .ZN(P2_U3239) );
  INV_X1 U19139 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19795) );
  OAI222_X1 U19140 ( .A1(n17226), .A2(n17227), .B1(n19795), .B2(n17237), .C1(
        n17228), .C2(n17230), .ZN(P2_U3240) );
  INV_X1 U19141 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19798) );
  OAI222_X1 U19142 ( .A1(n17230), .A2(n17229), .B1(n19798), .B2(n17237), .C1(
        n17228), .C2(n17226), .ZN(P2_U3241) );
  INV_X1 U19143 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U19144 ( .A1(n17237), .A2(n17232), .B1(n17231), .B2(n21736), .ZN(
        P2_U3588) );
  INV_X1 U19145 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U19146 ( .A1(n17237), .A2(n17234), .B1(n17233), .B2(n21736), .ZN(
        P2_U3587) );
  MUX2_X1 U19147 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n17237), .Z(P2_U3586) );
  INV_X1 U19148 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U19149 ( .A1(n17237), .A2(n17236), .B1(n17235), .B2(n21736), .ZN(
        P2_U3585) );
  NOR3_X1 U19150 ( .A1(n20649), .A2(n17239), .A3(n17238), .ZN(n17240) );
  INV_X1 U19151 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18881) );
  NAND3_X1 U19152 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17245) );
  NOR2_X1 U19153 ( .A1(n20153), .A2(n17245), .ZN(n17278) );
  NAND3_X1 U19154 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17611), .A3(n17278), .ZN(
        n17262) );
  OAI221_X1 U19155 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17611), .C1(
        P3_EBX_REG_4__SCAN_IN), .C2(n17278), .A(n17262), .ZN(n17242) );
  AOI22_X1 U19156 ( .A1(n17609), .A2(n18881), .B1(n17242), .B2(n17606), .ZN(
        P3_U2699) );
  NAND2_X1 U19157 ( .A1(n20585), .A2(n17611), .ZN(n17607) );
  OR2_X1 U19158 ( .A1(n17245), .A2(n17607), .ZN(n17244) );
  INV_X1 U19159 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18922) );
  NAND3_X1 U19160 ( .A1(n17244), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17606), .ZN(
        n17243) );
  OAI221_X1 U19161 ( .B1(n17244), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17606), 
        .C2(n18922), .A(n17243), .ZN(P3_U2700) );
  INV_X1 U19162 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20126) );
  INV_X1 U19163 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20125) );
  NOR2_X1 U19164 ( .A1(n20126), .A2(n20125), .ZN(n17604) );
  AOI21_X1 U19165 ( .B1(n17611), .B2(n17604), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17247) );
  OAI21_X1 U19166 ( .B1(n17245), .B2(n17607), .A(n17606), .ZN(n17246) );
  INV_X1 U19167 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18963) );
  OAI22_X1 U19168 ( .A1(n17247), .A2(n17246), .B1(n18963), .B2(n17606), .ZN(
        P3_U2701) );
  AOI22_X1 U19169 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U19170 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U19171 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U19172 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17248) );
  NAND4_X1 U19173 ( .A1(n17251), .A2(n17250), .A3(n17249), .A4(n17248), .ZN(
        n17257) );
  AOI22_X1 U19174 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U19175 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U19176 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U19177 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17252) );
  NAND4_X1 U19178 ( .A1(n17255), .A2(n17254), .A3(n17253), .A4(n17252), .ZN(
        n17256) );
  NOR2_X1 U19179 ( .A1(n17257), .A2(n17256), .ZN(n20725) );
  INV_X1 U19180 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20225) );
  NAND3_X1 U19181 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n17280) );
  NOR2_X1 U19182 ( .A1(n17280), .A2(n17262), .ZN(n17258) );
  INV_X1 U19183 ( .A(n17258), .ZN(n17260) );
  NOR2_X1 U19184 ( .A1(n20225), .A2(n17260), .ZN(n17377) );
  OAI21_X1 U19185 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17258), .A(n17606), .ZN(
        n17259) );
  OAI22_X1 U19186 ( .A1(n20725), .A2(n17606), .B1(n17377), .B2(n17259), .ZN(
        P3_U2695) );
  INV_X1 U19187 ( .A(n17262), .ZN(n17265) );
  AND3_X1 U19188 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17265), .A3(
        P3_EBX_REG_5__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U19189 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17264), .A(n17260), .ZN(
        n17261) );
  AOI22_X1 U19190 ( .A1(n17609), .A2(n18760), .B1(n17261), .B2(n17606), .ZN(
        P3_U2696) );
  NOR3_X1 U19191 ( .A1(n20649), .A2(n20181), .A3(n17262), .ZN(n17267) );
  AOI21_X1 U19192 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17606), .A(n17267), .ZN(
        n17263) );
  INV_X1 U19193 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18800) );
  OAI22_X1 U19194 ( .A1(n17264), .A2(n17263), .B1(n18800), .B2(n17606), .ZN(
        P3_U2697) );
  OAI21_X1 U19195 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17265), .A(n17606), .ZN(
        n17266) );
  OAI22_X1 U19196 ( .A1(n17267), .A2(n17266), .B1(n18841), .B2(n17606), .ZN(
        P3_U2698) );
  AOI22_X1 U19197 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U19198 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U19199 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U19200 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17268) );
  NAND4_X1 U19201 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17277) );
  AOI22_X1 U19202 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U19203 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U19204 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U19205 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17272) );
  NAND4_X1 U19206 ( .A1(n17275), .A2(n17274), .A3(n17273), .A4(n17272), .ZN(
        n17276) );
  NOR2_X1 U19207 ( .A1(n17277), .A2(n17276), .ZN(n20705) );
  NAND3_X1 U19208 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17571) );
  NAND4_X1 U19209 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_4__SCAN_IN), .A4(n17278), .ZN(n17279) );
  NOR4_X1 U19210 ( .A1(n20239), .A2(n20225), .A3(n17280), .A4(n17279), .ZN(
        n17297) );
  NAND2_X1 U19211 ( .A1(n17611), .A2(n17297), .ZN(n17348) );
  INV_X1 U19212 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17572) );
  INV_X1 U19213 ( .A(n17379), .ZN(n17281) );
  OAI33_X1 U19214 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20649), .A3(n17379), 
        .B1(n17572), .B2(n17609), .B3(n17281), .ZN(n17282) );
  INV_X1 U19215 ( .A(n17282), .ZN(n17283) );
  OAI21_X1 U19216 ( .B1(n20705), .B2(n17606), .A(n17283), .ZN(P3_U2687) );
  AOI22_X1 U19217 ( .A1(n10998), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U19218 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15360), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U19219 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17284) );
  OAI21_X1 U19220 ( .B1(n11387), .B2(n18760), .A(n17284), .ZN(n17290) );
  AOI22_X1 U19221 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U19222 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U19223 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U19224 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17285) );
  NAND4_X1 U19225 ( .A1(n17288), .A2(n17287), .A3(n17286), .A4(n17285), .ZN(
        n17289) );
  AOI211_X1 U19226 ( .C1(n10996), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17290), .B(n17289), .ZN(n17291) );
  NAND3_X1 U19227 ( .A1(n17293), .A2(n17292), .A3(n17291), .ZN(n20714) );
  INV_X1 U19228 ( .A(n20714), .ZN(n17296) );
  OAI211_X1 U19229 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17294), .A(n17379), .B(
        n17606), .ZN(n17295) );
  OAI21_X1 U19230 ( .B1(n17296), .B2(n17606), .A(n17295), .ZN(P3_U2688) );
  INV_X1 U19231 ( .A(n17607), .ZN(n17608) );
  INV_X1 U19232 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20282) );
  NAND2_X1 U19233 ( .A1(n17608), .A2(n20282), .ZN(n17323) );
  NAND2_X1 U19234 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17297), .ZN(n17309) );
  AOI22_X1 U19235 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U19236 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U19237 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U19238 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17298) );
  NAND4_X1 U19239 ( .A1(n17301), .A2(n17300), .A3(n17299), .A4(n17298), .ZN(
        n17307) );
  AOI22_X1 U19240 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U19241 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U19242 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U19243 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17302) );
  NAND4_X1 U19244 ( .A1(n17305), .A2(n17304), .A3(n17303), .A4(n17302), .ZN(
        n17306) );
  NOR2_X1 U19245 ( .A1(n17307), .A2(n17306), .ZN(n20559) );
  INV_X1 U19246 ( .A(n17611), .ZN(n17308) );
  AOI21_X1 U19247 ( .B1(n20585), .B2(n17309), .A(n17308), .ZN(n17322) );
  OAI222_X1 U19248 ( .A1(n17323), .A2(n17309), .B1(n17606), .B2(n20559), .C1(
        n20282), .C2(n17322), .ZN(P3_U2690) );
  INV_X1 U19249 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20305) );
  AOI22_X1 U19250 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U19251 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U19252 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U19253 ( .B1(n11387), .B2(n18800), .A(n17310), .ZN(n17316) );
  AOI22_X1 U19254 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U19255 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U19256 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U19257 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17311) );
  NAND4_X1 U19258 ( .A1(n17314), .A2(n17313), .A3(n17312), .A4(n17311), .ZN(
        n17315) );
  AOI211_X1 U19259 ( .C1(n17701), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17316), .B(n17315), .ZN(n17317) );
  NAND3_X1 U19260 ( .A1(n17319), .A2(n17318), .A3(n17317), .ZN(n20709) );
  NOR2_X1 U19261 ( .A1(n20649), .A2(n17348), .ZN(n17574) );
  INV_X1 U19262 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17334) );
  NOR3_X1 U19263 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20282), .A3(n17334), .ZN(
        n17320) );
  AOI22_X1 U19264 ( .A1(n17609), .A2(n20709), .B1(n17574), .B2(n17320), .ZN(
        n17321) );
  OAI221_X1 U19265 ( .B1(n20305), .B2(n17323), .C1(n20305), .C2(n17322), .A(
        n17321), .ZN(P3_U2689) );
  AOI22_X1 U19266 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U19267 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U19268 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U19269 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17324) );
  NAND4_X1 U19270 ( .A1(n17327), .A2(n17326), .A3(n17325), .A4(n17324), .ZN(
        n17333) );
  AOI22_X1 U19271 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U19272 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U19273 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19274 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17328) );
  NAND4_X1 U19275 ( .A1(n17331), .A2(n17330), .A3(n17329), .A4(n17328), .ZN(
        n17332) );
  NOR2_X1 U19276 ( .A1(n17333), .A2(n17332), .ZN(n20564) );
  AND2_X1 U19277 ( .A1(n17606), .A2(n17348), .ZN(n17335) );
  AOI22_X1 U19278 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17335), .B1(n17574), 
        .B2(n17334), .ZN(n17336) );
  OAI21_X1 U19279 ( .B1(n20564), .B2(n17606), .A(n17336), .ZN(P3_U2691) );
  AOI22_X1 U19280 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U19281 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U19282 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U19283 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17337) );
  NAND4_X1 U19284 ( .A1(n17340), .A2(n17339), .A3(n17338), .A4(n17337), .ZN(
        n17347) );
  AOI22_X1 U19285 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U19286 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U19287 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U19288 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17342) );
  NAND4_X1 U19289 ( .A1(n17345), .A2(n17344), .A3(n17343), .A4(n17342), .ZN(
        n17346) );
  NOR2_X1 U19290 ( .A1(n17347), .A2(n17346), .ZN(n20569) );
  INV_X1 U19291 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20249) );
  NAND2_X1 U19292 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17377), .ZN(n17376) );
  NOR2_X1 U19293 ( .A1(n20249), .A2(n17376), .ZN(n17362) );
  OAI211_X1 U19294 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17362), .A(n17348), .B(
        n17606), .ZN(n17349) );
  OAI21_X1 U19295 ( .B1(n20569), .B2(n17606), .A(n17349), .ZN(P3_U2692) );
  AOI22_X1 U19296 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U19297 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17662), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U19298 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17350) );
  OAI21_X1 U19299 ( .B1(n11387), .B2(n18963), .A(n17350), .ZN(n17356) );
  AOI22_X1 U19300 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U19301 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U19302 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U19303 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17351) );
  NAND4_X1 U19304 ( .A1(n17354), .A2(n17353), .A3(n17352), .A4(n17351), .ZN(
        n17355) );
  AOI211_X1 U19305 ( .C1(n15360), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17356), .B(n17355), .ZN(n17357) );
  NAND3_X1 U19306 ( .A1(n17359), .A2(n17358), .A3(n17357), .ZN(n20574) );
  INV_X1 U19307 ( .A(n20574), .ZN(n17363) );
  INV_X1 U19308 ( .A(n17376), .ZN(n17360) );
  OAI21_X1 U19309 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17360), .A(n17606), .ZN(
        n17361) );
  OAI22_X1 U19310 ( .A1(n17363), .A2(n17606), .B1(n17362), .B2(n17361), .ZN(
        P3_U2693) );
  AOI22_X1 U19311 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n10997), .ZN(n17368) );
  AOI22_X1 U19312 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17700), .ZN(n17367) );
  AOI22_X1 U19313 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10994), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17590), .ZN(n17366) );
  AOI22_X1 U19314 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20172), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17681), .ZN(n17365) );
  NAND4_X1 U19315 ( .A1(n17368), .A2(n17367), .A3(n17366), .A4(n17365), .ZN(
        n17375) );
  AOI22_X1 U19316 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15360), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17643), .ZN(n17373) );
  AOI22_X1 U19317 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U19318 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n10998), .ZN(n17371) );
  AOI22_X1 U19319 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17370) );
  NAND4_X1 U19320 ( .A1(n17373), .A2(n17372), .A3(n17371), .A4(n17370), .ZN(
        n17374) );
  NOR2_X1 U19321 ( .A1(n17375), .A2(n17374), .ZN(n20580) );
  OAI21_X1 U19322 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17377), .A(n17376), .ZN(
        n17378) );
  AOI22_X1 U19323 ( .A1(n17609), .A2(n20580), .B1(n17378), .B2(n17606), .ZN(
        P3_U2694) );
  INV_X1 U19324 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20533) );
  INV_X1 U19325 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20364) );
  NAND2_X1 U19326 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17588), .ZN(n17587) );
  INV_X1 U19327 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17381) );
  INV_X1 U19328 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20495) );
  INV_X1 U19329 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20404) );
  NAND4_X1 U19330 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n17380)
         );
  NOR4_X1 U19331 ( .A1(n17381), .A2(n20495), .A3(n20404), .A4(n17380), .ZN(
        n17382) );
  NAND4_X1 U19332 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17484), .A4(n17382), .ZN(n17481) );
  NOR2_X1 U19333 ( .A1(n20533), .A2(n17481), .ZN(n17480) );
  NAND2_X1 U19334 ( .A1(n17606), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U19335 ( .A1(n17480), .A2(n20585), .ZN(n17383) );
  OAI22_X1 U19336 ( .A1(n17480), .A2(n17384), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17383), .ZN(P3_U2672) );
  AOI22_X1 U19337 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U19338 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U19339 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U19340 ( .A1(n10998), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17385) );
  NAND4_X1 U19341 ( .A1(n17388), .A2(n17387), .A3(n17386), .A4(n17385), .ZN(
        n17394) );
  AOI22_X1 U19342 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17662), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U19343 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U19344 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U19345 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17389) );
  NAND4_X1 U19346 ( .A1(n17392), .A2(n17391), .A3(n17390), .A4(n17389), .ZN(
        n17393) );
  NOR2_X1 U19347 ( .A1(n17394), .A2(n17393), .ZN(n17479) );
  AOI22_X1 U19348 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U19349 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U19350 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U19351 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17395) );
  NAND4_X1 U19352 ( .A1(n17398), .A2(n17397), .A3(n17396), .A4(n17395), .ZN(
        n17404) );
  AOI22_X1 U19353 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U19354 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U19355 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U19356 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17399) );
  NAND4_X1 U19357 ( .A1(n17402), .A2(n17401), .A3(n17400), .A4(n17399), .ZN(
        n17403) );
  NOR2_X1 U19358 ( .A1(n17404), .A2(n17403), .ZN(n17504) );
  AOI22_X1 U19359 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U19360 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U19361 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U19362 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17405) );
  NAND4_X1 U19363 ( .A1(n17408), .A2(n17407), .A3(n17406), .A4(n17405), .ZN(
        n17415) );
  AOI22_X1 U19364 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U19365 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U19366 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U19367 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17410) );
  NAND4_X1 U19368 ( .A1(n17413), .A2(n17412), .A3(n17411), .A4(n17410), .ZN(
        n17414) );
  NOR2_X1 U19369 ( .A1(n17415), .A2(n17414), .ZN(n17498) );
  AOI22_X1 U19370 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U19371 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U19372 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U19373 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17416) );
  NAND4_X1 U19374 ( .A1(n17419), .A2(n17418), .A3(n17417), .A4(n17416), .ZN(
        n17425) );
  AOI22_X1 U19375 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U19376 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U19377 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U19378 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15360), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17420) );
  NAND4_X1 U19379 ( .A1(n17423), .A2(n17422), .A3(n17421), .A4(n17420), .ZN(
        n17424) );
  NOR2_X1 U19380 ( .A1(n17425), .A2(n17424), .ZN(n17519) );
  AOI22_X1 U19381 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U19382 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U19383 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U19384 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17426) );
  NAND4_X1 U19385 ( .A1(n17429), .A2(n17428), .A3(n17427), .A4(n17426), .ZN(
        n17435) );
  AOI22_X1 U19386 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U19387 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U19388 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U19389 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17430) );
  NAND4_X1 U19390 ( .A1(n17433), .A2(n17432), .A3(n17431), .A4(n17430), .ZN(
        n17434) );
  NOR2_X1 U19391 ( .A1(n17435), .A2(n17434), .ZN(n17529) );
  AOI22_X1 U19392 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U19393 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U19394 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U19395 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17436) );
  NAND4_X1 U19396 ( .A1(n17439), .A2(n17438), .A3(n17437), .A4(n17436), .ZN(
        n17445) );
  AOI22_X1 U19397 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U19398 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U19399 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U19400 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17440) );
  NAND4_X1 U19401 ( .A1(n17443), .A2(n17442), .A3(n17441), .A4(n17440), .ZN(
        n17444) );
  NOR2_X1 U19402 ( .A1(n17445), .A2(n17444), .ZN(n17530) );
  NOR2_X1 U19403 ( .A1(n17529), .A2(n17530), .ZN(n17528) );
  AOI22_X1 U19404 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10991), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U19405 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10997), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U19406 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10998), .ZN(n17446) );
  OAI21_X1 U19407 ( .B1(n17469), .B2(n19008), .A(n17446), .ZN(n17452) );
  AOI22_X1 U19408 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17650), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U19409 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15306), .ZN(n17449) );
  AOI22_X1 U19410 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17681), .ZN(n17448) );
  AOI22_X1 U19411 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17590), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17447) );
  NAND4_X1 U19412 ( .A1(n17450), .A2(n17449), .A3(n17448), .A4(n17447), .ZN(
        n17451) );
  AOI211_X1 U19413 ( .C1(n17671), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n17452), .B(n17451), .ZN(n17453) );
  NAND3_X1 U19414 ( .A1(n17455), .A2(n17454), .A3(n17453), .ZN(n17524) );
  NAND2_X1 U19415 ( .A1(n17528), .A2(n17524), .ZN(n17523) );
  NOR2_X1 U19416 ( .A1(n17519), .A2(n17523), .ZN(n17518) );
  AOI22_X1 U19417 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U19418 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U19419 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U19420 ( .B1(n17469), .B2(n18922), .A(n17457), .ZN(n17463) );
  AOI22_X1 U19421 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U19422 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U19423 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U19424 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17458) );
  NAND4_X1 U19425 ( .A1(n17461), .A2(n17460), .A3(n17459), .A4(n17458), .ZN(
        n17462) );
  AOI211_X1 U19426 ( .C1(n17701), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17463), .B(n17462), .ZN(n17464) );
  NAND3_X1 U19427 ( .A1(n17466), .A2(n17465), .A3(n17464), .ZN(n17514) );
  NAND2_X1 U19428 ( .A1(n17518), .A2(n17514), .ZN(n17513) );
  NOR2_X1 U19429 ( .A1(n17498), .A2(n17513), .ZN(n17510) );
  AOI22_X1 U19430 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U19431 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U19432 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U19433 ( .B1(n17469), .B2(n18841), .A(n17468), .ZN(n17475) );
  AOI22_X1 U19434 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U19435 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U19436 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19437 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17470) );
  NAND4_X1 U19438 ( .A1(n17473), .A2(n17472), .A3(n17471), .A4(n17470), .ZN(
        n17474) );
  AOI211_X1 U19439 ( .C1(n17671), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n17475), .B(n17474), .ZN(n17476) );
  NAND3_X1 U19440 ( .A1(n17478), .A2(n17477), .A3(n17476), .ZN(n17509) );
  NAND2_X1 U19441 ( .A1(n17510), .A2(n17509), .ZN(n17508) );
  NOR2_X1 U19442 ( .A1(n17504), .A2(n17508), .ZN(n17503) );
  XNOR2_X1 U19443 ( .A(n17479), .B(n17503), .ZN(n20663) );
  AOI211_X1 U19444 ( .C1(n20533), .C2(n17481), .A(n17480), .B(n17609), .ZN(
        n17482) );
  AOI21_X1 U19445 ( .B1(n17609), .B2(n20663), .A(n17482), .ZN(n17483) );
  INV_X1 U19446 ( .A(n17483), .ZN(P3_U2673) );
  NAND2_X1 U19447 ( .A1(n20585), .A2(n17484), .ZN(n17497) );
  NOR2_X1 U19448 ( .A1(n17609), .A2(n17484), .ZN(n17558) );
  AOI22_X1 U19449 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U19450 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U19451 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U19452 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17485) );
  NAND4_X1 U19453 ( .A1(n17488), .A2(n17487), .A3(n17486), .A4(n17485), .ZN(
        n17494) );
  AOI22_X1 U19454 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19455 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U19456 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U19457 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17489) );
  NAND4_X1 U19458 ( .A1(n17492), .A2(n17491), .A3(n17490), .A4(n17489), .ZN(
        n17493) );
  NOR2_X1 U19459 ( .A1(n17494), .A2(n17493), .ZN(n20619) );
  INV_X1 U19460 ( .A(n20619), .ZN(n17495) );
  AOI22_X1 U19461 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17558), .B1(n17609), 
        .B2(n17495), .ZN(n17496) );
  OAI21_X1 U19462 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17497), .A(n17496), .ZN(
        P3_U2682) );
  INV_X1 U19463 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20457) );
  INV_X1 U19464 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20435) );
  NAND2_X1 U19465 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17534), .ZN(n17527) );
  NAND2_X1 U19466 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17533), .ZN(n17517) );
  NAND2_X1 U19467 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17516), .ZN(n17512) );
  INV_X1 U19468 ( .A(n17512), .ZN(n17501) );
  AOI21_X1 U19469 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17606), .A(n17516), .ZN(
        n17500) );
  AOI21_X1 U19470 ( .B1(n17498), .B2(n17513), .A(n17510), .ZN(n20684) );
  INV_X1 U19471 ( .A(n20684), .ZN(n17499) );
  OAI22_X1 U19472 ( .A1(n17501), .A2(n17500), .B1(n17606), .B2(n17499), .ZN(
        P3_U2676) );
  NAND2_X1 U19473 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17501), .ZN(n17507) );
  NAND2_X1 U19474 ( .A1(n17606), .A2(n17512), .ZN(n17502) );
  OAI21_X1 U19475 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17607), .A(n17502), .ZN(
        n17505) );
  AOI21_X1 U19476 ( .B1(n17504), .B2(n17508), .A(n17503), .ZN(n20672) );
  AOI22_X1 U19477 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17505), .B1(n20672), 
        .B2(n17609), .ZN(n17506) );
  OAI21_X1 U19478 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17507), .A(n17506), .ZN(
        P3_U2674) );
  OAI21_X1 U19479 ( .B1(n17510), .B2(n17509), .A(n17508), .ZN(n20678) );
  NAND3_X1 U19480 ( .A1(n17512), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n17606), 
        .ZN(n17511) );
  OAI221_X1 U19481 ( .B1(n17512), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n17606), 
        .C2(n20678), .A(n17511), .ZN(P3_U2675) );
  AOI21_X1 U19482 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17606), .A(n17522), .ZN(
        n17515) );
  OAI21_X1 U19483 ( .B1(n17518), .B2(n17514), .A(n17513), .ZN(n20659) );
  OAI22_X1 U19484 ( .A1(n17516), .A2(n17515), .B1(n17606), .B2(n20659), .ZN(
        P3_U2677) );
  INV_X1 U19485 ( .A(n17517), .ZN(n17526) );
  AOI21_X1 U19486 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17606), .A(n17526), .ZN(
        n17521) );
  AOI21_X1 U19487 ( .B1(n17519), .B2(n17523), .A(n17518), .ZN(n20653) );
  INV_X1 U19488 ( .A(n20653), .ZN(n17520) );
  OAI22_X1 U19489 ( .A1(n17522), .A2(n17521), .B1(n17606), .B2(n17520), .ZN(
        P3_U2678) );
  AOI21_X1 U19490 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17606), .A(n17533), .ZN(
        n17525) );
  OAI21_X1 U19491 ( .B1(n17528), .B2(n17524), .A(n17523), .ZN(n20691) );
  OAI22_X1 U19492 ( .A1(n17526), .A2(n17525), .B1(n17606), .B2(n20691), .ZN(
        P3_U2679) );
  INV_X1 U19493 ( .A(n17527), .ZN(n17547) );
  AOI21_X1 U19494 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17606), .A(n17547), .ZN(
        n17532) );
  AOI21_X1 U19495 ( .B1(n17530), .B2(n17529), .A(n17528), .ZN(n20692) );
  INV_X1 U19496 ( .A(n20692), .ZN(n17531) );
  OAI22_X1 U19497 ( .A1(n17533), .A2(n17532), .B1(n17606), .B2(n17531), .ZN(
        P3_U2680) );
  AOI21_X1 U19498 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17606), .A(n17534), .ZN(
        n17546) );
  AOI22_X1 U19499 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U19500 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U19501 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U19502 ( .B1(n15367), .B2(n18800), .A(n17535), .ZN(n17541) );
  AOI22_X1 U19503 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U19504 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U19505 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U19506 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17536) );
  NAND4_X1 U19507 ( .A1(n17539), .A2(n17538), .A3(n17537), .A4(n17536), .ZN(
        n17540) );
  AOI211_X1 U19508 ( .C1(n17701), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17541), .B(n17540), .ZN(n17542) );
  NAND3_X1 U19509 ( .A1(n17544), .A2(n17543), .A3(n17542), .ZN(n20624) );
  INV_X1 U19510 ( .A(n20624), .ZN(n17545) );
  OAI22_X1 U19511 ( .A1(n17547), .A2(n17546), .B1(n17545), .B2(n17606), .ZN(
        P3_U2681) );
  AOI22_X1 U19512 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U19513 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U19514 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17549) );
  AOI22_X1 U19515 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17548) );
  NAND4_X1 U19516 ( .A1(n17551), .A2(n17550), .A3(n17549), .A4(n17548), .ZN(
        n17557) );
  AOI22_X1 U19517 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U19518 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U19519 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17553) );
  AOI22_X1 U19520 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17552) );
  NAND4_X1 U19521 ( .A1(n17555), .A2(n17554), .A3(n17553), .A4(n17552), .ZN(
        n17556) );
  NOR2_X1 U19522 ( .A1(n17557), .A2(n17556), .ZN(n20623) );
  OAI21_X1 U19523 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17559), .A(n17558), .ZN(
        n17560) );
  OAI21_X1 U19524 ( .B1(n20623), .B2(n17606), .A(n17560), .ZN(P3_U2683) );
  NAND2_X1 U19525 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17601), .ZN(n17576) );
  AOI22_X1 U19526 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17564) );
  AOI22_X1 U19527 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U19528 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17562) );
  AOI22_X1 U19529 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17561) );
  NAND4_X1 U19530 ( .A1(n17564), .A2(n17563), .A3(n17562), .A4(n17561), .ZN(
        n17570) );
  AOI22_X1 U19531 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U19532 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U19533 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U19534 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17565) );
  NAND4_X1 U19535 ( .A1(n17568), .A2(n17567), .A3(n17566), .A4(n17565), .ZN(
        n17569) );
  NOR2_X1 U19536 ( .A1(n17570), .A2(n17569), .ZN(n20640) );
  INV_X1 U19537 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20316) );
  NOR3_X1 U19538 ( .A1(n17572), .A2(n20316), .A3(n17571), .ZN(n17573) );
  NAND4_X1 U19539 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17574), .A3(n17573), 
        .A4(n20364), .ZN(n17575) );
  OAI221_X1 U19540 ( .B1(n17609), .B2(n17576), .C1(n17606), .C2(n20640), .A(
        n17575), .ZN(P3_U2685) );
  AOI22_X1 U19541 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17663), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U19542 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17579) );
  AOI22_X1 U19543 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U19544 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17577) );
  NAND4_X1 U19545 ( .A1(n17580), .A2(n17579), .A3(n17578), .A4(n17577), .ZN(
        n17586) );
  AOI22_X1 U19546 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U19547 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U19548 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U19549 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17581) );
  NAND4_X1 U19550 ( .A1(n17584), .A2(n17583), .A3(n17582), .A4(n17581), .ZN(
        n17585) );
  NOR2_X1 U19551 ( .A1(n17586), .A2(n17585), .ZN(n20635) );
  OAI21_X1 U19552 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17588), .A(n17587), .ZN(
        n17589) );
  AOI22_X1 U19553 ( .A1(n17609), .A2(n20635), .B1(n17589), .B2(n17606), .ZN(
        P3_U2684) );
  AOI22_X1 U19554 ( .A1(n17662), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17409), .ZN(n17594) );
  AOI22_X1 U19555 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17643), .ZN(n17593) );
  AOI22_X1 U19556 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17681), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n20172), .ZN(n17592) );
  AOI22_X1 U19557 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17590), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n10994), .ZN(n17591) );
  NAND4_X1 U19558 ( .A1(n17594), .A2(n17593), .A3(n17592), .A4(n17591), .ZN(
        n17600) );
  AOI22_X1 U19559 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17598) );
  AOI22_X1 U19560 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U19561 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10997), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19562 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17671), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17595) );
  NAND4_X1 U19563 ( .A1(n17598), .A2(n17597), .A3(n17596), .A4(n17595), .ZN(
        n17599) );
  NOR2_X1 U19564 ( .A1(n17600), .A2(n17599), .ZN(n20645) );
  OAI21_X1 U19565 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17602), .A(n17601), .ZN(
        n17603) );
  AOI22_X1 U19566 ( .A1(n17609), .A2(n20645), .B1(n17603), .B2(n17606), .ZN(
        P3_U2686) );
  INV_X1 U19567 ( .A(n17604), .ZN(n17605) );
  OAI21_X1 U19568 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17605), .ZN(n20124) );
  OAI222_X1 U19569 ( .A1(n20124), .A2(n17607), .B1(n20125), .B2(n17611), .C1(
        n19008), .C2(n17606), .ZN(P3_U2702) );
  AOI22_X1 U19570 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17609), .B1(
        n17608), .B2(n20126), .ZN(n17610) );
  OAI21_X1 U19571 ( .B1(n17611), .B2(n20126), .A(n17610), .ZN(P3_U2703) );
  INV_X1 U19572 ( .A(n17765), .ZN(n17613) );
  OAI21_X1 U19573 ( .B1(n21250), .B2(n20062), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17612) );
  OAI21_X1 U19574 ( .B1(n17613), .B2(n21277), .A(n17612), .ZN(P3_U2634) );
  NOR2_X1 U19575 ( .A1(n20058), .A2(n18178), .ZN(n17617) );
  AOI21_X1 U19576 ( .B1(n21284), .B2(n17615), .A(n17614), .ZN(n21269) );
  NOR2_X1 U19577 ( .A1(n21269), .A2(n18676), .ZN(n17616) );
  OAI22_X1 U19578 ( .A1(n18721), .A2(n17617), .B1(n18178), .B2(n17616), .ZN(
        P3_U2863) );
  AOI22_X1 U19579 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U19580 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U19581 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U19582 ( .B1(n11386), .B2(n18760), .A(n17619), .ZN(n17625) );
  AOI22_X1 U19583 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U19584 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U19585 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U19586 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17620) );
  NAND4_X1 U19587 ( .A1(n17623), .A2(n17622), .A3(n17621), .A4(n17620), .ZN(
        n17624) );
  AOI211_X1 U19588 ( .C1(n17590), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n17625), .B(n17624), .ZN(n17626) );
  AOI22_X1 U19589 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U19590 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U19591 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U19592 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10994), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17629) );
  NAND4_X1 U19593 ( .A1(n17632), .A2(n17631), .A3(n17630), .A4(n17629), .ZN(
        n17638) );
  AOI22_X1 U19594 ( .A1(n15306), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U19595 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17635) );
  AOI22_X1 U19596 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U19597 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10996), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17633) );
  NAND4_X1 U19598 ( .A1(n17636), .A2(n17635), .A3(n17634), .A4(n17633), .ZN(
        n17637) );
  AOI22_X1 U19599 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U19600 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17641) );
  AOI22_X1 U19601 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17640) );
  AOI22_X1 U19602 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17639) );
  NAND4_X1 U19603 ( .A1(n17642), .A2(n17641), .A3(n17640), .A4(n17639), .ZN(
        n17649) );
  AOI22_X1 U19604 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U19605 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19606 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U19607 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17644) );
  NAND4_X1 U19608 ( .A1(n17647), .A2(n17646), .A3(n17645), .A4(n17644), .ZN(
        n17648) );
  AOI22_X1 U19609 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17650), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U19610 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U19611 ( .A1(n15348), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17651) );
  OAI21_X1 U19612 ( .B1(n11386), .B2(n18963), .A(n17651), .ZN(n17656) );
  AOI22_X1 U19613 ( .A1(n17663), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17364), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17655) );
  AOI22_X1 U19614 ( .A1(n17661), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17467), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U19615 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17652), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17653) );
  NAND3_X1 U19616 ( .A1(n17659), .A2(n17658), .A3(n17657), .ZN(n20610) );
  AOI22_X1 U19617 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10994), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17681), .ZN(n17660) );
  AOI22_X1 U19618 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17661), .ZN(n17667) );
  AOI22_X1 U19619 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17456), .ZN(n17666) );
  AOI22_X1 U19620 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17662), .B1(
        n17467), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U19621 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17663), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U19622 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17652), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U19623 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U19624 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U19625 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17670) );
  OAI21_X1 U19626 ( .B1(n11386), .B2(n18881), .A(n17670), .ZN(n17677) );
  AOI22_X1 U19627 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U19628 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17702), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19629 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U19630 ( .A1(n10991), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17672) );
  NAND4_X1 U19631 ( .A1(n17675), .A2(n17674), .A3(n17673), .A4(n17672), .ZN(
        n17676) );
  AOI211_X1 U19632 ( .C1(n17590), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17677), .B(n17676), .ZN(n17678) );
  NAND3_X1 U19633 ( .A1(n17680), .A2(n17679), .A3(n17678), .ZN(n17737) );
  NAND2_X1 U19634 ( .A1(n17693), .A2(n17737), .ZN(n17720) );
  AOI22_X1 U19635 ( .A1(n17695), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U19636 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U19637 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17682) );
  OAI21_X1 U19638 ( .B1(n11386), .B2(n18800), .A(n17682), .ZN(n17688) );
  AOI22_X1 U19639 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U19640 ( .A1(n15365), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17685) );
  AOI22_X1 U19641 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U19642 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17683) );
  NAND4_X1 U19643 ( .A1(n17686), .A2(n17685), .A3(n17684), .A4(n17683), .ZN(
        n17687) );
  AOI211_X1 U19644 ( .C1(n17590), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17688), .B(n17687), .ZN(n17689) );
  NAND3_X1 U19645 ( .A1(n17691), .A2(n17690), .A3(n17689), .ZN(n17738) );
  INV_X1 U19646 ( .A(n17738), .ZN(n20592) );
  XNOR2_X1 U19647 ( .A(n20592), .B(n17692), .ZN(n17725) );
  NAND2_X1 U19648 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17725), .ZN(
        n17726) );
  INV_X1 U19649 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20880) );
  INV_X1 U19650 ( .A(n17737), .ZN(n20601) );
  XNOR2_X1 U19651 ( .A(n20601), .B(n17693), .ZN(n17718) );
  XNOR2_X1 U19652 ( .A(n20880), .B(n17718), .ZN(n18126) );
  NAND2_X1 U19653 ( .A1(n17694), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17709) );
  AOI22_X1 U19654 ( .A1(n10996), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17695), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U19655 ( .A1(n17409), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10998), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U19656 ( .A1(n20172), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n20777), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17697) );
  AOI22_X1 U19657 ( .A1(n10994), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17681), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17696) );
  NAND4_X1 U19658 ( .A1(n17699), .A2(n17698), .A3(n17697), .A4(n17696), .ZN(
        n17708) );
  AOI22_X1 U19659 ( .A1(n17671), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U19660 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10991), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19661 ( .A1(n17702), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10997), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U19662 ( .A1(n17650), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17467), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17703) );
  NAND4_X1 U19663 ( .A1(n17706), .A2(n17705), .A3(n17704), .A4(n17703), .ZN(
        n17707) );
  INV_X1 U19664 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20846) );
  NOR2_X1 U19665 ( .A1(n20740), .A2(n20846), .ZN(n18165) );
  NAND2_X1 U19666 ( .A1(n18159), .A2(n18165), .ZN(n18158) );
  NAND2_X1 U19667 ( .A1(n17709), .A2(n18158), .ZN(n18148) );
  INV_X1 U19668 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20856) );
  INV_X1 U19669 ( .A(n17710), .ZN(n17716) );
  NOR2_X1 U19670 ( .A1(n20610), .A2(n20726), .ZN(n17711) );
  XNOR2_X1 U19671 ( .A(n20856), .B(n17712), .ZN(n18149) );
  NAND2_X1 U19672 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17712), .ZN(
        n17713) );
  NAND2_X1 U19673 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17715), .ZN(
        n17717) );
  XNOR2_X1 U19674 ( .A(n20605), .B(n17716), .ZN(n18141) );
  NAND2_X1 U19675 ( .A1(n17717), .A2(n18140), .ZN(n18125) );
  NAND2_X1 U19676 ( .A1(n18126), .A2(n18125), .ZN(n18124) );
  NAND2_X1 U19677 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17718), .ZN(
        n17719) );
  XOR2_X1 U19678 ( .A(n20596), .B(n17720), .Z(n17723) );
  NAND2_X1 U19679 ( .A1(n17723), .A2(n17722), .ZN(n17724) );
  INV_X1 U19680 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20902) );
  XNOR2_X1 U19681 ( .A(n20902), .B(n17725), .ZN(n18106) );
  AOI21_X1 U19682 ( .B1(n20811), .B2(n21090), .A(n17976), .ZN(n17728) );
  NAND2_X1 U19683 ( .A1(n17728), .A2(n17792), .ZN(n17729) );
  INV_X1 U19684 ( .A(n20808), .ZN(n21225) );
  NOR2_X1 U19685 ( .A1(n17732), .A2(n17731), .ZN(n20782) );
  AND2_X1 U19686 ( .A1(n20796), .A2(n17733), .ZN(n20753) );
  INV_X1 U19687 ( .A(n17734), .ZN(n17736) );
  AOI21_X1 U19688 ( .B1(n17736), .B2(n17735), .A(n21249), .ZN(n21229) );
  NOR2_X2 U19689 ( .A1(n21086), .A2(n18170), .ZN(n18088) );
  NAND2_X2 U19690 ( .A1(n20800), .A2(n21282), .ZN(n18171) );
  INV_X1 U19691 ( .A(n20740), .ZN(n17750) );
  AOI21_X1 U19692 ( .B1(n20726), .B2(n17750), .A(n20610), .ZN(n17744) );
  NOR2_X1 U19693 ( .A1(n20605), .A2(n17744), .ZN(n17743) );
  NAND2_X1 U19694 ( .A1(n17743), .A2(n17737), .ZN(n17741) );
  NOR2_X1 U19695 ( .A1(n20596), .A2(n17741), .ZN(n17740) );
  NAND2_X1 U19696 ( .A1(n17740), .A2(n17738), .ZN(n17739) );
  NOR2_X1 U19697 ( .A1(n20811), .A2(n17739), .ZN(n17763) );
  XNOR2_X1 U19698 ( .A(n21086), .B(n17739), .ZN(n18098) );
  XNOR2_X1 U19699 ( .A(n20592), .B(n17740), .ZN(n17758) );
  XOR2_X1 U19700 ( .A(n20596), .B(n17741), .Z(n17742) );
  NAND2_X1 U19701 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17742), .ZN(
        n17756) );
  INV_X1 U19702 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20888) );
  XNOR2_X1 U19703 ( .A(n20888), .B(n17742), .ZN(n18120) );
  XNOR2_X1 U19704 ( .A(n20601), .B(n17743), .ZN(n17753) );
  INV_X1 U19705 ( .A(n17744), .ZN(n17746) );
  XNOR2_X1 U19706 ( .A(n20605), .B(n17746), .ZN(n17745) );
  NAND2_X1 U19707 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17745), .ZN(
        n17752) );
  XNOR2_X1 U19708 ( .A(n17714), .B(n17745), .ZN(n18138) );
  OAI21_X1 U19709 ( .B1(n20740), .B2(n17710), .A(n17746), .ZN(n17747) );
  NAND2_X1 U19710 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17747), .ZN(
        n17751) );
  XOR2_X1 U19711 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n17747), .Z(
        n18152) );
  AOI21_X1 U19712 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20726), .A(
        n17750), .ZN(n17749) );
  NOR2_X1 U19713 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20726), .ZN(
        n17748) );
  AOI221_X1 U19714 ( .B1(n17750), .B2(n20726), .C1(n17749), .C2(n20846), .A(
        n17748), .ZN(n18151) );
  NAND2_X1 U19715 ( .A1(n18152), .A2(n18151), .ZN(n18150) );
  NAND2_X1 U19716 ( .A1(n17753), .A2(n17754), .ZN(n17755) );
  NAND2_X1 U19717 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18132), .ZN(
        n18131) );
  NAND2_X1 U19718 ( .A1(n17758), .A2(n17757), .ZN(n17759) );
  NAND2_X1 U19719 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18108), .ZN(
        n18107) );
  INV_X1 U19720 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20903) );
  NAND2_X1 U19721 ( .A1(n17763), .A2(n17760), .ZN(n17764) );
  NAND2_X1 U19722 ( .A1(n17763), .A2(n17762), .ZN(n17761) );
  NAND2_X1 U19723 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18076), .ZN(
        n18075) );
  AOI22_X2 U19724 ( .A1(n20812), .A2(n18088), .B1(n18161), .B2(n20925), .ZN(
        n18074) );
  INV_X1 U19725 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17830) );
  INV_X1 U19726 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21214) );
  NOR2_X1 U19727 ( .A1(n21214), .A2(n21195), .ZN(n20927) );
  NAND3_X1 U19728 ( .A1(n20927), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20934) );
  NOR2_X1 U19729 ( .A1(n17830), .A2(n20934), .ZN(n20948) );
  NAND2_X1 U19730 ( .A1(n20948), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20969) );
  NOR2_X1 U19731 ( .A1(n17794), .A2(n20969), .ZN(n20994) );
  NAND2_X1 U19732 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21157) );
  INV_X1 U19733 ( .A(n20948), .ZN(n20947) );
  NAND2_X1 U19734 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18025), .ZN(
        n18024) );
  NAND2_X1 U19735 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18033), .ZN(
        n20964) );
  AOI22_X1 U19736 ( .A1(n21151), .A2(n18161), .B1(n20976), .B2(n18088), .ZN(
        n17810) );
  INV_X1 U19737 ( .A(n17810), .ZN(n17795) );
  AOI21_X1 U19738 ( .B1(n18014), .B2(n21157), .A(n17795), .ZN(n18018) );
  INV_X1 U19739 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17787) );
  NAND2_X1 U19740 ( .A1(n18129), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18117) );
  NAND4_X1 U19741 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18040) );
  NAND2_X1 U19742 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17833) );
  NAND2_X1 U19743 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17804) );
  NAND2_X1 U19744 ( .A1(n18011), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17767) );
  NOR2_X1 U19745 ( .A1(n17767), .A2(n20130), .ZN(n20355) );
  INV_X1 U19746 ( .A(n17877), .ZN(n18167) );
  INV_X1 U19747 ( .A(n18128), .ZN(n17812) );
  AOI21_X1 U19748 ( .B1(n17812), .B2(n17767), .A(n18156), .ZN(n18022) );
  OAI21_X1 U19749 ( .B1(n20355), .B2(n18167), .A(n18022), .ZN(n17785) );
  NOR3_X1 U19750 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17966), .A3(
        n17767), .ZN(n17786) );
  INV_X1 U19751 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21166) );
  NAND2_X1 U19752 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20353) );
  OAI21_X1 U19753 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20355), .A(
        n20353), .ZN(n20358) );
  OAI22_X1 U19754 ( .A1(n21199), .A2(n21166), .B1(n17894), .B2(n20358), .ZN(
        n17768) );
  AOI211_X1 U19755 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17785), .A(
        n17786), .B(n17768), .ZN(n17778) );
  NAND2_X1 U19756 ( .A1(n18051), .A2(n17787), .ZN(n17844) );
  INV_X1 U19757 ( .A(n17844), .ZN(n17867) );
  AOI21_X1 U19758 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17976), .A(
        n17867), .ZN(n17776) );
  AOI22_X1 U19759 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18051), .B1(
        n17976), .B2(n21208), .ZN(n18078) );
  NOR2_X1 U19760 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18061) );
  INV_X1 U19761 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21184) );
  AND2_X1 U19762 ( .A1(n18061), .A2(n21184), .ZN(n17770) );
  NOR2_X1 U19763 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17771) );
  INV_X1 U19764 ( .A(n17774), .ZN(n17773) );
  INV_X1 U19765 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21177) );
  INV_X1 U19766 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21170) );
  NOR2_X1 U19767 ( .A1(n17775), .A2(n17774), .ZN(n17800) );
  OR2_X1 U19768 ( .A1(n21157), .A2(n17800), .ZN(n17779) );
  NAND2_X1 U19769 ( .A1(n17902), .A2(n17779), .ZN(n17845) );
  XNOR2_X1 U19770 ( .A(n17776), .B(n17845), .ZN(n21164) );
  NOR2_X1 U19771 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21157), .ZN(
        n21163) );
  AOI22_X1 U19772 ( .A1(n18086), .A2(n21164), .B1(n18014), .B2(n21163), .ZN(
        n17777) );
  OAI211_X1 U19773 ( .C1(n18018), .C2(n17787), .A(n17778), .B(n17777), .ZN(
        P3_U2812) );
  NOR3_X1 U19774 ( .A1(n18051), .A2(n17787), .A3(n17779), .ZN(n17866) );
  NOR2_X1 U19775 ( .A1(n17844), .A2(n17845), .ZN(n17850) );
  NOR2_X1 U19776 ( .A1(n17866), .A2(n17850), .ZN(n17780) );
  XOR2_X1 U19777 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17780), .Z(
        n21140) );
  INV_X1 U19778 ( .A(n20353), .ZN(n17781) );
  NOR2_X1 U19779 ( .A1(n17863), .A2(n20130), .ZN(n20383) );
  INV_X1 U19780 ( .A(n20383), .ZN(n17861) );
  OAI21_X1 U19781 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17781), .A(
        n17861), .ZN(n20370) );
  NAND2_X1 U19782 ( .A1(n10990), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21137) );
  NAND3_X1 U19783 ( .A1(n17782), .A2(n11157), .A3(n17923), .ZN(n17783) );
  OAI211_X1 U19784 ( .C1(n17894), .C2(n20370), .A(n21137), .B(n17783), .ZN(
        n17784) );
  AOI221_X1 U19785 ( .B1(n17786), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(
        n17785), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17784), .ZN(
        n17789) );
  OR2_X1 U19786 ( .A1(n21157), .A2(n17787), .ZN(n20824) );
  INV_X1 U19787 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21136) );
  OR2_X1 U19788 ( .A1(n20824), .A2(n21136), .ZN(n20818) );
  NOR2_X1 U19789 ( .A1(n20976), .A2(n20818), .ZN(n21131) );
  NOR2_X1 U19790 ( .A1(n21151), .A2(n20818), .ZN(n21129) );
  OAI22_X1 U19791 ( .A1(n21131), .A2(n18034), .B1(n21129), .B2(n18171), .ZN(
        n17869) );
  NOR2_X1 U19792 ( .A1(n20824), .A2(n17958), .ZN(n17916) );
  AOI22_X1 U19793 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17869), .B1(
        n17916), .B2(n21136), .ZN(n17788) );
  OAI211_X1 U19794 ( .C1(n21140), .C2(n18035), .A(n17789), .B(n17788), .ZN(
        P3_U2811) );
  NOR2_X1 U19795 ( .A1(n17966), .A2(n17790), .ZN(n17805) );
  INV_X1 U19796 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20313) );
  NOR2_X1 U19797 ( .A1(n17790), .A2(n20130), .ZN(n20308) );
  AOI21_X1 U19798 ( .B1(n17812), .B2(n17790), .A(n18156), .ZN(n18028) );
  OAI21_X1 U19799 ( .B1(n20308), .B2(n18167), .A(n18028), .ZN(n17803) );
  INV_X1 U19800 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20322) );
  NAND2_X1 U19801 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20308), .ZN(
        n20310) );
  OAI21_X1 U19802 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20308), .A(
        n20310), .ZN(n20311) );
  OAI22_X1 U19803 ( .A1(n21199), .A2(n20322), .B1(n17894), .B2(n20311), .ZN(
        n17791) );
  AOI221_X1 U19804 ( .B1(n17805), .B2(n20313), .C1(n17803), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17791), .ZN(n17799) );
  NOR2_X1 U19805 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18024), .ZN(
        n20973) );
  NAND2_X1 U19806 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20813) );
  INV_X1 U19807 ( .A(n20813), .ZN(n20921) );
  AND3_X1 U19808 ( .A1(n17792), .A2(n17976), .A3(n20921), .ZN(n18064) );
  NAND2_X1 U19809 ( .A1(n20948), .A2(n18064), .ZN(n18030) );
  NAND2_X1 U19810 ( .A1(n18045), .A2(n11076), .ZN(n18031) );
  INV_X1 U19811 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20963) );
  AOI22_X1 U19812 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18030), .B1(
        n18031), .B2(n20963), .ZN(n17793) );
  XNOR2_X1 U19813 ( .A(n17794), .B(n17793), .ZN(n20974) );
  AOI22_X1 U19814 ( .A1(n18161), .A2(n20973), .B1(n18086), .B2(n20974), .ZN(
        n17798) );
  OAI21_X1 U19815 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17796), .A(
        n17795), .ZN(n17797) );
  NAND3_X1 U19816 ( .A1(n17799), .A2(n17798), .A3(n17797), .ZN(P3_U2815) );
  AOI22_X1 U19817 ( .A1(n17976), .A2(n21177), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18051), .ZN(n17801) );
  XNOR2_X1 U19818 ( .A(n17800), .B(n17801), .ZN(n21179) );
  INV_X1 U19819 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21181) );
  INV_X1 U19820 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17802) );
  AND2_X1 U19821 ( .A1(n18011), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20336) );
  AOI21_X1 U19822 ( .B1(n17802), .B2(n20310), .A(n20336), .ZN(n20330) );
  AOI22_X1 U19823 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17803), .B1(
        n18006), .B2(n20330), .ZN(n17807) );
  OAI211_X1 U19824 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17805), .B(n17804), .ZN(n17806) );
  OAI211_X1 U19825 ( .C1(n21181), .C2(n21199), .A(n17807), .B(n17806), .ZN(
        n17808) );
  AOI21_X1 U19826 ( .B1(n18086), .B2(n21179), .A(n17808), .ZN(n17809) );
  OAI221_X1 U19827 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17958), 
        .C1(n21177), .C2(n17810), .A(n17809), .ZN(P3_U2814) );
  NOR2_X1 U19828 ( .A1(n17811), .A2(n20130), .ZN(n18042) );
  NAND2_X1 U19829 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18042), .ZN(
        n17824) );
  OAI21_X1 U19830 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18042), .A(
        n17824), .ZN(n20272) );
  NOR2_X1 U19831 ( .A1(n17966), .A2(n17811), .ZN(n17834) );
  INV_X1 U19832 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20276) );
  AOI21_X1 U19833 ( .B1(n17812), .B2(n17811), .A(n17877), .ZN(n17813) );
  OAI21_X1 U19834 ( .B1(n18042), .B2(n17813), .A(n18166), .ZN(n17825) );
  NAND2_X1 U19835 ( .A1(n10990), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n20944) );
  INV_X1 U19836 ( .A(n20944), .ZN(n17814) );
  AOI221_X1 U19837 ( .B1(n17834), .B2(n20276), .C1(n17825), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17814), .ZN(n17823) );
  NAND2_X1 U19838 ( .A1(n20927), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20933) );
  NOR2_X1 U19839 ( .A1(n17815), .A2(n20933), .ZN(n17816) );
  MUX2_X1 U19840 ( .A(n17816), .B(n11329), .S(n18051), .Z(n17817) );
  XOR2_X1 U19841 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17817), .Z(
        n20943) );
  NOR2_X1 U19842 ( .A1(n18074), .A2(n20933), .ZN(n17820) );
  NOR2_X1 U19843 ( .A1(n21152), .A2(n20934), .ZN(n20936) );
  INV_X1 U19844 ( .A(n20936), .ZN(n17818) );
  INV_X1 U19845 ( .A(n20934), .ZN(n17829) );
  NAND2_X1 U19846 ( .A1(n17829), .A2(n20925), .ZN(n20938) );
  AOI22_X1 U19847 ( .A1(n18088), .A2(n17818), .B1(n18161), .B2(n20938), .ZN(
        n17831) );
  INV_X1 U19848 ( .A(n17831), .ZN(n17819) );
  MUX2_X1 U19849 ( .A(n17820), .B(n17819), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17821) );
  AOI21_X1 U19850 ( .B1(n18086), .B2(n20943), .A(n17821), .ZN(n17822) );
  OAI211_X1 U19851 ( .C1(n17894), .C2(n20272), .A(n17823), .B(n17822), .ZN(
        P3_U2818) );
  INV_X1 U19852 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20291) );
  AOI22_X1 U19853 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18027), .B1(
        n20291), .B2(n17824), .ZN(n20290) );
  AOI22_X1 U19854 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17825), .B1(
        n18006), .B2(n20290), .ZN(n17838) );
  INV_X1 U19855 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21185) );
  AOI22_X1 U19856 ( .A1(n17829), .A2(n18053), .B1(n18051), .B2(n21185), .ZN(
        n17826) );
  AOI21_X1 U19857 ( .B1(n17827), .B2(n18051), .A(n17826), .ZN(n17828) );
  XNOR2_X1 U19858 ( .A(n17828), .B(n17830), .ZN(n21183) );
  NAND2_X1 U19859 ( .A1(n17829), .A2(n17830), .ZN(n21194) );
  OAI22_X1 U19860 ( .A1(n18074), .A2(n21194), .B1(n17831), .B2(n17830), .ZN(
        n17832) );
  AOI21_X1 U19861 ( .B1(n18086), .B2(n21183), .A(n17832), .ZN(n17837) );
  NAND2_X1 U19862 ( .A1(n10990), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17836) );
  OAI211_X1 U19863 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17834), .B(n17833), .ZN(n17835) );
  NAND4_X1 U19864 ( .A1(n17838), .A2(n17837), .A3(n17836), .A4(n17835), .ZN(
        P3_U2817) );
  NAND2_X1 U19865 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20825) );
  INV_X1 U19866 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20826) );
  NOR2_X1 U19867 ( .A1(n20825), .A2(n20826), .ZN(n20983) );
  INV_X1 U19868 ( .A(n20983), .ZN(n20992) );
  NOR2_X1 U19869 ( .A1(n20824), .A2(n20992), .ZN(n17920) );
  NAND2_X1 U19870 ( .A1(n17920), .A2(n18014), .ZN(n17849) );
  INV_X1 U19871 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17841) );
  NAND3_X1 U19872 ( .A1(n11073), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17839) );
  NOR2_X1 U19873 ( .A1(n17882), .A2(n20130), .ZN(n17878) );
  AOI21_X1 U19874 ( .B1(n17841), .B2(n17839), .A(n17878), .ZN(n20409) );
  INV_X1 U19875 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20398) );
  NAND2_X1 U19876 ( .A1(n11073), .A2(n17923), .ZN(n17856) );
  AOI221_X1 U19877 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17841), .C2(n20398), .A(
        n17856), .ZN(n17843) );
  AOI21_X1 U19878 ( .B1(n17877), .B2(n17861), .A(n18156), .ZN(n17840) );
  OAI21_X1 U19879 ( .B1(n11073), .B2(n18128), .A(n17840), .ZN(n17865) );
  AOI21_X1 U19880 ( .B1(n17879), .B2(n17862), .A(n17865), .ZN(n17855) );
  INV_X1 U19881 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20420) );
  OAI22_X1 U19882 ( .A1(n17855), .A2(n17841), .B1(n21199), .B2(n20420), .ZN(
        n17842) );
  AOI211_X1 U19883 ( .C1(n20409), .C2(n18006), .A(n17843), .B(n17842), .ZN(
        n17848) );
  INV_X1 U19884 ( .A(n17920), .ZN(n17959) );
  NOR2_X1 U19885 ( .A1(n17959), .A2(n21151), .ZN(n20822) );
  NOR2_X1 U19886 ( .A1(n17959), .A2(n20976), .ZN(n20821) );
  OAI22_X1 U19887 ( .A1(n20822), .A2(n18171), .B1(n20821), .B2(n18034), .ZN(
        n17858) );
  NOR4_X1 U19888 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n17844), .ZN(n17885) );
  NAND3_X1 U19889 ( .A1(n20983), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17845), .ZN(n17903) );
  INV_X1 U19890 ( .A(n17903), .ZN(n17846) );
  OAI21_X1 U19891 ( .B1(n17885), .B2(n17846), .A(n17902), .ZN(n17886) );
  XNOR2_X1 U19892 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17886), .ZN(
        n20988) );
  AOI22_X1 U19893 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17858), .B1(
        n18086), .B2(n20988), .ZN(n17847) );
  OAI211_X1 U19894 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17849), .A(
        n17848), .B(n17847), .ZN(P3_U2808) );
  INV_X1 U19895 ( .A(n20825), .ZN(n17852) );
  NOR2_X1 U19896 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U19897 ( .A1(n17852), .A2(n17866), .B1(n17851), .B2(n17850), .ZN(
        n17853) );
  XNOR2_X1 U19898 ( .A(n17853), .B(n20826), .ZN(n20832) );
  NAND2_X1 U19899 ( .A1(n11073), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17854) );
  XNOR2_X1 U19900 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n17854), .ZN(
        n20396) );
  NAND2_X1 U19901 ( .A1(n10990), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n20830) );
  OAI221_X1 U19902 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17856), .C1(
        n20398), .C2(n17855), .A(n20830), .ZN(n17857) );
  AOI21_X1 U19903 ( .B1(n18006), .B2(n20396), .A(n17857), .ZN(n17860) );
  NOR2_X1 U19904 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n20825), .ZN(
        n20829) );
  AOI22_X1 U19905 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17858), .B1(
        n20829), .B2(n17916), .ZN(n17859) );
  OAI211_X1 U19906 ( .C1(n20832), .C2(n18035), .A(n17860), .B(n17859), .ZN(
        P3_U2809) );
  AOI22_X1 U19907 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11073), .B1(
        n17862), .B2(n17861), .ZN(n20386) );
  NAND2_X1 U19908 ( .A1(n17894), .A2(n17967), .ZN(n18015) );
  OAI21_X1 U19909 ( .B1(n17863), .B2(n18751), .A(n17862), .ZN(n17864) );
  AOI22_X1 U19910 ( .A1(n20386), .A2(n18015), .B1(n17865), .B2(n17864), .ZN(
        n17873) );
  OAI221_X1 U19911 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17867), 
        .C1(n21136), .C2(n17866), .A(n17902), .ZN(n17868) );
  XNOR2_X1 U19912 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17868), .ZN(
        n21143) );
  NOR2_X1 U19913 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21136), .ZN(
        n21141) );
  AOI22_X1 U19914 ( .A1(n18086), .A2(n21143), .B1(n17916), .B2(n21141), .ZN(
        n17872) );
  NAND2_X1 U19915 ( .A1(n10990), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17871) );
  NAND2_X1 U19916 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17869), .ZN(
        n17870) );
  NAND4_X1 U19917 ( .A1(n17873), .A2(n17872), .A3(n17871), .A4(n17870), .ZN(
        P3_U2810) );
  NAND3_X1 U19918 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17920), .ZN(n17900) );
  NOR2_X1 U19919 ( .A1(n17900), .A2(n21151), .ZN(n21110) );
  NOR2_X1 U19920 ( .A1(n21110), .A2(n18171), .ZN(n17875) );
  NOR2_X1 U19921 ( .A1(n17900), .A2(n20976), .ZN(n21109) );
  NOR2_X1 U19922 ( .A1(n21109), .A2(n18034), .ZN(n17874) );
  AOI22_X1 U19923 ( .A1(n20822), .A2(n17875), .B1(n20821), .B2(n17874), .ZN(
        n17890) );
  INV_X1 U19924 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21027) );
  INV_X1 U19925 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20429) );
  NAND2_X1 U19926 ( .A1(n17892), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17911) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17878), .A(
        n17911), .ZN(n17876) );
  INV_X1 U19928 ( .A(n17876), .ZN(n20423) );
  INV_X1 U19929 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20425) );
  NOR2_X1 U19930 ( .A1(n21199), .A2(n20425), .ZN(n21116) );
  NOR2_X1 U19931 ( .A1(n17892), .A2(n18751), .ZN(n17880) );
  AOI211_X1 U19932 ( .C1(n17877), .C2(n17911), .A(n18156), .B(n17880), .ZN(
        n17912) );
  AOI21_X1 U19933 ( .B1(n17879), .B2(n17878), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17883) );
  INV_X1 U19934 ( .A(n17880), .ZN(n17881) );
  OAI22_X1 U19935 ( .A1(n17912), .A2(n17883), .B1(n17882), .B2(n17881), .ZN(
        n17884) );
  AOI211_X1 U19936 ( .C1(n20423), .C2(n18006), .A(n21116), .B(n17884), .ZN(
        n17889) );
  OAI22_X1 U19937 ( .A1(n21110), .A2(n18171), .B1(n21109), .B2(n18034), .ZN(
        n17917) );
  NAND2_X1 U19938 ( .A1(n17885), .A2(n21027), .ZN(n17899) );
  AOI221_X1 U19939 ( .B1(n21027), .B2(n17899), .C1(n18051), .C2(n17899), .A(
        n17886), .ZN(n17887) );
  XOR2_X1 U19940 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17887), .Z(
        n21117) );
  AOI22_X1 U19941 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17917), .B1(
        n18086), .B2(n21117), .ZN(n17888) );
  OAI211_X1 U19942 ( .C1(n17890), .C2(n21027), .A(n17889), .B(n17888), .ZN(
        P3_U2807) );
  NAND2_X1 U19943 ( .A1(n21110), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17891) );
  INV_X1 U19944 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21012) );
  XNOR2_X1 U19945 ( .A(n17891), .B(n21012), .ZN(n21007) );
  INV_X1 U19946 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17895) );
  INV_X1 U19947 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20446) );
  NAND2_X1 U19948 ( .A1(n17892), .A2(n17923), .ZN(n17913) );
  AOI221_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n17895), .C2(n20446), .A(
        n17913), .ZN(n17897) );
  NOR2_X1 U19950 ( .A1(n20446), .A2(n17911), .ZN(n17910) );
  NOR2_X1 U19951 ( .A1(n17952), .A2(n20130), .ZN(n17949) );
  INV_X1 U19952 ( .A(n17949), .ZN(n17893) );
  OAI21_X1 U19953 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17910), .A(
        n17893), .ZN(n20451) );
  OAI22_X1 U19954 ( .A1(n17912), .A2(n17895), .B1(n17894), .B2(n20451), .ZN(
        n17896) );
  AOI211_X1 U19955 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n10990), .A(n17897), 
        .B(n17896), .ZN(n17907) );
  NAND2_X1 U19956 ( .A1(n21109), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17898) );
  XNOR2_X1 U19957 ( .A(n17898), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n20999) );
  OAI22_X1 U19958 ( .A1(n17800), .A2(n17900), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17899), .ZN(n17901) );
  NAND2_X1 U19959 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17915) );
  INV_X1 U19960 ( .A(n17931), .ZN(n17904) );
  AOI21_X1 U19961 ( .B1(n17976), .B2(n17932), .A(n17904), .ZN(n17905) );
  XNOR2_X1 U19962 ( .A(n17905), .B(n21012), .ZN(n21003) );
  AOI22_X1 U19963 ( .A1(n18088), .A2(n20999), .B1(n18086), .B2(n21003), .ZN(
        n17906) );
  OAI211_X1 U19964 ( .C1(n18171), .C2(n21007), .A(n17907), .B(n17906), .ZN(
        P3_U2805) );
  AOI21_X1 U19965 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17909), .A(
        n17908), .ZN(n21127) );
  AOI21_X1 U19966 ( .B1(n20446), .B2(n17911), .A(n17910), .ZN(n20442) );
  NAND2_X1 U19967 ( .A1(n10990), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n21125) );
  OAI221_X1 U19968 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17913), .C1(
        n20446), .C2(n17912), .A(n21125), .ZN(n17914) );
  AOI21_X1 U19969 ( .B1(n18006), .B2(n20442), .A(n17914), .ZN(n17919) );
  NOR3_X1 U19970 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n20992), .A3(
        n17915), .ZN(n21123) );
  AOI22_X1 U19971 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17917), .B1(
        n17916), .B2(n21123), .ZN(n17918) );
  OAI211_X1 U19972 ( .C1(n21127), .C2(n18035), .A(n17919), .B(n17918), .ZN(
        P3_U2806) );
  NAND2_X1 U19973 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21041) );
  NAND2_X1 U19974 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20991) );
  NOR2_X1 U19975 ( .A1(n21041), .A2(n20991), .ZN(n21028) );
  INV_X1 U19976 ( .A(n21028), .ZN(n21022) );
  NAND2_X1 U19977 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17920), .ZN(
        n20997) );
  OR2_X1 U19978 ( .A1(n21022), .A2(n20997), .ZN(n21051) );
  NOR2_X1 U19979 ( .A1(n21051), .A2(n17958), .ZN(n17938) );
  INV_X1 U19980 ( .A(n17938), .ZN(n17987) );
  INV_X1 U19981 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21057) );
  NAND2_X1 U19982 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21057), .ZN(
        n21092) );
  INV_X1 U19983 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17922) );
  NAND2_X1 U19984 ( .A1(n17939), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17927) );
  NOR2_X1 U19985 ( .A1(n17927), .A2(n20130), .ZN(n17940) );
  INV_X1 U19986 ( .A(n17940), .ZN(n17921) );
  NAND2_X1 U19987 ( .A1(n18002), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18004) );
  INV_X1 U19988 ( .A(n18004), .ZN(n17970) );
  AOI21_X1 U19989 ( .B1(n17922), .B2(n17921), .A(n17970), .ZN(n20491) );
  INV_X1 U19990 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21029) );
  OAI22_X1 U19991 ( .A1(n17989), .A2(n18171), .B1(n21046), .B2(n18034), .ZN(
        n17957) );
  NOR2_X1 U19992 ( .A1(n21029), .A2(n17957), .ZN(n17947) );
  AOI211_X1 U19993 ( .C1(n18034), .C2(n18171), .A(n17947), .B(n21057), .ZN(
        n17929) );
  NAND2_X1 U19994 ( .A1(n17922), .A2(n17923), .ZN(n17926) );
  NAND2_X1 U19995 ( .A1(n10990), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21103) );
  INV_X1 U19996 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20480) );
  AND3_X1 U19997 ( .A1(n20480), .A2(n17923), .A3(n17939), .ZN(n17941) );
  OAI22_X1 U19998 ( .A1(n17939), .A2(n18128), .B1(n17949), .B2(n18167), .ZN(
        n17924) );
  NOR2_X1 U19999 ( .A1(n18156), .A2(n17924), .ZN(n17951) );
  OAI21_X1 U20000 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17967), .A(
        n17951), .ZN(n17943) );
  OAI21_X1 U20001 ( .B1(n17941), .B2(n17943), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17925) );
  OAI211_X1 U20002 ( .C1(n17927), .C2(n17926), .A(n21103), .B(n17925), .ZN(
        n17928) );
  AOI211_X1 U20003 ( .C1(n18006), .C2(n20491), .A(n17929), .B(n17928), .ZN(
        n17937) );
  NOR2_X1 U20004 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17976), .ZN(
        n17973) );
  AOI21_X1 U20005 ( .B1(n17976), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17973), .ZN(n21101) );
  INV_X1 U20006 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17955) );
  INV_X1 U20007 ( .A(n21041), .ZN(n17933) );
  INV_X1 U20008 ( .A(n17974), .ZN(n21102) );
  NOR2_X1 U20009 ( .A1(n17934), .A2(n21029), .ZN(n17975) );
  NOR2_X1 U20010 ( .A1(n17974), .A2(n17975), .ZN(n17942) );
  OAI211_X1 U20011 ( .C1(n21101), .C2(n17935), .A(n18086), .B(n21089), .ZN(
        n17936) );
  OAI211_X1 U20012 ( .C1(n17987), .C2(n21092), .A(n17937), .B(n17936), .ZN(
        P3_U2802) );
  NOR2_X1 U20013 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17938), .ZN(
        n17946) );
  NAND2_X1 U20014 ( .A1(n17939), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17948) );
  AOI21_X1 U20015 ( .B1(n20480), .B2(n17948), .A(n17940), .ZN(n20478) );
  INV_X1 U20016 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20487) );
  NOR2_X1 U20017 ( .A1(n21199), .A2(n20487), .ZN(n21033) );
  AOI211_X1 U20018 ( .C1(n18006), .C2(n20478), .A(n21033), .B(n17941), .ZN(
        n17945) );
  AOI22_X1 U20019 ( .A1(n18086), .A2(n21034), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17943), .ZN(n17944) );
  OAI211_X1 U20020 ( .C1(n17947), .C2(n17946), .A(n17945), .B(n17944), .ZN(
        P3_U2803) );
  OAI21_X1 U20021 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17949), .A(
        n17948), .ZN(n17950) );
  INV_X1 U20022 ( .A(n17950), .ZN(n20468) );
  AOI221_X1 U20023 ( .B1(n17952), .B2(n20473), .C1(n18751), .C2(n20473), .A(
        n17951), .ZN(n17953) );
  AOI221_X1 U20024 ( .B1(n18006), .B2(n20468), .C1(n17879), .C2(n20468), .A(
        n17953), .ZN(n17962) );
  OAI21_X1 U20025 ( .B1(n17956), .B2(n17955), .A(n17954), .ZN(n21009) );
  AOI22_X1 U20026 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17957), .B1(
        n18086), .B2(n21009), .ZN(n17961) );
  INV_X1 U20027 ( .A(n20991), .ZN(n20998) );
  NAND3_X1 U20028 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n20998), .ZN(n21016) );
  NAND2_X1 U20029 ( .A1(n10990), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21019) );
  NAND4_X1 U20030 ( .A1(n17962), .A2(n17961), .A3(n17960), .A4(n21019), .ZN(
        P3_U2804) );
  INV_X1 U20031 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21059) );
  INV_X1 U20032 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17977) );
  NOR2_X1 U20033 ( .A1(n21059), .A2(n17977), .ZN(n21072) );
  NAND2_X1 U20034 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21040) );
  NOR2_X1 U20035 ( .A1(n21040), .A2(n21013), .ZN(n21095) );
  NAND2_X1 U20036 ( .A1(n21072), .A2(n21095), .ZN(n17963) );
  XOR2_X1 U20037 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n17963), .Z(
        n21079) );
  NAND2_X1 U20038 ( .A1(n18002), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17968) );
  NAND2_X1 U20039 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18003), .ZN(
        n17965) );
  INV_X1 U20040 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20530) );
  NOR2_X1 U20041 ( .A1(n21199), .A2(n20530), .ZN(n21083) );
  OR2_X1 U20042 ( .A1(n17968), .A2(n17966), .ZN(n17986) );
  XOR2_X1 U20043 ( .A(n17964), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17971) );
  NOR2_X1 U20044 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17967), .ZN(
        n18007) );
  AOI21_X1 U20045 ( .B1(n19011), .B2(n17968), .A(n18156), .ZN(n17969) );
  OAI21_X1 U20046 ( .B1(n17970), .B2(n18167), .A(n17969), .ZN(n18001) );
  NOR2_X1 U20047 ( .A1(n18007), .A2(n18001), .ZN(n17984) );
  OAI22_X1 U20048 ( .A1(n17986), .A2(n17971), .B1(n17984), .B2(n17964), .ZN(
        n17972) );
  AOI211_X1 U20049 ( .C1(n20354), .C2(n18006), .A(n21083), .B(n17972), .ZN(
        n17982) );
  NAND3_X1 U20050 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17976), .A3(
        n17975), .ZN(n21100) );
  OAI33_X1 U20051 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n17995), .B1(n17977), .B2(
        n21100), .B3(n21059), .ZN(n17979) );
  XNOR2_X1 U20052 ( .A(n17979), .B(n17978), .ZN(n21082) );
  INV_X1 U20053 ( .A(n21046), .ZN(n21023) );
  NOR2_X1 U20054 ( .A1(n21040), .A2(n21023), .ZN(n21096) );
  NAND2_X1 U20055 ( .A1(n21072), .A2(n21096), .ZN(n17980) );
  XNOR2_X1 U20056 ( .A(n17980), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n21075) );
  AOI22_X1 U20057 ( .A1(n18086), .A2(n21082), .B1(n18088), .B2(n21075), .ZN(
        n17981) );
  OAI211_X1 U20058 ( .C1(n21079), .C2(n18171), .A(n17982), .B(n17981), .ZN(
        P3_U2799) );
  AOI22_X1 U20059 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21100), .B1(
        n17995), .B2(n21059), .ZN(n17983) );
  XNOR2_X1 U20060 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n17983), .ZN(
        n21071) );
  XOR2_X1 U20061 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n18003), .Z(
        n20526) );
  INV_X1 U20062 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17985) );
  NAND2_X1 U20063 ( .A1(n10990), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21069) );
  OAI221_X1 U20064 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17986), .C1(
        n17985), .C2(n17984), .A(n21069), .ZN(n17993) );
  NOR2_X1 U20065 ( .A1(n21040), .A2(n21059), .ZN(n21065) );
  INV_X1 U20066 ( .A(n21065), .ZN(n17988) );
  NOR2_X1 U20067 ( .A1(n17988), .A2(n17987), .ZN(n17991) );
  NAND2_X1 U20068 ( .A1(n17989), .A2(n21065), .ZN(n21047) );
  AOI21_X1 U20069 ( .B1(n21046), .B2(n21065), .A(n18034), .ZN(n18000) );
  AOI21_X1 U20070 ( .B1(n18161), .B2(n21047), .A(n18000), .ZN(n17998) );
  INV_X1 U20071 ( .A(n17998), .ZN(n17990) );
  MUX2_X1 U20072 ( .A(n17991), .B(n17990), .S(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n17992) );
  AOI211_X1 U20073 ( .C1(n18006), .C2(n20526), .A(n17993), .B(n17992), .ZN(
        n17994) );
  OAI21_X1 U20074 ( .B1(n21071), .B2(n18035), .A(n17994), .ZN(P3_U2800) );
  AOI21_X1 U20075 ( .B1(n21095), .B2(n18161), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U20076 ( .A1(n17995), .A2(n21100), .ZN(n17996) );
  XNOR2_X1 U20077 ( .A(n17996), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21063) );
  OAI22_X1 U20078 ( .A1(n17998), .A2(n17997), .B1(n21063), .B2(n18035), .ZN(
        n17999) );
  AOI21_X1 U20079 ( .B1(n21096), .B2(n18000), .A(n17999), .ZN(n18010) );
  NAND2_X1 U20080 ( .A1(n10990), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21061) );
  OAI221_X1 U20081 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18002), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19011), .A(n18001), .ZN(
        n18009) );
  INV_X1 U20082 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18005) );
  AOI21_X1 U20083 ( .B1(n18005), .B2(n18004), .A(n18003), .ZN(n20508) );
  OAI21_X1 U20084 ( .B1(n18007), .B2(n18006), .A(n20508), .ZN(n18008) );
  NAND4_X1 U20085 ( .A1(n18010), .A2(n21061), .A3(n18009), .A4(n18008), .ZN(
        P3_U2801) );
  AOI21_X1 U20086 ( .B1(n18011), .B2(n19011), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18023) );
  OAI21_X1 U20087 ( .B1(n18013), .B2(n21170), .A(n18012), .ZN(n21168) );
  AOI21_X1 U20088 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18014), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18017) );
  INV_X1 U20089 ( .A(n20355), .ZN(n18016) );
  OAI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20336), .A(
        n18016), .ZN(n20338) );
  OAI22_X1 U20091 ( .A1(n18018), .A2(n18017), .B1(n18153), .B2(n20338), .ZN(
        n18019) );
  AOI21_X1 U20092 ( .B1(n18086), .B2(n21168), .A(n18019), .ZN(n18021) );
  NAND2_X1 U20093 ( .A1(n10990), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18020) );
  OAI211_X1 U20094 ( .C1(n18023), .C2(n18022), .A(n18021), .B(n18020), .ZN(
        P3_U2813) );
  OAI21_X1 U20095 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18025), .A(
        n18024), .ZN(n20956) );
  INV_X1 U20096 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18026) );
  NAND2_X1 U20097 ( .A1(n18027), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20280) );
  AOI21_X1 U20098 ( .B1(n18026), .B2(n20280), .A(n20308), .ZN(n20299) );
  AOI21_X1 U20099 ( .B1(n18027), .B2(n19011), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18029) );
  NAND2_X1 U20100 ( .A1(n10990), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n20961) );
  OAI21_X1 U20101 ( .B1(n18029), .B2(n18028), .A(n20961), .ZN(n18037) );
  NAND2_X1 U20102 ( .A1(n18031), .A2(n18030), .ZN(n18032) );
  XNOR2_X1 U20103 ( .A(n18032), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20957) );
  OAI21_X1 U20104 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18033), .A(
        n20964), .ZN(n20954) );
  OAI22_X1 U20105 ( .A1(n20957), .A2(n18035), .B1(n18034), .B2(n20954), .ZN(
        n18036) );
  AOI211_X1 U20106 ( .C1(n20299), .C2(n18015), .A(n18037), .B(n18036), .ZN(
        n18038) );
  OAI21_X1 U20107 ( .B1(n18171), .B2(n20956), .A(n18038), .ZN(P3_U2816) );
  AOI22_X1 U20108 ( .A1(n18161), .A2(n18039), .B1(n18088), .B2(n21152), .ZN(
        n18073) );
  NAND2_X1 U20109 ( .A1(n18166), .A2(n18128), .ZN(n18162) );
  INV_X1 U20110 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20263) );
  NAND3_X1 U20111 ( .A1(n18103), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19011), .ZN(n18094) );
  NOR2_X1 U20112 ( .A1(n18040), .A2(n18094), .ZN(n18058) );
  NOR2_X1 U20113 ( .A1(n20263), .A2(n18058), .ZN(n18044) );
  NAND2_X1 U20114 ( .A1(n18041), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18056) );
  INV_X1 U20115 ( .A(n18056), .ZN(n20254) );
  INV_X1 U20116 ( .A(n18042), .ZN(n20269) );
  OAI21_X1 U20117 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20254), .A(
        n20269), .ZN(n20256) );
  INV_X1 U20118 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20278) );
  OAI22_X1 U20119 ( .A1(n18153), .A2(n20256), .B1(n21199), .B2(n20278), .ZN(
        n18043) );
  AOI221_X1 U20120 ( .B1(n18162), .B2(n18044), .C1(n20263), .C2(n18058), .A(
        n18043), .ZN(n18050) );
  AND2_X1 U20121 ( .A1(n21208), .A2(n18045), .ZN(n18065) );
  AOI22_X1 U20122 ( .A1(n20927), .A2(n18064), .B1(n18061), .B2(n18065), .ZN(
        n18046) );
  XNOR2_X1 U20123 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18046), .ZN(
        n20923) );
  INV_X1 U20124 ( .A(n18074), .ZN(n18048) );
  NAND2_X1 U20125 ( .A1(n20927), .A2(n21184), .ZN(n20932) );
  OAI21_X1 U20126 ( .B1(n20927), .B2(n21184), .A(n20932), .ZN(n18047) );
  AOI22_X1 U20127 ( .A1(n18086), .A2(n20923), .B1(n18048), .B2(n18047), .ZN(
        n18049) );
  OAI211_X1 U20128 ( .C1(n18073), .C2(n21184), .A(n18050), .B(n18049), .ZN(
        P3_U2819) );
  AOI21_X1 U20129 ( .B1(n18051), .B2(n21214), .A(n18064), .ZN(n18052) );
  AOI21_X1 U20130 ( .B1(n21214), .B2(n18053), .A(n18052), .ZN(n18055) );
  AOI221_X1 U20131 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18064), .C1(
        n21214), .C2(n18065), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18054) );
  AOI21_X1 U20132 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18055), .A(
        n18054), .ZN(n21196) );
  INV_X1 U20133 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20246) );
  NOR2_X1 U20134 ( .A1(n21199), .A2(n20246), .ZN(n18060) );
  NAND2_X1 U20135 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18081) );
  INV_X1 U20136 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20229) );
  NOR3_X1 U20137 ( .A1(n18081), .A2(n20229), .A3(n18094), .ZN(n18070) );
  AOI21_X1 U20138 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18162), .A(
        n18070), .ZN(n18057) );
  INV_X1 U20139 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18093) );
  NOR3_X1 U20140 ( .A1(n18080), .A2(n18093), .A3(n20130), .ZN(n20217) );
  NAND2_X1 U20141 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20217), .ZN(
        n18079) );
  NOR2_X1 U20142 ( .A1(n20229), .A2(n18079), .ZN(n20228) );
  OAI21_X1 U20143 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20228), .A(
        n18056), .ZN(n20238) );
  OAI22_X1 U20144 ( .A1(n18058), .A2(n18057), .B1(n18153), .B2(n20238), .ZN(
        n18059) );
  AOI211_X1 U20145 ( .C1(n18086), .C2(n21196), .A(n18060), .B(n18059), .ZN(
        n18063) );
  OR3_X1 U20146 ( .A1(n20927), .A2(n18061), .A3(n18074), .ZN(n18062) );
  OAI211_X1 U20147 ( .C1(n18073), .C2(n21195), .A(n18063), .B(n18062), .ZN(
        P3_U2820) );
  NOR2_X1 U20148 ( .A1(n18065), .A2(n18064), .ZN(n18066) );
  XNOR2_X1 U20149 ( .A(n18066), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n21219) );
  INV_X1 U20150 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20245) );
  NOR2_X1 U20151 ( .A1(n21199), .A2(n20245), .ZN(n21218) );
  NOR2_X1 U20152 ( .A1(n18081), .A2(n18094), .ZN(n18067) );
  AOI21_X1 U20153 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18162), .A(
        n18067), .ZN(n18069) );
  AOI21_X1 U20154 ( .B1(n20229), .B2(n18079), .A(n20228), .ZN(n18068) );
  INV_X1 U20155 ( .A(n18068), .ZN(n20230) );
  OAI22_X1 U20156 ( .A1(n18070), .A2(n18069), .B1(n18153), .B2(n20230), .ZN(
        n18071) );
  AOI211_X1 U20157 ( .C1(n18086), .C2(n21219), .A(n21218), .B(n18071), .ZN(
        n18072) );
  OAI221_X1 U20158 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18074), .C1(
        n21214), .C2(n18073), .A(n18072), .ZN(P3_U2821) );
  OAI21_X1 U20159 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18076), .A(
        n18075), .ZN(n20919) );
  XOR2_X1 U20160 ( .A(n18078), .B(n18077), .Z(n20915) );
  INV_X1 U20161 ( .A(n20915), .ZN(n18087) );
  OAI21_X1 U20162 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20217), .A(
        n18079), .ZN(n20218) );
  INV_X1 U20163 ( .A(n18080), .ZN(n18092) );
  OAI21_X1 U20164 ( .B1(n18092), .B2(n18128), .A(n18166), .ZN(n18100) );
  AOI22_X1 U20165 ( .A1(n10990), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18100), .ZN(n18084) );
  NOR2_X1 U20166 ( .A1(n18080), .A2(n18093), .ZN(n18082) );
  OAI211_X1 U20167 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18082), .A(
        n19011), .B(n18081), .ZN(n18083) );
  OAI211_X1 U20168 ( .C1(n18153), .C2(n20218), .A(n18084), .B(n18083), .ZN(
        n18085) );
  AOI221_X1 U20169 ( .B1(n18088), .B2(n18087), .C1(n18086), .C2(n20915), .A(
        n18085), .ZN(n18089) );
  OAI21_X1 U20170 ( .B1(n18171), .B2(n20919), .A(n18089), .ZN(P3_U2822) );
  OAI21_X1 U20171 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18091), .A(
        n18090), .ZN(n20911) );
  NAND2_X1 U20172 ( .A1(n18092), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20192) );
  AOI21_X1 U20173 ( .B1(n18093), .B2(n20192), .A(n20217), .ZN(n20203) );
  OAI22_X1 U20174 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18094), .B1(
        n21199), .B2(n20898), .ZN(n18095) );
  AOI21_X1 U20175 ( .B1(n20203), .B2(n18015), .A(n18095), .ZN(n18102) );
  AOI21_X1 U20176 ( .B1(n18098), .B2(n18097), .A(n18096), .ZN(n18099) );
  XNOR2_X1 U20177 ( .A(n18099), .B(n20903), .ZN(n20900) );
  AOI22_X1 U20178 ( .A1(n18161), .A2(n20900), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18100), .ZN(n18101) );
  OAI211_X1 U20179 ( .C1(n18170), .C2(n20911), .A(n18102), .B(n18101), .ZN(
        P3_U2823) );
  AND2_X1 U20180 ( .A1(n18103), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18115) );
  OAI21_X1 U20181 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18115), .A(
        n20192), .ZN(n20200) );
  NAND2_X1 U20182 ( .A1(n18103), .A2(n19011), .ZN(n18109) );
  OAI21_X1 U20183 ( .B1(n18106), .B2(n18105), .A(n18104), .ZN(n20892) );
  OAI22_X1 U20184 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18109), .B1(
        n18170), .B2(n20892), .ZN(n18111) );
  OAI21_X1 U20185 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18108), .A(
        n18107), .ZN(n20891) );
  NAND2_X1 U20186 ( .A1(n18162), .A2(n18109), .ZN(n18116) );
  OAI22_X1 U20187 ( .A1(n18171), .A2(n20891), .B1(n11167), .B2(n18116), .ZN(
        n18110) );
  AOI211_X1 U20188 ( .C1(n10990), .C2(P3_REIP_REG_6__SCAN_IN), .A(n18111), .B(
        n18110), .ZN(n18112) );
  OAI21_X1 U20189 ( .B1(n18153), .B2(n20200), .A(n18112), .ZN(P3_U2824) );
  OAI21_X1 U20190 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18114), .A(
        n18113), .ZN(n20883) );
  INV_X1 U20191 ( .A(n18117), .ZN(n20169) );
  NAND2_X1 U20192 ( .A1(n20169), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18130) );
  AOI21_X1 U20193 ( .B1(n20180), .B2(n18130), .A(n18115), .ZN(n20176) );
  AOI221_X1 U20194 ( .B1(n18156), .B2(n20180), .C1(n18117), .C2(n20180), .A(
        n18116), .ZN(n18122) );
  INV_X1 U20195 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20179) );
  OAI21_X1 U20196 ( .B1(n18120), .B2(n18119), .A(n18118), .ZN(n20882) );
  OAI22_X1 U20197 ( .A1(n21199), .A2(n20179), .B1(n18171), .B2(n20882), .ZN(
        n18121) );
  AOI211_X1 U20198 ( .C1(n20176), .C2(n18015), .A(n18122), .B(n18121), .ZN(
        n18123) );
  OAI21_X1 U20199 ( .B1(n18170), .B2(n20883), .A(n18123), .ZN(P3_U2825) );
  OAI21_X1 U20200 ( .B1(n18126), .B2(n18125), .A(n18124), .ZN(n20869) );
  NOR2_X1 U20201 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18751), .ZN(
        n18127) );
  AOI22_X1 U20202 ( .A1(n10990), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18129), 
        .B2(n18127), .ZN(n18135) );
  OAI21_X1 U20203 ( .B1(n18129), .B2(n18128), .A(n18166), .ZN(n18145) );
  NAND2_X1 U20204 ( .A1(n18129), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18139) );
  INV_X1 U20205 ( .A(n18139), .ZN(n20160) );
  OAI21_X1 U20206 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20160), .A(
        n18130), .ZN(n20170) );
  OAI21_X1 U20207 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18132), .A(
        n18131), .ZN(n20868) );
  OAI22_X1 U20208 ( .A1(n18153), .A2(n20170), .B1(n18171), .B2(n20868), .ZN(
        n18133) );
  AOI21_X1 U20209 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18145), .A(
        n18133), .ZN(n18134) );
  OAI211_X1 U20210 ( .C1(n18170), .C2(n20869), .A(n18135), .B(n18134), .ZN(
        P3_U2826) );
  OAI21_X1 U20211 ( .B1(n18138), .B2(n18137), .A(n18136), .ZN(n20862) );
  NOR2_X1 U20212 ( .A1(n18156), .A2(n18155), .ZN(n18144) );
  NOR2_X1 U20213 ( .A1(n18155), .A2(n20130), .ZN(n20146) );
  OAI21_X1 U20214 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20146), .A(
        n18139), .ZN(n20148) );
  OAI21_X1 U20215 ( .B1(n18142), .B2(n18141), .A(n18140), .ZN(n20863) );
  OAI22_X1 U20216 ( .A1(n18153), .A2(n20148), .B1(n18170), .B2(n20863), .ZN(
        n18143) );
  AOI221_X1 U20217 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18145), .C1(
        n18144), .C2(n18145), .A(n18143), .ZN(n18146) );
  NAND2_X1 U20218 ( .A1(n10990), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n20866) );
  OAI211_X1 U20219 ( .C1(n18171), .C2(n20862), .A(n18146), .B(n20866), .ZN(
        P3_U2827) );
  OAI21_X1 U20220 ( .B1(n18149), .B2(n18148), .A(n18147), .ZN(n20851) );
  AOI21_X1 U20221 ( .B1(n18155), .B2(n20130), .A(n20146), .ZN(n20129) );
  INV_X1 U20222 ( .A(n20129), .ZN(n20134) );
  OAI21_X1 U20223 ( .B1(n18152), .B2(n18151), .A(n18150), .ZN(n20855) );
  OAI22_X1 U20224 ( .A1(n18153), .A2(n20134), .B1(n18171), .B2(n20855), .ZN(
        n18154) );
  AOI221_X1 U20225 ( .B1(n18156), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19011), .C2(n18155), .A(n18154), .ZN(n18157) );
  NAND2_X1 U20226 ( .A1(n10990), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n20853) );
  OAI211_X1 U20227 ( .C1(n18170), .C2(n20851), .A(n18157), .B(n20853), .ZN(
        P3_U2828) );
  OAI21_X1 U20228 ( .B1(n18159), .B2(n18165), .A(n18158), .ZN(n20845) );
  NAND2_X1 U20229 ( .A1(n20846), .A2(n20740), .ZN(n18160) );
  XNOR2_X1 U20230 ( .A(n18160), .B(n18159), .ZN(n20841) );
  AOI22_X1 U20231 ( .A1(n10990), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18161), 
        .B2(n20841), .ZN(n18164) );
  AOI22_X1 U20232 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18162), .B1(
        n18015), .B2(n20130), .ZN(n18163) );
  OAI211_X1 U20233 ( .C1(n18170), .C2(n20845), .A(n18164), .B(n18163), .ZN(
        P3_U2829) );
  AOI21_X1 U20234 ( .B1(n20740), .B2(n20846), .A(n18165), .ZN(n18172) );
  INV_X1 U20235 ( .A(n18172), .ZN(n20837) );
  NAND3_X1 U20236 ( .A1(n20750), .A2(n18167), .A3(n18166), .ZN(n18168) );
  AOI22_X1 U20237 ( .A1(n10990), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18168), .ZN(n18169) );
  OAI221_X1 U20238 ( .B1(n18172), .B2(n18171), .C1(n20837), .C2(n18170), .A(
        n18169), .ZN(P3_U2830) );
  NAND2_X1 U20239 ( .A1(n18674), .A2(n18683), .ZN(n18714) );
  INV_X1 U20240 ( .A(n18714), .ZN(n18707) );
  NOR2_X1 U20241 ( .A1(n21241), .A2(n18683), .ZN(n18689) );
  NAND2_X1 U20242 ( .A1(n21241), .A2(n18683), .ZN(n18741) );
  INV_X1 U20243 ( .A(n18741), .ZN(n18743) );
  INV_X1 U20244 ( .A(n18173), .ZN(n18736) );
  NOR3_X1 U20245 ( .A1(n18689), .A2(n18743), .A3(n18736), .ZN(n18174) );
  AOI21_X1 U20246 ( .B1(n18707), .B2(n18175), .A(n18174), .ZN(n18177) );
  OAI22_X1 U20247 ( .A1(n18178), .A2(n18177), .B1(n18176), .B2(n18683), .ZN(
        P3_U2866) );
  NOR4_X1 U20248 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18182) );
  NOR4_X1 U20249 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18181) );
  NOR4_X1 U20250 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18180) );
  NOR4_X1 U20251 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18179) );
  NAND4_X1 U20252 ( .A1(n18182), .A2(n18181), .A3(n18180), .A4(n18179), .ZN(
        n18188) );
  NOR4_X1 U20253 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18186) );
  AOI211_X1 U20254 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18185) );
  NOR4_X1 U20255 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18184) );
  NOR4_X1 U20256 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18183) );
  NAND4_X1 U20257 ( .A1(n18186), .A2(n18185), .A3(n18184), .A4(n18183), .ZN(
        n18187) );
  NOR2_X1 U20258 ( .A1(n18188), .A2(n18187), .ZN(n18196) );
  INV_X1 U20259 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18276) );
  OAI21_X1 U20260 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18196), .ZN(n18189) );
  OAI21_X1 U20261 ( .B1(n18196), .B2(n18276), .A(n18189), .ZN(P3_U3293) );
  INV_X1 U20262 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18280) );
  AOI21_X1 U20263 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18190) );
  INV_X1 U20264 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18239) );
  OAI221_X1 U20265 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18190), .C1(n18239), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18196), .ZN(n18191) );
  OAI21_X1 U20266 ( .B1(n18196), .B2(n18280), .A(n18191), .ZN(P3_U3292) );
  INV_X1 U20267 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18278) );
  NOR3_X1 U20268 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18193) );
  OAI21_X1 U20269 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18193), .A(n18196), .ZN(
        n18192) );
  OAI21_X1 U20270 ( .B1(n18196), .B2(n18278), .A(n18192), .ZN(P3_U2638) );
  INV_X1 U20271 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21705) );
  AOI21_X1 U20272 ( .B1(n18239), .B2(n21705), .A(n18193), .ZN(n18195) );
  INV_X1 U20273 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18282) );
  INV_X1 U20274 ( .A(n18196), .ZN(n18194) );
  AOI22_X1 U20275 ( .A1(n18196), .A2(n18195), .B1(n18282), .B2(n18194), .ZN(
        P3_U2639) );
  INV_X1 U20276 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18283) );
  AOI22_X1 U20277 ( .A1(n21713), .A2(n18197), .B1(n18283), .B2(n21765), .ZN(
        P3_U3297) );
  INV_X1 U20278 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18198) );
  AOI22_X1 U20279 ( .A1(n21713), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18198), 
        .B2(n21765), .ZN(P3_U3294) );
  AOI21_X1 U20280 ( .B1(n21767), .B2(n21709), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18199) );
  AOI22_X1 U20281 ( .A1(n21713), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18199), 
        .B2(n21765), .ZN(P3_U2635) );
  INV_X1 U20282 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20728) );
  AOI22_X1 U20283 ( .A1(n18233), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18200) );
  OAI21_X1 U20284 ( .B1(n20728), .B2(n18216), .A(n18200), .ZN(P3_U2767) );
  INV_X1 U20285 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20586) );
  AOI22_X1 U20286 ( .A1(n18233), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18201) );
  OAI21_X1 U20287 ( .B1(n20586), .B2(n18216), .A(n18201), .ZN(P3_U2766) );
  INV_X1 U20288 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U20289 ( .A1(n18233), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18202) );
  OAI21_X1 U20290 ( .B1(n20091), .B2(n18216), .A(n18202), .ZN(P3_U2765) );
  INV_X1 U20291 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20093) );
  AOI22_X1 U20292 ( .A1(n18233), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18203) );
  OAI21_X1 U20293 ( .B1(n20093), .B2(n18216), .A(n18203), .ZN(P3_U2764) );
  INV_X1 U20294 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20587) );
  AOI22_X1 U20295 ( .A1(n18233), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18204) );
  OAI21_X1 U20296 ( .B1(n20587), .B2(n18216), .A(n18204), .ZN(P3_U2763) );
  INV_X1 U20297 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20096) );
  AOI22_X1 U20298 ( .A1(n18233), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18205) );
  OAI21_X1 U20299 ( .B1(n20096), .B2(n18216), .A(n18205), .ZN(P3_U2762) );
  INV_X1 U20300 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U20301 ( .A1(n18233), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18206) );
  OAI21_X1 U20302 ( .B1(n20588), .B2(n18216), .A(n18206), .ZN(P3_U2761) );
  INV_X1 U20303 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20100) );
  AOI22_X1 U20304 ( .A1(n18233), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18207) );
  OAI21_X1 U20305 ( .B1(n20100), .B2(n18216), .A(n18207), .ZN(P3_U2760) );
  INV_X1 U20306 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20721) );
  AOI22_X1 U20307 ( .A1(n18233), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18208) );
  OAI21_X1 U20308 ( .B1(n20721), .B2(n18216), .A(n18208), .ZN(P3_U2759) );
  INV_X1 U20309 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20562) );
  AOI22_X1 U20310 ( .A1(n18233), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18209) );
  OAI21_X1 U20311 ( .B1(n20562), .B2(n18216), .A(n18209), .ZN(P3_U2758) );
  INV_X1 U20312 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U20313 ( .A1(n18233), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18210) );
  OAI21_X1 U20314 ( .B1(n20555), .B2(n18216), .A(n18210), .ZN(P3_U2757) );
  INV_X1 U20315 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20563) );
  AOI22_X1 U20316 ( .A1(n18233), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18211) );
  OAI21_X1 U20317 ( .B1(n20563), .B2(n18216), .A(n18211), .ZN(P3_U2756) );
  INV_X1 U20318 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20556) );
  AOI22_X1 U20319 ( .A1(n18233), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18212) );
  OAI21_X1 U20320 ( .B1(n20556), .B2(n18216), .A(n18212), .ZN(P3_U2755) );
  INV_X1 U20321 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U20322 ( .A1(n18233), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18213) );
  OAI21_X1 U20323 ( .B1(n20107), .B2(n18216), .A(n18213), .ZN(P3_U2754) );
  INV_X1 U20324 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U20325 ( .A1(n18233), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18214) );
  OAI21_X1 U20326 ( .B1(n20711), .B2(n18216), .A(n18214), .ZN(P3_U2753) );
  INV_X1 U20327 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20717) );
  AOI22_X1 U20328 ( .A1(n18233), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18215) );
  OAI21_X1 U20329 ( .B1(n20717), .B2(n18216), .A(n18215), .ZN(P3_U2752) );
  INV_X1 U20330 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U20331 ( .A1(n18233), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18218) );
  OAI21_X1 U20332 ( .B1(n20065), .B2(n18235), .A(n18218), .ZN(P3_U2751) );
  INV_X1 U20333 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20067) );
  AOI22_X1 U20334 ( .A1(n18233), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18219) );
  OAI21_X1 U20335 ( .B1(n20067), .B2(n18235), .A(n18219), .ZN(P3_U2750) );
  INV_X1 U20336 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20069) );
  AOI22_X1 U20337 ( .A1(n18233), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18220) );
  OAI21_X1 U20338 ( .B1(n20069), .B2(n18235), .A(n18220), .ZN(P3_U2749) );
  INV_X1 U20339 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20631) );
  AOI22_X1 U20340 ( .A1(n18233), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18221) );
  OAI21_X1 U20341 ( .B1(n20631), .B2(n18235), .A(n18221), .ZN(P3_U2748) );
  INV_X1 U20342 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20072) );
  AOI22_X1 U20343 ( .A1(n18233), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18222) );
  OAI21_X1 U20344 ( .B1(n20072), .B2(n18235), .A(n18222), .ZN(P3_U2747) );
  INV_X1 U20345 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20647) );
  AOI22_X1 U20346 ( .A1(n18233), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18223) );
  OAI21_X1 U20347 ( .B1(n20647), .B2(n18235), .A(n18223), .ZN(P3_U2746) );
  INV_X1 U20348 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20648) );
  AOI22_X1 U20349 ( .A1(n18233), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18224) );
  OAI21_X1 U20350 ( .B1(n20648), .B2(n18235), .A(n18224), .ZN(P3_U2745) );
  INV_X1 U20351 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20076) );
  AOI22_X1 U20352 ( .A1(n18233), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18225) );
  OAI21_X1 U20353 ( .B1(n20076), .B2(n18235), .A(n18225), .ZN(P3_U2744) );
  INV_X1 U20354 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20078) );
  AOI22_X1 U20355 ( .A1(n18233), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18227) );
  OAI21_X1 U20356 ( .B1(n20078), .B2(n18235), .A(n18227), .ZN(P3_U2743) );
  INV_X1 U20357 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U20358 ( .A1(n18233), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18228) );
  OAI21_X1 U20359 ( .B1(n20650), .B2(n18235), .A(n18228), .ZN(P3_U2742) );
  INV_X1 U20360 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20082) );
  AOI22_X1 U20361 ( .A1(n18233), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18229) );
  OAI21_X1 U20362 ( .B1(n20082), .B2(n18235), .A(n18229), .ZN(P3_U2741) );
  INV_X1 U20363 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20681) );
  AOI22_X1 U20364 ( .A1(n18233), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18230) );
  OAI21_X1 U20365 ( .B1(n20681), .B2(n18235), .A(n18230), .ZN(P3_U2740) );
  INV_X1 U20366 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20085) );
  AOI22_X1 U20367 ( .A1(n18233), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18231) );
  OAI21_X1 U20368 ( .B1(n20085), .B2(n18235), .A(n18231), .ZN(P3_U2739) );
  INV_X1 U20369 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U20370 ( .A1(n18233), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18232) );
  OAI21_X1 U20371 ( .B1(n20669), .B2(n18235), .A(n18232), .ZN(P3_U2738) );
  INV_X1 U20372 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20667) );
  AOI22_X1 U20373 ( .A1(n18233), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18226), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18234) );
  OAI21_X1 U20374 ( .B1(n20667), .B2(n18235), .A(n18234), .ZN(P3_U2737) );
  NOR2_X1 U20375 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18236), .ZN(n18237) );
  NOR2_X1 U20376 ( .A1(n21713), .A2(n18237), .ZN(P3_U2633) );
  INV_X1 U20377 ( .A(n18269), .ZN(n18274) );
  AOI22_X1 U20378 ( .A1(n18272), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n21765), .ZN(n18238) );
  OAI21_X1 U20379 ( .B1(n18274), .B2(n18239), .A(n18238), .ZN(P3_U3032) );
  INV_X1 U20380 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U20381 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n21765), .ZN(n18240) );
  OAI21_X1 U20382 ( .B1(n20150), .B2(n18271), .A(n18240), .ZN(P3_U3033) );
  AOI22_X1 U20383 ( .A1(n18272), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n21765), .ZN(n18241) );
  OAI21_X1 U20384 ( .B1(n18274), .B2(n20150), .A(n18241), .ZN(P3_U3034) );
  INV_X1 U20385 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20162) );
  AOI22_X1 U20386 ( .A1(n18272), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n21765), .ZN(n18242) );
  OAI21_X1 U20387 ( .B1(n18274), .B2(n20162), .A(n18242), .ZN(P3_U3035) );
  AOI22_X1 U20388 ( .A1(n18272), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n21765), .ZN(n18243) );
  OAI21_X1 U20389 ( .B1(n18274), .B2(n20179), .A(n18243), .ZN(P3_U3036) );
  AOI22_X1 U20390 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n21765), .ZN(n18244) );
  OAI21_X1 U20391 ( .B1(n20898), .B2(n18271), .A(n18244), .ZN(P3_U3037) );
  AOI22_X1 U20392 ( .A1(n18272), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n21765), .ZN(n18245) );
  OAI21_X1 U20393 ( .B1(n18274), .B2(n20898), .A(n18245), .ZN(P3_U3038) );
  AOI22_X1 U20394 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n21765), .ZN(n18246) );
  OAI21_X1 U20395 ( .B1(n20245), .B2(n18271), .A(n18246), .ZN(P3_U3039) );
  AOI22_X1 U20396 ( .A1(n18272), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n21765), .ZN(n18247) );
  OAI21_X1 U20397 ( .B1(n18274), .B2(n20245), .A(n18247), .ZN(P3_U3040) );
  AOI22_X1 U20398 ( .A1(n18272), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n21765), .ZN(n18248) );
  OAI21_X1 U20399 ( .B1(n18274), .B2(n20246), .A(n18248), .ZN(P3_U3041) );
  AOI22_X1 U20400 ( .A1(n18272), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n21765), .ZN(n18249) );
  OAI21_X1 U20401 ( .B1(n18274), .B2(n20278), .A(n18249), .ZN(P3_U3042) );
  INV_X1 U20402 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U20403 ( .A1(n18272), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n21765), .ZN(n18250) );
  OAI21_X1 U20404 ( .B1(n18274), .B2(n18251), .A(n18250), .ZN(P3_U3043) );
  INV_X1 U20405 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U20406 ( .A1(n18272), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n21765), .ZN(n18252) );
  OAI21_X1 U20407 ( .B1(n18274), .B2(n18253), .A(n18252), .ZN(P3_U3044) );
  AOI22_X1 U20408 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n21765), .ZN(n18254) );
  OAI21_X1 U20409 ( .B1(n20322), .B2(n18271), .A(n18254), .ZN(P3_U3045) );
  AOI22_X1 U20410 ( .A1(n18272), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n21765), .ZN(n18255) );
  OAI21_X1 U20411 ( .B1(n18274), .B2(n20322), .A(n18255), .ZN(P3_U3046) );
  AOI22_X1 U20412 ( .A1(n18272), .A2(P3_REIP_REG_17__SCAN_IN), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n21765), .ZN(n18256) );
  OAI21_X1 U20413 ( .B1(n18274), .B2(n21181), .A(n18256), .ZN(P3_U3047) );
  INV_X1 U20414 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20345) );
  AOI22_X1 U20415 ( .A1(n18272), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n21765), .ZN(n18257) );
  OAI21_X1 U20416 ( .B1(n18274), .B2(n20345), .A(n18257), .ZN(P3_U3048) );
  AOI22_X1 U20417 ( .A1(n18272), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n21765), .ZN(n18258) );
  OAI21_X1 U20418 ( .B1(n18274), .B2(n21166), .A(n18258), .ZN(P3_U3049) );
  INV_X1 U20419 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21150) );
  AOI22_X1 U20420 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n21765), .ZN(n18259) );
  OAI21_X1 U20421 ( .B1(n21150), .B2(n18271), .A(n18259), .ZN(P3_U3050) );
  AOI22_X1 U20422 ( .A1(n18272), .A2(P3_REIP_REG_21__SCAN_IN), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n21765), .ZN(n18260) );
  OAI21_X1 U20423 ( .B1(n18274), .B2(n21150), .A(n18260), .ZN(P3_U3051) );
  AOI22_X1 U20424 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n21765), .ZN(n18261) );
  OAI21_X1 U20425 ( .B1(n20420), .B2(n18271), .A(n18261), .ZN(P3_U3052) );
  AOI22_X1 U20426 ( .A1(n18272), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n21765), .ZN(n18262) );
  OAI21_X1 U20427 ( .B1(n18274), .B2(n20420), .A(n18262), .ZN(P3_U3053) );
  AOI22_X1 U20428 ( .A1(n18272), .A2(P3_REIP_REG_24__SCAN_IN), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n21765), .ZN(n18263) );
  OAI21_X1 U20429 ( .B1(n18274), .B2(n20425), .A(n18263), .ZN(P3_U3054) );
  INV_X1 U20430 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20466) );
  AOI22_X1 U20431 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n21765), .ZN(n18264) );
  OAI21_X1 U20432 ( .B1(n20466), .B2(n18271), .A(n18264), .ZN(P3_U3055) );
  AOI22_X1 U20433 ( .A1(n18272), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n21765), .ZN(n18265) );
  OAI21_X1 U20434 ( .B1(n18274), .B2(n20466), .A(n18265), .ZN(P3_U3056) );
  AOI22_X1 U20435 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n21765), .ZN(n18266) );
  OAI21_X1 U20436 ( .B1(n20487), .B2(n18271), .A(n18266), .ZN(P3_U3057) );
  AOI22_X1 U20437 ( .A1(n18272), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n21765), .ZN(n18267) );
  OAI21_X1 U20438 ( .B1(n18274), .B2(n20487), .A(n18267), .ZN(P3_U3058) );
  INV_X1 U20439 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20497) );
  AOI22_X1 U20440 ( .A1(n18272), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n21765), .ZN(n18268) );
  OAI21_X1 U20441 ( .B1(n18274), .B2(n20497), .A(n18268), .ZN(P3_U3059) );
  INV_X1 U20442 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20515) );
  AOI22_X1 U20443 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18269), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n21765), .ZN(n18270) );
  OAI21_X1 U20444 ( .B1(n20515), .B2(n18271), .A(n18270), .ZN(P3_U3060) );
  AOI22_X1 U20445 ( .A1(n18272), .A2(P3_REIP_REG_31__SCAN_IN), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n21765), .ZN(n18273) );
  OAI21_X1 U20446 ( .B1(n18274), .B2(n20515), .A(n18273), .ZN(P3_U3061) );
  INV_X1 U20447 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U20448 ( .A1(n21713), .A2(n18276), .B1(n18275), .B2(n21765), .ZN(
        P3_U3277) );
  INV_X1 U20449 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U20450 ( .A1(n21713), .A2(n18278), .B1(n18277), .B2(n21765), .ZN(
        P3_U3276) );
  INV_X1 U20451 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U20452 ( .A1(n21713), .A2(n18280), .B1(n18279), .B2(n21765), .ZN(
        P3_U3275) );
  INV_X1 U20453 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20454 ( .A1(n21713), .A2(n18282), .B1(n18281), .B2(n21765), .ZN(
        P3_U3274) );
  NOR4_X1 U20455 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18285)
         );
  NOR4_X1 U20456 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18283), .ZN(n18284) );
  NAND3_X1 U20457 ( .A1(n18285), .A2(n18284), .A3(U215), .ZN(U213) );
  NAND4_X1 U20458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n18286), .A4(n21735), .ZN(n18287) );
  OAI211_X1 U20459 ( .C1(n18634), .C2(n18289), .A(n18288), .B(n18287), .ZN(
        n18301) );
  INV_X1 U20460 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21745) );
  AOI211_X1 U20461 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n18292), .A(n18291), 
        .B(n18290), .ZN(n18299) );
  INV_X1 U20462 ( .A(n18293), .ZN(n18297) );
  NOR2_X1 U20463 ( .A1(n18630), .A2(n19335), .ZN(n18294) );
  OAI22_X1 U20464 ( .A1(n18297), .A2(n18296), .B1(n18295), .B2(n18294), .ZN(
        n18298) );
  OAI21_X1 U20465 ( .B1(n18299), .B2(n18298), .A(n18301), .ZN(n18300) );
  OAI21_X1 U20466 ( .B1(n18301), .B2(n21745), .A(n18300), .ZN(P2_U3610) );
  AOI22_X1 U20467 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18561), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18577), .ZN(n18316) );
  INV_X1 U20468 ( .A(n18302), .ZN(n18304) );
  OAI22_X1 U20469 ( .A1(n18562), .A2(n18304), .B1(n18522), .B2(n18303), .ZN(
        n18305) );
  AOI211_X1 U20470 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18576), .A(n16396), .B(
        n18305), .ZN(n18315) );
  OAI22_X1 U20471 ( .A1(n19399), .A2(n18307), .B1(n18578), .B2(n18306), .ZN(
        n18308) );
  INV_X1 U20472 ( .A(n18308), .ZN(n18314) );
  AND2_X1 U20473 ( .A1(n18584), .A2(n18309), .ZN(n18311) );
  AOI21_X1 U20474 ( .B1(n18312), .B2(n18311), .A(n18627), .ZN(n18310) );
  OAI21_X1 U20475 ( .B1(n18312), .B2(n18311), .A(n18310), .ZN(n18313) );
  NAND4_X1 U20476 ( .A1(n18316), .A2(n18315), .A3(n18314), .A4(n18313), .ZN(
        P2_U2851) );
  NOR2_X1 U20477 ( .A1(n18376), .A2(n18317), .ZN(n18318) );
  XOR2_X1 U20478 ( .A(n18319), .B(n18318), .Z(n18327) );
  INV_X1 U20479 ( .A(n18320), .ZN(n18321) );
  AOI22_X1 U20480 ( .A1(n13297), .A2(n18321), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18577), .ZN(n18322) );
  OAI211_X1 U20481 ( .C1(n15177), .C2(n18520), .A(n18322), .B(n18381), .ZN(
        n18325) );
  OAI22_X1 U20482 ( .A1(n19403), .A2(n18562), .B1(n18578), .B2(n18323), .ZN(
        n18324) );
  AOI211_X1 U20483 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n18561), .A(n18325), .B(
        n18324), .ZN(n18326) );
  OAI21_X1 U20484 ( .B1(n18627), .B2(n18327), .A(n18326), .ZN(P2_U2850) );
  NAND2_X1 U20485 ( .A1(n18584), .A2(n18328), .ZN(n18330) );
  XOR2_X1 U20486 ( .A(n18330), .B(n18329), .Z(n18341) );
  INV_X1 U20487 ( .A(n18331), .ZN(n18332) );
  AOI22_X1 U20488 ( .A1(n18561), .A2(P2_EBX_REG_6__SCAN_IN), .B1(n13297), .B2(
        n18332), .ZN(n18333) );
  OAI211_X1 U20489 ( .C1(n18334), .C2(n18520), .A(n18333), .B(n18381), .ZN(
        n18339) );
  INV_X1 U20490 ( .A(n18335), .ZN(n18336) );
  OAI22_X1 U20491 ( .A1(n18337), .A2(n18562), .B1(n18578), .B2(n18336), .ZN(
        n18338) );
  AOI211_X1 U20492 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18577), .A(
        n18339), .B(n18338), .ZN(n18340) );
  OAI21_X1 U20493 ( .B1(n18341), .B2(n18627), .A(n18340), .ZN(P2_U2849) );
  NOR2_X1 U20494 ( .A1(n18376), .A2(n18342), .ZN(n18343) );
  XOR2_X1 U20495 ( .A(n18344), .B(n18343), .Z(n18353) );
  AOI22_X1 U20496 ( .A1(n18561), .A2(P2_EBX_REG_7__SCAN_IN), .B1(n13297), .B2(
        n18345), .ZN(n18346) );
  OAI211_X1 U20497 ( .C1(n18347), .C2(n18520), .A(n18346), .B(n18381), .ZN(
        n18351) );
  OAI22_X1 U20498 ( .A1(n18349), .A2(n18562), .B1(n18578), .B2(n18348), .ZN(
        n18350) );
  AOI211_X1 U20499 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18577), .A(
        n18351), .B(n18350), .ZN(n18352) );
  OAI21_X1 U20500 ( .B1(n18627), .B2(n18353), .A(n18352), .ZN(P2_U2848) );
  OAI21_X1 U20501 ( .B1(n13042), .B2(n18520), .A(n18381), .ZN(n18357) );
  OAI22_X1 U20502 ( .A1(n18355), .A2(n18522), .B1(n18537), .B2(n18354), .ZN(
        n18356) );
  AOI211_X1 U20503 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18577), .A(
        n18357), .B(n18356), .ZN(n18365) );
  NOR2_X1 U20504 ( .A1(n18376), .A2(n18358), .ZN(n18360) );
  XNOR2_X1 U20505 ( .A(n18360), .B(n18359), .ZN(n18363) );
  AOI22_X1 U20506 ( .A1(n18363), .A2(n18362), .B1(n18551), .B2(n18361), .ZN(
        n18364) );
  OAI211_X1 U20507 ( .C1(n18562), .C2(n18366), .A(n18365), .B(n18364), .ZN(
        P2_U2846) );
  NAND2_X1 U20508 ( .A1(n18551), .A2(n18367), .ZN(n18369) );
  AOI22_X1 U20509 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18577), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n18561), .ZN(n18368) );
  NAND3_X1 U20510 ( .A1(n18369), .A2(n18368), .A3(n18381), .ZN(n18372) );
  OAI22_X1 U20511 ( .A1(n18562), .A2(n18370), .B1(n18520), .B2(n16663), .ZN(
        n18371) );
  NOR2_X1 U20512 ( .A1(n18372), .A2(n18371), .ZN(n18373) );
  OAI21_X1 U20513 ( .B1(n18374), .B2(n18522), .A(n18373), .ZN(n18375) );
  INV_X1 U20514 ( .A(n18375), .ZN(n18379) );
  NOR2_X1 U20515 ( .A1(n18376), .A2(n18627), .ZN(n18424) );
  OAI211_X1 U20516 ( .C1(n18377), .C2(n18380), .A(n18424), .B(n18386), .ZN(
        n18378) );
  OAI211_X1 U20517 ( .C1(n18407), .C2(n18380), .A(n18379), .B(n18378), .ZN(
        P2_U2844) );
  OAI21_X1 U20518 ( .B1(n13048), .B2(n18520), .A(n18381), .ZN(n18385) );
  OAI22_X1 U20519 ( .A1(n18383), .A2(n18522), .B1(n18488), .B2(n18382), .ZN(
        n18384) );
  AOI211_X1 U20520 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n18561), .A(n18385), .B(
        n18384), .ZN(n18392) );
  NAND2_X1 U20521 ( .A1(n18584), .A2(n18386), .ZN(n18387) );
  XNOR2_X1 U20522 ( .A(n18388), .B(n18387), .ZN(n18390) );
  AOI22_X1 U20523 ( .A1(n18390), .A2(n18362), .B1(n18551), .B2(n18389), .ZN(
        n18391) );
  OAI211_X1 U20524 ( .C1(n18562), .C2(n19124), .A(n18392), .B(n18391), .ZN(
        P2_U2843) );
  OAI21_X1 U20525 ( .B1(n18488), .B2(n16423), .A(n14035), .ZN(n18393) );
  AOI21_X1 U20526 ( .B1(n18576), .B2(P2_REIP_REG_13__SCAN_IN), .A(n18393), 
        .ZN(n18394) );
  OAI21_X1 U20527 ( .B1(n18537), .B2(n18395), .A(n18394), .ZN(n18400) );
  AND2_X1 U20528 ( .A1(n18584), .A2(n18396), .ZN(n18409) );
  OAI211_X1 U20529 ( .C1(n18397), .C2(n18408), .A(n18362), .B(n18409), .ZN(
        n18398) );
  INV_X1 U20530 ( .A(n18398), .ZN(n18399) );
  AOI211_X1 U20531 ( .C1(n13297), .C2(n18401), .A(n18400), .B(n18399), .ZN(
        n18406) );
  INV_X1 U20532 ( .A(n18402), .ZN(n18404) );
  AOI22_X1 U20533 ( .A1(n18580), .A2(n18404), .B1(n18551), .B2(n18403), .ZN(
        n18405) );
  OAI211_X1 U20534 ( .C1(n18408), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P2_U2842) );
  XNOR2_X1 U20535 ( .A(n18410), .B(n18409), .ZN(n18420) );
  AOI22_X1 U20536 ( .A1(n18411), .A2(n13297), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n18561), .ZN(n18412) );
  OAI21_X1 U20537 ( .B1(n18413), .B2(n18488), .A(n18412), .ZN(n18414) );
  AOI211_X1 U20538 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18576), .A(n16396), 
        .B(n18414), .ZN(n18419) );
  AOI21_X1 U20539 ( .B1(n18416), .B2(n18415), .A(n14934), .ZN(n19118) );
  INV_X1 U20540 ( .A(n18417), .ZN(n18599) );
  AOI22_X1 U20541 ( .A1(n18580), .A2(n19118), .B1(n18551), .B2(n18599), .ZN(
        n18418) );
  OAI211_X1 U20542 ( .C1(n18627), .C2(n18420), .A(n18419), .B(n18418), .ZN(
        P2_U2841) );
  OAI21_X1 U20543 ( .B1(n18488), .B2(n13190), .A(n14035), .ZN(n18421) );
  AOI21_X1 U20544 ( .B1(n18576), .B2(P2_REIP_REG_15__SCAN_IN), .A(n18421), 
        .ZN(n18422) );
  OAI21_X1 U20545 ( .B1(n18537), .B2(n13283), .A(n18422), .ZN(n18428) );
  OAI211_X1 U20546 ( .C1(n18425), .C2(n18430), .A(n18424), .B(n18423), .ZN(
        n18426) );
  INV_X1 U20547 ( .A(n18426), .ZN(n18427) );
  AOI211_X1 U20548 ( .C1(n13297), .C2(n18429), .A(n18428), .B(n18427), .ZN(
        n18435) );
  INV_X1 U20549 ( .A(n18430), .ZN(n18432) );
  AOI22_X1 U20550 ( .A1(n18433), .A2(n18551), .B1(n18432), .B2(n18431), .ZN(
        n18434) );
  OAI211_X1 U20551 ( .C1(n18562), .C2(n18436), .A(n18435), .B(n18434), .ZN(
        P2_U2840) );
  AOI22_X1 U20552 ( .A1(n18437), .A2(n13297), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18577), .ZN(n18438) );
  OAI211_X1 U20553 ( .C1(n18439), .C2(n18520), .A(n18438), .B(n18381), .ZN(
        n18444) );
  INV_X1 U20554 ( .A(n18440), .ZN(n18441) );
  OAI22_X1 U20555 ( .A1(n18442), .A2(n18578), .B1(n18441), .B2(n18562), .ZN(
        n18443) );
  AOI211_X1 U20556 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18561), .A(n18444), .B(
        n18443), .ZN(n18449) );
  OAI211_X1 U20557 ( .C1(n18447), .C2(n18446), .A(n18362), .B(n18445), .ZN(
        n18448) );
  NAND2_X1 U20558 ( .A1(n18449), .A2(n18448), .ZN(P2_U2838) );
  AOI22_X1 U20559 ( .A1(n18450), .A2(n13297), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18561), .ZN(n18451) );
  OAI211_X1 U20560 ( .C1(n18452), .C2(n18520), .A(n18451), .B(n14035), .ZN(
        n18456) );
  OAI22_X1 U20561 ( .A1(n18454), .A2(n18578), .B1(n18562), .B2(n18453), .ZN(
        n18455) );
  AOI211_X1 U20562 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18577), .A(
        n18456), .B(n18455), .ZN(n18461) );
  OAI211_X1 U20563 ( .C1(n18459), .C2(n18458), .A(n18362), .B(n18457), .ZN(
        n18460) );
  NAND2_X1 U20564 ( .A1(n18461), .A2(n18460), .ZN(P2_U2837) );
  AOI22_X1 U20565 ( .A1(n18561), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18577), .ZN(n18462) );
  OAI21_X1 U20566 ( .B1(n18463), .B2(n18522), .A(n18462), .ZN(n18464) );
  AOI211_X1 U20567 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n18576), .A(n16396), 
        .B(n18464), .ZN(n18473) );
  OAI22_X1 U20568 ( .A1(n18466), .A2(n18578), .B1(n18465), .B2(n18562), .ZN(
        n18467) );
  INV_X1 U20569 ( .A(n18467), .ZN(n18472) );
  OAI211_X1 U20570 ( .C1(n18470), .C2(n18469), .A(n18362), .B(n18468), .ZN(
        n18471) );
  NAND3_X1 U20571 ( .A1(n18473), .A2(n18472), .A3(n18471), .ZN(P2_U2836) );
  OAI22_X1 U20572 ( .A1(n13215), .A2(n18488), .B1(n18474), .B2(n18520), .ZN(
        n18476) );
  NOR2_X1 U20573 ( .A1(n18537), .A2(n13819), .ZN(n18475) );
  NOR2_X1 U20574 ( .A1(n18476), .A2(n18475), .ZN(n18477) );
  OAI21_X1 U20575 ( .B1(n18478), .B2(n18578), .A(n18477), .ZN(n18479) );
  AOI21_X1 U20576 ( .B1(n18480), .B2(n13297), .A(n18479), .ZN(n18485) );
  OAI211_X1 U20577 ( .C1(n18483), .C2(n18482), .A(n18362), .B(n18481), .ZN(
        n18484) );
  OAI211_X1 U20578 ( .C1(n18562), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P2_U2834) );
  INV_X1 U20579 ( .A(n18487), .ZN(n18493) );
  OAI22_X1 U20580 ( .A1(n18578), .A2(n18489), .B1(n18488), .B2(n13144), .ZN(
        n18490) );
  AOI21_X1 U20581 ( .B1(n18576), .B2(P2_REIP_REG_23__SCAN_IN), .A(n18490), 
        .ZN(n18491) );
  OAI21_X1 U20582 ( .B1(n18537), .B2(n13287), .A(n18491), .ZN(n18492) );
  AOI21_X1 U20583 ( .B1(n18493), .B2(n13297), .A(n18492), .ZN(n18498) );
  OAI211_X1 U20584 ( .C1(n18496), .C2(n18495), .A(n18362), .B(n18494), .ZN(
        n18497) );
  OAI211_X1 U20585 ( .C1(n18499), .C2(n18562), .A(n18498), .B(n18497), .ZN(
        P2_U2832) );
  AOI22_X1 U20586 ( .A1(n18500), .A2(n13297), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n18576), .ZN(n18509) );
  AOI22_X1 U20587 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18561), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18577), .ZN(n18508) );
  AOI22_X1 U20588 ( .A1(n18502), .A2(n18551), .B1(n18580), .B2(n18501), .ZN(
        n18507) );
  OAI211_X1 U20589 ( .C1(n18505), .C2(n18504), .A(n18362), .B(n18503), .ZN(
        n18506) );
  NAND4_X1 U20590 ( .A1(n18509), .A2(n18508), .A3(n18507), .A4(n18506), .ZN(
        P2_U2831) );
  AOI22_X1 U20591 ( .A1(n18510), .A2(n13297), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n18576), .ZN(n18519) );
  AOI22_X1 U20592 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18577), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18561), .ZN(n18518) );
  AOI22_X1 U20593 ( .A1(n18512), .A2(n18551), .B1(n18580), .B2(n18511), .ZN(
        n18517) );
  OAI211_X1 U20594 ( .C1(n18515), .C2(n18514), .A(n18362), .B(n18513), .ZN(
        n18516) );
  NAND4_X1 U20595 ( .A1(n18519), .A2(n18518), .A3(n18517), .A4(n18516), .ZN(
        P2_U2830) );
  OAI22_X1 U20596 ( .A1(n18523), .A2(n18522), .B1(n18521), .B2(n18520), .ZN(
        n18524) );
  INV_X1 U20597 ( .A(n18524), .ZN(n18534) );
  AOI22_X1 U20598 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18561), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18577), .ZN(n18533) );
  OAI22_X1 U20599 ( .A1(n18526), .A2(n18578), .B1(n18562), .B2(n18525), .ZN(
        n18527) );
  INV_X1 U20600 ( .A(n18527), .ZN(n18532) );
  OAI211_X1 U20601 ( .C1(n18530), .C2(n18529), .A(n18362), .B(n18528), .ZN(
        n18531) );
  NAND4_X1 U20602 ( .A1(n18534), .A2(n18533), .A3(n18532), .A4(n18531), .ZN(
        P2_U2829) );
  NOR2_X1 U20603 ( .A1(n18535), .A2(n18578), .ZN(n18539) );
  AOI22_X1 U20604 ( .A1(n18576), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18577), .ZN(n18536) );
  OAI21_X1 U20605 ( .B1(n18537), .B2(n13290), .A(n18536), .ZN(n18538) );
  AOI211_X1 U20606 ( .C1(n18540), .C2(n13297), .A(n18539), .B(n18538), .ZN(
        n18545) );
  OAI211_X1 U20607 ( .C1(n18543), .C2(n18542), .A(n18362), .B(n18541), .ZN(
        n18544) );
  OAI211_X1 U20608 ( .C1(n18562), .C2(n18546), .A(n18545), .B(n18544), .ZN(
        P2_U2828) );
  INV_X1 U20609 ( .A(n18547), .ZN(n18548) );
  AOI22_X1 U20610 ( .A1(n18548), .A2(n13297), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n18576), .ZN(n18559) );
  AOI22_X1 U20611 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18577), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18561), .ZN(n18558) );
  INV_X1 U20612 ( .A(n18549), .ZN(n18550) );
  AOI22_X1 U20613 ( .A1(n18552), .A2(n18551), .B1(n18550), .B2(n18580), .ZN(
        n18557) );
  OAI211_X1 U20614 ( .C1(n18555), .C2(n18554), .A(n18362), .B(n18553), .ZN(
        n18556) );
  NAND4_X1 U20615 ( .A1(n18559), .A2(n18558), .A3(n18557), .A4(n18556), .ZN(
        P2_U2827) );
  AOI22_X1 U20616 ( .A1(n18560), .A2(n13297), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n18576), .ZN(n18572) );
  AOI22_X1 U20617 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18561), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18577), .ZN(n18571) );
  OAI22_X1 U20618 ( .A1(n18564), .A2(n18578), .B1(n18563), .B2(n18562), .ZN(
        n18565) );
  INV_X1 U20619 ( .A(n18565), .ZN(n18570) );
  OAI211_X1 U20620 ( .C1(n18568), .C2(n18567), .A(n18362), .B(n18566), .ZN(
        n18569) );
  NAND4_X1 U20621 ( .A1(n18572), .A2(n18571), .A3(n18570), .A4(n18569), .ZN(
        P2_U2826) );
  NOR2_X1 U20622 ( .A1(n18573), .A2(n16091), .ZN(n18574) );
  AOI21_X1 U20623 ( .B1(n18575), .B2(n13297), .A(n18574), .ZN(n18589) );
  AOI22_X1 U20624 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18577), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18576), .ZN(n18588) );
  OR2_X1 U20625 ( .A1(n18579), .A2(n18578), .ZN(n18582) );
  NAND2_X1 U20626 ( .A1(n19115), .A2(n18580), .ZN(n18581) );
  AND2_X1 U20627 ( .A1(n18582), .A2(n18581), .ZN(n18587) );
  NAND4_X1 U20628 ( .A1(n18362), .A2(n18585), .A3(n18584), .A4(n18583), .ZN(
        n18586) );
  NAND4_X1 U20629 ( .A1(n18589), .A2(n18588), .A3(n18587), .A4(n18586), .ZN(
        P2_U2824) );
  NOR4_X1 U20630 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18592), .A3(
        n18591), .A4(n18590), .ZN(n18598) );
  NAND2_X1 U20631 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n16396), .ZN(n18593) );
  OAI221_X1 U20632 ( .B1(n18596), .B2(n18595), .C1(n18596), .C2(n18594), .A(
        n18593), .ZN(n18597) );
  AOI211_X1 U20633 ( .C1(n18606), .C2(n19118), .A(n18598), .B(n18597), .ZN(
        n18602) );
  AOI22_X1 U20634 ( .A1(n18600), .A2(n18609), .B1(n18611), .B2(n18599), .ZN(
        n18601) );
  OAI211_X1 U20635 ( .C1(n18604), .C2(n18603), .A(n18602), .B(n18601), .ZN(
        P2_U3032) );
  AOI22_X1 U20636 ( .A1(n18607), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18606), .B2(n18605), .ZN(n18619) );
  AOI222_X1 U20637 ( .A1(n18613), .A2(n18612), .B1(n18611), .B2(n18610), .C1(
        n18609), .C2(n18608), .ZN(n18618) );
  NAND2_X1 U20638 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16396), .ZN(n18617) );
  OAI211_X1 U20639 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n18615), .B(n18614), .ZN(n18616) );
  NAND4_X1 U20640 ( .A1(n18619), .A2(n18618), .A3(n18617), .A4(n18616), .ZN(
        P2_U3038) );
  NAND2_X1 U20641 ( .A1(n18633), .A2(n18620), .ZN(n18639) );
  OAI21_X1 U20642 ( .B1(n18622), .B2(n18621), .A(n18644), .ZN(n18626) );
  INV_X1 U20643 ( .A(n18629), .ZN(n18624) );
  NAND2_X1 U20644 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18630), .ZN(n18623) );
  AOI21_X1 U20645 ( .B1(n18624), .B2(n18639), .A(n18623), .ZN(n18625) );
  AOI21_X1 U20646 ( .B1(n18639), .B2(n18626), .A(n18625), .ZN(n18628) );
  NAND2_X1 U20647 ( .A1(n18628), .A2(n18627), .ZN(P2_U3177) );
  AOI22_X1 U20648 ( .A1(n18632), .A2(n18631), .B1(n18630), .B2(n18629), .ZN(
        n18643) );
  AOI22_X1 U20649 ( .A1(n18635), .A2(n18634), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n18633), .ZN(n18642) );
  OAI21_X1 U20650 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n18637), .A(n18636), 
        .ZN(n18638) );
  OAI21_X1 U20651 ( .B1(n18639), .B2(n21735), .A(n18638), .ZN(n18640) );
  NAND4_X1 U20652 ( .A1(n18643), .A2(n18642), .A3(n18641), .A4(n18640), .ZN(
        P2_U3176) );
  NOR2_X1 U20653 ( .A1(n18645), .A2(n18644), .ZN(n18648) );
  MUX2_X1 U20654 ( .A(P2_MORE_REG_SCAN_IN), .B(n18646), .S(n18648), .Z(
        P2_U3609) );
  OAI21_X1 U20655 ( .B1(n18648), .B2(n13888), .A(n18647), .ZN(P2_U2819) );
  INV_X1 U20656 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20051) );
  INV_X1 U20657 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18649) );
  AOI22_X1 U20658 ( .A1(n18964), .A2(n20051), .B1(n18649), .B2(U215), .ZN(U282) );
  OAI22_X1 U20659 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18964), .ZN(n18650) );
  INV_X1 U20660 ( .A(n18650), .ZN(U281) );
  OAI22_X1 U20661 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18964), .ZN(n18651) );
  INV_X1 U20662 ( .A(n18651), .ZN(U280) );
  OAI22_X1 U20663 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19010), .ZN(n18652) );
  INV_X1 U20664 ( .A(n18652), .ZN(U279) );
  OAI22_X1 U20665 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19010), .ZN(n18653) );
  INV_X1 U20666 ( .A(n18653), .ZN(U278) );
  OAI22_X1 U20667 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18964), .ZN(n18654) );
  INV_X1 U20668 ( .A(n18654), .ZN(U277) );
  OAI22_X1 U20669 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19010), .ZN(n18655) );
  INV_X1 U20670 ( .A(n18655), .ZN(U276) );
  OAI22_X1 U20671 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19010), .ZN(n18656) );
  INV_X1 U20672 ( .A(n18656), .ZN(U275) );
  OAI22_X1 U20673 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19010), .ZN(n18657) );
  INV_X1 U20674 ( .A(n18657), .ZN(U274) );
  OAI22_X1 U20675 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19010), .ZN(n18658) );
  INV_X1 U20676 ( .A(n18658), .ZN(U273) );
  OAI22_X1 U20677 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18964), .ZN(n18659) );
  INV_X1 U20678 ( .A(n18659), .ZN(U272) );
  OAI22_X1 U20679 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18964), .ZN(n18660) );
  INV_X1 U20680 ( .A(n18660), .ZN(U271) );
  OAI22_X1 U20681 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18964), .ZN(n18661) );
  INV_X1 U20682 ( .A(n18661), .ZN(U270) );
  OAI22_X1 U20683 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18964), .ZN(n18662) );
  INV_X1 U20684 ( .A(n18662), .ZN(U269) );
  OAI22_X1 U20685 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18964), .ZN(n18663) );
  INV_X1 U20686 ( .A(n18663), .ZN(U268) );
  OAI22_X1 U20687 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18964), .ZN(n18664) );
  INV_X1 U20688 ( .A(n18664), .ZN(U267) );
  OAI22_X1 U20689 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18964), .ZN(n18665) );
  INV_X1 U20690 ( .A(n18665), .ZN(U266) );
  OAI22_X1 U20691 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18964), .ZN(n18666) );
  INV_X1 U20692 ( .A(n18666), .ZN(U265) );
  INV_X1 U20693 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n18667) );
  INV_X1 U20694 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20561) );
  AOI22_X1 U20695 ( .A1(n18964), .A2(n18667), .B1(n20561), .B2(U215), .ZN(U264) );
  INV_X1 U20696 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18668) );
  INV_X1 U20697 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U20698 ( .A1(n18964), .A2(n18668), .B1(n20567), .B2(U215), .ZN(U263) );
  INV_X1 U20699 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n18669) );
  INV_X1 U20700 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20572) );
  AOI22_X1 U20701 ( .A1(n18964), .A2(n18669), .B1(n20572), .B2(U215), .ZN(U262) );
  INV_X1 U20702 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n18670) );
  INV_X1 U20703 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U20704 ( .A1(n19010), .A2(n18670), .B1(n20577), .B2(U215), .ZN(U261) );
  INV_X1 U20705 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18671) );
  INV_X1 U20706 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U20707 ( .A1(n19010), .A2(n18671), .B1(n20583), .B2(U215), .ZN(U260) );
  OAI22_X1 U20708 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18964), .ZN(n18672) );
  INV_X1 U20709 ( .A(n18672), .ZN(U259) );
  INV_X1 U20710 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18673) );
  INV_X1 U20711 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U20712 ( .A1(n18964), .A2(n18673), .B1(n20697), .B2(U215), .ZN(U258) );
  NAND2_X1 U20713 ( .A1(n21234), .A2(n18689), .ZN(n18687) );
  INV_X1 U20714 ( .A(n18687), .ZN(n18677) );
  NAND2_X1 U20715 ( .A1(n18677), .A2(n18721), .ZN(n18969) );
  NAND2_X1 U20716 ( .A1(n19011), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18735) );
  NAND2_X1 U20717 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19011), .ZN(n18748) );
  NOR2_X2 U20718 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21264), .ZN(n21273) );
  NAND2_X1 U20719 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18674), .ZN(
        n18675) );
  NOR2_X1 U20720 ( .A1(n21273), .A2(n18675), .ZN(n19014) );
  INV_X1 U20721 ( .A(n18966), .ZN(n19013) );
  NOR2_X2 U20722 ( .A1(n20697), .A2(n19013), .ZN(n18754) );
  AOI22_X1 U20723 ( .A1(n10969), .A2(n18755), .B1(n19014), .B2(n18754), .ZN(
        n18682) );
  INV_X1 U20724 ( .A(n18675), .ZN(n18745) );
  NOR2_X1 U20725 ( .A1(n18676), .A2(n19013), .ZN(n18688) );
  AOI22_X1 U20726 ( .A1(n19011), .A2(n18677), .B1(n18745), .B2(n18688), .ZN(
        n19017) );
  NAND2_X1 U20727 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21233) );
  INV_X1 U20728 ( .A(n21233), .ZN(n18700) );
  NAND2_X1 U20729 ( .A1(n18700), .A2(n18689), .ZN(n19094) );
  INV_X1 U20730 ( .A(n19094), .ZN(n19097) );
  INV_X1 U20731 ( .A(n18678), .ZN(n18679) );
  NAND2_X1 U20732 ( .A1(n18680), .A2(n18679), .ZN(n19015) );
  NOR2_X2 U20733 ( .A1(n20585), .A2(n19015), .ZN(n18756) );
  AOI22_X1 U20734 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18756), .ZN(n18681) );
  OAI211_X1 U20735 ( .C1(n18969), .C2(n18735), .A(n18682), .B(n18681), .ZN(
        P3_U2995) );
  NOR2_X1 U20736 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18683), .ZN(
        n18706) );
  NAND2_X1 U20737 ( .A1(n18700), .A2(n18706), .ZN(n19030) );
  INV_X1 U20738 ( .A(n18969), .ZN(n19032) );
  INV_X1 U20739 ( .A(n10969), .ZN(n19020) );
  NAND2_X1 U20740 ( .A1(n18745), .A2(n18721), .ZN(n19114) );
  AOI21_X1 U20741 ( .B1(n19020), .B2(n19114), .A(n21273), .ZN(n19021) );
  AOI22_X1 U20742 ( .A1(n19032), .A2(n18755), .B1(n18754), .B2(n19021), .ZN(
        n18686) );
  INV_X1 U20743 ( .A(n19114), .ZN(n19022) );
  INV_X1 U20744 ( .A(n19030), .ZN(n19038) );
  NOR2_X1 U20745 ( .A1(n19032), .A2(n19038), .ZN(n18692) );
  OAI22_X1 U20746 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19020), .B1(n18692), 
        .B2(n18736), .ZN(n18684) );
  OAI21_X1 U20747 ( .B1(n19022), .B2(n18684), .A(n18966), .ZN(n19023) );
  AOI22_X1 U20748 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19023), .B1(
        n18756), .B2(n19022), .ZN(n18685) );
  OAI211_X1 U20749 ( .C1(n18735), .C2(n19030), .A(n18686), .B(n18685), .ZN(
        P3_U2987) );
  NAND3_X1 U20750 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18706), .A3(
        n18721), .ZN(n19036) );
  NOR2_X1 U20751 ( .A1(n21273), .A2(n18687), .ZN(n19026) );
  AOI22_X1 U20752 ( .A1(n18755), .A2(n19038), .B1(n18754), .B2(n19026), .ZN(
        n18691) );
  INV_X1 U20753 ( .A(n18706), .ZN(n18705) );
  NOR2_X1 U20754 ( .A1(n21234), .A2(n18705), .ZN(n18696) );
  INV_X1 U20755 ( .A(n18688), .ZN(n18697) );
  NOR2_X1 U20756 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18697), .ZN(
        n18744) );
  AOI22_X1 U20757 ( .A1(n19011), .A2(n18696), .B1(n18689), .B2(n18744), .ZN(
        n19027) );
  AOI22_X1 U20758 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19027), .B1(
        n18756), .B2(n10969), .ZN(n18690) );
  OAI211_X1 U20759 ( .C1(n18735), .C2(n19036), .A(n18691), .B(n18690), .ZN(
        P3_U2979) );
  NOR2_X1 U20760 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18721), .ZN(
        n18726) );
  NAND2_X1 U20761 ( .A1(n18706), .A2(n18726), .ZN(n19042) );
  NOR2_X1 U20762 ( .A1(n21273), .A2(n18692), .ZN(n19031) );
  AOI22_X1 U20763 ( .A1(n18755), .A2(n19044), .B1(n18754), .B2(n19031), .ZN(
        n18695) );
  NOR2_X1 U20764 ( .A1(n19044), .A2(n19050), .ZN(n18702) );
  OAI22_X1 U20765 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19030), .B1(n18702), 
        .B2(n18736), .ZN(n18693) );
  OAI21_X1 U20766 ( .B1(n19032), .B2(n18693), .A(n18966), .ZN(n19033) );
  AOI22_X1 U20767 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18756), .ZN(n18694) );
  OAI211_X1 U20768 ( .C1(n18735), .C2(n19042), .A(n18695), .B(n18694), .ZN(
        P3_U2971) );
  INV_X1 U20769 ( .A(n18735), .ZN(n18757) );
  NOR2_X1 U20770 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21243) );
  NAND2_X1 U20771 ( .A1(n21243), .A2(n18706), .ZN(n18980) );
  INV_X1 U20772 ( .A(n21273), .ZN(n21259) );
  AND2_X1 U20773 ( .A1(n21259), .A2(n18696), .ZN(n19037) );
  AOI22_X1 U20774 ( .A1(n18757), .A2(n19056), .B1(n18754), .B2(n19037), .ZN(
        n18699) );
  AOI21_X1 U20775 ( .B1(n21234), .B2(n18736), .A(n18697), .ZN(n18732) );
  NAND2_X1 U20776 ( .A1(n18706), .A2(n18732), .ZN(n19039) );
  AOI22_X1 U20777 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19039), .B1(
        n18756), .B2(n19038), .ZN(n18698) );
  OAI211_X1 U20778 ( .C1(n18748), .C2(n19042), .A(n18699), .B(n18698), .ZN(
        P3_U2963) );
  NOR2_X1 U20779 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21241), .ZN(
        n18723) );
  NAND2_X1 U20780 ( .A1(n18700), .A2(n18723), .ZN(n19048) );
  NOR2_X1 U20781 ( .A1(n19056), .A2(n19062), .ZN(n18710) );
  OAI21_X1 U20782 ( .B1(n18710), .B2(n18736), .A(n18702), .ZN(n18701) );
  OAI211_X1 U20783 ( .C1(n19044), .C2(n21264), .A(n18966), .B(n18701), .ZN(
        n19045) );
  NOR2_X1 U20784 ( .A1(n21273), .A2(n18702), .ZN(n19043) );
  AOI22_X1 U20785 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19045), .B1(
        n18754), .B2(n19043), .ZN(n18704) );
  AOI22_X1 U20786 ( .A1(n18756), .A2(n19044), .B1(n18755), .B2(n19056), .ZN(
        n18703) );
  OAI211_X1 U20787 ( .C1(n18735), .C2(n19048), .A(n18704), .B(n18703), .ZN(
        P3_U2955) );
  NOR2_X2 U20788 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18714), .ZN(
        n19069) );
  NAND2_X1 U20789 ( .A1(n21234), .A2(n21259), .ZN(n18742) );
  NOR2_X1 U20790 ( .A1(n18705), .A2(n18742), .ZN(n19049) );
  AOI22_X1 U20791 ( .A1(n18757), .A2(n19069), .B1(n18754), .B2(n19049), .ZN(
        n18709) );
  AOI22_X1 U20792 ( .A1(n19011), .A2(n18707), .B1(n18706), .B2(n18744), .ZN(
        n19051) );
  AOI22_X1 U20793 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19051), .B1(
        n18756), .B2(n19050), .ZN(n18708) );
  OAI211_X1 U20794 ( .C1(n18748), .C2(n19048), .A(n18709), .B(n18708), .ZN(
        P3_U2947) );
  NAND2_X1 U20795 ( .A1(n18726), .A2(n18723), .ZN(n19060) );
  NOR2_X1 U20796 ( .A1(n21273), .A2(n18710), .ZN(n19055) );
  AOI22_X1 U20797 ( .A1(n18757), .A2(n19073), .B1(n18754), .B2(n19055), .ZN(
        n18713) );
  NAND2_X1 U20798 ( .A1(n19054), .A2(n19060), .ZN(n18718) );
  AOI21_X1 U20799 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19013), .ZN(n18749) );
  INV_X1 U20800 ( .A(n18710), .ZN(n18711) );
  AOI22_X1 U20801 ( .A1(n19011), .A2(n18718), .B1(n18749), .B2(n18711), .ZN(
        n19057) );
  AOI22_X1 U20802 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19057), .B1(
        n18756), .B2(n19056), .ZN(n18712) );
  OAI211_X1 U20803 ( .C1(n18748), .C2(n19054), .A(n18713), .B(n18712), .ZN(
        P3_U2939) );
  NAND2_X1 U20804 ( .A1(n21243), .A2(n18723), .ZN(n19066) );
  NOR2_X1 U20805 ( .A1(n21273), .A2(n18714), .ZN(n19061) );
  AOI22_X1 U20806 ( .A1(n18755), .A2(n19073), .B1(n18754), .B2(n19061), .ZN(
        n18716) );
  NAND2_X1 U20807 ( .A1(n18732), .A2(n18723), .ZN(n19063) );
  AOI22_X1 U20808 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19063), .B1(
        n18756), .B2(n19062), .ZN(n18715) );
  OAI211_X1 U20809 ( .C1(n18735), .C2(n19066), .A(n18716), .B(n18715), .ZN(
        P3_U2931) );
  NOR2_X2 U20810 ( .A1(n21233), .A2(n18741), .ZN(n19084) );
  NOR2_X1 U20811 ( .A1(n19079), .A2(n19084), .ZN(n18727) );
  OAI22_X1 U20812 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19060), .B1(n18727), 
        .B2(n18736), .ZN(n18717) );
  OAI21_X1 U20813 ( .B1(n19069), .B2(n18717), .A(n18966), .ZN(n19068) );
  AND2_X1 U20814 ( .A1(n21259), .A2(n18718), .ZN(n19067) );
  AOI22_X1 U20815 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19068), .B1(
        n18754), .B2(n19067), .ZN(n18720) );
  AOI22_X1 U20816 ( .A1(n18757), .A2(n19084), .B1(n18756), .B2(n19069), .ZN(
        n18719) );
  OAI211_X1 U20817 ( .C1(n18748), .C2(n19066), .A(n18720), .B(n18719), .ZN(
        P3_U2923) );
  NOR2_X1 U20818 ( .A1(n21234), .A2(n18741), .ZN(n18731) );
  NAND2_X1 U20819 ( .A1(n18731), .A2(n18721), .ZN(n18993) );
  INV_X1 U20820 ( .A(n18723), .ZN(n18722) );
  NOR2_X1 U20821 ( .A1(n18722), .A2(n18742), .ZN(n19072) );
  AOI22_X1 U20822 ( .A1(n18755), .A2(n19084), .B1(n18754), .B2(n19072), .ZN(
        n18725) );
  AOI22_X1 U20823 ( .A1(n19011), .A2(n18731), .B1(n18744), .B2(n18723), .ZN(
        n19074) );
  AOI22_X1 U20824 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19074), .B1(
        n18756), .B2(n19073), .ZN(n18724) );
  OAI211_X1 U20825 ( .C1(n18735), .C2(n18993), .A(n18725), .B(n18724), .ZN(
        P3_U2915) );
  NAND2_X1 U20826 ( .A1(n18726), .A2(n18743), .ZN(n19088) );
  NOR2_X1 U20827 ( .A1(n21273), .A2(n18727), .ZN(n19078) );
  AOI22_X1 U20828 ( .A1(n18755), .A2(n19091), .B1(n18754), .B2(n19078), .ZN(
        n18730) );
  NAND2_X1 U20829 ( .A1(n18993), .A2(n19088), .ZN(n18738) );
  INV_X1 U20830 ( .A(n18727), .ZN(n18728) );
  AOI22_X1 U20831 ( .A1(n19011), .A2(n18738), .B1(n18749), .B2(n18728), .ZN(
        n19080) );
  AOI22_X1 U20832 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19080), .B1(
        n18756), .B2(n19079), .ZN(n18729) );
  OAI211_X1 U20833 ( .C1(n18735), .C2(n19088), .A(n18730), .B(n18729), .ZN(
        P3_U2907) );
  NAND2_X1 U20834 ( .A1(n21243), .A2(n18743), .ZN(n18951) );
  INV_X1 U20835 ( .A(n19088), .ZN(n19098) );
  AND2_X1 U20836 ( .A1(n21259), .A2(n18731), .ZN(n19083) );
  AOI22_X1 U20837 ( .A1(n18755), .A2(n19098), .B1(n18754), .B2(n19083), .ZN(
        n18734) );
  NAND2_X1 U20838 ( .A1(n18732), .A2(n18743), .ZN(n19085) );
  AOI22_X1 U20839 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19085), .B1(
        n18756), .B2(n19084), .ZN(n18733) );
  OAI211_X1 U20840 ( .C1(n18735), .C2(n18951), .A(n18734), .B(n18733), .ZN(
        P3_U2899) );
  NOR2_X1 U20841 ( .A1(n19097), .A2(n19109), .ZN(n18753) );
  OAI22_X1 U20842 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19088), .B1(n18753), 
        .B2(n18736), .ZN(n18737) );
  OAI21_X1 U20843 ( .B1(n19091), .B2(n18737), .A(n18966), .ZN(n19090) );
  AND2_X1 U20844 ( .A1(n21259), .A2(n18738), .ZN(n19089) );
  AOI22_X1 U20845 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19090), .B1(
        n18754), .B2(n19089), .ZN(n18740) );
  AOI22_X1 U20846 ( .A1(n18757), .A2(n19097), .B1(n18756), .B2(n19091), .ZN(
        n18739) );
  OAI211_X1 U20847 ( .C1(n18748), .C2(n18951), .A(n18740), .B(n18739), .ZN(
        P3_U2891) );
  NOR2_X1 U20848 ( .A1(n18742), .A2(n18741), .ZN(n19095) );
  AOI22_X1 U20849 ( .A1(n18757), .A2(n19022), .B1(n18754), .B2(n19095), .ZN(
        n18747) );
  AOI22_X1 U20850 ( .A1(n19011), .A2(n18745), .B1(n18744), .B2(n18743), .ZN(
        n19099) );
  AOI22_X1 U20851 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19099), .B1(
        n18756), .B2(n19098), .ZN(n18746) );
  OAI211_X1 U20852 ( .C1(n19094), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        P3_U2883) );
  NOR2_X1 U20853 ( .A1(n10969), .A2(n19022), .ZN(n18752) );
  INV_X1 U20854 ( .A(n18749), .ZN(n18750) );
  OAI22_X1 U20855 ( .A1(n18752), .A2(n18751), .B1(n18753), .B2(n18750), .ZN(
        n19107) );
  NOR2_X1 U20856 ( .A1(n21273), .A2(n18753), .ZN(n19104) );
  AOI22_X1 U20857 ( .A1(n18755), .A2(n19022), .B1(n18754), .B2(n19104), .ZN(
        n18759) );
  AOI22_X1 U20858 ( .A1(n18757), .A2(n10969), .B1(n18756), .B2(n19109), .ZN(
        n18758) );
  OAI211_X1 U20859 ( .C1(n18760), .C2(n19107), .A(n18759), .B(n18758), .ZN(
        P3_U2875) );
  INV_X1 U20860 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n18761) );
  AOI22_X1 U20861 ( .A1(n19010), .A2(n18761), .B1(n20595), .B2(U215), .ZN(U257) );
  NAND2_X1 U20862 ( .A1(n19011), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18790) );
  NAND2_X1 U20863 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19011), .ZN(n18793) );
  INV_X1 U20864 ( .A(n18793), .ZN(n18795) );
  NOR2_X2 U20865 ( .A1(n19013), .A2(n20595), .ZN(n18794) );
  AOI22_X1 U20866 ( .A1(n19032), .A2(n18795), .B1(n19014), .B2(n18794), .ZN(
        n18763) );
  NOR2_X2 U20867 ( .A1(n20799), .A2(n19015), .ZN(n18796) );
  AOI22_X1 U20868 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18796), .ZN(n18762) );
  OAI211_X1 U20869 ( .C1(n19020), .C2(n18790), .A(n18763), .B(n18762), .ZN(
        P3_U2994) );
  AOI22_X1 U20870 ( .A1(n19038), .A2(n18795), .B1(n19021), .B2(n18794), .ZN(
        n18765) );
  AOI22_X1 U20871 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n18796), .ZN(n18764) );
  OAI211_X1 U20872 ( .C1(n18969), .C2(n18790), .A(n18765), .B(n18764), .ZN(
        P3_U2986) );
  INV_X1 U20873 ( .A(n18790), .ZN(n18797) );
  AOI22_X1 U20874 ( .A1(n19038), .A2(n18797), .B1(n19026), .B2(n18794), .ZN(
        n18767) );
  AOI22_X1 U20875 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n18796), .ZN(n18766) );
  OAI211_X1 U20876 ( .C1(n19036), .C2(n18793), .A(n18767), .B(n18766), .ZN(
        P3_U2978) );
  AOI22_X1 U20877 ( .A1(n19050), .A2(n18795), .B1(n19031), .B2(n18794), .ZN(
        n18769) );
  AOI22_X1 U20878 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18796), .ZN(n18768) );
  OAI211_X1 U20879 ( .C1(n19036), .C2(n18790), .A(n18769), .B(n18768), .ZN(
        P3_U2970) );
  AOI22_X1 U20880 ( .A1(n19056), .A2(n18795), .B1(n19037), .B2(n18794), .ZN(
        n18771) );
  AOI22_X1 U20881 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n18796), .ZN(n18770) );
  OAI211_X1 U20882 ( .C1(n19042), .C2(n18790), .A(n18771), .B(n18770), .ZN(
        P3_U2962) );
  AOI22_X1 U20883 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19045), .B1(
        n19043), .B2(n18794), .ZN(n18773) );
  AOI22_X1 U20884 ( .A1(n19044), .A2(n18796), .B1(n19056), .B2(n18797), .ZN(
        n18772) );
  OAI211_X1 U20885 ( .C1(n19048), .C2(n18793), .A(n18773), .B(n18772), .ZN(
        P3_U2954) );
  AOI22_X1 U20886 ( .A1(n19069), .A2(n18795), .B1(n19049), .B2(n18794), .ZN(
        n18775) );
  AOI22_X1 U20887 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n18796), .ZN(n18774) );
  OAI211_X1 U20888 ( .C1(n19048), .C2(n18790), .A(n18775), .B(n18774), .ZN(
        P3_U2946) );
  AOI22_X1 U20889 ( .A1(n19069), .A2(n18797), .B1(n19055), .B2(n18794), .ZN(
        n18777) );
  AOI22_X1 U20890 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18796), .ZN(n18776) );
  OAI211_X1 U20891 ( .C1(n19060), .C2(n18793), .A(n18777), .B(n18776), .ZN(
        P3_U2938) );
  AOI22_X1 U20892 ( .A1(n19073), .A2(n18797), .B1(n19061), .B2(n18794), .ZN(
        n18779) );
  AOI22_X1 U20893 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n18796), .ZN(n18778) );
  OAI211_X1 U20894 ( .C1(n19066), .C2(n18793), .A(n18779), .B(n18778), .ZN(
        P3_U2930) );
  AOI22_X1 U20895 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19068), .B1(
        n19067), .B2(n18794), .ZN(n18781) );
  AOI22_X1 U20896 ( .A1(n19069), .A2(n18796), .B1(n19084), .B2(n18795), .ZN(
        n18780) );
  OAI211_X1 U20897 ( .C1(n19066), .C2(n18790), .A(n18781), .B(n18780), .ZN(
        P3_U2922) );
  AOI22_X1 U20898 ( .A1(n19084), .A2(n18797), .B1(n19072), .B2(n18794), .ZN(
        n18783) );
  AOI22_X1 U20899 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n18796), .ZN(n18782) );
  OAI211_X1 U20900 ( .C1(n18993), .C2(n18793), .A(n18783), .B(n18782), .ZN(
        P3_U2914) );
  AOI22_X1 U20901 ( .A1(n19091), .A2(n18797), .B1(n19078), .B2(n18794), .ZN(
        n18785) );
  AOI22_X1 U20902 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18796), .ZN(n18784) );
  OAI211_X1 U20903 ( .C1(n19088), .C2(n18793), .A(n18785), .B(n18784), .ZN(
        P3_U2906) );
  AOI22_X1 U20904 ( .A1(n19098), .A2(n18797), .B1(n19083), .B2(n18794), .ZN(
        n18787) );
  AOI22_X1 U20905 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n18796), .ZN(n18786) );
  OAI211_X1 U20906 ( .C1(n18951), .C2(n18793), .A(n18787), .B(n18786), .ZN(
        P3_U2898) );
  AOI22_X1 U20907 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18794), .ZN(n18789) );
  AOI22_X1 U20908 ( .A1(n19097), .A2(n18795), .B1(n19091), .B2(n18796), .ZN(
        n18788) );
  OAI211_X1 U20909 ( .C1(n18951), .C2(n18790), .A(n18789), .B(n18788), .ZN(
        P3_U2890) );
  AOI22_X1 U20910 ( .A1(n19097), .A2(n18797), .B1(n19095), .B2(n18794), .ZN(
        n18792) );
  AOI22_X1 U20911 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n18796), .ZN(n18791) );
  OAI211_X1 U20912 ( .C1(n19114), .C2(n18793), .A(n18792), .B(n18791), .ZN(
        P3_U2882) );
  AOI22_X1 U20913 ( .A1(n10969), .A2(n18795), .B1(n19104), .B2(n18794), .ZN(
        n18799) );
  AOI22_X1 U20914 ( .A1(n19022), .A2(n18797), .B1(n19109), .B2(n18796), .ZN(
        n18798) );
  OAI211_X1 U20915 ( .C1(n18800), .C2(n19107), .A(n18799), .B(n18798), .ZN(
        P3_U2874) );
  INV_X1 U20916 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n18801) );
  INV_X1 U20917 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20599) );
  AOI22_X1 U20918 ( .A1(n18964), .A2(n18801), .B1(n20599), .B2(U215), .ZN(U256) );
  NAND2_X1 U20919 ( .A1(n19011), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18834) );
  NAND2_X1 U20920 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19011), .ZN(n18829) );
  INV_X1 U20921 ( .A(n18829), .ZN(n18836) );
  NOR2_X2 U20922 ( .A1(n19013), .A2(n20599), .ZN(n18835) );
  AOI22_X1 U20923 ( .A1(n19032), .A2(n18836), .B1(n19014), .B2(n18835), .ZN(
        n18804) );
  NOR2_X2 U20924 ( .A1(n18802), .A2(n19015), .ZN(n18837) );
  AOI22_X1 U20925 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18837), .ZN(n18803) );
  OAI211_X1 U20926 ( .C1(n19020), .C2(n18834), .A(n18804), .B(n18803), .ZN(
        P3_U2993) );
  AOI22_X1 U20927 ( .A1(n19032), .A2(n18838), .B1(n19021), .B2(n18835), .ZN(
        n18806) );
  AOI22_X1 U20928 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n18837), .ZN(n18805) );
  OAI211_X1 U20929 ( .C1(n19030), .C2(n18829), .A(n18806), .B(n18805), .ZN(
        P3_U2985) );
  AOI22_X1 U20930 ( .A1(n19044), .A2(n18836), .B1(n19026), .B2(n18835), .ZN(
        n18808) );
  AOI22_X1 U20931 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n18837), .ZN(n18807) );
  OAI211_X1 U20932 ( .C1(n19030), .C2(n18834), .A(n18808), .B(n18807), .ZN(
        P3_U2977) );
  AOI22_X1 U20933 ( .A1(n19044), .A2(n18838), .B1(n19031), .B2(n18835), .ZN(
        n18810) );
  AOI22_X1 U20934 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18837), .ZN(n18809) );
  OAI211_X1 U20935 ( .C1(n19042), .C2(n18829), .A(n18810), .B(n18809), .ZN(
        P3_U2969) );
  AOI22_X1 U20936 ( .A1(n19056), .A2(n18836), .B1(n19037), .B2(n18835), .ZN(
        n18812) );
  AOI22_X1 U20937 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n18837), .ZN(n18811) );
  OAI211_X1 U20938 ( .C1(n19042), .C2(n18834), .A(n18812), .B(n18811), .ZN(
        P3_U2961) );
  AOI22_X1 U20939 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19045), .B1(
        n19043), .B2(n18835), .ZN(n18814) );
  AOI22_X1 U20940 ( .A1(n19044), .A2(n18837), .B1(n19056), .B2(n18838), .ZN(
        n18813) );
  OAI211_X1 U20941 ( .C1(n19048), .C2(n18829), .A(n18814), .B(n18813), .ZN(
        P3_U2953) );
  AOI22_X1 U20942 ( .A1(n19069), .A2(n18836), .B1(n19049), .B2(n18835), .ZN(
        n18816) );
  AOI22_X1 U20943 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n18837), .ZN(n18815) );
  OAI211_X1 U20944 ( .C1(n19048), .C2(n18834), .A(n18816), .B(n18815), .ZN(
        P3_U2945) );
  AOI22_X1 U20945 ( .A1(n19069), .A2(n18838), .B1(n19055), .B2(n18835), .ZN(
        n18818) );
  AOI22_X1 U20946 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18837), .ZN(n18817) );
  OAI211_X1 U20947 ( .C1(n19060), .C2(n18829), .A(n18818), .B(n18817), .ZN(
        P3_U2937) );
  AOI22_X1 U20948 ( .A1(n19073), .A2(n18838), .B1(n19061), .B2(n18835), .ZN(
        n18820) );
  AOI22_X1 U20949 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n18837), .ZN(n18819) );
  OAI211_X1 U20950 ( .C1(n19066), .C2(n18829), .A(n18820), .B(n18819), .ZN(
        P3_U2929) );
  INV_X1 U20951 ( .A(n19084), .ZN(n19077) );
  AOI22_X1 U20952 ( .A1(n19079), .A2(n18838), .B1(n19067), .B2(n18835), .ZN(
        n18822) );
  AOI22_X1 U20953 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19068), .B1(
        n19069), .B2(n18837), .ZN(n18821) );
  OAI211_X1 U20954 ( .C1(n19077), .C2(n18829), .A(n18822), .B(n18821), .ZN(
        P3_U2921) );
  AOI22_X1 U20955 ( .A1(n19091), .A2(n18836), .B1(n19072), .B2(n18835), .ZN(
        n18824) );
  AOI22_X1 U20956 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n18837), .ZN(n18823) );
  OAI211_X1 U20957 ( .C1(n19077), .C2(n18834), .A(n18824), .B(n18823), .ZN(
        P3_U2913) );
  AOI22_X1 U20958 ( .A1(n19091), .A2(n18838), .B1(n19078), .B2(n18835), .ZN(
        n18826) );
  AOI22_X1 U20959 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18837), .ZN(n18825) );
  OAI211_X1 U20960 ( .C1(n19088), .C2(n18829), .A(n18826), .B(n18825), .ZN(
        P3_U2905) );
  AOI22_X1 U20961 ( .A1(n19098), .A2(n18838), .B1(n19083), .B2(n18835), .ZN(
        n18828) );
  AOI22_X1 U20962 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n18837), .ZN(n18827) );
  OAI211_X1 U20963 ( .C1(n18951), .C2(n18829), .A(n18828), .B(n18827), .ZN(
        P3_U2897) );
  AOI22_X1 U20964 ( .A1(n19097), .A2(n18836), .B1(n19089), .B2(n18835), .ZN(
        n18831) );
  AOI22_X1 U20965 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19090), .B1(
        n19091), .B2(n18837), .ZN(n18830) );
  OAI211_X1 U20966 ( .C1(n18951), .C2(n18834), .A(n18831), .B(n18830), .ZN(
        P3_U2889) );
  AOI22_X1 U20967 ( .A1(n19022), .A2(n18836), .B1(n19095), .B2(n18835), .ZN(
        n18833) );
  AOI22_X1 U20968 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n18837), .ZN(n18832) );
  OAI211_X1 U20969 ( .C1(n19094), .C2(n18834), .A(n18833), .B(n18832), .ZN(
        P3_U2881) );
  AOI22_X1 U20970 ( .A1(n10969), .A2(n18836), .B1(n19104), .B2(n18835), .ZN(
        n18840) );
  AOI22_X1 U20971 ( .A1(n19022), .A2(n18838), .B1(n19109), .B2(n18837), .ZN(
        n18839) );
  OAI211_X1 U20972 ( .C1(n18841), .C2(n19107), .A(n18840), .B(n18839), .ZN(
        P3_U2873) );
  INV_X1 U20973 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n18842) );
  AOI22_X1 U20974 ( .A1(n18964), .A2(n18842), .B1(n20604), .B2(U215), .ZN(U255) );
  NAND2_X1 U20975 ( .A1(n19011), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18871) );
  AND2_X1 U20976 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19011), .ZN(n18876) );
  NOR2_X2 U20977 ( .A1(n19013), .A2(n20604), .ZN(n18875) );
  AOI22_X1 U20978 ( .A1(n19032), .A2(n18876), .B1(n19014), .B2(n18875), .ZN(
        n18844) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18877), .ZN(n18843) );
  OAI211_X1 U20980 ( .C1(n19020), .C2(n18871), .A(n18844), .B(n18843), .ZN(
        P3_U2992) );
  AOI22_X1 U20981 ( .A1(n19038), .A2(n18876), .B1(n19021), .B2(n18875), .ZN(
        n18846) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n18877), .ZN(n18845) );
  OAI211_X1 U20983 ( .C1(n18969), .C2(n18871), .A(n18846), .B(n18845), .ZN(
        P3_U2984) );
  AOI22_X1 U20984 ( .A1(n19044), .A2(n18876), .B1(n19026), .B2(n18875), .ZN(
        n18848) );
  AOI22_X1 U20985 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19027), .B1(
        n18877), .B2(n10969), .ZN(n18847) );
  OAI211_X1 U20986 ( .C1(n19030), .C2(n18871), .A(n18848), .B(n18847), .ZN(
        P3_U2976) );
  AOI22_X1 U20987 ( .A1(n19050), .A2(n18876), .B1(n19031), .B2(n18875), .ZN(
        n18850) );
  AOI22_X1 U20988 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18877), .ZN(n18849) );
  OAI211_X1 U20989 ( .C1(n19036), .C2(n18871), .A(n18850), .B(n18849), .ZN(
        P3_U2968) );
  INV_X1 U20990 ( .A(n18877), .ZN(n18874) );
  INV_X1 U20991 ( .A(n18871), .ZN(n18878) );
  AOI22_X1 U20992 ( .A1(n19050), .A2(n18878), .B1(n19037), .B2(n18875), .ZN(
        n18852) );
  AOI22_X1 U20993 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19039), .B1(
        n19056), .B2(n18876), .ZN(n18851) );
  OAI211_X1 U20994 ( .C1(n19030), .C2(n18874), .A(n18852), .B(n18851), .ZN(
        P3_U2960) );
  AOI22_X1 U20995 ( .A1(n19056), .A2(n18878), .B1(n19043), .B2(n18875), .ZN(
        n18854) );
  AOI22_X1 U20996 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19045), .B1(
        n19062), .B2(n18876), .ZN(n18853) );
  OAI211_X1 U20997 ( .C1(n19036), .C2(n18874), .A(n18854), .B(n18853), .ZN(
        P3_U2952) );
  AOI22_X1 U20998 ( .A1(n19069), .A2(n18876), .B1(n19049), .B2(n18875), .ZN(
        n18856) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n18877), .ZN(n18855) );
  OAI211_X1 U21000 ( .C1(n19048), .C2(n18871), .A(n18856), .B(n18855), .ZN(
        P3_U2944) );
  AOI22_X1 U21001 ( .A1(n19073), .A2(n18876), .B1(n19055), .B2(n18875), .ZN(
        n18858) );
  AOI22_X1 U21002 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18877), .ZN(n18857) );
  OAI211_X1 U21003 ( .C1(n19054), .C2(n18871), .A(n18858), .B(n18857), .ZN(
        P3_U2936) );
  AOI22_X1 U21004 ( .A1(n19079), .A2(n18876), .B1(n19061), .B2(n18875), .ZN(
        n18860) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n18877), .ZN(n18859) );
  OAI211_X1 U21006 ( .C1(n19060), .C2(n18871), .A(n18860), .B(n18859), .ZN(
        P3_U2928) );
  AOI22_X1 U21007 ( .A1(n19079), .A2(n18878), .B1(n19067), .B2(n18875), .ZN(
        n18862) );
  AOI22_X1 U21008 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19068), .B1(
        n19084), .B2(n18876), .ZN(n18861) );
  OAI211_X1 U21009 ( .C1(n19054), .C2(n18874), .A(n18862), .B(n18861), .ZN(
        P3_U2920) );
  AOI22_X1 U21010 ( .A1(n19084), .A2(n18878), .B1(n19072), .B2(n18875), .ZN(
        n18864) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19074), .B1(
        n19091), .B2(n18876), .ZN(n18863) );
  OAI211_X1 U21012 ( .C1(n19060), .C2(n18874), .A(n18864), .B(n18863), .ZN(
        P3_U2912) );
  AOI22_X1 U21013 ( .A1(n19098), .A2(n18876), .B1(n19078), .B2(n18875), .ZN(
        n18866) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18877), .ZN(n18865) );
  OAI211_X1 U21015 ( .C1(n18993), .C2(n18871), .A(n18866), .B(n18865), .ZN(
        P3_U2904) );
  AOI22_X1 U21016 ( .A1(n19109), .A2(n18876), .B1(n19083), .B2(n18875), .ZN(
        n18868) );
  AOI22_X1 U21017 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n18877), .ZN(n18867) );
  OAI211_X1 U21018 ( .C1(n19088), .C2(n18871), .A(n18868), .B(n18867), .ZN(
        P3_U2896) );
  AOI22_X1 U21019 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18875), .ZN(n18870) );
  AOI22_X1 U21020 ( .A1(n19097), .A2(n18876), .B1(n19091), .B2(n18877), .ZN(
        n18869) );
  OAI211_X1 U21021 ( .C1(n18951), .C2(n18871), .A(n18870), .B(n18869), .ZN(
        P3_U2888) );
  AOI22_X1 U21022 ( .A1(n19097), .A2(n18878), .B1(n19095), .B2(n18875), .ZN(
        n18873) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19099), .B1(
        n19022), .B2(n18876), .ZN(n18872) );
  OAI211_X1 U21024 ( .C1(n19088), .C2(n18874), .A(n18873), .B(n18872), .ZN(
        P3_U2880) );
  AOI22_X1 U21025 ( .A1(n10969), .A2(n18876), .B1(n19104), .B2(n18875), .ZN(
        n18880) );
  AOI22_X1 U21026 ( .A1(n19022), .A2(n18878), .B1(n19109), .B2(n18877), .ZN(
        n18879) );
  OAI211_X1 U21027 ( .C1(n18881), .C2(n19107), .A(n18880), .B(n18879), .ZN(
        P3_U2872) );
  INV_X1 U21028 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n18882) );
  INV_X1 U21029 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20608) );
  AOI22_X1 U21030 ( .A1(n18964), .A2(n18882), .B1(n20608), .B2(U215), .ZN(U254) );
  NAND2_X1 U21031 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19011), .ZN(n18910) );
  NAND2_X1 U21032 ( .A1(n19011), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18915) );
  INV_X1 U21033 ( .A(n18915), .ZN(n18917) );
  NOR2_X2 U21034 ( .A1(n19013), .A2(n20608), .ZN(n18916) );
  AOI22_X1 U21035 ( .A1(n10969), .A2(n18917), .B1(n19014), .B2(n18916), .ZN(
        n18885) );
  NOR2_X2 U21036 ( .A1(n18883), .A2(n19015), .ZN(n18918) );
  AOI22_X1 U21037 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18918), .ZN(n18884) );
  OAI211_X1 U21038 ( .C1(n18969), .C2(n18910), .A(n18885), .B(n18884), .ZN(
        P3_U2991) );
  INV_X1 U21039 ( .A(n18910), .ZN(n18919) );
  AOI22_X1 U21040 ( .A1(n19038), .A2(n18919), .B1(n19021), .B2(n18916), .ZN(
        n18887) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n18918), .ZN(n18886) );
  OAI211_X1 U21042 ( .C1(n18969), .C2(n18915), .A(n18887), .B(n18886), .ZN(
        P3_U2983) );
  AOI22_X1 U21043 ( .A1(n19038), .A2(n18917), .B1(n19026), .B2(n18916), .ZN(
        n18889) );
  AOI22_X1 U21044 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n18918), .ZN(n18888) );
  OAI211_X1 U21045 ( .C1(n19036), .C2(n18910), .A(n18889), .B(n18888), .ZN(
        P3_U2975) );
  AOI22_X1 U21046 ( .A1(n19050), .A2(n18919), .B1(n19031), .B2(n18916), .ZN(
        n18891) );
  AOI22_X1 U21047 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18918), .ZN(n18890) );
  OAI211_X1 U21048 ( .C1(n19036), .C2(n18915), .A(n18891), .B(n18890), .ZN(
        P3_U2967) );
  AOI22_X1 U21049 ( .A1(n19056), .A2(n18919), .B1(n19037), .B2(n18916), .ZN(
        n18893) );
  AOI22_X1 U21050 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n18918), .ZN(n18892) );
  OAI211_X1 U21051 ( .C1(n19042), .C2(n18915), .A(n18893), .B(n18892), .ZN(
        P3_U2959) );
  AOI22_X1 U21052 ( .A1(n19062), .A2(n18919), .B1(n19043), .B2(n18916), .ZN(
        n18895) );
  AOI22_X1 U21053 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19045), .B1(
        n19044), .B2(n18918), .ZN(n18894) );
  OAI211_X1 U21054 ( .C1(n18980), .C2(n18915), .A(n18895), .B(n18894), .ZN(
        P3_U2951) );
  AOI22_X1 U21055 ( .A1(n19069), .A2(n18919), .B1(n19049), .B2(n18916), .ZN(
        n18897) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n18918), .ZN(n18896) );
  OAI211_X1 U21057 ( .C1(n19048), .C2(n18915), .A(n18897), .B(n18896), .ZN(
        P3_U2943) );
  AOI22_X1 U21058 ( .A1(n19073), .A2(n18919), .B1(n19055), .B2(n18916), .ZN(
        n18899) );
  AOI22_X1 U21059 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18918), .ZN(n18898) );
  OAI211_X1 U21060 ( .C1(n19054), .C2(n18915), .A(n18899), .B(n18898), .ZN(
        P3_U2935) );
  AOI22_X1 U21061 ( .A1(n19073), .A2(n18917), .B1(n19061), .B2(n18916), .ZN(
        n18901) );
  AOI22_X1 U21062 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n18918), .ZN(n18900) );
  OAI211_X1 U21063 ( .C1(n19066), .C2(n18910), .A(n18901), .B(n18900), .ZN(
        P3_U2927) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19068), .B1(
        n19067), .B2(n18916), .ZN(n18903) );
  AOI22_X1 U21065 ( .A1(n19069), .A2(n18918), .B1(n19084), .B2(n18919), .ZN(
        n18902) );
  OAI211_X1 U21066 ( .C1(n19066), .C2(n18915), .A(n18903), .B(n18902), .ZN(
        P3_U2919) );
  AOI22_X1 U21067 ( .A1(n19084), .A2(n18917), .B1(n19072), .B2(n18916), .ZN(
        n18905) );
  AOI22_X1 U21068 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n18918), .ZN(n18904) );
  OAI211_X1 U21069 ( .C1(n18993), .C2(n18910), .A(n18905), .B(n18904), .ZN(
        P3_U2911) );
  AOI22_X1 U21070 ( .A1(n19098), .A2(n18919), .B1(n19078), .B2(n18916), .ZN(
        n18907) );
  AOI22_X1 U21071 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18918), .ZN(n18906) );
  OAI211_X1 U21072 ( .C1(n18993), .C2(n18915), .A(n18907), .B(n18906), .ZN(
        P3_U2903) );
  AOI22_X1 U21073 ( .A1(n19098), .A2(n18917), .B1(n19083), .B2(n18916), .ZN(
        n18909) );
  AOI22_X1 U21074 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n18918), .ZN(n18908) );
  OAI211_X1 U21075 ( .C1(n18951), .C2(n18910), .A(n18909), .B(n18908), .ZN(
        P3_U2895) );
  AOI22_X1 U21076 ( .A1(n19097), .A2(n18919), .B1(n19089), .B2(n18916), .ZN(
        n18912) );
  AOI22_X1 U21077 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19090), .B1(
        n19091), .B2(n18918), .ZN(n18911) );
  OAI211_X1 U21078 ( .C1(n18951), .C2(n18915), .A(n18912), .B(n18911), .ZN(
        P3_U2887) );
  AOI22_X1 U21079 ( .A1(n19022), .A2(n18919), .B1(n19095), .B2(n18916), .ZN(
        n18914) );
  AOI22_X1 U21080 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n18918), .ZN(n18913) );
  OAI211_X1 U21081 ( .C1(n19094), .C2(n18915), .A(n18914), .B(n18913), .ZN(
        P3_U2879) );
  AOI22_X1 U21082 ( .A1(n19022), .A2(n18917), .B1(n19104), .B2(n18916), .ZN(
        n18921) );
  AOI22_X1 U21083 ( .A1(n10969), .A2(n18919), .B1(n19109), .B2(n18918), .ZN(
        n18920) );
  OAI211_X1 U21084 ( .C1(n18922), .C2(n19107), .A(n18921), .B(n18920), .ZN(
        P3_U2871) );
  INV_X1 U21085 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n18923) );
  INV_X1 U21086 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U21087 ( .A1(n18964), .A2(n18923), .B1(n20614), .B2(U215), .ZN(U253) );
  NAND2_X1 U21088 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19011), .ZN(n18956) );
  NAND2_X1 U21089 ( .A1(n19011), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18942) );
  INV_X1 U21090 ( .A(n18942), .ZN(n18960) );
  NOR2_X2 U21091 ( .A1(n19013), .A2(n20614), .ZN(n18957) );
  AOI22_X1 U21092 ( .A1(n10969), .A2(n18960), .B1(n19014), .B2(n18957), .ZN(
        n18925) );
  NOR2_X2 U21093 ( .A1(n20807), .A2(n19015), .ZN(n18959) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n18959), .ZN(n18924) );
  OAI211_X1 U21095 ( .C1(n18969), .C2(n18956), .A(n18925), .B(n18924), .ZN(
        P3_U2990) );
  INV_X1 U21096 ( .A(n18956), .ZN(n18958) );
  AOI22_X1 U21097 ( .A1(n19038), .A2(n18958), .B1(n19021), .B2(n18957), .ZN(
        n18927) );
  AOI22_X1 U21098 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n18959), .ZN(n18926) );
  OAI211_X1 U21099 ( .C1(n18969), .C2(n18942), .A(n18927), .B(n18926), .ZN(
        P3_U2982) );
  AOI22_X1 U21100 ( .A1(n19044), .A2(n18958), .B1(n19026), .B2(n18957), .ZN(
        n18929) );
  AOI22_X1 U21101 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n18959), .ZN(n18928) );
  OAI211_X1 U21102 ( .C1(n19030), .C2(n18942), .A(n18929), .B(n18928), .ZN(
        P3_U2974) );
  AOI22_X1 U21103 ( .A1(n19050), .A2(n18958), .B1(n19031), .B2(n18957), .ZN(
        n18931) );
  AOI22_X1 U21104 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n18959), .ZN(n18930) );
  OAI211_X1 U21105 ( .C1(n19036), .C2(n18942), .A(n18931), .B(n18930), .ZN(
        P3_U2966) );
  AOI22_X1 U21106 ( .A1(n19050), .A2(n18960), .B1(n19037), .B2(n18957), .ZN(
        n18933) );
  AOI22_X1 U21107 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n18959), .ZN(n18932) );
  OAI211_X1 U21108 ( .C1(n18980), .C2(n18956), .A(n18933), .B(n18932), .ZN(
        P3_U2958) );
  AOI22_X1 U21109 ( .A1(n19062), .A2(n18958), .B1(n19043), .B2(n18957), .ZN(
        n18935) );
  AOI22_X1 U21110 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19045), .B1(
        n19044), .B2(n18959), .ZN(n18934) );
  OAI211_X1 U21111 ( .C1(n18980), .C2(n18942), .A(n18935), .B(n18934), .ZN(
        P3_U2950) );
  AOI22_X1 U21112 ( .A1(n19062), .A2(n18960), .B1(n19049), .B2(n18957), .ZN(
        n18937) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n18959), .ZN(n18936) );
  OAI211_X1 U21114 ( .C1(n19054), .C2(n18956), .A(n18937), .B(n18936), .ZN(
        P3_U2942) );
  AOI22_X1 U21115 ( .A1(n19069), .A2(n18960), .B1(n19055), .B2(n18957), .ZN(
        n18939) );
  AOI22_X1 U21116 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n18959), .ZN(n18938) );
  OAI211_X1 U21117 ( .C1(n19060), .C2(n18956), .A(n18939), .B(n18938), .ZN(
        P3_U2934) );
  AOI22_X1 U21118 ( .A1(n19079), .A2(n18958), .B1(n19061), .B2(n18957), .ZN(
        n18941) );
  AOI22_X1 U21119 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n18959), .ZN(n18940) );
  OAI211_X1 U21120 ( .C1(n19060), .C2(n18942), .A(n18941), .B(n18940), .ZN(
        P3_U2926) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19068), .B1(
        n19067), .B2(n18957), .ZN(n18944) );
  AOI22_X1 U21122 ( .A1(n19069), .A2(n18959), .B1(n19079), .B2(n18960), .ZN(
        n18943) );
  OAI211_X1 U21123 ( .C1(n19077), .C2(n18956), .A(n18944), .B(n18943), .ZN(
        P3_U2918) );
  AOI22_X1 U21124 ( .A1(n19084), .A2(n18960), .B1(n19072), .B2(n18957), .ZN(
        n18946) );
  AOI22_X1 U21125 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n18959), .ZN(n18945) );
  OAI211_X1 U21126 ( .C1(n18993), .C2(n18956), .A(n18946), .B(n18945), .ZN(
        P3_U2910) );
  AOI22_X1 U21127 ( .A1(n19091), .A2(n18960), .B1(n19078), .B2(n18957), .ZN(
        n18948) );
  AOI22_X1 U21128 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n18959), .ZN(n18947) );
  OAI211_X1 U21129 ( .C1(n19088), .C2(n18956), .A(n18948), .B(n18947), .ZN(
        P3_U2902) );
  AOI22_X1 U21130 ( .A1(n19098), .A2(n18960), .B1(n19083), .B2(n18957), .ZN(
        n18950) );
  AOI22_X1 U21131 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n18959), .ZN(n18949) );
  OAI211_X1 U21132 ( .C1(n18951), .C2(n18956), .A(n18950), .B(n18949), .ZN(
        P3_U2894) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18957), .ZN(n18953) );
  AOI22_X1 U21134 ( .A1(n19091), .A2(n18959), .B1(n19109), .B2(n18960), .ZN(
        n18952) );
  OAI211_X1 U21135 ( .C1(n19094), .C2(n18956), .A(n18953), .B(n18952), .ZN(
        P3_U2886) );
  AOI22_X1 U21136 ( .A1(n19097), .A2(n18960), .B1(n19095), .B2(n18957), .ZN(
        n18955) );
  AOI22_X1 U21137 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n18959), .ZN(n18954) );
  OAI211_X1 U21138 ( .C1(n19114), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        P3_U2878) );
  AOI22_X1 U21139 ( .A1(n10969), .A2(n18958), .B1(n19104), .B2(n18957), .ZN(
        n18962) );
  AOI22_X1 U21140 ( .A1(n19022), .A2(n18960), .B1(n19109), .B2(n18959), .ZN(
        n18961) );
  OAI211_X1 U21141 ( .C1(n18963), .C2(n19107), .A(n18962), .B(n18961), .ZN(
        P3_U2870) );
  OAI22_X1 U21142 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18964), .ZN(n18965) );
  INV_X1 U21143 ( .A(n18965), .ZN(U252) );
  NAND2_X1 U21144 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19011), .ZN(n19001) );
  NAND2_X1 U21145 ( .A1(n19011), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18996) );
  INV_X1 U21146 ( .A(n18996), .ZN(n19005) );
  AND2_X1 U21147 ( .A1(n18966), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19002) );
  AOI22_X1 U21148 ( .A1(n10969), .A2(n19005), .B1(n19014), .B2(n19002), .ZN(
        n18968) );
  NOR2_X2 U21149 ( .A1(n20800), .A2(n19015), .ZN(n19004) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n19004), .ZN(n18967) );
  OAI211_X1 U21151 ( .C1(n18969), .C2(n19001), .A(n18968), .B(n18967), .ZN(
        P3_U2989) );
  AOI22_X1 U21152 ( .A1(n19032), .A2(n19005), .B1(n19021), .B2(n19002), .ZN(
        n18971) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n19004), .ZN(n18970) );
  OAI211_X1 U21154 ( .C1(n19030), .C2(n19001), .A(n18971), .B(n18970), .ZN(
        P3_U2981) );
  INV_X1 U21155 ( .A(n19001), .ZN(n19003) );
  AOI22_X1 U21156 ( .A1(n19044), .A2(n19003), .B1(n19026), .B2(n19002), .ZN(
        n18973) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n19004), .ZN(n18972) );
  OAI211_X1 U21158 ( .C1(n19030), .C2(n18996), .A(n18973), .B(n18972), .ZN(
        P3_U2973) );
  AOI22_X1 U21159 ( .A1(n19044), .A2(n19005), .B1(n19031), .B2(n19002), .ZN(
        n18975) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n19004), .ZN(n18974) );
  OAI211_X1 U21161 ( .C1(n19042), .C2(n19001), .A(n18975), .B(n18974), .ZN(
        P3_U2965) );
  AOI22_X1 U21162 ( .A1(n19056), .A2(n19003), .B1(n19037), .B2(n19002), .ZN(
        n18977) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n19004), .ZN(n18976) );
  OAI211_X1 U21164 ( .C1(n19042), .C2(n18996), .A(n18977), .B(n18976), .ZN(
        P3_U2957) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19045), .B1(
        n19043), .B2(n19002), .ZN(n18979) );
  AOI22_X1 U21166 ( .A1(n19044), .A2(n19004), .B1(n19062), .B2(n19003), .ZN(
        n18978) );
  OAI211_X1 U21167 ( .C1(n18980), .C2(n18996), .A(n18979), .B(n18978), .ZN(
        P3_U2949) );
  AOI22_X1 U21168 ( .A1(n19069), .A2(n19003), .B1(n19049), .B2(n19002), .ZN(
        n18982) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n19004), .ZN(n18981) );
  OAI211_X1 U21170 ( .C1(n19048), .C2(n18996), .A(n18982), .B(n18981), .ZN(
        P3_U2941) );
  AOI22_X1 U21171 ( .A1(n19073), .A2(n19003), .B1(n19055), .B2(n19002), .ZN(
        n18984) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n19004), .ZN(n18983) );
  OAI211_X1 U21173 ( .C1(n19054), .C2(n18996), .A(n18984), .B(n18983), .ZN(
        P3_U2933) );
  AOI22_X1 U21174 ( .A1(n19079), .A2(n19003), .B1(n19061), .B2(n19002), .ZN(
        n18986) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n19004), .ZN(n18985) );
  OAI211_X1 U21176 ( .C1(n19060), .C2(n18996), .A(n18986), .B(n18985), .ZN(
        P3_U2925) );
  AOI22_X1 U21177 ( .A1(n19079), .A2(n19005), .B1(n19067), .B2(n19002), .ZN(
        n18988) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19068), .B1(
        n19069), .B2(n19004), .ZN(n18987) );
  OAI211_X1 U21179 ( .C1(n19077), .C2(n19001), .A(n18988), .B(n18987), .ZN(
        P3_U2917) );
  AOI22_X1 U21180 ( .A1(n19091), .A2(n19003), .B1(n19072), .B2(n19002), .ZN(
        n18990) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n19004), .ZN(n18989) );
  OAI211_X1 U21182 ( .C1(n19077), .C2(n18996), .A(n18990), .B(n18989), .ZN(
        P3_U2909) );
  AOI22_X1 U21183 ( .A1(n19098), .A2(n19003), .B1(n19078), .B2(n19002), .ZN(
        n18992) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n19004), .ZN(n18991) );
  OAI211_X1 U21185 ( .C1(n18993), .C2(n18996), .A(n18992), .B(n18991), .ZN(
        P3_U2901) );
  AOI22_X1 U21186 ( .A1(n19109), .A2(n19003), .B1(n19083), .B2(n19002), .ZN(
        n18995) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n19004), .ZN(n18994) );
  OAI211_X1 U21188 ( .C1(n19088), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        P3_U2893) );
  AOI22_X1 U21189 ( .A1(n19109), .A2(n19005), .B1(n19089), .B2(n19002), .ZN(
        n18998) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19090), .B1(
        n19091), .B2(n19004), .ZN(n18997) );
  OAI211_X1 U21191 ( .C1(n19094), .C2(n19001), .A(n18998), .B(n18997), .ZN(
        P3_U2885) );
  AOI22_X1 U21192 ( .A1(n19097), .A2(n19005), .B1(n19095), .B2(n19002), .ZN(
        n19000) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n19004), .ZN(n18999) );
  OAI211_X1 U21194 ( .C1(n19114), .C2(n19001), .A(n19000), .B(n18999), .ZN(
        P3_U2877) );
  AOI22_X1 U21195 ( .A1(n10969), .A2(n19003), .B1(n19104), .B2(n19002), .ZN(
        n19007) );
  AOI22_X1 U21196 ( .A1(n19022), .A2(n19005), .B1(n19109), .B2(n19004), .ZN(
        n19006) );
  OAI211_X1 U21197 ( .C1(n19008), .C2(n19107), .A(n19007), .B(n19006), .ZN(
        P3_U2869) );
  INV_X1 U21198 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n19009) );
  AOI22_X1 U21199 ( .A1(n19010), .A2(n19009), .B1(n19012), .B2(U215), .ZN(U251) );
  NAND2_X1 U21200 ( .A1(n19011), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19113) );
  NAND2_X1 U21201 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19011), .ZN(n19102) );
  INV_X1 U21202 ( .A(n19102), .ZN(n19105) );
  NOR2_X2 U21203 ( .A1(n19013), .A2(n19012), .ZN(n19103) );
  AOI22_X1 U21204 ( .A1(n19032), .A2(n19105), .B1(n19014), .B2(n19103), .ZN(
        n19019) );
  NOR2_X2 U21205 ( .A1(n19016), .A2(n19015), .ZN(n19108) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19017), .B1(
        n19097), .B2(n19108), .ZN(n19018) );
  OAI211_X1 U21207 ( .C1(n19020), .C2(n19113), .A(n19019), .B(n19018), .ZN(
        P3_U2988) );
  INV_X1 U21208 ( .A(n19113), .ZN(n19096) );
  AOI22_X1 U21209 ( .A1(n19032), .A2(n19096), .B1(n19021), .B2(n19103), .ZN(
        n19025) );
  AOI22_X1 U21210 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19023), .B1(
        n19022), .B2(n19108), .ZN(n19024) );
  OAI211_X1 U21211 ( .C1(n19030), .C2(n19102), .A(n19025), .B(n19024), .ZN(
        P3_U2980) );
  AOI22_X1 U21212 ( .A1(n19044), .A2(n19105), .B1(n19026), .B2(n19103), .ZN(
        n19029) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19027), .B1(
        n10969), .B2(n19108), .ZN(n19028) );
  OAI211_X1 U21214 ( .C1(n19030), .C2(n19113), .A(n19029), .B(n19028), .ZN(
        P3_U2972) );
  AOI22_X1 U21215 ( .A1(n19050), .A2(n19105), .B1(n19031), .B2(n19103), .ZN(
        n19035) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19033), .B1(
        n19032), .B2(n19108), .ZN(n19034) );
  OAI211_X1 U21217 ( .C1(n19036), .C2(n19113), .A(n19035), .B(n19034), .ZN(
        P3_U2964) );
  AOI22_X1 U21218 ( .A1(n19056), .A2(n19105), .B1(n19037), .B2(n19103), .ZN(
        n19041) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19039), .B1(
        n19038), .B2(n19108), .ZN(n19040) );
  OAI211_X1 U21220 ( .C1(n19042), .C2(n19113), .A(n19041), .B(n19040), .ZN(
        P3_U2956) );
  AOI22_X1 U21221 ( .A1(n19056), .A2(n19096), .B1(n19043), .B2(n19103), .ZN(
        n19047) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19045), .B1(
        n19044), .B2(n19108), .ZN(n19046) );
  OAI211_X1 U21223 ( .C1(n19048), .C2(n19102), .A(n19047), .B(n19046), .ZN(
        P3_U2948) );
  AOI22_X1 U21224 ( .A1(n19062), .A2(n19096), .B1(n19049), .B2(n19103), .ZN(
        n19053) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19051), .B1(
        n19050), .B2(n19108), .ZN(n19052) );
  OAI211_X1 U21226 ( .C1(n19054), .C2(n19102), .A(n19053), .B(n19052), .ZN(
        P3_U2940) );
  AOI22_X1 U21227 ( .A1(n19069), .A2(n19096), .B1(n19055), .B2(n19103), .ZN(
        n19059) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19057), .B1(
        n19056), .B2(n19108), .ZN(n19058) );
  OAI211_X1 U21229 ( .C1(n19060), .C2(n19102), .A(n19059), .B(n19058), .ZN(
        P3_U2932) );
  AOI22_X1 U21230 ( .A1(n19073), .A2(n19096), .B1(n19061), .B2(n19103), .ZN(
        n19065) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19063), .B1(
        n19062), .B2(n19108), .ZN(n19064) );
  OAI211_X1 U21232 ( .C1(n19066), .C2(n19102), .A(n19065), .B(n19064), .ZN(
        P3_U2924) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19068), .B1(
        n19067), .B2(n19103), .ZN(n19071) );
  AOI22_X1 U21234 ( .A1(n19069), .A2(n19108), .B1(n19079), .B2(n19096), .ZN(
        n19070) );
  OAI211_X1 U21235 ( .C1(n19077), .C2(n19102), .A(n19071), .B(n19070), .ZN(
        P3_U2916) );
  AOI22_X1 U21236 ( .A1(n19091), .A2(n19105), .B1(n19072), .B2(n19103), .ZN(
        n19076) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19074), .B1(
        n19073), .B2(n19108), .ZN(n19075) );
  OAI211_X1 U21238 ( .C1(n19077), .C2(n19113), .A(n19076), .B(n19075), .ZN(
        P3_U2908) );
  AOI22_X1 U21239 ( .A1(n19091), .A2(n19096), .B1(n19078), .B2(n19103), .ZN(
        n19082) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19080), .B1(
        n19079), .B2(n19108), .ZN(n19081) );
  OAI211_X1 U21241 ( .C1(n19088), .C2(n19102), .A(n19082), .B(n19081), .ZN(
        P3_U2900) );
  AOI22_X1 U21242 ( .A1(n19109), .A2(n19105), .B1(n19083), .B2(n19103), .ZN(
        n19087) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19085), .B1(
        n19084), .B2(n19108), .ZN(n19086) );
  OAI211_X1 U21244 ( .C1(n19088), .C2(n19113), .A(n19087), .B(n19086), .ZN(
        P3_U2892) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n19103), .ZN(n19093) );
  AOI22_X1 U21246 ( .A1(n19091), .A2(n19108), .B1(n19109), .B2(n19096), .ZN(
        n19092) );
  OAI211_X1 U21247 ( .C1(n19094), .C2(n19102), .A(n19093), .B(n19092), .ZN(
        P3_U2884) );
  AOI22_X1 U21248 ( .A1(n19097), .A2(n19096), .B1(n19095), .B2(n19103), .ZN(
        n19101) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19099), .B1(
        n19098), .B2(n19108), .ZN(n19100) );
  OAI211_X1 U21250 ( .C1(n19114), .C2(n19102), .A(n19101), .B(n19100), .ZN(
        P3_U2876) );
  AOI22_X1 U21251 ( .A1(n10969), .A2(n19105), .B1(n19104), .B2(n19103), .ZN(
        n19112) );
  INV_X1 U21252 ( .A(n19107), .ZN(n19110) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19110), .B1(
        n19109), .B2(n19108), .ZN(n19111) );
  OAI211_X1 U21254 ( .C1(n19114), .C2(n19113), .A(n19112), .B(n19111), .ZN(
        P3_U2868) );
  AOI22_X1 U21255 ( .A1(n19616), .A2(BUF1_REG_31__SCAN_IN), .B1(n19619), .B2(
        n19115), .ZN(n19117) );
  AOI22_X1 U21256 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19613), .B1(n19617), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19116) );
  NAND2_X1 U21257 ( .A1(n19117), .A2(n19116), .ZN(P2_U2888) );
  INV_X1 U21258 ( .A(n19118), .ZN(n19121) );
  AOI22_X1 U21259 ( .A1(n19397), .A2(n19119), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19613), .ZN(n19120) );
  OAI21_X1 U21260 ( .B1(n19404), .B2(n19121), .A(n19120), .ZN(P2_U2905) );
  AOI22_X1 U21261 ( .A1(n19397), .A2(n19122), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19613), .ZN(n19123) );
  OAI21_X1 U21262 ( .B1(n19404), .B2(n19124), .A(n19123), .ZN(P2_U2907) );
  AOI22_X1 U21263 ( .A1(n19397), .A2(n19125), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19613), .ZN(n19126) );
  OAI21_X1 U21264 ( .B1(n19404), .B2(n19127), .A(n19126), .ZN(P2_U2909) );
  AOI22_X1 U21265 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19631), .ZN(n19319) );
  NAND2_X1 U21266 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19149), .ZN(
        n19130) );
  INV_X1 U21267 ( .A(n19135), .ZN(n19128) );
  INV_X1 U21268 ( .A(n19134), .ZN(n19629) );
  OAI21_X1 U21269 ( .B1(n19128), .B2(n19629), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19129) );
  OAI21_X1 U21270 ( .B1(n19130), .B2(n19307), .A(n19129), .ZN(n19630) );
  NOR2_X2 U21271 ( .A1(n19131), .A2(n19625), .ZN(n19340) );
  INV_X1 U21272 ( .A(n12425), .ZN(n19132) );
  NOR2_X2 U21273 ( .A1(n19132), .A2(n19627), .ZN(n19331) );
  AOI22_X1 U21274 ( .A1(n19630), .A2(n19340), .B1(n19629), .B2(n19331), .ZN(
        n19139) );
  INV_X1 U21275 ( .A(n19149), .ZN(n19143) );
  OAI22_X1 U21276 ( .A1(n19153), .A2(n19133), .B1(n19302), .B2(n19143), .ZN(
        n19137) );
  OAI211_X1 U21277 ( .C1(n19135), .C2(n19262), .A(n19307), .B(n19134), .ZN(
        n19136) );
  NAND3_X1 U21278 ( .A1(n19137), .A2(n19313), .A3(n19136), .ZN(n19633) );
  AOI22_X1 U21279 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19631), .ZN(n19301) );
  INV_X1 U21280 ( .A(n19301), .ZN(n19332) );
  NOR2_X2 U21281 ( .A1(n19153), .A2(n19282), .ZN(n19639) );
  AOI22_X1 U21282 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19633), .B1(
        n19332), .B2(n19639), .ZN(n19138) );
  OAI211_X1 U21283 ( .C1(n19319), .C2(n19636), .A(n19139), .B(n19138), .ZN(
        P2_U3175) );
  NOR2_X1 U21284 ( .A1(n19143), .A2(n19288), .ZN(n19637) );
  OAI21_X1 U21285 ( .B1(n13646), .B2(n19637), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19141) );
  OAI21_X1 U21286 ( .B1(n19143), .B2(n19142), .A(n19141), .ZN(n19638) );
  AOI22_X1 U21287 ( .A1(n19638), .A2(n19340), .B1(n19331), .B2(n19637), .ZN(
        n19148) );
  NOR2_X1 U21288 ( .A1(n19143), .A2(n19305), .ZN(n19643) );
  INV_X1 U21289 ( .A(n19643), .ZN(n19154) );
  OAI21_X1 U21290 ( .B1(n19153), .B2(n19292), .A(n19154), .ZN(n19146) );
  OAI21_X1 U21291 ( .B1(n19144), .B2(n19262), .A(n19325), .ZN(n19145) );
  AOI22_X1 U21292 ( .A1(n19146), .A2(n19145), .B1(n19637), .B2(n19313), .ZN(
        n19640) );
  AOI22_X1 U21293 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19339), .ZN(n19147) );
  OAI211_X1 U21294 ( .C1(n19301), .C2(n19648), .A(n19148), .B(n19147), .ZN(
        P2_U3167) );
  NAND2_X1 U21295 ( .A1(n19149), .A2(n19302), .ZN(n19164) );
  INV_X1 U21296 ( .A(n19155), .ZN(n19150) );
  OAI21_X1 U21297 ( .B1(n19150), .B2(n19643), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19151) );
  OAI21_X1 U21298 ( .B1(n19164), .B2(n19307), .A(n19151), .ZN(n19644) );
  AOI22_X1 U21299 ( .A1(n19644), .A2(n19340), .B1(n19331), .B2(n19643), .ZN(
        n19159) );
  NOR2_X2 U21300 ( .A1(n19153), .A2(n19316), .ZN(n19651) );
  AND2_X1 U21301 ( .A1(n19152), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19241) );
  INV_X1 U21302 ( .A(n19241), .ZN(n19308) );
  OAI21_X1 U21303 ( .B1(n19153), .B2(n19308), .A(n19164), .ZN(n19157) );
  OAI211_X1 U21304 ( .C1(n19155), .C2(n19262), .A(n19154), .B(n19307), .ZN(
        n19156) );
  NAND3_X1 U21305 ( .A1(n19157), .A2(n19313), .A3(n19156), .ZN(n19645) );
  AOI22_X1 U21306 ( .A1(n19651), .A2(n19332), .B1(n19645), .B2(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19158) );
  OAI211_X1 U21307 ( .C1(n19319), .C2(n19648), .A(n19159), .B(n19158), .ZN(
        P2_U3159) );
  INV_X1 U21308 ( .A(n19161), .ZN(n19167) );
  NAND2_X1 U21309 ( .A1(n19163), .A2(n19162), .ZN(n19260) );
  INV_X1 U21310 ( .A(n19170), .ZN(n19165) );
  NOR2_X1 U21311 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19164), .ZN(
        n19649) );
  OAI21_X1 U21312 ( .B1(n19165), .B2(n19649), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19166) );
  OAI21_X1 U21313 ( .B1(n19167), .B2(n19260), .A(n19166), .ZN(n19650) );
  AOI22_X1 U21314 ( .A1(n19650), .A2(n19340), .B1(n19331), .B2(n19649), .ZN(
        n19174) );
  INV_X1 U21315 ( .A(n19660), .ZN(n19362) );
  OAI21_X1 U21316 ( .B1(n19651), .B2(n19362), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19168) );
  OAI21_X1 U21317 ( .B1(n19260), .B2(n19175), .A(n19168), .ZN(n19172) );
  INV_X1 U21318 ( .A(n19649), .ZN(n19169) );
  OAI211_X1 U21319 ( .C1(n19170), .C2(n19262), .A(n19169), .B(n19307), .ZN(
        n19171) );
  NAND3_X1 U21320 ( .A1(n19172), .A2(n19171), .A3(n19313), .ZN(n19652) );
  AOI22_X1 U21321 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19651), .B2(n19339), .ZN(n19173) );
  OAI211_X1 U21322 ( .C1(n19301), .C2(n19660), .A(n19174), .B(n19173), .ZN(
        P2_U3151) );
  NOR2_X1 U21323 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19175), .ZN(
        n19200) );
  NAND2_X1 U21324 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19200), .ZN(
        n19177) );
  INV_X1 U21325 ( .A(n19200), .ZN(n19186) );
  NOR2_X1 U21326 ( .A1(n19272), .A2(n19186), .ZN(n19655) );
  OAI21_X1 U21327 ( .B1(n19178), .B2(n19655), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19176) );
  OAI21_X1 U21328 ( .B1(n19177), .B2(n19307), .A(n19176), .ZN(n19656) );
  AOI22_X1 U21329 ( .A1(n19656), .A2(n19340), .B1(n19331), .B2(n19655), .ZN(
        n19185) );
  INV_X1 U21330 ( .A(n19325), .ZN(n19182) );
  AOI21_X1 U21331 ( .B1(n19178), .B2(n19329), .A(n19655), .ZN(n19179) );
  INV_X1 U21332 ( .A(n19179), .ZN(n19181) );
  OAI22_X1 U21333 ( .A1(n19255), .A2(n19273), .B1(n19302), .B2(n19186), .ZN(
        n19180) );
  OAI211_X1 U21334 ( .C1(n19182), .C2(n19181), .A(n19180), .B(n19313), .ZN(
        n19657) );
  INV_X1 U21335 ( .A(n19206), .ZN(n19183) );
  NOR2_X2 U21336 ( .A1(n19183), .A2(n19282), .ZN(n19662) );
  AOI22_X1 U21337 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19332), .ZN(n19184) );
  OAI211_X1 U21338 ( .C1(n19319), .C2(n19660), .A(n19185), .B(n19184), .ZN(
        P2_U3143) );
  NOR2_X1 U21339 ( .A1(n19288), .A2(n19186), .ZN(n19661) );
  AOI22_X1 U21340 ( .A1(n19339), .A2(n19662), .B1(n19331), .B2(n19661), .ZN(
        n19198) );
  NOR2_X1 U21341 ( .A1(n19305), .A2(n19186), .ZN(n19667) );
  NOR2_X1 U21342 ( .A1(n19661), .A2(n19667), .ZN(n19196) );
  INV_X1 U21343 ( .A(n19196), .ZN(n19191) );
  OAI21_X1 U21344 ( .B1(n19188), .B2(n19187), .A(n19321), .ZN(n19195) );
  INV_X1 U21345 ( .A(n19661), .ZN(n19189) );
  OAI211_X1 U21346 ( .C1(n19192), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19189), 
        .B(n19325), .ZN(n19190) );
  OAI211_X1 U21347 ( .C1(n19191), .C2(n19195), .A(n19190), .B(n19313), .ZN(
        n19664) );
  INV_X1 U21348 ( .A(n19192), .ZN(n19193) );
  OAI21_X1 U21349 ( .B1(n19193), .B2(n19661), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19194) );
  OAI21_X1 U21350 ( .B1(n19196), .B2(n19195), .A(n19194), .ZN(n19663) );
  AOI22_X1 U21351 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19664), .B1(
        n19340), .B2(n19663), .ZN(n19197) );
  OAI211_X1 U21352 ( .C1(n19301), .C2(n19672), .A(n19198), .B(n19197), .ZN(
        P2_U3135) );
  NAND2_X1 U21353 ( .A1(n19206), .A2(n19241), .ZN(n19199) );
  NAND2_X1 U21354 ( .A1(n19199), .A2(n19321), .ZN(n19208) );
  NAND2_X1 U21355 ( .A1(n19200), .A2(n19302), .ZN(n19212) );
  INV_X1 U21356 ( .A(n19212), .ZN(n19201) );
  OR2_X1 U21357 ( .A1(n19208), .A2(n19201), .ZN(n19205) );
  INV_X1 U21358 ( .A(n19667), .ZN(n19203) );
  NAND2_X1 U21359 ( .A1(n13699), .A2(n19329), .ZN(n19202) );
  OAI211_X1 U21360 ( .C1(n19625), .C2(n19203), .A(n19202), .B(n19325), .ZN(
        n19204) );
  INV_X1 U21361 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n19211) );
  INV_X1 U21362 ( .A(n19316), .ZN(n19239) );
  AOI22_X1 U21363 ( .A1(n19332), .A2(n19674), .B1(n19667), .B2(n19331), .ZN(
        n19210) );
  OAI21_X1 U21364 ( .B1(n13699), .B2(n19667), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19207) );
  OAI21_X1 U21365 ( .B1(n19208), .B2(n19212), .A(n19207), .ZN(n19668) );
  AOI22_X1 U21366 ( .A1(n19340), .A2(n19668), .B1(n19462), .B2(n19339), .ZN(
        n19209) );
  OAI211_X1 U21367 ( .C1(n19367), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P2_U3127) );
  NOR2_X1 U21368 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19212), .ZN(
        n19673) );
  AOI22_X1 U21369 ( .A1(n19339), .A2(n19674), .B1(n19673), .B2(n19331), .ZN(
        n19226) );
  NAND2_X1 U21370 ( .A1(n19321), .A2(n19684), .ZN(n19213) );
  NAND2_X1 U21371 ( .A1(n19321), .A2(n21698), .ZN(n19322) );
  NOR2_X1 U21372 ( .A1(n19272), .A2(n19240), .ZN(n19679) );
  NOR2_X1 U21373 ( .A1(n19679), .A2(n19673), .ZN(n19222) );
  INV_X1 U21374 ( .A(n19222), .ZN(n19216) );
  INV_X1 U21375 ( .A(n19673), .ZN(n19217) );
  OAI211_X1 U21376 ( .C1(n19218), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19217), 
        .B(n19307), .ZN(n19215) );
  NAND2_X1 U21377 ( .A1(n19218), .A2(n19217), .ZN(n19219) );
  NAND2_X1 U21378 ( .A1(n19219), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19220) );
  NAND2_X1 U21379 ( .A1(n19221), .A2(n19220), .ZN(n19224) );
  NAND2_X1 U21380 ( .A1(n19335), .A2(n19222), .ZN(n19223) );
  AOI22_X1 U21381 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19340), .ZN(n19225) );
  OAI211_X1 U21382 ( .C1(n19301), .C2(n19684), .A(n19226), .B(n19225), .ZN(
        P2_U3119) );
  NAND2_X1 U21383 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19243), .ZN(
        n19229) );
  INV_X1 U21384 ( .A(n19231), .ZN(n19227) );
  OAI21_X1 U21385 ( .B1(n19227), .B2(n19679), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19228) );
  OAI21_X1 U21386 ( .B1(n19229), .B2(n19307), .A(n19228), .ZN(n19680) );
  AOI22_X1 U21387 ( .A1(n19680), .A2(n19340), .B1(n19679), .B2(n19331), .ZN(
        n19236) );
  INV_X1 U21388 ( .A(n19229), .ZN(n19233) );
  INV_X1 U21389 ( .A(n19679), .ZN(n19230) );
  OAI211_X1 U21390 ( .C1(n19231), .C2(n19262), .A(n19307), .B(n19230), .ZN(
        n19232) );
  OAI211_X1 U21391 ( .C1(n19234), .C2(n19233), .A(n19313), .B(n19232), .ZN(
        n19681) );
  AOI22_X1 U21392 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n19332), .B2(n19688), .ZN(n19235) );
  OAI211_X1 U21393 ( .C1(n19319), .C2(n19684), .A(n19236), .B(n19235), .ZN(
        P2_U3111) );
  AOI22_X1 U21394 ( .A1(n19686), .A2(n19340), .B1(n19331), .B2(n19685), .ZN(
        n19238) );
  AOI22_X1 U21395 ( .A1(n19339), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19237) );
  OAI211_X1 U21396 ( .C1(n19301), .C2(n19696), .A(n19238), .B(n19237), .ZN(
        P2_U3103) );
  NOR2_X1 U21397 ( .A1(n19305), .A2(n19240), .ZN(n19691) );
  AOI22_X1 U21398 ( .A1(n19332), .A2(n19698), .B1(n19691), .B2(n19331), .ZN(
        n19253) );
  AOI21_X1 U21399 ( .B1(n19242), .B2(n19241), .A(n19307), .ZN(n19249) );
  INV_X1 U21400 ( .A(n19249), .ZN(n19246) );
  NAND2_X1 U21401 ( .A1(n19243), .A2(n19302), .ZN(n19257) );
  INV_X1 U21402 ( .A(n19248), .ZN(n19244) );
  OAI21_X1 U21403 ( .B1(n19244), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19245) );
  INV_X1 U21404 ( .A(n19691), .ZN(n19247) );
  OAI211_X1 U21405 ( .C1(n19248), .C2(n19262), .A(n19307), .B(n19247), .ZN(
        n19251) );
  NAND2_X1 U21406 ( .A1(n19249), .A2(n19257), .ZN(n19250) );
  NAND3_X1 U21407 ( .A1(n19251), .A2(n19313), .A3(n19250), .ZN(n19692) );
  AOI22_X1 U21408 ( .A1(n19693), .A2(n19340), .B1(
        P2_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n19692), .ZN(n19252) );
  OAI211_X1 U21409 ( .C1(n19319), .C2(n19696), .A(n19253), .B(n19252), .ZN(
        P2_U3095) );
  NOR2_X1 U21410 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19257), .ZN(
        n19697) );
  AOI22_X1 U21411 ( .A1(n19339), .A2(n19698), .B1(n19697), .B2(n19331), .ZN(
        n19271) );
  NOR3_X1 U21412 ( .A1(n19705), .A2(n19698), .A3(n19307), .ZN(n19259) );
  INV_X1 U21413 ( .A(n19322), .ZN(n19258) );
  NOR2_X1 U21414 ( .A1(n19259), .A2(n19258), .ZN(n19269) );
  OR2_X1 U21415 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19260), .ZN(
        n19268) );
  INV_X1 U21416 ( .A(n19268), .ZN(n19265) );
  INV_X1 U21417 ( .A(n19697), .ZN(n19261) );
  OAI211_X1 U21418 ( .C1(n19263), .C2(n19262), .A(n19261), .B(n19325), .ZN(
        n19264) );
  OAI211_X1 U21419 ( .C1(n19269), .C2(n19265), .A(n19313), .B(n19264), .ZN(
        n19700) );
  OAI21_X1 U21420 ( .B1(n19266), .B2(n19697), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19267) );
  AOI22_X1 U21421 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19700), .B1(
        n19340), .B2(n19699), .ZN(n19270) );
  OAI211_X1 U21422 ( .C1(n19301), .C2(n19703), .A(n19271), .B(n19270), .ZN(
        P2_U3087) );
  NAND2_X1 U21423 ( .A1(n13698), .A2(n19329), .ZN(n19278) );
  NOR2_X1 U21424 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19303) );
  INV_X1 U21425 ( .A(n19303), .ZN(n19304) );
  NOR2_X1 U21426 ( .A1(n19272), .A2(n19304), .ZN(n19704) );
  OAI21_X1 U21427 ( .B1(n19321), .B2(n19704), .A(n19313), .ZN(n19277) );
  NOR2_X1 U21428 ( .A1(n19274), .A2(n19273), .ZN(n19275) );
  AND2_X1 U21429 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19303), .ZN(
        n19279) );
  NOR2_X1 U21430 ( .A1(n19275), .A2(n19279), .ZN(n19276) );
  INV_X1 U21431 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n19285) );
  AOI22_X1 U21432 ( .A1(n19339), .A2(n19705), .B1(n19704), .B2(n19331), .ZN(
        n19284) );
  OAI21_X1 U21433 ( .B1(n13698), .B2(n19704), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19281) );
  NAND2_X1 U21434 ( .A1(n19321), .A2(n19279), .ZN(n19280) );
  NAND2_X1 U21435 ( .A1(n19281), .A2(n19280), .ZN(n19706) );
  NOR2_X2 U21436 ( .A1(n19315), .A2(n19282), .ZN(n19713) );
  AOI22_X1 U21437 ( .A1(n19340), .A2(n19706), .B1(n19713), .B2(n19332), .ZN(
        n19283) );
  OAI211_X1 U21438 ( .C1(n19710), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        P2_U3079) );
  NOR2_X1 U21439 ( .A1(n19288), .A2(n19304), .ZN(n19711) );
  OAI21_X1 U21440 ( .B1(n19294), .B2(n19711), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19290) );
  NAND2_X1 U21441 ( .A1(n19289), .A2(n19303), .ZN(n19291) );
  NAND2_X1 U21442 ( .A1(n19290), .A2(n19291), .ZN(n19712) );
  AOI22_X1 U21443 ( .A1(n19712), .A2(n19340), .B1(n19331), .B2(n19711), .ZN(
        n19300) );
  OAI211_X1 U21444 ( .C1(n19315), .C2(n19292), .A(n19321), .B(n19291), .ZN(
        n19298) );
  OAI21_X1 U21445 ( .B1(n19294), .B2(n19335), .A(n19293), .ZN(n19296) );
  INV_X1 U21446 ( .A(n19711), .ZN(n19295) );
  AOI21_X1 U21447 ( .B1(n19296), .B2(n19295), .A(n19327), .ZN(n19297) );
  NAND2_X1 U21448 ( .A1(n19298), .A2(n19297), .ZN(n19714) );
  AOI22_X1 U21449 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19339), .ZN(n19299) );
  OAI211_X1 U21450 ( .C1(n19301), .C2(n19723), .A(n19300), .B(n19299), .ZN(
        P2_U3071) );
  NAND2_X1 U21451 ( .A1(n19303), .A2(n19302), .ZN(n19324) );
  NOR2_X1 U21452 ( .A1(n19305), .A2(n19304), .ZN(n19718) );
  OAI21_X1 U21453 ( .B1(n19309), .B2(n19718), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19306) );
  OAI21_X1 U21454 ( .B1(n19324), .B2(n19307), .A(n19306), .ZN(n19719) );
  AOI22_X1 U21455 ( .A1(n19719), .A2(n19340), .B1(n19331), .B2(n19718), .ZN(
        n19318) );
  OAI21_X1 U21456 ( .B1(n19315), .B2(n19308), .A(n19324), .ZN(n19314) );
  NAND2_X1 U21457 ( .A1(n19309), .A2(n19329), .ZN(n19311) );
  INV_X1 U21458 ( .A(n19718), .ZN(n19310) );
  NAND3_X1 U21459 ( .A1(n19311), .A2(n19325), .A3(n19310), .ZN(n19312) );
  NAND3_X1 U21460 ( .A1(n19314), .A2(n19313), .A3(n19312), .ZN(n19720) );
  AOI22_X1 U21461 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19332), .ZN(n19317) );
  OAI211_X1 U21462 ( .C1(n19319), .C2(n19723), .A(n19318), .B(n19317), .ZN(
        P2_U3063) );
  INV_X1 U21463 ( .A(n19732), .ZN(n19320) );
  NAND2_X1 U21464 ( .A1(n19321), .A2(n19320), .ZN(n19323) );
  OAI21_X1 U21465 ( .B1(n19727), .B2(n19323), .A(n19322), .ZN(n19333) );
  NOR2_X1 U21466 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19324), .ZN(
        n19726) );
  NOR2_X1 U21467 ( .A1(n19629), .A2(n19726), .ZN(n19336) );
  INV_X1 U21468 ( .A(n19726), .ZN(n19326) );
  OAI21_X1 U21469 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19328) );
  AOI21_X1 U21470 ( .B1(n19334), .B2(n19329), .A(n19328), .ZN(n19330) );
  AOI22_X1 U21471 ( .A1(n19332), .A2(n19727), .B1(n19726), .B2(n19331), .ZN(
        n19342) );
  INV_X1 U21472 ( .A(n19333), .ZN(n19338) );
  OAI21_X1 U21473 ( .B1(n19334), .B2(n19726), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19337) );
  AOI22_X1 U21474 ( .A1(n19340), .A2(n19730), .B1(n19732), .B2(n19339), .ZN(
        n19341) );
  OAI211_X1 U21475 ( .C1(n19735), .C2(n19343), .A(n19342), .B(n19341), .ZN(
        P2_U3055) );
  AOI22_X1 U21476 ( .A1(n19615), .A2(n19344), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19613), .ZN(n19351) );
  AOI22_X1 U21477 ( .A1(n19617), .A2(BUF2_REG_22__SCAN_IN), .B1(n19616), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19350) );
  INV_X1 U21478 ( .A(n19345), .ZN(n19348) );
  INV_X1 U21479 ( .A(n19346), .ZN(n19347) );
  AOI22_X1 U21480 ( .A1(n19348), .A2(n19620), .B1(n19619), .B2(n19347), .ZN(
        n19349) );
  NAND3_X1 U21481 ( .A1(n19351), .A2(n19350), .A3(n19349), .ZN(P2_U2897) );
  AOI22_X1 U21482 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19631), .ZN(n19388) );
  NOR2_X2 U21483 ( .A1(n19352), .A2(n19625), .ZN(n19391) );
  NOR2_X2 U21484 ( .A1(n19353), .A2(n19627), .ZN(n19389) );
  AOI22_X1 U21485 ( .A1(n19630), .A2(n19391), .B1(n19629), .B2(n19389), .ZN(
        n19355) );
  AOI22_X1 U21486 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19632), .ZN(n19385) );
  INV_X1 U21487 ( .A(n19385), .ZN(n19390) );
  AOI22_X1 U21488 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19633), .B1(
        n19390), .B2(n19639), .ZN(n19354) );
  OAI211_X1 U21489 ( .C1(n19388), .C2(n19636), .A(n19355), .B(n19354), .ZN(
        P2_U3174) );
  AOI22_X1 U21490 ( .A1(n19638), .A2(n19391), .B1(n19389), .B2(n19637), .ZN(
        n19357) );
  INV_X1 U21491 ( .A(n19388), .ZN(n19392) );
  AOI22_X1 U21492 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19392), .ZN(n19356) );
  OAI211_X1 U21493 ( .C1(n19385), .C2(n19648), .A(n19357), .B(n19356), .ZN(
        P2_U3166) );
  AOI22_X1 U21494 ( .A1(n19644), .A2(n19391), .B1(n19389), .B2(n19643), .ZN(
        n19359) );
  AOI22_X1 U21495 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19645), .B1(
        n19390), .B2(n19651), .ZN(n19358) );
  OAI211_X1 U21496 ( .C1(n19388), .C2(n19648), .A(n19359), .B(n19358), .ZN(
        P2_U3158) );
  AOI22_X1 U21497 ( .A1(n19650), .A2(n19391), .B1(n19389), .B2(n19649), .ZN(
        n19361) );
  AOI22_X1 U21498 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n19651), .B2(n19392), .ZN(n19360) );
  OAI211_X1 U21499 ( .C1(n19385), .C2(n19660), .A(n19361), .B(n19360), .ZN(
        P2_U3150) );
  INV_X1 U21500 ( .A(n19662), .ZN(n19465) );
  AOI22_X1 U21501 ( .A1(n19656), .A2(n19391), .B1(n19389), .B2(n19655), .ZN(
        n19364) );
  AOI22_X1 U21502 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19657), .B1(
        n19362), .B2(n19392), .ZN(n19363) );
  OAI211_X1 U21503 ( .C1(n19385), .C2(n19465), .A(n19364), .B(n19363), .ZN(
        P2_U3142) );
  AOI22_X1 U21504 ( .A1(n19390), .A2(n19462), .B1(n19389), .B2(n19661), .ZN(
        n19366) );
  AOI22_X1 U21505 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19664), .B1(
        n19391), .B2(n19663), .ZN(n19365) );
  OAI211_X1 U21506 ( .C1(n19388), .C2(n19465), .A(n19366), .B(n19365), .ZN(
        P2_U3134) );
  AOI22_X1 U21507 ( .A1(n19390), .A2(n19674), .B1(n19667), .B2(n19389), .ZN(
        n19369) );
  AOI22_X1 U21508 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19669), .B1(
        n19391), .B2(n19668), .ZN(n19368) );
  OAI211_X1 U21509 ( .C1(n19388), .C2(n19672), .A(n19369), .B(n19368), .ZN(
        P2_U3126) );
  AOI22_X1 U21510 ( .A1(n19392), .A2(n19674), .B1(n19673), .B2(n19389), .ZN(
        n19371) );
  AOI22_X1 U21511 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19391), .ZN(n19370) );
  OAI211_X1 U21512 ( .C1(n19385), .C2(n19684), .A(n19371), .B(n19370), .ZN(
        P2_U3118) );
  AOI22_X1 U21513 ( .A1(n19680), .A2(n19391), .B1(n19679), .B2(n19389), .ZN(
        n19373) );
  AOI22_X1 U21514 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n19390), .B2(n19688), .ZN(n19372) );
  OAI211_X1 U21515 ( .C1(n19388), .C2(n19684), .A(n19373), .B(n19372), .ZN(
        P2_U3110) );
  AOI22_X1 U21516 ( .A1(n19686), .A2(n19391), .B1(n19389), .B2(n19685), .ZN(
        n19375) );
  AOI22_X1 U21517 ( .A1(n19392), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n19374) );
  OAI211_X1 U21518 ( .C1(n19385), .C2(n19696), .A(n19375), .B(n19374), .ZN(
        P2_U3102) );
  AOI22_X1 U21519 ( .A1(n19390), .A2(n19698), .B1(n19691), .B2(n19389), .ZN(
        n19377) );
  AOI22_X1 U21520 ( .A1(n19693), .A2(n19391), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n19692), .ZN(n19376) );
  OAI211_X1 U21521 ( .C1(n19388), .C2(n19696), .A(n19377), .B(n19376), .ZN(
        P2_U3094) );
  AOI22_X1 U21522 ( .A1(n19392), .A2(n19698), .B1(n19697), .B2(n19389), .ZN(
        n19379) );
  AOI22_X1 U21523 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19700), .B1(
        n19391), .B2(n19699), .ZN(n19378) );
  OAI211_X1 U21524 ( .C1(n19385), .C2(n19703), .A(n19379), .B(n19378), .ZN(
        P2_U3086) );
  INV_X1 U21525 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n19382) );
  AOI22_X1 U21526 ( .A1(n19392), .A2(n19705), .B1(n19704), .B2(n19389), .ZN(
        n19381) );
  AOI22_X1 U21527 ( .A1(n19391), .A2(n19706), .B1(n19713), .B2(n19390), .ZN(
        n19380) );
  OAI211_X1 U21528 ( .C1(n19710), .C2(n19382), .A(n19381), .B(n19380), .ZN(
        P2_U3078) );
  AOI22_X1 U21529 ( .A1(n19712), .A2(n19391), .B1(n19389), .B2(n19711), .ZN(
        n19384) );
  AOI22_X1 U21530 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19392), .ZN(n19383) );
  OAI211_X1 U21531 ( .C1(n19385), .C2(n19723), .A(n19384), .B(n19383), .ZN(
        P2_U3070) );
  AOI22_X1 U21532 ( .A1(n19719), .A2(n19391), .B1(n19389), .B2(n19718), .ZN(
        n19387) );
  AOI22_X1 U21533 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19390), .ZN(n19386) );
  OAI211_X1 U21534 ( .C1(n19388), .C2(n19723), .A(n19387), .B(n19386), .ZN(
        P2_U3062) );
  AOI22_X1 U21535 ( .A1(n19390), .A2(n19727), .B1(n19726), .B2(n19389), .ZN(
        n19394) );
  AOI22_X1 U21536 ( .A1(n19732), .A2(n19392), .B1(n19730), .B2(n19391), .ZN(
        n19393) );
  OAI211_X1 U21537 ( .C1(n19735), .C2(n19395), .A(n19394), .B(n19393), .ZN(
        P2_U3054) );
  INV_X1 U21538 ( .A(n19405), .ZN(n19396) );
  AOI22_X1 U21539 ( .A1(n19397), .A2(n19396), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19613), .ZN(n19402) );
  OR3_X1 U21540 ( .A1(n19400), .A2(n19399), .A3(n19398), .ZN(n19401) );
  OAI211_X1 U21541 ( .C1(n19404), .C2(n19403), .A(n19402), .B(n19401), .ZN(
        P2_U2914) );
  AOI22_X1 U21542 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19631), .ZN(n19438) );
  NOR2_X2 U21543 ( .A1(n19405), .A2(n19625), .ZN(n19441) );
  NOR2_X2 U21544 ( .A1(n13989), .A2(n19627), .ZN(n19439) );
  AOI22_X1 U21545 ( .A1(n19630), .A2(n19441), .B1(n19629), .B2(n19439), .ZN(
        n19407) );
  AOI22_X1 U21546 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19632), .ZN(n19435) );
  AOI22_X1 U21547 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19633), .B1(
        n19440), .B2(n19639), .ZN(n19406) );
  OAI211_X1 U21548 ( .C1(n19438), .C2(n19636), .A(n19407), .B(n19406), .ZN(
        P2_U3173) );
  AOI22_X1 U21549 ( .A1(n19638), .A2(n19441), .B1(n19439), .B2(n19637), .ZN(
        n19409) );
  INV_X1 U21550 ( .A(n19438), .ZN(n19442) );
  AOI22_X1 U21551 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19442), .ZN(n19408) );
  OAI211_X1 U21552 ( .C1(n19435), .C2(n19648), .A(n19409), .B(n19408), .ZN(
        P2_U3165) );
  AOI22_X1 U21553 ( .A1(n19644), .A2(n19441), .B1(n19439), .B2(n19643), .ZN(
        n19411) );
  AOI22_X1 U21554 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19645), .B1(
        n19440), .B2(n19651), .ZN(n19410) );
  OAI211_X1 U21555 ( .C1(n19438), .C2(n19648), .A(n19411), .B(n19410), .ZN(
        P2_U3157) );
  AOI22_X1 U21556 ( .A1(n19650), .A2(n19441), .B1(n19439), .B2(n19649), .ZN(
        n19413) );
  AOI22_X1 U21557 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n19651), .B2(n19442), .ZN(n19412) );
  OAI211_X1 U21558 ( .C1(n19435), .C2(n19660), .A(n19413), .B(n19412), .ZN(
        P2_U3149) );
  AOI22_X1 U21559 ( .A1(n19656), .A2(n19441), .B1(n19439), .B2(n19655), .ZN(
        n19415) );
  AOI22_X1 U21560 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19440), .ZN(n19414) );
  OAI211_X1 U21561 ( .C1(n19438), .C2(n19660), .A(n19415), .B(n19414), .ZN(
        P2_U3141) );
  AOI22_X1 U21562 ( .A1(n19440), .A2(n19462), .B1(n19439), .B2(n19661), .ZN(
        n19417) );
  AOI22_X1 U21563 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19664), .B1(
        n19441), .B2(n19663), .ZN(n19416) );
  OAI211_X1 U21564 ( .C1(n19438), .C2(n19465), .A(n19417), .B(n19416), .ZN(
        P2_U3133) );
  AOI22_X1 U21565 ( .A1(n19440), .A2(n19674), .B1(n19667), .B2(n19439), .ZN(
        n19419) );
  AOI22_X1 U21566 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19669), .B1(
        n19441), .B2(n19668), .ZN(n19418) );
  OAI211_X1 U21567 ( .C1(n19438), .C2(n19672), .A(n19419), .B(n19418), .ZN(
        P2_U3125) );
  AOI22_X1 U21568 ( .A1(n19442), .A2(n19674), .B1(n19439), .B2(n19673), .ZN(
        n19421) );
  AOI22_X1 U21569 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19441), .ZN(n19420) );
  OAI211_X1 U21570 ( .C1(n19435), .C2(n19684), .A(n19421), .B(n19420), .ZN(
        P2_U3117) );
  AOI22_X1 U21571 ( .A1(n19680), .A2(n19441), .B1(n19679), .B2(n19439), .ZN(
        n19423) );
  AOI22_X1 U21572 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n19688), .B2(n19440), .ZN(n19422) );
  OAI211_X1 U21573 ( .C1(n19438), .C2(n19684), .A(n19423), .B(n19422), .ZN(
        P2_U3109) );
  AOI22_X1 U21574 ( .A1(n19686), .A2(n19441), .B1(n19439), .B2(n19685), .ZN(
        n19425) );
  AOI22_X1 U21575 ( .A1(n19442), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n19424) );
  OAI211_X1 U21576 ( .C1(n19435), .C2(n19696), .A(n19425), .B(n19424), .ZN(
        P2_U3101) );
  AOI22_X1 U21577 ( .A1(n19440), .A2(n19698), .B1(n19439), .B2(n19691), .ZN(
        n19427) );
  AOI22_X1 U21578 ( .A1(n19693), .A2(n19441), .B1(
        P2_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n19692), .ZN(n19426) );
  OAI211_X1 U21579 ( .C1(n19438), .C2(n19696), .A(n19427), .B(n19426), .ZN(
        P2_U3093) );
  AOI22_X1 U21580 ( .A1(n19442), .A2(n19698), .B1(n19439), .B2(n19697), .ZN(
        n19429) );
  AOI22_X1 U21581 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19700), .B1(
        n19441), .B2(n19699), .ZN(n19428) );
  OAI211_X1 U21582 ( .C1(n19435), .C2(n19703), .A(n19429), .B(n19428), .ZN(
        P2_U3085) );
  INV_X1 U21583 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n19432) );
  AOI22_X1 U21584 ( .A1(n19442), .A2(n19705), .B1(n19439), .B2(n19704), .ZN(
        n19431) );
  AOI22_X1 U21585 ( .A1(n19441), .A2(n19706), .B1(n19713), .B2(n19440), .ZN(
        n19430) );
  OAI211_X1 U21586 ( .C1(n19710), .C2(n19432), .A(n19431), .B(n19430), .ZN(
        P2_U3077) );
  AOI22_X1 U21587 ( .A1(n19712), .A2(n19441), .B1(n19439), .B2(n19711), .ZN(
        n19434) );
  AOI22_X1 U21588 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19442), .ZN(n19433) );
  OAI211_X1 U21589 ( .C1(n19435), .C2(n19723), .A(n19434), .B(n19433), .ZN(
        P2_U3069) );
  AOI22_X1 U21590 ( .A1(n19719), .A2(n19441), .B1(n19439), .B2(n19718), .ZN(
        n19437) );
  AOI22_X1 U21591 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19440), .ZN(n19436) );
  OAI211_X1 U21592 ( .C1(n19438), .C2(n19723), .A(n19437), .B(n19436), .ZN(
        P2_U3061) );
  AOI22_X1 U21593 ( .A1(n19440), .A2(n19727), .B1(n19726), .B2(n19439), .ZN(
        n19444) );
  AOI22_X1 U21594 ( .A1(n19732), .A2(n19442), .B1(n19730), .B2(n19441), .ZN(
        n19443) );
  OAI211_X1 U21595 ( .C1(n19735), .C2(n14610), .A(n19444), .B(n19443), .ZN(
        P2_U3053) );
  AOI22_X1 U21596 ( .A1(n19615), .A2(n19445), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19613), .ZN(n19450) );
  AOI22_X1 U21597 ( .A1(n19617), .A2(BUF2_REG_20__SCAN_IN), .B1(n19616), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n19449) );
  AOI22_X1 U21598 ( .A1(n19447), .A2(n19620), .B1(n19619), .B2(n19446), .ZN(
        n19448) );
  NAND3_X1 U21599 ( .A1(n19450), .A2(n19449), .A3(n19448), .ZN(P2_U2899) );
  AOI22_X1 U21600 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19631), .ZN(n19486) );
  NOR2_X2 U21601 ( .A1(n19451), .A2(n19625), .ZN(n19489) );
  NOR2_X2 U21602 ( .A1(n12419), .A2(n19627), .ZN(n19487) );
  AOI22_X1 U21603 ( .A1(n19630), .A2(n19489), .B1(n19629), .B2(n19487), .ZN(
        n19453) );
  AOI22_X1 U21604 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19632), .ZN(n19483) );
  AOI22_X1 U21605 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19633), .B1(
        n19488), .B2(n19639), .ZN(n19452) );
  OAI211_X1 U21606 ( .C1(n19486), .C2(n19636), .A(n19453), .B(n19452), .ZN(
        P2_U3172) );
  AOI22_X1 U21607 ( .A1(n19638), .A2(n19489), .B1(n19487), .B2(n19637), .ZN(
        n19455) );
  INV_X1 U21608 ( .A(n19486), .ZN(n19490) );
  AOI22_X1 U21609 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19490), .ZN(n19454) );
  OAI211_X1 U21610 ( .C1(n19483), .C2(n19648), .A(n19455), .B(n19454), .ZN(
        P2_U3164) );
  AOI22_X1 U21611 ( .A1(n19644), .A2(n19489), .B1(n19487), .B2(n19643), .ZN(
        n19457) );
  AOI22_X1 U21612 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19645), .B1(
        n19488), .B2(n19651), .ZN(n19456) );
  OAI211_X1 U21613 ( .C1(n19486), .C2(n19648), .A(n19457), .B(n19456), .ZN(
        P2_U3156) );
  AOI22_X1 U21614 ( .A1(n19650), .A2(n19489), .B1(n19487), .B2(n19649), .ZN(
        n19459) );
  AOI22_X1 U21615 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n19651), .B2(n19490), .ZN(n19458) );
  OAI211_X1 U21616 ( .C1(n19483), .C2(n19660), .A(n19459), .B(n19458), .ZN(
        P2_U3148) );
  AOI22_X1 U21617 ( .A1(n19656), .A2(n19489), .B1(n19487), .B2(n19655), .ZN(
        n19461) );
  AOI22_X1 U21618 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19488), .ZN(n19460) );
  OAI211_X1 U21619 ( .C1(n19486), .C2(n19660), .A(n19461), .B(n19460), .ZN(
        P2_U3140) );
  AOI22_X1 U21620 ( .A1(n19488), .A2(n19462), .B1(n19487), .B2(n19661), .ZN(
        n19464) );
  AOI22_X1 U21621 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19664), .B1(
        n19489), .B2(n19663), .ZN(n19463) );
  OAI211_X1 U21622 ( .C1(n19486), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P2_U3132) );
  AOI22_X1 U21623 ( .A1(n19488), .A2(n19674), .B1(n19667), .B2(n19487), .ZN(
        n19467) );
  AOI22_X1 U21624 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19669), .B1(
        n19489), .B2(n19668), .ZN(n19466) );
  OAI211_X1 U21625 ( .C1(n19486), .C2(n19672), .A(n19467), .B(n19466), .ZN(
        P2_U3124) );
  AOI22_X1 U21626 ( .A1(n19490), .A2(n19674), .B1(n19487), .B2(n19673), .ZN(
        n19469) );
  AOI22_X1 U21627 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19489), .ZN(n19468) );
  OAI211_X1 U21628 ( .C1(n19483), .C2(n19684), .A(n19469), .B(n19468), .ZN(
        P2_U3116) );
  AOI22_X1 U21629 ( .A1(n19680), .A2(n19489), .B1(n19679), .B2(n19487), .ZN(
        n19471) );
  AOI22_X1 U21630 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n19688), .B2(n19488), .ZN(n19470) );
  OAI211_X1 U21631 ( .C1(n19486), .C2(n19684), .A(n19471), .B(n19470), .ZN(
        P2_U3108) );
  AOI22_X1 U21632 ( .A1(n19686), .A2(n19489), .B1(n19487), .B2(n19685), .ZN(
        n19473) );
  AOI22_X1 U21633 ( .A1(n19490), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n19472) );
  OAI211_X1 U21634 ( .C1(n19483), .C2(n19696), .A(n19473), .B(n19472), .ZN(
        P2_U3100) );
  AOI22_X1 U21635 ( .A1(n19488), .A2(n19698), .B1(n19487), .B2(n19691), .ZN(
        n19475) );
  AOI22_X1 U21636 ( .A1(n19693), .A2(n19489), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n19692), .ZN(n19474) );
  OAI211_X1 U21637 ( .C1(n19486), .C2(n19696), .A(n19475), .B(n19474), .ZN(
        P2_U3092) );
  AOI22_X1 U21638 ( .A1(n19490), .A2(n19698), .B1(n19697), .B2(n19487), .ZN(
        n19477) );
  AOI22_X1 U21639 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19700), .B1(
        n19489), .B2(n19699), .ZN(n19476) );
  OAI211_X1 U21640 ( .C1(n19483), .C2(n19703), .A(n19477), .B(n19476), .ZN(
        P2_U3084) );
  INV_X1 U21641 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n19480) );
  AOI22_X1 U21642 ( .A1(n19490), .A2(n19705), .B1(n19487), .B2(n19704), .ZN(
        n19479) );
  AOI22_X1 U21643 ( .A1(n19489), .A2(n19706), .B1(n19713), .B2(n19488), .ZN(
        n19478) );
  OAI211_X1 U21644 ( .C1(n19710), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P2_U3076) );
  AOI22_X1 U21645 ( .A1(n19712), .A2(n19489), .B1(n19487), .B2(n19711), .ZN(
        n19482) );
  AOI22_X1 U21646 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19490), .ZN(n19481) );
  OAI211_X1 U21647 ( .C1(n19483), .C2(n19723), .A(n19482), .B(n19481), .ZN(
        P2_U3068) );
  AOI22_X1 U21648 ( .A1(n19719), .A2(n19489), .B1(n19487), .B2(n19718), .ZN(
        n19485) );
  AOI22_X1 U21649 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19488), .ZN(n19484) );
  OAI211_X1 U21650 ( .C1(n19486), .C2(n19723), .A(n19485), .B(n19484), .ZN(
        P2_U3060) );
  AOI22_X1 U21651 ( .A1(n19488), .A2(n19727), .B1(n19726), .B2(n19487), .ZN(
        n19492) );
  AOI22_X1 U21652 ( .A1(n19732), .A2(n19490), .B1(n19730), .B2(n19489), .ZN(
        n19491) );
  OAI211_X1 U21653 ( .C1(n19735), .C2(n19493), .A(n19492), .B(n19491), .ZN(
        P2_U3052) );
  AOI22_X1 U21654 ( .A1(n19630), .A2(n19527), .B1(n19629), .B2(n19525), .ZN(
        n19495) );
  INV_X1 U21655 ( .A(n19521), .ZN(n19526) );
  AOI22_X1 U21656 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19633), .B1(
        n19526), .B2(n19639), .ZN(n19494) );
  OAI211_X1 U21657 ( .C1(n19524), .C2(n19636), .A(n19495), .B(n19494), .ZN(
        P2_U3171) );
  AOI22_X1 U21658 ( .A1(n19638), .A2(n19527), .B1(n19525), .B2(n19637), .ZN(
        n19497) );
  AOI22_X1 U21659 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19528), .ZN(n19496) );
  OAI211_X1 U21660 ( .C1(n19521), .C2(n19648), .A(n19497), .B(n19496), .ZN(
        P2_U3163) );
  AOI22_X1 U21661 ( .A1(n19644), .A2(n19527), .B1(n19525), .B2(n19643), .ZN(
        n19499) );
  AOI22_X1 U21662 ( .A1(n19651), .A2(n19526), .B1(n19645), .B2(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n19498) );
  OAI211_X1 U21663 ( .C1(n19524), .C2(n19648), .A(n19499), .B(n19498), .ZN(
        P2_U3155) );
  AOI22_X1 U21664 ( .A1(n19650), .A2(n19527), .B1(n19525), .B2(n19649), .ZN(
        n19501) );
  AOI22_X1 U21665 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19651), .B2(n19528), .ZN(n19500) );
  OAI211_X1 U21666 ( .C1(n19521), .C2(n19660), .A(n19501), .B(n19500), .ZN(
        P2_U3147) );
  AOI22_X1 U21667 ( .A1(n19656), .A2(n19527), .B1(n19525), .B2(n19655), .ZN(
        n19503) );
  AOI22_X1 U21668 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19526), .ZN(n19502) );
  OAI211_X1 U21669 ( .C1(n19524), .C2(n19660), .A(n19503), .B(n19502), .ZN(
        P2_U3139) );
  AOI22_X1 U21670 ( .A1(n19528), .A2(n19662), .B1(n19525), .B2(n19661), .ZN(
        n19505) );
  AOI22_X1 U21671 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19664), .B1(
        n19527), .B2(n19663), .ZN(n19504) );
  OAI211_X1 U21672 ( .C1(n19521), .C2(n19672), .A(n19505), .B(n19504), .ZN(
        P2_U3131) );
  AOI22_X1 U21673 ( .A1(n19526), .A2(n19674), .B1(n19667), .B2(n19525), .ZN(
        n19507) );
  AOI22_X1 U21674 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19669), .B1(
        n19527), .B2(n19668), .ZN(n19506) );
  OAI211_X1 U21675 ( .C1(n19524), .C2(n19672), .A(n19507), .B(n19506), .ZN(
        P2_U3123) );
  AOI22_X1 U21676 ( .A1(n19528), .A2(n19674), .B1(n19673), .B2(n19525), .ZN(
        n19509) );
  AOI22_X1 U21677 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19527), .ZN(n19508) );
  OAI211_X1 U21678 ( .C1(n19521), .C2(n19684), .A(n19509), .B(n19508), .ZN(
        P2_U3115) );
  AOI22_X1 U21679 ( .A1(n19680), .A2(n19527), .B1(n19679), .B2(n19525), .ZN(
        n19511) );
  AOI22_X1 U21680 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n19526), .B2(n19688), .ZN(n19510) );
  OAI211_X1 U21681 ( .C1(n19524), .C2(n19684), .A(n19511), .B(n19510), .ZN(
        P2_U3107) );
  AOI22_X1 U21682 ( .A1(n19526), .A2(n19698), .B1(n19525), .B2(n19691), .ZN(
        n19513) );
  AOI22_X1 U21683 ( .A1(n19693), .A2(n19527), .B1(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n19692), .ZN(n19512) );
  OAI211_X1 U21684 ( .C1(n19524), .C2(n19696), .A(n19513), .B(n19512), .ZN(
        P2_U3091) );
  AOI22_X1 U21685 ( .A1(n19528), .A2(n19698), .B1(n19697), .B2(n19525), .ZN(
        n19515) );
  AOI22_X1 U21686 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19700), .B1(
        n19527), .B2(n19699), .ZN(n19514) );
  OAI211_X1 U21687 ( .C1(n19521), .C2(n19703), .A(n19515), .B(n19514), .ZN(
        P2_U3083) );
  INV_X1 U21688 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n19518) );
  AOI22_X1 U21689 ( .A1(n19528), .A2(n19705), .B1(n19704), .B2(n19525), .ZN(
        n19517) );
  AOI22_X1 U21690 ( .A1(n19527), .A2(n19706), .B1(n19713), .B2(n19526), .ZN(
        n19516) );
  OAI211_X1 U21691 ( .C1(n19710), .C2(n19518), .A(n19517), .B(n19516), .ZN(
        P2_U3075) );
  AOI22_X1 U21692 ( .A1(n19712), .A2(n19527), .B1(n19525), .B2(n19711), .ZN(
        n19520) );
  AOI22_X1 U21693 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19528), .ZN(n19519) );
  OAI211_X1 U21694 ( .C1(n19521), .C2(n19723), .A(n19520), .B(n19519), .ZN(
        P2_U3067) );
  AOI22_X1 U21695 ( .A1(n19719), .A2(n19527), .B1(n19525), .B2(n19718), .ZN(
        n19523) );
  AOI22_X1 U21696 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19526), .ZN(n19522) );
  OAI211_X1 U21697 ( .C1(n19524), .C2(n19723), .A(n19523), .B(n19522), .ZN(
        P2_U3059) );
  AOI22_X1 U21698 ( .A1(n19526), .A2(n19727), .B1(n19726), .B2(n19525), .ZN(
        n19530) );
  AOI22_X1 U21699 ( .A1(n19732), .A2(n19528), .B1(n19730), .B2(n19527), .ZN(
        n19529) );
  OAI211_X1 U21700 ( .C1(n19735), .C2(n19531), .A(n19530), .B(n19529), .ZN(
        P2_U3051) );
  AOI22_X1 U21701 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19631), .ZN(n19565) );
  NOR2_X2 U21702 ( .A1(n19532), .A2(n19625), .ZN(n19568) );
  NOR2_X2 U21703 ( .A1(n12397), .A2(n19627), .ZN(n19566) );
  AOI22_X1 U21704 ( .A1(n19630), .A2(n19568), .B1(n19629), .B2(n19566), .ZN(
        n19534) );
  AOI22_X1 U21705 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19632), .ZN(n19562) );
  INV_X1 U21706 ( .A(n19562), .ZN(n19567) );
  AOI22_X1 U21707 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19633), .B1(
        n19567), .B2(n19639), .ZN(n19533) );
  OAI211_X1 U21708 ( .C1(n19565), .C2(n19636), .A(n19534), .B(n19533), .ZN(
        P2_U3170) );
  AOI22_X1 U21709 ( .A1(n19638), .A2(n19568), .B1(n19566), .B2(n19637), .ZN(
        n19536) );
  AOI22_X1 U21710 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19569), .ZN(n19535) );
  OAI211_X1 U21711 ( .C1(n19562), .C2(n19648), .A(n19536), .B(n19535), .ZN(
        P2_U3162) );
  AOI22_X1 U21712 ( .A1(n19644), .A2(n19568), .B1(n19566), .B2(n19643), .ZN(
        n19538) );
  AOI22_X1 U21713 ( .A1(n19651), .A2(n19567), .B1(n19645), .B2(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19537) );
  OAI211_X1 U21714 ( .C1(n19565), .C2(n19648), .A(n19538), .B(n19537), .ZN(
        P2_U3154) );
  AOI22_X1 U21715 ( .A1(n19650), .A2(n19568), .B1(n19566), .B2(n19649), .ZN(
        n19540) );
  AOI22_X1 U21716 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n19651), .B2(n19569), .ZN(n19539) );
  OAI211_X1 U21717 ( .C1(n19562), .C2(n19660), .A(n19540), .B(n19539), .ZN(
        P2_U3146) );
  AOI22_X1 U21718 ( .A1(n19656), .A2(n19568), .B1(n19566), .B2(n19655), .ZN(
        n19542) );
  AOI22_X1 U21719 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19567), .ZN(n19541) );
  OAI211_X1 U21720 ( .C1(n19565), .C2(n19660), .A(n19542), .B(n19541), .ZN(
        P2_U3138) );
  AOI22_X1 U21721 ( .A1(n19569), .A2(n19662), .B1(n19566), .B2(n19661), .ZN(
        n19544) );
  AOI22_X1 U21722 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19664), .B1(
        n19568), .B2(n19663), .ZN(n19543) );
  OAI211_X1 U21723 ( .C1(n19562), .C2(n19672), .A(n19544), .B(n19543), .ZN(
        P2_U3130) );
  AOI22_X1 U21724 ( .A1(n19567), .A2(n19674), .B1(n19667), .B2(n19566), .ZN(
        n19546) );
  AOI22_X1 U21725 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19669), .B1(
        n19568), .B2(n19668), .ZN(n19545) );
  OAI211_X1 U21726 ( .C1(n19565), .C2(n19672), .A(n19546), .B(n19545), .ZN(
        P2_U3122) );
  AOI22_X1 U21727 ( .A1(n19569), .A2(n19674), .B1(n19673), .B2(n19566), .ZN(
        n19548) );
  AOI22_X1 U21728 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19568), .ZN(n19547) );
  OAI211_X1 U21729 ( .C1(n19562), .C2(n19684), .A(n19548), .B(n19547), .ZN(
        P2_U3114) );
  AOI22_X1 U21730 ( .A1(n19680), .A2(n19568), .B1(n19679), .B2(n19566), .ZN(
        n19550) );
  AOI22_X1 U21731 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n19567), .B2(n19688), .ZN(n19549) );
  OAI211_X1 U21732 ( .C1(n19565), .C2(n19684), .A(n19550), .B(n19549), .ZN(
        P2_U3106) );
  AOI22_X1 U21733 ( .A1(n19686), .A2(n19568), .B1(n19566), .B2(n19685), .ZN(
        n19552) );
  AOI22_X1 U21734 ( .A1(n19569), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n19551) );
  OAI211_X1 U21735 ( .C1(n19562), .C2(n19696), .A(n19552), .B(n19551), .ZN(
        P2_U3098) );
  AOI22_X1 U21736 ( .A1(n19567), .A2(n19698), .B1(n19691), .B2(n19566), .ZN(
        n19554) );
  AOI22_X1 U21737 ( .A1(n19693), .A2(n19568), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n19692), .ZN(n19553) );
  OAI211_X1 U21738 ( .C1(n19565), .C2(n19696), .A(n19554), .B(n19553), .ZN(
        P2_U3090) );
  AOI22_X1 U21739 ( .A1(n19569), .A2(n19698), .B1(n19697), .B2(n19566), .ZN(
        n19556) );
  AOI22_X1 U21740 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19700), .B1(
        n19568), .B2(n19699), .ZN(n19555) );
  OAI211_X1 U21741 ( .C1(n19562), .C2(n19703), .A(n19556), .B(n19555), .ZN(
        P2_U3082) );
  INV_X1 U21742 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19559) );
  AOI22_X1 U21743 ( .A1(n19569), .A2(n19705), .B1(n19704), .B2(n19566), .ZN(
        n19558) );
  AOI22_X1 U21744 ( .A1(n19568), .A2(n19706), .B1(n19713), .B2(n19567), .ZN(
        n19557) );
  OAI211_X1 U21745 ( .C1(n19710), .C2(n19559), .A(n19558), .B(n19557), .ZN(
        P2_U3074) );
  AOI22_X1 U21746 ( .A1(n19712), .A2(n19568), .B1(n19566), .B2(n19711), .ZN(
        n19561) );
  AOI22_X1 U21747 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19569), .ZN(n19560) );
  OAI211_X1 U21748 ( .C1(n19562), .C2(n19723), .A(n19561), .B(n19560), .ZN(
        P2_U3066) );
  AOI22_X1 U21749 ( .A1(n19719), .A2(n19568), .B1(n19566), .B2(n19718), .ZN(
        n19564) );
  AOI22_X1 U21750 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19567), .ZN(n19563) );
  OAI211_X1 U21751 ( .C1(n19565), .C2(n19723), .A(n19564), .B(n19563), .ZN(
        P2_U3058) );
  AOI22_X1 U21752 ( .A1(n19567), .A2(n19727), .B1(n19726), .B2(n19566), .ZN(
        n19571) );
  AOI22_X1 U21753 ( .A1(n19732), .A2(n19569), .B1(n19730), .B2(n19568), .ZN(
        n19570) );
  OAI211_X1 U21754 ( .C1(n19735), .C2(n19572), .A(n19571), .B(n19570), .ZN(
        P2_U3050) );
  AOI22_X1 U21755 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19631), .ZN(n19606) );
  NOR2_X2 U21756 ( .A1(n19573), .A2(n19625), .ZN(n19609) );
  NOR2_X2 U21757 ( .A1(n19574), .A2(n19627), .ZN(n19607) );
  AOI22_X1 U21758 ( .A1(n19630), .A2(n19609), .B1(n19629), .B2(n19607), .ZN(
        n19576) );
  AOI22_X1 U21759 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19631), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19632), .ZN(n19603) );
  INV_X1 U21760 ( .A(n19603), .ZN(n19608) );
  AOI22_X1 U21761 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19633), .B1(
        n19608), .B2(n19639), .ZN(n19575) );
  OAI211_X1 U21762 ( .C1(n19606), .C2(n19636), .A(n19576), .B(n19575), .ZN(
        P2_U3169) );
  AOI22_X1 U21763 ( .A1(n19638), .A2(n19609), .B1(n19607), .B2(n19637), .ZN(
        n19578) );
  AOI22_X1 U21764 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19610), .ZN(n19577) );
  OAI211_X1 U21765 ( .C1(n19603), .C2(n19648), .A(n19578), .B(n19577), .ZN(
        P2_U3161) );
  AOI22_X1 U21766 ( .A1(n19644), .A2(n19609), .B1(n19607), .B2(n19643), .ZN(
        n19580) );
  AOI22_X1 U21767 ( .A1(n19651), .A2(n19608), .B1(n19645), .B2(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n19579) );
  OAI211_X1 U21768 ( .C1(n19606), .C2(n19648), .A(n19580), .B(n19579), .ZN(
        P2_U3153) );
  AOI22_X1 U21769 ( .A1(n19650), .A2(n19609), .B1(n19607), .B2(n19649), .ZN(
        n19582) );
  AOI22_X1 U21770 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n19651), .B2(n19610), .ZN(n19581) );
  OAI211_X1 U21771 ( .C1(n19603), .C2(n19660), .A(n19582), .B(n19581), .ZN(
        P2_U3145) );
  AOI22_X1 U21772 ( .A1(n19656), .A2(n19609), .B1(n19607), .B2(n19655), .ZN(
        n19584) );
  AOI22_X1 U21773 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19608), .ZN(n19583) );
  OAI211_X1 U21774 ( .C1(n19606), .C2(n19660), .A(n19584), .B(n19583), .ZN(
        P2_U3137) );
  AOI22_X1 U21775 ( .A1(n19610), .A2(n19662), .B1(n19607), .B2(n19661), .ZN(
        n19586) );
  AOI22_X1 U21776 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19664), .B1(
        n19609), .B2(n19663), .ZN(n19585) );
  OAI211_X1 U21777 ( .C1(n19603), .C2(n19672), .A(n19586), .B(n19585), .ZN(
        P2_U3129) );
  AOI22_X1 U21778 ( .A1(n19608), .A2(n19674), .B1(n19667), .B2(n19607), .ZN(
        n19588) );
  AOI22_X1 U21779 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19669), .B1(
        n19609), .B2(n19668), .ZN(n19587) );
  OAI211_X1 U21780 ( .C1(n19606), .C2(n19672), .A(n19588), .B(n19587), .ZN(
        P2_U3121) );
  AOI22_X1 U21781 ( .A1(n19610), .A2(n19674), .B1(n19673), .B2(n19607), .ZN(
        n19590) );
  AOI22_X1 U21782 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19609), .ZN(n19589) );
  OAI211_X1 U21783 ( .C1(n19603), .C2(n19684), .A(n19590), .B(n19589), .ZN(
        P2_U3113) );
  AOI22_X1 U21784 ( .A1(n19680), .A2(n19609), .B1(n19679), .B2(n19607), .ZN(
        n19592) );
  AOI22_X1 U21785 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n19608), .B2(n19688), .ZN(n19591) );
  OAI211_X1 U21786 ( .C1(n19606), .C2(n19684), .A(n19592), .B(n19591), .ZN(
        P2_U3105) );
  AOI22_X1 U21787 ( .A1(n19686), .A2(n19609), .B1(n19607), .B2(n19685), .ZN(
        n19594) );
  AOI22_X1 U21788 ( .A1(n19610), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19593) );
  OAI211_X1 U21789 ( .C1(n19603), .C2(n19696), .A(n19594), .B(n19593), .ZN(
        P2_U3097) );
  AOI22_X1 U21790 ( .A1(n19608), .A2(n19698), .B1(n19691), .B2(n19607), .ZN(
        n19596) );
  AOI22_X1 U21791 ( .A1(n19693), .A2(n19609), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n19692), .ZN(n19595) );
  OAI211_X1 U21792 ( .C1(n19606), .C2(n19696), .A(n19596), .B(n19595), .ZN(
        P2_U3089) );
  AOI22_X1 U21793 ( .A1(n19610), .A2(n19698), .B1(n19697), .B2(n19607), .ZN(
        n19598) );
  AOI22_X1 U21794 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19700), .B1(
        n19609), .B2(n19699), .ZN(n19597) );
  OAI211_X1 U21795 ( .C1(n19603), .C2(n19703), .A(n19598), .B(n19597), .ZN(
        P2_U3081) );
  AOI22_X1 U21796 ( .A1(n19610), .A2(n19705), .B1(n19704), .B2(n19607), .ZN(
        n19600) );
  AOI22_X1 U21797 ( .A1(n19609), .A2(n19706), .B1(n19713), .B2(n19608), .ZN(
        n19599) );
  OAI211_X1 U21798 ( .C1(n19710), .C2(n13647), .A(n19600), .B(n19599), .ZN(
        P2_U3073) );
  AOI22_X1 U21799 ( .A1(n19712), .A2(n19609), .B1(n19607), .B2(n19711), .ZN(
        n19602) );
  AOI22_X1 U21800 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19610), .ZN(n19601) );
  OAI211_X1 U21801 ( .C1(n19603), .C2(n19723), .A(n19602), .B(n19601), .ZN(
        P2_U3065) );
  AOI22_X1 U21802 ( .A1(n19719), .A2(n19609), .B1(n19607), .B2(n19718), .ZN(
        n19605) );
  AOI22_X1 U21803 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19608), .ZN(n19604) );
  OAI211_X1 U21804 ( .C1(n19606), .C2(n19723), .A(n19605), .B(n19604), .ZN(
        P2_U3057) );
  AOI22_X1 U21805 ( .A1(n19608), .A2(n19727), .B1(n19726), .B2(n19607), .ZN(
        n19612) );
  AOI22_X1 U21806 ( .A1(n19732), .A2(n19610), .B1(n19730), .B2(n19609), .ZN(
        n19611) );
  OAI211_X1 U21807 ( .C1(n19735), .C2(n13651), .A(n19612), .B(n19611), .ZN(
        P2_U3049) );
  AOI22_X1 U21808 ( .A1(n19615), .A2(n19614), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19613), .ZN(n19624) );
  AOI22_X1 U21809 ( .A1(n19617), .A2(BUF2_REG_16__SCAN_IN), .B1(n19616), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U21810 ( .A1(n19621), .A2(n19620), .B1(n19619), .B2(n19618), .ZN(
        n19622) );
  NAND3_X1 U21811 ( .A1(n19624), .A2(n19623), .A3(n19622), .ZN(P2_U2903) );
  AOI22_X1 U21812 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19631), .ZN(n19724) );
  NOR2_X2 U21813 ( .A1(n19626), .A2(n19625), .ZN(n19729) );
  NOR2_X2 U21814 ( .A1(n19628), .A2(n19627), .ZN(n19725) );
  AOI22_X1 U21815 ( .A1(n19630), .A2(n19729), .B1(n19629), .B2(n19725), .ZN(
        n19635) );
  AOI22_X1 U21816 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19632), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19631), .ZN(n19717) );
  INV_X1 U21817 ( .A(n19717), .ZN(n19728) );
  AOI22_X1 U21818 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19633), .B1(
        n19728), .B2(n19639), .ZN(n19634) );
  OAI211_X1 U21819 ( .C1(n19724), .C2(n19636), .A(n19635), .B(n19634), .ZN(
        P2_U3168) );
  AOI22_X1 U21820 ( .A1(n19638), .A2(n19729), .B1(n19725), .B2(n19637), .ZN(
        n19642) );
  AOI22_X1 U21821 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19731), .ZN(n19641) );
  OAI211_X1 U21822 ( .C1(n19717), .C2(n19648), .A(n19642), .B(n19641), .ZN(
        P2_U3160) );
  AOI22_X1 U21823 ( .A1(n19644), .A2(n19729), .B1(n19725), .B2(n19643), .ZN(
        n19647) );
  AOI22_X1 U21824 ( .A1(n19651), .A2(n19728), .B1(n19645), .B2(
        P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19646) );
  OAI211_X1 U21825 ( .C1(n19724), .C2(n19648), .A(n19647), .B(n19646), .ZN(
        P2_U3152) );
  AOI22_X1 U21826 ( .A1(n19650), .A2(n19729), .B1(n19725), .B2(n19649), .ZN(
        n19654) );
  AOI22_X1 U21827 ( .A1(n19652), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n19651), .B2(n19731), .ZN(n19653) );
  OAI211_X1 U21828 ( .C1(n19717), .C2(n19660), .A(n19654), .B(n19653), .ZN(
        P2_U3144) );
  AOI22_X1 U21829 ( .A1(n19656), .A2(n19729), .B1(n19725), .B2(n19655), .ZN(
        n19659) );
  AOI22_X1 U21830 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19657), .B1(
        n19662), .B2(n19728), .ZN(n19658) );
  OAI211_X1 U21831 ( .C1(n19724), .C2(n19660), .A(n19659), .B(n19658), .ZN(
        P2_U3136) );
  AOI22_X1 U21832 ( .A1(n19731), .A2(n19662), .B1(n19725), .B2(n19661), .ZN(
        n19666) );
  AOI22_X1 U21833 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19664), .B1(
        n19729), .B2(n19663), .ZN(n19665) );
  OAI211_X1 U21834 ( .C1(n19717), .C2(n19672), .A(n19666), .B(n19665), .ZN(
        P2_U3128) );
  AOI22_X1 U21835 ( .A1(n19728), .A2(n19674), .B1(n19667), .B2(n19725), .ZN(
        n19671) );
  AOI22_X1 U21836 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19669), .B1(
        n19729), .B2(n19668), .ZN(n19670) );
  OAI211_X1 U21837 ( .C1(n19724), .C2(n19672), .A(n19671), .B(n19670), .ZN(
        P2_U3120) );
  AOI22_X1 U21838 ( .A1(n19731), .A2(n19674), .B1(n19673), .B2(n19725), .ZN(
        n19678) );
  AOI22_X1 U21839 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19676), .B1(
        n19675), .B2(n19729), .ZN(n19677) );
  OAI211_X1 U21840 ( .C1(n19717), .C2(n19684), .A(n19678), .B(n19677), .ZN(
        P2_U3112) );
  AOI22_X1 U21841 ( .A1(n19680), .A2(n19729), .B1(n19679), .B2(n19725), .ZN(
        n19683) );
  AOI22_X1 U21842 ( .A1(n19681), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n19728), .B2(n19688), .ZN(n19682) );
  OAI211_X1 U21843 ( .C1(n19724), .C2(n19684), .A(n19683), .B(n19682), .ZN(
        P2_U3104) );
  AOI22_X1 U21844 ( .A1(n19686), .A2(n19729), .B1(n19725), .B2(n19685), .ZN(
        n19690) );
  AOI22_X1 U21845 ( .A1(n19731), .A2(n19688), .B1(n19687), .B2(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19689) );
  OAI211_X1 U21846 ( .C1(n19717), .C2(n19696), .A(n19690), .B(n19689), .ZN(
        P2_U3096) );
  AOI22_X1 U21847 ( .A1(n19728), .A2(n19698), .B1(n19691), .B2(n19725), .ZN(
        n19695) );
  AOI22_X1 U21848 ( .A1(n19693), .A2(n19729), .B1(
        P2_INSTQUEUE_REG_5__0__SCAN_IN), .B2(n19692), .ZN(n19694) );
  OAI211_X1 U21849 ( .C1(n19724), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P2_U3088) );
  AOI22_X1 U21850 ( .A1(n19731), .A2(n19698), .B1(n19697), .B2(n19725), .ZN(
        n19702) );
  AOI22_X1 U21851 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19700), .B1(
        n19729), .B2(n19699), .ZN(n19701) );
  OAI211_X1 U21852 ( .C1(n19717), .C2(n19703), .A(n19702), .B(n19701), .ZN(
        P2_U3080) );
  INV_X1 U21853 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U21854 ( .A1(n19731), .A2(n19705), .B1(n19704), .B2(n19725), .ZN(
        n19708) );
  AOI22_X1 U21855 ( .A1(n19729), .A2(n19706), .B1(n19713), .B2(n19728), .ZN(
        n19707) );
  OAI211_X1 U21856 ( .C1(n19710), .C2(n19709), .A(n19708), .B(n19707), .ZN(
        P2_U3072) );
  AOI22_X1 U21857 ( .A1(n19712), .A2(n19729), .B1(n19725), .B2(n19711), .ZN(
        n19716) );
  AOI22_X1 U21858 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19731), .ZN(n19715) );
  OAI211_X1 U21859 ( .C1(n19717), .C2(n19723), .A(n19716), .B(n19715), .ZN(
        P2_U3064) );
  AOI22_X1 U21860 ( .A1(n19719), .A2(n19729), .B1(n19725), .B2(n19718), .ZN(
        n19722) );
  AOI22_X1 U21861 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19720), .B1(
        n19732), .B2(n19728), .ZN(n19721) );
  OAI211_X1 U21862 ( .C1(n19724), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P2_U3056) );
  AOI22_X1 U21863 ( .A1(n19728), .A2(n19727), .B1(n19726), .B2(n19725), .ZN(
        n19734) );
  AOI22_X1 U21864 ( .A1(n19732), .A2(n19731), .B1(n19730), .B2(n19729), .ZN(
        n19733) );
  OAI211_X1 U21865 ( .C1(n19735), .C2(n12715), .A(n19734), .B(n19733), .ZN(
        P2_U3048) );
  INV_X1 U21866 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20048) );
  INV_X1 U21867 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19736) );
  AOI222_X1 U21868 ( .A1(n20048), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20051), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19736), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19737) );
  INV_X1 U21869 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U21870 ( .A1(n19786), .A2(n19739), .B1(n19738), .B2(n19797), .ZN(
        U376) );
  INV_X1 U21871 ( .A(n19797), .ZN(n19800) );
  INV_X1 U21872 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U21873 ( .A1(n19800), .A2(n19741), .B1(n19740), .B2(n19797), .ZN(
        U365) );
  INV_X1 U21874 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U21875 ( .A1(n19786), .A2(n19743), .B1(n19742), .B2(n19797), .ZN(
        U354) );
  INV_X1 U21876 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U21877 ( .A1(n19786), .A2(n19745), .B1(n19744), .B2(n19797), .ZN(
        U353) );
  INV_X1 U21878 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U21879 ( .A1(n19786), .A2(n19747), .B1(n19746), .B2(n19797), .ZN(
        U352) );
  INV_X1 U21880 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U21881 ( .A1(n19786), .A2(n19749), .B1(n19748), .B2(n19797), .ZN(
        U351) );
  INV_X1 U21882 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U21883 ( .A1(n19800), .A2(n19751), .B1(n19750), .B2(n19797), .ZN(
        U350) );
  INV_X1 U21884 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U21885 ( .A1(n19786), .A2(n19753), .B1(n19752), .B2(n19797), .ZN(
        U349) );
  INV_X1 U21886 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U21887 ( .A1(n19786), .A2(n19755), .B1(n19754), .B2(n19797), .ZN(
        U348) );
  INV_X1 U21888 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U21889 ( .A1(n19786), .A2(n19757), .B1(n19756), .B2(n19797), .ZN(
        U347) );
  INV_X1 U21890 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U21891 ( .A1(n19786), .A2(n19759), .B1(n19758), .B2(n19797), .ZN(
        U375) );
  INV_X1 U21892 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U21893 ( .A1(n19786), .A2(n19761), .B1(n19760), .B2(n19797), .ZN(
        U374) );
  INV_X1 U21894 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U21895 ( .A1(n19786), .A2(n19763), .B1(n19762), .B2(n19797), .ZN(
        U373) );
  INV_X1 U21896 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U21897 ( .A1(n19786), .A2(n19765), .B1(n19764), .B2(n19797), .ZN(
        U372) );
  INV_X1 U21898 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U21899 ( .A1(n19786), .A2(n19767), .B1(n19766), .B2(n19797), .ZN(
        U371) );
  INV_X1 U21900 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U21901 ( .A1(n19786), .A2(n19769), .B1(n19768), .B2(n19797), .ZN(
        U370) );
  INV_X1 U21902 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U21903 ( .A1(n19786), .A2(n19771), .B1(n19770), .B2(n19797), .ZN(
        U369) );
  INV_X1 U21904 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U21905 ( .A1(n19786), .A2(n19773), .B1(n19772), .B2(n19797), .ZN(
        U368) );
  INV_X1 U21906 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U21907 ( .A1(n19786), .A2(n19775), .B1(n19774), .B2(n19797), .ZN(
        U367) );
  INV_X1 U21908 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U21909 ( .A1(n19786), .A2(n19777), .B1(n19776), .B2(n19797), .ZN(
        U366) );
  INV_X1 U21910 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U21911 ( .A1(n19786), .A2(n19779), .B1(n19778), .B2(n19797), .ZN(
        U364) );
  INV_X1 U21912 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U21913 ( .A1(n19786), .A2(n19781), .B1(n19780), .B2(n19797), .ZN(
        U363) );
  INV_X1 U21914 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19783) );
  AOI22_X1 U21915 ( .A1(n19786), .A2(n19783), .B1(n19782), .B2(n19797), .ZN(
        U362) );
  INV_X1 U21916 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U21917 ( .A1(n19786), .A2(n19785), .B1(n19784), .B2(n19797), .ZN(
        U361) );
  INV_X1 U21918 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U21919 ( .A1(n19800), .A2(n19788), .B1(n19787), .B2(n19797), .ZN(
        U360) );
  INV_X1 U21920 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U21921 ( .A1(n19800), .A2(n19790), .B1(n19789), .B2(n19797), .ZN(
        U359) );
  INV_X1 U21922 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U21923 ( .A1(n19800), .A2(n19792), .B1(n19791), .B2(n19797), .ZN(
        U358) );
  INV_X1 U21924 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U21925 ( .A1(n19800), .A2(n19794), .B1(n19793), .B2(n19797), .ZN(
        U357) );
  INV_X1 U21926 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U21927 ( .A1(n19800), .A2(n19796), .B1(n19795), .B2(n19797), .ZN(
        U356) );
  INV_X1 U21928 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U21929 ( .A1(n19800), .A2(n19799), .B1(n19798), .B2(n19797), .ZN(
        U355) );
  AOI22_X1 U21930 ( .A1(n21288), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19802) );
  OAI21_X1 U21931 ( .B1(n21780), .B2(n19820), .A(n19802), .ZN(P1_U2936) );
  AOI22_X1 U21932 ( .A1(n19811), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U21933 ( .B1(n21786), .B2(n19820), .A(n19803), .ZN(P1_U2935) );
  AOI22_X1 U21934 ( .A1(n19811), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19804) );
  OAI21_X1 U21935 ( .B1(n21792), .B2(n19820), .A(n19804), .ZN(P1_U2934) );
  AOI22_X1 U21936 ( .A1(n19811), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U21937 ( .B1(n21798), .B2(n19820), .A(n19805), .ZN(P1_U2933) );
  AOI22_X1 U21938 ( .A1(n19811), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19806) );
  OAI21_X1 U21939 ( .B1(n21804), .B2(n19820), .A(n19806), .ZN(P1_U2932) );
  INV_X1 U21940 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n21811) );
  AOI22_X1 U21941 ( .A1(n19811), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U21942 ( .B1(n21811), .B2(n19820), .A(n19807), .ZN(P1_U2931) );
  AOI22_X1 U21943 ( .A1(n19811), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U21944 ( .B1(n11794), .B2(n19820), .A(n19809), .ZN(P1_U2930) );
  AOI22_X1 U21945 ( .A1(n21288), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19810) );
  OAI21_X1 U21946 ( .B1(n11816), .B2(n19820), .A(n19810), .ZN(P1_U2929) );
  AOI22_X1 U21947 ( .A1(n19811), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19812) );
  OAI21_X1 U21948 ( .B1(n15032), .B2(n19820), .A(n19812), .ZN(P1_U2928) );
  AOI22_X1 U21949 ( .A1(n21288), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U21950 ( .B1(n15018), .B2(n19820), .A(n19813), .ZN(P1_U2927) );
  INV_X1 U21951 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21837) );
  AOI22_X1 U21952 ( .A1(n21288), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19814) );
  OAI21_X1 U21953 ( .B1(n21837), .B2(n19820), .A(n19814), .ZN(P1_U2926) );
  AOI22_X1 U21954 ( .A1(n21288), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19815) );
  OAI21_X1 U21955 ( .B1(n15205), .B2(n19820), .A(n19815), .ZN(P1_U2925) );
  AOI22_X1 U21956 ( .A1(n21288), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19816) );
  OAI21_X1 U21957 ( .B1(n15226), .B2(n19820), .A(n19816), .ZN(P1_U2924) );
  INV_X1 U21958 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21854) );
  AOI22_X1 U21959 ( .A1(n21288), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19817) );
  OAI21_X1 U21960 ( .B1(n21854), .B2(n19820), .A(n19817), .ZN(P1_U2923) );
  INV_X1 U21961 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21864) );
  AOI22_X1 U21962 ( .A1(n21288), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19818) );
  OAI21_X1 U21963 ( .B1(n21864), .B2(n19820), .A(n19818), .ZN(P1_U2922) );
  AOI22_X1 U21964 ( .A1(n21288), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19808), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19819) );
  OAI21_X1 U21965 ( .B1(n14216), .B2(n19820), .A(n19819), .ZN(P1_U2921) );
  OAI222_X1 U21966 ( .A1(n19860), .A2(n14718), .B1(n19821), .B2(n22339), .C1(
        n14367), .C2(n21720), .ZN(P1_U3197) );
  AOI222_X1 U21967 ( .A1(n19855), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n19858), .ZN(n19822) );
  INV_X1 U21968 ( .A(n19822), .ZN(P1_U3198) );
  AOI222_X1 U21969 ( .A1(n19855), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n19858), .ZN(n19823) );
  INV_X1 U21970 ( .A(n19823), .ZN(P1_U3199) );
  INV_X1 U21971 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n19824) );
  INV_X1 U21972 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21488) );
  OAI222_X1 U21973 ( .A1(n19860), .A2(n21506), .B1(n19824), .B2(n22339), .C1(
        n21488), .C2(n21720), .ZN(P1_U3200) );
  AOI22_X1 U21974 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19855), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n22337), .ZN(n19825) );
  OAI21_X1 U21975 ( .B1(n21506), .B2(n21720), .A(n19825), .ZN(P1_U3201) );
  AOI22_X1 U21976 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19858), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n22337), .ZN(n19826) );
  OAI21_X1 U21977 ( .B1(n21529), .B2(n19860), .A(n19826), .ZN(P1_U3202) );
  AOI22_X1 U21978 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19855), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n22337), .ZN(n19827) );
  OAI21_X1 U21979 ( .B1(n21529), .B2(n21720), .A(n19827), .ZN(P1_U3203) );
  AOI22_X1 U21980 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19858), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n22337), .ZN(n19828) );
  OAI21_X1 U21981 ( .B1(n21552), .B2(n19860), .A(n19828), .ZN(P1_U3204) );
  AOI22_X1 U21982 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19855), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22337), .ZN(n19829) );
  OAI21_X1 U21983 ( .B1(n21552), .B2(n21720), .A(n19829), .ZN(P1_U3205) );
  AOI22_X1 U21984 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19858), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n22337), .ZN(n19830) );
  OAI21_X1 U21985 ( .B1(n21576), .B2(n19860), .A(n19830), .ZN(P1_U3206) );
  INV_X1 U21986 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n19831) );
  OAI222_X1 U21987 ( .A1(n19860), .A2(n21580), .B1(n19831), .B2(n22339), .C1(
        n21576), .C2(n21720), .ZN(P1_U3207) );
  AOI222_X1 U21988 ( .A1(n19858), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n19855), .ZN(n19832) );
  INV_X1 U21989 ( .A(n19832), .ZN(P1_U3208) );
  AOI222_X1 U21990 ( .A1(n19858), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n19855), .ZN(n19833) );
  INV_X1 U21991 ( .A(n19833), .ZN(P1_U3209) );
  AOI22_X1 U21992 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19855), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n22337), .ZN(n19834) );
  OAI21_X1 U21993 ( .B1(n21310), .B2(n21720), .A(n19834), .ZN(P1_U3210) );
  AOI22_X1 U21994 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19858), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22337), .ZN(n19835) );
  OAI21_X1 U21995 ( .B1(n21600), .B2(n19860), .A(n19835), .ZN(P1_U3211) );
  INV_X1 U21996 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n19836) );
  OAI222_X1 U21997 ( .A1(n19860), .A2(n15841), .B1(n19836), .B2(n22339), .C1(
        n21600), .C2(n21720), .ZN(P1_U3212) );
  INV_X1 U21998 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n19837) );
  OAI222_X1 U21999 ( .A1(n19860), .A2(n21428), .B1(n19837), .B2(n22339), .C1(
        n15841), .C2(n21720), .ZN(P1_U3213) );
  INV_X1 U22000 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n19839) );
  OAI222_X1 U22001 ( .A1(n21720), .A2(n21428), .B1(n19839), .B2(n22339), .C1(
        n19838), .C2(n19860), .ZN(P1_U3214) );
  AOI222_X1 U22002 ( .A1(n19855), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n19858), .ZN(n19840) );
  INV_X1 U22003 ( .A(n19840), .ZN(P1_U3215) );
  AOI222_X1 U22004 ( .A1(n19855), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n22337), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n19858), .ZN(n19841) );
  INV_X1 U22005 ( .A(n19841), .ZN(P1_U3216) );
  INV_X1 U22006 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n19843) );
  OAI222_X1 U22007 ( .A1(n19860), .A2(n21635), .B1(n19843), .B2(n22339), .C1(
        n19842), .C2(n21720), .ZN(P1_U3217) );
  INV_X1 U22008 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n19844) );
  OAI222_X1 U22009 ( .A1(n19860), .A2(n19846), .B1(n19844), .B2(n22339), .C1(
        n21635), .C2(n21720), .ZN(P1_U3218) );
  INV_X1 U22010 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n19845) );
  OAI222_X1 U22011 ( .A1(n21720), .A2(n19846), .B1(n19845), .B2(n22339), .C1(
        n21655), .C2(n19860), .ZN(P1_U3219) );
  INV_X1 U22012 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n19847) );
  OAI222_X1 U22013 ( .A1(n21720), .A2(n21655), .B1(n19847), .B2(n22339), .C1(
        n19849), .C2(n19860), .ZN(P1_U3220) );
  INV_X1 U22014 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U22015 ( .A1(n21720), .A2(n19849), .B1(n19848), .B2(n22339), .C1(
        n15543), .C2(n19860), .ZN(P1_U3221) );
  INV_X1 U22016 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n19850) );
  OAI222_X1 U22017 ( .A1(n21720), .A2(n15543), .B1(n19850), .B2(n22339), .C1(
        n19851), .C2(n19860), .ZN(P1_U3222) );
  INV_X1 U22018 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n19852) );
  OAI222_X1 U22019 ( .A1(n19860), .A2(n19854), .B1(n19852), .B2(n22339), .C1(
        n19851), .C2(n21720), .ZN(P1_U3223) );
  INV_X1 U22020 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n19853) );
  OAI222_X1 U22021 ( .A1(n21720), .A2(n19854), .B1(n19853), .B2(n22339), .C1(
        n19857), .C2(n19860), .ZN(P1_U3224) );
  AOI22_X1 U22022 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19855), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n22337), .ZN(n19856) );
  OAI21_X1 U22023 ( .B1(n19857), .B2(n21720), .A(n19856), .ZN(P1_U3225) );
  AOI22_X1 U22024 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19858), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22337), .ZN(n19859) );
  OAI21_X1 U22025 ( .B1(n19861), .B2(n19860), .A(n19859), .ZN(P1_U3226) );
  OAI22_X1 U22026 ( .A1(n22337), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22339), .ZN(n19862) );
  INV_X1 U22027 ( .A(n19862), .ZN(P1_U3458) );
  NOR4_X1 U22028 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19866) );
  NOR4_X1 U22029 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19865) );
  NOR4_X1 U22030 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19864) );
  NOR4_X1 U22031 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19863) );
  NAND4_X1 U22032 ( .A1(n19866), .A2(n19865), .A3(n19864), .A4(n19863), .ZN(
        n19872) );
  NOR4_X1 U22033 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19870) );
  AOI211_X1 U22034 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19869) );
  NOR4_X1 U22035 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19868) );
  NOR4_X1 U22036 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19867) );
  NAND4_X1 U22037 ( .A1(n19870), .A2(n19869), .A3(n19868), .A4(n19867), .ZN(
        n19871) );
  NOR2_X1 U22038 ( .A1(n19872), .A2(n19871), .ZN(n19884) );
  NAND2_X1 U22039 ( .A1(n19884), .A2(n14367), .ZN(n19877) );
  INV_X1 U22040 ( .A(n19884), .ZN(n19887) );
  NAND2_X1 U22041 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(n19887), .ZN(n19873) );
  NOR2_X1 U22042 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19876) );
  NAND3_X1 U22043 ( .A1(n19884), .A2(n19876), .A3(n14291), .ZN(n19882) );
  OAI211_X1 U22044 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(n19877), .A(n19873), 
        .B(n19882), .ZN(P1_U2808) );
  INV_X1 U22045 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U22046 ( .A1(n22339), .A2(n19875), .B1(n19874), .B2(n22337), .ZN(
        P1_U3459) );
  AOI22_X1 U22047 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n19876), .B2(n14367), .ZN(n19880) );
  NOR2_X1 U22048 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n19877), .ZN(n19886) );
  NAND2_X1 U22049 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(n19886), .ZN(n19879)
         );
  NAND2_X1 U22050 ( .A1(n19887), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19878) );
  OAI211_X1 U22051 ( .C1(n19887), .C2(n19880), .A(n19879), .B(n19878), .ZN(
        P1_U3481) );
  INV_X1 U22052 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U22053 ( .A1(n22339), .A2(n19883), .B1(n19881), .B2(n22337), .ZN(
        P1_U3460) );
  OAI221_X1 U22054 ( .B1(n19884), .B2(n19883), .C1(n19887), .C2(n14367), .A(
        n19882), .ZN(P1_U2807) );
  INV_X1 U22055 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U22056 ( .A1(n22339), .A2(n19888), .B1(n19885), .B2(n22337), .ZN(
        P1_U3461) );
  AOI21_X1 U22057 ( .B1(n19888), .B2(n19887), .A(n19886), .ZN(P1_U3482) );
  INV_X1 U22058 ( .A(n19889), .ZN(n21583) );
  XNOR2_X1 U22059 ( .A(n19891), .B(n19890), .ZN(n21578) );
  AOI22_X1 U22060 ( .A1(n21583), .A2(n19908), .B1(n13472), .B2(n21578), .ZN(
        n19892) );
  OAI21_X1 U22061 ( .B1(n19911), .B2(n21581), .A(n19892), .ZN(P1_U2860) );
  XOR2_X1 U22062 ( .A(n19894), .B(n19893), .Z(n21555) );
  AOI22_X1 U22063 ( .A1(n19940), .A2(n19908), .B1(n13472), .B2(n21555), .ZN(
        n19895) );
  OAI21_X1 U22064 ( .B1(n19911), .B2(n21566), .A(n19895), .ZN(P1_U2862) );
  INV_X1 U22065 ( .A(n19907), .ZN(n19898) );
  AOI21_X1 U22066 ( .B1(n19898), .B2(n19897), .A(n19896), .ZN(n19900) );
  OR2_X1 U22067 ( .A1(n19900), .A2(n19899), .ZN(n21520) );
  NOR2_X1 U22068 ( .A1(n21520), .A2(n15657), .ZN(n19901) );
  AOI21_X1 U22069 ( .B1(n21526), .B2(n19908), .A(n19901), .ZN(n19902) );
  OAI21_X1 U22070 ( .B1(n19911), .B2(n19903), .A(n19902), .ZN(P1_U2865) );
  NAND2_X1 U22071 ( .A1(n19905), .A2(n19904), .ZN(n19906) );
  AND2_X1 U22072 ( .A1(n19907), .A2(n19906), .ZN(n21496) );
  AOI22_X1 U22073 ( .A1(n21498), .A2(n19908), .B1(n13472), .B2(n21496), .ZN(
        n19909) );
  OAI21_X1 U22074 ( .B1(n19911), .B2(n19910), .A(n19909), .ZN(P1_U2867) );
  AOI22_X1 U22075 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19916) );
  XOR2_X1 U22076 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n19912), .Z(
        n19913) );
  XNOR2_X1 U22077 ( .A(n19914), .B(n19913), .ZN(n21331) );
  AOI22_X1 U22078 ( .A1(n21331), .A2(n19978), .B1(n19979), .B2(n21490), .ZN(
        n19915) );
  OAI211_X1 U22079 ( .C1(n21493), .C2(n19982), .A(n19916), .B(n19915), .ZN(
        P1_U2995) );
  AOI22_X1 U22080 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n19922) );
  INV_X1 U22081 ( .A(n19918), .ZN(n19919) );
  AOI21_X1 U22082 ( .B1(n19920), .B2(n19917), .A(n19919), .ZN(n21364) );
  AOI22_X1 U22083 ( .A1(n21364), .A2(n19978), .B1(n19979), .B2(n21498), .ZN(
        n19921) );
  OAI211_X1 U22084 ( .C1(n21499), .C2(n19982), .A(n19922), .B(n19921), .ZN(
        P1_U2994) );
  AOI22_X1 U22085 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n19928) );
  NAND2_X1 U22086 ( .A1(n19924), .A2(n19923), .ZN(n19925) );
  NAND2_X1 U22087 ( .A1(n19926), .A2(n19925), .ZN(n21354) );
  AOI22_X1 U22088 ( .A1(n21354), .A2(n19978), .B1(n19979), .B2(n21514), .ZN(
        n19927) );
  OAI211_X1 U22089 ( .C1(n21512), .C2(n19982), .A(n19928), .B(n19927), .ZN(
        P1_U2993) );
  AOI22_X1 U22090 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n19934) );
  INV_X1 U22091 ( .A(n19929), .ZN(n19930) );
  AOI21_X1 U22092 ( .B1(n19932), .B2(n19931), .A(n19930), .ZN(n21373) );
  AOI22_X1 U22093 ( .A1(n21373), .A2(n19978), .B1(n19979), .B2(n21526), .ZN(
        n19933) );
  OAI211_X1 U22094 ( .C1(n21524), .C2(n19982), .A(n19934), .B(n19933), .ZN(
        P1_U2992) );
  MUX2_X1 U22095 ( .A(n11346), .B(n15870), .S(n10972), .Z(n19937) );
  INV_X1 U22096 ( .A(n19937), .ZN(n19939) );
  INV_X1 U22097 ( .A(n19943), .ZN(n19938) );
  OAI21_X1 U22098 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19939), .A(
        n19938), .ZN(n21404) );
  AOI22_X1 U22099 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n19942) );
  AOI22_X1 U22100 ( .A1(n19940), .A2(n19979), .B1(n19965), .B2(n21560), .ZN(
        n19941) );
  OAI211_X1 U22101 ( .C1(n21667), .C2(n21404), .A(n19942), .B(n19941), .ZN(
        P1_U2989) );
  NOR2_X1 U22102 ( .A1(n21616), .A2(n21576), .ZN(n21416) );
  OAI22_X1 U22103 ( .A1(n21422), .A2(n21667), .B1(n21575), .B2(n19982), .ZN(
        n19944) );
  OAI21_X1 U22104 ( .B1(n19947), .B2(n19946), .A(n19945), .ZN(P1_U2988) );
  INV_X1 U22105 ( .A(n19948), .ZN(n19953) );
  OAI21_X1 U22106 ( .B1(n13559), .B2(n19950), .A(n19949), .ZN(n19952) );
  AOI21_X1 U22107 ( .B1(n19953), .B2(n19952), .A(n19951), .ZN(n21415) );
  AOI22_X1 U22108 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U22109 ( .A1(n21584), .A2(n19965), .B1(n19979), .B2(n21583), .ZN(
        n19954) );
  OAI211_X1 U22110 ( .C1(n21415), .C2(n21667), .A(n19955), .B(n19954), .ZN(
        P1_U2987) );
  MUX2_X1 U22111 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n13561), .S(
        n13550), .Z(n19963) );
  INV_X1 U22112 ( .A(n19956), .ZN(n19958) );
  NAND3_X1 U22113 ( .A1(n19959), .A2(n19958), .A3(n19957), .ZN(n19961) );
  NAND2_X1 U22114 ( .A1(n19961), .A2(n19960), .ZN(n19962) );
  XOR2_X1 U22115 ( .A(n19963), .B(n19962), .Z(n21318) );
  AOI22_X1 U22116 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U22117 ( .A1(n19966), .A2(n19979), .B1(n19965), .B2(n19964), .ZN(
        n19967) );
  OAI211_X1 U22118 ( .C1(n21318), .C2(n21667), .A(n19968), .B(n19967), .ZN(
        P1_U2985) );
  AOI22_X1 U22119 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U22120 ( .A1(n19969), .A2(n19978), .B1(n19979), .B2(n21612), .ZN(
        n19970) );
  OAI211_X1 U22121 ( .C1(n21605), .C2(n19982), .A(n19971), .B(n19970), .ZN(
        P1_U2983) );
  AOI22_X1 U22122 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n19974) );
  AOI22_X1 U22123 ( .A1(n19972), .A2(n19978), .B1(n19979), .B2(n21631), .ZN(
        n19973) );
  OAI211_X1 U22124 ( .C1(n19975), .C2(n19982), .A(n19974), .B(n19973), .ZN(
        P1_U2979) );
  AOI22_X1 U22125 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19976), .B1(
        n21457), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22126 ( .A1(n21646), .A2(n19979), .B1(n19978), .B2(n19977), .ZN(
        n19980) );
  OAI211_X1 U22127 ( .C1(n21643), .C2(n19982), .A(n19981), .B(n19980), .ZN(
        P1_U2977) );
  INV_X1 U22128 ( .A(n19983), .ZN(n19984) );
  OAI21_X1 U22129 ( .B1(n19984), .B2(n21692), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19985) );
  OAI21_X1 U22130 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19986), .A(n19985), 
        .ZN(P1_U2803) );
  NOR2_X1 U22131 ( .A1(n22339), .A2(n21715), .ZN(n19987) );
  AOI22_X1 U22132 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22339), .B1(n19988), 
        .B2(n19987), .ZN(P1_U2804) );
  AOI22_X1 U22133 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10993), .ZN(n19990) );
  OAI21_X1 U22134 ( .B1(n19991), .B2(n20050), .A(n19990), .ZN(U247) );
  AOI22_X1 U22135 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10993), .ZN(n19992) );
  OAI21_X1 U22136 ( .B1(n14511), .B2(n20050), .A(n19992), .ZN(U246) );
  INV_X1 U22137 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n19994) );
  AOI22_X1 U22138 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10993), .ZN(n19993) );
  OAI21_X1 U22139 ( .B1(n19994), .B2(n20050), .A(n19993), .ZN(U245) );
  AOI22_X1 U22140 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10993), .ZN(n19995) );
  OAI21_X1 U22141 ( .B1(n14583), .B2(n20050), .A(n19995), .ZN(U244) );
  AOI22_X1 U22142 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10993), .ZN(n19996) );
  OAI21_X1 U22143 ( .B1(n19997), .B2(n20050), .A(n19996), .ZN(U243) );
  INV_X1 U22144 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U22145 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10993), .ZN(n19998) );
  OAI21_X1 U22146 ( .B1(n19999), .B2(n20050), .A(n19998), .ZN(U242) );
  AOI22_X1 U22147 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10993), .ZN(n20000) );
  OAI21_X1 U22148 ( .B1(n20001), .B2(n20050), .A(n20000), .ZN(U241) );
  AOI22_X1 U22149 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10993), .ZN(n20002) );
  OAI21_X1 U22150 ( .B1(n14575), .B2(n20050), .A(n20002), .ZN(U240) );
  INV_X1 U22151 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U22152 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10993), .ZN(n20003) );
  OAI21_X1 U22153 ( .B1(n20004), .B2(n20050), .A(n20003), .ZN(U239) );
  INV_X1 U22154 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U22155 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10993), .ZN(n20005) );
  OAI21_X1 U22156 ( .B1(n20006), .B2(n20050), .A(n20005), .ZN(U238) );
  AOI22_X1 U22157 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10993), .ZN(n20007) );
  OAI21_X1 U22158 ( .B1(n20008), .B2(n20050), .A(n20007), .ZN(U237) );
  AOI22_X1 U22159 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10993), .ZN(n20009) );
  OAI21_X1 U22160 ( .B1(n20010), .B2(n20050), .A(n20009), .ZN(U236) );
  AOI22_X1 U22161 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10993), .ZN(n20011) );
  OAI21_X1 U22162 ( .B1(n20012), .B2(n20050), .A(n20011), .ZN(U235) );
  AOI22_X1 U22163 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10993), .ZN(n20013) );
  OAI21_X1 U22164 ( .B1(n20014), .B2(n20050), .A(n20013), .ZN(U234) );
  AOI22_X1 U22165 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10993), .ZN(n20015) );
  OAI21_X1 U22166 ( .B1(n20016), .B2(n20050), .A(n20015), .ZN(U233) );
  AOI22_X1 U22167 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10993), .ZN(n20017) );
  OAI21_X1 U22168 ( .B1(n14209), .B2(n20050), .A(n20017), .ZN(U232) );
  AOI22_X1 U22169 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10993), .ZN(n20018) );
  OAI21_X1 U22170 ( .B1(n20019), .B2(n20050), .A(n20018), .ZN(U231) );
  AOI22_X1 U22171 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10993), .ZN(n20020) );
  OAI21_X1 U22172 ( .B1(n20021), .B2(n20050), .A(n20020), .ZN(U230) );
  AOI22_X1 U22173 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10993), .ZN(n20022) );
  OAI21_X1 U22174 ( .B1(n20023), .B2(n20050), .A(n20022), .ZN(U229) );
  AOI22_X1 U22175 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10993), .ZN(n20024) );
  OAI21_X1 U22176 ( .B1(n20025), .B2(n20050), .A(n20024), .ZN(U228) );
  AOI22_X1 U22177 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10993), .ZN(n20026) );
  OAI21_X1 U22178 ( .B1(n20027), .B2(n20050), .A(n20026), .ZN(U227) );
  AOI22_X1 U22179 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10993), .ZN(n20028) );
  OAI21_X1 U22180 ( .B1(n20029), .B2(n20050), .A(n20028), .ZN(U226) );
  AOI22_X1 U22181 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10993), .ZN(n20030) );
  OAI21_X1 U22182 ( .B1(n20031), .B2(n20050), .A(n20030), .ZN(U225) );
  AOI22_X1 U22183 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10993), .ZN(n20032) );
  OAI21_X1 U22184 ( .B1(n20033), .B2(n20050), .A(n20032), .ZN(U224) );
  AOI22_X1 U22185 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10993), .ZN(n20034) );
  OAI21_X1 U22186 ( .B1(n20035), .B2(n20050), .A(n20034), .ZN(U223) );
  AOI22_X1 U22187 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10993), .ZN(n20036) );
  OAI21_X1 U22188 ( .B1(n20037), .B2(n20050), .A(n20036), .ZN(U222) );
  AOI22_X1 U22189 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10993), .ZN(n20039) );
  OAI21_X1 U22190 ( .B1(n20040), .B2(n20050), .A(n20039), .ZN(U221) );
  AOI22_X1 U22191 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10993), .ZN(n20041) );
  OAI21_X1 U22192 ( .B1(n20042), .B2(n20050), .A(n20041), .ZN(U220) );
  AOI22_X1 U22193 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10993), .ZN(n20043) );
  OAI21_X1 U22194 ( .B1(n20044), .B2(n20050), .A(n20043), .ZN(U219) );
  AOI22_X1 U22195 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10993), .ZN(n20045) );
  OAI21_X1 U22196 ( .B1(n20046), .B2(n20050), .A(n20045), .ZN(U218) );
  AOI22_X1 U22197 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20038), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10993), .ZN(n20047) );
  OAI21_X1 U22198 ( .B1(n14066), .B2(n20050), .A(n20047), .ZN(U217) );
  OAI222_X1 U22199 ( .A1(U212), .A2(n20051), .B1(n20050), .B2(n20049), .C1(
        U214), .C2(n20048), .ZN(U216) );
  AOI22_X1 U22200 ( .A1(n22339), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20052), 
        .B2(n22337), .ZN(P1_U3483) );
  OAI21_X1 U22201 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20796), .A(n20801), 
        .ZN(n20053) );
  AOI211_X1 U22202 ( .C1(n20054), .C2(n20053), .A(n21710), .B(n21144), .ZN(
        n20055) );
  OAI21_X1 U22203 ( .B1(n20055), .B2(n21277), .A(n21267), .ZN(n20060) );
  AOI21_X1 U22204 ( .B1(n21764), .B2(n18233), .A(n20116), .ZN(n20056) );
  INV_X1 U22205 ( .A(n20056), .ZN(n20057) );
  AOI21_X1 U22206 ( .B1(n20058), .B2(n21279), .A(n20057), .ZN(n20059) );
  MUX2_X1 U22207 ( .A(n20060), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20059), 
        .Z(P3_U3296) );
  AOI22_X1 U22208 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20080), .ZN(n20064) );
  OAI21_X1 U22209 ( .B1(n20065), .B2(n20112), .A(n20064), .ZN(P3_U2768) );
  AOI22_X1 U22210 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20080), .ZN(n20066) );
  OAI21_X1 U22211 ( .B1(n20067), .B2(n20112), .A(n20066), .ZN(P3_U2769) );
  AOI22_X1 U22212 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20080), .ZN(n20068) );
  OAI21_X1 U22213 ( .B1(n20069), .B2(n20112), .A(n20068), .ZN(P3_U2770) );
  AOI22_X1 U22214 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20080), .ZN(n20070) );
  OAI21_X1 U22215 ( .B1(n20631), .B2(n20112), .A(n20070), .ZN(P3_U2771) );
  AOI22_X1 U22216 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20080), .ZN(n20071) );
  OAI21_X1 U22217 ( .B1(n20072), .B2(n20112), .A(n20071), .ZN(P3_U2772) );
  AOI22_X1 U22218 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20080), .ZN(n20073) );
  OAI21_X1 U22219 ( .B1(n20647), .B2(n20112), .A(n20073), .ZN(P3_U2773) );
  AOI22_X1 U22220 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20080), .ZN(n20074) );
  OAI21_X1 U22221 ( .B1(n20648), .B2(n20112), .A(n20074), .ZN(P3_U2774) );
  AOI22_X1 U22222 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20080), .ZN(n20075) );
  OAI21_X1 U22223 ( .B1(n20076), .B2(n20112), .A(n20075), .ZN(P3_U2775) );
  AOI22_X1 U22224 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20080), .ZN(n20077) );
  OAI21_X1 U22225 ( .B1(n20078), .B2(n20112), .A(n20077), .ZN(P3_U2776) );
  AOI22_X1 U22226 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20080), .ZN(n20079) );
  OAI21_X1 U22227 ( .B1(n20650), .B2(n20112), .A(n20079), .ZN(P3_U2777) );
  AOI22_X1 U22228 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20109), .ZN(n20081) );
  OAI21_X1 U22229 ( .B1(n20082), .B2(n20112), .A(n20081), .ZN(P3_U2778) );
  AOI22_X1 U22230 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20109), .ZN(n20083) );
  OAI21_X1 U22231 ( .B1(n20681), .B2(n20112), .A(n20083), .ZN(P3_U2779) );
  AOI22_X1 U22232 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20110), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20109), .ZN(n20084) );
  OAI21_X1 U22233 ( .B1(n20085), .B2(n20112), .A(n20084), .ZN(P3_U2780) );
  AOI22_X1 U22234 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20098), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20109), .ZN(n20086) );
  OAI21_X1 U22235 ( .B1(n20669), .B2(n20112), .A(n20086), .ZN(P3_U2781) );
  AOI22_X1 U22236 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20098), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20109), .ZN(n20087) );
  OAI21_X1 U22237 ( .B1(n20667), .B2(n20112), .A(n20087), .ZN(P3_U2782) );
  AOI22_X1 U22238 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20109), .ZN(n20088) );
  OAI21_X1 U22239 ( .B1(n20728), .B2(n20112), .A(n20088), .ZN(P3_U2783) );
  AOI22_X1 U22240 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20109), .ZN(n20089) );
  OAI21_X1 U22241 ( .B1(n20586), .B2(n20112), .A(n20089), .ZN(P3_U2784) );
  AOI22_X1 U22242 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20109), .ZN(n20090) );
  OAI21_X1 U22243 ( .B1(n20091), .B2(n20112), .A(n20090), .ZN(P3_U2785) );
  AOI22_X1 U22244 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20109), .ZN(n20092) );
  OAI21_X1 U22245 ( .B1(n20093), .B2(n20112), .A(n20092), .ZN(P3_U2786) );
  AOI22_X1 U22246 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20109), .ZN(n20094) );
  OAI21_X1 U22247 ( .B1(n20587), .B2(n20112), .A(n20094), .ZN(P3_U2787) );
  AOI22_X1 U22248 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20109), .ZN(n20095) );
  OAI21_X1 U22249 ( .B1(n20096), .B2(n20112), .A(n20095), .ZN(P3_U2788) );
  AOI22_X1 U22250 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20109), .ZN(n20097) );
  OAI21_X1 U22251 ( .B1(n20588), .B2(n20112), .A(n20097), .ZN(P3_U2789) );
  AOI22_X1 U22252 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20098), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20109), .ZN(n20099) );
  OAI21_X1 U22253 ( .B1(n20100), .B2(n20112), .A(n20099), .ZN(P3_U2790) );
  AOI22_X1 U22254 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20109), .ZN(n20101) );
  OAI21_X1 U22255 ( .B1(n20721), .B2(n20112), .A(n20101), .ZN(P3_U2791) );
  AOI22_X1 U22256 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20109), .ZN(n20102) );
  OAI21_X1 U22257 ( .B1(n20562), .B2(n20112), .A(n20102), .ZN(P3_U2792) );
  AOI22_X1 U22258 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20109), .ZN(n20103) );
  OAI21_X1 U22259 ( .B1(n20555), .B2(n20112), .A(n20103), .ZN(P3_U2793) );
  AOI22_X1 U22260 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20109), .ZN(n20104) );
  OAI21_X1 U22261 ( .B1(n20563), .B2(n20112), .A(n20104), .ZN(P3_U2794) );
  AOI22_X1 U22262 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20109), .ZN(n20105) );
  OAI21_X1 U22263 ( .B1(n20556), .B2(n20112), .A(n20105), .ZN(P3_U2795) );
  AOI22_X1 U22264 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20109), .ZN(n20106) );
  OAI21_X1 U22265 ( .B1(n20107), .B2(n20112), .A(n20106), .ZN(P3_U2796) );
  AOI22_X1 U22266 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20109), .ZN(n20108) );
  OAI21_X1 U22267 ( .B1(n20711), .B2(n20112), .A(n20108), .ZN(P3_U2797) );
  AOI22_X1 U22268 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20110), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20109), .ZN(n20111) );
  OAI21_X1 U22269 ( .B1(n20717), .B2(n20112), .A(n20111), .ZN(P3_U2798) );
  NAND2_X1 U22270 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20796), .ZN(n20114) );
  AOI211_X4 U22271 ( .C1(n21764), .C2(n21703), .A(n20118), .B(n20114), .ZN(
        n20504) );
  NAND4_X1 U22272 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21277), .A3(n21144), 
        .A4(n21703), .ZN(n21261) );
  INV_X1 U22273 ( .A(n21261), .ZN(n20368) );
  NAND2_X1 U22274 ( .A1(n21199), .A2(n20525), .ZN(n20115) );
  INV_X1 U22275 ( .A(n20775), .ZN(n20769) );
  NAND2_X1 U22276 ( .A1(n20117), .A2(n20769), .ZN(n20748) );
  INV_X1 U22277 ( .A(n20748), .ZN(n20751) );
  AOI22_X1 U22278 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20340), .B1(n20751), 
        .B2(n20171), .ZN(n20123) );
  INV_X1 U22279 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20335) );
  NAND2_X1 U22280 ( .A1(n20354), .A2(n20368), .ZN(n20131) );
  OAI21_X1 U22281 ( .B1(n20335), .B2(n20131), .A(n20479), .ZN(n20121) );
  AOI21_X1 U22282 ( .B1(n20354), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n20525), .ZN(n20289) );
  OAI211_X1 U22283 ( .C1(n20801), .C2(n20796), .A(n21764), .B(n21703), .ZN(
        n21258) );
  INV_X1 U22284 ( .A(n21258), .ZN(n20119) );
  AOI211_X4 U22285 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20796), .A(n20119), .B(
        n20118), .ZN(n20522) );
  OAI22_X1 U22286 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20463), .B1(n20544), 
        .B2(n20125), .ZN(n20120) );
  AOI221_X1 U22287 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20121), .C1(
        n20130), .C2(n20289), .A(n20120), .ZN(n20122) );
  OAI211_X1 U22288 ( .C1(n20543), .C2(n20124), .A(n20123), .B(n20122), .ZN(
        P3_U2670) );
  INV_X1 U22289 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20141) );
  NAND2_X1 U22290 ( .A1(n20126), .A2(n20125), .ZN(n20127) );
  NOR3_X1 U22291 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20154) );
  AOI211_X1 U22292 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20127), .A(n20154), .B(
        n20543), .ZN(n20138) );
  OAI21_X1 U22293 ( .B1(n21240), .B2(n20775), .A(n20764), .ZN(n20128) );
  INV_X1 U22294 ( .A(n20128), .ZN(n20762) );
  NOR2_X1 U22295 ( .A1(n20354), .A2(n20525), .ZN(n20309) );
  AOI22_X1 U22296 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n20340), .B1(n20129), 
        .B2(n20309), .ZN(n20136) );
  NOR2_X1 U22297 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20130), .ZN(
        n20168) );
  INV_X1 U22298 ( .A(n20131), .ZN(n20133) );
  NAND2_X1 U22299 ( .A1(n20146), .A2(n20335), .ZN(n20132) );
  OAI211_X1 U22300 ( .C1(n20168), .C2(n20134), .A(n20133), .B(n20132), .ZN(
        n20135) );
  OAI211_X1 U22301 ( .C1(n20762), .C2(n20550), .A(n20136), .B(n20135), .ZN(
        n20137) );
  AOI211_X1 U22302 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20138), .B(n20137), .ZN(n20140) );
  NAND2_X1 U22303 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20144) );
  OAI211_X1 U22304 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20363), .B(n20144), .ZN(n20139) );
  OAI211_X1 U22305 ( .C1(n20141), .C2(n20544), .A(n20140), .B(n20139), .ZN(
        P3_U2669) );
  INV_X1 U22306 ( .A(n20758), .ZN(n20780) );
  OAI21_X1 U22307 ( .B1(n20772), .B2(n20780), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20783) );
  NAND2_X1 U22308 ( .A1(n20783), .A2(n20142), .ZN(n20791) );
  NOR2_X1 U22309 ( .A1(n20150), .A2(n20144), .ZN(n20178) );
  NOR2_X1 U22310 ( .A1(n20463), .A2(n20178), .ZN(n20145) );
  INV_X1 U22311 ( .A(n20145), .ZN(n20143) );
  OAI22_X1 U22312 ( .A1(n20544), .A2(n20153), .B1(n20144), .B2(n20143), .ZN(
        n20152) );
  NOR2_X1 U22313 ( .A1(n20340), .A2(n20145), .ZN(n20163) );
  AOI21_X1 U22314 ( .B1(n20335), .B2(n20146), .A(n20528), .ZN(n20147) );
  XOR2_X1 U22315 ( .A(n20148), .B(n20147), .Z(n20149) );
  OAI22_X1 U22316 ( .A1(n20163), .A2(n20150), .B1(n21261), .B2(n20149), .ZN(
        n20151) );
  AOI211_X1 U22317 ( .C1(n20171), .C2(n20791), .A(n20152), .B(n20151), .ZN(
        n20156) );
  NAND2_X1 U22318 ( .A1(n20154), .A2(n20153), .ZN(n20158) );
  OAI211_X1 U22319 ( .C1(n20154), .C2(n20153), .A(n20504), .B(n20158), .ZN(
        n20155) );
  OAI211_X1 U22320 ( .C1(n20479), .C2(n20157), .A(n20156), .B(n20155), .ZN(
        P3_U2668) );
  AND3_X1 U22321 ( .A1(n20162), .A2(n20363), .A3(n20178), .ZN(n20167) );
  NOR2_X1 U22322 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20158), .ZN(n20182) );
  AOI211_X1 U22323 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20158), .A(n20182), .B(
        n20543), .ZN(n20166) );
  AOI22_X1 U22324 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n20159) );
  INV_X1 U22325 ( .A(n20159), .ZN(n20165) );
  NOR2_X1 U22326 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20525), .ZN(
        n20307) );
  AOI21_X1 U22327 ( .B1(n20160), .B2(n20307), .A(n20309), .ZN(n20161) );
  OAI22_X1 U22328 ( .A1(n20163), .A2(n20162), .B1(n20161), .B2(n20170), .ZN(
        n20164) );
  NOR4_X1 U22329 ( .A1(n20167), .A2(n20166), .A3(n20165), .A4(n20164), .ZN(
        n20175) );
  AOI21_X1 U22330 ( .B1(n20169), .B2(n20168), .A(n20528), .ZN(n20177) );
  NAND3_X1 U22331 ( .A1(n20368), .A2(n20177), .A3(n20170), .ZN(n20174) );
  OAI21_X1 U22332 ( .B1(n20172), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20171), .ZN(n20173) );
  NAND4_X1 U22333 ( .A1(n20175), .A2(n21199), .A3(n20174), .A4(n20173), .ZN(
        P3_U2667) );
  XNOR2_X1 U22334 ( .A(n20177), .B(n20176), .ZN(n20189) );
  NAND2_X1 U22335 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20178), .ZN(n20185) );
  NOR2_X1 U22336 ( .A1(n20179), .A2(n20185), .ZN(n20201) );
  OAI21_X1 U22337 ( .B1(n20201), .B2(n20463), .A(n20547), .ZN(n20207) );
  OAI22_X1 U22338 ( .A1(n20180), .A2(n20479), .B1(n20544), .B2(n20181), .ZN(
        n20187) );
  INV_X1 U22339 ( .A(n20201), .ZN(n20190) );
  NAND2_X1 U22340 ( .A1(n20363), .A2(n20190), .ZN(n20184) );
  NAND2_X1 U22341 ( .A1(n20182), .A2(n20181), .ZN(n20194) );
  OAI211_X1 U22342 ( .C1(n20182), .C2(n20181), .A(n20504), .B(n20194), .ZN(
        n20183) );
  OAI211_X1 U22343 ( .C1(n20185), .C2(n20184), .A(n21199), .B(n20183), .ZN(
        n20186) );
  AOI211_X1 U22344 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n20207), .A(n20187), .B(
        n20186), .ZN(n20188) );
  OAI21_X1 U22345 ( .B1(n21261), .B2(n20189), .A(n20188), .ZN(P3_U2666) );
  OAI21_X1 U22346 ( .B1(n11019), .B2(n11167), .A(n20289), .ZN(n20199) );
  NOR3_X1 U22347 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20463), .A3(n20190), .ZN(
        n20208) );
  OAI21_X1 U22348 ( .B1(n11167), .B2(n20479), .A(n21199), .ZN(n20191) );
  AOI211_X1 U22349 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20522), .A(n20208), .B(
        n20191), .ZN(n20198) );
  INV_X1 U22350 ( .A(n20200), .ZN(n20193) );
  OAI21_X1 U22351 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20192), .A(
        n20354), .ZN(n20202) );
  NOR3_X1 U22352 ( .A1(n20193), .A2(n20525), .A3(n20202), .ZN(n20196) );
  AOI211_X1 U22353 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20194), .A(n20210), .B(
        n20543), .ZN(n20195) );
  AOI211_X1 U22354 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n20207), .A(n20196), .B(
        n20195), .ZN(n20197) );
  OAI211_X1 U22355 ( .C1(n20200), .C2(n20199), .A(n20198), .B(n20197), .ZN(
        P3_U2665) );
  NAND2_X1 U22356 ( .A1(n20363), .A2(n20898), .ZN(n20213) );
  NAND2_X1 U22357 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20201), .ZN(n20215) );
  XOR2_X1 U22358 ( .A(n20203), .B(n20202), .Z(n20205) );
  AOI22_X1 U22359 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n20204) );
  OAI211_X1 U22360 ( .C1(n21261), .C2(n20205), .A(n20204), .B(n21199), .ZN(
        n20206) );
  AOI221_X1 U22361 ( .B1(n20208), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n20207), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n20206), .ZN(n20212) );
  INV_X1 U22362 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U22363 ( .A1(n20210), .A2(n20209), .ZN(n20214) );
  OAI211_X1 U22364 ( .C1(n20210), .C2(n20209), .A(n20504), .B(n20214), .ZN(
        n20211) );
  OAI211_X1 U22365 ( .C1(n20213), .C2(n20215), .A(n20212), .B(n20211), .ZN(
        P3_U2664) );
  AOI211_X1 U22366 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20214), .A(n20240), .B(
        n20543), .ZN(n20223) );
  NOR2_X1 U22367 ( .A1(n20898), .A2(n20215), .ZN(n20216) );
  NAND2_X1 U22368 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20216), .ZN(n20244) );
  AOI21_X1 U22369 ( .B1(n20244), .B2(n20363), .A(n20340), .ZN(n20227) );
  AOI21_X1 U22370 ( .B1(n20363), .B2(n20216), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n20221) );
  AOI21_X1 U22371 ( .B1(n20217), .B2(n20335), .A(n20528), .ZN(n20219) );
  XOR2_X1 U22372 ( .A(n20219), .B(n20218), .Z(n20220) );
  OAI22_X1 U22373 ( .A1(n20227), .A2(n20221), .B1(n21261), .B2(n20220), .ZN(
        n20222) );
  AOI211_X1 U22374 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20223), .B(n20222), .ZN(n20224) );
  OAI211_X1 U22375 ( .C1(n20544), .C2(n20225), .A(n20224), .B(n21199), .ZN(
        P3_U2663) );
  AOI21_X1 U22376 ( .B1(n20504), .B2(n20240), .A(n20522), .ZN(n20236) );
  NOR2_X1 U22377 ( .A1(n20240), .A2(n20543), .ZN(n20226) );
  NOR3_X1 U22378 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20463), .A3(n20244), .ZN(
        n20243) );
  AOI211_X1 U22379 ( .C1(n20226), .C2(n20239), .A(n10990), .B(n20243), .ZN(
        n20235) );
  INV_X1 U22380 ( .A(n20227), .ZN(n20242) );
  AOI21_X1 U22381 ( .B1(n20335), .B2(n20228), .A(n20528), .ZN(n20237) );
  AND3_X1 U22382 ( .A1(n20230), .A2(n20368), .A3(n20237), .ZN(n20233) );
  AOI21_X1 U22383 ( .B1(n20307), .B2(n20229), .A(n20309), .ZN(n20231) );
  OAI22_X1 U22384 ( .A1(n20231), .A2(n20230), .B1(n20229), .B2(n20479), .ZN(
        n20232) );
  AOI211_X1 U22385 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n20242), .A(n20233), .B(
        n20232), .ZN(n20234) );
  OAI211_X1 U22386 ( .C1(n20239), .C2(n20236), .A(n20235), .B(n20234), .ZN(
        P3_U2662) );
  XOR2_X1 U22387 ( .A(n20238), .B(n20237), .Z(n20253) );
  NAND2_X1 U22388 ( .A1(n20240), .A2(n20239), .ZN(n20241) );
  AOI211_X1 U22389 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20241), .A(n20260), .B(
        n20543), .ZN(n20251) );
  OAI21_X1 U22390 ( .B1(n20243), .B2(n20242), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20248) );
  NOR2_X1 U22391 ( .A1(n20245), .A2(n20244), .ZN(n20257) );
  NAND3_X1 U22392 ( .A1(n20363), .A2(n20257), .A3(n20246), .ZN(n20247) );
  OAI211_X1 U22393 ( .C1(n20249), .C2(n20544), .A(n20248), .B(n20247), .ZN(
        n20250) );
  AOI211_X1 U22394 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20251), .B(n20250), .ZN(n20252) );
  OAI211_X1 U22395 ( .C1(n20253), .C2(n21261), .A(n20252), .B(n21199), .ZN(
        P3_U2661) );
  AOI21_X1 U22396 ( .B1(n20254), .B2(n20335), .A(n20528), .ZN(n20255) );
  XOR2_X1 U22397 ( .A(n20256), .B(n20255), .Z(n20266) );
  NAND2_X1 U22398 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20257), .ZN(n20277) );
  NOR2_X1 U22399 ( .A1(n20463), .A2(n20277), .ZN(n20258) );
  NOR2_X1 U22400 ( .A1(n20278), .A2(n20277), .ZN(n20297) );
  OAI21_X1 U22401 ( .B1(n20297), .B2(n20463), .A(n20547), .ZN(n20287) );
  OAI21_X1 U22402 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n20258), .A(n20287), 
        .ZN(n20262) );
  INV_X1 U22403 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20259) );
  NAND2_X1 U22404 ( .A1(n20260), .A2(n20259), .ZN(n20267) );
  OAI211_X1 U22405 ( .C1(n20260), .C2(n20259), .A(n20504), .B(n20267), .ZN(
        n20261) );
  OAI211_X1 U22406 ( .C1(n20479), .C2(n20263), .A(n20262), .B(n20261), .ZN(
        n20264) );
  AOI211_X1 U22407 ( .C1(n20522), .C2(P3_EBX_REG_11__SCAN_IN), .A(n10990), .B(
        n20264), .ZN(n20265) );
  OAI21_X1 U22408 ( .B1(n21261), .B2(n20266), .A(n20265), .ZN(P3_U2660) );
  AOI211_X1 U22409 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20267), .A(n20283), .B(
        n20543), .ZN(n20268) );
  AOI211_X1 U22410 ( .C1(n20522), .C2(P3_EBX_REG_12__SCAN_IN), .A(n10990), .B(
        n20268), .ZN(n20275) );
  NOR4_X1 U22411 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20463), .A3(n20278), 
        .A4(n20277), .ZN(n20288) );
  OAI21_X1 U22412 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20269), .A(
        n20354), .ZN(n20271) );
  OAI21_X1 U22413 ( .B1(n20272), .B2(n20271), .A(n20368), .ZN(n20270) );
  AOI21_X1 U22414 ( .B1(n20272), .B2(n20271), .A(n20270), .ZN(n20273) );
  AOI211_X1 U22415 ( .C1(P3_REIP_REG_12__SCAN_IN), .C2(n20287), .A(n20288), 
        .B(n20273), .ZN(n20274) );
  OAI211_X1 U22416 ( .C1(n20276), .C2(n20479), .A(n20275), .B(n20274), .ZN(
        P3_U2659) );
  NOR3_X1 U22417 ( .A1(n20463), .A2(n20278), .A3(n20277), .ZN(n20279) );
  NAND2_X1 U22418 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20279), .ZN(n20295) );
  OAI21_X1 U22419 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20280), .A(
        n20354), .ZN(n20298) );
  NOR3_X1 U22420 ( .A1(n20290), .A2(n20525), .A3(n20298), .ZN(n20281) );
  AOI211_X1 U22421 ( .C1(n20522), .C2(P3_EBX_REG_13__SCAN_IN), .A(n10990), .B(
        n20281), .ZN(n20285) );
  NAND2_X1 U22422 ( .A1(n20283), .A2(n20282), .ZN(n20294) );
  OAI211_X1 U22423 ( .C1(n20283), .C2(n20282), .A(n20504), .B(n20294), .ZN(
        n20284) );
  OAI211_X1 U22424 ( .C1(n20479), .C2(n20291), .A(n20285), .B(n20284), .ZN(
        n20286) );
  AOI221_X1 U22425 ( .B1(n20288), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n20287), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n20286), .ZN(n20293) );
  OAI211_X1 U22426 ( .C1(n20309), .C2(n20291), .A(n20290), .B(n20289), .ZN(
        n20292) );
  OAI211_X1 U22427 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n20295), .A(n20293), 
        .B(n20292), .ZN(P3_U2658) );
  AOI211_X1 U22428 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20294), .A(n20317), .B(
        n20543), .ZN(n20303) );
  INV_X1 U22429 ( .A(n20295), .ZN(n20296) );
  AOI21_X1 U22430 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n20296), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n20301) );
  NAND4_X1 U22431 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .A3(P3_REIP_REG_12__SCAN_IN), .A4(n20297), .ZN(n20321) );
  AOI21_X1 U22432 ( .B1(n20363), .B2(n20321), .A(n20340), .ZN(n20306) );
  XOR2_X1 U22433 ( .A(n20299), .B(n20298), .Z(n20300) );
  OAI22_X1 U22434 ( .A1(n20301), .A2(n20306), .B1(n21261), .B2(n20300), .ZN(
        n20302) );
  AOI211_X1 U22435 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20303), .B(n20302), .ZN(n20304) );
  OAI211_X1 U22436 ( .C1(n20544), .C2(n20305), .A(n20304), .B(n21199), .ZN(
        P3_U2657) );
  INV_X1 U22437 ( .A(n20306), .ZN(n20327) );
  AOI22_X1 U22438 ( .A1(n20368), .A2(n20311), .B1(n20308), .B2(n20307), .ZN(
        n20312) );
  INV_X1 U22439 ( .A(n20309), .ZN(n20357) );
  NOR2_X1 U22440 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20310), .ZN(
        n20382) );
  NOR2_X1 U22441 ( .A1(n20382), .A2(n20528), .ZN(n20352) );
  INV_X1 U22442 ( .A(n20352), .ZN(n20328) );
  AOI22_X1 U22443 ( .A1(n20312), .A2(n20357), .B1(n20311), .B2(n20328), .ZN(
        n20315) );
  OAI22_X1 U22444 ( .A1(n20313), .A2(n20479), .B1(n20544), .B2(n20316), .ZN(
        n20314) );
  AOI211_X1 U22445 ( .C1(n20327), .C2(P3_REIP_REG_15__SCAN_IN), .A(n20315), 
        .B(n20314), .ZN(n20320) );
  NOR3_X1 U22446 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20463), .A3(n20321), 
        .ZN(n20326) );
  INV_X1 U22447 ( .A(n20326), .ZN(n20319) );
  NAND2_X1 U22448 ( .A1(n20317), .A2(n20316), .ZN(n20323) );
  OAI211_X1 U22449 ( .C1(n20317), .C2(n20316), .A(n20504), .B(n20323), .ZN(
        n20318) );
  NAND4_X1 U22450 ( .A1(n20320), .A2(n21199), .A3(n20319), .A4(n20318), .ZN(
        P3_U2656) );
  AOI22_X1 U22451 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n20334) );
  NOR2_X1 U22452 ( .A1(n20322), .A2(n20321), .ZN(n20339) );
  NOR2_X1 U22453 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20463), .ZN(n20325) );
  AOI211_X1 U22454 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20323), .A(n20348), .B(
        n20543), .ZN(n20324) );
  AOI211_X1 U22455 ( .C1(n20339), .C2(n20325), .A(n10990), .B(n20324), .ZN(
        n20333) );
  OAI21_X1 U22456 ( .B1(n20327), .B2(n20326), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n20332) );
  INV_X1 U22457 ( .A(n20330), .ZN(n20329) );
  OAI221_X1 U22458 ( .B1(n20330), .B2(n20352), .C1(n20329), .C2(n20328), .A(
        n20368), .ZN(n20331) );
  NAND4_X1 U22459 ( .A1(n20334), .A2(n20333), .A3(n20332), .A4(n20331), .ZN(
        P3_U2655) );
  INV_X1 U22460 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20351) );
  AOI21_X1 U22461 ( .B1(n20336), .B2(n20335), .A(n20528), .ZN(n20337) );
  XNOR2_X1 U22462 ( .A(n20338), .B(n20337), .ZN(n20347) );
  NAND2_X1 U22463 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20339), .ZN(n20341) );
  NOR2_X1 U22464 ( .A1(n20345), .A2(n20341), .ZN(n20362) );
  NOR2_X1 U22465 ( .A1(n20362), .A2(n20463), .ZN(n20342) );
  NOR2_X1 U22466 ( .A1(n20340), .A2(n20342), .ZN(n20421) );
  INV_X1 U22467 ( .A(n20341), .ZN(n20343) );
  AOI22_X1 U22468 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20523), .B1(
        n20343), .B2(n20342), .ZN(n20344) );
  OAI211_X1 U22469 ( .C1(n20421), .C2(n20345), .A(n20344), .B(n21199), .ZN(
        n20346) );
  AOI21_X1 U22470 ( .B1(n20347), .B2(n20368), .A(n20346), .ZN(n20350) );
  NAND2_X1 U22471 ( .A1(n20348), .A2(n20351), .ZN(n20359) );
  OAI211_X1 U22472 ( .C1(n20348), .C2(n20351), .A(n20504), .B(n20359), .ZN(
        n20349) );
  OAI211_X1 U22473 ( .C1(n20351), .C2(n20544), .A(n20350), .B(n20349), .ZN(
        P3_U2654) );
  AOI21_X1 U22474 ( .B1(n20354), .B2(n20353), .A(n20352), .ZN(n20371) );
  OAI221_X1 U22475 ( .B1(n20358), .B2(n20382), .C1(n20358), .C2(n20355), .A(
        n20368), .ZN(n20356) );
  AOI22_X1 U22476 ( .A1(n20371), .A2(n20358), .B1(n20357), .B2(n20356), .ZN(
        n20361) );
  AOI211_X1 U22477 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20359), .A(n20377), .B(
        n20543), .ZN(n20360) );
  AOI211_X1 U22478 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20361), .B(n20360), .ZN(n20367) );
  INV_X1 U22479 ( .A(n20421), .ZN(n20375) );
  OAI22_X1 U22480 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20428), .B1(n20544), 
        .B2(n20364), .ZN(n20365) );
  AOI211_X1 U22481 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n20375), .A(n10990), 
        .B(n20365), .ZN(n20366) );
  NAND2_X1 U22482 ( .A1(n20367), .A2(n20366), .ZN(P3_U2653) );
  OAI21_X1 U22483 ( .B1(n20371), .B2(n20370), .A(n20368), .ZN(n20369) );
  AOI21_X1 U22484 ( .B1(n20371), .B2(n20370), .A(n20369), .ZN(n20374) );
  INV_X1 U22485 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20376) );
  NAND2_X1 U22486 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20387) );
  OAI211_X1 U22487 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n20438), .B(n20387), .ZN(n20372) );
  OAI211_X1 U22488 ( .C1(n20544), .C2(n20376), .A(n21199), .B(n20372), .ZN(
        n20373) );
  AOI211_X1 U22489 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n20375), .A(n20374), 
        .B(n20373), .ZN(n20379) );
  NAND2_X1 U22490 ( .A1(n20377), .A2(n20376), .ZN(n20380) );
  OAI211_X1 U22491 ( .C1(n20377), .C2(n20376), .A(n20504), .B(n20380), .ZN(
        n20378) );
  OAI211_X1 U22492 ( .C1(n20479), .C2(n11157), .A(n20379), .B(n20378), .ZN(
        P3_U2652) );
  NOR2_X1 U22493 ( .A1(n21150), .A2(n20387), .ZN(n20410) );
  OAI21_X1 U22494 ( .B1(n20410), .B2(n20463), .A(n20421), .ZN(n20414) );
  INV_X1 U22495 ( .A(n20414), .ZN(n20392) );
  AOI211_X1 U22496 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20380), .A(n20401), .B(
        n20543), .ZN(n20381) );
  AOI21_X1 U22497 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n20522), .A(n20381), .ZN(
        n20391) );
  AOI211_X1 U22498 ( .C1(n20386), .C2(n20385), .A(n20394), .B(n21261), .ZN(
        n20389) );
  NOR3_X1 U22499 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20387), .A3(n20428), 
        .ZN(n20388) );
  AOI211_X1 U22500 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n20389), .B(n20388), .ZN(n20390) );
  OAI211_X1 U22501 ( .C1(n20392), .C2(n21150), .A(n20391), .B(n20390), .ZN(
        P3_U2651) );
  AOI211_X1 U22502 ( .C1(n20396), .C2(n20395), .A(n20407), .B(n21261), .ZN(
        n20400) );
  INV_X1 U22503 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20397) );
  NAND3_X1 U22504 ( .A1(n20397), .A2(n20410), .A3(n20438), .ZN(n20413) );
  OAI21_X1 U22505 ( .B1(n20479), .B2(n20398), .A(n20413), .ZN(n20399) );
  AOI211_X1 U22506 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n20414), .A(n20400), 
        .B(n20399), .ZN(n20403) );
  NAND2_X1 U22507 ( .A1(n20401), .A2(n20404), .ZN(n20405) );
  OAI211_X1 U22508 ( .C1(n20401), .C2(n20404), .A(n20504), .B(n20405), .ZN(
        n20402) );
  OAI211_X1 U22509 ( .C1(n20404), .C2(n20544), .A(n20403), .B(n20402), .ZN(
        P3_U2650) );
  AOI211_X1 U22510 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20405), .A(n20432), .B(
        n20543), .ZN(n20406) );
  AOI21_X1 U22511 ( .B1(n20523), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n20406), .ZN(n20418) );
  NOR2_X1 U22512 ( .A1(n20409), .A2(n20408), .ZN(n20422) );
  AOI211_X1 U22513 ( .C1(n20409), .C2(n20408), .A(n20422), .B(n21261), .ZN(
        n20412) );
  NAND2_X1 U22514 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20410), .ZN(n20419) );
  NOR3_X1 U22515 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20419), .A3(n20428), 
        .ZN(n20411) );
  AOI211_X1 U22516 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20522), .A(n20412), .B(
        n20411), .ZN(n20417) );
  INV_X1 U22517 ( .A(n20413), .ZN(n20415) );
  OAI21_X1 U22518 ( .B1(n20415), .B2(n20414), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n20416) );
  NAND3_X1 U22519 ( .A1(n20418), .A2(n20417), .A3(n20416), .ZN(P3_U2649) );
  NOR2_X1 U22520 ( .A1(n20420), .A2(n20419), .ZN(n20426) );
  AND2_X1 U22521 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20426), .ZN(n20439) );
  OAI21_X1 U22522 ( .B1(n20439), .B2(n20463), .A(n20421), .ZN(n20449) );
  NOR2_X1 U22523 ( .A1(n20422), .A2(n20528), .ZN(n20424) );
  NOR2_X1 U22524 ( .A1(n20424), .A2(n20423), .ZN(n20440) );
  AOI211_X1 U22525 ( .C1(n20424), .C2(n20423), .A(n20440), .B(n21261), .ZN(
        n20431) );
  NAND2_X1 U22526 ( .A1(n20426), .A2(n20425), .ZN(n20427) );
  OAI22_X1 U22527 ( .A1(n20429), .A2(n20479), .B1(n20428), .B2(n20427), .ZN(
        n20430) );
  AOI211_X1 U22528 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n20449), .A(n20431), 
        .B(n20430), .ZN(n20434) );
  NAND2_X1 U22529 ( .A1(n20432), .A2(n20435), .ZN(n20436) );
  OAI211_X1 U22530 ( .C1(n20432), .C2(n20435), .A(n20504), .B(n20436), .ZN(
        n20433) );
  OAI211_X1 U22531 ( .C1(n20435), .C2(n20544), .A(n20434), .B(n20433), .ZN(
        P3_U2648) );
  NOR2_X1 U22532 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20436), .ZN(n20455) );
  AOI211_X1 U22533 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20436), .A(n20455), .B(
        n20543), .ZN(n20437) );
  AOI21_X1 U22534 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n20522), .A(n20437), .ZN(
        n20445) );
  NAND2_X1 U22535 ( .A1(n20439), .A2(n20438), .ZN(n20447) );
  NOR2_X1 U22536 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20447), .ZN(n20450) );
  NOR2_X1 U22537 ( .A1(n20440), .A2(n20528), .ZN(n20441) );
  NOR2_X1 U22538 ( .A1(n20442), .A2(n20441), .ZN(n20452) );
  AOI211_X1 U22539 ( .C1(n20442), .C2(n20441), .A(n20452), .B(n20525), .ZN(
        n20443) );
  AOI211_X1 U22540 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n20449), .A(n20450), 
        .B(n20443), .ZN(n20444) );
  OAI211_X1 U22541 ( .C1(n20446), .C2(n20479), .A(n20445), .B(n20444), .ZN(
        P3_U2647) );
  INV_X1 U22542 ( .A(n20447), .ZN(n20448) );
  NAND2_X1 U22543 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20448), .ZN(n20475) );
  NOR2_X1 U22544 ( .A1(n20450), .A2(n20449), .ZN(n20464) );
  INV_X1 U22545 ( .A(n20451), .ZN(n20454) );
  AOI211_X1 U22546 ( .C1(n20454), .C2(n20453), .A(n11042), .B(n20525), .ZN(
        n20459) );
  NAND2_X1 U22547 ( .A1(n20455), .A2(n20457), .ZN(n20461) );
  OAI211_X1 U22548 ( .C1(n20455), .C2(n20457), .A(n20504), .B(n20461), .ZN(
        n20456) );
  OAI21_X1 U22549 ( .B1(n20457), .B2(n20544), .A(n20456), .ZN(n20458) );
  AOI211_X1 U22550 ( .C1(n20523), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20459), .B(n20458), .ZN(n20460) );
  OAI221_X1 U22551 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n20475), .C1(n20466), 
        .C2(n20464), .A(n20460), .ZN(P3_U2646) );
  NOR2_X1 U22552 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20461), .ZN(n20484) );
  AOI211_X1 U22553 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20461), .A(n20484), .B(
        n20543), .ZN(n20462) );
  AOI21_X1 U22554 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n20522), .A(n20462), .ZN(
        n20472) );
  NAND2_X1 U22555 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n20474) );
  NAND2_X1 U22556 ( .A1(n20463), .A2(n20547), .ZN(n20545) );
  INV_X1 U22557 ( .A(n20464), .ZN(n20465) );
  AOI21_X1 U22558 ( .B1(n20474), .B2(n20545), .A(n20465), .ZN(n20488) );
  INV_X1 U22559 ( .A(n20488), .ZN(n20502) );
  NOR3_X1 U22560 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n20466), .A3(n20475), 
        .ZN(n20470) );
  AOI211_X1 U22561 ( .C1(n20468), .C2(n20467), .A(n20476), .B(n21261), .ZN(
        n20469) );
  AOI211_X1 U22562 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n20502), .A(n20470), 
        .B(n20469), .ZN(n20471) );
  OAI211_X1 U22563 ( .C1(n20473), .C2(n20479), .A(n20472), .B(n20471), .ZN(
        P3_U2645) );
  AND2_X1 U22564 ( .A1(n20487), .A2(n20514), .ZN(n20493) );
  NOR2_X1 U22565 ( .A1(n20476), .A2(n20528), .ZN(n20477) );
  NOR2_X1 U22566 ( .A1(n20478), .A2(n20477), .ZN(n20489) );
  AOI211_X1 U22567 ( .C1(n20478), .C2(n20477), .A(n20489), .B(n20525), .ZN(
        n20482) );
  INV_X1 U22568 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20483) );
  OAI22_X1 U22569 ( .A1(n20480), .A2(n20479), .B1(n20544), .B2(n20483), .ZN(
        n20481) );
  NOR3_X1 U22570 ( .A1(n20493), .A2(n20482), .A3(n20481), .ZN(n20486) );
  NAND2_X1 U22571 ( .A1(n20484), .A2(n20483), .ZN(n20494) );
  OAI211_X1 U22572 ( .C1(n20484), .C2(n20483), .A(n20504), .B(n20494), .ZN(
        n20485) );
  OAI211_X1 U22573 ( .C1(n20488), .C2(n20487), .A(n20486), .B(n20485), .ZN(
        P3_U2644) );
  AOI22_X1 U22574 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20501) );
  NOR2_X1 U22575 ( .A1(n20489), .A2(n20528), .ZN(n20490) );
  NOR2_X1 U22576 ( .A1(n20491), .A2(n20490), .ZN(n20506) );
  AOI211_X1 U22577 ( .C1(n20491), .C2(n20490), .A(n20506), .B(n20525), .ZN(
        n20492) );
  AOI221_X1 U22578 ( .B1(n20493), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n20502), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n20492), .ZN(n20500) );
  INV_X1 U22579 ( .A(n20494), .ZN(n20496) );
  NAND2_X1 U22580 ( .A1(n20495), .A2(n20496), .ZN(n20505) );
  OAI211_X1 U22581 ( .C1(n20496), .C2(n20495), .A(n20504), .B(n20505), .ZN(
        n20499) );
  NAND3_X1 U22582 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20514), .A3(n20497), 
        .ZN(n20498) );
  NAND4_X1 U22583 ( .A1(n20501), .A2(n20500), .A3(n20499), .A4(n20498), .ZN(
        P3_U2643) );
  NAND3_X1 U22584 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n20514), .ZN(n20512) );
  AOI22_X1 U22585 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20523), .B1(
        n20522), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n20511) );
  NAND3_X1 U22586 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n20503) );
  AOI21_X1 U22587 ( .B1(n20503), .B2(n20545), .A(n20502), .ZN(n20532) );
  INV_X1 U22588 ( .A(n20532), .ZN(n20510) );
  NAND2_X1 U22589 ( .A1(n20504), .A2(n20518), .ZN(n20516) );
  AOI21_X1 U22590 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n20505), .A(n20516), .ZN(
        n20509) );
  NOR2_X1 U22591 ( .A1(n20506), .A2(n20528), .ZN(n20507) );
  NOR2_X1 U22592 ( .A1(n20513), .A2(n11019), .ZN(n20524) );
  XNOR2_X1 U22593 ( .A(n20526), .B(n20524), .ZN(n20521) );
  NAND4_X1 U22594 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n20514), .ZN(n20542) );
  NOR2_X1 U22595 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20542), .ZN(n20529) );
  OAI22_X1 U22596 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n20516), .B1(n20532), 
        .B2(n20515), .ZN(n20517) );
  AOI211_X1 U22597 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n20523), .A(
        n20529), .B(n20517), .ZN(n20520) );
  NOR2_X1 U22598 ( .A1(n20543), .A2(n20518), .ZN(n20534) );
  OAI21_X1 U22599 ( .B1(n20522), .B2(n20534), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20519) );
  OAI211_X1 U22600 ( .C1(n21261), .C2(n20521), .A(n20520), .B(n20519), .ZN(
        P3_U2641) );
  NAND2_X1 U22601 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20530), .ZN(n20541) );
  AOI22_X1 U22602 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n20523), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n20522), .ZN(n20540) );
  INV_X1 U22603 ( .A(n20524), .ZN(n20538) );
  OR2_X1 U22604 ( .A1(n20526), .A2(n20525), .ZN(n20527) );
  NOR2_X1 U22605 ( .A1(n20528), .A2(n20527), .ZN(n20537) );
  INV_X1 U22606 ( .A(n20529), .ZN(n20531) );
  AOI21_X1 U22607 ( .B1(n20532), .B2(n20531), .A(n20530), .ZN(n20536) );
  AND2_X1 U22608 ( .A1(n20534), .A2(n20533), .ZN(n20535) );
  OAI211_X1 U22609 ( .C1(n20542), .C2(n20541), .A(n20540), .B(n20539), .ZN(
        P3_U2640) );
  NAND2_X1 U22610 ( .A1(n20544), .A2(n20543), .ZN(n20546) );
  AOI22_X1 U22611 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n20546), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n20545), .ZN(n20549) );
  NAND3_X1 U22612 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20547), .A3(
        n20767), .ZN(n20548) );
  OAI211_X1 U22613 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20550), .A(
        n20549), .B(n20548), .ZN(P3_U2671) );
  OAI22_X2 U22614 ( .A1(n11033), .A2(n20553), .B1(n20552), .B2(n20551), .ZN(
        n20584) );
  NAND2_X1 U22615 ( .A1(n20584), .A2(n20554), .ZN(n20708) );
  NOR4_X1 U22616 ( .A1(n20556), .A2(n20563), .A3(n20562), .A4(n20555), .ZN(
        n20616) );
  NAND2_X1 U22617 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n20584), .ZN(n20730) );
  NAND4_X1 U22618 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n20557) );
  NOR2_X1 U22619 ( .A1(n20730), .A2(n20557), .ZN(n20558) );
  NAND4_X1 U22620 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(n20558), .ZN(n20722) );
  NOR2_X1 U22621 ( .A1(n20649), .A2(n20722), .ZN(n20590) );
  AND3_X1 U22622 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20616), .A3(n20590), .ZN(
        n20566) );
  NAND2_X1 U22623 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20566), .ZN(n20712) );
  INV_X1 U22624 ( .A(n20712), .ZN(n20713) );
  AOI21_X1 U22625 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n20707), .A(n20566), .ZN(
        n20560) );
  INV_X1 U22626 ( .A(n20584), .ZN(n20734) );
  OAI222_X1 U22627 ( .A1(n20708), .A2(n20561), .B1(n20713), .B2(n20560), .C1(
        n20739), .C2(n20559), .ZN(P3_U2722) );
  NAND2_X1 U22628 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20590), .ZN(n20578) );
  NOR2_X1 U22629 ( .A1(n20562), .A2(n20578), .ZN(n20582) );
  NAND2_X1 U22630 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20582), .ZN(n20573) );
  NOR2_X1 U22631 ( .A1(n20563), .A2(n20573), .ZN(n20571) );
  AOI21_X1 U22632 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20707), .A(n20571), .ZN(
        n20565) );
  OAI222_X1 U22633 ( .A1(n20708), .A2(n20567), .B1(n20566), .B2(n20565), .C1(
        n20739), .C2(n20564), .ZN(P3_U2723) );
  INV_X1 U22634 ( .A(n20573), .ZN(n20568) );
  AOI21_X1 U22635 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20707), .A(n20568), .ZN(
        n20570) );
  OAI222_X1 U22636 ( .A1(n20708), .A2(n20572), .B1(n20571), .B2(n20570), .C1(
        n20739), .C2(n20569), .ZN(P3_U2724) );
  OAI211_X1 U22637 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n20582), .A(n20707), .B(
        n20573), .ZN(n20576) );
  NAND2_X1 U22638 ( .A1(n20727), .A2(n20574), .ZN(n20575) );
  OAI211_X1 U22639 ( .C1(n20708), .C2(n20577), .A(n20576), .B(n20575), .ZN(
        P3_U2725) );
  INV_X1 U22640 ( .A(n20578), .ZN(n20579) );
  AOI21_X1 U22641 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20707), .A(n20579), .ZN(
        n20581) );
  OAI222_X1 U22642 ( .A1(n20708), .A2(n20583), .B1(n20582), .B2(n20581), .C1(
        n20739), .C2(n20580), .ZN(P3_U2726) );
  NAND2_X1 U22643 ( .A1(n20585), .A2(n20584), .ZN(n20729) );
  NOR3_X1 U22644 ( .A1(n20586), .A2(n20728), .A3(n20729), .ZN(n20609) );
  NAND2_X1 U22645 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n20613), .ZN(n20600) );
  NOR2_X1 U22646 ( .A1(n20587), .A2(n20600), .ZN(n20603) );
  NAND2_X1 U22647 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20603), .ZN(n20591) );
  NOR2_X1 U22648 ( .A1(n20588), .A2(n20591), .ZN(n20594) );
  AOI21_X1 U22649 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20707), .A(n20594), .ZN(
        n20589) );
  OAI222_X1 U22650 ( .A1(n20697), .A2(n20708), .B1(n20590), .B2(n20589), .C1(
        n20739), .C2(n20811), .ZN(P3_U2728) );
  INV_X1 U22651 ( .A(n20591), .ZN(n20598) );
  AOI21_X1 U22652 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20707), .A(n20598), .ZN(
        n20593) );
  OAI222_X1 U22653 ( .A1(n20595), .A2(n20708), .B1(n20594), .B2(n20593), .C1(
        n20739), .C2(n20592), .ZN(P3_U2729) );
  AOI21_X1 U22654 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20707), .A(n20603), .ZN(
        n20597) );
  OAI222_X1 U22655 ( .A1(n20599), .A2(n20708), .B1(n20598), .B2(n20597), .C1(
        n20739), .C2(n20596), .ZN(P3_U2730) );
  INV_X1 U22656 ( .A(n20600), .ZN(n20607) );
  AOI21_X1 U22657 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20707), .A(n20607), .ZN(
        n20602) );
  OAI222_X1 U22658 ( .A1(n20604), .A2(n20708), .B1(n20603), .B2(n20602), .C1(
        n20739), .C2(n20601), .ZN(P3_U2731) );
  AOI21_X1 U22659 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20707), .A(n20613), .ZN(
        n20606) );
  OAI222_X1 U22660 ( .A1(n20608), .A2(n20708), .B1(n20607), .B2(n20606), .C1(
        n20739), .C2(n20605), .ZN(P3_U2732) );
  AOI21_X1 U22661 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n20707), .A(n20609), .ZN(
        n20612) );
  INV_X1 U22662 ( .A(n20610), .ZN(n20611) );
  OAI222_X1 U22663 ( .A1(n20614), .A2(n20708), .B1(n20613), .B2(n20612), .C1(
        n20739), .C2(n20611), .ZN(P3_U2733) );
  NOR2_X2 U22664 ( .A1(n20615), .A2(n20707), .ZN(n20700) );
  NOR2_X2 U22665 ( .A1(n20799), .A2(n20707), .ZN(n20699) );
  AOI22_X1 U22666 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20699), .ZN(n20618) );
  NAND4_X1 U22667 ( .A1(n20719), .A2(n20616), .A3(P3_EAX_REG_13__SCAN_IN), 
        .A4(P3_EAX_REG_14__SCAN_IN), .ZN(n20706) );
  NOR2_X1 U22668 ( .A1(n20649), .A2(n20701), .ZN(n20642) );
  NAND2_X1 U22669 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n20642), .ZN(n20641) );
  NAND2_X1 U22670 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20630), .ZN(n20620) );
  NAND2_X1 U22671 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20625), .ZN(n20629) );
  OAI211_X1 U22672 ( .C1(n20625), .C2(P3_EAX_REG_21__SCAN_IN), .A(n20707), .B(
        n20629), .ZN(n20617) );
  OAI211_X1 U22673 ( .C1(n20619), .C2(n20739), .A(n20618), .B(n20617), .ZN(
        P3_U2714) );
  AOI22_X1 U22674 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20699), .ZN(n20622) );
  OAI211_X1 U22675 ( .C1(n20630), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20707), .B(
        n20620), .ZN(n20621) );
  OAI211_X1 U22676 ( .C1(n20623), .C2(n20739), .A(n20622), .B(n20621), .ZN(
        P3_U2715) );
  AOI22_X1 U22677 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20699), .B1(n20727), .B2(
        n20624), .ZN(n20628) );
  OAI22_X1 U22678 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20729), .B1(n20720), 
        .B2(n20625), .ZN(n20626) );
  AOI22_X1 U22679 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20700), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n20626), .ZN(n20627) );
  OAI211_X1 U22680 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n20629), .A(n20628), .B(
        n20627), .ZN(P3_U2713) );
  AOI22_X1 U22681 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20699), .ZN(n20634) );
  AOI211_X1 U22682 ( .C1(n20631), .C2(n20636), .A(n20630), .B(n20720), .ZN(
        n20632) );
  INV_X1 U22683 ( .A(n20632), .ZN(n20633) );
  OAI211_X1 U22684 ( .C1(n20635), .C2(n20739), .A(n20634), .B(n20633), .ZN(
        P3_U2716) );
  AOI22_X1 U22685 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20699), .ZN(n20639) );
  OAI211_X1 U22686 ( .C1(n20637), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20707), .B(
        n20636), .ZN(n20638) );
  OAI211_X1 U22687 ( .C1(n20640), .C2(n20739), .A(n20639), .B(n20638), .ZN(
        P3_U2717) );
  AOI22_X1 U22688 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20699), .ZN(n20644) );
  OAI211_X1 U22689 ( .C1(n20642), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20707), .B(
        n20641), .ZN(n20643) );
  OAI211_X1 U22690 ( .C1(n20645), .C2(n20739), .A(n20644), .B(n20643), .ZN(
        P3_U2718) );
  NAND4_X1 U22691 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_20__SCAN_IN), .ZN(n20646)
         );
  NOR4_X2 U22692 ( .A1(n20701), .A2(n20648), .A3(n20647), .A4(n20646), .ZN(
        n20694) );
  NAND2_X1 U22693 ( .A1(n20694), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20693) );
  INV_X1 U22694 ( .A(n20656), .ZN(n20652) );
  OAI21_X1 U22695 ( .B1(n20720), .B2(n20650), .A(n20687), .ZN(n20651) );
  AOI22_X1 U22696 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20699), .B1(n20652), .B2(
        n20651), .ZN(n20655) );
  AOI22_X1 U22697 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20700), .B1(n20727), .B2(
        n20653), .ZN(n20654) );
  NAND2_X1 U22698 ( .A1(n20655), .A2(n20654), .ZN(P3_U2710) );
  AOI22_X1 U22699 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20699), .ZN(n20658) );
  OAI211_X1 U22700 ( .C1(n20656), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20707), .B(
        n20680), .ZN(n20657) );
  OAI211_X1 U22701 ( .C1(n20659), .C2(n20739), .A(n20658), .B(n20657), .ZN(
        P3_U2709) );
  NAND2_X1 U22702 ( .A1(n20664), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20662) );
  OAI21_X1 U22703 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20729), .A(n20668), .ZN(
        n20660) );
  AOI22_X1 U22704 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20699), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20660), .ZN(n20661) );
  OAI21_X1 U22705 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n20662), .A(n20661), .ZN(
        P3_U2704) );
  AOI22_X1 U22706 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20699), .B1(n20727), .B2(
        n20663), .ZN(n20666) );
  AOI22_X1 U22707 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20700), .B1(n20664), .B2(
        n20667), .ZN(n20665) );
  OAI211_X1 U22708 ( .C1(n20668), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        P3_U2705) );
  OAI21_X1 U22709 ( .B1(n20720), .B2(n20669), .A(n20675), .ZN(n20670) );
  AOI22_X1 U22710 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20699), .B1(n20671), .B2(
        n20670), .ZN(n20674) );
  AOI22_X1 U22711 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20700), .B1(n20727), .B2(
        n20672), .ZN(n20673) );
  NAND2_X1 U22712 ( .A1(n20674), .A2(n20673), .ZN(P3_U2706) );
  AOI22_X1 U22713 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20699), .ZN(n20677) );
  OAI211_X1 U22714 ( .C1(n20679), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20707), .B(
        n20675), .ZN(n20676) );
  OAI211_X1 U22715 ( .C1(n20678), .C2(n20739), .A(n20677), .B(n20676), .ZN(
        P3_U2707) );
  INV_X1 U22716 ( .A(n20679), .ZN(n20683) );
  OAI21_X1 U22717 ( .B1(n20720), .B2(n20681), .A(n20680), .ZN(n20682) );
  AOI22_X1 U22718 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20699), .B1(n20683), .B2(
        n20682), .ZN(n20686) );
  AOI22_X1 U22719 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20700), .B1(n20727), .B2(
        n20684), .ZN(n20685) );
  NAND2_X1 U22720 ( .A1(n20686), .A2(n20685), .ZN(P3_U2708) );
  AOI22_X1 U22721 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20699), .ZN(n20690) );
  OAI211_X1 U22722 ( .C1(n20688), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20707), .B(
        n20687), .ZN(n20689) );
  OAI211_X1 U22723 ( .C1(n20691), .C2(n20739), .A(n20690), .B(n20689), .ZN(
        P3_U2711) );
  INV_X1 U22724 ( .A(n20700), .ZN(n20698) );
  AOI22_X1 U22725 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n20699), .B1(n20727), .B2(
        n20692), .ZN(n20696) );
  OAI211_X1 U22726 ( .C1(n20694), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20707), .B(
        n20693), .ZN(n20695) );
  OAI211_X1 U22727 ( .C1(n20698), .C2(n20697), .A(n20696), .B(n20695), .ZN(
        P3_U2712) );
  AOI22_X1 U22728 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20700), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20699), .ZN(n20704) );
  OAI211_X1 U22729 ( .C1(n20702), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20707), .B(
        n20701), .ZN(n20703) );
  OAI211_X1 U22730 ( .C1(n20705), .C2(n20739), .A(n20704), .B(n20703), .ZN(
        P3_U2719) );
  NAND2_X1 U22731 ( .A1(n20707), .A2(n20706), .ZN(n20716) );
  INV_X1 U22732 ( .A(n20708), .ZN(n20735) );
  AOI22_X1 U22733 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20735), .B1(n20727), .B2(
        n20709), .ZN(n20710) );
  OAI221_X1 U22734 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n20712), .C1(n20711), 
        .C2(n20716), .A(n20710), .ZN(P3_U2721) );
  NAND2_X1 U22735 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20713), .ZN(n20718) );
  AOI22_X1 U22736 ( .A1(n20727), .A2(n20714), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n20735), .ZN(n20715) );
  OAI221_X1 U22737 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n20718), .C1(n20717), 
        .C2(n20716), .A(n20715), .ZN(P3_U2720) );
  AOI211_X1 U22738 ( .C1(n20722), .C2(n20721), .A(n20720), .B(n20719), .ZN(
        n20723) );
  AOI21_X1 U22739 ( .B1(n20735), .B2(BUF2_REG_8__SCAN_IN), .A(n20723), .ZN(
        n20724) );
  OAI21_X1 U22740 ( .B1(n20725), .B2(n20739), .A(n20724), .ZN(P3_U2727) );
  AOI22_X1 U22741 ( .A1(n20735), .A2(BUF2_REG_1__SCAN_IN), .B1(n20727), .B2(
        n20726), .ZN(n20733) );
  NOR2_X1 U22742 ( .A1(n20728), .A2(n20729), .ZN(n20731) );
  NOR2_X1 U22743 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20729), .ZN(n20736) );
  OAI22_X1 U22744 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n20731), .B1(n20736), .B2(
        n20730), .ZN(n20732) );
  NAND2_X1 U22745 ( .A1(n20733), .A2(n20732), .ZN(P3_U2734) );
  AOI22_X1 U22746 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20735), .B1(n20734), .B2(
        P3_EAX_REG_0__SCAN_IN), .ZN(n20738) );
  INV_X1 U22747 ( .A(n20736), .ZN(n20737) );
  OAI211_X1 U22748 ( .C1(n20740), .C2(n20739), .A(n20738), .B(n20737), .ZN(
        P3_U2735) );
  INV_X1 U22749 ( .A(n20741), .ZN(n20742) );
  INV_X1 U22750 ( .A(n20743), .ZN(n20745) );
  OAI21_X1 U22751 ( .B1(n20745), .B2(n20744), .A(n20779), .ZN(n21207) );
  INV_X1 U22752 ( .A(n21207), .ZN(n21054) );
  AND2_X1 U22753 ( .A1(n20746), .A2(n21054), .ZN(n20749) );
  AOI22_X1 U22754 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21188), .B1(
        n20749), .B2(n20772), .ZN(n21236) );
  AOI222_X1 U22755 ( .A1(n20846), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21236), 
        .B2(n20790), .C1(n20772), .C2(n20792), .ZN(n20747) );
  AOI22_X1 U22756 ( .A1(n20795), .A2(n20772), .B1(n20747), .B2(n20793), .ZN(
        P3_U3290) );
  INV_X1 U22757 ( .A(n21206), .ZN(n20907) );
  AOI21_X1 U22758 ( .B1(n21188), .B2(n20772), .A(n20907), .ZN(n20787) );
  INV_X1 U22759 ( .A(n20787), .ZN(n20757) );
  OAI22_X1 U22760 ( .A1(n20749), .A2(n20748), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20757), .ZN(n21235) );
  AOI22_X1 U22761 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17978), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11313), .ZN(n20766) );
  NOR2_X1 U22762 ( .A1(n20750), .A2(n20846), .ZN(n20763) );
  AOI222_X1 U22763 ( .A1(n21235), .A2(n20790), .B1(n20751), .B2(n20792), .C1(
        n20766), .C2(n20763), .ZN(n20752) );
  AOI22_X1 U22764 ( .A1(n20795), .A2(n20759), .B1(n20752), .B2(n20793), .ZN(
        P3_U3289) );
  AOI22_X1 U22765 ( .A1(n20756), .A2(n20755), .B1(n20754), .B2(n20753), .ZN(
        n20784) );
  AOI211_X1 U22766 ( .C1(n20779), .C2(n20784), .A(n20775), .B(n21240), .ZN(
        n20761) );
  AOI211_X1 U22767 ( .C1(n21240), .C2(n20759), .A(n20758), .B(n20757), .ZN(
        n20760) );
  AOI211_X1 U22768 ( .C1(n21224), .C2(n20762), .A(n20761), .B(n20760), .ZN(
        n21239) );
  INV_X1 U22769 ( .A(n20763), .ZN(n20765) );
  INV_X1 U22770 ( .A(n20792), .ZN(n21266) );
  OAI222_X1 U22771 ( .A1(n21239), .A2(n20767), .B1(n20766), .B2(n20765), .C1(
        n20764), .C2(n21266), .ZN(n20768) );
  INV_X1 U22772 ( .A(n20768), .ZN(n20771) );
  AOI21_X1 U22773 ( .B1(n20792), .B2(n20769), .A(n20795), .ZN(n20770) );
  OAI22_X1 U22774 ( .A1(n20795), .A2(n20771), .B1(n20770), .B2(n21240), .ZN(
        P3_U3288) );
  NOR2_X1 U22775 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20780), .ZN(
        n20788) );
  NAND2_X1 U22776 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20772), .ZN(
        n20778) );
  OAI211_X1 U22777 ( .C1(n20775), .C2(n20774), .A(n21224), .B(n20773), .ZN(
        n20776) );
  OAI22_X1 U22778 ( .A1(n20779), .A2(n20778), .B1(n20777), .B2(n20776), .ZN(
        n20786) );
  NAND2_X1 U22779 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20780), .ZN(
        n20781) );
  OAI22_X1 U22780 ( .A1(n20784), .A2(n20783), .B1(n20782), .B2(n20781), .ZN(
        n20785) );
  AOI211_X1 U22781 ( .C1(n20788), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        n21231) );
  INV_X1 U22782 ( .A(n21231), .ZN(n20789) );
  AOI22_X1 U22783 ( .A1(n20792), .A2(n20791), .B1(n20790), .B2(n20789), .ZN(
        n20794) );
  AOI22_X1 U22784 ( .A1(n20795), .A2(n21232), .B1(n20794), .B2(n20793), .ZN(
        P3_U3285) );
  NAND2_X1 U22785 ( .A1(n21229), .A2(n20796), .ZN(n20798) );
  OAI22_X1 U22786 ( .A1(n20799), .A2(n20798), .B1(n20808), .B2(n20797), .ZN(
        n20806) );
  XOR2_X1 U22787 ( .A(n20800), .B(n20807), .Z(n20802) );
  OAI21_X1 U22788 ( .B1(n20802), .B2(n20801), .A(n21764), .ZN(n21248) );
  NOR3_X1 U22789 ( .A1(n20803), .A2(n21249), .A3(n21248), .ZN(n20805) );
  AOI211_X1 U22790 ( .C1(n20807), .C2(n20806), .A(n20805), .B(n20804), .ZN(
        n20809) );
  AOI221_X4 U22791 ( .B1(n20810), .B2(n20809), .C1(n20808), .C2(n20809), .A(
        n21279), .ZN(n21216) );
  INV_X1 U22792 ( .A(n21087), .ZN(n21230) );
  AOI22_X1 U22793 ( .A1(n21153), .A2(n20812), .B1(n21223), .B2(n20925), .ZN(
        n20922) );
  NOR2_X1 U22794 ( .A1(n21162), .A2(n20824), .ZN(n20814) );
  INV_X1 U22795 ( .A(n20814), .ZN(n20816) );
  NOR2_X1 U22796 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21213), .ZN(
        n20838) );
  NOR2_X1 U22797 ( .A1(n20907), .A2(n20838), .ZN(n20857) );
  NOR3_X1 U22798 ( .A1(n20880), .A2(n17714), .A3(n20888), .ZN(n20890) );
  NAND3_X1 U22799 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20890), .ZN(n20878) );
  NOR2_X1 U22800 ( .A1(n20902), .A2(n20878), .ZN(n20906) );
  NAND2_X1 U22801 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20906), .ZN(
        n21212) );
  NOR2_X1 U22802 ( .A1(n21208), .A2(n21212), .ZN(n20951) );
  NAND2_X1 U22803 ( .A1(n20994), .A2(n20951), .ZN(n21036) );
  NOR2_X1 U22804 ( .A1(n20824), .A2(n21036), .ZN(n20815) );
  INV_X1 U22805 ( .A(n21224), .ZN(n20950) );
  OAI21_X1 U22806 ( .B1(n11313), .B2(n20846), .A(n20856), .ZN(n20858) );
  AND2_X1 U22807 ( .A1(n20858), .A2(n20890), .ZN(n20877) );
  NAND2_X1 U22808 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20877), .ZN(
        n20904) );
  NOR2_X1 U22809 ( .A1(n20813), .A2(n20904), .ZN(n20993) );
  NAND2_X1 U22810 ( .A1(n20814), .A2(n20993), .ZN(n20817) );
  NOR2_X1 U22811 ( .A1(n20950), .A2(n20817), .ZN(n21039) );
  AOI21_X1 U22812 ( .B1(n20857), .B2(n20815), .A(n21039), .ZN(n21002) );
  OAI21_X1 U22813 ( .B1(n20922), .B2(n20816), .A(n21002), .ZN(n20982) );
  AND2_X1 U22814 ( .A1(n21216), .A2(n20982), .ZN(n21142) );
  NOR2_X1 U22815 ( .A1(n21224), .A2(n21213), .ZN(n21197) );
  INV_X1 U22816 ( .A(n21197), .ZN(n20968) );
  INV_X1 U22817 ( .A(n20817), .ZN(n20820) );
  OAI21_X1 U22818 ( .B1(n21036), .B2(n20818), .A(n21213), .ZN(n20819) );
  OAI21_X1 U22819 ( .B1(n20820), .B2(n20950), .A(n20819), .ZN(n21132) );
  OAI22_X1 U22820 ( .A1(n20822), .A2(n21128), .B1(n20821), .B2(n21130), .ZN(
        n20823) );
  AOI211_X1 U22821 ( .C1(n20825), .C2(n20968), .A(n21132), .B(n20823), .ZN(
        n20985) );
  NAND2_X1 U22822 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20951), .ZN(
        n21205) );
  NOR2_X1 U22823 ( .A1(n21162), .A2(n21205), .ZN(n20965) );
  INV_X1 U22824 ( .A(n20965), .ZN(n21050) );
  NOR2_X1 U22825 ( .A1(n20824), .A2(n21050), .ZN(n21038) );
  OAI21_X1 U22826 ( .B1(n21054), .B2(n21038), .A(n21216), .ZN(n21133) );
  AOI21_X1 U22827 ( .B1(n20825), .B2(n21207), .A(n21133), .ZN(n20827) );
  AOI211_X1 U22828 ( .C1(n20985), .C2(n20827), .A(n10990), .B(n20826), .ZN(
        n20828) );
  AOI21_X1 U22829 ( .B1(n21142), .B2(n20829), .A(n20828), .ZN(n20831) );
  OAI211_X1 U22830 ( .C1(n20832), .C2(n21139), .A(n20831), .B(n20830), .ZN(
        P3_U2841) );
  NOR2_X1 U22831 ( .A1(n21224), .A2(n21207), .ZN(n21145) );
  AOI22_X1 U22832 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21213), .B1(
        n21223), .B2(n20837), .ZN(n20833) );
  OAI21_X1 U22833 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21145), .A(
        n20833), .ZN(n20834) );
  AOI22_X1 U22834 ( .A1(n21216), .A2(n20834), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21113), .ZN(n20836) );
  NAND2_X1 U22835 ( .A1(n10990), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20835) );
  OAI211_X1 U22836 ( .C1(n20910), .C2(n20837), .A(n20836), .B(n20835), .ZN(
        P3_U2862) );
  AOI22_X1 U22837 ( .A1(n10990), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21113), .ZN(n20844) );
  NOR2_X1 U22838 ( .A1(n21122), .A2(n20838), .ZN(n20840) );
  NOR2_X1 U22839 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21145), .ZN(
        n20839) );
  MUX2_X1 U22840 ( .A(n20840), .B(n20839), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n20842) );
  AOI22_X1 U22841 ( .A1(n21216), .A2(n20842), .B1(n21014), .B2(n20841), .ZN(
        n20843) );
  OAI211_X1 U22842 ( .C1(n20910), .C2(n20845), .A(n20844), .B(n20843), .ZN(
        P3_U2861) );
  INV_X1 U22843 ( .A(n20858), .ZN(n20861) );
  NAND3_X1 U22844 ( .A1(n21224), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U22845 ( .A1(n20846), .A2(n21207), .ZN(n20995) );
  OAI211_X1 U22846 ( .C1(n20907), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20847), .B(n20995), .ZN(n20848) );
  AOI22_X1 U22847 ( .A1(n21224), .A2(n20861), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20848), .ZN(n20850) );
  NAND3_X1 U22848 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20857), .A3(
        n20856), .ZN(n20849) );
  OAI211_X1 U22849 ( .C1(n20851), .C2(n21230), .A(n20850), .B(n20849), .ZN(
        n20852) );
  AOI22_X1 U22850 ( .A1(n21216), .A2(n20852), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21113), .ZN(n20854) );
  OAI211_X1 U22851 ( .C1(n20855), .C2(n21008), .A(n20854), .B(n20853), .ZN(
        P3_U2860) );
  NOR2_X1 U22852 ( .A1(n20856), .A2(n11313), .ZN(n20859) );
  AOI22_X1 U22853 ( .A1(n20858), .A2(n21224), .B1(n20857), .B2(n20859), .ZN(
        n20881) );
  AOI21_X1 U22854 ( .B1(n20859), .B2(n20995), .A(n20907), .ZN(n20860) );
  AOI211_X1 U22855 ( .C1(n21224), .C2(n20861), .A(n20860), .B(n17714), .ZN(
        n20870) );
  AOI211_X1 U22856 ( .C1(n20881), .C2(n17714), .A(n20870), .B(n21154), .ZN(
        n20865) );
  OAI22_X1 U22857 ( .A1(n20910), .A2(n20863), .B1(n21008), .B2(n20862), .ZN(
        n20864) );
  NOR2_X1 U22858 ( .A1(n20865), .A2(n20864), .ZN(n20867) );
  OAI211_X1 U22859 ( .C1(n21186), .C2(n17714), .A(n20867), .B(n20866), .ZN(
        P3_U2859) );
  NAND2_X1 U22860 ( .A1(n10990), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n20876) );
  OAI22_X1 U22861 ( .A1(n21230), .A2(n20869), .B1(n21128), .B2(n20868), .ZN(
        n20874) );
  INV_X1 U22862 ( .A(n20881), .ZN(n20889) );
  AND2_X1 U22863 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20889), .ZN(
        n20872) );
  NOR2_X1 U22864 ( .A1(n21122), .A2(n20870), .ZN(n20871) );
  MUX2_X1 U22865 ( .A(n20872), .B(n20871), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n20873) );
  OAI21_X1 U22866 ( .B1(n20874), .B2(n20873), .A(n21216), .ZN(n20875) );
  OAI211_X1 U22867 ( .C1(n21186), .C2(n20880), .A(n20876), .B(n20875), .ZN(
        P3_U2858) );
  OAI211_X1 U22868 ( .C1(n20877), .C2(n20950), .A(n21216), .B(n20995), .ZN(
        n20879) );
  OAI221_X1 U22869 ( .B1(n20879), .B2(n21206), .C1(n20879), .C2(n20878), .A(
        n21199), .ZN(n20897) );
  NOR4_X1 U22870 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20881), .A3(
        n17714), .A4(n20880), .ZN(n20885) );
  OAI22_X1 U22871 ( .A1(n20910), .A2(n20883), .B1(n21008), .B2(n20882), .ZN(
        n20884) );
  AOI21_X1 U22872 ( .B1(n21216), .B2(n20885), .A(n20884), .ZN(n20887) );
  NAND2_X1 U22873 ( .A1(n10990), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n20886) );
  OAI211_X1 U22874 ( .C1(n20888), .C2(n20897), .A(n20887), .B(n20886), .ZN(
        P3_U2857) );
  NAND2_X1 U22875 ( .A1(n20890), .A2(n20889), .ZN(n20901) );
  NOR2_X1 U22876 ( .A1(n20901), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20894) );
  OAI22_X1 U22877 ( .A1(n20910), .A2(n20892), .B1(n21008), .B2(n20891), .ZN(
        n20893) );
  AOI21_X1 U22878 ( .B1(n20894), .B2(n21216), .A(n20893), .ZN(n20896) );
  NAND2_X1 U22879 ( .A1(n10990), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n20895) );
  OAI211_X1 U22880 ( .C1(n20902), .C2(n20897), .A(n20896), .B(n20895), .ZN(
        P3_U2856) );
  OAI22_X1 U22881 ( .A1(n21199), .A2(n20898), .B1(n20903), .B2(n21186), .ZN(
        n20899) );
  AOI21_X1 U22882 ( .B1(n21014), .B2(n20900), .A(n20899), .ZN(n20909) );
  NOR2_X1 U22883 ( .A1(n20902), .A2(n20901), .ZN(n20920) );
  AOI21_X1 U22884 ( .B1(n21224), .B2(n20904), .A(n20903), .ZN(n20905) );
  OAI211_X1 U22885 ( .C1(n20907), .C2(n20906), .A(n20905), .B(n20995), .ZN(
        n20912) );
  OAI211_X1 U22886 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n20920), .A(
        n21216), .B(n20912), .ZN(n20908) );
  OAI211_X1 U22887 ( .C1(n20911), .C2(n20910), .A(n20909), .B(n20908), .ZN(
        P3_U2855) );
  AOI22_X1 U22888 ( .A1(n10990), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21113), .ZN(n20918) );
  NAND3_X1 U22889 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20920), .A3(
        n21208), .ZN(n20914) );
  NAND3_X1 U22890 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21175), .A3(
        n20912), .ZN(n20913) );
  OAI211_X1 U22891 ( .C1(n20915), .C2(n21130), .A(n20914), .B(n20913), .ZN(
        n20916) );
  AOI22_X1 U22892 ( .A1(n21216), .A2(n20916), .B1(n21220), .B2(n20915), .ZN(
        n20917) );
  OAI211_X1 U22893 ( .C1(n21008), .C2(n20919), .A(n20918), .B(n20917), .ZN(
        P3_U2854) );
  NAND2_X1 U22894 ( .A1(n20921), .A2(n20920), .ZN(n20970) );
  NAND2_X1 U22895 ( .A1(n20922), .A2(n20970), .ZN(n20941) );
  NAND2_X1 U22896 ( .A1(n21216), .A2(n20941), .ZN(n21222) );
  AOI22_X1 U22897 ( .A1(n10990), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n21220), 
        .B2(n20923), .ZN(n20931) );
  NOR2_X1 U22898 ( .A1(n21153), .A2(n21223), .ZN(n21161) );
  NAND2_X1 U22899 ( .A1(n21153), .A2(n21152), .ZN(n20924) );
  OR2_X1 U22900 ( .A1(n20950), .A2(n20993), .ZN(n20952) );
  OAI211_X1 U22901 ( .C1(n20925), .C2(n21128), .A(n20924), .B(n20952), .ZN(
        n21210) );
  AOI221_X1 U22902 ( .B1(n21214), .B2(n21207), .C1(n21205), .C2(n21207), .A(
        n21210), .ZN(n20926) );
  OAI211_X1 U22903 ( .C1(n20927), .C2(n21161), .A(n20926), .B(n21186), .ZN(
        n21200) );
  AOI21_X1 U22904 ( .B1(n20927), .B2(n20951), .A(n21188), .ZN(n20928) );
  AOI21_X1 U22905 ( .B1(n21224), .B2(n20933), .A(n20928), .ZN(n20935) );
  OAI21_X1 U22906 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n21054), .A(
        n20935), .ZN(n20929) );
  OAI211_X1 U22907 ( .C1(n21200), .C2(n20929), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n21199), .ZN(n20930) );
  OAI211_X1 U22908 ( .C1(n20932), .C2(n21222), .A(n20931), .B(n20930), .ZN(
        P3_U2851) );
  INV_X1 U22909 ( .A(n20933), .ZN(n20942) );
  NOR2_X1 U22910 ( .A1(n20934), .A2(n21205), .ZN(n20949) );
  AOI211_X1 U22911 ( .C1(n21184), .C2(n21213), .A(n21185), .B(n21207), .ZN(
        n20939) );
  OAI211_X1 U22912 ( .C1(n20936), .C2(n21130), .A(n20935), .B(n20952), .ZN(
        n20937) );
  AOI21_X1 U22913 ( .B1(n21223), .B2(n20938), .A(n20937), .ZN(n21187) );
  OAI21_X1 U22914 ( .B1(n20949), .B2(n20939), .A(n21187), .ZN(n20940) );
  OAI221_X1 U22915 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n20942), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n20941), .A(n20940), .ZN(
        n20946) );
  AOI22_X1 U22916 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21113), .B1(
        n21220), .B2(n20943), .ZN(n20945) );
  OAI211_X1 U22917 ( .C1(n21154), .C2(n20946), .A(n20945), .B(n20944), .ZN(
        P3_U2850) );
  NOR3_X1 U22918 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n20947), .A3(
        n20970), .ZN(n20960) );
  AOI21_X1 U22919 ( .B1(n21188), .B2(n21145), .A(n20948), .ZN(n20953) );
  OAI22_X1 U22920 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n20950), .B1(
        n21054), .B2(n20949), .ZN(n21191) );
  OR2_X1 U22921 ( .A1(n21188), .A2(n20951), .ZN(n21198) );
  NAND2_X1 U22922 ( .A1(n20952), .A2(n21198), .ZN(n20966) );
  NOR3_X1 U22923 ( .A1(n20953), .A2(n21191), .A3(n20966), .ZN(n20955) );
  OAI22_X1 U22924 ( .A1(n20955), .A2(n20963), .B1(n21130), .B2(n20954), .ZN(
        n20959) );
  OAI22_X1 U22925 ( .A1(n20957), .A2(n21139), .B1(n21008), .B2(n20956), .ZN(
        n20958) );
  AOI221_X1 U22926 ( .B1(n20960), .B2(n21216), .C1(n20959), .C2(n21216), .A(
        n20958), .ZN(n20962) );
  OAI211_X1 U22927 ( .C1(n21186), .C2(n20963), .A(n20962), .B(n20961), .ZN(
        P3_U2848) );
  NOR3_X1 U22928 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21130), .A3(
        n20964), .ZN(n20972) );
  AOI21_X1 U22929 ( .B1(n21054), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n20965), .ZN(n20967) );
  AOI211_X1 U22930 ( .C1(n20968), .C2(n20969), .A(n20967), .B(n20966), .ZN(
        n20975) );
  NOR3_X1 U22931 ( .A1(n20975), .A2(n20970), .A3(n20969), .ZN(n20971) );
  AOI211_X1 U22932 ( .C1(n21223), .C2(n20973), .A(n20972), .B(n20971), .ZN(
        n20981) );
  AOI22_X1 U22933 ( .A1(n10990), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n21220), 
        .B2(n20974), .ZN(n20980) );
  INV_X1 U22934 ( .A(n20975), .ZN(n21174) );
  NAND2_X1 U22935 ( .A1(n21153), .A2(n20976), .ZN(n20977) );
  OAI211_X1 U22936 ( .C1(n20978), .C2(n21128), .A(n21216), .B(n20977), .ZN(
        n21176) );
  OAI211_X1 U22937 ( .C1(n21174), .C2(n21176), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21199), .ZN(n20979) );
  OAI211_X1 U22938 ( .C1(n20981), .C2(n21154), .A(n20980), .B(n20979), .ZN(
        P3_U2847) );
  NAND2_X1 U22939 ( .A1(n20983), .A2(n20982), .ZN(n21026) );
  AOI21_X1 U22940 ( .B1(n21027), .B2(n21026), .A(n21154), .ZN(n20987) );
  OAI22_X1 U22941 ( .A1(n21027), .A2(n21207), .B1(n20997), .B2(n21050), .ZN(
        n20984) );
  OAI211_X1 U22942 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21197), .A(
        n20985), .B(n20984), .ZN(n20986) );
  AOI22_X1 U22943 ( .A1(n21220), .A2(n20988), .B1(n20987), .B2(n20986), .ZN(
        n20990) );
  NAND2_X1 U22944 ( .A1(n10990), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n20989) );
  OAI211_X1 U22945 ( .C1(n21186), .C2(n21027), .A(n20990), .B(n20989), .ZN(
        P3_U2840) );
  AOI22_X1 U22946 ( .A1(n10990), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21113), .ZN(n21006) );
  NOR3_X1 U22947 ( .A1(n21027), .A2(n20992), .A3(n20991), .ZN(n21037) );
  NAND2_X1 U22948 ( .A1(n21012), .A2(n21037), .ZN(n21001) );
  NAND2_X1 U22949 ( .A1(n20994), .A2(n20993), .ZN(n21156) );
  OAI21_X1 U22950 ( .B1(n20997), .B2(n21156), .A(n21224), .ZN(n21114) );
  INV_X1 U22951 ( .A(n21036), .ZN(n20996) );
  NAND2_X1 U22952 ( .A1(n20996), .A2(n20995), .ZN(n21155) );
  OAI21_X1 U22953 ( .B1(n20997), .B2(n21155), .A(n21206), .ZN(n21108) );
  OAI211_X1 U22954 ( .C1(n21122), .C2(n20998), .A(n21114), .B(n21108), .ZN(
        n21010) );
  AOI22_X1 U22955 ( .A1(n21153), .A2(n20999), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21010), .ZN(n21000) );
  OAI21_X1 U22956 ( .B1(n21002), .B2(n21001), .A(n21000), .ZN(n21004) );
  AOI22_X1 U22957 ( .A1(n21216), .A2(n21004), .B1(n21220), .B2(n21003), .ZN(
        n21005) );
  OAI211_X1 U22958 ( .C1(n21008), .C2(n21007), .A(n21006), .B(n21005), .ZN(
        P3_U2837) );
  INV_X1 U22959 ( .A(n21009), .ZN(n21021) );
  NOR2_X1 U22960 ( .A1(n21046), .A2(n21130), .ZN(n21011) );
  AOI211_X1 U22961 ( .C1(n21175), .C2(n21012), .A(n21011), .B(n21010), .ZN(
        n21015) );
  NAND2_X1 U22962 ( .A1(n21014), .A2(n21013), .ZN(n21030) );
  OAI221_X1 U22963 ( .B1(n21154), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n21154), .C2(n21015), .A(n21030), .ZN(n21018) );
  NOR2_X1 U22964 ( .A1(n21026), .A2(n21016), .ZN(n21017) );
  AOI222_X1 U22965 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21018), 
        .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21113), .C1(n21018), 
        .C2(n21017), .ZN(n21020) );
  OAI211_X1 U22966 ( .C1(n21021), .C2(n21139), .A(n21020), .B(n21019), .ZN(
        P3_U2836) );
  AOI22_X1 U22967 ( .A1(n21153), .A2(n21023), .B1(n21206), .B2(n21022), .ZN(
        n21024) );
  OAI21_X1 U22968 ( .B1(n21051), .B2(n21156), .A(n21224), .ZN(n21052) );
  NAND4_X1 U22969 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21024), .A3(
        n21108), .A4(n21052), .ZN(n21025) );
  AOI22_X1 U22970 ( .A1(n21216), .A2(n21025), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21113), .ZN(n21031) );
  NOR2_X1 U22971 ( .A1(n21027), .A2(n21026), .ZN(n21107) );
  NAND2_X1 U22972 ( .A1(n21107), .A2(n21028), .ZN(n21091) );
  AOI22_X1 U22973 ( .A1(n21031), .A2(n21030), .B1(n21029), .B2(n21091), .ZN(
        n21032) );
  AOI211_X1 U22974 ( .C1(n21220), .C2(n21034), .A(n21033), .B(n21032), .ZN(
        n21035) );
  INV_X1 U22975 ( .A(n21035), .ZN(P3_U2835) );
  INV_X1 U22976 ( .A(n21095), .ZN(n21045) );
  NOR2_X1 U22977 ( .A1(n21036), .A2(n21051), .ZN(n21049) );
  NAND2_X1 U22978 ( .A1(n21049), .A2(n21213), .ZN(n21043) );
  OAI221_X1 U22979 ( .B1(n21039), .B2(n21038), .C1(n21039), .C2(n21207), .A(
        n21037), .ZN(n21042) );
  AOI211_X1 U22980 ( .C1(n21043), .C2(n21042), .A(n21041), .B(n21040), .ZN(
        n21073) );
  AOI21_X1 U22981 ( .B1(n21153), .B2(n21096), .A(n21073), .ZN(n21044) );
  NAND2_X1 U22982 ( .A1(n21046), .A2(n21065), .ZN(n21048) );
  AOI22_X1 U22983 ( .A1(n21153), .A2(n21048), .B1(n21223), .B2(n21047), .ZN(
        n21067) );
  INV_X1 U22984 ( .A(n21049), .ZN(n21056) );
  NOR2_X1 U22985 ( .A1(n21051), .A2(n21050), .ZN(n21053) );
  OAI221_X1 U22986 ( .B1(n21054), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n21054), .C2(n21053), .A(n21052), .ZN(n21055) );
  AOI21_X1 U22987 ( .B1(n21213), .B2(n21056), .A(n21055), .ZN(n21064) );
  OAI211_X1 U22988 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n21197), .A(
        n21064), .B(n21186), .ZN(n21098) );
  AOI21_X1 U22989 ( .B1(n21057), .B2(n21175), .A(n21098), .ZN(n21058) );
  AOI21_X1 U22990 ( .B1(n21067), .B2(n21058), .A(n10990), .ZN(n21060) );
  OAI222_X1 U22991 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21216), 
        .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21066), .C1(n21060), 
        .C2(n21059), .ZN(n21062) );
  OAI211_X1 U22992 ( .C1(n21063), .C2(n21139), .A(n21062), .B(n21061), .ZN(
        P3_U2833) );
  OAI211_X1 U22993 ( .C1(n21122), .C2(n21065), .A(n21064), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21076) );
  INV_X1 U22994 ( .A(n21076), .ZN(n21068) );
  OAI211_X1 U22995 ( .C1(n21071), .C2(n21139), .A(n21070), .B(n21069), .ZN(
        P3_U2832) );
  AND2_X1 U22996 ( .A1(n17978), .A2(n21072), .ZN(n21074) );
  AOI22_X1 U22997 ( .A1(n21153), .A2(n21075), .B1(n21074), .B2(n21073), .ZN(
        n21078) );
  NAND3_X1 U22998 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21175), .A3(
        n21076), .ZN(n21077) );
  OAI211_X1 U22999 ( .C1(n21079), .C2(n21128), .A(n21078), .B(n21077), .ZN(
        n21080) );
  AOI21_X1 U23000 ( .B1(n21082), .B2(n21220), .A(n21081), .ZN(n21085) );
  INV_X1 U23001 ( .A(n21083), .ZN(n21084) );
  OAI211_X1 U23002 ( .C1(n17978), .C2(n21186), .A(n21085), .B(n21084), .ZN(
        P3_U2831) );
  AND2_X1 U23003 ( .A1(n21087), .A2(n21086), .ZN(n21088) );
  OAI22_X1 U23004 ( .A1(n21092), .A2(n21091), .B1(n21090), .B2(n21094), .ZN(
        n21093) );
  AOI22_X1 U23005 ( .A1(n21216), .A2(n21093), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21199), .ZN(n21106) );
  NAND2_X1 U23006 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21094), .ZN(
        n21099) );
  OAI22_X1 U23007 ( .A1(n21096), .A2(n21130), .B1(n21095), .B2(n21128), .ZN(
        n21097) );
  OR3_X1 U23008 ( .A1(n21102), .A2(n21139), .A3(n21101), .ZN(n21104) );
  AOI21_X1 U23009 ( .B1(n21107), .B2(n21186), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21119) );
  INV_X1 U23010 ( .A(n21108), .ZN(n21112) );
  OAI22_X1 U23011 ( .A1(n21110), .A2(n21128), .B1(n21109), .B2(n21130), .ZN(
        n21111) );
  NOR3_X1 U23012 ( .A1(n21113), .A2(n21112), .A3(n21111), .ZN(n21121) );
  NAND3_X1 U23013 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21121), .A3(
        n21114), .ZN(n21115) );
  NAND2_X1 U23014 ( .A1(n21199), .A2(n21115), .ZN(n21120) );
  AOI21_X1 U23015 ( .B1(n21117), .B2(n21220), .A(n21116), .ZN(n21118) );
  OAI21_X1 U23016 ( .B1(n21119), .B2(n21120), .A(n21118), .ZN(P3_U2839) );
  AOI21_X1 U23017 ( .B1(n21122), .B2(n21121), .A(n21120), .ZN(n21124) );
  AOI22_X1 U23018 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21124), .B1(
        n21142), .B2(n21123), .ZN(n21126) );
  OAI211_X1 U23019 ( .C1(n21127), .C2(n21139), .A(n21126), .B(n21125), .ZN(
        P3_U2838) );
  OAI22_X1 U23020 ( .A1(n21131), .A2(n21130), .B1(n21129), .B2(n21128), .ZN(
        n21134) );
  NOR3_X1 U23021 ( .A1(n21134), .A2(n21133), .A3(n21132), .ZN(n21135) );
  NOR2_X1 U23022 ( .A1(n21135), .A2(n10990), .ZN(n21147) );
  AOI22_X1 U23023 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21147), .B1(
        n21142), .B2(n21136), .ZN(n21138) );
  OAI211_X1 U23024 ( .C1(n21140), .C2(n21139), .A(n21138), .B(n21137), .ZN(
        P3_U2843) );
  AOI22_X1 U23025 ( .A1(n21220), .A2(n21143), .B1(n21142), .B2(n21141), .ZN(
        n21149) );
  NOR3_X1 U23026 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21145), .A3(
        n21144), .ZN(n21146) );
  OAI21_X1 U23027 ( .B1(n21147), .B2(n21146), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21148) );
  OAI211_X1 U23028 ( .C1(n21150), .C2(n21199), .A(n21149), .B(n21148), .ZN(
        P3_U2842) );
  AOI211_X1 U23029 ( .C1(n21153), .C2(n21152), .A(n21157), .B(n21151), .ZN(
        n21160) );
  AOI221_X1 U23030 ( .B1(n21177), .B2(n21206), .C1(n21155), .C2(n21206), .A(
        n21154), .ZN(n21159) );
  OAI21_X1 U23031 ( .B1(n21157), .B2(n21156), .A(n21224), .ZN(n21158) );
  OAI211_X1 U23032 ( .C1(n21161), .C2(n21160), .A(n21159), .B(n21158), .ZN(
        n21169) );
  OAI221_X1 U23033 ( .B1(n21169), .B2(n21206), .C1(n21169), .C2(n21170), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21167) );
  NOR2_X1 U23034 ( .A1(n21162), .A2(n21222), .ZN(n21178) );
  AOI22_X1 U23035 ( .A1(n21220), .A2(n21164), .B1(n21178), .B2(n21163), .ZN(
        n21165) );
  OAI221_X1 U23036 ( .B1(n10990), .B2(n21167), .C1(n21199), .C2(n21166), .A(
        n21165), .ZN(P3_U2844) );
  AOI22_X1 U23037 ( .A1(n10990), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n21220), 
        .B2(n21168), .ZN(n21173) );
  NAND3_X1 U23038 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21199), .A3(
        n21169), .ZN(n21172) );
  NAND3_X1 U23039 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21178), .A3(
        n21170), .ZN(n21171) );
  NAND3_X1 U23040 ( .A1(n21173), .A2(n21172), .A3(n21171), .ZN(P3_U2845) );
  OAI221_X1 U23041 ( .B1(n21176), .B2(n21175), .C1(n21176), .C2(n21174), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21182) );
  AOI22_X1 U23042 ( .A1(n21179), .A2(n21220), .B1(n21178), .B2(n21177), .ZN(
        n21180) );
  OAI221_X1 U23043 ( .B1(n10990), .B2(n21182), .C1(n21199), .C2(n21181), .A(
        n21180), .ZN(P3_U2846) );
  AOI22_X1 U23044 ( .A1(n10990), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21220), 
        .B2(n21183), .ZN(n21193) );
  NOR2_X1 U23045 ( .A1(n21185), .A2(n21184), .ZN(n21189) );
  OAI211_X1 U23046 ( .C1(n21189), .C2(n21188), .A(n21187), .B(n21186), .ZN(
        n21190) );
  OAI211_X1 U23047 ( .C1(n21191), .C2(n21190), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21199), .ZN(n21192) );
  OAI211_X1 U23048 ( .C1(n21194), .C2(n21222), .A(n21193), .B(n21192), .ZN(
        P3_U2849) );
  NAND2_X1 U23049 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21195), .ZN(
        n21204) );
  AOI22_X1 U23050 ( .A1(n10990), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21220), 
        .B2(n21196), .ZN(n21203) );
  AOI21_X1 U23051 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21198), .A(
        n21197), .ZN(n21201) );
  OAI211_X1 U23052 ( .C1(n21201), .C2(n21200), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21199), .ZN(n21202) );
  OAI211_X1 U23053 ( .C1(n21204), .C2(n21222), .A(n21203), .B(n21202), .ZN(
        P3_U2852) );
  OAI211_X1 U23054 ( .C1(n21208), .C2(n21207), .A(n21206), .B(n21205), .ZN(
        n21209) );
  INV_X1 U23055 ( .A(n21209), .ZN(n21211) );
  AOI211_X1 U23056 ( .C1(n21213), .C2(n21212), .A(n21211), .B(n21210), .ZN(
        n21215) );
  AOI211_X1 U23057 ( .C1(n21216), .C2(n21215), .A(n10990), .B(n21214), .ZN(
        n21217) );
  AOI211_X1 U23058 ( .C1(n21220), .C2(n21219), .A(n21218), .B(n21217), .ZN(
        n21221) );
  OAI21_X1 U23059 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21222), .A(
        n21221), .ZN(P3_U2853) );
  NOR2_X1 U23060 ( .A1(n21224), .A2(n21223), .ZN(n21226) );
  OAI222_X1 U23061 ( .A1(n21230), .A2(n21229), .B1(n21228), .B2(n21227), .C1(
        n21226), .C2(n21225), .ZN(n21281) );
  AOI22_X1 U23062 ( .A1(n21256), .A2(n21232), .B1(n21231), .B2(n21238), .ZN(
        n21247) );
  AOI222_X1 U23063 ( .A1(n21236), .A2(n21235), .B1(n21236), .B2(n21234), .C1(
        n21235), .C2(n21233), .ZN(n21237) );
  NOR2_X1 U23064 ( .A1(n21256), .A2(n21237), .ZN(n21242) );
  AOI22_X1 U23065 ( .A1(n21256), .A2(n21240), .B1(n21239), .B2(n21238), .ZN(
        n21244) );
  INV_X1 U23066 ( .A(n21244), .ZN(n21245) );
  NOR2_X1 U23067 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21246) );
  INV_X1 U23068 ( .A(n21248), .ZN(n21251) );
  NOR3_X1 U23069 ( .A1(n21251), .A2(n21250), .A3(n21249), .ZN(n21280) );
  OAI21_X1 U23070 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21280), .ZN(n21252) );
  AOI211_X1 U23071 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21256), .A(
        n21281), .B(n21255), .ZN(n21270) );
  OAI211_X1 U23072 ( .C1(n21258), .C2(n21257), .A(n21272), .B(n21270), .ZN(
        n21263) );
  OAI221_X1 U23073 ( .B1(n21264), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21264), 
        .C2(n21263), .A(n21262), .ZN(P3_U3282) );
  OAI22_X1 U23074 ( .A1(n21267), .A2(n21266), .B1(n21764), .B2(n21265), .ZN(
        n21278) );
  NOR2_X1 U23075 ( .A1(n21269), .A2(n21268), .ZN(n21276) );
  INV_X1 U23076 ( .A(n21270), .ZN(n21271) );
  AOI22_X1 U23077 ( .A1(n21274), .A2(n21273), .B1(n21272), .B2(n21271), .ZN(
        n21275) );
  OAI221_X1 U23078 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n21278), .C1(n21277), 
        .C2(n21276), .A(n21275), .ZN(P3_U2996) );
  NOR2_X1 U23079 ( .A1(n21280), .A2(n21279), .ZN(n21285) );
  MUX2_X1 U23080 ( .A(P3_MORE_REG_SCAN_IN), .B(n21281), .S(n21285), .Z(
        P3_U3295) );
  INV_X1 U23081 ( .A(n21282), .ZN(n21283) );
  OAI21_X1 U23082 ( .B1(n21285), .B2(n21284), .A(n21283), .ZN(P3_U2637) );
  AOI211_X1 U23083 ( .C1(n21288), .C2(n21716), .A(n21287), .B(n21286), .ZN(
        n21295) );
  INV_X1 U23084 ( .A(n21289), .ZN(n21290) );
  OAI211_X1 U23085 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21291), .A(n21290), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21292) );
  AOI21_X1 U23086 ( .B1(n21292), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21687), 
        .ZN(n21294) );
  NAND2_X1 U23087 ( .A1(n21295), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21293) );
  OAI21_X1 U23088 ( .B1(n21295), .B2(n21294), .A(n21293), .ZN(P1_U3485) );
  AOI21_X1 U23089 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21304), .A(
        n21296), .ZN(n21303) );
  OAI22_X1 U23090 ( .A1(n21298), .A2(n21334), .B1(n21304), .B2(n21297), .ZN(
        n21299) );
  NOR3_X1 U23091 ( .A1(n21303), .A2(n21300), .A3(n21299), .ZN(n21309) );
  AND2_X1 U23092 ( .A1(n21457), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n21302) );
  AND2_X1 U23093 ( .A1(n13552), .A2(n21301), .ZN(n21313) );
  AOI211_X1 U23094 ( .C1(n21304), .C2(n21303), .A(n21302), .B(n21313), .ZN(
        n21308) );
  AOI22_X1 U23095 ( .A1(n21306), .A2(n21462), .B1(n21461), .B2(n21305), .ZN(
        n21307) );
  OAI211_X1 U23096 ( .C1(n21309), .C2(n13552), .A(n21308), .B(n21307), .ZN(
        P1_U3018) );
  INV_X1 U23097 ( .A(n21309), .ZN(n21312) );
  NOR2_X1 U23098 ( .A1(n21616), .A2(n21310), .ZN(n21311) );
  AOI221_X1 U23099 ( .B1(n21313), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n21312), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n21311), .ZN(
        n21317) );
  AOI22_X1 U23100 ( .A1(n21315), .A2(n13561), .B1(n21461), .B2(n21314), .ZN(
        n21316) );
  OAI211_X1 U23101 ( .C1(n21318), .C2(n21430), .A(n21317), .B(n21316), .ZN(
        P1_U3017) );
  INV_X1 U23102 ( .A(n21319), .ZN(n21405) );
  NAND2_X1 U23103 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21405), .ZN(
        n21333) );
  NAND3_X1 U23104 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21407), .ZN(n21335) );
  INV_X1 U23105 ( .A(n21335), .ZN(n21320) );
  OAI21_X1 U23106 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21349), .A(
        n21348), .ZN(n21328) );
  NOR2_X1 U23107 ( .A1(n21320), .A2(n21328), .ZN(n21327) );
  NOR2_X1 U23108 ( .A1(n21321), .A2(n21430), .ZN(n21325) );
  AND2_X1 U23109 ( .A1(n21407), .A2(n21322), .ZN(n21329) );
  OAI22_X1 U23110 ( .A1(n21323), .A2(n21429), .B1(n14718), .B2(n21616), .ZN(
        n21324) );
  AOI211_X1 U23111 ( .C1(n21325), .C2(n14622), .A(n21329), .B(n21324), .ZN(
        n21326) );
  OAI221_X1 U23112 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21333), .C1(
        n21336), .C2(n21327), .A(n21326), .ZN(P1_U3029) );
  AOI211_X1 U23113 ( .C1(n21336), .C2(n21330), .A(n21329), .B(n21328), .ZN(
        n21347) );
  AOI222_X1 U23114 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21457), .B1(n21461), 
        .B2(n21332), .C1(n21462), .C2(n21331), .ZN(n21339) );
  AOI22_X1 U23115 ( .A1(n21336), .A2(n21335), .B1(n21334), .B2(n21333), .ZN(
        n21342) );
  OAI211_X1 U23116 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21342), .B(n21337), .ZN(n21338) );
  OAI211_X1 U23117 ( .C1(n21347), .C2(n13509), .A(n21339), .B(n21338), .ZN(
        P1_U3027) );
  AOI21_X1 U23118 ( .B1(n21341), .B2(n21461), .A(n21340), .ZN(n21345) );
  AOI22_X1 U23119 ( .A1(n21343), .A2(n21462), .B1(n21342), .B2(n21346), .ZN(
        n21344) );
  OAI211_X1 U23120 ( .C1(n21347), .C2(n21346), .A(n21345), .B(n21344), .ZN(
        P1_U3028) );
  NAND2_X1 U23121 ( .A1(n21407), .A2(n21351), .ZN(n21361) );
  OAI211_X1 U23122 ( .C1(n21349), .C2(n21366), .A(n21348), .B(n21361), .ZN(
        n21363) );
  OAI21_X1 U23123 ( .B1(n21351), .B2(n21363), .A(n21350), .ZN(n21391) );
  INV_X1 U23124 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21352) );
  OAI22_X1 U23125 ( .A1(n21509), .A2(n21429), .B1(n21616), .B2(n21352), .ZN(
        n21353) );
  INV_X1 U23126 ( .A(n21353), .ZN(n21356) );
  AOI22_X1 U23127 ( .A1(n21354), .A2(n21462), .B1(n21396), .B2(n21357), .ZN(
        n21355) );
  OAI211_X1 U23128 ( .C1(n21391), .C2(n21357), .A(n21356), .B(n21355), .ZN(
        P1_U3025) );
  INV_X1 U23129 ( .A(n21358), .ZN(n21360) );
  INV_X1 U23130 ( .A(n21496), .ZN(n21359) );
  OAI22_X1 U23131 ( .A1(n21361), .A2(n21360), .B1(n21429), .B2(n21359), .ZN(
        n21362) );
  INV_X1 U23132 ( .A(n21362), .ZN(n21370) );
  AOI22_X1 U23133 ( .A1(n21364), .A2(n21462), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21363), .ZN(n21369) );
  NAND2_X1 U23134 ( .A1(n21457), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n21368) );
  NAND3_X1 U23135 ( .A1(n21366), .A2(n21405), .A3(n21365), .ZN(n21367) );
  NAND4_X1 U23136 ( .A1(n21370), .A2(n21369), .A3(n21368), .A4(n21367), .ZN(
        P1_U3026) );
  NAND2_X1 U23137 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21396), .ZN(
        n21376) );
  OAI22_X1 U23138 ( .A1(n21520), .A2(n21429), .B1(n21616), .B2(n21529), .ZN(
        n21371) );
  INV_X1 U23139 ( .A(n21371), .ZN(n21375) );
  OAI21_X1 U23140 ( .B1(n21372), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n21391), .ZN(n21382) );
  AOI22_X1 U23141 ( .A1(n21373), .A2(n21462), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21382), .ZN(n21374) );
  OAI211_X1 U23142 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n21376), .A(
        n21375), .B(n21374), .ZN(P1_U3024) );
  NOR2_X1 U23143 ( .A1(n21378), .A2(n21377), .ZN(n21387) );
  OAI211_X1 U23144 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n21396), .ZN(n21386) );
  INV_X1 U23145 ( .A(n21531), .ZN(n21381) );
  INV_X1 U23146 ( .A(n21379), .ZN(n21380) );
  AOI21_X1 U23147 ( .B1(n21381), .B2(n21461), .A(n21380), .ZN(n21385) );
  AOI22_X1 U23148 ( .A1(n21383), .A2(n21462), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21382), .ZN(n21384) );
  OAI211_X1 U23149 ( .C1(n21387), .C2(n21386), .A(n21385), .B(n21384), .ZN(
        P1_U3023) );
  INV_X1 U23150 ( .A(n21543), .ZN(n21390) );
  INV_X1 U23151 ( .A(n21388), .ZN(n21389) );
  AOI21_X1 U23152 ( .B1(n21390), .B2(n21461), .A(n21389), .ZN(n21395) );
  OAI21_X1 U23153 ( .B1(n21426), .B2(n21397), .A(n21391), .ZN(n21401) );
  AOI22_X1 U23154 ( .A1(n21392), .A2(n21462), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21401), .ZN(n21394) );
  NAND3_X1 U23155 ( .A1(n21397), .A2(n21398), .A3(n21396), .ZN(n21393) );
  NAND3_X1 U23156 ( .A1(n21395), .A2(n21394), .A3(n21393), .ZN(P1_U3022) );
  AOI22_X1 U23157 ( .A1(n21555), .A2(n21461), .B1(n21457), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n21403) );
  AND2_X1 U23158 ( .A1(n21397), .A2(n21396), .ZN(n21400) );
  XNOR2_X1 U23159 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21398), .ZN(
        n21399) );
  AOI22_X1 U23160 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21401), .B1(
        n21400), .B2(n21399), .ZN(n21402) );
  OAI211_X1 U23161 ( .C1(n21430), .C2(n21404), .A(n21403), .B(n21402), .ZN(
        P1_U3021) );
  NOR2_X1 U23162 ( .A1(n21616), .A2(n21580), .ZN(n21411) );
  AOI22_X1 U23163 ( .A1(n21407), .A2(n21406), .B1(n21405), .B2(n21417), .ZN(
        n21408) );
  AOI21_X1 U23164 ( .B1(n21409), .B2(n21408), .A(n13559), .ZN(n21410) );
  AOI211_X1 U23165 ( .C1(n21461), .C2(n21578), .A(n21411), .B(n21410), .ZN(
        n21414) );
  INV_X1 U23166 ( .A(n21412), .ZN(n21418) );
  NAND3_X1 U23167 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21418), .A3(
        n13559), .ZN(n21413) );
  OAI211_X1 U23168 ( .C1(n21415), .C2(n21430), .A(n21414), .B(n21413), .ZN(
        P1_U3019) );
  AOI21_X1 U23169 ( .B1(n21568), .B2(n21461), .A(n21416), .ZN(n21421) );
  AOI22_X1 U23170 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21419), .B1(
        n21418), .B2(n21417), .ZN(n21420) );
  OAI211_X1 U23171 ( .C1(n21422), .C2(n21430), .A(n21421), .B(n21420), .ZN(
        P1_U3020) );
  NOR2_X1 U23172 ( .A1(n21424), .A2(n21423), .ZN(n21439) );
  NAND2_X1 U23173 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21439), .ZN(
        n21435) );
  OAI21_X1 U23174 ( .B1(n21427), .B2(n21426), .A(n21425), .ZN(n21438) );
  NOR2_X1 U23175 ( .A1(n21616), .A2(n21428), .ZN(n21433) );
  OAI22_X1 U23176 ( .A1(n21431), .A2(n21430), .B1(n21429), .B2(n21624), .ZN(
        n21432) );
  AOI211_X1 U23177 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n21438), .A(
        n21433), .B(n21432), .ZN(n21434) );
  OAI21_X1 U23178 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21435), .A(
        n21434), .ZN(P1_U3013) );
  AOI22_X1 U23179 ( .A1(n21437), .A2(n21462), .B1(n21461), .B2(n21436), .ZN(
        n21441) );
  OAI21_X1 U23180 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21439), .A(
        n21438), .ZN(n21440) );
  OAI211_X1 U23181 ( .C1(n15841), .C2(n21616), .A(n21441), .B(n21440), .ZN(
        P1_U3014) );
  AOI22_X1 U23182 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21442), .B1(
        n21457), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n21447) );
  INV_X1 U23183 ( .A(n21443), .ZN(n21445) );
  AOI22_X1 U23184 ( .A1(n21445), .A2(n21462), .B1(n21461), .B2(n21444), .ZN(
        n21446) );
  OAI211_X1 U23185 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21448), .A(
        n21447), .B(n21446), .ZN(P1_U3012) );
  AOI21_X1 U23186 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21457), .A(n21449), 
        .ZN(n21454) );
  INV_X1 U23187 ( .A(n21450), .ZN(n21452) );
  AOI22_X1 U23188 ( .A1(n21452), .A2(n21462), .B1(n21461), .B2(n21451), .ZN(
        n21453) );
  OAI211_X1 U23189 ( .C1(n21456), .C2(n21455), .A(n21454), .B(n21453), .ZN(
        P1_U3010) );
  AOI22_X1 U23190 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21458), .B1(
        n21457), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n21465) );
  INV_X1 U23191 ( .A(n21459), .ZN(n21463) );
  AOI22_X1 U23192 ( .A1(n21463), .A2(n21462), .B1(n21461), .B2(n21460), .ZN(
        n21464) );
  OAI211_X1 U23193 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21466), .A(
        n21465), .B(n21464), .ZN(P1_U3008) );
  NAND2_X1 U23194 ( .A1(n21651), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n21468) );
  AOI22_X1 U23195 ( .A1(n21652), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21553), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n21467) );
  OAI211_X1 U23196 ( .C1(n14973), .C2(n21483), .A(n21468), .B(n21467), .ZN(
        n21469) );
  INV_X1 U23197 ( .A(n21469), .ZN(n21470) );
  OAI21_X1 U23198 ( .B1(n21472), .B2(n21471), .A(n21470), .ZN(n21473) );
  AOI21_X1 U23199 ( .B1(n21659), .B2(n21474), .A(n21473), .ZN(n21476) );
  NAND2_X1 U23200 ( .A1(n21562), .A2(n14367), .ZN(n21475) );
  OAI211_X1 U23201 ( .C1(n21665), .C2(n21477), .A(n21476), .B(n21475), .ZN(
        P1_U2839) );
  AOI21_X1 U23202 ( .B1(n21562), .B2(n21494), .A(n21553), .ZN(n21507) );
  NAND3_X1 U23203 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21480) );
  NAND2_X1 U23204 ( .A1(n21562), .A2(n21494), .ZN(n21479) );
  AOI22_X1 U23205 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n21652), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(n21651), .ZN(n21478) );
  OAI211_X1 U23206 ( .C1(n21480), .C2(n21479), .A(n21478), .B(n21616), .ZN(
        n21481) );
  INV_X1 U23207 ( .A(n21481), .ZN(n21487) );
  OAI22_X1 U23208 ( .A1(n21484), .A2(n21483), .B1(n21665), .B2(n21482), .ZN(
        n21485) );
  INV_X1 U23209 ( .A(n21485), .ZN(n21486) );
  OAI211_X1 U23210 ( .C1(n21488), .C2(n21507), .A(n21487), .B(n21486), .ZN(
        n21489) );
  INV_X1 U23211 ( .A(n21489), .ZN(n21492) );
  NAND2_X1 U23212 ( .A1(n21490), .A2(n21497), .ZN(n21491) );
  OAI211_X1 U23213 ( .C1(n21642), .C2(n21493), .A(n21492), .B(n21491), .ZN(
        P1_U2836) );
  NOR3_X1 U23214 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21494), .A3(n21539), .ZN(
        n21495) );
  AOI211_X1 U23215 ( .C1(n21652), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21457), .B(n21495), .ZN(n21504) );
  AOI22_X1 U23216 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n21651), .B1(n21628), .B2(
        n21496), .ZN(n21503) );
  NAND2_X1 U23217 ( .A1(n21498), .A2(n21497), .ZN(n21502) );
  INV_X1 U23218 ( .A(n21499), .ZN(n21500) );
  NAND2_X1 U23219 ( .A1(n21659), .A2(n21500), .ZN(n21501) );
  AND4_X1 U23220 ( .A1(n21504), .A2(n21503), .A3(n21502), .A4(n21501), .ZN(
        n21505) );
  OAI21_X1 U23221 ( .B1(n21507), .B2(n21506), .A(n21505), .ZN(P1_U2835) );
  AOI21_X1 U23222 ( .B1(n21508), .B2(n21562), .A(P1_REIP_REG_6__SCAN_IN), .ZN(
        n21517) );
  AOI21_X1 U23223 ( .B1(n21562), .B2(n21518), .A(n21553), .ZN(n21528) );
  OAI22_X1 U23224 ( .A1(n21510), .A2(n21570), .B1(n21665), .B2(n21509), .ZN(
        n21511) );
  AOI211_X1 U23225 ( .C1(n21651), .C2(P1_EBX_REG_6__SCAN_IN), .A(n21457), .B(
        n21511), .ZN(n21516) );
  INV_X1 U23226 ( .A(n21512), .ZN(n21513) );
  AOI22_X1 U23227 ( .A1(n21514), .A2(n21661), .B1(n21513), .B2(n21659), .ZN(
        n21515) );
  OAI211_X1 U23228 ( .C1(n21517), .C2(n21528), .A(n21516), .B(n21515), .ZN(
        P1_U2834) );
  NOR3_X1 U23229 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21518), .A3(n21539), .ZN(
        n21519) );
  AOI211_X1 U23230 ( .C1(n21652), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21457), .B(n21519), .ZN(n21523) );
  INV_X1 U23231 ( .A(n21520), .ZN(n21521) );
  AOI22_X1 U23232 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n21651), .B1(n21628), .B2(
        n21521), .ZN(n21522) );
  OAI211_X1 U23233 ( .C1(n21524), .C2(n21642), .A(n21523), .B(n21522), .ZN(
        n21525) );
  AOI21_X1 U23234 ( .B1(n21661), .B2(n21526), .A(n21525), .ZN(n21527) );
  OAI21_X1 U23235 ( .B1(n21529), .B2(n21528), .A(n21527), .ZN(P1_U2833) );
  AOI21_X1 U23236 ( .B1(n21530), .B2(n21562), .A(P1_REIP_REG_8__SCAN_IN), .ZN(
        n21538) );
  AOI21_X1 U23237 ( .B1(n21562), .B2(n21540), .A(n21553), .ZN(n21551) );
  OAI22_X1 U23238 ( .A1(n15245), .A2(n21570), .B1(n21665), .B2(n21531), .ZN(
        n21532) );
  AOI211_X1 U23239 ( .C1(n21651), .C2(P1_EBX_REG_8__SCAN_IN), .A(n21457), .B(
        n21532), .ZN(n21537) );
  INV_X1 U23240 ( .A(n21533), .ZN(n21535) );
  AOI22_X1 U23241 ( .A1(n21535), .A2(n21661), .B1(n21659), .B2(n21534), .ZN(
        n21536) );
  OAI211_X1 U23242 ( .C1(n21538), .C2(n21551), .A(n21537), .B(n21536), .ZN(
        P1_U2832) );
  NOR3_X1 U23243 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21540), .A3(n21539), .ZN(
        n21545) );
  AOI21_X1 U23244 ( .B1(n21652), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n21457), .ZN(n21542) );
  NAND2_X1 U23245 ( .A1(n21651), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n21541) );
  OAI211_X1 U23246 ( .C1(n21543), .C2(n21665), .A(n21542), .B(n21541), .ZN(
        n21544) );
  AOI211_X1 U23247 ( .C1(n21546), .C2(n21661), .A(n21545), .B(n21544), .ZN(
        n21547) );
  INV_X1 U23248 ( .A(n21547), .ZN(n21548) );
  AOI21_X1 U23249 ( .B1(n21549), .B2(n21659), .A(n21548), .ZN(n21550) );
  OAI21_X1 U23250 ( .B1(n21552), .B2(n21551), .A(n21550), .ZN(P1_U2831) );
  AND2_X1 U23251 ( .A1(n21553), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n21554) );
  AOI211_X1 U23252 ( .C1(n21652), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21457), .B(n21554), .ZN(n21557) );
  NAND2_X1 U23253 ( .A1(n21555), .A2(n21628), .ZN(n21556) );
  OAI211_X1 U23254 ( .C1(n21558), .C2(n21591), .A(n21557), .B(n21556), .ZN(
        n21559) );
  AOI21_X1 U23255 ( .B1(n21560), .B2(n21659), .A(n21559), .ZN(n21565) );
  OAI211_X1 U23256 ( .C1(n21563), .C2(P1_REIP_REG_10__SCAN_IN), .A(n21562), 
        .B(n21561), .ZN(n21564) );
  OAI211_X1 U23257 ( .C1(n21649), .C2(n21566), .A(n21565), .B(n21564), .ZN(
        P1_U2830) );
  OAI21_X1 U23258 ( .B1(n21576), .B2(n21567), .A(n21594), .ZN(n21579) );
  AOI21_X1 U23259 ( .B1(n21576), .B2(n21638), .A(n21579), .ZN(n21572) );
  AOI22_X1 U23260 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n21651), .B1(n21628), 
        .B2(n21568), .ZN(n21569) );
  OAI211_X1 U23261 ( .C1(n21570), .C2(n11870), .A(n21569), .B(n21616), .ZN(
        n21571) );
  AOI211_X1 U23262 ( .C1(n21573), .C2(n21661), .A(n21572), .B(n21571), .ZN(
        n21574) );
  OAI21_X1 U23263 ( .B1(n21575), .B2(n21642), .A(n21574), .ZN(P1_U2829) );
  NOR2_X1 U23264 ( .A1(n21576), .A2(n21638), .ZN(n21577) );
  AOI22_X1 U23265 ( .A1(n21628), .A2(n21578), .B1(n21577), .B2(n21580), .ZN(
        n21587) );
  OAI22_X1 U23266 ( .A1(n21581), .A2(n21649), .B1(n21580), .B2(n21579), .ZN(
        n21582) );
  AOI21_X1 U23267 ( .B1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n21652), .A(
        n21582), .ZN(n21586) );
  AOI22_X1 U23268 ( .A1(n21584), .A2(n21659), .B1(n21661), .B2(n21583), .ZN(
        n21585) );
  NAND4_X1 U23269 ( .A1(n21587), .A2(n21586), .A3(n21585), .A4(n21616), .ZN(
        P1_U2828) );
  AOI22_X1 U23270 ( .A1(n21588), .A2(n21659), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n21651), .ZN(n21590) );
  AOI21_X1 U23271 ( .B1(n21652), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21457), .ZN(n21589) );
  OAI211_X1 U23272 ( .C1(n21592), .C2(n21591), .A(n21590), .B(n21589), .ZN(
        n21593) );
  INV_X1 U23273 ( .A(n21593), .ZN(n21597) );
  OAI211_X1 U23274 ( .C1(n21595), .C2(P1_REIP_REG_15__SCAN_IN), .A(n21594), 
        .B(n21599), .ZN(n21596) );
  OAI211_X1 U23275 ( .C1(n21598), .C2(n21665), .A(n21597), .B(n21596), .ZN(
        P1_U2825) );
  OAI21_X1 U23276 ( .B1(n21601), .B2(n21600), .A(n21599), .ZN(n21604) );
  INV_X1 U23277 ( .A(n21602), .ZN(n21603) );
  NAND2_X1 U23278 ( .A1(n21604), .A2(n21603), .ZN(n21610) );
  INV_X1 U23279 ( .A(n21605), .ZN(n21608) );
  AOI22_X1 U23280 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21652), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(n21651), .ZN(n21606) );
  NAND2_X1 U23281 ( .A1(n21616), .A2(n21606), .ZN(n21607) );
  AOI21_X1 U23282 ( .B1(n21659), .B2(n21608), .A(n21607), .ZN(n21609) );
  NAND2_X1 U23283 ( .A1(n21610), .A2(n21609), .ZN(n21611) );
  AOI21_X1 U23284 ( .B1(n21612), .B2(n21661), .A(n21611), .ZN(n21613) );
  OAI21_X1 U23285 ( .B1(n21665), .B2(n21614), .A(n21613), .ZN(P1_U2824) );
  NAND2_X1 U23286 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n21652), .ZN(
        n21615) );
  OAI211_X1 U23287 ( .C1(n21642), .C2(n21617), .A(n21616), .B(n21615), .ZN(
        n21618) );
  AOI211_X1 U23288 ( .C1(n21651), .C2(P1_EBX_REG_18__SCAN_IN), .A(n21619), .B(
        n21618), .ZN(n21623) );
  AOI22_X1 U23289 ( .A1(n21621), .A2(n21661), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n21620), .ZN(n21622) );
  OAI211_X1 U23290 ( .C1(n21665), .C2(n21624), .A(n21623), .B(n21622), .ZN(
        P1_U2822) );
  AOI21_X1 U23291 ( .B1(n21626), .B2(n21625), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n21634) );
  AOI22_X1 U23292 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21652), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(n21651), .ZN(n21633) );
  INV_X1 U23293 ( .A(n21627), .ZN(n21629) );
  AOI222_X1 U23294 ( .A1(n21631), .A2(n21661), .B1(n21630), .B2(n21659), .C1(
        n21629), .C2(n21628), .ZN(n21632) );
  OAI211_X1 U23295 ( .C1(n21634), .C2(n21637), .A(n21633), .B(n21632), .ZN(
        P1_U2820) );
  AOI21_X1 U23296 ( .B1(n21637), .B2(n21636), .A(n21635), .ZN(n21641) );
  NOR3_X1 U23297 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n21639), .A3(n21638), 
        .ZN(n21640) );
  AOI211_X1 U23298 ( .C1(n21652), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n21641), .B(n21640), .ZN(n21648) );
  OAI22_X1 U23299 ( .A1(n21644), .A2(n21665), .B1(n21643), .B2(n21642), .ZN(
        n21645) );
  AOI21_X1 U23300 ( .B1(n21646), .B2(n21661), .A(n21645), .ZN(n21647) );
  OAI211_X1 U23301 ( .C1(n21650), .C2(n21649), .A(n21648), .B(n21647), .ZN(
        P1_U2818) );
  AOI22_X1 U23302 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21652), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(n21651), .ZN(n21653) );
  INV_X1 U23303 ( .A(n21653), .ZN(n21654) );
  AOI221_X1 U23304 ( .B1(n21657), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n21656), 
        .C2(n21655), .A(n21654), .ZN(n21664) );
  INV_X1 U23305 ( .A(n21658), .ZN(n21660) );
  AOI22_X1 U23306 ( .A1(n21662), .A2(n21661), .B1(n21660), .B2(n21659), .ZN(
        n21663) );
  OAI211_X1 U23307 ( .C1(n21666), .C2(n21665), .A(n21664), .B(n21663), .ZN(
        P1_U2816) );
  OAI21_X1 U23308 ( .B1(n21669), .B2(n21668), .A(n21667), .ZN(P1_U2806) );
  INV_X1 U23309 ( .A(n21670), .ZN(n21672) );
  OAI22_X1 U23310 ( .A1(n21674), .A2(n21673), .B1(n21672), .B2(n21671), .ZN(
        n21676) );
  MUX2_X1 U23311 ( .A(n21676), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21675), .Z(P1_U3469) );
  AOI21_X1 U23312 ( .B1(n21679), .B2(n21678), .A(n21677), .ZN(n21681) );
  OAI211_X1 U23313 ( .C1(n21684), .C2(n22008), .A(n21681), .B(n21680), .ZN(
        P1_U3163) );
  OAI22_X1 U23314 ( .A1(n21684), .A2(n21930), .B1(n21683), .B2(n21682), .ZN(
        P1_U3466) );
  AOI21_X1 U23315 ( .B1(n21687), .B2(n21686), .A(n21685), .ZN(n21688) );
  OAI22_X1 U23316 ( .A1(n21690), .A2(n21689), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21688), .ZN(n21691) );
  OAI21_X1 U23317 ( .B1(n21693), .B2(n21692), .A(n21691), .ZN(P1_U3161) );
  OAI21_X1 U23318 ( .B1(n21696), .B2(n21936), .A(n21694), .ZN(P1_U2805) );
  INV_X1 U23319 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21695) );
  OAI21_X1 U23320 ( .B1(n21696), .B2(n21695), .A(n21694), .ZN(P1_U3465) );
  INV_X1 U23321 ( .A(n21697), .ZN(n21699) );
  OAI21_X1 U23322 ( .B1(n21701), .B2(n21698), .A(n21699), .ZN(P2_U2818) );
  OAI21_X1 U23323 ( .B1(n21701), .B2(n21700), .A(n21699), .ZN(P2_U3592) );
  INV_X1 U23324 ( .A(n21702), .ZN(n21704) );
  OAI21_X1 U23325 ( .B1(n21706), .B2(n21703), .A(n21704), .ZN(P3_U2636) );
  OAI21_X1 U23326 ( .B1(n21706), .B2(n21705), .A(n21704), .ZN(P3_U3281) );
  INV_X1 U23327 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21707) );
  AOI21_X1 U23328 ( .B1(HOLD), .B2(n21708), .A(n21707), .ZN(n21712) );
  AOI21_X1 U23329 ( .B1(n21710), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21709), 
        .ZN(n21772) );
  OAI21_X1 U23330 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21768), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n21771) );
  INV_X1 U23331 ( .A(n21771), .ZN(n21711) );
  OAI22_X1 U23332 ( .A1(n21713), .A2(n21712), .B1(n21772), .B2(n21711), .ZN(
        P3_U3029) );
  INV_X1 U23333 ( .A(HOLD), .ZN(n21766) );
  OAI21_X1 U23334 ( .B1(NA), .B2(n21716), .A(n21724), .ZN(n21714) );
  OAI211_X1 U23335 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21723), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n21714), .ZN(n21721) );
  AOI211_X1 U23336 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21723), .A(NA), .B(
        n21715), .ZN(n21718) );
  NOR2_X1 U23337 ( .A1(n21722), .A2(n21716), .ZN(n21717) );
  INV_X1 U23338 ( .A(n21717), .ZN(n21725) );
  NAND2_X1 U23339 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21725), .ZN(n21728) );
  OAI221_X1 U23340 ( .B1(n21718), .B2(n21717), .C1(n21718), .C2(
        P1_STATE_REG_2__SCAN_IN), .A(n21728), .ZN(n21719) );
  OAI211_X1 U23341 ( .C1(n21766), .C2(n21721), .A(n21720), .B(n21719), .ZN(
        P1_U3196) );
  NOR2_X1 U23342 ( .A1(n21722), .A2(n21766), .ZN(n21731) );
  AOI21_X1 U23343 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21723), .ZN(
        n21729) );
  AOI22_X1 U23344 ( .A1(n21724), .A2(n21731), .B1(P1_STATE_REG_0__SCAN_IN), 
        .B2(n21729), .ZN(n21727) );
  NAND3_X1 U23345 ( .A1(n21727), .A2(n21726), .A3(n21725), .ZN(P1_U3195) );
  INV_X1 U23346 ( .A(n21728), .ZN(n21734) );
  INV_X1 U23347 ( .A(n21729), .ZN(n21730) );
  AOI211_X1 U23348 ( .C1(NA), .C2(n21732), .A(n21731), .B(n21730), .ZN(n21733)
         );
  OAI22_X1 U23349 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21734), .B1(n22339), 
        .B2(n21733), .ZN(P1_U3194) );
  NOR2_X1 U23350 ( .A1(n21735), .A2(n21746), .ZN(n21747) );
  OR2_X1 U23351 ( .A1(n21755), .A2(n21747), .ZN(n21748) );
  AOI22_X1 U23352 ( .A1(NA), .A2(n21749), .B1(n21752), .B2(n21748), .ZN(n21738) );
  OAI211_X1 U23353 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(P2_STATE_REG_1__SCAN_IN), .A(HOLD), .B(n21736), .ZN(n21737) );
  OAI211_X1 U23354 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21739), .A(
        n21738), .B(n21737), .ZN(P2_U3209) );
  NOR2_X1 U23355 ( .A1(HOLD), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21754)
         );
  INV_X1 U23356 ( .A(n21754), .ZN(n21741) );
  AOI211_X1 U23357 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21755), .B(
        n21745), .ZN(n21740) );
  AOI211_X1 U23358 ( .C1(n21742), .C2(n21741), .A(n21747), .B(n21740), .ZN(
        n21743) );
  NAND2_X1 U23359 ( .A1(n21744), .A2(n21743), .ZN(P2_U3210) );
  AOI22_X1 U23360 ( .A1(n21747), .A2(n21768), .B1(n21746), .B2(n21745), .ZN(
        n21753) );
  NOR2_X1 U23361 ( .A1(HOLD), .A2(n21748), .ZN(n21751) );
  AND2_X1 U23362 ( .A1(n21749), .A2(NA), .ZN(n21750) );
  OAI33_X1 U23363 ( .A1(n21755), .A2(n21754), .A3(n21753), .B1(n21752), .B2(
        n21751), .B3(n21750), .ZN(P2_U3211) );
  NOR2_X1 U23364 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21774)
         );
  OAI21_X1 U23365 ( .B1(n21767), .B2(n21766), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21758) );
  NOR2_X1 U23366 ( .A1(n21764), .A2(n21756), .ZN(n21769) );
  INV_X1 U23367 ( .A(n21769), .ZN(n21757) );
  OAI21_X1 U23368 ( .B1(n21774), .B2(n21758), .A(n21757), .ZN(n21761) );
  OAI211_X1 U23369 ( .C1(n21767), .C2(n21766), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21759) );
  AOI21_X1 U23370 ( .B1(n21759), .B2(n21762), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21760) );
  AOI21_X1 U23371 ( .B1(n21762), .B2(n21761), .A(n21760), .ZN(n21763) );
  OAI221_X1 U23372 ( .B1(n21765), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n21765), 
        .C2(n21764), .A(n21763), .ZN(P3_U3030) );
  OAI22_X1 U23373 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21767), .B2(n21766), .ZN(n21770)
         );
  OAI221_X1 U23374 ( .B1(n21770), .B2(n21769), .C1(n21770), .C2(n21768), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21773) );
  OAI22_X1 U23375 ( .A1(n21774), .A2(n21773), .B1(n21772), .B2(n21771), .ZN(
        P3_U3031) );
  NOR2_X1 U23376 ( .A1(n21857), .A2(n21775), .ZN(n21778) );
  AOI21_X1 U23377 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n21858), .A(n21778), 
        .ZN(n21776) );
  OAI21_X1 U23378 ( .B1(n21777), .B2(n21863), .A(n21776), .ZN(P1_U2937) );
  AOI21_X1 U23379 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n21858), .A(n21778), 
        .ZN(n21779) );
  OAI21_X1 U23380 ( .B1(n21780), .B2(n21863), .A(n21779), .ZN(P1_U2952) );
  NOR2_X1 U23381 ( .A1(n21857), .A2(n21781), .ZN(n21784) );
  AOI21_X1 U23382 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n21858), .A(n21784), 
        .ZN(n21782) );
  OAI21_X1 U23383 ( .B1(n21783), .B2(n21863), .A(n21782), .ZN(P1_U2938) );
  AOI21_X1 U23384 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n21858), .A(n21784), 
        .ZN(n21785) );
  OAI21_X1 U23385 ( .B1(n21786), .B2(n21863), .A(n21785), .ZN(P1_U2953) );
  NOR2_X1 U23386 ( .A1(n21857), .A2(n21787), .ZN(n21790) );
  AOI21_X1 U23387 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n21858), .A(n21790), 
        .ZN(n21788) );
  OAI21_X1 U23388 ( .B1(n21789), .B2(n21863), .A(n21788), .ZN(P1_U2939) );
  AOI21_X1 U23389 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n21858), .A(n21790), 
        .ZN(n21791) );
  OAI21_X1 U23390 ( .B1(n21792), .B2(n21863), .A(n21791), .ZN(P1_U2954) );
  NOR2_X1 U23391 ( .A1(n21857), .A2(n21793), .ZN(n21796) );
  AOI21_X1 U23392 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n21858), .A(n21796), 
        .ZN(n21794) );
  OAI21_X1 U23393 ( .B1(n21795), .B2(n21863), .A(n21794), .ZN(P1_U2940) );
  AOI21_X1 U23394 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n21858), .A(n21796), 
        .ZN(n21797) );
  OAI21_X1 U23395 ( .B1(n21798), .B2(n21863), .A(n21797), .ZN(P1_U2955) );
  NOR2_X1 U23396 ( .A1(n21857), .A2(n21799), .ZN(n21802) );
  AOI21_X1 U23397 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n21858), .A(n21802), 
        .ZN(n21800) );
  OAI21_X1 U23398 ( .B1(n12026), .B2(n21863), .A(n21800), .ZN(P1_U2941) );
  AOI21_X1 U23399 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n21843), .A(n21802), 
        .ZN(n21803) );
  OAI21_X1 U23400 ( .B1(n21804), .B2(n21863), .A(n21803), .ZN(P1_U2956) );
  INV_X1 U23401 ( .A(n21805), .ZN(n21806) );
  NOR2_X1 U23402 ( .A1(n21857), .A2(n21806), .ZN(n21809) );
  AOI21_X1 U23403 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n21843), .A(n21809), 
        .ZN(n21807) );
  OAI21_X1 U23404 ( .B1(n21808), .B2(n21863), .A(n21807), .ZN(P1_U2942) );
  AOI21_X1 U23405 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n21843), .A(n21809), 
        .ZN(n21810) );
  OAI21_X1 U23406 ( .B1(n21811), .B2(n21863), .A(n21810), .ZN(P1_U2957) );
  NOR2_X1 U23407 ( .A1(n21857), .A2(n21812), .ZN(n21814) );
  AOI21_X1 U23408 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n21843), .A(n21814), 
        .ZN(n21813) );
  OAI21_X1 U23409 ( .B1(n12064), .B2(n21863), .A(n21813), .ZN(P1_U2943) );
  AOI21_X1 U23410 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n21843), .A(n21814), 
        .ZN(n21815) );
  OAI21_X1 U23411 ( .B1(n11794), .B2(n21863), .A(n21815), .ZN(P1_U2958) );
  NOR2_X1 U23412 ( .A1(n21857), .A2(n21816), .ZN(n21819) );
  AOI21_X1 U23413 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n21843), .A(n21819), 
        .ZN(n21817) );
  OAI21_X1 U23414 ( .B1(n21818), .B2(n21863), .A(n21817), .ZN(P1_U2944) );
  AOI21_X1 U23415 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n21843), .A(n21819), 
        .ZN(n21820) );
  OAI21_X1 U23416 ( .B1(n11816), .B2(n21863), .A(n21820), .ZN(P1_U2959) );
  NOR2_X1 U23417 ( .A1(n21857), .A2(n21821), .ZN(n21824) );
  AOI21_X1 U23418 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21843), .A(n21824), 
        .ZN(n21822) );
  OAI21_X1 U23419 ( .B1(n21823), .B2(n21863), .A(n21822), .ZN(P1_U2945) );
  AOI21_X1 U23420 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21843), .A(n21824), 
        .ZN(n21825) );
  OAI21_X1 U23421 ( .B1(n15032), .B2(n21863), .A(n21825), .ZN(P1_U2960) );
  NOR2_X1 U23422 ( .A1(n21857), .A2(n21826), .ZN(n21829) );
  AOI21_X1 U23423 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n21858), .A(n21829), 
        .ZN(n21827) );
  OAI21_X1 U23424 ( .B1(n21828), .B2(n21863), .A(n21827), .ZN(P1_U2946) );
  AOI21_X1 U23425 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n21843), .A(n21829), 
        .ZN(n21830) );
  OAI21_X1 U23426 ( .B1(n15018), .B2(n21863), .A(n21830), .ZN(P1_U2961) );
  INV_X1 U23427 ( .A(n21831), .ZN(n21832) );
  NOR2_X1 U23428 ( .A1(n21857), .A2(n21832), .ZN(n21835) );
  AOI21_X1 U23429 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21843), .A(n21835), 
        .ZN(n21833) );
  OAI21_X1 U23430 ( .B1(n21834), .B2(n21863), .A(n21833), .ZN(P1_U2947) );
  AOI21_X1 U23431 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n21843), .A(n21835), 
        .ZN(n21836) );
  OAI21_X1 U23432 ( .B1(n21837), .B2(n21863), .A(n21836), .ZN(P1_U2962) );
  NOR2_X1 U23433 ( .A1(n21857), .A2(n21838), .ZN(n21840) );
  AOI21_X1 U23434 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21843), .A(n21840), 
        .ZN(n21839) );
  OAI21_X1 U23435 ( .B1(n12162), .B2(n21863), .A(n21839), .ZN(P1_U2948) );
  AOI21_X1 U23436 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n21843), .A(n21840), 
        .ZN(n21841) );
  OAI21_X1 U23437 ( .B1(n15205), .B2(n21863), .A(n21841), .ZN(P1_U2963) );
  NOR2_X1 U23438 ( .A1(n21857), .A2(n21842), .ZN(n21846) );
  AOI21_X1 U23439 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21843), .A(n21846), 
        .ZN(n21844) );
  OAI21_X1 U23440 ( .B1(n21845), .B2(n21863), .A(n21844), .ZN(P1_U2949) );
  AOI21_X1 U23441 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n21843), .A(n21846), 
        .ZN(n21847) );
  OAI21_X1 U23442 ( .B1(n15226), .B2(n21863), .A(n21847), .ZN(P1_U2964) );
  INV_X1 U23443 ( .A(n21848), .ZN(n21849) );
  NOR2_X1 U23444 ( .A1(n21857), .A2(n21849), .ZN(n21852) );
  AOI21_X1 U23445 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21858), .A(n21852), 
        .ZN(n21850) );
  OAI21_X1 U23446 ( .B1(n21851), .B2(n21863), .A(n21850), .ZN(P1_U2950) );
  AOI21_X1 U23447 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n21843), .A(n21852), 
        .ZN(n21853) );
  OAI21_X1 U23448 ( .B1(n21854), .B2(n21863), .A(n21853), .ZN(P1_U2965) );
  INV_X1 U23449 ( .A(n21855), .ZN(n21856) );
  NOR2_X1 U23450 ( .A1(n21857), .A2(n21856), .ZN(n21861) );
  AOI21_X1 U23451 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n21858), .A(n21861), 
        .ZN(n21859) );
  OAI21_X1 U23452 ( .B1(n21860), .B2(n21863), .A(n21859), .ZN(P1_U2951) );
  AOI21_X1 U23453 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n21843), .A(n21861), 
        .ZN(n21862) );
  OAI21_X1 U23454 ( .B1(n21864), .B2(n21863), .A(n21862), .ZN(P1_U2966) );
  INV_X1 U23455 ( .A(n21866), .ZN(n21867) );
  NAND3_X1 U23456 ( .A1(n21876), .A2(n21982), .A3(n22247), .ZN(n21869) );
  NOR2_X1 U23457 ( .A1(n22015), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21979) );
  INV_X1 U23458 ( .A(n21979), .ZN(n21868) );
  NAND2_X1 U23459 ( .A1(n21869), .A2(n21868), .ZN(n21874) );
  OR2_X1 U23460 ( .A1(n21961), .A2(n14445), .ZN(n21899) );
  NOR2_X1 U23461 ( .A1(n21899), .A2(n21962), .ZN(n21872) );
  NAND3_X1 U23462 ( .A1(n21965), .A2(n21922), .A3(n12217), .ZN(n21880) );
  OR2_X1 U23463 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21880), .ZN(
        n22246) );
  OAI22_X1 U23464 ( .A1(n22247), .A2(n22022), .B1(n21966), .B2(n22246), .ZN(
        n21870) );
  INV_X1 U23465 ( .A(n21870), .ZN(n21878) );
  NOR2_X1 U23466 ( .A1(n21991), .A2(n21871), .ZN(n21952) );
  INV_X1 U23467 ( .A(n21872), .ZN(n21873) );
  AOI22_X1 U23468 ( .A1(n21874), .A2(n21873), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22246), .ZN(n21875) );
  OAI211_X1 U23469 ( .C1(n11391), .C2(n22008), .A(n21952), .B(n21875), .ZN(
        n22249) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22019), .ZN(n21877) );
  OAI211_X1 U23471 ( .C1(n22252), .C2(n21974), .A(n21878), .B(n21877), .ZN(
        P1_U3033) );
  OR2_X1 U23472 ( .A1(n14520), .A2(n11020), .ZN(n21983) );
  INV_X1 U23473 ( .A(n21899), .ZN(n21879) );
  NOR2_X1 U23474 ( .A1(n21975), .A2(n21880), .ZN(n22253) );
  AOI21_X1 U23475 ( .B1(n21879), .B2(n21976), .A(n22253), .ZN(n21881) );
  OAI22_X1 U23476 ( .A1(n21881), .A2(n22015), .B1(n21880), .B2(n22008), .ZN(
        n22254) );
  AOI22_X1 U23477 ( .A1(n22254), .A2(n22011), .B1(n22010), .B2(n22253), .ZN(
        n21885) );
  INV_X1 U23478 ( .A(n21880), .ZN(n21883) );
  OAI211_X1 U23479 ( .C1(n21894), .C2(n21936), .A(n21982), .B(n21881), .ZN(
        n21882) );
  OAI211_X1 U23480 ( .C1(n21982), .C2(n21883), .A(n22017), .B(n21882), .ZN(
        n22256) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22000), .ZN(n21884) );
  OAI211_X1 U23482 ( .C1(n22003), .C2(n22259), .A(n21885), .B(n21884), .ZN(
        P1_U3041) );
  NOR3_X1 U23483 ( .A1(n22263), .A2(n22271), .A3(n22015), .ZN(n21886) );
  NOR2_X1 U23484 ( .A1(n21886), .A2(n21979), .ZN(n21891) );
  INV_X1 U23485 ( .A(n21891), .ZN(n21887) );
  NOR2_X1 U23486 ( .A1(n21899), .A2(n14973), .ZN(n21890) );
  NOR2_X1 U23487 ( .A1(n21923), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21911) );
  NAND3_X1 U23488 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21922), .A3(
        n12217), .ZN(n21897) );
  OR2_X1 U23489 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21897), .ZN(
        n22260) );
  OAI22_X1 U23490 ( .A1(n22261), .A2(n22003), .B1(n21966), .B2(n22260), .ZN(
        n21888) );
  INV_X1 U23491 ( .A(n21888), .ZN(n21893) );
  NOR2_X1 U23492 ( .A1(n21911), .A2(n22008), .ZN(n21914) );
  AOI21_X1 U23493 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22260), .A(n21914), 
        .ZN(n21889) );
  OAI211_X1 U23494 ( .C1(n21891), .C2(n21890), .A(n21952), .B(n21889), .ZN(
        n22264) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22000), .ZN(n21892) );
  OAI211_X1 U23496 ( .C1(n22267), .C2(n21974), .A(n21893), .B(n21892), .ZN(
        P1_U3049) );
  INV_X1 U23497 ( .A(n21897), .ZN(n21902) );
  INV_X1 U23498 ( .A(n21894), .ZN(n21896) );
  OAI21_X1 U23499 ( .B1(n21896), .B2(n22015), .A(n21895), .ZN(n21905) );
  OR2_X1 U23500 ( .A1(n21975), .A2(n21897), .ZN(n22268) );
  OAI21_X1 U23501 ( .B1(n21899), .B2(n21898), .A(n22268), .ZN(n21901) );
  AOI22_X1 U23502 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21902), .B1(n21905), 
        .B2(n21901), .ZN(n22275) );
  OAI22_X1 U23503 ( .A1(n22261), .A2(n22022), .B1(n21966), .B2(n22268), .ZN(
        n21900) );
  INV_X1 U23504 ( .A(n21900), .ZN(n21908) );
  INV_X1 U23505 ( .A(n21901), .ZN(n21904) );
  OAI21_X1 U23506 ( .B1(n21982), .B2(n21902), .A(n22017), .ZN(n21903) );
  AOI21_X1 U23507 ( .B1(n21905), .B2(n21904), .A(n21903), .ZN(n21906) );
  INV_X1 U23508 ( .A(n22269), .ZN(n22069) );
  AOI22_X1 U23509 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22069), .B2(n22019), .ZN(n21907) );
  OAI211_X1 U23510 ( .C1(n22275), .C2(n21974), .A(n21908), .B(n21907), .ZN(
        P1_U3057) );
  NOR2_X1 U23511 ( .A1(n22279), .A2(n22015), .ZN(n21909) );
  AOI21_X1 U23512 ( .B1(n21909), .B2(n22277), .A(n21979), .ZN(n21917) );
  INV_X1 U23513 ( .A(n21917), .ZN(n21912) );
  OR3_X1 U23514 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n22007), .ZN(n22276) );
  OAI22_X1 U23515 ( .A1(n22277), .A2(n22022), .B1(n21966), .B2(n22276), .ZN(
        n21913) );
  INV_X1 U23516 ( .A(n21913), .ZN(n21919) );
  AOI21_X1 U23517 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22276), .A(n21914), 
        .ZN(n21915) );
  OAI211_X1 U23518 ( .C1(n21917), .C2(n21916), .A(n21998), .B(n21915), .ZN(
        n22280) );
  AOI22_X1 U23519 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22019), .B2(n22279), .ZN(n21918) );
  OAI211_X1 U23520 ( .C1(n22283), .C2(n21974), .A(n21919), .B(n21918), .ZN(
        P1_U3081) );
  NAND3_X1 U23521 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21965), .A3(
        n21922), .ZN(n21933) );
  NOR2_X1 U23522 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21933), .ZN(
        n22284) );
  AOI21_X1 U23523 ( .B1(n21943), .B2(n14973), .A(n22284), .ZN(n21927) );
  NAND2_X1 U23524 ( .A1(n21924), .A2(n21923), .ZN(n21968) );
  INV_X1 U23525 ( .A(n21945), .ZN(n21925) );
  OAI22_X1 U23526 ( .A1(n21927), .A2(n22015), .B1(n21968), .B2(n21925), .ZN(
        n22285) );
  AOI22_X1 U23527 ( .A1(n22285), .A2(n22011), .B1(n22010), .B2(n22284), .ZN(
        n21932) );
  INV_X1 U23528 ( .A(n22295), .ZN(n21926) );
  OAI21_X1 U23529 ( .B1(n21926), .B2(n22286), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21928) );
  NAND2_X1 U23530 ( .A1(n21928), .A2(n21927), .ZN(n21929) );
  AOI22_X1 U23531 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22000), .B2(n22286), .ZN(n21931) );
  OAI211_X1 U23532 ( .C1(n22003), .C2(n22295), .A(n21932), .B(n21931), .ZN(
        P1_U3097) );
  NOR2_X1 U23533 ( .A1(n21975), .A2(n21933), .ZN(n22290) );
  AOI21_X1 U23534 ( .B1(n21943), .B2(n21976), .A(n22290), .ZN(n21934) );
  OAI22_X1 U23535 ( .A1(n21934), .A2(n22015), .B1(n21933), .B2(n22008), .ZN(
        n22291) );
  AOI22_X1 U23536 ( .A1(n22291), .A2(n22011), .B1(n22010), .B2(n22290), .ZN(
        n21941) );
  INV_X1 U23537 ( .A(n21933), .ZN(n21938) );
  OAI211_X1 U23538 ( .C1(n21939), .C2(n21936), .A(n21935), .B(n21934), .ZN(
        n21937) );
  OAI211_X1 U23539 ( .C1(n21982), .C2(n21938), .A(n22017), .B(n21937), .ZN(
        n22292) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22019), .ZN(n21940) );
  OAI211_X1 U23541 ( .C1(n22022), .C2(n22295), .A(n21941), .B(n21940), .ZN(
        P1_U3105) );
  NOR3_X1 U23542 ( .A1(n22298), .A2(n22297), .A3(n22015), .ZN(n21942) );
  NOR2_X1 U23543 ( .A1(n21942), .A2(n21979), .ZN(n21954) );
  INV_X1 U23544 ( .A(n21954), .ZN(n21946) );
  NAND2_X1 U23545 ( .A1(n21944), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21948) );
  INV_X1 U23546 ( .A(n21948), .ZN(n21992) );
  NOR2_X1 U23547 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21947), .ZN(
        n22296) );
  AOI22_X1 U23548 ( .A1(n22298), .A2(n22000), .B1(n22010), .B2(n22296), .ZN(
        n21956) );
  INV_X1 U23549 ( .A(n22296), .ZN(n21950) );
  NAND2_X1 U23550 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21948), .ZN(n21997) );
  INV_X1 U23551 ( .A(n21997), .ZN(n21949) );
  AOI21_X1 U23552 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21950), .A(n21949), 
        .ZN(n21951) );
  OAI211_X1 U23553 ( .C1(n21954), .C2(n21953), .A(n21952), .B(n21951), .ZN(
        n22299) );
  AOI22_X1 U23554 ( .A1(n22299), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22019), .B2(n22297), .ZN(n21955) );
  OAI211_X1 U23555 ( .C1(n22302), .C2(n21974), .A(n21956), .B(n21955), .ZN(
        P1_U3113) );
  INV_X1 U23556 ( .A(n22317), .ZN(n21958) );
  NOR3_X1 U23557 ( .A1(n22306), .A2(n21958), .A3(n22015), .ZN(n21959) );
  NOR2_X1 U23558 ( .A1(n21959), .A2(n21979), .ZN(n21971) );
  INV_X1 U23559 ( .A(n21971), .ZN(n21964) );
  NAND2_X1 U23560 ( .A1(n21961), .A2(n21960), .ZN(n21990) );
  NOR2_X1 U23561 ( .A1(n21990), .A2(n21962), .ZN(n21970) );
  INV_X1 U23562 ( .A(n21968), .ZN(n21963) );
  NAND3_X1 U23563 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21965), .ZN(n21977) );
  OR2_X1 U23564 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21977), .ZN(
        n22303) );
  OAI22_X1 U23565 ( .A1(n22317), .A2(n22003), .B1(n21966), .B2(n22303), .ZN(
        n21967) );
  INV_X1 U23566 ( .A(n21967), .ZN(n21973) );
  AOI22_X1 U23567 ( .A1(n21968), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22303), .ZN(n21969) );
  OAI211_X1 U23568 ( .C1(n21971), .C2(n21970), .A(n21998), .B(n21969), .ZN(
        n22307) );
  AOI22_X1 U23569 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22000), .B2(n22306), .ZN(n21972) );
  OAI211_X1 U23570 ( .C1(n22311), .C2(n21974), .A(n21973), .B(n21972), .ZN(
        P1_U3129) );
  NOR2_X1 U23571 ( .A1(n21975), .A2(n21977), .ZN(n22313) );
  INV_X1 U23572 ( .A(n21990), .ZN(n22006) );
  AOI21_X1 U23573 ( .B1(n22006), .B2(n21976), .A(n22313), .ZN(n21978) );
  OAI22_X1 U23574 ( .A1(n21978), .A2(n22015), .B1(n21977), .B2(n22008), .ZN(
        n22312) );
  AOI22_X1 U23575 ( .A1(n22010), .A2(n22313), .B1(n22312), .B2(n22011), .ZN(
        n21986) );
  INV_X1 U23576 ( .A(n21977), .ZN(n21981) );
  OAI21_X1 U23577 ( .B1(n21984), .B2(n21979), .A(n21978), .ZN(n21980) );
  OAI211_X1 U23578 ( .C1(n21982), .C2(n21981), .A(n22017), .B(n21980), .ZN(
        n22314) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22019), .ZN(n21985) );
  OAI211_X1 U23580 ( .C1(n22022), .C2(n22317), .A(n21986), .B(n21985), .ZN(
        P1_U3137) );
  INV_X1 U23581 ( .A(n21987), .ZN(n21988) );
  NOR3_X2 U23582 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22007), .A3(
        n12217), .ZN(n22319) );
  OR2_X1 U23583 ( .A1(n21990), .A2(n14973), .ZN(n21995) );
  NAND2_X1 U23584 ( .A1(n21992), .A2(n21991), .ZN(n21993) );
  OAI21_X1 U23585 ( .B1(n21995), .B2(n22015), .A(n21993), .ZN(n22318) );
  AOI22_X1 U23586 ( .A1(n22010), .A2(n22319), .B1(n22011), .B2(n22318), .ZN(
        n22002) );
  INV_X1 U23587 ( .A(n22335), .ZN(n21994) );
  OAI21_X1 U23588 ( .B1(n21994), .B2(n22321), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21996) );
  AOI21_X1 U23589 ( .B1(n21996), .B2(n21995), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21999) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22000), .ZN(n22001) );
  OAI211_X1 U23591 ( .C1(n22003), .C2(n22335), .A(n22002), .B(n22001), .ZN(
        P1_U3145) );
  NOR2_X1 U23592 ( .A1(n22004), .A2(n12217), .ZN(n22326) );
  AOI21_X1 U23593 ( .B1(n22006), .B2(n22005), .A(n22326), .ZN(n22012) );
  NOR2_X1 U23594 ( .A1(n22007), .A2(n12217), .ZN(n22018) );
  INV_X1 U23595 ( .A(n22018), .ZN(n22009) );
  OAI22_X1 U23596 ( .A1(n22012), .A2(n22015), .B1(n22009), .B2(n22008), .ZN(
        n22328) );
  AOI22_X1 U23597 ( .A1(n22011), .A2(n22328), .B1(n22010), .B2(n22326), .ZN(
        n22021) );
  NAND2_X1 U23598 ( .A1(n22013), .A2(n22012), .ZN(n22014) );
  OR2_X1 U23599 ( .A1(n22015), .A2(n22014), .ZN(n22016) );
  OAI211_X1 U23600 ( .C1(n21982), .C2(n22018), .A(n22017), .B(n22016), .ZN(
        n22330) );
  AOI22_X1 U23601 ( .A1(n22019), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n22020) );
  OAI211_X1 U23602 ( .C1(n22022), .C2(n22335), .A(n22021), .B(n22020), .ZN(
        P1_U3153) );
  OAI22_X1 U23603 ( .A1(n22247), .A2(n22059), .B1(n22043), .B2(n22246), .ZN(
        n22023) );
  INV_X1 U23604 ( .A(n22023), .ZN(n22025) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22056), .ZN(n22024) );
  OAI211_X1 U23606 ( .C1(n22252), .C2(n22047), .A(n22025), .B(n22024), .ZN(
        P1_U3034) );
  AOI22_X1 U23607 ( .A1(n22254), .A2(n22055), .B1(n22054), .B2(n22253), .ZN(
        n22027) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22050), .ZN(n22026) );
  OAI211_X1 U23609 ( .C1(n22053), .C2(n22259), .A(n22027), .B(n22026), .ZN(
        P1_U3042) );
  OAI22_X1 U23610 ( .A1(n22261), .A2(n22053), .B1(n22043), .B2(n22260), .ZN(
        n22028) );
  INV_X1 U23611 ( .A(n22028), .ZN(n22030) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22050), .ZN(n22029) );
  OAI211_X1 U23613 ( .C1(n22267), .C2(n22047), .A(n22030), .B(n22029), .ZN(
        P1_U3050) );
  OAI22_X1 U23614 ( .A1(n22261), .A2(n22059), .B1(n22043), .B2(n22268), .ZN(
        n22031) );
  INV_X1 U23615 ( .A(n22031), .ZN(n22033) );
  AOI22_X1 U23616 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22069), .B2(n22056), .ZN(n22032) );
  OAI211_X1 U23617 ( .C1(n22275), .C2(n22047), .A(n22033), .B(n22032), .ZN(
        P1_U3058) );
  OAI22_X1 U23618 ( .A1(n22277), .A2(n22059), .B1(n22043), .B2(n22276), .ZN(
        n22034) );
  INV_X1 U23619 ( .A(n22034), .ZN(n22036) );
  AOI22_X1 U23620 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22056), .B2(n22279), .ZN(n22035) );
  OAI211_X1 U23621 ( .C1(n22283), .C2(n22047), .A(n22036), .B(n22035), .ZN(
        P1_U3082) );
  AOI22_X1 U23622 ( .A1(n22285), .A2(n22055), .B1(n22054), .B2(n22284), .ZN(
        n22038) );
  AOI22_X1 U23623 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22050), .B2(n22286), .ZN(n22037) );
  OAI211_X1 U23624 ( .C1(n22053), .C2(n22295), .A(n22038), .B(n22037), .ZN(
        P1_U3098) );
  AOI22_X1 U23625 ( .A1(n22291), .A2(n22055), .B1(n22054), .B2(n22290), .ZN(
        n22040) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22056), .ZN(n22039) );
  OAI211_X1 U23627 ( .C1(n22059), .C2(n22295), .A(n22040), .B(n22039), .ZN(
        P1_U3106) );
  AOI22_X1 U23628 ( .A1(n22297), .A2(n22056), .B1(n22054), .B2(n22296), .ZN(
        n22042) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22299), .B1(
        n22298), .B2(n22050), .ZN(n22041) );
  OAI211_X1 U23630 ( .C1(n22302), .C2(n22047), .A(n22042), .B(n22041), .ZN(
        P1_U3114) );
  OAI22_X1 U23631 ( .A1(n22317), .A2(n22053), .B1(n22043), .B2(n22303), .ZN(
        n22044) );
  INV_X1 U23632 ( .A(n22044), .ZN(n22046) );
  AOI22_X1 U23633 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22050), .B2(n22306), .ZN(n22045) );
  OAI211_X1 U23634 ( .C1(n22311), .C2(n22047), .A(n22046), .B(n22045), .ZN(
        P1_U3130) );
  AOI22_X1 U23635 ( .A1(n22054), .A2(n22313), .B1(n22312), .B2(n22055), .ZN(
        n22049) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22056), .ZN(n22048) );
  OAI211_X1 U23637 ( .C1(n22059), .C2(n22317), .A(n22049), .B(n22048), .ZN(
        P1_U3138) );
  AOI22_X1 U23638 ( .A1(n22054), .A2(n22319), .B1(n22055), .B2(n22318), .ZN(
        n22052) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22050), .ZN(n22051) );
  OAI211_X1 U23640 ( .C1(n22053), .C2(n22335), .A(n22052), .B(n22051), .ZN(
        P1_U3146) );
  AOI22_X1 U23641 ( .A1(n22055), .A2(n22328), .B1(n22054), .B2(n22326), .ZN(
        n22058) );
  AOI22_X1 U23642 ( .A1(n22056), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n22057) );
  OAI211_X1 U23643 ( .C1(n22059), .C2(n22335), .A(n22058), .B(n22057), .ZN(
        P1_U3154) );
  OAI22_X1 U23644 ( .A1(n22247), .A2(n22097), .B1(n22081), .B2(n22246), .ZN(
        n22060) );
  INV_X1 U23645 ( .A(n22060), .ZN(n22062) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22094), .ZN(n22061) );
  OAI211_X1 U23647 ( .C1(n22252), .C2(n22085), .A(n22062), .B(n22061), .ZN(
        P1_U3035) );
  AOI22_X1 U23648 ( .A1(n22254), .A2(n22093), .B1(n22092), .B2(n22253), .ZN(
        n22064) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22088), .ZN(n22063) );
  OAI211_X1 U23650 ( .C1(n22091), .C2(n22259), .A(n22064), .B(n22063), .ZN(
        P1_U3043) );
  OAI22_X1 U23651 ( .A1(n22261), .A2(n22091), .B1(n22081), .B2(n22260), .ZN(
        n22065) );
  INV_X1 U23652 ( .A(n22065), .ZN(n22067) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22088), .ZN(n22066) );
  OAI211_X1 U23654 ( .C1(n22267), .C2(n22085), .A(n22067), .B(n22066), .ZN(
        P1_U3051) );
  OAI22_X1 U23655 ( .A1(n22261), .A2(n22097), .B1(n22081), .B2(n22268), .ZN(
        n22068) );
  INV_X1 U23656 ( .A(n22068), .ZN(n22071) );
  AOI22_X1 U23657 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22069), .B2(n22094), .ZN(n22070) );
  OAI211_X1 U23658 ( .C1(n22275), .C2(n22085), .A(n22071), .B(n22070), .ZN(
        P1_U3059) );
  OAI22_X1 U23659 ( .A1(n22277), .A2(n22097), .B1(n22081), .B2(n22276), .ZN(
        n22072) );
  INV_X1 U23660 ( .A(n22072), .ZN(n22074) );
  AOI22_X1 U23661 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22094), .B2(n22279), .ZN(n22073) );
  OAI211_X1 U23662 ( .C1(n22283), .C2(n22085), .A(n22074), .B(n22073), .ZN(
        P1_U3083) );
  AOI22_X1 U23663 ( .A1(n22285), .A2(n22093), .B1(n22092), .B2(n22284), .ZN(
        n22076) );
  AOI22_X1 U23664 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22088), .B2(n22286), .ZN(n22075) );
  OAI211_X1 U23665 ( .C1(n22091), .C2(n22295), .A(n22076), .B(n22075), .ZN(
        P1_U3099) );
  AOI22_X1 U23666 ( .A1(n22291), .A2(n22093), .B1(n22092), .B2(n22290), .ZN(
        n22078) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22094), .ZN(n22077) );
  OAI211_X1 U23668 ( .C1(n22097), .C2(n22295), .A(n22078), .B(n22077), .ZN(
        P1_U3107) );
  AOI22_X1 U23669 ( .A1(n22297), .A2(n22094), .B1(n22092), .B2(n22296), .ZN(
        n22080) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22299), .B1(
        n22298), .B2(n22088), .ZN(n22079) );
  OAI211_X1 U23671 ( .C1(n22302), .C2(n22085), .A(n22080), .B(n22079), .ZN(
        P1_U3115) );
  OAI22_X1 U23672 ( .A1(n22317), .A2(n22091), .B1(n22081), .B2(n22303), .ZN(
        n22082) );
  INV_X1 U23673 ( .A(n22082), .ZN(n22084) );
  AOI22_X1 U23674 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22088), .B2(n22306), .ZN(n22083) );
  OAI211_X1 U23675 ( .C1(n22311), .C2(n22085), .A(n22084), .B(n22083), .ZN(
        P1_U3131) );
  AOI22_X1 U23676 ( .A1(n22092), .A2(n22313), .B1(n22312), .B2(n22093), .ZN(
        n22087) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22094), .ZN(n22086) );
  OAI211_X1 U23678 ( .C1(n22097), .C2(n22317), .A(n22087), .B(n22086), .ZN(
        P1_U3139) );
  AOI22_X1 U23679 ( .A1(n22092), .A2(n22319), .B1(n22093), .B2(n22318), .ZN(
        n22090) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22088), .ZN(n22089) );
  OAI211_X1 U23681 ( .C1(n22091), .C2(n22335), .A(n22090), .B(n22089), .ZN(
        P1_U3147) );
  AOI22_X1 U23682 ( .A1(n22093), .A2(n22328), .B1(n22092), .B2(n22326), .ZN(
        n22096) );
  AOI22_X1 U23683 ( .A1(n22094), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n22095) );
  OAI211_X1 U23684 ( .C1(n22097), .C2(n22335), .A(n22096), .B(n22095), .ZN(
        P1_U3155) );
  OAI22_X1 U23685 ( .A1(n22247), .A2(n22134), .B1(n22118), .B2(n22246), .ZN(
        n22098) );
  INV_X1 U23686 ( .A(n22098), .ZN(n22100) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22131), .ZN(n22099) );
  OAI211_X1 U23688 ( .C1(n22252), .C2(n22122), .A(n22100), .B(n22099), .ZN(
        P1_U3036) );
  AOI22_X1 U23689 ( .A1(n22254), .A2(n22130), .B1(n22129), .B2(n22253), .ZN(
        n22102) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22125), .ZN(n22101) );
  OAI211_X1 U23691 ( .C1(n22128), .C2(n22259), .A(n22102), .B(n22101), .ZN(
        P1_U3044) );
  OAI22_X1 U23692 ( .A1(n22261), .A2(n22128), .B1(n22118), .B2(n22260), .ZN(
        n22103) );
  INV_X1 U23693 ( .A(n22103), .ZN(n22105) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22125), .ZN(n22104) );
  OAI211_X1 U23695 ( .C1(n22267), .C2(n22122), .A(n22105), .B(n22104), .ZN(
        P1_U3052) );
  OAI22_X1 U23696 ( .A1(n22269), .A2(n22128), .B1(n22118), .B2(n22268), .ZN(
        n22106) );
  INV_X1 U23697 ( .A(n22106), .ZN(n22108) );
  AOI22_X1 U23698 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22125), .B2(n22271), .ZN(n22107) );
  OAI211_X1 U23699 ( .C1(n22275), .C2(n22122), .A(n22108), .B(n22107), .ZN(
        P1_U3060) );
  OAI22_X1 U23700 ( .A1(n22277), .A2(n22134), .B1(n22118), .B2(n22276), .ZN(
        n22109) );
  INV_X1 U23701 ( .A(n22109), .ZN(n22111) );
  AOI22_X1 U23702 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22131), .B2(n22279), .ZN(n22110) );
  OAI211_X1 U23703 ( .C1(n22283), .C2(n22122), .A(n22111), .B(n22110), .ZN(
        P1_U3084) );
  AOI22_X1 U23704 ( .A1(n22285), .A2(n22130), .B1(n22129), .B2(n22284), .ZN(
        n22113) );
  AOI22_X1 U23705 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22125), .B2(n22286), .ZN(n22112) );
  OAI211_X1 U23706 ( .C1(n22128), .C2(n22295), .A(n22113), .B(n22112), .ZN(
        P1_U3100) );
  AOI22_X1 U23707 ( .A1(n22291), .A2(n22130), .B1(n22129), .B2(n22290), .ZN(
        n22115) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22131), .ZN(n22114) );
  OAI211_X1 U23709 ( .C1(n22134), .C2(n22295), .A(n22115), .B(n22114), .ZN(
        P1_U3108) );
  AOI22_X1 U23710 ( .A1(n22298), .A2(n22125), .B1(n22129), .B2(n22296), .ZN(
        n22117) );
  AOI22_X1 U23711 ( .A1(n22299), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22131), .B2(n22297), .ZN(n22116) );
  OAI211_X1 U23712 ( .C1(n22302), .C2(n22122), .A(n22117), .B(n22116), .ZN(
        P1_U3116) );
  OAI22_X1 U23713 ( .A1(n22317), .A2(n22128), .B1(n22118), .B2(n22303), .ZN(
        n22119) );
  INV_X1 U23714 ( .A(n22119), .ZN(n22121) );
  AOI22_X1 U23715 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22125), .B2(n22306), .ZN(n22120) );
  OAI211_X1 U23716 ( .C1(n22311), .C2(n22122), .A(n22121), .B(n22120), .ZN(
        P1_U3132) );
  AOI22_X1 U23717 ( .A1(n22129), .A2(n22313), .B1(n22312), .B2(n22130), .ZN(
        n22124) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22131), .ZN(n22123) );
  OAI211_X1 U23719 ( .C1(n22134), .C2(n22317), .A(n22124), .B(n22123), .ZN(
        P1_U3140) );
  AOI22_X1 U23720 ( .A1(n22129), .A2(n22319), .B1(n22130), .B2(n22318), .ZN(
        n22127) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22125), .ZN(n22126) );
  OAI211_X1 U23722 ( .C1(n22128), .C2(n22335), .A(n22127), .B(n22126), .ZN(
        P1_U3148) );
  AOI22_X1 U23723 ( .A1(n22130), .A2(n22328), .B1(n22129), .B2(n22326), .ZN(
        n22133) );
  AOI22_X1 U23724 ( .A1(n22131), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n22132) );
  OAI211_X1 U23725 ( .C1(n22134), .C2(n22335), .A(n22133), .B(n22132), .ZN(
        P1_U3156) );
  OAI22_X1 U23726 ( .A1(n22247), .A2(n22171), .B1(n22155), .B2(n22246), .ZN(
        n22135) );
  INV_X1 U23727 ( .A(n22135), .ZN(n22137) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22168), .ZN(n22136) );
  OAI211_X1 U23729 ( .C1(n22252), .C2(n22159), .A(n22137), .B(n22136), .ZN(
        P1_U3037) );
  AOI22_X1 U23730 ( .A1(n22254), .A2(n22167), .B1(n22166), .B2(n22253), .ZN(
        n22139) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22162), .ZN(n22138) );
  OAI211_X1 U23732 ( .C1(n22165), .C2(n22259), .A(n22139), .B(n22138), .ZN(
        P1_U3045) );
  OAI22_X1 U23733 ( .A1(n22259), .A2(n22171), .B1(n22155), .B2(n22260), .ZN(
        n22140) );
  INV_X1 U23734 ( .A(n22140), .ZN(n22142) );
  AOI22_X1 U23735 ( .A1(n22264), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22168), .B2(n22271), .ZN(n22141) );
  OAI211_X1 U23736 ( .C1(n22267), .C2(n22159), .A(n22142), .B(n22141), .ZN(
        P1_U3053) );
  OAI22_X1 U23737 ( .A1(n22269), .A2(n22165), .B1(n22155), .B2(n22268), .ZN(
        n22143) );
  INV_X1 U23738 ( .A(n22143), .ZN(n22145) );
  AOI22_X1 U23739 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22162), .B2(n22271), .ZN(n22144) );
  OAI211_X1 U23740 ( .C1(n22275), .C2(n22159), .A(n22145), .B(n22144), .ZN(
        P1_U3061) );
  OAI22_X1 U23741 ( .A1(n22277), .A2(n22171), .B1(n22155), .B2(n22276), .ZN(
        n22146) );
  INV_X1 U23742 ( .A(n22146), .ZN(n22148) );
  AOI22_X1 U23743 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22168), .B2(n22279), .ZN(n22147) );
  OAI211_X1 U23744 ( .C1(n22283), .C2(n22159), .A(n22148), .B(n22147), .ZN(
        P1_U3085) );
  AOI22_X1 U23745 ( .A1(n22285), .A2(n22167), .B1(n22166), .B2(n22284), .ZN(
        n22150) );
  AOI22_X1 U23746 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22162), .B2(n22286), .ZN(n22149) );
  OAI211_X1 U23747 ( .C1(n22165), .C2(n22295), .A(n22150), .B(n22149), .ZN(
        P1_U3101) );
  AOI22_X1 U23748 ( .A1(n22291), .A2(n22167), .B1(n22166), .B2(n22290), .ZN(
        n22152) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22168), .ZN(n22151) );
  OAI211_X1 U23750 ( .C1(n22171), .C2(n22295), .A(n22152), .B(n22151), .ZN(
        P1_U3109) );
  AOI22_X1 U23751 ( .A1(n22297), .A2(n22168), .B1(n22166), .B2(n22296), .ZN(
        n22154) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22299), .B1(
        n22298), .B2(n22162), .ZN(n22153) );
  OAI211_X1 U23753 ( .C1(n22302), .C2(n22159), .A(n22154), .B(n22153), .ZN(
        P1_U3117) );
  OAI22_X1 U23754 ( .A1(n22317), .A2(n22165), .B1(n22155), .B2(n22303), .ZN(
        n22156) );
  INV_X1 U23755 ( .A(n22156), .ZN(n22158) );
  AOI22_X1 U23756 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22162), .B2(n22306), .ZN(n22157) );
  OAI211_X1 U23757 ( .C1(n22311), .C2(n22159), .A(n22158), .B(n22157), .ZN(
        P1_U3133) );
  AOI22_X1 U23758 ( .A1(n22166), .A2(n22313), .B1(n22312), .B2(n22167), .ZN(
        n22161) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22168), .ZN(n22160) );
  OAI211_X1 U23760 ( .C1(n22171), .C2(n22317), .A(n22161), .B(n22160), .ZN(
        P1_U3141) );
  AOI22_X1 U23761 ( .A1(n22166), .A2(n22319), .B1(n22167), .B2(n22318), .ZN(
        n22164) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22162), .ZN(n22163) );
  OAI211_X1 U23763 ( .C1(n22165), .C2(n22335), .A(n22164), .B(n22163), .ZN(
        P1_U3149) );
  AOI22_X1 U23764 ( .A1(n22167), .A2(n22328), .B1(n22166), .B2(n22326), .ZN(
        n22170) );
  AOI22_X1 U23765 ( .A1(n22168), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n22169) );
  OAI211_X1 U23766 ( .C1(n22171), .C2(n22335), .A(n22170), .B(n22169), .ZN(
        P1_U3157) );
  OAI22_X1 U23767 ( .A1(n22247), .A2(n22208), .B1(n22192), .B2(n22246), .ZN(
        n22172) );
  INV_X1 U23768 ( .A(n22172), .ZN(n22174) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22205), .ZN(n22173) );
  OAI211_X1 U23770 ( .C1(n22252), .C2(n22196), .A(n22174), .B(n22173), .ZN(
        P1_U3038) );
  AOI22_X1 U23771 ( .A1(n22254), .A2(n22204), .B1(n22203), .B2(n22253), .ZN(
        n22176) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22199), .ZN(n22175) );
  OAI211_X1 U23773 ( .C1(n22202), .C2(n22259), .A(n22176), .B(n22175), .ZN(
        P1_U3046) );
  OAI22_X1 U23774 ( .A1(n22261), .A2(n22202), .B1(n22192), .B2(n22260), .ZN(
        n22177) );
  INV_X1 U23775 ( .A(n22177), .ZN(n22179) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22199), .ZN(n22178) );
  OAI211_X1 U23777 ( .C1(n22267), .C2(n22196), .A(n22179), .B(n22178), .ZN(
        P1_U3054) );
  OAI22_X1 U23778 ( .A1(n22269), .A2(n22202), .B1(n22192), .B2(n22268), .ZN(
        n22180) );
  INV_X1 U23779 ( .A(n22180), .ZN(n22182) );
  AOI22_X1 U23780 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22199), .B2(n22271), .ZN(n22181) );
  OAI211_X1 U23781 ( .C1(n22275), .C2(n22196), .A(n22182), .B(n22181), .ZN(
        P1_U3062) );
  OAI22_X1 U23782 ( .A1(n22277), .A2(n22208), .B1(n22192), .B2(n22276), .ZN(
        n22183) );
  INV_X1 U23783 ( .A(n22183), .ZN(n22185) );
  AOI22_X1 U23784 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22205), .B2(n22279), .ZN(n22184) );
  OAI211_X1 U23785 ( .C1(n22283), .C2(n22196), .A(n22185), .B(n22184), .ZN(
        P1_U3086) );
  AOI22_X1 U23786 ( .A1(n22285), .A2(n22204), .B1(n22203), .B2(n22284), .ZN(
        n22187) );
  AOI22_X1 U23787 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22199), .B2(n22286), .ZN(n22186) );
  OAI211_X1 U23788 ( .C1(n22202), .C2(n22295), .A(n22187), .B(n22186), .ZN(
        P1_U3102) );
  AOI22_X1 U23789 ( .A1(n22291), .A2(n22204), .B1(n22203), .B2(n22290), .ZN(
        n22189) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22205), .ZN(n22188) );
  OAI211_X1 U23791 ( .C1(n22208), .C2(n22295), .A(n22189), .B(n22188), .ZN(
        P1_U3110) );
  AOI22_X1 U23792 ( .A1(n22298), .A2(n22199), .B1(n22203), .B2(n22296), .ZN(
        n22191) );
  AOI22_X1 U23793 ( .A1(n22299), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22205), .B2(n22297), .ZN(n22190) );
  OAI211_X1 U23794 ( .C1(n22302), .C2(n22196), .A(n22191), .B(n22190), .ZN(
        P1_U3118) );
  OAI22_X1 U23795 ( .A1(n22317), .A2(n22202), .B1(n22192), .B2(n22303), .ZN(
        n22193) );
  INV_X1 U23796 ( .A(n22193), .ZN(n22195) );
  AOI22_X1 U23797 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22199), .B2(n22306), .ZN(n22194) );
  OAI211_X1 U23798 ( .C1(n22311), .C2(n22196), .A(n22195), .B(n22194), .ZN(
        P1_U3134) );
  AOI22_X1 U23799 ( .A1(n22203), .A2(n22313), .B1(n22312), .B2(n22204), .ZN(
        n22198) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22205), .ZN(n22197) );
  OAI211_X1 U23801 ( .C1(n22208), .C2(n22317), .A(n22198), .B(n22197), .ZN(
        P1_U3142) );
  AOI22_X1 U23802 ( .A1(n22203), .A2(n22319), .B1(n22204), .B2(n22318), .ZN(
        n22201) );
  AOI22_X1 U23803 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22199), .ZN(n22200) );
  OAI211_X1 U23804 ( .C1(n22202), .C2(n22335), .A(n22201), .B(n22200), .ZN(
        P1_U3150) );
  AOI22_X1 U23805 ( .A1(n22204), .A2(n22328), .B1(n22203), .B2(n22326), .ZN(
        n22207) );
  AOI22_X1 U23806 ( .A1(n22205), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n22206) );
  OAI211_X1 U23807 ( .C1(n22208), .C2(n22335), .A(n22207), .B(n22206), .ZN(
        P1_U3158) );
  OAI22_X1 U23808 ( .A1(n22247), .A2(n22245), .B1(n22229), .B2(n22246), .ZN(
        n22209) );
  INV_X1 U23809 ( .A(n22209), .ZN(n22211) );
  AOI22_X1 U23810 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22242), .ZN(n22210) );
  OAI211_X1 U23811 ( .C1(n22252), .C2(n22233), .A(n22211), .B(n22210), .ZN(
        P1_U3039) );
  AOI22_X1 U23812 ( .A1(n22254), .A2(n22241), .B1(n22240), .B2(n22253), .ZN(
        n22213) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22236), .ZN(n22212) );
  OAI211_X1 U23814 ( .C1(n22239), .C2(n22259), .A(n22213), .B(n22212), .ZN(
        P1_U3047) );
  OAI22_X1 U23815 ( .A1(n22261), .A2(n22239), .B1(n22229), .B2(n22260), .ZN(
        n22214) );
  INV_X1 U23816 ( .A(n22214), .ZN(n22216) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22236), .ZN(n22215) );
  OAI211_X1 U23818 ( .C1(n22267), .C2(n22233), .A(n22216), .B(n22215), .ZN(
        P1_U3055) );
  OAI22_X1 U23819 ( .A1(n22269), .A2(n22239), .B1(n22229), .B2(n22268), .ZN(
        n22217) );
  INV_X1 U23820 ( .A(n22217), .ZN(n22219) );
  AOI22_X1 U23821 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22236), .B2(n22271), .ZN(n22218) );
  OAI211_X1 U23822 ( .C1(n22275), .C2(n22233), .A(n22219), .B(n22218), .ZN(
        P1_U3063) );
  OAI22_X1 U23823 ( .A1(n22277), .A2(n22245), .B1(n22229), .B2(n22276), .ZN(
        n22220) );
  INV_X1 U23824 ( .A(n22220), .ZN(n22222) );
  AOI22_X1 U23825 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22242), .B2(n22279), .ZN(n22221) );
  OAI211_X1 U23826 ( .C1(n22283), .C2(n22233), .A(n22222), .B(n22221), .ZN(
        P1_U3087) );
  AOI22_X1 U23827 ( .A1(n22285), .A2(n22241), .B1(n22240), .B2(n22284), .ZN(
        n22224) );
  AOI22_X1 U23828 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22236), .B2(n22286), .ZN(n22223) );
  OAI211_X1 U23829 ( .C1(n22239), .C2(n22295), .A(n22224), .B(n22223), .ZN(
        P1_U3103) );
  AOI22_X1 U23830 ( .A1(n22291), .A2(n22241), .B1(n22240), .B2(n22290), .ZN(
        n22226) );
  AOI22_X1 U23831 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22242), .ZN(n22225) );
  OAI211_X1 U23832 ( .C1(n22245), .C2(n22295), .A(n22226), .B(n22225), .ZN(
        P1_U3111) );
  AOI22_X1 U23833 ( .A1(n22297), .A2(n22242), .B1(n22240), .B2(n22296), .ZN(
        n22228) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22299), .B1(
        n22298), .B2(n22236), .ZN(n22227) );
  OAI211_X1 U23835 ( .C1(n22302), .C2(n22233), .A(n22228), .B(n22227), .ZN(
        P1_U3119) );
  OAI22_X1 U23836 ( .A1(n22317), .A2(n22239), .B1(n22229), .B2(n22303), .ZN(
        n22230) );
  INV_X1 U23837 ( .A(n22230), .ZN(n22232) );
  AOI22_X1 U23838 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22236), .B2(n22306), .ZN(n22231) );
  OAI211_X1 U23839 ( .C1(n22311), .C2(n22233), .A(n22232), .B(n22231), .ZN(
        P1_U3135) );
  AOI22_X1 U23840 ( .A1(n22240), .A2(n22313), .B1(n22312), .B2(n22241), .ZN(
        n22235) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22242), .ZN(n22234) );
  OAI211_X1 U23842 ( .C1(n22245), .C2(n22317), .A(n22235), .B(n22234), .ZN(
        P1_U3143) );
  AOI22_X1 U23843 ( .A1(n22240), .A2(n22319), .B1(n22241), .B2(n22318), .ZN(
        n22238) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22236), .ZN(n22237) );
  OAI211_X1 U23845 ( .C1(n22239), .C2(n22335), .A(n22238), .B(n22237), .ZN(
        P1_U3151) );
  AOI22_X1 U23846 ( .A1(n22241), .A2(n22328), .B1(n22240), .B2(n22326), .ZN(
        n22244) );
  AOI22_X1 U23847 ( .A1(n22242), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n22243) );
  OAI211_X1 U23848 ( .C1(n22245), .C2(n22335), .A(n22244), .B(n22243), .ZN(
        P1_U3159) );
  OAI22_X1 U23849 ( .A1(n22247), .A2(n22336), .B1(n22304), .B2(n22246), .ZN(
        n22248) );
  INV_X1 U23850 ( .A(n22248), .ZN(n22251) );
  AOI22_X1 U23851 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22249), .B1(
        n22255), .B2(n22332), .ZN(n22250) );
  OAI211_X1 U23852 ( .C1(n22252), .C2(n22310), .A(n22251), .B(n22250), .ZN(
        P1_U3040) );
  AOI22_X1 U23853 ( .A1(n22254), .A2(n22329), .B1(n22327), .B2(n22253), .ZN(
        n22258) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22256), .B1(
        n22255), .B2(n22320), .ZN(n22257) );
  OAI211_X1 U23855 ( .C1(n22325), .C2(n22259), .A(n22258), .B(n22257), .ZN(
        P1_U3048) );
  OAI22_X1 U23856 ( .A1(n22261), .A2(n22325), .B1(n22304), .B2(n22260), .ZN(
        n22262) );
  INV_X1 U23857 ( .A(n22262), .ZN(n22266) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22264), .B1(
        n22263), .B2(n22320), .ZN(n22265) );
  OAI211_X1 U23859 ( .C1(n22267), .C2(n22310), .A(n22266), .B(n22265), .ZN(
        P1_U3056) );
  OAI22_X1 U23860 ( .A1(n22269), .A2(n22325), .B1(n22304), .B2(n22268), .ZN(
        n22270) );
  INV_X1 U23861 ( .A(n22270), .ZN(n22274) );
  AOI22_X1 U23862 ( .A1(n22272), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22320), .B2(n22271), .ZN(n22273) );
  OAI211_X1 U23863 ( .C1(n22275), .C2(n22310), .A(n22274), .B(n22273), .ZN(
        P1_U3064) );
  OAI22_X1 U23864 ( .A1(n22277), .A2(n22336), .B1(n22304), .B2(n22276), .ZN(
        n22278) );
  INV_X1 U23865 ( .A(n22278), .ZN(n22282) );
  AOI22_X1 U23866 ( .A1(n22280), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22332), .B2(n22279), .ZN(n22281) );
  OAI211_X1 U23867 ( .C1(n22283), .C2(n22310), .A(n22282), .B(n22281), .ZN(
        P1_U3088) );
  AOI22_X1 U23868 ( .A1(n22285), .A2(n22329), .B1(n22327), .B2(n22284), .ZN(
        n22289) );
  AOI22_X1 U23869 ( .A1(n22287), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n22320), .B2(n22286), .ZN(n22288) );
  OAI211_X1 U23870 ( .C1(n22325), .C2(n22295), .A(n22289), .B(n22288), .ZN(
        P1_U3104) );
  AOI22_X1 U23871 ( .A1(n22291), .A2(n22329), .B1(n22327), .B2(n22290), .ZN(
        n22294) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22292), .B1(
        n22298), .B2(n22332), .ZN(n22293) );
  OAI211_X1 U23873 ( .C1(n22336), .C2(n22295), .A(n22294), .B(n22293), .ZN(
        P1_U3112) );
  AOI22_X1 U23874 ( .A1(n22297), .A2(n22332), .B1(n22327), .B2(n22296), .ZN(
        n22301) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22299), .B1(
        n22298), .B2(n22320), .ZN(n22300) );
  OAI211_X1 U23876 ( .C1(n22302), .C2(n22310), .A(n22301), .B(n22300), .ZN(
        P1_U3120) );
  OAI22_X1 U23877 ( .A1(n22317), .A2(n22325), .B1(n22304), .B2(n22303), .ZN(
        n22305) );
  INV_X1 U23878 ( .A(n22305), .ZN(n22309) );
  AOI22_X1 U23879 ( .A1(n22307), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n22320), .B2(n22306), .ZN(n22308) );
  OAI211_X1 U23880 ( .C1(n22311), .C2(n22310), .A(n22309), .B(n22308), .ZN(
        P1_U3136) );
  AOI22_X1 U23881 ( .A1(n22327), .A2(n22313), .B1(n22312), .B2(n22329), .ZN(
        n22316) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22314), .B1(
        n22321), .B2(n22332), .ZN(n22315) );
  OAI211_X1 U23883 ( .C1(n22336), .C2(n22317), .A(n22316), .B(n22315), .ZN(
        P1_U3144) );
  AOI22_X1 U23884 ( .A1(n22327), .A2(n22319), .B1(n22329), .B2(n22318), .ZN(
        n22324) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22322), .B1(
        n22321), .B2(n22320), .ZN(n22323) );
  OAI211_X1 U23886 ( .C1(n22325), .C2(n22335), .A(n22324), .B(n22323), .ZN(
        P1_U3152) );
  AOI22_X1 U23887 ( .A1(n22329), .A2(n22328), .B1(n22327), .B2(n22326), .ZN(
        n22334) );
  AOI22_X1 U23888 ( .A1(n22332), .A2(n22331), .B1(n22330), .B2(
        P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n22333) );
  OAI211_X1 U23889 ( .C1(n22336), .C2(n22335), .A(n22334), .B(n22333), .ZN(
        P1_U3160) );
  AOI22_X1 U23890 ( .A1(n22339), .A2(n14113), .B1(n22338), .B2(n22337), .ZN(
        P1_U3486) );
  NAND2_X1 U15474 ( .A1(n13918), .A2(n13672), .ZN(n14919) );
  NAND2_X1 U11194 ( .A1(n13691), .A2(n13919), .ZN(n13722) );
  XNOR2_X1 U12674 ( .A(n13921), .B(n13920), .ZN(n13923) );
  XNOR2_X1 U11193 ( .A(n13722), .B(n13723), .ZN(n13926) );
  NOR2_X2 U11145 ( .A1(n22337), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19855) );
  CLKBUF_X1 U11183 ( .A(n11547), .Z(n11635) );
  CLKBUF_X1 U11184 ( .A(n13918), .Z(n13921) );
  AND2_X1 U11226 ( .A1(n13621), .A2(n15096), .ZN(n13616) );
  CLKBUF_X1 U11488 ( .A(n13482), .Z(n11020) );
  AND2_X1 U11714 ( .A1(n11201), .A2(n15128), .ZN(n19334) );
  CLKBUF_X1 U11892 ( .A(n19327), .Z(n19625) );
  CLKBUF_X1 U12376 ( .A(n15540), .Z(n15541) );
  CLKBUF_X1 U12562 ( .A(n16280), .Z(n16329) );
  CLKBUF_X1 U12627 ( .A(n20393), .Z(n11019) );
  CLKBUF_X1 U12675 ( .A(n19010), .Z(n18964) );
endmodule

