

module b21_C_SARLock_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167;

  NAND2_X1 U4900 ( .A1(n7232), .A2(n7233), .ZN(n7316) );
  BUF_X1 U4901 ( .A(n5668), .Z(n5790) );
  CLKBUF_X1 U4902 ( .A(n6818), .Z(n9703) );
  BUF_X2 U4903 ( .A(n5177), .Z(n5516) );
  INV_X1 U4904 ( .A(n6081), .ZN(n6548) );
  CLKBUF_X2 U4905 ( .A(n6310), .Z(n7905) );
  CLKBUF_X2 U4906 ( .A(n6095), .Z(n7477) );
  CLKBUF_X1 U4907 ( .A(n6203), .Z(n6583) );
  AND2_X1 U4908 ( .A1(n7896), .A2(n8730), .ZN(n6111) );
  NAND2_X1 U4909 ( .A1(n7896), .A2(n6069), .ZN(n6095) );
  XNOR2_X1 U4910 ( .A(n5909), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6070) );
  NOR3_X1 U4911 ( .A1(n9513), .A2(n5543), .A3(n5611), .ZN(n4394) );
  NAND2_X1 U4912 ( .A1(n5599), .A2(n5598), .ZN(n5611) );
  CLKBUF_X3 U4913 ( .A(P1_U4006), .Z(n10144) );
  INV_X2 U4914 ( .A(n8145), .ZN(n8179) );
  INV_X1 U4915 ( .A(n7905), .ZN(n7370) );
  AND2_X2 U4916 ( .A1(n6070), .A2(n6069), .ZN(n6145) );
  NAND2_X1 U4917 ( .A1(n7918), .A2(n9606), .ZN(n9629) );
  OR2_X1 U4918 ( .A1(n8732), .A2(n8735), .ZN(n4546) );
  AOI21_X1 U4919 ( .B1(n5619), .B2(n8758), .A(n5618), .ZN(n6159) );
  INV_X1 U4920 ( .A(n8753), .ZN(n5761) );
  INV_X1 U4921 ( .A(n6145), .ZN(n7480) );
  INV_X1 U4922 ( .A(n6583), .ZN(n7907) );
  AND4_X1 U4923 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n7853)
         );
  OAI211_X1 U4924 ( .C1(n5168), .C2(n9407), .A(n5175), .B(n5174), .ZN(n7869)
         );
  OR2_X1 U4925 ( .A1(n5131), .A2(n9218), .ZN(n5111) );
  INV_X1 U4926 ( .A(n6905), .ZN(n8885) );
  INV_X2 U4927 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI211_X1 U4928 ( .C1(n6423), .C2(n6422), .A(n6421), .B(n6420), .ZN(n9583)
         );
  AOI21_X2 U4929 ( .B1(n9042), .B2(n5586), .A(n5585), .ZN(n9022) );
  AOI21_X2 U4930 ( .B1(n9055), .B2(n9054), .A(n5584), .ZN(n9042) );
  OAI21_X2 U4931 ( .B1(n9099), .B2(n7641), .A(n7677), .ZN(n9085) );
  BUF_X2 U4932 ( .A(n9614), .Z(n4395) );
  AND2_X4 U4933 ( .A1(n5138), .A2(n7512), .ZN(n5193) );
  AND3_X2 U4934 ( .A1(n6082), .A2(n6081), .A3(n6138), .ZN(n8046) );
  NAND2_X1 U4935 ( .A1(n6082), .A2(n6548), .ZN(n6752) );
  XNOR2_X2 U4936 ( .A(n5938), .B(n5937), .ZN(n6082) );
  NAND2_X2 U4937 ( .A1(n5524), .A2(n9368), .ZN(n5168) );
  XNOR2_X2 U4938 ( .A(n5111), .B(n5130), .ZN(n5524) );
  OAI21_X2 U4939 ( .B1(n6883), .B2(n4918), .A(n4916), .ZN(n7075) );
  OAI22_X2 U4940 ( .A1(n6990), .A2(n6991), .B1(n9763), .B2(n6888), .ZN(n6883)
         );
  NAND2_X1 U4941 ( .A1(n8443), .A2(n8024), .ZN(n8425) );
  AOI21_X1 U4942 ( .B1(n4900), .B2(n4902), .A(n4446), .ZN(n4898) );
  NAND2_X1 U4943 ( .A1(n4925), .A2(n4926), .ZN(n8550) );
  NAND2_X1 U4944 ( .A1(n5590), .A2(n4975), .ZN(n8993) );
  NAND2_X1 U4945 ( .A1(n5747), .A2(n5746), .ZN(n8834) );
  NAND2_X1 U4946 ( .A1(n8799), .A2(n8800), .ZN(n8798) );
  NAND2_X1 U4947 ( .A1(n4792), .A2(n4790), .ZN(n8998) );
  NAND3_X1 U4948 ( .A1(n4877), .A2(n4876), .A3(n8597), .ZN(n8596) );
  AOI21_X1 U4949 ( .B1(n4881), .B2(n6885), .A(n4532), .ZN(n7081) );
  NAND2_X1 U4950 ( .A1(n5191), .A2(n7757), .ZN(n6726) );
  NAND4_X1 U4951 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n8277)
         );
  NAND2_X1 U4952 ( .A1(n8281), .A2(n6776), .ZN(n6814) );
  XNOR2_X1 U4953 ( .A(n4774), .B(n4773), .ZN(n6429) );
  XNOR2_X1 U4954 ( .A(n6754), .B(n4631), .ZN(n6815) );
  NAND4_X1 U4955 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n8281)
         );
  AND4_X1 U4956 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n6824)
         );
  AND3_X1 U4957 ( .A1(n6315), .A2(n6314), .A3(n6313), .ZN(n9717) );
  AND4_X1 U4958 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n6556)
         );
  BUF_X2 U4959 ( .A(n5615), .Z(n8756) );
  NAND4_X1 U4960 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n9253)
         );
  AND4_X1 U4961 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5178), .ZN(n7867)
         );
  AND4_X1 U4962 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n6905)
         );
  NOR2_X1 U4963 ( .A1(n5974), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X2 U4964 ( .A(n5520), .ZN(n5496) );
  OR2_X1 U4965 ( .A1(n6095), .A2(n6071), .ZN(n6072) );
  NAND4_X1 U4966 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n5631)
         );
  AND2_X2 U4967 ( .A1(n8759), .A2(n5612), .ZN(n8753) );
  AND2_X2 U4968 ( .A1(n5610), .A2(n5611), .ZN(n8759) );
  AND2_X1 U4969 ( .A1(n8106), .A2(n5139), .ZN(n5268) );
  AND2_X1 U4970 ( .A1(n6070), .A2(n8730), .ZN(n6096) );
  NAND2_X2 U4971 ( .A1(n6142), .A2(n8095), .ZN(n6423) );
  NAND2_X1 U4972 ( .A1(n9219), .A2(n5137), .ZN(n7512) );
  OAI21_X1 U4973 ( .B1(n5939), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U4974 ( .A1(n4970), .A2(n5935), .ZN(n8095) );
  NAND2_X1 U4975 ( .A1(n8723), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U4976 ( .A(n5911), .B(n5907), .ZN(n8730) );
  NAND2_X1 U4977 ( .A1(n5910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  NAND3_X1 U4978 ( .A1(n4924), .A2(n5906), .A3(n4657), .ZN(n5910) );
  INV_X1 U4979 ( .A(n5904), .ZN(n4924) );
  INV_X2 U4980 ( .A(n7259), .ZN(n4396) );
  INV_X2 U4981 ( .A(n5893), .ZN(n5834) );
  NAND2_X2 U4982 ( .A1(n4803), .A2(n4802), .ZN(n7555) );
  AND2_X1 U4983 ( .A1(n4422), .A2(n5835), .ZN(n4922) );
  AND2_X1 U4984 ( .A1(n5831), .A2(n5830), .ZN(n5881) );
  AND2_X1 U4985 ( .A1(n4772), .A2(n5240), .ZN(n4771) );
  AND2_X1 U4986 ( .A1(n5102), .A2(n5101), .ZN(n4969) );
  NOR2_X1 U4987 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5102) );
  INV_X1 U4988 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5504) );
  INV_X1 U4989 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5860) );
  INV_X1 U4990 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5937) );
  INV_X1 U4991 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6079) );
  INV_X1 U4992 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4614) );
  INV_X1 U4993 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5845) );
  INV_X1 U4994 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5348) );
  NOR2_X1 U4995 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5830) );
  INV_X1 U4996 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5833) );
  NOR2_X1 U4997 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5831) );
  INV_X4 U4998 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X2 U4999 ( .A1(n5168), .A2(n7555), .ZN(n5185) );
  AOI21_X1 U5000 ( .B1(n9680), .B2(n9688), .A(n9689), .ZN(n8622) );
  INV_X1 U5001 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5927) );
  INV_X1 U5002 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5853) );
  OR2_X1 U5003 ( .A1(n5611), .A2(n5609), .ZN(n5668) );
  NAND2_X1 U5004 ( .A1(n4743), .A2(n8854), .ZN(n4742) );
  NAND2_X1 U5005 ( .A1(n5065), .A2(n5064), .ZN(n5425) );
  NAND2_X1 U5006 ( .A1(n5414), .A2(n5413), .ZN(n5065) );
  NAND2_X1 U5007 ( .A1(n5361), .A2(n4966), .ZN(n4965) );
  INV_X1 U5008 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4966) );
  AOI21_X1 U5009 ( .B1(n4515), .B2(n4518), .A(n5016), .ZN(n4513) );
  OR2_X1 U5010 ( .A1(n4536), .A2(n5730), .ZN(n4535) );
  INV_X1 U5011 ( .A(n8004), .ZN(n4643) );
  OR2_X1 U5012 ( .A1(n6754), .A2(n4631), .ZN(n6839) );
  INV_X1 U5013 ( .A(SI_16_), .ZN(n9901) );
  INV_X1 U5014 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5043) );
  OR2_X1 U5015 ( .A1(n4674), .A2(n4671), .ZN(n4670) );
  INV_X1 U5016 ( .A(n8191), .ZN(n4671) );
  NAND2_X1 U5017 ( .A1(n4658), .A2(n6087), .ZN(n6191) );
  AND2_X1 U5018 ( .A1(n6133), .A2(n6749), .ZN(n4658) );
  INV_X1 U5019 ( .A(n6102), .ZN(n8145) );
  OR2_X1 U5020 ( .A1(n8653), .A2(n8161), .ZN(n8017) );
  NOR2_X1 U5021 ( .A1(n8663), .A2(n4626), .ZN(n4625) );
  INV_X1 U5022 ( .A(n4627), .ZN(n4626) );
  OR2_X1 U5023 ( .A1(n8663), .A2(n8195), .ZN(n8007) );
  INV_X1 U5024 ( .A(n4933), .ZN(n4930) );
  INV_X1 U5025 ( .A(n7367), .ZN(n4932) );
  OAI21_X1 U5026 ( .B1(n7118), .B2(n4445), .A(n4955), .ZN(n4536) );
  NAND2_X1 U5027 ( .A1(n4957), .A2(n4956), .ZN(n4955) );
  INV_X1 U5028 ( .A(n7131), .ZN(n4957) );
  NAND2_X1 U5029 ( .A1(n4552), .A2(n4551), .ZN(n5682) );
  OR2_X1 U5030 ( .A1(n6943), .A2(n5687), .ZN(n4551) );
  OR2_X1 U5031 ( .A1(n7006), .A2(n5686), .ZN(n4552) );
  AOI21_X1 U5032 ( .B1(n4398), .B2(n4939), .A(n4440), .ZN(n4934) );
  NAND2_X1 U5033 ( .A1(n8745), .A2(n4398), .ZN(n4537) );
  AND2_X1 U5034 ( .A1(n4825), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5035 ( .A1(n4818), .A2(n4820), .ZN(n4817) );
  NOR2_X1 U5036 ( .A1(n8926), .A2(n4826), .ZN(n4825) );
  INV_X1 U5037 ( .A(n4823), .ZN(n4818) );
  NOR2_X1 U5038 ( .A1(n7693), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U5039 ( .A1(n4811), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5040 ( .A1(n6451), .A2(n6450), .ZN(n6449) );
  NAND2_X1 U5041 ( .A1(n4854), .A2(n4855), .ZN(n5414) );
  AOI21_X1 U5042 ( .B1(n4863), .B2(n4857), .A(n4856), .ZN(n4855) );
  INV_X1 U5043 ( .A(n5059), .ZN(n4856) );
  INV_X1 U5044 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U5045 ( .A1(n4483), .A2(n5151), .ZN(n4985) );
  NAND2_X1 U5046 ( .A1(n7555), .A2(n4435), .ZN(n4483) );
  NAND2_X1 U5047 ( .A1(n4630), .A2(n6191), .ZN(n6093) );
  INV_X1 U5048 ( .A(n6754), .ZN(n4630) );
  AND2_X1 U5049 ( .A1(n9581), .A2(n4425), .ZN(n4666) );
  NAND2_X1 U5050 ( .A1(n6417), .A2(n6416), .ZN(n4667) );
  OR2_X1 U5051 ( .A1(n8700), .A2(n6741), .ZN(n6139) );
  NAND2_X1 U5052 ( .A1(n4524), .A2(n4523), .ZN(n7897) );
  INV_X1 U5053 ( .A(n8040), .ZN(n4523) );
  INV_X1 U5054 ( .A(n7507), .ZN(n4524) );
  OR2_X1 U5055 ( .A1(n8638), .A2(n8419), .ZN(n7452) );
  XNOR2_X1 U5056 ( .A(n8638), .B(n7912), .ZN(n8430) );
  NAND2_X1 U5057 ( .A1(n8431), .A2(n8430), .ZN(n8429) );
  AOI21_X1 U5058 ( .B1(n4913), .B2(n4642), .A(n4444), .ZN(n4911) );
  AND2_X1 U5059 ( .A1(n8695), .A2(n8265), .ZN(n7367) );
  AND2_X1 U5060 ( .A1(n8063), .A2(n7937), .ZN(n4884) );
  NAND2_X1 U5061 ( .A1(n6744), .A2(n6743), .ZN(n6753) );
  AND2_X1 U5062 ( .A1(n8700), .A2(n6742), .ZN(n6743) );
  AND2_X1 U5063 ( .A1(n6121), .A2(n6118), .ZN(n9680) );
  OR2_X1 U5064 ( .A1(n7174), .A2(n6117), .ZN(n6118) );
  NAND2_X1 U5065 ( .A1(n5930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  INV_X1 U5066 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5067 ( .A1(n4536), .A2(n5730), .ZN(n7281) );
  NAND2_X1 U5068 ( .A1(n4481), .A2(n4943), .ZN(n8799) );
  AOI21_X1 U5069 ( .B1(n4945), .B2(n4947), .A(n4436), .ZN(n4943) );
  NAND2_X1 U5070 ( .A1(n5733), .A2(n4945), .ZN(n4481) );
  AOI21_X1 U5071 ( .B1(n7561), .B2(n9342), .A(n7786), .ZN(n7821) );
  NAND2_X1 U5072 ( .A1(n4962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5509) );
  INV_X1 U5073 ( .A(n5268), .ZN(n5520) );
  CLKBUF_X2 U5074 ( .A(n5176), .Z(n5472) );
  INV_X1 U5075 ( .A(n5499), .ZN(n5176) );
  AND2_X1 U5076 ( .A1(n5138), .A2(n5139), .ZN(n5177) );
  AND2_X1 U5077 ( .A1(n4952), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5078 ( .A1(n7516), .A2(n7515), .ZN(n8919) );
  INV_X1 U5079 ( .A(n7816), .ZN(n5595) );
  AND2_X1 U5080 ( .A1(n7781), .A2(n7731), .ZN(n8932) );
  OR2_X1 U5081 ( .A1(n9169), .A2(n9046), .ZN(n9035) );
  INV_X1 U5082 ( .A(n4752), .ZN(n4751) );
  OAI21_X1 U5083 ( .B1(n7207), .B2(n4397), .A(n4420), .ZN(n4752) );
  INV_X1 U5084 ( .A(n5229), .ZN(n7560) );
  NAND2_X1 U5085 ( .A1(n5168), .A2(n4895), .ZN(n5229) );
  OR2_X1 U5086 ( .A1(n7746), .A2(n7831), .ZN(n9534) );
  AND2_X1 U5087 ( .A1(n5545), .A2(n5544), .ZN(n5536) );
  XNOR2_X1 U5088 ( .A(n7558), .B(n7557), .ZN(n8721) );
  NAND2_X1 U5089 ( .A1(n4833), .A2(n4834), .ZN(n5262) );
  AOI21_X1 U5090 ( .B1(n4835), .B2(n4406), .A(n4448), .ZN(n4834) );
  OAI211_X1 U5091 ( .C1(n4700), .C2(n4695), .A(n4694), .B(n4468), .ZN(n4693)
         );
  INV_X1 U5092 ( .A(n4698), .ZN(n4695) );
  NAND2_X1 U5093 ( .A1(n4700), .A2(n4433), .ZN(n4694) );
  AOI21_X1 U5094 ( .B1(n8387), .B2(n8388), .A(n8386), .ZN(n8389) );
  NAND2_X1 U5095 ( .A1(n7914), .A2(n9660), .ZN(n4648) );
  NAND2_X1 U5096 ( .A1(n7946), .A2(n7947), .ZN(n4635) );
  MUX2_X1 U5097 ( .A(n7945), .B(n7944), .S(n8046), .Z(n7946) );
  NOR2_X1 U5098 ( .A1(n4637), .A2(n6835), .ZN(n4636) );
  INV_X1 U5099 ( .A(n7939), .ZN(n4637) );
  MUX2_X1 U5100 ( .A(n4494), .B(n4493), .S(n7746), .Z(n7705) );
  OAI21_X1 U5101 ( .B1(n4442), .B2(n4643), .A(n8046), .ZN(n4640) );
  OAI21_X1 U5102 ( .B1(n7716), .B2(n7715), .A(n4508), .ZN(n7722) );
  AND2_X1 U5103 ( .A1(n4829), .A2(n4455), .ZN(n4508) );
  NAND2_X1 U5104 ( .A1(n4832), .A2(n7735), .ZN(n7749) );
  NAND2_X1 U5105 ( .A1(n7734), .A2(n7733), .ZN(n4832) );
  OAI21_X1 U5106 ( .B1(n7522), .B2(n7521), .A(n7520), .ZN(n7552) );
  NAND2_X1 U5107 ( .A1(n5026), .A2(n5025), .ZN(n5029) );
  AOI21_X1 U5108 ( .B1(n4520), .B2(n5007), .A(n5273), .ZN(n4519) );
  NAND2_X1 U5109 ( .A1(n4677), .A2(n8191), .ZN(n4673) );
  OR2_X1 U5110 ( .A1(n7909), .A2(n7908), .ZN(n8048) );
  OR2_X1 U5111 ( .A1(n8415), .A2(n8426), .ZN(n8034) );
  NAND2_X1 U5112 ( .A1(n4527), .A2(n4526), .ZN(n8496) );
  AND2_X1 U5113 ( .A1(n7502), .A2(n8003), .ZN(n4526) );
  OR2_X1 U5114 ( .A1(n7353), .A2(n9963), .ZN(n7395) );
  OR2_X1 U5115 ( .A1(n8692), .A2(n8598), .ZN(n7984) );
  OR2_X1 U5116 ( .A1(n7222), .A2(n7244), .ZN(n7971) );
  OR2_X1 U5117 ( .A1(n7026), .A2(n6974), .ZN(n7961) );
  AND2_X1 U5118 ( .A1(n6991), .A2(n7947), .ZN(n4882) );
  OR2_X1 U5119 ( .A1(n8277), .A2(n9717), .ZN(n7918) );
  NAND2_X1 U5120 ( .A1(n5931), .A2(n4678), .ZN(n6077) );
  AND2_X1 U5121 ( .A1(n4464), .A2(n4679), .ZN(n4678) );
  INV_X1 U5122 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4679) );
  AND2_X1 U5123 ( .A1(n5838), .A2(n5954), .ZN(n5839) );
  INV_X1 U5124 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5838) );
  INV_X1 U5125 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5126 ( .A1(n6869), .A2(n5672), .ZN(n5673) );
  AND2_X1 U5127 ( .A1(n5662), .A2(n5661), .ZN(n5686) );
  INV_X1 U5128 ( .A(n8861), .ZN(n4950) );
  INV_X1 U5129 ( .A(n8808), .ZN(n4548) );
  OR2_X1 U5130 ( .A1(n4545), .A2(n8735), .ZN(n4544) );
  INV_X1 U5131 ( .A(n5784), .ZN(n4545) );
  OAI21_X1 U5132 ( .B1(n4548), .B2(n4545), .A(n8782), .ZN(n4543) );
  NAND2_X1 U5133 ( .A1(n7742), .A2(n7622), .ZN(n7819) );
  NOR2_X1 U5134 ( .A1(n7724), .A2(n4824), .ZN(n4823) );
  AND2_X1 U5135 ( .A1(n8944), .A2(n8959), .ZN(n7790) );
  INV_X1 U5136 ( .A(n9150), .ZN(n5779) );
  NAND2_X1 U5137 ( .A1(n5458), .A2(n4405), .ZN(n7772) );
  NAND2_X1 U5138 ( .A1(n9043), .A2(n9044), .ZN(n4799) );
  OR2_X1 U5139 ( .A1(n5418), .A2(n5417), .ZN(n5429) );
  NOR2_X1 U5140 ( .A1(n9186), .A2(n9191), .ZN(n4574) );
  NOR2_X1 U5141 ( .A1(n4591), .A2(n7276), .ZN(n4590) );
  INV_X1 U5142 ( .A(n4592), .ZN(n4591) );
  INV_X1 U5143 ( .A(n7209), .ZN(n4812) );
  INV_X1 U5144 ( .A(n7586), .ZN(n4778) );
  AOI21_X1 U5145 ( .B1(n4782), .B2(n4781), .A(n4780), .ZN(n4779) );
  INV_X1 U5146 ( .A(n7632), .ZN(n4780) );
  INV_X1 U5147 ( .A(n4788), .ZN(n4781) );
  NOR2_X1 U5148 ( .A1(n4579), .A2(n7018), .ZN(n4578) );
  NAND2_X1 U5149 ( .A1(n4505), .A2(n7758), .ZN(n4504) );
  INV_X1 U5150 ( .A(n7657), .ZN(n4505) );
  XNOR2_X1 U5151 ( .A(n5162), .B(n5613), .ZN(n4724) );
  NOR2_X1 U5152 ( .A1(n5619), .A2(n6452), .ZN(n6455) );
  NOR2_X1 U5153 ( .A1(n9106), .A2(n9196), .ZN(n9105) );
  INV_X1 U5154 ( .A(n4724), .ZN(n6451) );
  INV_X1 U5155 ( .A(n5322), .ZN(n4498) );
  OAI21_X1 U5156 ( .B1(n5466), .B2(n5465), .A(n5086), .ZN(n5477) );
  NAND2_X1 U5157 ( .A1(n5078), .A2(n5077), .ZN(n5456) );
  NAND2_X1 U5158 ( .A1(n5446), .A2(n5445), .ZN(n5078) );
  AND2_X1 U5159 ( .A1(n5064), .A2(n5063), .ZN(n5413) );
  AOI21_X1 U5160 ( .B1(n4864), .B2(n4862), .A(n4471), .ZN(n4861) );
  INV_X1 U5161 ( .A(n5052), .ZN(n4862) );
  NAND2_X1 U5162 ( .A1(n5048), .A2(n5047), .ZN(n5374) );
  NAND2_X1 U5163 ( .A1(n4839), .A2(n4837), .ZN(n5334) );
  AOI21_X1 U5164 ( .B1(n4840), .B2(n4410), .A(n4838), .ZN(n4837) );
  INV_X1 U5165 ( .A(n4978), .ZN(n4838) );
  NOR2_X1 U5166 ( .A1(n5024), .A2(n4845), .ZN(n4844) );
  INV_X1 U5167 ( .A(n5017), .ZN(n4845) );
  INV_X1 U5168 ( .A(n4519), .ZN(n4518) );
  AOI21_X1 U5169 ( .B1(n4519), .B2(n4517), .A(n4516), .ZN(n4515) );
  INV_X1 U5170 ( .A(n5012), .ZN(n4516) );
  INV_X1 U5171 ( .A(n5007), .ZN(n4517) );
  INV_X1 U5172 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5173 ( .A1(n4866), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4803) );
  INV_X1 U5174 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4867) );
  OAI21_X2 U5175 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n4865), .ZN(n4802) );
  INV_X1 U5176 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4865) );
  AOI22_X1 U5177 ( .A1(n7231), .A2(n7230), .B1(n7229), .B2(n7228), .ZN(n7232)
         );
  INV_X1 U5178 ( .A(n8184), .ZN(n4704) );
  AND2_X1 U5179 ( .A1(n4421), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U5180 ( .A1(n8178), .A2(n8251), .ZN(n4701) );
  AOI21_X1 U5181 ( .B1(n4675), .B2(n4677), .A(n4443), .ZN(n4674) );
  INV_X1 U5182 ( .A(n8167), .ZN(n4675) );
  NAND2_X1 U5183 ( .A1(n4718), .A2(n4711), .ZN(n4710) );
  NOR2_X1 U5184 ( .A1(n4717), .A2(n4715), .ZN(n4711) );
  OR2_X1 U5185 ( .A1(n6961), .A2(n4717), .ZN(n4709) );
  NAND2_X1 U5186 ( .A1(n4720), .A2(n4706), .ZN(n4705) );
  NOR2_X1 U5187 ( .A1(n4716), .A2(n6653), .ZN(n4706) );
  NAND2_X1 U5188 ( .A1(n8168), .A2(n8167), .ZN(n8166) );
  INV_X1 U5189 ( .A(n6961), .ZN(n4716) );
  NAND2_X1 U5190 ( .A1(n6961), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5191 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  INV_X1 U5192 ( .A(n4687), .ZN(n4684) );
  OR2_X1 U5193 ( .A1(n8200), .A2(n8201), .ZN(n8138) );
  NAND2_X1 U5194 ( .A1(n7103), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7190) );
  INV_X1 U5195 ( .A(n7104), .ZN(n7103) );
  AND2_X1 U5196 ( .A1(n7224), .A2(n7223), .ZN(n7310) );
  NAND2_X1 U5197 ( .A1(n7897), .A2(n4522), .ZN(n7902) );
  INV_X1 U5198 ( .A(n8039), .ZN(n4522) );
  AND2_X1 U5199 ( .A1(n8048), .A2(n8038), .ZN(n8083) );
  AND3_X1 U5200 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(n8161) );
  INV_X1 U5201 ( .A(n6111), .ZN(n7389) );
  NOR2_X1 U5202 ( .A1(n6284), .A2(n4605), .ZN(n6261) );
  AND2_X1 U5203 ( .A1(n6244), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4605) );
  OR2_X1 U5204 ( .A1(n6261), .A2(n6260), .ZN(n4604) );
  OR2_X1 U5205 ( .A1(n6239), .A2(n6238), .ZN(n4601) );
  AND2_X1 U5206 ( .A1(n4601), .A2(n4600), .ZN(n8288) );
  NAND2_X1 U5207 ( .A1(n6275), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4600) );
  OR2_X1 U5208 ( .A1(n8288), .A2(n8289), .ZN(n4599) );
  NOR2_X1 U5209 ( .A1(n6390), .A2(n4470), .ZN(n8300) );
  NOR2_X1 U5210 ( .A1(n8300), .A2(n8301), .ZN(n8299) );
  NAND2_X1 U5211 ( .A1(n8320), .A2(n4593), .ZN(n8333) );
  OR2_X1 U5212 ( .A1(n8322), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4593) );
  NOR2_X1 U5213 ( .A1(n8374), .A2(n4594), .ZN(n8387) );
  AND2_X1 U5214 ( .A1(n8375), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4594) );
  OR2_X1 U5215 ( .A1(n7457), .A2(n7456), .ZN(n7482) );
  AND2_X1 U5216 ( .A1(n8466), .A2(n4456), .ZN(n8403) );
  NAND2_X1 U5217 ( .A1(n8466), .A2(n4617), .ZN(n8411) );
  NAND2_X1 U5218 ( .A1(n8034), .A2(n8035), .ZN(n8416) );
  AND2_X1 U5219 ( .A1(n8416), .A2(n4901), .ZN(n4900) );
  OR2_X1 U5220 ( .A1(n8430), .A2(n4902), .ZN(n4901) );
  INV_X1 U5221 ( .A(n7452), .ZN(n4902) );
  OR2_X1 U5222 ( .A1(n8645), .A2(n8427), .ZN(n7439) );
  NAND2_X1 U5223 ( .A1(n7504), .A2(n4874), .ZN(n8443) );
  NOR2_X1 U5224 ( .A1(n8446), .A2(n4875), .ZN(n4874) );
  INV_X1 U5225 ( .A(n8019), .ZN(n4875) );
  NAND2_X1 U5226 ( .A1(n8463), .A2(n8462), .ZN(n7504) );
  NAND2_X1 U5227 ( .A1(n8483), .A2(n8017), .ZN(n8463) );
  NAND2_X1 U5228 ( .A1(n4910), .A2(n4909), .ZN(n8458) );
  AOI21_X1 U5229 ( .B1(n4911), .B2(n4912), .A(n8462), .ZN(n4909) );
  OR2_X1 U5230 ( .A1(n8490), .A2(n8653), .ZN(n8474) );
  AND2_X1 U5231 ( .A1(n8017), .A2(n8014), .ZN(n8480) );
  NAND2_X1 U5232 ( .A1(n8489), .A2(n8497), .ZN(n8488) );
  NAND2_X1 U5233 ( .A1(n7501), .A2(n4525), .ZN(n4527) );
  NOR2_X1 U5234 ( .A1(n8526), .A2(n4528), .ZN(n4525) );
  INV_X1 U5235 ( .A(n8001), .ZN(n4528) );
  OR2_X1 U5236 ( .A1(n8675), .A2(n8555), .ZN(n8001) );
  NOR2_X1 U5237 ( .A1(n8553), .A2(n4886), .ZN(n4885) );
  INV_X1 U5238 ( .A(n7992), .ZN(n4886) );
  AND2_X1 U5239 ( .A1(n7992), .A2(n7990), .ZN(n8569) );
  OR2_X1 U5240 ( .A1(n8692), .A2(n8572), .ZN(n4933) );
  INV_X1 U5241 ( .A(n8603), .ZN(n4931) );
  NOR2_X1 U5242 ( .A1(n7198), .A2(n7222), .ZN(n7199) );
  OR2_X1 U5243 ( .A1(n7087), .A2(n9325), .ZN(n7198) );
  AOI21_X1 U5244 ( .B1(n4441), .B2(n7029), .A(n4407), .ZN(n4916) );
  AND2_X1 U5245 ( .A1(n7957), .A2(n7963), .ZN(n8072) );
  NAND2_X1 U5246 ( .A1(n7029), .A2(n7027), .ZN(n4918) );
  INV_X1 U5247 ( .A(n7028), .ZN(n4920) );
  INV_X1 U5248 ( .A(n7027), .ZN(n4919) );
  NAND2_X1 U5249 ( .A1(n6883), .A2(n8068), .ZN(n7028) );
  NAND2_X1 U5250 ( .A1(n6847), .A2(n6846), .ZN(n7885) );
  OAI211_X1 U5251 ( .C1(n6423), .C2(n6369), .A(n6368), .B(n6367), .ZN(n9614)
         );
  AND2_X1 U5252 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6320) );
  INV_X1 U5253 ( .A(n9613), .ZN(n8573) );
  AND2_X1 U5254 ( .A1(n8086), .A2(n7911), .ZN(n9644) );
  NAND2_X1 U5255 ( .A1(n7901), .A2(n7900), .ZN(n8625) );
  NAND2_X1 U5256 ( .A1(n7394), .A2(n7393), .ZN(n8663) );
  NAND2_X1 U5257 ( .A1(n7360), .A2(n7359), .ZN(n8682) );
  AND2_X1 U5258 ( .A1(n6087), .A2(n6133), .ZN(n9752) );
  NAND2_X1 U5259 ( .A1(n9683), .A2(n6120), .ZN(n8700) );
  OR2_X1 U5260 ( .A1(n6199), .A2(n9684), .ZN(n8702) );
  NOR2_X1 U5261 ( .A1(n8623), .A2(n8622), .ZN(n8704) );
  XNOR2_X1 U5262 ( .A(n5855), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6121) );
  OR2_X1 U5263 ( .A1(n4940), .A2(n4938), .ZN(n4937) );
  INV_X1 U5264 ( .A(n4476), .ZN(n4938) );
  INV_X1 U5265 ( .A(n4941), .ZN(n4940) );
  OAI21_X1 U5266 ( .B1(n8746), .B2(n4942), .A(n8816), .ZN(n4941) );
  NAND2_X1 U5267 ( .A1(n8834), .A2(n8837), .ZN(n4539) );
  NAND2_X1 U5268 ( .A1(n4476), .A2(n5754), .ZN(n4939) );
  NAND2_X1 U5269 ( .A1(n8806), .A2(n5784), .ZN(n8781) );
  INV_X1 U5270 ( .A(n4948), .ZN(n4947) );
  INV_X1 U5271 ( .A(n4946), .ZN(n4945) );
  OAI21_X1 U5272 ( .B1(n4949), .B2(n4947), .A(n8792), .ZN(n4946) );
  OR2_X1 U5273 ( .A1(n5732), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5274 ( .A1(n5732), .A2(n4950), .ZN(n4948) );
  OAI21_X1 U5275 ( .B1(n5776), .B2(n8825), .A(n5775), .ZN(n8734) );
  OAI22_X1 U5276 ( .A1(n6556), .A2(n5790), .B1(n9524), .B2(n5788), .ZN(n5647)
         );
  NAND2_X1 U5277 ( .A1(n6949), .A2(n8759), .ZN(n5666) );
  NAND2_X1 U5278 ( .A1(n4480), .A2(n4479), .ZN(n4538) );
  INV_X1 U5279 ( .A(n5746), .ZN(n4479) );
  INV_X1 U5280 ( .A(n5747), .ZN(n4480) );
  OR2_X1 U5281 ( .A1(n5864), .A2(n7832), .ZN(n5815) );
  NAND2_X1 U5282 ( .A1(n7281), .A2(n7284), .ZN(n4534) );
  INV_X1 U5283 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5506) );
  AND4_X1 U5284 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n7143)
         );
  NAND2_X1 U5285 ( .A1(n6012), .A2(n6013), .ZN(n6011) );
  OR2_X1 U5286 ( .A1(n9450), .A2(n9449), .ZN(n4564) );
  AND2_X1 U5287 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  INV_X1 U5288 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4968) );
  OR2_X1 U5289 ( .A1(n7161), .A2(n7160), .ZN(n4557) );
  NOR2_X1 U5290 ( .A1(n8940), .A2(n4580), .ZN(n8917) );
  INV_X1 U5291 ( .A(n4582), .ZN(n4580) );
  NAND2_X1 U5292 ( .A1(n7619), .A2(n4582), .ZN(n4581) );
  NOR2_X1 U5293 ( .A1(n7790), .A2(n4821), .ZN(n4820) );
  NOR2_X1 U5294 ( .A1(n7790), .A2(n4826), .ZN(n8946) );
  AOI21_X1 U5295 ( .B1(n4761), .B2(n4765), .A(n4439), .ZN(n4759) );
  AOI21_X1 U5296 ( .B1(n4399), .B2(n4764), .A(n4451), .ZN(n4763) );
  AND2_X1 U5297 ( .A1(n7709), .A2(n7772), .ZN(n8967) );
  AOI21_X1 U5298 ( .B1(n4793), .B2(n4796), .A(n4791), .ZN(n4790) );
  INV_X1 U5299 ( .A(n7703), .ZN(n4791) );
  AND2_X1 U5300 ( .A1(n4800), .A2(n4794), .ZN(n4793) );
  AND2_X1 U5301 ( .A1(n9014), .A2(n9035), .ZN(n4800) );
  NAND2_X1 U5302 ( .A1(n4797), .A2(n4795), .ZN(n4794) );
  INV_X1 U5303 ( .A(n9044), .ZN(n4795) );
  INV_X1 U5304 ( .A(n4797), .ZN(n4796) );
  OR2_X1 U5305 ( .A1(n9023), .A2(n9165), .ZN(n9008) );
  NAND2_X1 U5306 ( .A1(n4799), .A2(n4797), .ZN(n9030) );
  AND4_X1 U5307 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n9046)
         );
  OAI22_X1 U5308 ( .A1(n9070), .A2(n5583), .B1(n9088), .B2(n9079), .ZN(n9055)
         );
  OR2_X1 U5309 ( .A1(n5367), .A2(n5121), .ZN(n5378) );
  NAND2_X1 U5310 ( .A1(n4804), .A2(n4807), .ZN(n9099) );
  INV_X1 U5311 ( .A(n4808), .ZN(n4807) );
  OAI21_X1 U5312 ( .B1(n4415), .B2(n4809), .A(n7644), .ZN(n4808) );
  AOI21_X1 U5313 ( .B1(n4751), .B2(n4397), .A(n4754), .ZN(n4750) );
  AND2_X1 U5314 ( .A1(n7579), .A2(n7585), .ZN(n7807) );
  NAND2_X1 U5315 ( .A1(n5579), .A2(n5578), .ZN(n7208) );
  OAI21_X1 U5316 ( .B1(n4734), .B2(n4731), .A(n4730), .ZN(n7141) );
  NOR2_X1 U5317 ( .A1(n4733), .A2(n4427), .ZN(n4730) );
  INV_X1 U5318 ( .A(n5185), .ZN(n5404) );
  AOI21_X1 U5319 ( .B1(n5574), .B2(n4739), .A(n4738), .ZN(n4737) );
  INV_X1 U5320 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5321 ( .B1(n4728), .B2(n5566), .A(n6537), .ZN(n4726) );
  NAND2_X1 U5322 ( .A1(n4729), .A2(n5566), .ZN(n6709) );
  INV_X1 U5323 ( .A(n6711), .ZN(n4729) );
  NAND2_X1 U5324 ( .A1(n4723), .A2(n6451), .ZN(n4722) );
  INV_X1 U5325 ( .A(n6455), .ZN(n4723) );
  INV_X1 U5326 ( .A(n9256), .ZN(n9065) );
  INV_X1 U5327 ( .A(n9104), .ZN(n9251) );
  NAND2_X1 U5328 ( .A1(n4744), .A2(n4412), .ZN(n8902) );
  NAND2_X1 U5329 ( .A1(n4744), .A2(n4742), .ZN(n5596) );
  INV_X1 U5330 ( .A(n8944), .ZN(n9139) );
  NAND2_X1 U5331 ( .A1(n5468), .A2(n5467), .ZN(n9144) );
  INV_X1 U5332 ( .A(n9546), .ZN(n9529) );
  OR2_X1 U5333 ( .A1(n6603), .A2(n7832), .ZN(n9546) );
  NAND2_X1 U5334 ( .A1(n5560), .A2(n9217), .ZN(n6461) );
  NAND2_X1 U5335 ( .A1(n5815), .A2(n7835), .ZN(n6462) );
  XNOR2_X1 U5336 ( .A(n7522), .B(n7472), .ZN(n7513) );
  NAND2_X1 U5337 ( .A1(n5098), .A2(n5097), .ZN(n7467) );
  NAND2_X1 U5338 ( .A1(n5488), .A2(n5489), .ZN(n5098) );
  XNOR2_X1 U5339 ( .A(n5532), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5558) );
  NOR2_X1 U5340 ( .A1(n4430), .A2(n4965), .ZN(n4964) );
  OAI21_X1 U5341 ( .B1(n5018), .B2(n4410), .A(n4840), .ZN(n5321) );
  XNOR2_X1 U5342 ( .A(n5302), .B(n5301), .ZN(n6655) );
  NAND2_X1 U5343 ( .A1(n5018), .A2(n5017), .ZN(n5302) );
  AND2_X1 U5344 ( .A1(n5001), .A2(SI_6_), .ZN(n4406) );
  INV_X1 U5345 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U5346 ( .A1(n4487), .A2(n4999), .ZN(n5214) );
  NAND2_X1 U5347 ( .A1(n5100), .A2(n4488), .ZN(n4954) );
  INV_X1 U5348 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4488) );
  XNOR2_X1 U5349 ( .A(n4985), .B(n4984), .ZN(n5157) );
  NAND2_X1 U5350 ( .A1(n7443), .A2(n7442), .ZN(n8638) );
  NAND2_X1 U5351 ( .A1(n9566), .A2(n6576), .ZN(n6654) );
  NOR2_X1 U5352 ( .A1(n4703), .A2(n4699), .ZN(n4698) );
  INV_X1 U5353 ( .A(n8185), .ZN(n4699) );
  INV_X1 U5354 ( .A(n8186), .ZN(n4703) );
  OAI211_X1 U5355 ( .C1(n4667), .C2(n4402), .A(n4668), .B(n4665), .ZN(n6568)
         );
  OR2_X1 U5356 ( .A1(n6499), .A2(n6498), .ZN(n4668) );
  OR2_X1 U5357 ( .A1(n4402), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U5358 ( .A1(n7383), .A2(n7382), .ZN(n8668) );
  NAND2_X1 U5359 ( .A1(n7418), .A2(n7417), .ZN(n8650) );
  NAND2_X1 U5360 ( .A1(n7307), .A2(n7306), .ZN(n8695) );
  NAND2_X1 U5361 ( .A1(n9568), .A2(n9567), .ZN(n9566) );
  NAND2_X1 U5362 ( .A1(n7372), .A2(n7371), .ZN(n8685) );
  NAND2_X1 U5363 ( .A1(n6746), .A2(n6143), .ZN(n9611) );
  NAND2_X1 U5364 ( .A1(n7451), .A2(n7450), .ZN(n8419) );
  NAND2_X1 U5365 ( .A1(n6145), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U5366 ( .A(n4602), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U5367 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4602) );
  NAND2_X1 U5368 ( .A1(n8393), .A2(n4611), .ZN(n4610) );
  INV_X1 U5369 ( .A(n4612), .ZN(n4611) );
  OAI21_X1 U5370 ( .B1(n8395), .B2(n8394), .A(n9595), .ZN(n4612) );
  NAND2_X1 U5371 ( .A1(n4609), .A2(n4608), .ZN(n4607) );
  INV_X1 U5372 ( .A(n8397), .ZN(n4608) );
  NAND2_X1 U5373 ( .A1(n9600), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4609) );
  AND2_X1 U5374 ( .A1(n4972), .A2(n4890), .ZN(n4889) );
  OAI21_X1 U5375 ( .B1(n7897), .B2(n8039), .A(n4892), .ZN(n4891) );
  NAND2_X1 U5376 ( .A1(n8399), .A2(n8261), .ZN(n4890) );
  OR2_X1 U5377 ( .A1(n9669), .A2(n6751), .ZN(n9676) );
  AND2_X1 U5378 ( .A1(n6197), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9690) );
  NAND2_X1 U5379 ( .A1(n4659), .A2(n4663), .ZN(n6084) );
  NAND2_X1 U5380 ( .A1(n4662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  INV_X1 U5381 ( .A(n5168), .ZN(n5866) );
  NAND2_X1 U5382 ( .A1(n5448), .A2(n5447), .ZN(n9156) );
  AND2_X1 U5383 ( .A1(n5515), .A2(n5129), .ZN(n8766) );
  AND4_X1 U5384 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n8984)
         );
  AND2_X1 U5385 ( .A1(n5487), .A2(n5486), .ZN(n8786) );
  INV_X1 U5386 ( .A(n9028), .ZN(n9169) );
  AND3_X1 U5387 ( .A1(n5475), .A2(n5474), .A3(n5473), .ZN(n8853) );
  INV_X1 U5388 ( .A(n5598), .ZN(n7831) );
  INV_X1 U5389 ( .A(n8853), .ZN(n8969) );
  OAI21_X1 U5390 ( .B1(n7541), .B2(n9488), .A(n4567), .ZN(n4566) );
  AOI21_X1 U5391 ( .B1(n7542), .B2(n9496), .A(n9483), .ZN(n4567) );
  NOR2_X1 U5392 ( .A1(n9481), .A2(n7544), .ZN(n4569) );
  INV_X1 U5393 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7544) );
  AOI21_X1 U5394 ( .B1(n8721), .B2(n7560), .A(n7559), .ZN(n9116) );
  NAND2_X1 U5395 ( .A1(n7524), .A2(n7523), .ZN(n9342) );
  OR2_X1 U5396 ( .A1(n9133), .A2(n9114), .ZN(n5606) );
  OR2_X1 U5397 ( .A1(n9534), .A2(n5542), .ZN(n9506) );
  OAI21_X1 U5398 ( .B1(n7929), .B2(n8046), .A(n4486), .ZN(n7930) );
  NAND2_X1 U5399 ( .A1(n7919), .A2(n8046), .ZN(n4486) );
  NAND2_X1 U5400 ( .A1(n4647), .A2(n4646), .ZN(n7925) );
  NOR2_X1 U5401 ( .A1(n7915), .A2(n8046), .ZN(n4646) );
  NAND2_X1 U5402 ( .A1(n4648), .A2(n7924), .ZN(n4647) );
  NAND2_X1 U5403 ( .A1(n7950), .A2(n7951), .ZN(n4633) );
  OAI21_X1 U5404 ( .B1(n7995), .B2(n7991), .A(n4485), .ZN(n4484) );
  INV_X1 U5405 ( .A(n7994), .ZN(n4485) );
  OAI21_X1 U5406 ( .B1(n7705), .B2(n7704), .A(n7703), .ZN(n4492) );
  NAND2_X1 U5407 ( .A1(n4830), .A2(n7746), .ZN(n4829) );
  OR2_X1 U5408 ( .A1(n7714), .A2(n7713), .ZN(n4830) );
  NOR2_X1 U5409 ( .A1(n4643), .A2(n4437), .ZN(n4641) );
  OAI22_X1 U5410 ( .A1(n7722), .A2(n9139), .B1(n7750), .B2(n7717), .ZN(n7718)
         );
  OR2_X1 U5411 ( .A1(n6837), .A2(n9750), .ZN(n7948) );
  INV_X1 U5412 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5413 ( .A1(n7130), .A2(n5717), .ZN(n4956) );
  INV_X1 U5414 ( .A(n8774), .ZN(n4935) );
  AND2_X1 U5415 ( .A1(n7583), .A2(n8878), .ZN(n5580) );
  INV_X1 U5416 ( .A(n9249), .ZN(n4736) );
  NAND2_X1 U5417 ( .A1(n8997), .A2(n8990), .ZN(n4588) );
  INV_X1 U5418 ( .A(n4861), .ZN(n4858) );
  AND2_X1 U5419 ( .A1(n5335), .A2(n5333), .ZN(n5034) );
  INV_X1 U5420 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5019) );
  INV_X1 U5421 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5020) );
  INV_X1 U5422 ( .A(SI_10_), .ZN(n9948) );
  INV_X1 U5423 ( .A(n4414), .ZN(n4715) );
  AND2_X1 U5424 ( .A1(n8032), .A2(n4460), .ZN(n4656) );
  NAND2_X1 U5425 ( .A1(n8038), .A2(n4652), .ZN(n4651) );
  NOR2_X1 U5426 ( .A1(n8043), .A2(n8041), .ZN(n4652) );
  NOR2_X1 U5427 ( .A1(n8081), .A2(n4654), .ZN(n4653) );
  INV_X1 U5428 ( .A(n8036), .ZN(n4654) );
  OR2_X1 U5429 ( .A1(n7477), .A2(n6144), .ZN(n6148) );
  NOR2_X1 U5430 ( .A1(n4621), .A2(n4618), .ZN(n4617) );
  INV_X1 U5431 ( .A(n4619), .ZN(n4618) );
  INV_X1 U5432 ( .A(n8419), .ZN(n7912) );
  NOR2_X1 U5433 ( .A1(n8638), .A2(n8645), .ZN(n4619) );
  NOR2_X1 U5434 ( .A1(n8480), .A2(n4915), .ZN(n4913) );
  NOR2_X1 U5435 ( .A1(n8668), .A2(n8675), .ZN(n4627) );
  NAND2_X1 U5436 ( .A1(n7337), .A2(n7336), .ZN(n7353) );
  INV_X1 U5437 ( .A(n7373), .ZN(n7337) );
  NOR2_X1 U5438 ( .A1(n8610), .A2(n8695), .ZN(n4616) );
  NAND2_X1 U5439 ( .A1(n7101), .A2(n4878), .ZN(n4877) );
  AND2_X1 U5440 ( .A1(n7973), .A2(n7100), .ZN(n4878) );
  AND2_X1 U5441 ( .A1(n4879), .A2(n7975), .ZN(n4876) );
  NAND2_X1 U5442 ( .A1(n7973), .A2(n4880), .ZN(n4879) );
  INV_X1 U5443 ( .A(n7971), .ZN(n4880) );
  AND2_X1 U5444 ( .A1(n8054), .A2(n9606), .ZN(n7929) );
  NAND2_X1 U5445 ( .A1(n8278), .A2(n9709), .ZN(n7928) );
  NAND2_X1 U5446 ( .A1(n6754), .A2(n4631), .ZN(n6840) );
  OR2_X1 U5447 ( .A1(n8474), .A2(n8650), .ZN(n8451) );
  INV_X1 U5448 ( .A(n8451), .ZN(n8466) );
  AOI21_X1 U5449 ( .B1(n6836), .B2(n6835), .A(n4979), .ZN(n6838) );
  INV_X1 U5450 ( .A(n6077), .ZN(n6076) );
  INV_X1 U5451 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5949) );
  OR2_X1 U5452 ( .A1(n5886), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5890) );
  INV_X1 U5453 ( .A(n7847), .ZN(n4549) );
  INV_X1 U5454 ( .A(n5682), .ZN(n4550) );
  XNOR2_X1 U5455 ( .A(n5616), .B(n5777), .ZN(n5627) );
  OAI21_X1 U5456 ( .B1(n5788), .B2(n9507), .A(n5614), .ZN(n5616) );
  NAND2_X1 U5457 ( .A1(n5768), .A2(n5767), .ZN(n5774) );
  AOI21_X1 U5458 ( .B1(n7749), .B2(n9122), .A(n4831), .ZN(n7744) );
  NAND2_X1 U5459 ( .A1(n7783), .A2(n7739), .ZN(n4831) );
  OAI21_X1 U5460 ( .B1(n7749), .B2(n4507), .A(n7788), .ZN(n7751) );
  NAND2_X1 U5461 ( .A1(n7783), .A2(n8874), .ZN(n4507) );
  INV_X1 U5462 ( .A(SI_15_), .ZN(n10047) );
  INV_X1 U5463 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5464 ( .A1(n4583), .A2(n9130), .ZN(n4582) );
  OR2_X1 U5465 ( .A1(n8919), .A2(n9134), .ZN(n4583) );
  OR2_X1 U5466 ( .A1(n9130), .A2(n8904), .ZN(n8907) );
  OAI21_X1 U5467 ( .B1(n4759), .B2(n7814), .A(n4469), .ZN(n4757) );
  NAND2_X1 U5468 ( .A1(n4587), .A2(n5779), .ZN(n4586) );
  INV_X1 U5469 ( .A(n4588), .ZN(n4587) );
  AND2_X1 U5470 ( .A1(n9159), .A2(n8984), .ZN(n7791) );
  OR2_X1 U5471 ( .A1(n9159), .A2(n8984), .ZN(n7792) );
  INV_X1 U5472 ( .A(n4809), .ZN(n4805) );
  INV_X1 U5473 ( .A(n5580), .ZN(n4749) );
  NOR2_X1 U5474 ( .A1(n4751), .A2(n5580), .ZN(n4747) );
  NAND2_X1 U5475 ( .A1(n4450), .A2(n7579), .ZN(n4811) );
  NOR2_X1 U5476 ( .A1(n7215), .A2(n7151), .ZN(n4592) );
  NOR2_X1 U5477 ( .A1(n4736), .A2(n5576), .ZN(n4735) );
  NOR2_X1 U5478 ( .A1(n4737), .A2(n4736), .ZN(n4733) );
  NOR2_X1 U5479 ( .A1(n4789), .A2(n6759), .ZN(n4788) );
  INV_X1 U5480 ( .A(n7627), .ZN(n4789) );
  INV_X1 U5481 ( .A(n6912), .ZN(n4577) );
  NAND2_X1 U5482 ( .A1(n7625), .A2(n7796), .ZN(n5246) );
  NAND2_X1 U5483 ( .A1(n8883), .A2(n7857), .ZN(n7661) );
  NAND2_X1 U5484 ( .A1(n7857), .A2(n6914), .ZN(n4579) );
  NAND2_X1 U5485 ( .A1(n8884), .A2(n6914), .ZN(n7660) );
  NOR2_X1 U5486 ( .A1(n9008), .A2(n4588), .ZN(n8985) );
  NAND2_X1 U5487 ( .A1(n9105), .A2(n9095), .ZN(n9089) );
  NAND2_X1 U5488 ( .A1(n7755), .A2(n5403), .ZN(n7746) );
  NAND2_X1 U5489 ( .A1(n6726), .A2(n7657), .ZN(n4503) );
  NAND2_X1 U5490 ( .A1(n7550), .A2(SI_30_), .ZN(n7554) );
  XNOR2_X1 U5491 ( .A(n7552), .B(n7551), .ZN(n7549) );
  NAND2_X1 U5492 ( .A1(n7471), .A2(n7470), .ZN(n7522) );
  NAND2_X1 U5493 ( .A1(n7467), .A2(n7466), .ZN(n7471) );
  NAND2_X1 U5494 ( .A1(n4452), .A2(n4769), .ZN(n4768) );
  INV_X1 U5495 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4769) );
  INV_X1 U5496 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5110) );
  NOR2_X1 U5497 ( .A1(n4768), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4497) );
  INV_X1 U5498 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5530) );
  AND2_X1 U5499 ( .A1(n5091), .A2(n5090), .ZN(n5476) );
  OAI21_X1 U5500 ( .B1(n5456), .B2(n5082), .A(n5081), .ZN(n5466) );
  AND2_X1 U5501 ( .A1(n5109), .A2(n5539), .ZN(n4495) );
  INV_X1 U5502 ( .A(n5068), .ZN(n4851) );
  INV_X1 U5503 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5505) );
  OAI21_X1 U5504 ( .B1(n5347), .B2(n5346), .A(n5042), .ZN(n5360) );
  AND2_X1 U5505 ( .A1(n5047), .A2(n5046), .ZN(n5359) );
  INV_X1 U5506 ( .A(n5023), .ZN(n4842) );
  INV_X1 U5507 ( .A(n4841), .ZN(n4840) );
  OAI21_X1 U5508 ( .B1(n4844), .B2(n4410), .A(n5029), .ZN(n4841) );
  INV_X1 U5509 ( .A(n4836), .ZN(n4835) );
  OAI21_X1 U5510 ( .B1(n5215), .B2(n4406), .A(n5242), .ZN(n4836) );
  OR2_X1 U5511 ( .A1(n8168), .A2(n4673), .ZN(n4672) );
  AOI21_X1 U5512 ( .B1(n4690), .B2(n4688), .A(n8109), .ZN(n4687) );
  INV_X1 U5513 ( .A(n7315), .ZN(n4688) );
  AOI22_X1 U5514 ( .A1(n6213), .A2(n6212), .B1(n6211), .B2(n6210), .ZN(n6308)
         );
  OR2_X1 U5515 ( .A1(n7062), .A2(n7061), .ZN(n7104) );
  AND2_X1 U5516 ( .A1(n6132), .A2(n9681), .ZN(n6141) );
  XNOR2_X1 U5517 ( .A(n9229), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9226) );
  AND2_X1 U5518 ( .A1(n4604), .A2(n4603), .ZN(n6297) );
  NAND2_X1 U5519 ( .A1(n6234), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U5520 ( .A1(n6297), .A2(n6296), .ZN(n6295) );
  NOR2_X1 U5521 ( .A1(n8299), .A2(n4475), .ZN(n8313) );
  NOR2_X1 U5522 ( .A1(n8313), .A2(n8314), .ZN(n8312) );
  NOR2_X1 U5523 ( .A1(n8336), .A2(n8335), .ZN(n8338) );
  NAND2_X1 U5524 ( .A1(n8359), .A2(n4595), .ZN(n8362) );
  NAND2_X1 U5525 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  INV_X1 U5526 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n4596) );
  INV_X1 U5527 ( .A(n8360), .ZN(n4597) );
  NOR2_X1 U5528 ( .A1(n8362), .A2(n8361), .ZN(n8374) );
  AND2_X1 U5529 ( .A1(n7485), .A2(n8418), .ZN(n8039) );
  AND2_X1 U5530 ( .A1(n7482), .A2(n7458), .ZN(n8413) );
  OR2_X1 U5531 ( .A1(n7444), .A2(n8150), .ZN(n7457) );
  OR2_X1 U5532 ( .A1(n7419), .A2(n8204), .ZN(n7431) );
  INV_X1 U5533 ( .A(n4913), .ZN(n4912) );
  NAND2_X1 U5534 ( .A1(n8499), .A2(n4883), .ZN(n8483) );
  AND2_X1 U5535 ( .A1(n8480), .A2(n8013), .ZN(n4883) );
  AND2_X1 U5536 ( .A1(n8495), .A2(n4625), .ZN(n4624) );
  AND2_X1 U5537 ( .A1(n8668), .A2(n8537), .ZN(n4482) );
  NAND2_X1 U5538 ( .A1(n8556), .A2(n4627), .ZN(n8521) );
  AND2_X1 U5539 ( .A1(n8565), .A2(n8561), .ZN(n8556) );
  NAND2_X1 U5540 ( .A1(n8556), .A2(n8546), .ZN(n8541) );
  INV_X1 U5541 ( .A(n4927), .ZN(n4926) );
  OAI21_X1 U5542 ( .B1(n4403), .B2(n4928), .A(n4428), .ZN(n4927) );
  NAND2_X1 U5543 ( .A1(n7188), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7319) );
  NAND2_X1 U5544 ( .A1(n4616), .A2(n4615), .ZN(n8582) );
  INV_X1 U5545 ( .A(n4616), .ZN(n8612) );
  NAND2_X1 U5546 ( .A1(n7199), .A2(n9312), .ZN(n8610) );
  NAND2_X1 U5547 ( .A1(n7186), .A2(n7971), .ZN(n7494) );
  NAND2_X1 U5548 ( .A1(n7096), .A2(n7095), .ZN(n7222) );
  NAND2_X1 U5549 ( .A1(n7101), .A2(n7100), .ZN(n7186) );
  NAND2_X1 U5550 ( .A1(n6663), .A2(n6662), .ZN(n6968) );
  AND2_X1 U5551 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n6662) );
  INV_X1 U5552 ( .A(n6661), .ZN(n6663) );
  OR2_X1 U5553 ( .A1(n6968), .A2(n6967), .ZN(n7062) );
  AND2_X1 U5554 ( .A1(n4882), .A2(n7958), .ZN(n4881) );
  OAI21_X1 U5555 ( .B1(n7955), .B2(n4533), .A(n7957), .ZN(n4532) );
  INV_X1 U5556 ( .A(n7958), .ZN(n4533) );
  NAND2_X1 U5557 ( .A1(n7021), .A2(n7955), .ZN(n7080) );
  INV_X1 U5558 ( .A(n8269), .ZN(n7082) );
  NAND2_X1 U5559 ( .A1(n6885), .A2(n4882), .ZN(n7021) );
  NAND2_X1 U5560 ( .A1(n6506), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6577) );
  AND2_X1 U5561 ( .A1(n6438), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U5562 ( .A1(n9744), .A2(n7888), .ZN(n7045) );
  AND2_X1 U5563 ( .A1(n7887), .A2(n7891), .ZN(n7888) );
  AND2_X1 U5564 ( .A1(n6432), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6438) );
  NOR2_X1 U5565 ( .A1(n6833), .A2(n4908), .ZN(n4907) );
  INV_X1 U5566 ( .A(n6830), .ZN(n4908) );
  NOR2_X1 U5567 ( .A1(n6371), .A2(n10027), .ZN(n6432) );
  NOR2_X1 U5568 ( .A1(n9615), .A2(n9583), .ZN(n7887) );
  OR2_X1 U5569 ( .A1(n9755), .A2(n6081), .ZN(n8620) );
  NAND2_X1 U5570 ( .A1(n4623), .A2(n4622), .ZN(n9615) );
  NOR2_X1 U5571 ( .A1(n9630), .A2(n4395), .ZN(n4622) );
  INV_X1 U5572 ( .A(n9651), .ZN(n4623) );
  NAND2_X1 U5573 ( .A1(n7928), .A2(n6841), .ZN(n9643) );
  NAND2_X1 U5574 ( .A1(n8060), .A2(n7923), .ZN(n9660) );
  INV_X1 U5575 ( .A(n6815), .ZN(n6773) );
  INV_X1 U5576 ( .A(n9752), .ZN(n9778) );
  AND2_X1 U5577 ( .A1(n4463), .A2(n5905), .ZN(n4657) );
  INV_X1 U5578 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5907) );
  NOR2_X1 U5579 ( .A1(n5932), .A2(n8722), .ZN(n5933) );
  AND2_X1 U5580 ( .A1(n5932), .A2(n5905), .ZN(n4629) );
  NAND2_X1 U5581 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U5582 ( .A1(n5938), .A2(n5937), .ZN(n5841) );
  NAND2_X1 U5583 ( .A1(n5955), .A2(n5839), .ZN(n6188) );
  AND3_X1 U5584 ( .A1(n5949), .A2(n5966), .A3(n5837), .ZN(n5954) );
  INV_X1 U5585 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U5586 ( .A1(n5904), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5955) );
  AND2_X1 U5587 ( .A1(n5834), .A2(n4422), .ZN(n5923) );
  AND2_X1 U5588 ( .A1(n4897), .A2(n4896), .ZN(n5832) );
  NOR2_X1 U5589 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4897) );
  NOR2_X1 U5590 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4896) );
  CLKBUF_X1 U5591 ( .A(n5881), .Z(n5882) );
  AOI21_X1 U5592 ( .B1(n5631), .B2(n8753), .A(n5635), .ZN(n5637) );
  XNOR2_X1 U5593 ( .A(n5634), .B(n8756), .ZN(n5636) );
  OR2_X1 U5594 ( .A1(n5494), .A2(n5128), .ZN(n5515) );
  NAND2_X1 U5595 ( .A1(n5655), .A2(n5654), .ZN(n5672) );
  AND2_X1 U5596 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  INV_X1 U5597 ( .A(n6525), .ZN(n5650) );
  NAND2_X1 U5598 ( .A1(n6406), .A2(n6405), .ZN(n4951) );
  INV_X1 U5599 ( .A(n7119), .ZN(n4958) );
  NAND2_X1 U5600 ( .A1(n5124), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5439) );
  NAND3_X1 U5601 ( .A1(n4541), .A2(n4540), .A3(n4542), .ZN(n8780) );
  INV_X1 U5602 ( .A(n4543), .ZN(n4542) );
  OR2_X1 U5603 ( .A1(n8734), .A2(n4545), .ZN(n4540) );
  OR2_X1 U5604 ( .A1(n7828), .A2(n5403), .ZN(n4873) );
  NAND2_X1 U5605 ( .A1(n6011), .A2(n6000), .ZN(n9414) );
  NAND2_X1 U5606 ( .A1(n4555), .A2(n4554), .ZN(n9416) );
  INV_X1 U5607 ( .A(n9413), .ZN(n4554) );
  INV_X1 U5608 ( .A(n9414), .ZN(n4555) );
  AOI21_X1 U5609 ( .B1(n9416), .B2(n6002), .A(n6003), .ZN(n6024) );
  NAND2_X1 U5610 ( .A1(n4564), .A2(n4563), .ZN(n9461) );
  NAND2_X1 U5611 ( .A1(n9444), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4563) );
  OAI22_X1 U5612 ( .A1(n9461), .A2(n9462), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9457), .ZN(n6174) );
  NOR2_X1 U5613 ( .A1(n6473), .A2(n4562), .ZN(n6477) );
  AND2_X1 U5614 ( .A1(n6474), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4562) );
  NOR2_X1 U5615 ( .A1(n6477), .A2(n6476), .ZN(n6919) );
  NOR2_X1 U5616 ( .A1(n6919), .A2(n4559), .ZN(n6920) );
  NOR2_X1 U5617 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  AOI21_X1 U5618 ( .B1(n4816), .B2(n4819), .A(n4815), .ZN(n4814) );
  INV_X1 U5619 ( .A(n4820), .ZN(n4819) );
  AND2_X1 U5620 ( .A1(n8907), .A2(n8909), .ZN(n7816) );
  INV_X1 U5621 ( .A(n8932), .ZN(n8926) );
  OR2_X1 U5622 ( .A1(n8953), .A2(n9139), .ZN(n8940) );
  INV_X1 U5623 ( .A(n4755), .ZN(n8939) );
  OAI21_X1 U5624 ( .B1(n8993), .B2(n4758), .A(n4756), .ZN(n4755) );
  NAND2_X1 U5625 ( .A1(n4761), .A2(n8957), .ZN(n4758) );
  INV_X1 U5626 ( .A(n4757), .ZN(n4756) );
  NOR2_X1 U5627 ( .A1(n9008), .A2(n9159), .ZN(n8994) );
  AND2_X1 U5628 ( .A1(n4799), .A2(n4801), .ZN(n9033) );
  AND2_X1 U5629 ( .A1(n9105), .A2(n4570), .ZN(n9047) );
  NOR2_X1 U5630 ( .A1(n9176), .A2(n4572), .ZN(n4570) );
  OR2_X1 U5631 ( .A1(n5392), .A2(n5391), .ZN(n5407) );
  AND2_X1 U5632 ( .A1(n9179), .A2(n8875), .ZN(n5584) );
  NAND2_X1 U5633 ( .A1(n9105), .A2(n4574), .ZN(n4981) );
  NAND2_X1 U5634 ( .A1(n5122), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5392) );
  INV_X1 U5635 ( .A(n5378), .ZN(n5122) );
  AOI21_X1 U5636 ( .B1(n9085), .B2(n7679), .A(n7610), .ZN(n9072) );
  OR2_X1 U5637 ( .A1(n7641), .A2(n7640), .ZN(n9100) );
  INV_X1 U5638 ( .A(n4753), .ZN(n9098) );
  OAI21_X1 U5639 ( .B1(n7208), .B2(n4748), .A(n4746), .ZN(n4753) );
  AOI21_X1 U5640 ( .B1(n4750), .B2(n4747), .A(n4400), .ZN(n4746) );
  NAND2_X1 U5641 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5642 ( .A1(n9265), .A2(n4589), .ZN(n9106) );
  AND2_X1 U5643 ( .A1(n4590), .A2(n9345), .ZN(n4589) );
  NAND2_X1 U5644 ( .A1(n4806), .A2(n4811), .ZN(n7292) );
  NAND2_X1 U5645 ( .A1(n4812), .A2(n4415), .ZN(n4806) );
  OR2_X1 U5646 ( .A1(n5327), .A2(n5326), .ZN(n5340) );
  NAND2_X1 U5647 ( .A1(n9265), .A2(n4590), .ZN(n7296) );
  NAND2_X1 U5648 ( .A1(n4812), .A2(n7667), .ZN(n7266) );
  NAND2_X1 U5649 ( .A1(n9265), .A2(n4592), .ZN(n7273) );
  AOI21_X1 U5650 ( .B1(n4779), .B2(n4783), .A(n4778), .ZN(n4777) );
  NAND2_X1 U5651 ( .A1(n5118), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5315) );
  INV_X1 U5652 ( .A(n5294), .ZN(n5118) );
  AND2_X1 U5653 ( .A1(n9265), .A2(n7249), .ZN(n7213) );
  NAND2_X1 U5654 ( .A1(n4776), .A2(n4779), .ZN(n7142) );
  OR2_X1 U5655 ( .A1(n6699), .A2(n4783), .ZN(n4776) );
  NAND2_X1 U5656 ( .A1(n4784), .A2(n4401), .ZN(n9250) );
  NAND2_X1 U5657 ( .A1(n6699), .A2(n4788), .ZN(n4784) );
  NOR2_X1 U5658 ( .A1(n9264), .A2(n9263), .ZN(n9265) );
  NAND2_X1 U5659 ( .A1(n4785), .A2(n7627), .ZN(n6760) );
  OR2_X1 U5660 ( .A1(n6699), .A2(n5264), .ZN(n4785) );
  AND4_X1 U5661 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), .ZN(n6801)
         );
  NAND2_X1 U5662 ( .A1(n4577), .A2(n4578), .ZN(n6765) );
  AND2_X1 U5663 ( .A1(n7629), .A2(n7627), .ZN(n7801) );
  OR2_X1 U5664 ( .A1(n5571), .A2(n6896), .ZN(n6792) );
  NAND2_X1 U5665 ( .A1(n7661), .A2(n7625), .ZN(n7796) );
  NOR2_X1 U5666 ( .A1(n4579), .A2(n6912), .ZN(n6804) );
  OR2_X1 U5667 ( .A1(n6733), .A2(n5247), .ZN(n6912) );
  NOR2_X1 U5668 ( .A1(n6912), .A2(n5527), .ZN(n6911) );
  AOI21_X1 U5669 ( .B1(n4404), .B2(n4506), .A(n5248), .ZN(n4502) );
  AND4_X1 U5670 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n6904)
         );
  AND2_X1 U5671 ( .A1(n7761), .A2(n7656), .ZN(n6902) );
  OR2_X1 U5672 ( .A1(n6717), .A2(n7869), .ZN(n6719) );
  NOR2_X1 U5673 ( .A1(n6719), .A2(n5190), .ZN(n6734) );
  OR2_X1 U5674 ( .A1(n6462), .A2(n5562), .ZN(n6732) );
  NAND2_X1 U5675 ( .A1(n5377), .A2(n5376), .ZN(n9186) );
  INV_X1 U5676 ( .A(n9263), .ZN(n9274) );
  OAI211_X1 U5677 ( .C1(P1_B_REG_SCAN_IN), .C2(n6989), .A(n5558), .B(n5546), 
        .ZN(n6342) );
  XNOR2_X1 U5678 ( .A(n7549), .B(SI_30_), .ZN(n7898) );
  AND2_X1 U5679 ( .A1(n5537), .A2(n4766), .ZN(n5131) );
  NOR2_X1 U5680 ( .A1(n4768), .A2(n4767), .ZN(n4766) );
  NAND2_X1 U5681 ( .A1(n5112), .A2(n5539), .ZN(n4767) );
  INV_X1 U5682 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5683 ( .A1(n5092), .A2(n5091), .ZN(n5488) );
  NAND2_X1 U5684 ( .A1(n5477), .A2(n5476), .ZN(n5092) );
  AND2_X1 U5685 ( .A1(n5097), .A2(n5096), .ZN(n5489) );
  XNOR2_X1 U5686 ( .A(n4576), .B(n5112), .ZN(n9368) );
  NAND2_X1 U5687 ( .A1(n4500), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5688 ( .A1(n4498), .A2(n4496), .ZN(n4500) );
  AND2_X1 U5689 ( .A1(n4497), .A2(n5109), .ZN(n4496) );
  XNOR2_X1 U5690 ( .A(n5466), .B(n5465), .ZN(n7415) );
  NAND2_X1 U5691 ( .A1(n4846), .A2(n4847), .ZN(n5446) );
  INV_X1 U5692 ( .A(n4848), .ZN(n4847) );
  NAND2_X1 U5693 ( .A1(n5425), .A2(n4850), .ZN(n4846) );
  OAI21_X1 U5694 ( .B1(n5424), .B2(n4849), .A(n5072), .ZN(n4848) );
  AND2_X1 U5695 ( .A1(n5077), .A2(n5076), .ZN(n5445) );
  NAND2_X1 U5696 ( .A1(n4852), .A2(n5068), .ZN(n5436) );
  NAND2_X1 U5697 ( .A1(n4853), .A2(n5424), .ZN(n4852) );
  INV_X1 U5698 ( .A(n5425), .ZN(n4853) );
  NAND2_X1 U5699 ( .A1(n4859), .A2(n4861), .ZN(n5399) );
  NAND2_X1 U5700 ( .A1(n4860), .A2(n4864), .ZN(n4859) );
  INV_X1 U5701 ( .A(n5374), .ZN(n4860) );
  INV_X1 U5702 ( .A(n4965), .ZN(n4963) );
  NAND2_X1 U5703 ( .A1(n5362), .A2(n5361), .ZN(n5375) );
  NAND2_X1 U5704 ( .A1(n4843), .A2(n5023), .ZN(n5311) );
  NAND2_X1 U5705 ( .A1(n5018), .A2(n4844), .ZN(n4843) );
  AND2_X1 U5706 ( .A1(n5275), .A2(n5101), .ZN(n5288) );
  OAI21_X1 U5707 ( .B1(n5262), .B2(n4518), .A(n4515), .ZN(n5290) );
  INV_X1 U5708 ( .A(n4411), .ZN(n4520) );
  NAND2_X1 U5709 ( .A1(n4993), .A2(n4992), .ZN(n5202) );
  NAND2_X1 U5710 ( .A1(n5157), .A2(n5158), .ZN(n4521) );
  NAND2_X1 U5711 ( .A1(n9579), .A2(n6427), .ZN(n6501) );
  OR2_X1 U5712 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NOR2_X1 U5713 ( .A1(n6356), .A2(n6355), .ZN(n6354) );
  NAND2_X1 U5714 ( .A1(n4669), .A2(n4674), .ZN(n8192) );
  OR2_X1 U5715 ( .A1(n8168), .A2(n4676), .ZN(n4669) );
  NAND2_X1 U5716 ( .A1(n4705), .A2(n4712), .ZN(n7056) );
  NAND2_X1 U5717 ( .A1(n4710), .A2(n4709), .ZN(n6963) );
  NAND2_X1 U5718 ( .A1(n8136), .A2(n8135), .ZN(n8200) );
  NAND2_X1 U5719 ( .A1(n4691), .A2(n4690), .ZN(n8110) );
  NAND2_X1 U5720 ( .A1(n7316), .A2(n7315), .ZN(n4691) );
  NOR2_X1 U5721 ( .A1(n6364), .A2(n6363), .ZN(n6417) );
  NAND2_X1 U5722 ( .A1(n4685), .A2(n4687), .ZN(n8210) );
  NAND2_X1 U5723 ( .A1(n4686), .A2(n4690), .ZN(n4685) );
  INV_X1 U5724 ( .A(n7316), .ZN(n4686) );
  NAND2_X1 U5725 ( .A1(n7407), .A2(n7406), .ZN(n8653) );
  OAI22_X1 U5726 ( .A1(n6308), .A2(n6307), .B1(n6306), .B2(n6305), .ZN(n6319)
         );
  NOR2_X1 U5727 ( .A1(n6319), .A2(n6318), .ZN(n6364) );
  AOI22_X1 U5728 ( .A1(n6568), .A2(n6567), .B1(n6566), .B2(n6565), .ZN(n9568)
         );
  NAND2_X1 U5729 ( .A1(n8166), .A2(n8120), .ZN(n8225) );
  NAND2_X1 U5730 ( .A1(n4713), .A2(n7055), .ZN(n4707) );
  NAND2_X1 U5731 ( .A1(n7055), .A2(n4719), .ZN(n4708) );
  NAND2_X1 U5732 ( .A1(n4718), .A2(n4414), .ZN(n6962) );
  NAND2_X1 U5733 ( .A1(n4681), .A2(n4682), .ZN(n8242) );
  AOI21_X1 U5734 ( .B1(n4689), .B2(n4683), .A(n4409), .ZN(n4682) );
  NAND2_X1 U5735 ( .A1(n7316), .A2(n4683), .ZN(n4681) );
  NAND2_X1 U5736 ( .A1(n4667), .A2(n4666), .ZN(n9579) );
  AND2_X1 U5737 ( .A1(n4667), .A2(n4425), .ZN(n9580) );
  INV_X1 U5738 ( .A(n8250), .ZN(n9589) );
  NAND2_X1 U5739 ( .A1(n6136), .A2(n6135), .ZN(n9573) );
  INV_X1 U5740 ( .A(n9593), .ZN(n8258) );
  NAND2_X1 U5741 ( .A1(n7185), .A2(n7184), .ZN(n7364) );
  INV_X1 U5742 ( .A(n9573), .ZN(n9584) );
  XNOR2_X1 U5743 ( .A(n4531), .B(n6749), .ZN(n4530) );
  AOI21_X1 U5744 ( .B1(n7910), .B2(n8083), .A(n8042), .ZN(n4531) );
  INV_X1 U5745 ( .A(n7902), .ZN(n7904) );
  NAND2_X1 U5746 ( .A1(n8140), .A2(n7911), .ZN(n8093) );
  INV_X1 U5747 ( .A(n6824), .ZN(n8278) );
  CLKBUF_X1 U5748 ( .A(n6820), .Z(n8279) );
  INV_X2 U5749 ( .A(P2_U3966), .ZN(n8280) );
  AND2_X1 U5750 ( .A1(n5879), .A2(n5878), .ZN(n9240) );
  INV_X1 U5751 ( .A(n4604), .ZN(n6259) );
  INV_X1 U5752 ( .A(n4601), .ZN(n6270) );
  INV_X1 U5753 ( .A(n4599), .ZN(n8287) );
  NAND2_X1 U5754 ( .A1(n6428), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4598) );
  XNOR2_X1 U5755 ( .A(n8333), .B(n8334), .ZN(n8321) );
  NOR2_X1 U5756 ( .A1(n8321), .A2(n9317), .ZN(n8335) );
  INV_X1 U5757 ( .A(n8390), .ZN(n9598) );
  AOI21_X1 U5758 ( .B1(n8721), .B2(n7907), .A(n7906), .ZN(n8619) );
  INV_X1 U5759 ( .A(n8625), .ZN(n8404) );
  NAND2_X1 U5760 ( .A1(n8429), .A2(n7452), .ZN(n8409) );
  NAND2_X1 U5761 ( .A1(n7504), .A2(n8019), .ZN(n8445) );
  NAND2_X1 U5762 ( .A1(n8488), .A2(n4914), .ZN(n8473) );
  NAND2_X1 U5763 ( .A1(n4527), .A2(n8003), .ZN(n8512) );
  NAND2_X1 U5764 ( .A1(n7501), .A2(n8001), .ZN(n8527) );
  NAND2_X1 U5765 ( .A1(n7497), .A2(n7992), .ZN(n8552) );
  NAND2_X1 U5766 ( .A1(n8579), .A2(n4933), .ZN(n8564) );
  NOR2_X1 U5767 ( .A1(n8603), .A2(n7367), .ZN(n8580) );
  NAND2_X1 U5768 ( .A1(n7060), .A2(n7059), .ZN(n9325) );
  NAND2_X1 U5769 ( .A1(n7028), .A2(n4921), .ZN(n7074) );
  NOR2_X1 U5770 ( .A1(n4920), .A2(n4919), .ZN(n7030) );
  INV_X1 U5771 ( .A(n4918), .ZN(n4921) );
  NAND2_X1 U5772 ( .A1(n4529), .A2(n6657), .ZN(n7026) );
  NAND2_X1 U5773 ( .A1(n6655), .A2(n7907), .ZN(n4529) );
  NAND2_X1 U5774 ( .A1(n7885), .A2(n7937), .ZN(n7042) );
  NAND2_X1 U5775 ( .A1(n6831), .A2(n6830), .ZN(n7874) );
  OAI22_X1 U5776 ( .A1(n6089), .A2(n4895), .B1(n6090), .B2(n7555), .ZN(n4894)
         );
  INV_X1 U5777 ( .A(n9676), .ZN(n9638) );
  INV_X1 U5778 ( .A(n9673), .ZN(n9631) );
  AND2_X2 U5779 ( .A1(n8704), .A2(n8624), .ZN(n9803) );
  AND2_X2 U5780 ( .A1(n8704), .A2(n8703), .ZN(n9785) );
  NAND2_X1 U5781 ( .A1(n9682), .A2(n9681), .ZN(n9687) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7416) );
  XNOR2_X1 U5783 ( .A(n5858), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7174) );
  XNOR2_X1 U5784 ( .A(n5843), .B(n5845), .ZN(n7053) );
  NAND2_X1 U5785 ( .A1(n5842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U5786 ( .A1(n5861), .A2(n5860), .ZN(n5842) );
  INV_X1 U5787 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7392) );
  INV_X1 U5788 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7381) );
  INV_X1 U5789 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U5790 ( .A1(n4661), .A2(n4660), .ZN(n6080) );
  AOI21_X1 U5791 ( .B1(n4663), .B2(n8722), .A(n8722), .ZN(n4660) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6482) );
  INV_X1 U5793 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5970) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5953) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10108) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5946) );
  INV_X1 U5797 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5926) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10084) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5892) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6419) );
  OR2_X1 U5801 ( .A1(n5610), .A2(n5863), .ZN(n5974) );
  INV_X1 U5802 ( .A(n8877), .ZN(n9087) );
  INV_X1 U5803 ( .A(n4535), .ZN(n7283) );
  NAND2_X1 U5804 ( .A1(n5810), .A2(n4960), .ZN(n4959) );
  INV_X1 U5805 ( .A(n5796), .ZN(n4960) );
  AND2_X1 U5806 ( .A1(n5263), .A2(n4461), .ZN(n4553) );
  OR2_X1 U5807 ( .A1(n8745), .A2(n4939), .ZN(n4936) );
  NAND2_X1 U5808 ( .A1(n5427), .A2(n5426), .ZN(n9165) );
  INV_X1 U5809 ( .A(n8879), .ZN(n7126) );
  CLKBUF_X1 U5810 ( .A(n7118), .Z(n7119) );
  NAND2_X1 U5811 ( .A1(n4944), .A2(n4948), .ZN(n8791) );
  NAND2_X1 U5812 ( .A1(n5733), .A2(n4949), .ZN(n4944) );
  NAND2_X1 U5813 ( .A1(n4546), .A2(n8734), .ZN(n8809) );
  INV_X1 U5814 ( .A(n8852), .ZN(n8865) );
  NAND2_X1 U5815 ( .A1(n4951), .A2(n5646), .ZN(n6524) );
  AND4_X1 U5816 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n7144)
         );
  AND2_X1 U5817 ( .A1(n5278), .A2(n4977), .ZN(n5279) );
  NAND2_X1 U5818 ( .A1(n8744), .A2(n5754), .ZN(n8818) );
  NAND2_X1 U5819 ( .A1(n5325), .A2(n5324), .ZN(n7276) );
  AND4_X1 U5820 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n9029)
         );
  INV_X1 U5821 ( .A(n9063), .ZN(n9088) );
  INV_X1 U5822 ( .A(n4538), .ZN(n8836) );
  AND2_X1 U5823 ( .A1(n5821), .A2(n6156), .ZN(n8812) );
  AND2_X1 U5824 ( .A1(n5813), .A2(n9506), .ZN(n8859) );
  NAND2_X1 U5825 ( .A1(n8780), .A2(n5796), .ZN(n8848) );
  AND3_X1 U5826 ( .A1(n5822), .A2(n5864), .A3(n9546), .ZN(n8849) );
  AND2_X1 U5827 ( .A1(n5492), .A2(n5481), .ZN(n8942) );
  AND4_X1 U5828 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n9103)
         );
  INV_X1 U5829 ( .A(n8839), .ZN(n8868) );
  INV_X1 U5830 ( .A(n8849), .ZN(n8872) );
  NOR2_X1 U5831 ( .A1(n5733), .A2(n5732), .ZN(n8860) );
  NAND2_X1 U5832 ( .A1(n5354), .A2(n5353), .ZN(n9196) );
  INV_X1 U5833 ( .A(n8859), .ZN(n8870) );
  OAI21_X1 U5834 ( .B1(n4429), .B2(n7831), .A(n4870), .ZN(n4869) );
  NAND2_X1 U5835 ( .A1(n7833), .A2(n7832), .ZN(n4870) );
  XNOR2_X1 U5836 ( .A(n5508), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U5837 ( .A1(n5507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5508) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10146) );
  INV_X1 U5839 ( .A(n6801), .ZN(n8882) );
  INV_X1 U5840 ( .A(n6904), .ZN(n8883) );
  XNOR2_X1 U5841 ( .A(n4558), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U5842 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4558) );
  INV_X1 U5843 ( .A(n4564), .ZN(n9448) );
  XNOR2_X1 U5844 ( .A(n6920), .B(n9469), .ZN(n9472) );
  NOR2_X1 U5845 ( .A1(n7157), .A2(n7158), .ZN(n7161) );
  INV_X1 U5846 ( .A(n4557), .ZN(n7530) );
  NOR2_X1 U5847 ( .A1(n8890), .A2(n8889), .ZN(n8888) );
  AND2_X1 U5848 ( .A1(n4557), .A2(n4556), .ZN(n8890) );
  NAND2_X1 U5849 ( .A1(n7538), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5850 ( .A1(n4741), .A2(n4740), .ZN(n8906) );
  AOI21_X1 U5851 ( .B1(n4412), .B2(n8932), .A(n4408), .ZN(n4740) );
  NAND2_X1 U5852 ( .A1(n4827), .A2(n7789), .ZN(n8933) );
  NAND2_X1 U5853 ( .A1(n4822), .A2(n4820), .ZN(n4827) );
  NAND2_X1 U5854 ( .A1(n4822), .A2(n7779), .ZN(n8945) );
  AND2_X1 U5855 ( .A1(n5479), .A2(n5478), .ZN(n8944) );
  OAI21_X1 U5856 ( .B1(n8993), .B2(n4760), .A(n4759), .ZN(n8952) );
  NAND2_X1 U5857 ( .A1(n5458), .A2(n5457), .ZN(n9150) );
  NAND2_X1 U5858 ( .A1(n4762), .A2(n4763), .ZN(n8964) );
  NAND2_X1 U5859 ( .A1(n8993), .A2(n4764), .ZN(n4762) );
  OAI21_X1 U5860 ( .B1(n8993), .B2(n4399), .A(n5591), .ZN(n8978) );
  OAI21_X1 U5861 ( .B1(n9043), .B2(n4796), .A(n4793), .ZN(n9013) );
  AND2_X1 U5862 ( .A1(n5416), .A2(n5415), .ZN(n9028) );
  INV_X1 U5863 ( .A(n9196), .ZN(n9111) );
  NAND2_X1 U5864 ( .A1(n4745), .A2(n4750), .ZN(n7291) );
  NAND2_X1 U5865 ( .A1(n7208), .A2(n4751), .ZN(n4745) );
  AOI21_X1 U5866 ( .B1(n7208), .B2(n7207), .A(n4397), .ZN(n7265) );
  OAI21_X1 U5867 ( .B1(n4731), .B2(n4732), .A(n4737), .ZN(n9248) );
  NAND2_X1 U5868 ( .A1(n6695), .A2(n4739), .ZN(n4732) );
  NAND2_X1 U5869 ( .A1(n9081), .A2(n9504), .ZN(n9110) );
  NAND2_X1 U5870 ( .A1(n6709), .A2(n5567), .ZN(n6532) );
  NAND2_X1 U5871 ( .A1(n6454), .A2(n4722), .ZN(n6456) );
  INV_X1 U5872 ( .A(n9110), .ZN(n9262) );
  AND2_X2 U5873 ( .A1(n6464), .A2(n6463), .ZN(n9565) );
  OAI21_X1 U5874 ( .B1(n9116), .B2(n9546), .A(n9338), .ZN(n9117) );
  AOI211_X1 U5875 ( .C1(n9529), .C2(n9342), .A(n9341), .B(n9340), .ZN(n9362)
         );
  INV_X1 U5876 ( .A(n9556), .ZN(n9554) );
  AND2_X1 U5877 ( .A1(n5610), .A2(n5541), .ZN(n7835) );
  NAND2_X1 U5878 ( .A1(n7835), .A2(n6342), .ZN(n9515) );
  OR2_X1 U5879 ( .A1(n5134), .A2(n9218), .ZN(n5133) );
  XNOR2_X1 U5880 ( .A(n7467), .B(n7466), .ZN(n8102) );
  XNOR2_X1 U5881 ( .A(n5488), .B(n5489), .ZN(n7440) );
  INV_X1 U5882 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6988) );
  INV_X1 U5883 ( .A(n5544), .ZN(n6989) );
  INV_X1 U5884 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6813) );
  XNOR2_X1 U5885 ( .A(n5446), .B(n5445), .ZN(n7333) );
  INV_X1 U5886 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6673) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6547) );
  INV_X1 U5888 ( .A(n5599), .ZN(n7825) );
  INV_X1 U5889 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U5890 ( .A1(n5510), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5512) );
  INV_X1 U5891 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7546) );
  INV_X1 U5892 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5972) );
  INV_X1 U5893 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9934) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10120) );
  INV_X1 U5895 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5943) );
  INV_X1 U5896 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5917) );
  INV_X1 U5897 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5898) );
  XNOR2_X1 U5898 ( .A(n5262), .B(n4411), .ZN(n6502) );
  INV_X1 U5899 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5889) );
  INV_X1 U5900 ( .A(n5242), .ZN(n4773) );
  AOI21_X1 U5901 ( .B1(n5214), .B2(n5215), .A(n4406), .ZN(n4774) );
  AND2_X1 U5902 ( .A1(n4953), .A2(n4952), .ZN(n5239) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5888) );
  NOR2_X1 U5904 ( .A1(n5198), .A2(n4954), .ZN(n5211) );
  NOR2_X1 U5905 ( .A1(n9305), .A2(n10157), .ZN(n9832) );
  AOI21_X1 U5906 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9830), .ZN(n9829) );
  NOR2_X1 U5907 ( .A1(n9829), .A2(n9828), .ZN(n9827) );
  AOI21_X1 U5908 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9827), .ZN(n9826) );
  NAND2_X1 U5909 ( .A1(n4698), .A2(n8178), .ZN(n4697) );
  INV_X1 U5910 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U5911 ( .A1(n8280), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5912 ( .A1(n4613), .A2(n4606), .ZN(P2_U3264) );
  NAND2_X1 U5913 ( .A1(n8396), .A2(n6749), .ZN(n4613) );
  AOI21_X1 U5914 ( .B1(n4610), .B2(n6138), .A(n4607), .ZN(n4606) );
  AOI211_X1 U5915 ( .C1(n8630), .C2(n9668), .A(n7510), .B(n7509), .ZN(n7511)
         );
  OAI211_X1 U5916 ( .C1(n7543), .C2(n5403), .A(n4568), .B(n4565), .ZN(P1_U3260) );
  NOR2_X1 U5917 ( .A1(n4569), .A2(n4478), .ZN(n4568) );
  NAND2_X1 U5918 ( .A1(n4566), .A2(n5403), .ZN(n4565) );
  INV_X1 U5919 ( .A(n5564), .ZN(n5608) );
  AND2_X1 U5920 ( .A1(n5606), .A2(n4971), .ZN(n5607) );
  INV_X1 U5921 ( .A(n7758), .ZN(n4506) );
  INV_X1 U5922 ( .A(n5543), .ZN(n5403) );
  AND2_X1 U5923 ( .A1(n7215), .A2(n8880), .ZN(n4397) );
  NAND2_X1 U5924 ( .A1(n5100), .A2(n4953), .ZN(n5200) );
  AND2_X1 U5925 ( .A1(n4937), .A2(n4935), .ZN(n4398) );
  NOR2_X1 U5926 ( .A1(n8997), .A2(n8984), .ZN(n4399) );
  NOR2_X1 U5927 ( .A1(n7583), .A2(n8878), .ZN(n4400) );
  INV_X1 U5928 ( .A(n6749), .ZN(n6138) );
  INV_X1 U5929 ( .A(n8497), .ZN(n4642) );
  AND2_X1 U5930 ( .A1(n4786), .A2(n7630), .ZN(n4401) );
  OR2_X1 U5931 ( .A1(n6426), .A2(n6500), .ZN(n4402) );
  AND2_X1 U5932 ( .A1(n8589), .A2(n4932), .ZN(n4403) );
  AND2_X1 U5933 ( .A1(n6902), .A2(n4504), .ZN(n4404) );
  AND2_X1 U5934 ( .A1(n4868), .A2(n5457), .ZN(n4405) );
  NAND2_X1 U5935 ( .A1(n5406), .A2(n5405), .ZN(n9176) );
  INV_X1 U5936 ( .A(n4765), .ZN(n4764) );
  NAND2_X1 U5937 ( .A1(n4424), .A2(n5591), .ZN(n4765) );
  NAND2_X1 U5938 ( .A1(n7779), .A2(n7717), .ZN(n8957) );
  NOR2_X1 U5939 ( .A1(n7073), .A2(n8269), .ZN(n4407) );
  AND2_X1 U5940 ( .A1(n9130), .A2(n8934), .ZN(n4408) );
  NOR2_X1 U5941 ( .A1(n8112), .A2(n8111), .ZN(n4409) );
  INV_X1 U5942 ( .A(n9130), .ZN(n8903) );
  NAND2_X1 U5943 ( .A1(n5114), .A2(n5113), .ZN(n9130) );
  AND2_X1 U5944 ( .A1(n9176), .A2(n5748), .ZN(n7693) );
  INV_X1 U5945 ( .A(n7693), .ZN(n4801) );
  NAND2_X1 U5946 ( .A1(n5491), .A2(n5490), .ZN(n9134) );
  INV_X1 U5947 ( .A(n9134), .ZN(n4743) );
  AND2_X1 U5948 ( .A1(n7317), .A2(n4417), .ZN(n4690) );
  INV_X1 U5949 ( .A(n6191), .ZN(n6193) );
  INV_X1 U5950 ( .A(n7555), .ZN(n5868) );
  OR2_X1 U5951 ( .A1(n5310), .A2(n4842), .ZN(n4410) );
  NOR2_X1 U5952 ( .A1(n5135), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U5953 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n5613)
         );
  AND2_X1 U5954 ( .A1(n5007), .A2(n5006), .ZN(n4411) );
  AND2_X1 U5955 ( .A1(n5595), .A2(n4742), .ZN(n4412) );
  NAND4_X1 U5956 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n5619)
         );
  NAND2_X1 U5957 ( .A1(n5834), .A2(n5833), .ZN(n5895) );
  AND2_X1 U5958 ( .A1(n4891), .A2(n4889), .ZN(n4413) );
  NAND4_X1 U5959 ( .A1(n4952), .A2(n4969), .A3(n4953), .A4(n4771), .ZN(n5322)
         );
  OR2_X1 U5960 ( .A1(n6652), .A2(n6651), .ZN(n4414) );
  INV_X1 U5961 ( .A(n5615), .ZN(n5777) );
  AND2_X1 U5962 ( .A1(n7667), .A2(n7579), .ZN(n4415) );
  AND2_X1 U5963 ( .A1(n4704), .A2(n8185), .ZN(n4416) );
  OR2_X1 U5964 ( .A1(n7364), .A2(n8599), .ZN(n7975) );
  XNOR2_X1 U5965 ( .A(n5940), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U5966 ( .A1(n7314), .A2(n7313), .ZN(n4417) );
  INV_X1 U5967 ( .A(n4783), .ZN(n4782) );
  NAND2_X1 U5968 ( .A1(n4401), .A2(n7634), .ZN(n4783) );
  NAND2_X1 U5969 ( .A1(n4936), .A2(n4937), .ZN(n8773) );
  OR2_X1 U5970 ( .A1(n8028), .A2(n8046), .ZN(n4418) );
  INV_X1 U5971 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5880) );
  INV_X1 U5972 ( .A(n8063), .ZN(n6835) );
  INV_X1 U5973 ( .A(n7789), .ZN(n4826) );
  OR2_X1 U5974 ( .A1(n8940), .A2(n4581), .ZN(n4419) );
  NAND2_X1 U5975 ( .A1(n5365), .A2(n5364), .ZN(n9191) );
  NAND2_X1 U5976 ( .A1(n7344), .A2(n7343), .ZN(n8675) );
  INV_X1 U5977 ( .A(n7794), .ZN(n4798) );
  NOR2_X1 U5978 ( .A1(n8040), .A2(n8039), .ZN(n8037) );
  AND2_X1 U5979 ( .A1(n4770), .A2(n4953), .ZN(n5275) );
  OR2_X1 U5980 ( .A1(n7276), .A2(n8879), .ZN(n4420) );
  OR2_X1 U5981 ( .A1(n8174), .A2(n8177), .ZN(n4421) );
  AND2_X1 U5982 ( .A1(n5833), .A2(n4923), .ZN(n4422) );
  AND2_X1 U5983 ( .A1(n4599), .A2(n4598), .ZN(n4423) );
  OR2_X1 U5984 ( .A1(n9144), .A2(n8853), .ZN(n7779) );
  INV_X1 U5985 ( .A(n7779), .ZN(n4821) );
  NAND2_X1 U5986 ( .A1(n5536), .A2(n5558), .ZN(n5610) );
  AOI21_X1 U5987 ( .B1(n7513), .B2(n7907), .A(n7473), .ZN(n7485) );
  OR2_X1 U5988 ( .A1(n9156), .A2(n9000), .ZN(n4424) );
  NAND2_X1 U5989 ( .A1(n6414), .A2(n6415), .ZN(n4425) );
  XNOR2_X1 U5990 ( .A(n7816), .B(n8910), .ZN(n4426) );
  NAND2_X1 U5991 ( .A1(n4498), .A2(n4495), .ZN(n5534) );
  AND2_X1 U5992 ( .A1(n7144), .A2(n9274), .ZN(n4427) );
  INV_X1 U5993 ( .A(n7151), .ZN(n7249) );
  NAND2_X1 U5994 ( .A1(n5308), .A2(n5307), .ZN(n7151) );
  NAND2_X1 U5995 ( .A1(n7429), .A2(n7428), .ZN(n8645) );
  NOR2_X1 U5996 ( .A1(n4684), .A2(n8209), .ZN(n4683) );
  NAND2_X1 U5997 ( .A1(n8466), .A2(n4619), .ZN(n4620) );
  NAND2_X1 U5998 ( .A1(n8556), .A2(n4625), .ZN(n4628) );
  INV_X1 U5999 ( .A(n4953), .ZN(n5198) );
  AND2_X1 U6000 ( .A1(n5099), .A2(n5169), .ZN(n4953) );
  OR2_X1 U6001 ( .A1(n8568), .A2(n8593), .ZN(n4428) );
  OR2_X1 U6002 ( .A1(n7833), .A2(n5543), .ZN(n4429) );
  NAND3_X1 U6003 ( .A1(n5505), .A2(n5504), .A3(n5503), .ZN(n4430) );
  NAND2_X1 U6004 ( .A1(n4514), .A2(n4513), .ZN(n5018) );
  OR2_X1 U6005 ( .A1(n9134), .A2(n8854), .ZN(n7781) );
  INV_X1 U6006 ( .A(n7781), .ZN(n4815) );
  OR2_X1 U6007 ( .A1(n6936), .A2(n5682), .ZN(n4431) );
  INV_X1 U6008 ( .A(n4915), .ZN(n4914) );
  NAND2_X1 U6009 ( .A1(n8499), .A2(n8013), .ZN(n4432) );
  AND2_X1 U6010 ( .A1(n4416), .A2(n4702), .ZN(n4433) );
  AND2_X1 U6011 ( .A1(n7455), .A2(n7454), .ZN(n8415) );
  NAND2_X1 U6012 ( .A1(n8124), .A2(n8125), .ZN(n4434) );
  AND2_X1 U6013 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4435) );
  NOR2_X1 U6014 ( .A1(n5738), .A2(n5737), .ZN(n4436) );
  INV_X1 U6015 ( .A(n5576), .ZN(n4739) );
  OR2_X1 U6016 ( .A1(n4645), .A2(n4644), .ZN(n4437) );
  NAND2_X1 U6017 ( .A1(n5362), .A2(n4963), .ZN(n4438) );
  NOR2_X1 U6018 ( .A1(n9150), .A2(n4868), .ZN(n4439) );
  NOR2_X1 U6019 ( .A1(n5763), .A2(n5762), .ZN(n4440) );
  AND2_X1 U6020 ( .A1(n4917), .A2(n7027), .ZN(n4441) );
  INV_X1 U6021 ( .A(n4572), .ZN(n4571) );
  NAND2_X1 U6022 ( .A1(n4574), .A2(n4573), .ZN(n4572) );
  AND2_X1 U6023 ( .A1(n8007), .A2(n8000), .ZN(n4442) );
  AND3_X1 U6024 ( .A1(n5464), .A2(n5463), .A3(n5462), .ZN(n8738) );
  INV_X1 U6025 ( .A(n8738), .ZN(n4868) );
  NOR2_X1 U6026 ( .A1(n8122), .A2(n8121), .ZN(n4443) );
  NOR2_X1 U6027 ( .A1(n8653), .A2(n8501), .ZN(n4444) );
  INV_X1 U6028 ( .A(n8997), .ZN(n9159) );
  AND2_X1 U6029 ( .A1(n5438), .A2(n5437), .ZN(n8997) );
  INV_X1 U6030 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6031 ( .A1(n4957), .A2(n5716), .ZN(n4445) );
  AND2_X1 U6032 ( .A1(n8415), .A2(n7465), .ZN(n4446) );
  OR2_X1 U6033 ( .A1(n5534), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4447) );
  AND2_X1 U6034 ( .A1(n5003), .A2(SI_7_), .ZN(n4448) );
  OR2_X1 U6035 ( .A1(n4716), .A2(n4708), .ZN(n4449) );
  INV_X1 U6036 ( .A(n4677), .ZN(n4676) );
  NOR2_X1 U6037 ( .A1(n8119), .A2(n8224), .ZN(n4677) );
  INV_X1 U6038 ( .A(n5016), .ZN(n5289) );
  NAND2_X1 U6039 ( .A1(n7635), .A2(n7585), .ZN(n4450) );
  INV_X1 U6040 ( .A(n4864), .ZN(n4863) );
  INV_X1 U6041 ( .A(n4690), .ZN(n4689) );
  NOR2_X1 U6042 ( .A1(n8990), .A2(n10145), .ZN(n4451) );
  NOR2_X1 U6043 ( .A1(n9350), .A2(n7126), .ZN(n4754) );
  INV_X1 U6044 ( .A(n4713), .ZN(n4712) );
  INV_X1 U6045 ( .A(n4761), .ZN(n4760) );
  AND2_X1 U6046 ( .A1(n4454), .A2(n4763), .ZN(n4761) );
  INV_X1 U6047 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5112) );
  AND2_X1 U6048 ( .A1(n5530), .A2(n5110), .ZN(n4452) );
  AND2_X1 U6049 ( .A1(n5810), .A2(n8782), .ZN(n4453) );
  OR2_X1 U6050 ( .A1(n5779), .A2(n8738), .ZN(n4454) );
  OR2_X1 U6051 ( .A1(n7775), .A2(n7746), .ZN(n4455) );
  INV_X1 U6052 ( .A(n6759), .ZN(n4787) );
  AND2_X1 U6053 ( .A1(n4617), .A2(n7485), .ZN(n4456) );
  AND2_X1 U6054 ( .A1(n4964), .A2(n5511), .ZN(n4457) );
  AND2_X1 U6055 ( .A1(n5906), .A2(n5905), .ZN(n4458) );
  AND2_X1 U6056 ( .A1(n6834), .A2(n7891), .ZN(n4459) );
  AND2_X1 U6057 ( .A1(n8033), .A2(n4418), .ZN(n4460) );
  OR2_X1 U6058 ( .A1(n5168), .A2(n6165), .ZN(n4461) );
  NOR2_X1 U6059 ( .A1(n4858), .A2(n5398), .ZN(n4857) );
  INV_X1 U6060 ( .A(n5567), .ZN(n4728) );
  AND2_X1 U6061 ( .A1(n4700), .A2(n4416), .ZN(n4462) );
  AND2_X1 U6062 ( .A1(n5927), .A2(n5932), .ZN(n4463) );
  INV_X1 U6063 ( .A(n4929), .ZN(n4928) );
  NOR2_X1 U6064 ( .A1(n7378), .A2(n4930), .ZN(n4929) );
  AND2_X1 U6065 ( .A1(n5839), .A2(n4680), .ZN(n4464) );
  AND2_X1 U6066 ( .A1(n4670), .A2(n4434), .ZN(n4465) );
  OAI21_X1 U6067 ( .B1(n4640), .B2(n4641), .A(n4642), .ZN(n4639) );
  INV_X1 U6068 ( .A(n6991), .ZN(n8067) );
  AND2_X1 U6069 ( .A1(n7951), .A2(n7952), .ZN(n6991) );
  INV_X1 U6070 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5932) );
  INV_X1 U6071 ( .A(n6654), .ZN(n4720) );
  NAND2_X1 U6072 ( .A1(n5390), .A2(n5389), .ZN(n9179) );
  INV_X1 U6073 ( .A(n9179), .ZN(n4573) );
  OAI21_X1 U6074 ( .B1(n6502), .B2(n5229), .A(n4553), .ZN(n7018) );
  INV_X1 U6075 ( .A(n8878), .ZN(n9102) );
  NAND2_X1 U6076 ( .A1(n6077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6402) );
  AND2_X1 U6077 ( .A1(n5733), .A2(n5732), .ZN(n4466) );
  NAND2_X1 U6078 ( .A1(n4958), .A2(n5716), .ZN(n7120) );
  NAND2_X1 U6079 ( .A1(n4931), .A2(n4403), .ZN(n8579) );
  NAND2_X1 U6080 ( .A1(n5834), .A2(n4922), .ZN(n5918) );
  NAND2_X1 U6081 ( .A1(n5339), .A2(n5338), .ZN(n7583) );
  INV_X1 U6082 ( .A(n8904), .ZN(n8934) );
  INV_X1 U6083 ( .A(n8251), .ZN(n8143) );
  OR2_X1 U6084 ( .A1(n8546), .A2(n8555), .ZN(n4467) );
  NOR3_X1 U6085 ( .A1(n9008), .A2(n9144), .A3(n4586), .ZN(n4584) );
  NAND2_X1 U6086 ( .A1(n9105), .A2(n4571), .ZN(n4575) );
  INV_X1 U6087 ( .A(n8854), .ZN(n8947) );
  AND2_X1 U6088 ( .A1(n5502), .A2(n5501), .ZN(n8854) );
  AND2_X1 U6089 ( .A1(n8189), .A2(n8190), .ZN(n4468) );
  INV_X1 U6090 ( .A(n8178), .ZN(n4702) );
  INV_X1 U6091 ( .A(n4585), .ZN(n8971) );
  NOR2_X1 U6092 ( .A1(n9008), .A2(n4586), .ZN(n4585) );
  INV_X1 U6093 ( .A(n4850), .ZN(n4849) );
  NOR2_X1 U6094 ( .A1(n5435), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U6095 ( .A1(n5280), .A2(n5279), .ZN(n6949) );
  INV_X1 U6096 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5511) );
  OR2_X1 U6097 ( .A1(n9144), .A2(n8969), .ZN(n4469) );
  AND2_X1 U6098 ( .A1(n6503), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4470) );
  AND2_X1 U6099 ( .A1(n5054), .A2(SI_18_), .ZN(n4471) );
  AND2_X1 U6100 ( .A1(n7120), .A2(n5717), .ZN(n4472) );
  NAND2_X1 U6101 ( .A1(n7335), .A2(n7334), .ZN(n8658) );
  AND2_X1 U6102 ( .A1(n4877), .A2(n4876), .ZN(n4473) );
  AND2_X1 U6103 ( .A1(n4691), .A2(n4417), .ZN(n4474) );
  INV_X1 U6104 ( .A(n7809), .ZN(n4810) );
  XNOR2_X1 U6105 ( .A(n5509), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5599) );
  INV_X1 U6106 ( .A(n5193), .ZN(n5296) );
  AND2_X1 U6107 ( .A1(n6570), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U6108 ( .A1(n4906), .A2(n6832), .ZN(n7882) );
  NAND2_X1 U6109 ( .A1(n7363), .A2(n7362), .ZN(n8692) );
  INV_X1 U6110 ( .A(n8692), .ZN(n4615) );
  OR2_X1 U6111 ( .A1(n5757), .A2(n5756), .ZN(n4476) );
  NOR2_X1 U6112 ( .A1(n4499), .A2(n5322), .ZN(n5537) );
  INV_X1 U6113 ( .A(n6653), .ZN(n4719) );
  AND2_X1 U6114 ( .A1(n6885), .A2(n7947), .ZN(n4477) );
  NAND2_X1 U6115 ( .A1(n4724), .A2(n6455), .ZN(n6454) );
  NAND2_X1 U6116 ( .A1(n7921), .A2(n7924), .ZN(n9675) );
  INV_X1 U6117 ( .A(n9675), .ZN(n4888) );
  AND2_X1 U6118 ( .A1(n5630), .A2(n6331), .ZN(n7862) );
  INV_X1 U6119 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n4560) );
  INV_X1 U6120 ( .A(n6925), .ZN(n4561) );
  AND2_X1 U6121 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n4478) );
  NAND2_X1 U6122 ( .A1(n6085), .A2(n6084), .ZN(n6749) );
  XNOR2_X1 U6123 ( .A(n5133), .B(n5132), .ZN(n8106) );
  AND2_X2 U6124 ( .A1(n4539), .A2(n4538), .ZN(n8745) );
  NAND2_X1 U6125 ( .A1(n4537), .A2(n4934), .ZN(n5765) );
  NOR2_X2 U6126 ( .A1(n8824), .A2(n8826), .ZN(n5776) );
  NAND2_X1 U6127 ( .A1(n4961), .A2(n4959), .ZN(n8762) );
  NAND2_X1 U6128 ( .A1(n5691), .A2(n5690), .ZN(n6642) );
  NAND2_X1 U6129 ( .A1(n4867), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4866) );
  OAI21_X1 U6130 ( .B1(n8027), .B2(n8029), .A(n4656), .ZN(n4655) );
  AOI21_X1 U6131 ( .B1(n7940), .B2(n4636), .A(n4635), .ZN(n4634) );
  OAI21_X1 U6132 ( .B1(n4650), .B2(n8089), .A(n8088), .ZN(n4649) );
  OAI21_X1 U6133 ( .B1(n8051), .B2(n8050), .A(n8049), .ZN(n8090) );
  OAI211_X1 U6134 ( .C1(n8023), .C2(n8022), .A(n8030), .B(n8021), .ZN(n8031)
         );
  AOI21_X1 U6135 ( .B1(n7978), .B2(n7977), .A(n8600), .ZN(n7983) );
  NOR2_X1 U6136 ( .A1(n7989), .A2(n7988), .ZN(n7995) );
  INV_X2 U6137 ( .A(n7555), .ZN(n4895) );
  AOI21_X2 U6138 ( .B1(n8520), .B2(n7390), .A(n4482), .ZN(n8506) );
  NAND2_X2 U6139 ( .A1(n8673), .A2(n4467), .ZN(n8520) );
  XNOR2_X1 U6140 ( .A(n7481), .B(n8037), .ZN(n8632) );
  NAND2_X2 U6141 ( .A1(n6829), .A2(n4980), .ZN(n6831) );
  NAND2_X1 U6142 ( .A1(n8441), .A2(n8446), .ZN(n8440) );
  NOR2_X2 U6143 ( .A1(n7093), .A2(n4973), .ZN(n7097) );
  AOI21_X1 U6144 ( .B1(n7366), .B2(n8075), .A(n7365), .ZN(n8601) );
  AOI21_X1 U6145 ( .B1(n8243), .B2(n8561), .A(n7379), .ZN(n8540) );
  NAND3_X1 U6146 ( .A1(n4484), .A2(n7999), .A3(n8534), .ZN(n7998) );
  AOI22_X1 U6147 ( .A1(n4649), .A2(n8092), .B1(n8093), .B2(n4530), .ZN(n8101)
         );
  NAND2_X1 U6148 ( .A1(n5173), .A2(n5172), .ZN(n4828) );
  INV_X1 U6149 ( .A(n8090), .ZN(n4650) );
  OAI21_X1 U6150 ( .B1(n4634), .B2(n4633), .A(n7956), .ZN(n7962) );
  AOI21_X1 U6151 ( .B1(n4655), .B2(n4653), .A(n4651), .ZN(n8051) );
  NOR2_X1 U6152 ( .A1(n8002), .A2(n4640), .ZN(n4638) );
  NAND2_X2 U6153 ( .A1(n8440), .A2(n7439), .ZN(n8431) );
  NAND2_X1 U6154 ( .A1(n9699), .A2(n6754), .ZN(n6816) );
  NAND3_X1 U6155 ( .A1(n8061), .A2(n6831), .A3(n4907), .ZN(n4904) );
  NAND3_X1 U6156 ( .A1(n4509), .A2(n4511), .A3(n5227), .ZN(n4487) );
  NAND2_X1 U6157 ( .A1(n6882), .A2(n6881), .ZN(n6990) );
  INV_X1 U6158 ( .A(n6832), .ZN(n4905) );
  NAND2_X1 U6159 ( .A1(n4872), .A2(n4489), .ZN(n4871) );
  NAND2_X1 U6160 ( .A1(n4490), .A2(n4873), .ZN(n4489) );
  NAND2_X1 U6161 ( .A1(n4491), .A2(n7827), .ZN(n4490) );
  NAND2_X1 U6162 ( .A1(n7830), .A2(n7824), .ZN(n4491) );
  AOI21_X1 U6163 ( .B1(n4492), .B2(n7792), .A(n7791), .ZN(n7706) );
  AOI21_X1 U6164 ( .B1(n7698), .B2(n7697), .A(n7696), .ZN(n4493) );
  AOI21_X1 U6165 ( .B1(n7698), .B2(n7695), .A(n7694), .ZN(n4494) );
  INV_X1 U6166 ( .A(n5109), .ZN(n4499) );
  NAND2_X1 U6167 ( .A1(n6726), .A2(n4404), .ZN(n4501) );
  NAND2_X1 U6168 ( .A1(n4501), .A2(n4502), .ZN(n6903) );
  NAND2_X1 U6169 ( .A1(n4503), .A2(n7758), .ZN(n6555) );
  NAND2_X1 U6170 ( .A1(n4996), .A2(n4510), .ZN(n4509) );
  INV_X1 U6171 ( .A(n5203), .ZN(n4510) );
  NAND3_X1 U6172 ( .A1(n4996), .A2(n4993), .A3(n4992), .ZN(n4511) );
  NAND2_X1 U6173 ( .A1(n4512), .A2(n4996), .ZN(n5228) );
  NAND2_X1 U6174 ( .A1(n5202), .A2(n5203), .ZN(n4512) );
  NAND2_X1 U6175 ( .A1(n5262), .A2(n4515), .ZN(n4514) );
  OAI21_X1 U6176 ( .B1(n5262), .B2(n4520), .A(n5007), .ZN(n5274) );
  NAND2_X1 U6177 ( .A1(n4521), .A2(n4986), .ZN(n5173) );
  MUX2_X1 U6178 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n7555), .Z(n5158) );
  MUX2_X1 U6179 ( .A(n5871), .B(n6105), .S(n7555), .Z(n4987) );
  AND2_X2 U6180 ( .A1(n4535), .A2(n4534), .ZN(n5733) );
  OR2_X1 U6181 ( .A1(n8732), .A2(n4544), .ZN(n4541) );
  AND2_X1 U6182 ( .A1(n8734), .A2(n4548), .ZN(n4547) );
  NAND2_X2 U6183 ( .A1(n4546), .A2(n4547), .ZN(n8806) );
  NAND3_X1 U6184 ( .A1(n6675), .A2(n6935), .A3(n5683), .ZN(n5685) );
  NAND2_X1 U6185 ( .A1(n4550), .A2(n4549), .ZN(n5683) );
  MUX2_X1 U6186 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5993), .S(n9386), .Z(n9388)
         );
  NOR2_X2 U6187 ( .A1(n4954), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4952) );
  INV_X1 U6188 ( .A(n4575), .ZN(n9056) );
  NAND3_X1 U6189 ( .A1(n4577), .A2(n4578), .A3(n9547), .ZN(n9264) );
  OR3_X1 U6190 ( .A1(n8940), .A2(n9134), .A3(n9130), .ZN(n8918) );
  NOR2_X1 U6191 ( .A1(n8940), .A2(n9134), .ZN(n8928) );
  INV_X1 U6192 ( .A(n4584), .ZN(n8953) );
  NAND2_X1 U6193 ( .A1(n4614), .A2(n6079), .ZN(n5844) );
  OAI21_X1 U6194 ( .B1(n8722), .B2(n6078), .A(n4614), .ZN(n4664) );
  OR2_X1 U6195 ( .A1(n6083), .A2(n4614), .ZN(n6085) );
  NAND2_X1 U6196 ( .A1(n8466), .A2(n8455), .ZN(n8449) );
  INV_X1 U6197 ( .A(n4620), .ZN(n8432) );
  INV_X1 U6198 ( .A(n8415), .ZN(n4621) );
  NAND2_X1 U6199 ( .A1(n8556), .A2(n4624), .ZN(n8490) );
  INV_X1 U6200 ( .A(n4628), .ZN(n8507) );
  NAND3_X1 U6201 ( .A1(n4924), .A2(n5906), .A3(n4629), .ZN(n5930) );
  INV_X1 U6202 ( .A(n9699), .ZN(n4631) );
  OAI21_X1 U6203 ( .B1(n6754), .B2(n8280), .A(n4632), .ZN(P2_U3553) );
  AND4_X2 U6204 ( .A1(n6074), .A2(n6075), .A3(n6072), .A4(n6073), .ZN(n6754)
         );
  NOR2_X1 U6205 ( .A1(n4638), .A2(n4639), .ZN(n8010) );
  INV_X1 U6206 ( .A(n7999), .ZN(n4644) );
  INV_X1 U6207 ( .A(n8003), .ZN(n4645) );
  NAND2_X1 U6208 ( .A1(n6773), .A2(n6772), .ZN(n8060) );
  NAND3_X2 U6209 ( .A1(n5834), .A2(n5836), .A3(n4922), .ZN(n5904) );
  OR2_X1 U6210 ( .A1(n6402), .A2(n8722), .ZN(n4659) );
  NAND2_X1 U6211 ( .A1(n6402), .A2(n4663), .ZN(n4661) );
  NAND2_X1 U6212 ( .A1(n6402), .A2(n6078), .ZN(n4662) );
  AND2_X2 U6213 ( .A1(n4672), .A2(n4465), .ZN(n8128) );
  NAND2_X1 U6214 ( .A1(n8144), .A2(n4462), .ZN(n4696) );
  OAI211_X1 U6215 ( .C1(n8144), .C2(n4697), .A(n4696), .B(n4692), .ZN(P2_U3222) );
  NAND2_X1 U6216 ( .A1(n8144), .A2(n8143), .ZN(n8253) );
  OAI21_X2 U6217 ( .B1(n6654), .B2(n4449), .A(n4707), .ZN(n7231) );
  NAND3_X1 U6218 ( .A1(n6964), .A2(n4721), .A3(n4714), .ZN(n4713) );
  INV_X1 U6219 ( .A(n4721), .ZN(n4717) );
  NAND2_X1 U6220 ( .A1(n6959), .A2(n6960), .ZN(n4721) );
  NAND4_X1 U6221 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n4724), .ZN(n7804)
         );
  NAND2_X1 U6222 ( .A1(n6711), .A2(n5567), .ZN(n4727) );
  NAND2_X1 U6223 ( .A1(n4727), .A2(n4725), .ZN(n6531) );
  INV_X1 U6224 ( .A(n5575), .ZN(n4731) );
  NAND2_X1 U6225 ( .A1(n6695), .A2(n4735), .ZN(n4734) );
  AOI21_X1 U6226 ( .B1(n5575), .B2(n6695), .A(n5574), .ZN(n6758) );
  NOR2_X1 U6227 ( .A1(n9253), .A2(n6949), .ZN(n4738) );
  NAND2_X1 U6228 ( .A1(n8927), .A2(n4412), .ZN(n4741) );
  OR2_X1 U6229 ( .A1(n8927), .A2(n8932), .ZN(n4744) );
  NAND3_X1 U6230 ( .A1(n4953), .A2(n4952), .A3(n5240), .ZN(n5260) );
  NAND2_X1 U6231 ( .A1(n4775), .A2(n4777), .ZN(n5309) );
  NAND2_X1 U6232 ( .A1(n6699), .A2(n4779), .ZN(n4775) );
  NAND3_X1 U6233 ( .A1(n4787), .A2(n7627), .A3(n5264), .ZN(n4786) );
  NAND2_X1 U6234 ( .A1(n9043), .A2(n4793), .ZN(n4792) );
  NAND3_X1 U6235 ( .A1(n4803), .A2(n4802), .A3(n4983), .ZN(n5151) );
  NAND2_X1 U6236 ( .A1(n7209), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U6237 ( .A1(n8966), .A2(n4816), .ZN(n4813) );
  NAND2_X1 U6238 ( .A1(n4813), .A2(n4814), .ZN(n8910) );
  NAND2_X1 U6239 ( .A1(n8966), .A2(n4823), .ZN(n4822) );
  NAND2_X1 U6240 ( .A1(n8966), .A2(n7709), .ZN(n8958) );
  INV_X1 U6241 ( .A(n7709), .ZN(n4824) );
  NAND2_X1 U6242 ( .A1(n4828), .A2(n4989), .ZN(n5186) );
  NAND2_X1 U6243 ( .A1(n5214), .A2(n4835), .ZN(n4833) );
  NAND2_X1 U6244 ( .A1(n5018), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U6245 ( .A1(n5374), .A2(n4857), .ZN(n4854) );
  OAI21_X1 U6246 ( .B1(n5374), .B2(n5053), .A(n5052), .ZN(n5385) );
  AOI21_X1 U6247 ( .B1(n5053), .B2(n5052), .A(n5386), .ZN(n4864) );
  AOI21_X1 U6248 ( .B1(n4871), .B2(n7831), .A(n4869), .ZN(n7841) );
  OR2_X1 U6249 ( .A1(n7830), .A2(n7829), .ZN(n4872) );
  NAND2_X1 U6250 ( .A1(n8496), .A2(n7503), .ZN(n8499) );
  NAND2_X1 U6251 ( .A1(n4884), .A2(n7885), .ZN(n7040) );
  NAND2_X1 U6252 ( .A1(n7497), .A2(n4885), .ZN(n8551) );
  NAND2_X1 U6253 ( .A1(n8551), .A2(n7500), .ZN(n7501) );
  INV_X1 U6254 ( .A(n8551), .ZN(n7498) );
  NAND2_X1 U6255 ( .A1(n4887), .A2(n7921), .ZN(n9642) );
  NAND3_X1 U6256 ( .A1(n8060), .A2(n7923), .A3(n4888), .ZN(n4887) );
  AOI21_X1 U6257 ( .B1(n7507), .B2(n8081), .A(n9644), .ZN(n4892) );
  NAND2_X1 U6258 ( .A1(n6423), .A2(n4895), .ZN(n6310) );
  NAND2_X1 U6259 ( .A1(n6423), .A2(n7555), .ZN(n6203) );
  NAND2_X1 U6260 ( .A1(n6423), .A2(n4894), .ZN(n4893) );
  AND2_X2 U6261 ( .A1(n6091), .A2(n4893), .ZN(n9699) );
  OAI21_X1 U6262 ( .B1(n8431), .B2(n4902), .A(n4900), .ZN(n8408) );
  NAND2_X1 U6263 ( .A1(n4899), .A2(n4898), .ZN(n7481) );
  NAND2_X1 U6264 ( .A1(n8431), .A2(n4900), .ZN(n4899) );
  NAND2_X1 U6265 ( .A1(n6831), .A2(n4907), .ZN(n4906) );
  NAND2_X1 U6266 ( .A1(n4904), .A2(n4903), .ZN(n7039) );
  AOI21_X1 U6267 ( .B1(n4905), .B2(n8061), .A(n4459), .ZN(n4903) );
  NAND2_X1 U6268 ( .A1(n8489), .A2(n4911), .ZN(n4910) );
  OAI21_X1 U6269 ( .B1(n8489), .B2(n4912), .A(n4911), .ZN(n8460) );
  NOR2_X1 U6270 ( .A1(n8495), .A2(n7403), .ZN(n4915) );
  INV_X1 U6271 ( .A(n8068), .ZN(n4917) );
  NAND2_X1 U6272 ( .A1(n8603), .A2(n4929), .ZN(n4925) );
  INV_X1 U6273 ( .A(n5754), .ZN(n4942) );
  NAND2_X1 U6274 ( .A1(n8745), .A2(n8746), .ZN(n8744) );
  OAI21_X1 U6275 ( .B1(n5733), .B2(n4947), .A(n4945), .ZN(n8790) );
  NAND3_X1 U6276 ( .A1(n5650), .A2(n4951), .A3(n5646), .ZN(n6522) );
  NAND2_X1 U6277 ( .A1(n8781), .A2(n4453), .ZN(n4961) );
  OR4_X2 U6278 ( .A1(n8762), .A2(n8768), .A3(n8872), .A4(n8767), .ZN(n8772) );
  NAND2_X1 U6279 ( .A1(n5362), .A2(n4964), .ZN(n5510) );
  NAND2_X1 U6280 ( .A1(n5362), .A2(n4457), .ZN(n4962) );
  NAND2_X1 U6281 ( .A1(n5275), .A2(n4967), .ZN(n5337) );
  NAND2_X1 U6282 ( .A1(n9119), .A2(n9118), .ZN(n9201) );
  NAND2_X1 U6283 ( .A1(n9115), .A2(n9530), .ZN(n9119) );
  OAI222_X1 U6284 ( .A1(n4426), .A2(n9256), .B1(n7563), .B2(n9104), .C1(n8854), 
        .C2(n5525), .ZN(n5526) );
  OAI22_X1 U6285 ( .A1(n6814), .A2(n6193), .B1(n6776), .B2(n6102), .ZN(n6355)
         );
  NAND2_X1 U6286 ( .A1(n6093), .A2(n6092), .ZN(n6103) );
  XNOR2_X1 U6287 ( .A(n6102), .B(n9699), .ZN(n6092) );
  NAND2_X1 U6288 ( .A1(n6088), .A2(n6750), .ZN(n6102) );
  INV_X4 U6289 ( .A(n6193), .ZN(n8140) );
  OR2_X1 U6290 ( .A1(n8603), .A2(n8602), .ZN(n8699) );
  NAND2_X1 U6291 ( .A1(n6823), .A2(n6824), .ZN(n6841) );
  NAND2_X1 U6292 ( .A1(n5177), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6293 ( .A1(n7862), .A2(n7864), .ZN(n7863) );
  INV_X1 U6294 ( .A(n6070), .ZN(n7896) );
  INV_X1 U6295 ( .A(n6157), .ZN(n6158) );
  NAND2_X1 U6296 ( .A1(n6522), .A2(n5653), .ZN(n6675) );
  XNOR2_X1 U6297 ( .A(n5656), .B(n8756), .ZN(n6869) );
  NOR2_X1 U6298 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5099) );
  OAI22_X1 U6299 ( .A1(n6905), .A2(n5668), .B1(n6553), .B2(n5788), .ZN(n5656)
         );
  NAND2_X1 U6300 ( .A1(n6145), .A2(n6146), .ZN(n6147) );
  OR2_X1 U6301 ( .A1(n5229), .A2(n6089), .ZN(n5160) );
  INV_X1 U6302 ( .A(n8730), .ZN(n6069) );
  INV_X4 U6303 ( .A(n7477), .ZN(n7488) );
  NAND2_X1 U6304 ( .A1(n5543), .A2(n5598), .ZN(n6602) );
  NAND2_X1 U6305 ( .A1(n5177), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5155) );
  AOI21_X1 U6306 ( .B1(n8417), .B2(n8033), .A(n7506), .ZN(n7507) );
  INV_X1 U6307 ( .A(n7512), .ZN(n5139) );
  INV_X1 U6308 ( .A(n7838), .ZN(n7755) );
  INV_X1 U6309 ( .A(n7093), .ZN(n7077) );
  NAND2_X1 U6310 ( .A1(n8106), .A2(n7512), .ZN(n5499) );
  INV_X1 U6311 ( .A(n8106), .ZN(n5138) );
  AND2_X2 U6312 ( .A1(n6753), .A2(n9666), .ZN(n9669) );
  NAND2_X1 U6313 ( .A1(n6732), .A2(n9506), .ZN(n9081) );
  INV_X1 U6314 ( .A(n9513), .ZN(n5603) );
  AND2_X1 U6315 ( .A1(n5930), .A2(n5929), .ZN(n4970) );
  NAND2_X1 U6316 ( .A1(n7464), .A2(n7463), .ZN(n8426) );
  INV_X1 U6317 ( .A(n8426), .ZN(n7465) );
  NOR2_X1 U6318 ( .A1(n5605), .A2(n5604), .ZN(n4971) );
  OR2_X1 U6319 ( .A1(n7465), .A2(n9611), .ZN(n4972) );
  AND2_X1 U6320 ( .A1(n9325), .A2(n8268), .ZN(n4973) );
  OR2_X1 U6321 ( .A1(n9111), .A2(n9087), .ZN(n4974) );
  OR2_X1 U6322 ( .A1(n9012), .A2(n9029), .ZN(n4975) );
  OR2_X1 U6323 ( .A1(n9122), .A2(n9546), .ZN(n4976) );
  OR2_X1 U6324 ( .A1(n5168), .A2(n5899), .ZN(n4977) );
  AND2_X1 U6325 ( .A1(n4895), .A2(P1_U3084), .ZN(n7259) );
  AND2_X1 U6326 ( .A1(n5333), .A2(n5033), .ZN(n4978) );
  AND2_X1 U6327 ( .A1(n6350), .A2(n5598), .ZN(n9530) );
  INV_X1 U6328 ( .A(n9530), .ZN(n9548) );
  AND2_X1 U6329 ( .A1(n7824), .A2(n7834), .ZN(n9254) );
  AND2_X1 U6330 ( .A1(n8273), .A2(n7941), .ZN(n4979) );
  OR2_X1 U6331 ( .A1(n8276), .A2(n4395), .ZN(n4980) );
  INV_X1 U6332 ( .A(n7583), .ZN(n9345) );
  OR2_X1 U6333 ( .A1(n7151), .A2(n9252), .ZN(n4982) );
  INV_X1 U6334 ( .A(n6096), .ZN(n7448) );
  INV_X1 U6335 ( .A(n7795), .ZN(n5566) );
  INV_X1 U6336 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5103) );
  NOR2_X1 U6337 ( .A1(n8625), .A2(n7508), .ZN(n8043) );
  INV_X1 U6338 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5905) );
  INV_X1 U6339 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5835) );
  INV_X1 U6340 ( .A(n5766), .ZN(n5767) );
  AOI21_X1 U6341 ( .B1(n7826), .B2(n7825), .A(n5543), .ZN(n7827) );
  INV_X1 U6342 ( .A(n7410), .ZN(n7408) );
  INV_X1 U6343 ( .A(n7395), .ZN(n7339) );
  INV_X1 U6344 ( .A(n8446), .ZN(n7505) );
  INV_X1 U6345 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5966) );
  INV_X1 U6346 ( .A(n6936), .ZN(n6937) );
  INV_X1 U6347 ( .A(n5429), .ZN(n5124) );
  INV_X1 U6348 ( .A(n7823), .ZN(n7828) );
  INV_X1 U6349 ( .A(n5340), .ZN(n5120) );
  INV_X1 U6350 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5602) );
  INV_X1 U6351 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6352 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  NAND2_X1 U6353 ( .A1(n7408), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7419) );
  NAND2_X1 U6354 ( .A1(n7339), .A2(n7338), .ZN(n7396) );
  OR2_X1 U6355 ( .A1(n6577), .A2(n6594), .ZN(n6661) );
  NAND2_X1 U6356 ( .A1(n8470), .A2(n8217), .ZN(n7425) );
  INV_X1 U6357 ( .A(n6752), .ZN(n6133) );
  INV_X1 U6358 ( .A(n5407), .ZN(n5123) );
  INV_X1 U6359 ( .A(n6869), .ZN(n6676) );
  INV_X1 U6360 ( .A(n7122), .ZN(n5716) );
  NAND2_X1 U6361 ( .A1(n5120), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5367) );
  NOR2_X1 U6362 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  OR2_X1 U6363 ( .A1(n5266), .A2(n5265), .ZN(n5282) );
  OR2_X1 U6364 ( .A1(n6791), .A2(n6902), .ZN(n6897) );
  INV_X1 U6365 ( .A(n5190), .ZN(n6535) );
  NAND2_X1 U6366 ( .A1(n5044), .A2(n9901), .ZN(n5047) );
  INV_X1 U6367 ( .A(SI_8_), .ZN(n10066) );
  INV_X1 U6368 ( .A(n6423), .ZN(n7369) );
  OAI21_X1 U6369 ( .B1(n8159), .B2(n8131), .A(n8130), .ZN(n8134) );
  OR2_X1 U6370 ( .A1(n7319), .A2(n8358), .ZN(n7373) );
  NAND2_X1 U6371 ( .A1(n6141), .A2(n6140), .ZN(n9586) );
  INV_X1 U6372 ( .A(n8187), .ZN(n8245) );
  OR2_X1 U6373 ( .A1(n7396), .A2(n8160), .ZN(n7410) );
  INV_X1 U6374 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10027) );
  INV_X1 U6375 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6594) );
  INV_X1 U6376 ( .A(n8528), .ZN(n8555) );
  INV_X1 U6377 ( .A(n8264), .ZN(n8593) );
  NOR2_X1 U6378 ( .A1(n7075), .A2(n8070), .ZN(n7093) );
  INV_X1 U6379 ( .A(n8702), .ZN(n6744) );
  AND2_X1 U6380 ( .A1(n8094), .A2(n6133), .ZN(n9751) );
  INV_X1 U6381 ( .A(n8271), .ZN(n6888) );
  XNOR2_X1 U6382 ( .A(n6080), .B(n6079), .ZN(n6087) );
  INV_X1 U6383 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8722) );
  AOI21_X1 U6384 ( .B1(n5805), .B2(n5804), .A(n8767), .ZN(n5806) );
  OR2_X1 U6385 ( .A1(n5449), .A2(n8737), .ZN(n5460) );
  NAND2_X1 U6386 ( .A1(n5123), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6387 ( .A1(n5627), .A2(n5626), .ZN(n6332) );
  INV_X1 U6388 ( .A(n5672), .ZN(n6678) );
  OR2_X1 U6389 ( .A1(n5439), .A2(n8829), .ZN(n5449) );
  OR2_X1 U6390 ( .A1(n5480), .A2(n8851), .ZN(n5492) );
  AND2_X1 U6391 ( .A1(n5816), .A2(n7835), .ZN(n5822) );
  OR2_X1 U6392 ( .A1(n8929), .A2(n5495), .ZN(n5502) );
  NAND2_X1 U6393 ( .A1(n5177), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5164) );
  INV_X1 U6394 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6643) );
  INV_X1 U6395 ( .A(n9156), .ZN(n8990) );
  AND2_X1 U6396 ( .A1(n9191), .A2(n8876), .ZN(n5582) );
  OR2_X1 U6397 ( .A1(n5282), .A2(n6643), .ZN(n5294) );
  OR2_X1 U6398 ( .A1(n5864), .A2(n7834), .ZN(n9104) );
  AND2_X1 U6399 ( .A1(n5514), .A2(n5513), .ZN(n9256) );
  OR2_X1 U6400 ( .A1(n6453), .A2(n5403), .ZN(n6906) );
  INV_X1 U6401 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5539) );
  OR2_X1 U6402 ( .A1(n7053), .A2(n5859), .ZN(n6226) );
  NOR2_X1 U6403 ( .A1(n6354), .A2(n6104), .ZN(n6213) );
  INV_X1 U6404 ( .A(n6082), .ZN(n8097) );
  OR2_X1 U6405 ( .A1(n8434), .A2(n7480), .ZN(n7451) );
  OR2_X1 U6406 ( .A1(n6237), .A2(n6253), .ZN(n9596) );
  INV_X1 U6407 ( .A(n9596), .ZN(n9594) );
  INV_X1 U6408 ( .A(n9611), .ZN(n8571) );
  INV_X1 U6409 ( .A(n9669), .ZN(n9618) );
  INV_X1 U6410 ( .A(n9644), .ZN(n9662) );
  INV_X1 U6411 ( .A(n9751), .ZN(n9776) );
  AND2_X1 U6412 ( .A1(n9640), .A2(n9755), .ZN(n9740) );
  INV_X1 U6413 ( .A(n9740), .ZN(n9783) );
  AND2_X1 U6414 ( .A1(n6226), .A2(n9690), .ZN(n9681) );
  NAND2_X1 U6415 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  AND2_X1 U6416 ( .A1(n5814), .A2(n5822), .ZN(n8839) );
  INV_X1 U6417 ( .A(n8812), .ZN(n8863) );
  AND2_X1 U6418 ( .A1(n5144), .A2(n5143), .ZN(n8904) );
  AND4_X1 U6419 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n9074)
         );
  INV_X1 U6420 ( .A(n9488), .ZN(n9477) );
  INV_X1 U6421 ( .A(n9496), .ZN(n9381) );
  AND2_X1 U6422 ( .A1(n5978), .A2(n5977), .ZN(n9496) );
  INV_X1 U6423 ( .A(n9342), .ZN(n7619) );
  AND2_X1 U6424 ( .A1(n7568), .A2(n7577), .ZN(n9071) );
  INV_X1 U6425 ( .A(n9506), .ZN(n9261) );
  AND2_X1 U6426 ( .A1(n9081), .A2(n6604), .ZN(n9068) );
  NAND2_X1 U6427 ( .A1(n7755), .A2(n7825), .ZN(n6603) );
  INV_X1 U6428 ( .A(n9117), .ZN(n9118) );
  INV_X1 U6429 ( .A(n9537), .ZN(n9198) );
  AND2_X1 U6430 ( .A1(n6346), .A2(n6345), .ZN(n6464) );
  XNOR2_X1 U6431 ( .A(n5512), .B(n5511), .ZN(n5598) );
  NOR2_X1 U6432 ( .A1(n10150), .A2(n9294), .ZN(n9295) );
  NAND2_X1 U6433 ( .A1(n5942), .A2(n5941), .ZN(n9600) );
  INV_X1 U6434 ( .A(n8682), .ZN(n8561) );
  INV_X1 U6435 ( .A(n8188), .ZN(n8244) );
  NAND2_X1 U6436 ( .A1(n6202), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9593) );
  NAND2_X1 U6437 ( .A1(n6141), .A2(n6134), .ZN(n8250) );
  OR2_X1 U6438 ( .A1(n8394), .A2(n6142), .ZN(n8390) );
  OR2_X1 U6439 ( .A1(n9669), .A2(n9617), .ZN(n9673) );
  NAND2_X1 U6440 ( .A1(n9681), .A2(n6745), .ZN(n9666) );
  INV_X1 U6441 ( .A(n9803), .ZN(n9801) );
  INV_X1 U6442 ( .A(n9785), .ZN(n9784) );
  INV_X1 U6443 ( .A(n9687), .ZN(n9685) );
  INV_X1 U6444 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7405) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10038) );
  INV_X1 U6446 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5903) );
  INV_X1 U6447 ( .A(n9176), .ZN(n9051) );
  INV_X1 U6448 ( .A(n9191), .ZN(n9095) );
  INV_X1 U6449 ( .A(n9186), .ZN(n9079) );
  INV_X1 U6450 ( .A(n8786), .ZN(n8959) );
  OR2_X1 U6451 ( .A1(P1_U3083), .A2(n9401), .ZN(n9481) );
  NAND2_X1 U6452 ( .A1(n9081), .A2(n5601), .ZN(n9114) );
  INV_X2 U6453 ( .A(n9081), .ZN(n9513) );
  INV_X1 U6454 ( .A(n9565), .ZN(n9563) );
  AND2_X1 U6455 ( .A1(n9544), .A2(n9543), .ZN(n9562) );
  AND2_X2 U6456 ( .A1(n6464), .A2(n6348), .ZN(n9556) );
  INV_X1 U6457 ( .A(n9515), .ZN(n9514) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7178) );
  INV_X1 U6459 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5947) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5897) );
  INV_X1 U6461 ( .A(n9221), .ZN(n8108) );
  NOR2_X1 U6462 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  NOR2_X1 U6463 ( .A1(n9832), .A2(n9831), .ZN(n9830) );
  AND2_X1 U6464 ( .A1(n5862), .A2(n9690), .ZN(P2_U3966) );
  NAND2_X1 U6465 ( .A1(n5608), .A2(n5607), .ZN(P1_U3263) );
  AND2_X1 U6466 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4983) );
  INV_X1 U6467 ( .A(SI_1_), .ZN(n4984) );
  NAND2_X1 U6468 ( .A1(n4985), .A2(SI_1_), .ZN(n4986) );
  INV_X1 U6469 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6105) );
  INV_X1 U6470 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5871) );
  XNOR2_X1 U6471 ( .A(n4987), .B(SI_2_), .ZN(n5172) );
  INV_X1 U6472 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6473 ( .A1(n4988), .A2(SI_2_), .ZN(n4989) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6205) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9921) );
  MUX2_X1 U6476 ( .A(n6205), .B(n9921), .S(n5868), .Z(n4990) );
  XNOR2_X1 U6477 ( .A(n4990), .B(SI_3_), .ZN(n5187) );
  NAND2_X1 U6478 ( .A1(n5186), .A2(n5187), .ZN(n4993) );
  INV_X1 U6479 ( .A(n4990), .ZN(n4991) );
  NAND2_X1 U6480 ( .A1(n4991), .A2(SI_3_), .ZN(n4992) );
  INV_X1 U6481 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6311) );
  INV_X1 U6482 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5872) );
  MUX2_X1 U6483 ( .A(n6311), .B(n5872), .S(n5868), .Z(n4994) );
  XNOR2_X1 U6484 ( .A(n4994), .B(SI_4_), .ZN(n5203) );
  INV_X1 U6485 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6486 ( .A1(n4995), .A2(SI_4_), .ZN(n4996) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6366) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5884) );
  MUX2_X1 U6489 ( .A(n6366), .B(n5884), .S(n4895), .Z(n4997) );
  XNOR2_X1 U6490 ( .A(n4997), .B(SI_5_), .ZN(n5227) );
  INV_X1 U6491 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6492 ( .A1(n4998), .A2(SI_5_), .ZN(n4999) );
  MUX2_X1 U6493 ( .A(n6419), .B(n5888), .S(n4895), .Z(n5000) );
  XNOR2_X1 U6494 ( .A(n5000), .B(SI_6_), .ZN(n5215) );
  INV_X1 U6495 ( .A(n5000), .ZN(n5001) );
  MUX2_X1 U6496 ( .A(n5892), .B(n5889), .S(n4895), .Z(n5002) );
  XNOR2_X1 U6497 ( .A(n5002), .B(SI_7_), .ZN(n5242) );
  INV_X1 U6498 ( .A(n5002), .ZN(n5003) );
  MUX2_X1 U6499 ( .A(n10084), .B(n5897), .S(n4895), .Z(n5004) );
  NAND2_X1 U6500 ( .A1(n5004), .A2(n10066), .ZN(n5007) );
  INV_X1 U6501 ( .A(n5004), .ZN(n5005) );
  NAND2_X1 U6502 ( .A1(n5005), .A2(SI_8_), .ZN(n5006) );
  MUX2_X1 U6503 ( .A(n5903), .B(n5898), .S(n4895), .Z(n5009) );
  INV_X1 U6504 ( .A(SI_9_), .ZN(n5008) );
  NAND2_X1 U6505 ( .A1(n5009), .A2(n5008), .ZN(n5012) );
  INV_X1 U6506 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6507 ( .A1(n5010), .A2(SI_9_), .ZN(n5011) );
  NAND2_X1 U6508 ( .A1(n5012), .A2(n5011), .ZN(n5273) );
  MUX2_X1 U6509 ( .A(n5926), .B(n5917), .S(n4895), .Z(n5013) );
  NAND2_X1 U6510 ( .A1(n5013), .A2(n9948), .ZN(n5017) );
  INV_X1 U6511 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6512 ( .A1(n5014), .A2(SI_10_), .ZN(n5015) );
  NAND2_X1 U6513 ( .A1(n5017), .A2(n5015), .ZN(n5016) );
  MUX2_X1 U6514 ( .A(n5020), .B(n5019), .S(n4895), .Z(n5021) );
  XNOR2_X1 U6515 ( .A(n5021), .B(SI_11_), .ZN(n5301) );
  INV_X1 U6516 ( .A(n5301), .ZN(n5024) );
  INV_X1 U6517 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6518 ( .A1(n5022), .A2(SI_11_), .ZN(n5023) );
  MUX2_X1 U6519 ( .A(n5946), .B(n5943), .S(n4895), .Z(n5026) );
  INV_X1 U6520 ( .A(SI_12_), .ZN(n5025) );
  INV_X1 U6521 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6522 ( .A1(n5027), .A2(SI_12_), .ZN(n5028) );
  NAND2_X1 U6523 ( .A1(n5029), .A2(n5028), .ZN(n5310) );
  MUX2_X1 U6524 ( .A(n10108), .B(n10120), .S(n4895), .Z(n5031) );
  INV_X1 U6525 ( .A(SI_13_), .ZN(n5030) );
  NAND2_X1 U6526 ( .A1(n5031), .A2(n5030), .ZN(n5333) );
  INV_X1 U6527 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6528 ( .A1(n5032), .A2(SI_13_), .ZN(n5033) );
  MUX2_X1 U6529 ( .A(n5953), .B(n5947), .S(n4895), .Z(n5035) );
  XNOR2_X1 U6530 ( .A(n5035), .B(SI_14_), .ZN(n5335) );
  NAND2_X1 U6531 ( .A1(n5334), .A2(n5034), .ZN(n5038) );
  INV_X1 U6532 ( .A(n5035), .ZN(n5036) );
  NAND2_X1 U6533 ( .A1(n5036), .A2(SI_14_), .ZN(n5037) );
  NAND2_X1 U6534 ( .A1(n5038), .A2(n5037), .ZN(n5347) );
  MUX2_X1 U6535 ( .A(n5970), .B(n9934), .S(n4895), .Z(n5039) );
  NAND2_X1 U6536 ( .A1(n5039), .A2(n10047), .ZN(n5042) );
  INV_X1 U6537 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6538 ( .A1(n5040), .A2(SI_15_), .ZN(n5041) );
  NAND2_X1 U6539 ( .A1(n5042), .A2(n5041), .ZN(n5346) );
  MUX2_X1 U6540 ( .A(n5043), .B(n5972), .S(n4895), .Z(n5044) );
  INV_X1 U6541 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6542 ( .A1(n5045), .A2(SI_16_), .ZN(n5046) );
  NAND2_X1 U6543 ( .A1(n5360), .A2(n5359), .ZN(n5048) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5049) );
  MUX2_X1 U6545 ( .A(n10038), .B(n5049), .S(n5868), .Z(n5050) );
  XNOR2_X1 U6546 ( .A(n5050), .B(SI_17_), .ZN(n5373) );
  INV_X1 U6547 ( .A(n5373), .ZN(n5053) );
  INV_X1 U6548 ( .A(n5050), .ZN(n5051) );
  NAND2_X1 U6549 ( .A1(n5051), .A2(SI_17_), .ZN(n5052) );
  MUX2_X1 U6550 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4895), .Z(n5054) );
  XNOR2_X1 U6551 ( .A(n5054), .B(SI_18_), .ZN(n5386) );
  MUX2_X1 U6552 ( .A(n6482), .B(n7546), .S(n4895), .Z(n5056) );
  INV_X1 U6553 ( .A(SI_19_), .ZN(n5055) );
  NAND2_X1 U6554 ( .A1(n5056), .A2(n5055), .ZN(n5059) );
  INV_X1 U6555 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6556 ( .A1(n5057), .A2(SI_19_), .ZN(n5058) );
  NAND2_X1 U6557 ( .A1(n5059), .A2(n5058), .ZN(n5398) );
  MUX2_X1 U6558 ( .A(n7846), .B(n9951), .S(n5868), .Z(n5061) );
  INV_X1 U6559 ( .A(SI_20_), .ZN(n5060) );
  NAND2_X1 U6560 ( .A1(n5061), .A2(n5060), .ZN(n5064) );
  INV_X1 U6561 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6562 ( .A1(n5062), .A2(SI_20_), .ZN(n5063) );
  MUX2_X1 U6563 ( .A(n7381), .B(n6547), .S(n4895), .Z(n5066) );
  XNOR2_X1 U6564 ( .A(n5066), .B(SI_21_), .ZN(n5424) );
  INV_X1 U6565 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6566 ( .A1(n5067), .A2(SI_21_), .ZN(n5068) );
  MUX2_X1 U6567 ( .A(n7392), .B(n6673), .S(n5868), .Z(n5069) );
  INV_X1 U6568 ( .A(SI_22_), .ZN(n10040) );
  NAND2_X1 U6569 ( .A1(n5069), .A2(n10040), .ZN(n5072) );
  INV_X1 U6570 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6571 ( .A1(n5070), .A2(SI_22_), .ZN(n5071) );
  NAND2_X1 U6572 ( .A1(n5072), .A2(n5071), .ZN(n5435) );
  MUX2_X1 U6573 ( .A(n10146), .B(n6813), .S(n4895), .Z(n5074) );
  INV_X1 U6574 ( .A(SI_23_), .ZN(n5073) );
  NAND2_X1 U6575 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  INV_X1 U6576 ( .A(n5074), .ZN(n5075) );
  NAND2_X1 U6577 ( .A1(n5075), .A2(SI_23_), .ZN(n5076) );
  MUX2_X1 U6578 ( .A(n7405), .B(n6988), .S(n4895), .Z(n5079) );
  XNOR2_X1 U6579 ( .A(n5079), .B(SI_24_), .ZN(n5455) );
  INV_X1 U6580 ( .A(n5455), .ZN(n5082) );
  INV_X1 U6581 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6582 ( .A1(n5080), .A2(SI_24_), .ZN(n5081) );
  MUX2_X1 U6583 ( .A(n7416), .B(n7178), .S(n5868), .Z(n5083) );
  INV_X1 U6584 ( .A(SI_25_), .ZN(n10050) );
  NAND2_X1 U6585 ( .A1(n5083), .A2(n10050), .ZN(n5086) );
  INV_X1 U6586 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6587 ( .A1(n5084), .A2(SI_25_), .ZN(n5085) );
  NAND2_X1 U6588 ( .A1(n5086), .A2(n5085), .ZN(n5465) );
  INV_X1 U6589 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7427) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7179) );
  MUX2_X1 U6591 ( .A(n7427), .B(n7179), .S(n4895), .Z(n5088) );
  INV_X1 U6592 ( .A(SI_26_), .ZN(n5087) );
  NAND2_X1 U6593 ( .A1(n5088), .A2(n5087), .ZN(n5091) );
  INV_X1 U6594 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6595 ( .A1(n5089), .A2(SI_26_), .ZN(n5090) );
  INV_X1 U6596 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7441) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7262) );
  MUX2_X1 U6598 ( .A(n7441), .B(n7262), .S(n4895), .Z(n5094) );
  INV_X1 U6599 ( .A(SI_27_), .ZN(n5093) );
  NAND2_X1 U6600 ( .A1(n5094), .A2(n5093), .ZN(n5097) );
  INV_X1 U6601 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6602 ( .A1(n5095), .A2(SI_27_), .ZN(n5096) );
  INV_X1 U6603 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7453) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8104) );
  MUX2_X1 U6605 ( .A(n7453), .B(n8104), .S(n4895), .Z(n7469) );
  XNOR2_X1 U6606 ( .A(n7469), .B(SI_28_), .ZN(n7466) );
  NOR2_X2 U6607 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5169) );
  NOR2_X1 U6608 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5106) );
  NOR2_X1 U6609 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5105) );
  NOR2_X1 U6610 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5104) );
  NAND4_X1 U6611 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n5108)
         );
  NAND4_X1 U6612 ( .A1(n5348), .A2(n5504), .A3(n5511), .A4(n5506), .ZN(n5107)
         );
  NOR2_X1 U6613 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  NAND2_X1 U6614 ( .A1(n8102), .A2(n7560), .ZN(n5114) );
  OR2_X1 U6615 ( .A1(n5185), .A2(n8104), .ZN(n5113) );
  NAND3_X1 U6616 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5221) );
  INV_X1 U6617 ( .A(n5221), .ZN(n5115) );
  NAND2_X1 U6618 ( .A1(n5115), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5233) );
  INV_X1 U6619 ( .A(n5233), .ZN(n5116) );
  NAND2_X1 U6620 ( .A1(n5116), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5254) );
  INV_X1 U6621 ( .A(n5254), .ZN(n5117) );
  NAND2_X1 U6622 ( .A1(n5117), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5266) );
  INV_X1 U6623 ( .A(n5315), .ZN(n5119) );
  NAND2_X1 U6624 ( .A1(n5119), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5327) );
  INV_X1 U6625 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6626 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5121) );
  INV_X1 U6627 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5391) );
  INV_X1 U6628 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5417) );
  INV_X1 U6629 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8829) );
  INV_X1 U6630 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8737) );
  INV_X1 U6631 ( .A(n5460), .ZN(n5125) );
  NAND2_X1 U6632 ( .A1(n5125), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5470) );
  INV_X1 U6633 ( .A(n5470), .ZN(n5126) );
  NAND2_X1 U6634 ( .A1(n5126), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5480) );
  INV_X1 U6635 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8851) );
  INV_X1 U6636 ( .A(n5492), .ZN(n5127) );
  NAND2_X1 U6637 ( .A1(n5127), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5494) );
  INV_X1 U6638 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6639 ( .A1(n5494), .A2(n5128), .ZN(n5129) );
  NAND2_X1 U6640 ( .A1(n5131), .A2(n5130), .ZN(n5135) );
  INV_X1 U6641 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5132) );
  INV_X1 U6642 ( .A(n5134), .ZN(n9219) );
  NAND2_X1 U6643 ( .A1(n5135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5136) );
  MUX2_X1 U6644 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5136), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5137) );
  NAND2_X1 U6645 ( .A1(n8766), .A2(n5516), .ZN(n5144) );
  NAND2_X1 U6646 ( .A1(n5176), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6647 ( .A1(n5496), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5140) );
  OAI211_X1 U6648 ( .C1(n5602), .C2(n5296), .A(n5141), .B(n5140), .ZN(n5142)
         );
  INV_X1 U6649 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6650 ( .A1(n9130), .A2(n8904), .ZN(n8909) );
  NAND2_X1 U6651 ( .A1(n5193), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6652 ( .A1(n5176), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6653 ( .A1(n5268), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5145) );
  INV_X1 U6654 ( .A(SI_0_), .ZN(n5150) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5149) );
  OAI21_X1 U6656 ( .B1(n7555), .B2(n5150), .A(n5149), .ZN(n5152) );
  AND2_X1 U6657 ( .A1(n5152), .A2(n5151), .ZN(n9224) );
  MUX2_X1 U6658 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9224), .S(n5168), .Z(n6605) );
  INV_X1 U6659 ( .A(n6605), .ZN(n6452) );
  NAND2_X1 U6660 ( .A1(n5193), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6661 ( .A1(n5176), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6662 ( .A1(n5268), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5153) );
  INV_X1 U6663 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5870) );
  OR2_X1 U6664 ( .A1(n5185), .A2(n5870), .ZN(n5161) );
  XNOR2_X1 U6665 ( .A(n5157), .B(n5158), .ZN(n6089) );
  INV_X1 U6666 ( .A(n9386), .ZN(n5869) );
  OR2_X1 U6667 ( .A1(n5168), .A2(n5869), .ZN(n5159) );
  AND3_X2 U6668 ( .A1(n5161), .A2(n5160), .A3(n5159), .ZN(n9507) );
  INV_X1 U6669 ( .A(n9507), .ZN(n5162) );
  INV_X1 U6670 ( .A(n5613), .ZN(n7866) );
  NAND2_X1 U6671 ( .A1(n7866), .A2(n5162), .ZN(n5163) );
  NAND2_X1 U6672 ( .A1(n6454), .A2(n5163), .ZN(n7597) );
  NAND2_X1 U6673 ( .A1(n5176), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6674 ( .A1(n5268), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6675 ( .A1(n5193), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5165) );
  OR2_X1 U6676 ( .A1(n5169), .A2(n9218), .ZN(n5171) );
  INV_X1 U6677 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6678 ( .A1(n5171), .A2(n5170), .ZN(n5182) );
  OAI21_X1 U6679 ( .B1(n5171), .B2(n5170), .A(n5182), .ZN(n9407) );
  OR2_X1 U6680 ( .A1(n5185), .A2(n5871), .ZN(n5175) );
  XNOR2_X1 U6681 ( .A(n5173), .B(n5172), .ZN(n6106) );
  OR2_X1 U6682 ( .A1(n5229), .A2(n6106), .ZN(n5174) );
  XNOR2_X1 U6683 ( .A(n5631), .B(n7869), .ZN(n7795) );
  NAND2_X1 U6684 ( .A1(n7597), .A2(n7795), .ZN(n6712) );
  INV_X1 U6685 ( .A(n5631), .ZN(n7596) );
  NAND2_X1 U6686 ( .A1(n7596), .A2(n7869), .ZN(n7599) );
  NAND2_X1 U6687 ( .A1(n6712), .A2(n7599), .ZN(n6536) );
  NAND2_X1 U6688 ( .A1(n5472), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6689 ( .A1(n5193), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6690 ( .A1(n5268), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5179) );
  INV_X1 U6691 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U6692 ( .A1(n5177), .A2(n6686), .ZN(n5178) );
  INV_X1 U6693 ( .A(n7867), .ZN(n8887) );
  NAND2_X1 U6694 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5184) );
  INV_X1 U6695 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U6696 ( .A(n5184), .B(n5183), .ZN(n5998) );
  OR2_X1 U6697 ( .A1(n5185), .A2(n9921), .ZN(n5189) );
  XNOR2_X1 U6698 ( .A(n5186), .B(n5187), .ZN(n6204) );
  OR2_X1 U6699 ( .A1(n5229), .A2(n6204), .ZN(n5188) );
  OAI211_X1 U6700 ( .C1(n5168), .C2(n5998), .A(n5189), .B(n5188), .ZN(n5190)
         );
  NAND2_X1 U6701 ( .A1(n8887), .A2(n6535), .ZN(n7591) );
  NAND2_X1 U6702 ( .A1(n6536), .A2(n7591), .ZN(n5191) );
  NAND2_X1 U6703 ( .A1(n7867), .A2(n5190), .ZN(n7757) );
  NAND2_X1 U6704 ( .A1(n5496), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6705 ( .A1(n5472), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5196) );
  INV_X1 U6706 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5192) );
  XNOR2_X1 U6707 ( .A(n5192), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U6708 ( .A1(n5516), .A2(n6526), .ZN(n5195) );
  NAND2_X1 U6709 ( .A1(n5193), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5194) );
  INV_X1 U6710 ( .A(n6556), .ZN(n8886) );
  NAND2_X1 U6711 ( .A1(n5198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5199) );
  MUX2_X1 U6712 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5199), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5201) );
  NAND2_X1 U6713 ( .A1(n5201), .A2(n5200), .ZN(n9417) );
  OR2_X1 U6714 ( .A1(n5185), .A2(n5872), .ZN(n5205) );
  XNOR2_X1 U6715 ( .A(n5202), .B(n5203), .ZN(n6309) );
  OR2_X1 U6716 ( .A1(n5229), .A2(n6309), .ZN(n5204) );
  OAI211_X1 U6717 ( .C1(n5168), .C2(n9417), .A(n5205), .B(n5204), .ZN(n6737)
         );
  INV_X1 U6718 ( .A(n6737), .ZN(n9524) );
  NAND2_X1 U6719 ( .A1(n8886), .A2(n9524), .ZN(n7657) );
  NAND2_X1 U6720 ( .A1(n6556), .A2(n6737), .ZN(n7758) );
  NAND2_X1 U6721 ( .A1(n5193), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6722 ( .A1(n5472), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5209) );
  INV_X1 U6723 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U6724 ( .A1(n5221), .A2(n10002), .ZN(n5206) );
  AND2_X1 U6725 ( .A1(n5233), .A2(n5206), .ZN(n6874) );
  NAND2_X1 U6726 ( .A1(n5516), .A2(n6874), .ZN(n5208) );
  NAND2_X1 U6727 ( .A1(n5268), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5207) );
  INV_X1 U6728 ( .A(n7853), .ZN(n8884) );
  INV_X1 U6729 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9218) );
  OR2_X1 U6730 ( .A1(n5211), .A2(n9218), .ZN(n5213) );
  XNOR2_X1 U6731 ( .A(n5213), .B(n5212), .ZN(n6039) );
  OR2_X1 U6732 ( .A1(n5185), .A2(n5888), .ZN(n5217) );
  XNOR2_X1 U6733 ( .A(n5214), .B(n5215), .ZN(n6418) );
  OR2_X1 U6734 ( .A1(n5229), .A2(n6418), .ZN(n5216) );
  OAI211_X1 U6735 ( .C1(n5168), .C2(n6039), .A(n5217), .B(n5216), .ZN(n5527)
         );
  INV_X1 U6736 ( .A(n5527), .ZN(n6914) );
  NAND2_X1 U6737 ( .A1(n5472), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6738 ( .A1(n5193), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5224) );
  INV_X1 U6739 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6740 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5218) );
  NAND2_X1 U6741 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  AND2_X1 U6742 ( .A1(n5221), .A2(n5220), .ZN(n6679) );
  NAND2_X1 U6743 ( .A1(n5516), .A2(n6679), .ZN(n5223) );
  NAND2_X1 U6744 ( .A1(n5268), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6745 ( .A1(n5200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6746 ( .A(n5226), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6023) );
  INV_X1 U6747 ( .A(n6023), .ZN(n6030) );
  XNOR2_X1 U6748 ( .A(n5228), .B(n5227), .ZN(n6365) );
  OR2_X1 U6749 ( .A1(n5229), .A2(n6365), .ZN(n5231) );
  OR2_X1 U6750 ( .A1(n5185), .A2(n5884), .ZN(n5230) );
  OAI211_X1 U6751 ( .C1(n5168), .C2(n6030), .A(n5231), .B(n5230), .ZN(n5247)
         );
  INV_X1 U6752 ( .A(n5247), .ZN(n6553) );
  NAND2_X1 U6753 ( .A1(n8885), .A2(n6553), .ZN(n7656) );
  AND2_X1 U6754 ( .A1(n7660), .A2(n7656), .ZN(n7601) );
  NAND2_X1 U6755 ( .A1(n5496), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6756 ( .A1(n5472), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5237) );
  INV_X1 U6757 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6758 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  AND2_X1 U6759 ( .A1(n5254), .A2(n5234), .ZN(n7859) );
  NAND2_X1 U6760 ( .A1(n5516), .A2(n7859), .ZN(n5236) );
  NAND2_X1 U6761 ( .A1(n5193), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5235) );
  OR2_X1 U6762 ( .A1(n5239), .A2(n9218), .ZN(n5241) );
  XNOR2_X1 U6763 ( .A(n5241), .B(n5240), .ZN(n6061) );
  OR2_X1 U6764 ( .A1(n5185), .A2(n5889), .ZN(n5244) );
  OR2_X1 U6765 ( .A1(n5229), .A2(n6429), .ZN(n5243) );
  OAI211_X1 U6766 ( .C1(n5168), .C2(n6061), .A(n5244), .B(n5243), .ZN(n6981)
         );
  NAND2_X1 U6767 ( .A1(n6904), .A2(n6981), .ZN(n7625) );
  INV_X1 U6768 ( .A(n6981), .ZN(n7857) );
  AND2_X1 U6769 ( .A1(n7601), .A2(n5246), .ZN(n5245) );
  NAND2_X1 U6770 ( .A1(n6555), .A2(n5245), .ZN(n5253) );
  INV_X1 U6771 ( .A(n5246), .ZN(n5251) );
  NAND2_X1 U6772 ( .A1(n6905), .A2(n5247), .ZN(n7761) );
  INV_X1 U6773 ( .A(n7761), .ZN(n5248) );
  NAND2_X1 U6774 ( .A1(n7601), .A2(n5248), .ZN(n5249) );
  NAND2_X1 U6775 ( .A1(n7853), .A2(n5527), .ZN(n7762) );
  AND2_X1 U6776 ( .A1(n5249), .A2(n7762), .ZN(n7602) );
  AND2_X1 U6777 ( .A1(n7602), .A2(n7625), .ZN(n5250) );
  OR2_X1 U6778 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  NAND2_X1 U6779 ( .A1(n5253), .A2(n5252), .ZN(n6699) );
  NAND2_X1 U6780 ( .A1(n5496), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6781 ( .A1(n5472), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5258) );
  INV_X1 U6782 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U6783 ( .A1(n5254), .A2(n6052), .ZN(n5255) );
  AND2_X1 U6784 ( .A1(n5266), .A2(n5255), .ZN(n7012) );
  NAND2_X1 U6785 ( .A1(n5516), .A2(n7012), .ZN(n5257) );
  NAND2_X1 U6786 ( .A1(n5193), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6787 ( .A1(n5260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6788 ( .A(n5261), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6180) );
  INV_X1 U6789 ( .A(n6180), .ZN(n6165) );
  OR2_X1 U6790 ( .A1(n5185), .A2(n5897), .ZN(n5263) );
  NAND2_X1 U6791 ( .A1(n6801), .A2(n7018), .ZN(n7629) );
  INV_X1 U6792 ( .A(n7629), .ZN(n5264) );
  INV_X1 U6793 ( .A(n7018), .ZN(n9539) );
  NAND2_X1 U6794 ( .A1(n8882), .A2(n9539), .ZN(n7627) );
  NAND2_X1 U6795 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  AND2_X1 U6796 ( .A1(n5282), .A2(n5267), .ZN(n6945) );
  NAND2_X1 U6797 ( .A1(n5516), .A2(n6945), .ZN(n5272) );
  NAND2_X1 U6798 ( .A1(n5472), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6799 ( .A1(n5193), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6800 ( .A1(n5268), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5269) );
  XNOR2_X1 U6801 ( .A(n5274), .B(n5273), .ZN(n6569) );
  OR2_X1 U6802 ( .A1(n5229), .A2(n6569), .ZN(n5280) );
  OR2_X1 U6803 ( .A1(n5185), .A2(n5898), .ZN(n5278) );
  INV_X1 U6804 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6805 ( .A1(n5276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5277) );
  XNOR2_X1 U6806 ( .A(n5277), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9441) );
  INV_X1 U6807 ( .A(n9441), .ZN(n5899) );
  INV_X1 U6808 ( .A(n6949), .ZN(n9547) );
  AND2_X1 U6809 ( .A1(n9253), .A2(n9547), .ZN(n6759) );
  INV_X1 U6810 ( .A(n9253), .ZN(n5281) );
  NAND2_X1 U6811 ( .A1(n5281), .A2(n6949), .ZN(n7630) );
  NAND2_X1 U6812 ( .A1(n5496), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6813 ( .A1(n5472), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6814 ( .A1(n5282), .A2(n6643), .ZN(n5283) );
  AND2_X1 U6815 ( .A1(n5294), .A2(n5283), .ZN(n9260) );
  NAND2_X1 U6816 ( .A1(n5516), .A2(n9260), .ZN(n5285) );
  NAND2_X1 U6817 ( .A1(n5193), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6818 ( .A1(n5288), .A2(n9218), .ZN(n5304) );
  XNOR2_X1 U6819 ( .A(n5304), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9444) );
  AOI22_X1 U6820 ( .A1(n5404), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5866), .B2(
        n9444), .ZN(n5292) );
  XNOR2_X1 U6821 ( .A(n5290), .B(n5289), .ZN(n6584) );
  NAND2_X1 U6822 ( .A1(n6584), .A2(n7560), .ZN(n5291) );
  NAND2_X1 U6823 ( .A1(n5292), .A2(n5291), .ZN(n9263) );
  NAND2_X1 U6824 ( .A1(n7144), .A2(n9263), .ZN(n7634) );
  INV_X1 U6825 ( .A(n7144), .ZN(n8881) );
  NAND2_X1 U6826 ( .A1(n8881), .A2(n9274), .ZN(n7632) );
  NAND2_X1 U6827 ( .A1(n5472), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6828 ( .A1(n5496), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5299) );
  INV_X1 U6829 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6830 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  AND2_X1 U6831 ( .A1(n5315), .A2(n5295), .ZN(n7150) );
  NAND2_X1 U6832 ( .A1(n5516), .A2(n7150), .ZN(n5298) );
  NAND2_X1 U6833 ( .A1(n5193), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5297) );
  NAND4_X1 U6834 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n9252)
         );
  INV_X1 U6835 ( .A(n9252), .ZN(n6646) );
  NAND2_X1 U6836 ( .A1(n6655), .A2(n7560), .ZN(n5308) );
  INV_X1 U6837 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6838 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6839 ( .A1(n5305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5306) );
  XNOR2_X1 U6840 ( .A(n5306), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9457) );
  AOI22_X1 U6841 ( .A1(n5404), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5866), .B2(
        n9457), .ZN(n5307) );
  NAND2_X1 U6842 ( .A1(n6646), .A2(n7151), .ZN(n7586) );
  NAND2_X1 U6843 ( .A1(n7249), .A2(n9252), .ZN(n7580) );
  NAND2_X1 U6844 ( .A1(n5309), .A2(n7580), .ZN(n7209) );
  XNOR2_X1 U6845 ( .A(n5311), .B(n5310), .ZN(n6952) );
  NAND2_X1 U6846 ( .A1(n6952), .A2(n7560), .ZN(n5314) );
  NAND2_X1 U6847 ( .A1(n5322), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6848 ( .A(n5312), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6474) );
  AOI22_X1 U6849 ( .A1(n5404), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5866), .B2(
        n6474), .ZN(n5313) );
  NAND2_X1 U6850 ( .A1(n5314), .A2(n5313), .ZN(n7215) );
  NAND2_X1 U6851 ( .A1(n5472), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6852 ( .A1(n5193), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5319) );
  INV_X1 U6853 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U6854 ( .A1(n5315), .A2(n6162), .ZN(n5316) );
  AND2_X1 U6855 ( .A1(n5327), .A2(n5316), .ZN(n7214) );
  NAND2_X1 U6856 ( .A1(n5516), .A2(n7214), .ZN(n5318) );
  NAND2_X1 U6857 ( .A1(n5496), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6858 ( .A1(n7215), .A2(n7143), .ZN(n7667) );
  NAND2_X1 U6859 ( .A1(n7215), .A2(n7143), .ZN(n7635) );
  XNOR2_X1 U6860 ( .A(n5321), .B(n4978), .ZN(n7057) );
  NAND2_X1 U6861 ( .A1(n7057), .A2(n7560), .ZN(n5325) );
  NAND2_X1 U6862 ( .A1(n5337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5323) );
  XNOR2_X1 U6863 ( .A(n5323), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U6864 ( .A1(n5404), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5866), .B2(
        n6925), .ZN(n5324) );
  NAND2_X1 U6865 ( .A1(n5496), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6866 ( .A1(n5472), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6867 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  AND2_X1 U6868 ( .A1(n5340), .A2(n5328), .ZN(n7275) );
  NAND2_X1 U6869 ( .A1(n5516), .A2(n7275), .ZN(n5330) );
  NAND2_X1 U6870 ( .A1(n5193), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5329) );
  NAND4_X1 U6871 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8879)
         );
  NAND2_X1 U6872 ( .A1(n7276), .A2(n7126), .ZN(n7585) );
  OR2_X1 U6873 ( .A1(n7276), .A2(n7126), .ZN(n7579) );
  NAND2_X1 U6874 ( .A1(n5334), .A2(n5333), .ZN(n5336) );
  XNOR2_X1 U6875 ( .A(n5336), .B(n5335), .ZN(n7094) );
  NAND2_X1 U6876 ( .A1(n7094), .A2(n7560), .ZN(n5339) );
  NOR2_X2 U6877 ( .A1(n5337), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6878 ( .A1(n5362), .A2(n9218), .ZN(n5349) );
  XNOR2_X1 U6879 ( .A(n5349), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U6880 ( .A1(n5404), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5866), .B2(
        n9469), .ZN(n5338) );
  NAND2_X1 U6881 ( .A1(n5472), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6882 ( .A1(n5193), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5344) );
  INV_X1 U6883 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U6884 ( .A1(n5340), .A2(n9996), .ZN(n5341) );
  AND2_X1 U6885 ( .A1(n5367), .A2(n5341), .ZN(n7298) );
  NAND2_X1 U6886 ( .A1(n5516), .A2(n7298), .ZN(n5343) );
  NAND2_X1 U6887 ( .A1(n5496), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5342) );
  NAND4_X1 U6888 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n8878)
         );
  XNOR2_X1 U6889 ( .A(n7583), .B(n9102), .ZN(n7809) );
  OR2_X1 U6890 ( .A1(n7583), .A2(n9102), .ZN(n7644) );
  XNOR2_X1 U6891 ( .A(n5347), .B(n5346), .ZN(n7183) );
  NAND2_X1 U6892 ( .A1(n7183), .A2(n7560), .ZN(n5354) );
  NAND2_X1 U6893 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  NAND2_X1 U6894 ( .A1(n5350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5352) );
  INV_X1 U6895 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5351) );
  XNOR2_X1 U6896 ( .A(n5352), .B(n5351), .ZN(n7163) );
  INV_X1 U6897 ( .A(n7163), .ZN(n6929) );
  AOI22_X1 U6898 ( .A1(n5404), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5866), .B2(
        n6929), .ZN(n5353) );
  NAND2_X1 U6899 ( .A1(n5472), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6900 ( .A1(n5496), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5357) );
  XNOR2_X1 U6901 ( .A(n5367), .B(P1_REG3_REG_15__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U6902 ( .A1(n5516), .A2(n9107), .ZN(n5356) );
  NAND2_X1 U6903 ( .A1(n5193), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5355) );
  NAND4_X1 U6904 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n8877)
         );
  AND2_X1 U6905 ( .A1(n9111), .A2(n8877), .ZN(n7641) );
  NAND2_X1 U6906 ( .A1(n9196), .A2(n9087), .ZN(n7677) );
  XNOR2_X1 U6907 ( .A(n5360), .B(n5359), .ZN(n7305) );
  NAND2_X1 U6908 ( .A1(n7305), .A2(n7560), .ZN(n5365) );
  NOR2_X1 U6909 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5361) );
  NAND2_X1 U6910 ( .A1(n5375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U6911 ( .A(n5363), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7538) );
  AOI22_X1 U6912 ( .A1(n5404), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5866), .B2(
        n7538), .ZN(n5364) );
  NAND2_X1 U6913 ( .A1(n5496), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6914 ( .A1(n5472), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5371) );
  INV_X1 U6915 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6928) );
  INV_X1 U6916 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5366) );
  OAI21_X1 U6917 ( .B1(n5367), .B2(n6928), .A(n5366), .ZN(n5368) );
  AND2_X1 U6918 ( .A1(n5368), .A2(n5378), .ZN(n9092) );
  NAND2_X1 U6919 ( .A1(n5516), .A2(n9092), .ZN(n5370) );
  NAND2_X1 U6920 ( .A1(n5193), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6921 ( .A1(n9191), .A2(n9103), .ZN(n7682) );
  NAND2_X1 U6922 ( .A1(n9191), .A2(n9103), .ZN(n7681) );
  NAND2_X1 U6923 ( .A1(n7682), .A2(n7681), .ZN(n9084) );
  INV_X1 U6924 ( .A(n9084), .ZN(n7679) );
  INV_X1 U6925 ( .A(n7681), .ZN(n7610) );
  XNOR2_X1 U6926 ( .A(n5374), .B(n5373), .ZN(n7361) );
  NAND2_X1 U6927 ( .A1(n7361), .A2(n7560), .ZN(n5377) );
  NAND2_X1 U6928 ( .A1(n4438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6929 ( .A(n5401), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8891) );
  AOI22_X1 U6930 ( .A1(n5404), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5866), .B2(
        n8891), .ZN(n5376) );
  NAND2_X1 U6931 ( .A1(n5472), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6932 ( .A1(n5193), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5382) );
  INV_X1 U6933 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U6934 ( .A1(n5378), .A2(n10033), .ZN(n5379) );
  AND2_X1 U6935 ( .A1(n5392), .A2(n5379), .ZN(n9076) );
  NAND2_X1 U6936 ( .A1(n5516), .A2(n9076), .ZN(n5381) );
  NAND2_X1 U6937 ( .A1(n5496), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5380) );
  NAND4_X1 U6938 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n9063)
         );
  OR2_X1 U6939 ( .A1(n9186), .A2(n9088), .ZN(n7568) );
  NAND2_X1 U6940 ( .A1(n9186), .A2(n9088), .ZN(n7577) );
  INV_X1 U6941 ( .A(n7568), .ZN(n5384) );
  AOI21_X2 U6942 ( .B1(n9072), .B2(n9071), .A(n5384), .ZN(n9060) );
  XNOR2_X1 U6943 ( .A(n5385), .B(n5386), .ZN(n7368) );
  NAND2_X1 U6944 ( .A1(n7368), .A2(n7560), .ZN(n5390) );
  NAND2_X1 U6945 ( .A1(n5401), .A2(n5505), .ZN(n5387) );
  NAND2_X1 U6946 ( .A1(n5387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5388) );
  XNOR2_X1 U6947 ( .A(n5388), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9482) );
  AOI22_X1 U6948 ( .A1(n5404), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5866), .B2(
        n9482), .ZN(n5389) );
  NAND2_X1 U6949 ( .A1(n5472), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6950 ( .A1(n5193), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6951 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  AND2_X1 U6952 ( .A1(n5407), .A2(n5393), .ZN(n9057) );
  NAND2_X1 U6953 ( .A1(n5516), .A2(n9057), .ZN(n5395) );
  NAND2_X1 U6954 ( .A1(n5496), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6955 ( .A1(n9179), .A2(n9074), .ZN(n7690) );
  NAND2_X1 U6956 ( .A1(n9179), .A2(n9074), .ZN(n7578) );
  NAND2_X1 U6957 ( .A1(n7690), .A2(n7578), .ZN(n9054) );
  INV_X1 U6958 ( .A(n9054), .ZN(n9061) );
  NAND2_X1 U6959 ( .A1(n9060), .A2(n9061), .ZN(n9059) );
  NAND2_X1 U6960 ( .A1(n9059), .A2(n7578), .ZN(n9043) );
  XNOR2_X1 U6961 ( .A(n5399), .B(n5398), .ZN(n7358) );
  NAND2_X1 U6962 ( .A1(n7358), .A2(n7560), .ZN(n5406) );
  OAI21_X1 U6963 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6964 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  XNOR2_X2 U6965 ( .A(n5402), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5543) );
  AOI22_X1 U6966 ( .A1(n5404), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5866), .B2(
        n5403), .ZN(n5405) );
  NAND2_X1 U6967 ( .A1(n5496), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6968 ( .A1(n5472), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5411) );
  INV_X1 U6969 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U6970 ( .A1(n5407), .A2(n8748), .ZN(n5408) );
  AND2_X1 U6971 ( .A1(n5418), .A2(n5408), .ZN(n9048) );
  NAND2_X1 U6972 ( .A1(n5516), .A2(n9048), .ZN(n5410) );
  NAND2_X1 U6973 ( .A1(n5193), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5409) );
  NAND4_X1 U6974 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n9062)
         );
  INV_X1 U6975 ( .A(n9062), .ZN(n5748) );
  NOR2_X1 U6976 ( .A1(n9176), .A2(n5748), .ZN(n7692) );
  NOR2_X1 U6977 ( .A1(n7692), .A2(n7693), .ZN(n9044) );
  XNOR2_X1 U6978 ( .A(n5414), .B(n5413), .ZN(n7529) );
  NAND2_X1 U6979 ( .A1(n7529), .A2(n7560), .ZN(n5416) );
  OR2_X1 U6980 ( .A1(n5185), .A2(n9951), .ZN(n5415) );
  NAND2_X1 U6981 ( .A1(n5472), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6982 ( .A1(n5496), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6983 ( .A1(n5418), .A2(n5417), .ZN(n5419) );
  AND2_X1 U6984 ( .A1(n5429), .A2(n5419), .ZN(n9026) );
  NAND2_X1 U6985 ( .A1(n5516), .A2(n9026), .ZN(n5421) );
  NAND2_X1 U6986 ( .A1(n5193), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6987 ( .A1(n9169), .A2(n9046), .ZN(n7794) );
  XNOR2_X1 U6988 ( .A(n5425), .B(n5424), .ZN(n7380) );
  NAND2_X1 U6989 ( .A1(n7380), .A2(n7560), .ZN(n5427) );
  OR2_X1 U6990 ( .A1(n5185), .A2(n6547), .ZN(n5426) );
  NAND2_X1 U6991 ( .A1(n5472), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6992 ( .A1(n5193), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5433) );
  INV_X1 U6993 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6994 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  AND2_X1 U6995 ( .A1(n5439), .A2(n5430), .ZN(n9010) );
  NAND2_X1 U6996 ( .A1(n5516), .A2(n9010), .ZN(n5432) );
  NAND2_X1 U6997 ( .A1(n5496), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6998 ( .A1(n9165), .A2(n9029), .ZN(n7702) );
  NAND2_X1 U6999 ( .A1(n9165), .A2(n9029), .ZN(n7703) );
  NAND2_X1 U7000 ( .A1(n7702), .A2(n7703), .ZN(n9006) );
  INV_X1 U7001 ( .A(n9006), .ZN(n9014) );
  XNOR2_X1 U7002 ( .A(n5436), .B(n5435), .ZN(n7391) );
  NAND2_X1 U7003 ( .A1(n7391), .A2(n7560), .ZN(n5438) );
  OR2_X1 U7004 ( .A1(n5185), .A2(n6673), .ZN(n5437) );
  NAND2_X1 U7005 ( .A1(n5472), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7006 ( .A1(n5496), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7007 ( .A1(n5439), .A2(n8829), .ZN(n5440) );
  AND2_X1 U7008 ( .A1(n5449), .A2(n5440), .ZN(n8995) );
  NAND2_X1 U7009 ( .A1(n5516), .A2(n8995), .ZN(n5442) );
  NAND2_X1 U7010 ( .A1(n5193), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5441) );
  AOI21_X1 U7011 ( .B1(n8998), .B2(n7792), .A(n7791), .ZN(n8981) );
  NAND2_X1 U7012 ( .A1(n7333), .A2(n7560), .ZN(n5448) );
  OR2_X1 U7013 ( .A1(n5185), .A2(n6813), .ZN(n5447) );
  NAND2_X1 U7014 ( .A1(n5449), .A2(n8737), .ZN(n5450) );
  AND2_X1 U7015 ( .A1(n5460), .A2(n5450), .ZN(n8987) );
  NAND2_X1 U7016 ( .A1(n8987), .A2(n5516), .ZN(n5454) );
  NAND2_X1 U7017 ( .A1(n5472), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U7018 ( .A1(n5496), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7019 ( .A1(n5193), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5451) );
  NAND4_X1 U7020 ( .A1(n5454), .A2(n5453), .A3(n5452), .A4(n5451), .ZN(n9000)
         );
  XNOR2_X1 U7021 ( .A(n9156), .B(n9000), .ZN(n8980) );
  NAND2_X1 U7022 ( .A1(n8981), .A2(n8980), .ZN(n8979) );
  XNOR2_X1 U7023 ( .A(n5456), .B(n5455), .ZN(n7404) );
  NAND2_X1 U7024 ( .A1(n7404), .A2(n7560), .ZN(n5458) );
  OR2_X1 U7025 ( .A1(n5185), .A2(n6988), .ZN(n5457) );
  INV_X1 U7026 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7027 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U7028 ( .A1(n5470), .A2(n5461), .ZN(n8974) );
  INV_X1 U7029 ( .A(n5516), .ZN(n5495) );
  OR2_X1 U7030 ( .A1(n8974), .A2(n5495), .ZN(n5464) );
  AOI22_X1 U7031 ( .A1(n5472), .A2(P1_REG0_REG_24__SCAN_IN), .B1(n5193), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U7032 ( .A1(n5496), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7033 ( .A1(n9150), .A2(n8738), .ZN(n7709) );
  INV_X1 U7034 ( .A(n9000), .ZN(n10145) );
  OR2_X1 U7035 ( .A1(n9156), .A2(n10145), .ZN(n8965) );
  NAND3_X1 U7036 ( .A1(n8979), .A2(n8967), .A3(n8965), .ZN(n8966) );
  NAND2_X1 U7037 ( .A1(n7415), .A2(n7560), .ZN(n5468) );
  OR2_X1 U7038 ( .A1(n5185), .A2(n7178), .ZN(n5467) );
  INV_X1 U7039 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7040 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7041 ( .A1(n5480), .A2(n5471), .ZN(n8784) );
  OR2_X1 U7042 ( .A1(n8784), .A2(n5495), .ZN(n5475) );
  AOI22_X1 U7043 ( .A1(n5496), .A2(P1_REG1_REG_25__SCAN_IN), .B1(n5472), .B2(
        P1_REG0_REG_25__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7044 ( .A1(n5193), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7045 ( .A1(n9144), .A2(n8853), .ZN(n7717) );
  INV_X1 U7046 ( .A(n7717), .ZN(n7724) );
  XNOR2_X1 U7047 ( .A(n5477), .B(n5476), .ZN(n7426) );
  NAND2_X1 U7048 ( .A1(n7426), .A2(n7560), .ZN(n5479) );
  OR2_X1 U7049 ( .A1(n5185), .A2(n7179), .ZN(n5478) );
  NAND2_X1 U7050 ( .A1(n5480), .A2(n8851), .ZN(n5481) );
  NAND2_X1 U7051 ( .A1(n8942), .A2(n5516), .ZN(n5487) );
  INV_X1 U7052 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7053 ( .A1(n5472), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7054 ( .A1(n5193), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U7055 ( .C1(n5520), .C2(n5484), .A(n5483), .B(n5482), .ZN(n5485)
         );
  INV_X1 U7056 ( .A(n5485), .ZN(n5486) );
  NAND2_X1 U7057 ( .A1(n9139), .A2(n8786), .ZN(n7789) );
  NAND2_X1 U7058 ( .A1(n7440), .A2(n7560), .ZN(n5491) );
  OR2_X1 U7059 ( .A1(n5185), .A2(n7262), .ZN(n5490) );
  INV_X1 U7060 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U7061 ( .A1(n5492), .A2(n10090), .ZN(n5493) );
  NAND2_X1 U7062 ( .A1(n5494), .A2(n5493), .ZN(n8929) );
  INV_X1 U7063 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U7064 ( .A1(n5496), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7065 ( .A1(n5193), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5497) );
  OAI211_X1 U7066 ( .C1(n5499), .C2(n9952), .A(n5498), .B(n5497), .ZN(n5500)
         );
  INV_X1 U7067 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U7068 ( .A1(n9134), .A2(n8854), .ZN(n7731) );
  INV_X1 U7069 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7070 ( .A1(n5509), .A2(n5506), .ZN(n5507) );
  NAND2_X1 U7071 ( .A1(n7838), .A2(n5403), .ZN(n5514) );
  NAND2_X1 U7072 ( .A1(n5599), .A2(n7831), .ZN(n5513) );
  INV_X1 U7073 ( .A(n5515), .ZN(n8920) );
  NAND2_X1 U7074 ( .A1(n8920), .A2(n5516), .ZN(n5523) );
  INV_X1 U7075 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7076 ( .A1(n5472), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7077 ( .A1(n5193), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U7078 ( .C1(n5520), .C2(n5519), .A(n5518), .B(n5517), .ZN(n5521)
         );
  INV_X1 U7079 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7080 ( .A1(n5523), .A2(n5522), .ZN(n8874) );
  NAND2_X1 U7081 ( .A1(n7838), .A2(n5599), .ZN(n5864) );
  INV_X1 U7082 ( .A(n5524), .ZN(n7834) );
  INV_X1 U7083 ( .A(n5864), .ZN(n7824) );
  INV_X1 U7084 ( .A(n9254), .ZN(n5525) );
  INV_X1 U7085 ( .A(n5526), .ZN(n9132) );
  NAND2_X1 U7086 ( .A1(n9507), .A2(n6452), .ZN(n6717) );
  NAND2_X1 U7087 ( .A1(n6734), .A2(n9524), .ZN(n6733) );
  INV_X1 U7088 ( .A(n7215), .ZN(n9357) );
  NAND2_X1 U7089 ( .A1(n9047), .A2(n9028), .ZN(n9023) );
  INV_X1 U7090 ( .A(n8928), .ZN(n5529) );
  INV_X1 U7091 ( .A(n6603), .ZN(n6350) );
  INV_X1 U7092 ( .A(n8918), .ZN(n5528) );
  AOI211_X1 U7093 ( .C1(n9130), .C2(n5529), .A(n9548), .B(n5528), .ZN(n9129)
         );
  NAND2_X1 U7094 ( .A1(n4447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7095 ( .A1(n5533), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U7096 ( .A1(n5531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5532) );
  XNOR2_X1 U7097 ( .A(n5533), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7098 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5535) );
  XNOR2_X1 U7099 ( .A(n5535), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5544) );
  INV_X1 U7100 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U7101 ( .A1(n5538), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5540) );
  XNOR2_X1 U7102 ( .A(n5540), .B(n5539), .ZN(n6811) );
  AND2_X1 U7103 ( .A1(n6811), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7104 ( .A1(n7825), .A2(n7835), .ZN(n5542) );
  AOI22_X1 U7105 ( .A1(n9129), .A2(n5543), .B1(n8766), .B2(n9261), .ZN(n5563)
         );
  INV_X1 U7106 ( .A(n6602), .ZN(n7832) );
  INV_X1 U7107 ( .A(n5545), .ZN(n7176) );
  NAND3_X1 U7108 ( .A1(n7176), .A2(P1_B_REG_SCAN_IN), .A3(n6989), .ZN(n5546)
         );
  NOR4_X1 U7109 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5550) );
  NOR4_X1 U7110 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5549) );
  NOR4_X1 U7111 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5548) );
  NOR4_X1 U7112 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U7113 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n5556)
         );
  NOR2_X1 U7114 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n5554) );
  NOR4_X1 U7115 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5553) );
  NOR4_X1 U7116 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5552) );
  NOR4_X1 U7117 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5551) );
  NAND4_X1 U7118 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .ZN(n5555)
         );
  NOR2_X1 U7119 ( .A1(n5556), .A2(n5555), .ZN(n6341) );
  AND2_X1 U7120 ( .A1(n6341), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5557) );
  OR2_X1 U7121 ( .A1(n6342), .A2(n5557), .ZN(n5559) );
  INV_X1 U7122 ( .A(n5558), .ZN(n7180) );
  NAND2_X1 U7123 ( .A1(n7180), .A2(n7176), .ZN(n6340) );
  NAND2_X1 U7124 ( .A1(n5559), .A2(n6340), .ZN(n5811) );
  INV_X1 U7125 ( .A(n5811), .ZN(n5561) );
  OR2_X1 U7126 ( .A1(n6342), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7127 ( .A1(n7180), .A2(n6989), .ZN(n9217) );
  NAND2_X1 U7128 ( .A1(n5561), .A2(n6461), .ZN(n5562) );
  AOI21_X1 U7129 ( .B1(n9132), .B2(n5563), .A(n9513), .ZN(n5564) );
  AND2_X1 U7130 ( .A1(n5619), .A2(n6605), .ZN(n6450) );
  NAND2_X1 U7131 ( .A1(n5613), .A2(n5162), .ZN(n5565) );
  NAND2_X1 U7132 ( .A1(n6449), .A2(n5565), .ZN(n6711) );
  INV_X1 U7133 ( .A(n7869), .ZN(n9517) );
  NAND2_X1 U7134 ( .A1(n7596), .A2(n9517), .ZN(n5567) );
  NAND2_X1 U7135 ( .A1(n7757), .A2(n7591), .ZN(n6537) );
  NAND2_X1 U7136 ( .A1(n7867), .A2(n6535), .ZN(n5568) );
  NAND2_X1 U7137 ( .A1(n6531), .A2(n5568), .ZN(n6725) );
  NAND2_X1 U7138 ( .A1(n7758), .A2(n7657), .ZN(n6727) );
  NAND2_X1 U7139 ( .A1(n6725), .A2(n6727), .ZN(n6724) );
  AND2_X1 U7140 ( .A1(n7853), .A2(n6914), .ZN(n5571) );
  OR2_X1 U7141 ( .A1(n6902), .A2(n5571), .ZN(n6790) );
  AND2_X1 U7142 ( .A1(n6904), .A2(n7857), .ZN(n5572) );
  NOR2_X1 U7143 ( .A1(n6790), .A2(n5572), .ZN(n5569) );
  NAND2_X1 U7144 ( .A1(n6556), .A2(n9524), .ZN(n6550) );
  AND2_X1 U7145 ( .A1(n5569), .A2(n6550), .ZN(n5570) );
  NAND2_X1 U7146 ( .A1(n6724), .A2(n5570), .ZN(n6695) );
  NAND2_X1 U7147 ( .A1(n7762), .A2(n7660), .ZN(n6901) );
  NAND2_X1 U7148 ( .A1(n8885), .A2(n5247), .ZN(n6895) );
  AND2_X1 U7149 ( .A1(n6901), .A2(n6895), .ZN(n6896) );
  AND2_X1 U7150 ( .A1(n6792), .A2(n7796), .ZN(n6793) );
  OR2_X1 U7151 ( .A1(n5572), .A2(n6793), .ZN(n6694) );
  NAND2_X1 U7152 ( .A1(n8882), .A2(n7018), .ZN(n5573) );
  AND2_X1 U7153 ( .A1(n6694), .A2(n5573), .ZN(n5575) );
  AND2_X1 U7154 ( .A1(n5573), .A2(n7801), .ZN(n5574) );
  AND2_X1 U7155 ( .A1(n9253), .A2(n6949), .ZN(n5576) );
  NAND2_X1 U7156 ( .A1(n7634), .A2(n7632), .ZN(n9249) );
  INV_X1 U7157 ( .A(n7141), .ZN(n5577) );
  NAND2_X1 U7158 ( .A1(n5577), .A2(n4982), .ZN(n5579) );
  NAND2_X1 U7159 ( .A1(n7151), .A2(n9252), .ZN(n5578) );
  NAND2_X1 U7160 ( .A1(n7667), .A2(n7635), .ZN(n7207) );
  INV_X1 U7161 ( .A(n7143), .ZN(n8880) );
  INV_X1 U7162 ( .A(n7276), .ZN(n9350) );
  OAI21_X1 U7163 ( .B1(n9196), .B2(n8877), .A(n9098), .ZN(n5581) );
  NAND2_X1 U7164 ( .A1(n5581), .A2(n4974), .ZN(n9083) );
  INV_X1 U7165 ( .A(n9103), .ZN(n8876) );
  AOI21_X1 U7166 ( .B1(n9083), .B2(n9084), .A(n5582), .ZN(n9070) );
  NOR2_X1 U7167 ( .A1(n9186), .A2(n9063), .ZN(n5583) );
  INV_X1 U7168 ( .A(n9074), .ZN(n8875) );
  NAND2_X1 U7169 ( .A1(n9176), .A2(n9062), .ZN(n5586) );
  NOR2_X1 U7170 ( .A1(n9176), .A2(n9062), .ZN(n5585) );
  NAND2_X1 U7171 ( .A1(n9028), .A2(n9046), .ZN(n5587) );
  NAND2_X1 U7172 ( .A1(n9022), .A2(n5587), .ZN(n5589) );
  INV_X1 U7173 ( .A(n9046), .ZN(n9016) );
  NAND2_X1 U7174 ( .A1(n9169), .A2(n9016), .ZN(n5588) );
  NAND2_X1 U7175 ( .A1(n5589), .A2(n5588), .ZN(n9007) );
  NAND2_X1 U7176 ( .A1(n9007), .A2(n9006), .ZN(n5590) );
  INV_X1 U7177 ( .A(n9165), .ZN(n9012) );
  NAND2_X1 U7178 ( .A1(n8997), .A2(n8984), .ZN(n5591) );
  NAND2_X1 U7179 ( .A1(n8944), .A2(n8786), .ZN(n5592) );
  NAND2_X1 U7180 ( .A1(n8939), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7181 ( .A1(n9139), .A2(n8959), .ZN(n5593) );
  NAND2_X1 U7182 ( .A1(n5594), .A2(n5593), .ZN(n8927) );
  NAND2_X1 U7183 ( .A1(n5596), .A2(n7816), .ZN(n5597) );
  NAND2_X1 U7184 ( .A1(n8902), .A2(n5597), .ZN(n9133) );
  NAND2_X1 U7185 ( .A1(n7838), .A2(n5543), .ZN(n5600) );
  OR2_X1 U7186 ( .A1(n5600), .A2(n5611), .ZN(n6349) );
  NAND2_X1 U7187 ( .A1(n5600), .A2(n5611), .ZN(n5615) );
  NAND2_X1 U7188 ( .A1(n6349), .A2(n8756), .ZN(n6453) );
  INV_X1 U7189 ( .A(n6453), .ZN(n5601) );
  NOR2_X1 U7190 ( .A1(n6603), .A2(n5598), .ZN(n9504) );
  NOR2_X1 U7191 ( .A1(n8903), .A2(n9110), .ZN(n5605) );
  INV_X1 U7192 ( .A(n5610), .ZN(n5609) );
  INV_X4 U7193 ( .A(n5668), .ZN(n8758) );
  OR2_X1 U7194 ( .A1(n7838), .A2(n6602), .ZN(n5612) );
  AOI22_X1 U7195 ( .A1(n9156), .A2(n8758), .B1(n8753), .B2(n9000), .ZN(n8735)
         );
  OAI22_X1 U7196 ( .A1(n9111), .A2(n5790), .B1(n9087), .B2(n5761), .ZN(n8861)
         );
  OAI22_X1 U7197 ( .A1(n9345), .A2(n5790), .B1(n9102), .B2(n5761), .ZN(n7284)
         );
  NAND2_X1 U7198 ( .A1(n5613), .A2(n8758), .ZN(n5614) );
  INV_X1 U7199 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U7200 ( .A1(n6605), .A2(n8759), .ZN(n5617) );
  OAI21_X1 U7201 ( .B1(n9377), .B2(n5610), .A(n5617), .ZN(n5618) );
  NAND2_X1 U7202 ( .A1(n5619), .A2(n8753), .ZN(n5622) );
  INV_X1 U7203 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9370) );
  NOR2_X1 U7204 ( .A1(n5610), .A2(n9370), .ZN(n5620) );
  AOI21_X1 U7205 ( .B1(n8758), .B2(n6605), .A(n5620), .ZN(n5621) );
  NAND2_X1 U7206 ( .A1(n5622), .A2(n5621), .ZN(n6157) );
  NAND2_X1 U7207 ( .A1(n6159), .A2(n8756), .ZN(n5623) );
  OAI21_X1 U7208 ( .B1(n6159), .B2(n6157), .A(n5623), .ZN(n5626) );
  NAND2_X1 U7209 ( .A1(n5613), .A2(n8753), .ZN(n5625) );
  NAND2_X1 U7210 ( .A1(n5162), .A2(n8758), .ZN(n5624) );
  NAND2_X1 U7211 ( .A1(n5625), .A2(n5624), .ZN(n6333) );
  NAND2_X1 U7212 ( .A1(n6332), .A2(n6333), .ZN(n5630) );
  INV_X1 U7213 ( .A(n5626), .ZN(n5629) );
  INV_X1 U7214 ( .A(n5627), .ZN(n5628) );
  NAND2_X1 U7215 ( .A1(n5629), .A2(n5628), .ZN(n6331) );
  NAND2_X1 U7216 ( .A1(n7869), .A2(n8759), .ZN(n5633) );
  NAND2_X1 U7217 ( .A1(n5631), .A2(n8758), .ZN(n5632) );
  NAND2_X1 U7218 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  AND2_X1 U7219 ( .A1(n8758), .A2(n7869), .ZN(n5635) );
  XNOR2_X1 U7220 ( .A(n5636), .B(n5637), .ZN(n7864) );
  INV_X1 U7221 ( .A(n5636), .ZN(n5638) );
  NAND2_X1 U7222 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U7223 ( .A1(n7863), .A2(n5639), .ZN(n6406) );
  INV_X2 U7224 ( .A(n8759), .ZN(n5788) );
  OAI22_X1 U7225 ( .A1(n7867), .A2(n5790), .B1(n6535), .B2(n5788), .ZN(n5640)
         );
  XNOR2_X1 U7226 ( .A(n5640), .B(n5777), .ZN(n5645) );
  OR2_X1 U7227 ( .A1(n7867), .A2(n5761), .ZN(n5642) );
  NAND2_X1 U7228 ( .A1(n8758), .A2(n5190), .ZN(n5641) );
  NAND2_X1 U7229 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  XNOR2_X1 U7230 ( .A(n5645), .B(n5643), .ZN(n6405) );
  INV_X1 U7231 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7232 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  XNOR2_X1 U7233 ( .A(n5647), .B(n8756), .ZN(n5652) );
  OR2_X1 U7234 ( .A1(n6556), .A2(n5761), .ZN(n5649) );
  NAND2_X1 U7235 ( .A1(n8758), .A2(n6737), .ZN(n5648) );
  NAND2_X1 U7236 ( .A1(n5649), .A2(n5648), .ZN(n5651) );
  XNOR2_X1 U7237 ( .A(n5652), .B(n5651), .ZN(n6525) );
  NAND2_X1 U7238 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  OR2_X1 U7239 ( .A1(n6905), .A2(n5761), .ZN(n5655) );
  NAND2_X1 U7240 ( .A1(n8758), .A2(n5247), .ZN(n5654) );
  OAI22_X1 U7241 ( .A1(n7853), .A2(n5790), .B1(n6914), .B2(n5788), .ZN(n5657)
         );
  XNOR2_X1 U7242 ( .A(n5657), .B(n5777), .ZN(n6871) );
  OR2_X1 U7243 ( .A1(n7853), .A2(n5761), .ZN(n5659) );
  NAND2_X1 U7244 ( .A1(n8758), .A2(n5527), .ZN(n5658) );
  AND2_X1 U7245 ( .A1(n5659), .A2(n5658), .ZN(n5674) );
  AOI22_X1 U7246 ( .A1(n6678), .A2(n6676), .B1(n6871), .B2(n5674), .ZN(n6935)
         );
  OAI22_X1 U7247 ( .A1(n6801), .A2(n5790), .B1(n9539), .B2(n5788), .ZN(n5660)
         );
  XNOR2_X1 U7248 ( .A(n5660), .B(n5777), .ZN(n7006) );
  OR2_X1 U7249 ( .A1(n6801), .A2(n5761), .ZN(n5662) );
  NAND2_X1 U7250 ( .A1(n8758), .A2(n7018), .ZN(n5661) );
  NAND2_X1 U7251 ( .A1(n9253), .A2(n8753), .ZN(n5664) );
  NAND2_X1 U7252 ( .A1(n8758), .A2(n6949), .ZN(n5663) );
  AND2_X1 U7253 ( .A1(n5664), .A2(n5663), .ZN(n5687) );
  NAND2_X1 U7254 ( .A1(n9253), .A2(n8758), .ZN(n5665) );
  NAND2_X1 U7255 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  XNOR2_X1 U7256 ( .A(n5667), .B(n5777), .ZN(n6943) );
  OAI22_X1 U7257 ( .A1(n6904), .A2(n5668), .B1(n7857), .B2(n5788), .ZN(n5669)
         );
  XNOR2_X1 U7258 ( .A(n5669), .B(n5777), .ZN(n5678) );
  OR2_X1 U7259 ( .A1(n6904), .A2(n5761), .ZN(n5671) );
  NAND2_X1 U7260 ( .A1(n8758), .A2(n6981), .ZN(n5670) );
  AND2_X1 U7261 ( .A1(n5671), .A2(n5670), .ZN(n5679) );
  NAND2_X1 U7262 ( .A1(n5678), .A2(n5679), .ZN(n7847) );
  INV_X1 U7263 ( .A(n6871), .ZN(n5677) );
  NAND2_X1 U7264 ( .A1(n5673), .A2(n5674), .ZN(n5676) );
  INV_X1 U7265 ( .A(n5673), .ZN(n5675) );
  INV_X1 U7266 ( .A(n5674), .ZN(n6870) );
  AOI22_X1 U7267 ( .A1(n5677), .A2(n5676), .B1(n5675), .B2(n6870), .ZN(n7849)
         );
  INV_X1 U7268 ( .A(n5678), .ZN(n5681) );
  INV_X1 U7269 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7270 ( .A1(n5681), .A2(n5680), .ZN(n7848) );
  NAND2_X1 U7271 ( .A1(n7849), .A2(n7848), .ZN(n6936) );
  NAND2_X1 U7272 ( .A1(n5683), .A2(n4431), .ZN(n5684) );
  NAND2_X1 U7273 ( .A1(n5685), .A2(n5684), .ZN(n5691) );
  INV_X1 U7274 ( .A(n7006), .ZN(n6939) );
  INV_X1 U7275 ( .A(n5686), .ZN(n6940) );
  INV_X1 U7276 ( .A(n5687), .ZN(n6942) );
  OAI21_X1 U7277 ( .B1(n6939), .B2(n6940), .A(n6942), .ZN(n5689) );
  NOR2_X1 U7278 ( .A1(n6940), .A2(n6942), .ZN(n5688) );
  AOI22_X1 U7279 ( .A1(n5689), .A2(n6943), .B1(n7006), .B2(n5688), .ZN(n5690)
         );
  OAI22_X1 U7280 ( .A1(n7144), .A2(n5790), .B1(n9274), .B2(n5788), .ZN(n5692)
         );
  XNOR2_X1 U7281 ( .A(n5692), .B(n5777), .ZN(n6640) );
  OR2_X1 U7282 ( .A1(n7144), .A2(n5761), .ZN(n5694) );
  NAND2_X1 U7283 ( .A1(n9263), .A2(n8758), .ZN(n5693) );
  AND2_X1 U7284 ( .A1(n5694), .A2(n5693), .ZN(n6639) );
  AND2_X1 U7285 ( .A1(n6640), .A2(n6639), .ZN(n5695) );
  OAI22_X1 U7286 ( .A1(n6642), .A2(n5695), .B1(n6640), .B2(n6639), .ZN(n6783)
         );
  NAND2_X1 U7287 ( .A1(n7151), .A2(n8759), .ZN(n5697) );
  NAND2_X1 U7288 ( .A1(n9252), .A2(n8758), .ZN(n5696) );
  NAND2_X1 U7289 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  XNOR2_X1 U7290 ( .A(n5698), .B(n5777), .ZN(n5701) );
  NAND2_X1 U7291 ( .A1(n7151), .A2(n8758), .ZN(n5700) );
  NAND2_X1 U7292 ( .A1(n9252), .A2(n8753), .ZN(n5699) );
  NAND2_X1 U7293 ( .A1(n5700), .A2(n5699), .ZN(n5702) );
  XNOR2_X1 U7294 ( .A(n5701), .B(n5702), .ZN(n6782) );
  NAND2_X1 U7295 ( .A1(n6783), .A2(n6782), .ZN(n5705) );
  INV_X1 U7296 ( .A(n5701), .ZN(n5703) );
  NAND2_X1 U7297 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7298 ( .A1(n5705), .A2(n5704), .ZN(n7118) );
  NAND2_X1 U7299 ( .A1(n7215), .A2(n8759), .ZN(n5707) );
  OR2_X1 U7300 ( .A1(n7143), .A2(n5790), .ZN(n5706) );
  NAND2_X1 U7301 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  XNOR2_X1 U7302 ( .A(n5708), .B(n5777), .ZN(n5711) );
  NAND2_X1 U7303 ( .A1(n7215), .A2(n8758), .ZN(n5710) );
  OR2_X1 U7304 ( .A1(n7143), .A2(n5761), .ZN(n5709) );
  AND2_X1 U7305 ( .A1(n5710), .A2(n5709), .ZN(n5712) );
  NAND2_X1 U7306 ( .A1(n5711), .A2(n5712), .ZN(n5717) );
  INV_X1 U7307 ( .A(n5711), .ZN(n5714) );
  INV_X1 U7308 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7309 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U7310 ( .A1(n5717), .A2(n5715), .ZN(n7122) );
  NAND2_X1 U7311 ( .A1(n7276), .A2(n8759), .ZN(n5719) );
  NAND2_X1 U7312 ( .A1(n8879), .A2(n8758), .ZN(n5718) );
  NAND2_X1 U7313 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  XNOR2_X1 U7314 ( .A(n5720), .B(n8756), .ZN(n5726) );
  INV_X1 U7315 ( .A(n5726), .ZN(n5724) );
  NAND2_X1 U7316 ( .A1(n7276), .A2(n8758), .ZN(n5722) );
  NAND2_X1 U7317 ( .A1(n8879), .A2(n8753), .ZN(n5721) );
  NAND2_X1 U7318 ( .A1(n5722), .A2(n5721), .ZN(n5725) );
  INV_X1 U7319 ( .A(n5725), .ZN(n5723) );
  NAND2_X1 U7320 ( .A1(n5724), .A2(n5723), .ZN(n7130) );
  AND2_X1 U7321 ( .A1(n5726), .A2(n5725), .ZN(n7131) );
  NAND2_X1 U7322 ( .A1(n7583), .A2(n8759), .ZN(n5728) );
  NAND2_X1 U7323 ( .A1(n8878), .A2(n8758), .ZN(n5727) );
  NAND2_X1 U7324 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  XNOR2_X1 U7325 ( .A(n5729), .B(n5777), .ZN(n5730) );
  OAI22_X1 U7326 ( .A1(n9111), .A2(n5788), .B1(n9087), .B2(n5790), .ZN(n5731)
         );
  XOR2_X1 U7327 ( .A(n8756), .B(n5731), .Z(n5732) );
  OAI22_X1 U7328 ( .A1(n9095), .A2(n5790), .B1(n9103), .B2(n5761), .ZN(n5737)
         );
  NAND2_X1 U7329 ( .A1(n9191), .A2(n8759), .ZN(n5735) );
  OR2_X1 U7330 ( .A1(n9103), .A2(n5790), .ZN(n5734) );
  NAND2_X1 U7331 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  XNOR2_X1 U7332 ( .A(n5736), .B(n8756), .ZN(n5738) );
  XOR2_X1 U7333 ( .A(n5737), .B(n5738), .Z(n8792) );
  OAI22_X1 U7334 ( .A1(n9079), .A2(n5790), .B1(n9088), .B2(n5761), .ZN(n5742)
         );
  NAND2_X1 U7335 ( .A1(n9186), .A2(n8759), .ZN(n5740) );
  NAND2_X1 U7336 ( .A1(n9063), .A2(n8758), .ZN(n5739) );
  NAND2_X1 U7337 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  XNOR2_X1 U7338 ( .A(n5741), .B(n8756), .ZN(n5743) );
  XOR2_X1 U7339 ( .A(n5742), .B(n5743), .Z(n8800) );
  OR2_X1 U7340 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  NAND2_X1 U7341 ( .A1(n8798), .A2(n5744), .ZN(n5747) );
  AOI22_X1 U7342 ( .A1(n9179), .A2(n8759), .B1(n8758), .B2(n8875), .ZN(n5745)
         );
  XNOR2_X1 U7343 ( .A(n5745), .B(n8756), .ZN(n5746) );
  OAI22_X1 U7344 ( .A1(n4573), .A2(n5790), .B1(n9074), .B2(n5761), .ZN(n8837)
         );
  OAI22_X1 U7345 ( .A1(n9051), .A2(n5790), .B1(n5748), .B2(n5761), .ZN(n5752)
         );
  NAND2_X1 U7346 ( .A1(n9176), .A2(n8759), .ZN(n5750) );
  NAND2_X1 U7347 ( .A1(n9062), .A2(n8758), .ZN(n5749) );
  NAND2_X1 U7348 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  XNOR2_X1 U7349 ( .A(n5751), .B(n8756), .ZN(n5753) );
  XOR2_X1 U7350 ( .A(n5752), .B(n5753), .Z(n8746) );
  OR2_X1 U7351 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  OAI22_X1 U7352 ( .A1(n9028), .A2(n5788), .B1(n9046), .B2(n5790), .ZN(n5755)
         );
  XNOR2_X1 U7353 ( .A(n5755), .B(n8756), .ZN(n5757) );
  OAI22_X1 U7354 ( .A1(n9028), .A2(n5790), .B1(n9046), .B2(n5761), .ZN(n5756)
         );
  NAND2_X1 U7355 ( .A1(n5757), .A2(n5756), .ZN(n8816) );
  NAND2_X1 U7356 ( .A1(n9165), .A2(n8759), .ZN(n5759) );
  OR2_X1 U7357 ( .A1(n9029), .A2(n5790), .ZN(n5758) );
  NAND2_X1 U7358 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  XNOR2_X1 U7359 ( .A(n5760), .B(n8756), .ZN(n5763) );
  OAI22_X1 U7360 ( .A1(n9012), .A2(n5790), .B1(n9029), .B2(n5761), .ZN(n5762)
         );
  XNOR2_X1 U7361 ( .A(n5763), .B(n5762), .ZN(n8774) );
  INV_X1 U7362 ( .A(n8984), .ZN(n9017) );
  AOI22_X1 U7363 ( .A1(n9159), .A2(n8758), .B1(n8753), .B2(n9017), .ZN(n5766)
         );
  AND2_X1 U7364 ( .A1(n5765), .A2(n5766), .ZN(n8824) );
  OAI22_X1 U7365 ( .A1(n8997), .A2(n5788), .B1(n8984), .B2(n5790), .ZN(n5764)
         );
  XOR2_X1 U7366 ( .A(n8756), .B(n5764), .Z(n8826) );
  INV_X1 U7367 ( .A(n5765), .ZN(n5768) );
  NAND2_X1 U7368 ( .A1(n9156), .A2(n8759), .ZN(n5770) );
  NAND2_X1 U7369 ( .A1(n9000), .A2(n8758), .ZN(n5769) );
  NAND2_X1 U7370 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  XNOR2_X1 U7371 ( .A(n5771), .B(n8756), .ZN(n5775) );
  INV_X1 U7372 ( .A(n5775), .ZN(n5772) );
  NAND2_X1 U7373 ( .A1(n5774), .A2(n5772), .ZN(n5773) );
  NOR2_X1 U7374 ( .A1(n5776), .A2(n5773), .ZN(n8732) );
  INV_X1 U7375 ( .A(n5774), .ZN(n8825) );
  OAI22_X1 U7376 ( .A1(n5779), .A2(n5788), .B1(n8738), .B2(n5790), .ZN(n5778)
         );
  XNOR2_X1 U7377 ( .A(n5778), .B(n5777), .ZN(n5783) );
  OR2_X1 U7378 ( .A1(n5779), .A2(n5790), .ZN(n5781) );
  NAND2_X1 U7379 ( .A1(n4868), .A2(n8753), .ZN(n5780) );
  NAND2_X1 U7380 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  OAI21_X1 U7381 ( .B1(n5783), .B2(n5782), .A(n5784), .ZN(n8808) );
  NAND2_X1 U7382 ( .A1(n9144), .A2(n8759), .ZN(n5786) );
  NAND2_X1 U7383 ( .A1(n8969), .A2(n8758), .ZN(n5785) );
  NAND2_X1 U7384 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  XNOR2_X1 U7385 ( .A(n5787), .B(n8756), .ZN(n5795) );
  AOI22_X1 U7386 ( .A1(n9144), .A2(n8758), .B1(n8753), .B2(n8969), .ZN(n5793)
         );
  XNOR2_X1 U7387 ( .A(n5795), .B(n5793), .ZN(n8782) );
  OAI22_X1 U7388 ( .A1(n8944), .A2(n5788), .B1(n8786), .B2(n5790), .ZN(n5789)
         );
  XNOR2_X1 U7389 ( .A(n5789), .B(n8756), .ZN(n5798) );
  OR2_X1 U7390 ( .A1(n8944), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U7391 ( .A1(n8959), .A2(n8753), .ZN(n5791) );
  NAND2_X1 U7392 ( .A1(n5792), .A2(n5791), .ZN(n5797) );
  XNOR2_X1 U7393 ( .A(n5798), .B(n5797), .ZN(n8845) );
  INV_X1 U7394 ( .A(n5793), .ZN(n5794) );
  NOR2_X1 U7395 ( .A1(n5795), .A2(n5794), .ZN(n8846) );
  NOR2_X1 U7396 ( .A1(n8845), .A2(n8846), .ZN(n5796) );
  NAND2_X1 U7397 ( .A1(n5798), .A2(n5797), .ZN(n5807) );
  NAND2_X1 U7398 ( .A1(n9134), .A2(n8759), .ZN(n5800) );
  NAND2_X1 U7399 ( .A1(n8947), .A2(n8758), .ZN(n5799) );
  NAND2_X1 U7400 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  XNOR2_X1 U7401 ( .A(n5801), .B(n8756), .ZN(n5805) );
  NAND2_X1 U7402 ( .A1(n9134), .A2(n8758), .ZN(n5803) );
  NAND2_X1 U7403 ( .A1(n8947), .A2(n8753), .ZN(n5802) );
  NAND2_X1 U7404 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  NOR2_X1 U7405 ( .A1(n5805), .A2(n5804), .ZN(n8767) );
  AOI21_X1 U7406 ( .B1(n8848), .B2(n5807), .A(n5806), .ZN(n5812) );
  INV_X1 U7407 ( .A(n5806), .ZN(n5809) );
  INV_X1 U7408 ( .A(n5807), .ZN(n5808) );
  NOR2_X1 U7409 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NOR2_X1 U7410 ( .A1(n6461), .A2(n5811), .ZN(n5816) );
  OAI21_X1 U7411 ( .B1(n5812), .B2(n8762), .A(n8849), .ZN(n5829) );
  NAND2_X1 U7412 ( .A1(n9504), .A2(n5822), .ZN(n5813) );
  NOR2_X1 U7413 ( .A1(n9104), .A2(n6602), .ZN(n5814) );
  AND3_X1 U7414 ( .A1(n5815), .A2(n5610), .A3(n6811), .ZN(n5817) );
  INV_X1 U7415 ( .A(n5816), .ZN(n5819) );
  NAND2_X1 U7416 ( .A1(n9546), .A2(n5819), .ZN(n6154) );
  NAND2_X1 U7417 ( .A1(n5817), .A2(n6154), .ZN(n5818) );
  NAND2_X1 U7418 ( .A1(n5818), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5821) );
  AND2_X1 U7419 ( .A1(n5819), .A2(n7835), .ZN(n5820) );
  NAND2_X1 U7420 ( .A1(n9504), .A2(n5820), .ZN(n6156) );
  NOR2_X1 U7421 ( .A1(n8929), .A2(n8812), .ZN(n5825) );
  NOR2_X1 U7422 ( .A1(n6349), .A2(n5524), .ZN(n5823) );
  NAND2_X1 U7423 ( .A1(n5823), .A2(n5822), .ZN(n8852) );
  OAI22_X1 U7424 ( .A1(n8786), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10090), .ZN(n5824) );
  AOI211_X1 U7425 ( .C1(n8934), .C2(n8839), .A(n5825), .B(n5824), .ZN(n5826)
         );
  OAI21_X1 U7426 ( .B1(n4743), .B2(n8859), .A(n5826), .ZN(n5827) );
  INV_X1 U7427 ( .A(n5827), .ZN(n5828) );
  NAND2_X1 U7428 ( .A1(n5829), .A2(n5828), .ZN(P1_U3212) );
  INV_X1 U7429 ( .A(n6811), .ZN(n5863) );
  NAND2_X1 U7430 ( .A1(n5881), .A2(n5832), .ZN(n5893) );
  INV_X1 U7431 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5836) );
  NOR2_X1 U7432 ( .A1(n5844), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7433 ( .A1(n6076), .A2(n5840), .ZN(n5939) );
  INV_X1 U7434 ( .A(n5904), .ZN(n5931) );
  INV_X1 U7435 ( .A(n5844), .ZN(n5846) );
  NAND4_X1 U7436 ( .A1(n5846), .A2(n5845), .A3(n5937), .A4(n5860), .ZN(n5852)
         );
  NOR2_X1 U7437 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5850) );
  NOR2_X1 U7438 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U7439 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5848) );
  NOR2_X1 U7440 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5847) );
  NAND4_X1 U7441 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n5851)
         );
  NOR2_X2 U7442 ( .A1(n5852), .A2(n5851), .ZN(n5856) );
  AND2_X2 U7443 ( .A1(n5856), .A2(n5853), .ZN(n5906) );
  NAND2_X1 U7444 ( .A1(n5931), .A2(n5906), .ZN(n5854) );
  NAND2_X1 U7445 ( .A1(n5854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7446 ( .A1(n5931), .A2(n5856), .ZN(n5857) );
  NAND2_X1 U7447 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7448 ( .A1(n6121), .A2(n7174), .ZN(n5859) );
  INV_X1 U7449 ( .A(n6226), .ZN(n5862) );
  XNOR2_X1 U7450 ( .A(n5861), .B(n5860), .ZN(n6197) );
  OR2_X1 U7451 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NAND2_X1 U7452 ( .A1(n5865), .A2(n5974), .ZN(n9374) );
  OR2_X1 U7453 ( .A1(n9374), .A2(n5866), .ZN(n5867) );
  NAND2_X1 U7454 ( .A1(n5867), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U7455 ( .A1(n7555), .A2(P1_U3084), .ZN(n8103) );
  OAI222_X1 U7456 ( .A1(n8103), .A2(n5870), .B1(n4396), .B2(n6089), .C1(
        P1_U3084), .C2(n5869), .ZN(P1_U3352) );
  OAI222_X1 U7457 ( .A1(n8103), .A2(n5871), .B1(n4396), .B2(n6106), .C1(
        P1_U3084), .C2(n9407), .ZN(P1_U3351) );
  OAI222_X1 U7458 ( .A1(n8103), .A2(n5872), .B1(n4396), .B2(n6309), .C1(
        P1_U3084), .C2(n9417), .ZN(P1_U3349) );
  INV_X1 U7459 ( .A(n8103), .ZN(n9221) );
  OAI222_X1 U7460 ( .A1(n8108), .A2(n9921), .B1(n4396), .B2(n6204), .C1(
        P1_U3084), .C2(n5998), .ZN(P1_U3350) );
  NOR2_X1 U7461 ( .A1(n7555), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8725) );
  INV_X2 U7462 ( .A(n8725), .ZN(n8727) );
  INV_X1 U7463 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6090) );
  AND2_X1 U7464 ( .A1(n7555), .A2(P2_U3152), .ZN(n7330) );
  INV_X2 U7465 ( .A(n7330), .ZN(n7895) );
  INV_X1 U7466 ( .A(n9229), .ZN(n6247) );
  OAI222_X1 U7467 ( .A1(n8727), .A2(n6090), .B1(n7895), .B2(n6089), .C1(
        P2_U3152), .C2(n6247), .ZN(P2_U3357) );
  INV_X1 U7468 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5876) );
  NOR2_X1 U7469 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5874) );
  NAND2_X1 U7470 ( .A1(n5876), .A2(n5874), .ZN(n5878) );
  NAND2_X1 U7471 ( .A1(n5878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U7472 ( .A(n5873), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6244) );
  INV_X1 U7473 ( .A(n6244), .ZN(n6294) );
  OAI222_X1 U7474 ( .A1(n8727), .A2(n6205), .B1(n7895), .B2(n6204), .C1(
        P2_U3152), .C2(n6294), .ZN(P2_U3355) );
  INV_X1 U7475 ( .A(n5874), .ZN(n5875) );
  NAND2_X1 U7476 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5875), .ZN(n5877) );
  MUX2_X1 U7477 ( .A(n5877), .B(P2_IR_REG_31__SCAN_IN), .S(n5876), .Z(n5879)
         );
  INV_X1 U7478 ( .A(n9240), .ZN(n6109) );
  OAI222_X1 U7479 ( .A1(n8727), .A2(n6105), .B1(n7895), .B2(n6106), .C1(
        P2_U3152), .C2(n6109), .ZN(P2_U3356) );
  OR2_X1 U7480 ( .A1(n5882), .A2(n8722), .ZN(n5883) );
  XNOR2_X1 U7481 ( .A(n5880), .B(n5883), .ZN(n6312) );
  OAI222_X1 U7482 ( .A1(n8727), .A2(n6311), .B1(n7895), .B2(n6309), .C1(
        P2_U3152), .C2(n6312), .ZN(P2_U3354) );
  OAI222_X1 U7483 ( .A1(n8103), .A2(n5884), .B1(n4396), .B2(n6365), .C1(
        P1_U3084), .C2(n6030), .ZN(P1_U3348) );
  NAND2_X1 U7484 ( .A1(n5882), .A2(n5880), .ZN(n5886) );
  NAND2_X1 U7485 ( .A1(n5886), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5885) );
  XNOR2_X1 U7486 ( .A(n5885), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6241) );
  INV_X1 U7487 ( .A(n6241), .ZN(n6369) );
  OAI222_X1 U7488 ( .A1(n8727), .A2(n6366), .B1(n7895), .B2(n6365), .C1(
        P2_U3152), .C2(n6369), .ZN(P2_U3353) );
  NAND2_X1 U7489 ( .A1(n5890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7490 ( .A(n5887), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6275) );
  INV_X1 U7491 ( .A(n6275), .ZN(n6422) );
  OAI222_X1 U7492 ( .A1(n8727), .A2(n6419), .B1(n7895), .B2(n6418), .C1(
        P2_U3152), .C2(n6422), .ZN(P2_U3352) );
  OAI222_X1 U7493 ( .A1(n8103), .A2(n5888), .B1(n4396), .B2(n6418), .C1(
        P1_U3084), .C2(n6039), .ZN(P1_U3347) );
  OAI222_X1 U7494 ( .A1(n8103), .A2(n5889), .B1(n4396), .B2(n6429), .C1(
        P1_U3084), .C2(n6061), .ZN(P1_U3346) );
  OAI21_X1 U7495 ( .B1(n5890), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U7496 ( .A(n5891), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6428) );
  INV_X1 U7497 ( .A(n6428), .ZN(n8286) );
  OAI222_X1 U7498 ( .A1(n8727), .A2(n5892), .B1(n7895), .B2(n6429), .C1(
        P2_U3152), .C2(n8286), .ZN(P2_U3351) );
  NAND2_X1 U7499 ( .A1(n5893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5894) );
  MUX2_X1 U7500 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5894), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5896) );
  NAND2_X1 U7501 ( .A1(n5896), .A2(n5895), .ZN(n6389) );
  OAI222_X1 U7502 ( .A1(n8727), .A2(n10084), .B1(n7895), .B2(n6502), .C1(
        P2_U3152), .C2(n6389), .ZN(P2_U3350) );
  OAI222_X1 U7503 ( .A1(n8108), .A2(n5897), .B1(n4396), .B2(n6502), .C1(
        P1_U3084), .C2(n6165), .ZN(P1_U3345) );
  OAI222_X1 U7504 ( .A1(n4396), .A2(n6569), .B1(n5899), .B2(P1_U3084), .C1(
        n5898), .C2(n8108), .ZN(P1_U3344) );
  INV_X1 U7505 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5901) );
  INV_X1 U7506 ( .A(n6340), .ZN(n5900) );
  AOI22_X1 U7507 ( .A1(n9515), .A2(n5901), .B1(n7835), .B2(n5900), .ZN(
        P1_U3441) );
  NAND2_X1 U7508 ( .A1(n5895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5902) );
  XNOR2_X1 U7509 ( .A(n5902), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6570) );
  INV_X1 U7510 ( .A(n6570), .ZN(n8298) );
  OAI222_X1 U7511 ( .A1(n8727), .A2(n5903), .B1(n7895), .B2(n6569), .C1(n8298), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7512 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5916) );
  INV_X1 U7513 ( .A(n5910), .ZN(n5908) );
  NAND2_X1 U7514 ( .A1(n5908), .A2(n5907), .ZN(n8723) );
  NAND2_X1 U7515 ( .A1(n7490), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5914) );
  INV_X2 U7516 ( .A(n7448), .ZN(n7459) );
  NAND2_X1 U7517 ( .A1(n7459), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7518 ( .A1(n7488), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5912) );
  NAND3_X1 U7519 ( .A1(n5914), .A2(n5913), .A3(n5912), .ZN(n8398) );
  NAND2_X1 U7520 ( .A1(n8398), .A2(P2_U3966), .ZN(n5915) );
  OAI21_X1 U7521 ( .B1(n5916), .B2(P2_U3966), .A(n5915), .ZN(P2_U3583) );
  INV_X1 U7522 ( .A(n6584), .ZN(n5925) );
  INV_X1 U7523 ( .A(n9444), .ZN(n6178) );
  OAI222_X1 U7524 ( .A1(n4396), .A2(n5925), .B1(n6178), .B2(P1_U3084), .C1(
        n5917), .C2(n8108), .ZN(P1_U3343) );
  INV_X1 U7525 ( .A(n6655), .ZN(n5922) );
  NAND2_X1 U7526 ( .A1(n5918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U7527 ( .A(n5919), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6656) );
  AOI22_X1 U7528 ( .A1(n6656), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8725), .ZN(n5920) );
  OAI21_X1 U7529 ( .B1(n5922), .B2(n7895), .A(n5920), .ZN(P2_U3347) );
  AOI22_X1 U7530 ( .A1(n9457), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9221), .ZN(n5921) );
  OAI21_X1 U7531 ( .B1(n5922), .B2(n4396), .A(n5921), .ZN(P1_U3342) );
  OR2_X1 U7532 ( .A1(n5923), .A2(n8722), .ZN(n5924) );
  XNOR2_X1 U7533 ( .A(n5924), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6585) );
  INV_X1 U7534 ( .A(n6585), .ZN(n8311) );
  OAI222_X1 U7535 ( .A1(n8727), .A2(n5926), .B1(n7895), .B2(n5925), .C1(n8311), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  OR2_X1 U7536 ( .A1(n6197), .A2(P2_U3152), .ZN(n8100) );
  INV_X1 U7537 ( .A(n8100), .ZN(n5936) );
  XNOR2_X2 U7538 ( .A(n5928), .B(n5927), .ZN(n6142) );
  NAND2_X1 U7539 ( .A1(n5932), .A2(n8722), .ZN(n5929) );
  NAND2_X1 U7540 ( .A1(n5931), .A2(n4458), .ZN(n5934) );
  OAI21_X1 U7541 ( .B1(n9681), .B2(n5936), .A(n7369), .ZN(n5942) );
  NAND2_X1 U7542 ( .A1(n5939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  AND2_X1 U7543 ( .A1(n8097), .A2(n6081), .ZN(n6746) );
  NAND2_X1 U7544 ( .A1(n9681), .A2(n6746), .ZN(n5941) );
  NOR2_X1 U7545 ( .A1(n9600), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7546 ( .A(n6952), .ZN(n5945) );
  INV_X1 U7547 ( .A(n6474), .ZN(n6164) );
  OAI222_X1 U7548 ( .A1(n8108), .A2(n5943), .B1(n4396), .B2(n5945), .C1(
        P1_U3084), .C2(n6164), .ZN(P1_U3341) );
  NAND2_X1 U7549 ( .A1(n5904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5944) );
  XNOR2_X1 U7550 ( .A(n5944), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6953) );
  INV_X1 U7551 ( .A(n6953), .ZN(n6497) );
  OAI222_X1 U7552 ( .A1(n8727), .A2(n5946), .B1(n7895), .B2(n5945), .C1(
        P2_U3152), .C2(n6497), .ZN(P2_U3346) );
  INV_X1 U7553 ( .A(n7057), .ZN(n5948) );
  OR2_X1 U7554 ( .A1(n5955), .A2(n8722), .ZN(n5950) );
  XNOR2_X1 U7555 ( .A(n5950), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7058) );
  INV_X1 U7556 ( .A(n7058), .ZN(n6629) );
  OAI222_X1 U7557 ( .A1(n8727), .A2(n10108), .B1(n7895), .B2(n5948), .C1(n6629), .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7558 ( .A(n7094), .ZN(n5952) );
  INV_X1 U7559 ( .A(n9469), .ZN(n6923) );
  OAI222_X1 U7560 ( .A1(n4396), .A2(n5952), .B1(n6923), .B2(P1_U3084), .C1(
        n5947), .C2(n8108), .ZN(P1_U3339) );
  OAI222_X1 U7561 ( .A1(n8108), .A2(n10120), .B1(n4561), .B2(P1_U3084), .C1(
        n4396), .C2(n5948), .ZN(P1_U3340) );
  NAND2_X1 U7562 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U7563 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  XNOR2_X1 U7564 ( .A(n5967), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8322) );
  INV_X1 U7565 ( .A(n8322), .ZN(n6630) );
  OAI222_X1 U7566 ( .A1(n8727), .A2(n5953), .B1(n7895), .B2(n5952), .C1(n6630), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7567 ( .A(n7305), .ZN(n5973) );
  AND2_X1 U7568 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  OR2_X1 U7569 ( .A1(n5956), .A2(n8722), .ZN(n5957) );
  XNOR2_X1 U7570 ( .A(n5957), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8360) );
  AOI22_X1 U7571 ( .A1(n8360), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8725), .ZN(n5958) );
  OAI21_X1 U7572 ( .B1(n5973), .B2(n7895), .A(n5958), .ZN(P2_U3342) );
  INV_X1 U7573 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7574 ( .A1(n5496), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7575 ( .A1(n5193), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7576 ( .A1(n5176), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5959) );
  NAND3_X1 U7577 ( .A1(n5961), .A2(n5960), .A3(n5959), .ZN(n7740) );
  NAND2_X1 U7578 ( .A1(n7740), .A2(n10144), .ZN(n5962) );
  OAI21_X1 U7579 ( .B1(n10144), .B2(n5963), .A(n5962), .ZN(P1_U3586) );
  INV_X1 U7580 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7581 ( .A1(n5619), .A2(n10144), .ZN(n5964) );
  OAI21_X1 U7582 ( .B1(n10144), .B2(n5965), .A(n5964), .ZN(P1_U3555) );
  INV_X1 U7583 ( .A(n7183), .ZN(n5971) );
  NAND2_X1 U7584 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  NAND2_X1 U7585 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  XNOR2_X1 U7586 ( .A(n5969), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8342) );
  INV_X1 U7587 ( .A(n8342), .ZN(n8334) );
  OAI222_X1 U7588 ( .A1(n8727), .A2(n5970), .B1(n7895), .B2(n5971), .C1(
        P2_U3152), .C2(n8334), .ZN(P2_U3343) );
  OAI222_X1 U7589 ( .A1(n8108), .A2(n9934), .B1(n4396), .B2(n5971), .C1(
        P1_U3084), .C2(n7163), .ZN(P1_U3338) );
  INV_X1 U7590 ( .A(n7538), .ZN(n7170) );
  OAI222_X1 U7591 ( .A1(n4396), .A2(n5973), .B1(n7170), .B2(P1_U3084), .C1(
        n5972), .C2(n8108), .ZN(P1_U3337) );
  INV_X1 U7592 ( .A(n5974), .ZN(n9401) );
  INV_X1 U7593 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7594 ( .A1(n9368), .A2(P1_U3084), .ZN(n7260) );
  NOR2_X1 U7595 ( .A1(n9374), .A2(n7260), .ZN(n6004) );
  INV_X1 U7596 ( .A(n6004), .ZN(n5975) );
  NOR2_X2 U7597 ( .A1(n5975), .A2(n7834), .ZN(n9483) );
  INV_X1 U7598 ( .A(n9374), .ZN(n5978) );
  NAND2_X1 U7599 ( .A1(n9368), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5976) );
  NOR2_X1 U7600 ( .A1(n5524), .A2(n5976), .ZN(n5977) );
  XNOR2_X1 U7601 ( .A(n9407), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U7602 ( .A1(n9386), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5980) );
  XNOR2_X1 U7603 ( .A(n9386), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9383) );
  NOR3_X1 U7604 ( .A1(n9370), .A2(n9377), .A3(n9383), .ZN(n9382) );
  INV_X1 U7605 ( .A(n9382), .ZN(n5979) );
  NAND2_X1 U7606 ( .A1(n5980), .A2(n5979), .ZN(n9393) );
  NAND2_X1 U7607 ( .A1(n9394), .A2(n9393), .ZN(n9392) );
  INV_X1 U7608 ( .A(n9407), .ZN(n5995) );
  NAND2_X1 U7609 ( .A1(n5995), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7610 ( .A1(n9392), .A2(n5981), .ZN(n6016) );
  XNOR2_X1 U7611 ( .A(n5998), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7612 ( .A1(n6016), .A2(n6017), .ZN(n6015) );
  INV_X1 U7613 ( .A(n5998), .ZN(n6014) );
  NAND2_X1 U7614 ( .A1(n6014), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7615 ( .A1(n6015), .A2(n5982), .ZN(n9420) );
  INV_X1 U7616 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9559) );
  MUX2_X1 U7617 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9559), .S(n9417), .Z(n9419)
         );
  OR2_X1 U7618 ( .A1(n9420), .A2(n9419), .ZN(n9422) );
  NAND2_X1 U7619 ( .A1(n9417), .A2(n9559), .ZN(n5983) );
  AND2_X1 U7620 ( .A1(n9422), .A2(n5983), .ZN(n5986) );
  OR2_X1 U7621 ( .A1(n6023), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7622 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6023), .ZN(n5984) );
  AND2_X1 U7623 ( .A1(n5985), .A2(n5984), .ZN(n5987) );
  NAND2_X1 U7624 ( .A1(n5986), .A2(n5987), .ZN(n6028) );
  INV_X1 U7625 ( .A(n5986), .ZN(n5989) );
  INV_X1 U7626 ( .A(n5987), .ZN(n5988) );
  NAND2_X1 U7627 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NAND3_X1 U7628 ( .A1(n9496), .A2(n6028), .A3(n5990), .ZN(n5992) );
  AND2_X1 U7629 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6680) );
  INV_X1 U7630 ( .A(n6680), .ZN(n5991) );
  NAND2_X1 U7631 ( .A1(n5992), .A2(n5991), .ZN(n6008) );
  NAND2_X1 U7632 ( .A1(n9386), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5994) );
  INV_X1 U7633 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5993) );
  NAND3_X1 U7634 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n9388), .ZN(n9387) );
  NAND2_X1 U7635 ( .A1(n5994), .A2(n9387), .ZN(n9403) );
  XNOR2_X1 U7636 ( .A(n9407), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U7637 ( .A1(n9403), .A2(n9404), .ZN(n5997) );
  NAND2_X1 U7638 ( .A1(n5995), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7639 ( .A1(n5997), .A2(n5996), .ZN(n6012) );
  INV_X1 U7640 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5999) );
  MUX2_X1 U7641 ( .A(n5999), .B(P1_REG2_REG_3__SCAN_IN), .S(n5998), .Z(n6013)
         );
  NAND2_X1 U7642 ( .A1(n6014), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6000) );
  INV_X1 U7643 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6001) );
  MUX2_X1 U7644 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6001), .S(n9417), .Z(n9413)
         );
  NAND2_X1 U7645 ( .A1(n9417), .A2(n6001), .ZN(n6002) );
  INV_X1 U7646 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6863) );
  MUX2_X1 U7647 ( .A(n6863), .B(P1_REG2_REG_5__SCAN_IN), .S(n6023), .Z(n6003)
         );
  INV_X1 U7648 ( .A(n6024), .ZN(n6006) );
  NAND3_X1 U7649 ( .A1(n9416), .A2(n6003), .A3(n6002), .ZN(n6005) );
  NAND2_X1 U7650 ( .A1(n6004), .A2(n7834), .ZN(n9488) );
  AOI21_X1 U7651 ( .B1(n6006), .B2(n6005), .A(n9488), .ZN(n6007) );
  AOI211_X1 U7652 ( .C1(n9483), .C2(n6023), .A(n6008), .B(n6007), .ZN(n6009)
         );
  OAI21_X1 U7653 ( .B1(n9481), .B2(n6010), .A(n6009), .ZN(P1_U3246) );
  INV_X1 U7654 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10110) );
  OAI211_X1 U7655 ( .C1(n6013), .C2(n6012), .A(n9477), .B(n6011), .ZN(n6021)
         );
  AND2_X1 U7656 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6407) );
  INV_X1 U7657 ( .A(n6407), .ZN(n6020) );
  NAND2_X1 U7658 ( .A1(n9483), .A2(n6014), .ZN(n6019) );
  OAI211_X1 U7659 ( .C1(n6017), .C2(n6016), .A(n9496), .B(n6015), .ZN(n6018)
         );
  AND4_X1 U7660 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n6022)
         );
  OAI21_X1 U7661 ( .B1(n10110), .B2(n9481), .A(n6022), .ZN(P1_U3244) );
  INV_X1 U7662 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6910) );
  NOR2_X1 U7663 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6023), .ZN(n6025) );
  NOR2_X1 U7664 ( .A1(n6025), .A2(n6024), .ZN(n6048) );
  MUX2_X1 U7665 ( .A(n6910), .B(P1_REG2_REG_6__SCAN_IN), .S(n6039), .Z(n6047)
         );
  NAND2_X1 U7666 ( .A1(n6048), .A2(n6047), .ZN(n6046) );
  OAI21_X1 U7667 ( .B1(n6039), .B2(n6910), .A(n6046), .ZN(n6027) );
  INV_X1 U7668 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6803) );
  MUX2_X1 U7669 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6803), .S(n6061), .Z(n6026)
         );
  NOR2_X1 U7670 ( .A1(n6026), .A2(n6027), .ZN(n6060) );
  AOI21_X1 U7671 ( .B1(n6027), .B2(n6026), .A(n6060), .ZN(n6038) );
  INV_X1 U7672 ( .A(n6061), .ZN(n6055) );
  AND2_X1 U7673 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7855) );
  INV_X1 U7674 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6985) );
  MUX2_X1 U7675 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6985), .S(n6061), .Z(n6033)
         );
  INV_X1 U7676 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6031) );
  INV_X1 U7677 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7678 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6041) );
  XOR2_X1 U7679 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6039), .Z(n6042) );
  NOR2_X1 U7680 ( .A1(n6041), .A2(n6042), .ZN(n6040) );
  AOI21_X1 U7681 ( .B1(n6031), .B2(n6039), .A(n6040), .ZN(n6032) );
  NOR2_X1 U7682 ( .A1(n6032), .A2(n6033), .ZN(n6053) );
  AOI21_X1 U7683 ( .B1(n6033), .B2(n6032), .A(n6053), .ZN(n6034) );
  NOR2_X1 U7684 ( .A1(n9381), .A2(n6034), .ZN(n6035) );
  AOI211_X1 U7685 ( .C1(n9483), .C2(n6055), .A(n7855), .B(n6035), .ZN(n6037)
         );
  INV_X1 U7686 ( .A(n9481), .ZN(n9495) );
  NAND2_X1 U7687 ( .A1(n9495), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7688 ( .C1(n6038), .C2(n9488), .A(n6037), .B(n6036), .ZN(P1_U3248) );
  INV_X1 U7689 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6051) );
  INV_X1 U7690 ( .A(n6039), .ZN(n6045) );
  NOR2_X1 U7691 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10002), .ZN(n6875) );
  AOI21_X1 U7692 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6043) );
  NOR2_X1 U7693 ( .A1(n9381), .A2(n6043), .ZN(n6044) );
  AOI211_X1 U7694 ( .C1(n9483), .C2(n6045), .A(n6875), .B(n6044), .ZN(n6050)
         );
  OAI211_X1 U7695 ( .C1(n6048), .C2(n6047), .A(n9477), .B(n6046), .ZN(n6049)
         );
  OAI211_X1 U7696 ( .C1(n6051), .C2(n9481), .A(n6050), .B(n6049), .ZN(P1_U3247) );
  INV_X1 U7697 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6067) );
  NOR2_X1 U7698 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6052), .ZN(n7013) );
  INV_X1 U7699 ( .A(n6053), .ZN(n6054) );
  OAI21_X1 U7700 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6055), .A(n6054), .ZN(
        n6058) );
  INV_X1 U7701 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6056) );
  MUX2_X1 U7702 ( .A(n6056), .B(P1_REG1_REG_8__SCAN_IN), .S(n6180), .Z(n6057)
         );
  NOR2_X1 U7703 ( .A1(n6057), .A2(n6058), .ZN(n6179) );
  AOI211_X1 U7704 ( .C1(n6058), .C2(n6057), .A(n6179), .B(n9381), .ZN(n6059)
         );
  AOI211_X1 U7705 ( .C1(n9483), .C2(n6180), .A(n7013), .B(n6059), .ZN(n6066)
         );
  AOI21_X1 U7706 ( .B1(n6061), .B2(n6803), .A(n6060), .ZN(n6169) );
  INV_X1 U7707 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6062) );
  MUX2_X1 U7708 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6062), .S(n6180), .Z(n6064)
         );
  NAND2_X1 U7709 ( .A1(n6180), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6166) );
  OAI211_X1 U7710 ( .C1(n6180), .C2(P1_REG2_REG_8__SCAN_IN), .A(n6169), .B(
        n6166), .ZN(n6063) );
  OAI211_X1 U7711 ( .C1(n6169), .C2(n6064), .A(n9477), .B(n6063), .ZN(n6065)
         );
  OAI211_X1 U7712 ( .C1(n6067), .C2(n9481), .A(n6066), .B(n6065), .ZN(P1_U3249) );
  INV_X1 U7713 ( .A(n7361), .ZN(n6190) );
  AOI22_X1 U7714 ( .A1(n8891), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9221), .ZN(n6068) );
  OAI21_X1 U7715 ( .B1(n6190), .B2(n4396), .A(n6068), .ZN(P1_U3336) );
  NAND2_X1 U7716 ( .A1(n6111), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7717 ( .A1(n6096), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6073) );
  INV_X1 U7718 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6071) );
  INV_X1 U7719 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6078) );
  AND2_X1 U7720 ( .A1(n6548), .A2(n6749), .ZN(n6086) );
  NAND2_X1 U7721 ( .A1(n6752), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7722 ( .A1(n6087), .A2(n6081), .ZN(n6750) );
  OR2_X1 U7723 ( .A1(n6423), .A2(n6247), .ZN(n6091) );
  NAND2_X1 U7724 ( .A1(n6103), .A2(n6094), .ZN(n6356) );
  INV_X1 U7725 ( .A(n6095), .ZN(n6110) );
  NAND2_X1 U7726 ( .A1(n6110), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7727 ( .A1(n6096), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7728 ( .A1(n6145), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7729 ( .A1(n6111), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7730 ( .A1(n7555), .A2(SI_0_), .ZN(n6101) );
  XNOR2_X1 U7731 ( .A(n6101), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8731) );
  MUX2_X1 U7732 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8731), .S(n6423), .Z(n6776) );
  INV_X1 U7733 ( .A(n6103), .ZN(n6104) );
  OR2_X1 U7734 ( .A1(n6310), .A2(n6105), .ZN(n6108) );
  OR2_X1 U7735 ( .A1(n6203), .A2(n6106), .ZN(n6107) );
  OAI211_X1 U7736 ( .C1(n6423), .C2(n6109), .A(n6108), .B(n6107), .ZN(n6818)
         );
  XNOR2_X1 U7737 ( .A(n6102), .B(n9703), .ZN(n6210) );
  NAND2_X1 U7738 ( .A1(n6110), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7739 ( .A1(n6111), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7740 ( .A1(n6145), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6112) );
  AND3_X1 U7741 ( .A1(n6114), .A2(n6113), .A3(n6112), .ZN(n6116) );
  NAND2_X1 U7742 ( .A1(n6096), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7743 ( .A1(n6116), .A2(n6115), .ZN(n6820) );
  NAND2_X1 U7744 ( .A1(n8279), .A2(n6191), .ZN(n6209) );
  XNOR2_X1 U7745 ( .A(n6210), .B(n6209), .ZN(n6212) );
  XNOR2_X1 U7746 ( .A(n6213), .B(n6212), .ZN(n6153) );
  INV_X1 U7747 ( .A(n6121), .ZN(n7221) );
  NAND2_X1 U7748 ( .A1(n7053), .A2(n7221), .ZN(n9683) );
  XOR2_X1 U7749 ( .A(n7053), .B(P2_B_REG_SCAN_IN), .Z(n6117) );
  INV_X1 U7750 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7751 ( .A1(n9680), .A2(n6119), .ZN(n6120) );
  INV_X1 U7752 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9688) );
  NOR2_X1 U7753 ( .A1(n7174), .A2(n6121), .ZN(n9689) );
  NOR4_X1 U7754 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6125) );
  NOR4_X1 U7755 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6124) );
  NOR4_X1 U7756 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6123) );
  NOR4_X1 U7757 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6122) );
  NAND4_X1 U7758 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(n6131)
         );
  NOR2_X1 U7759 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .ZN(
        n6129) );
  NOR4_X1 U7760 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6128) );
  NOR4_X1 U7761 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6127) );
  NOR4_X1 U7762 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6126) );
  NAND4_X1 U7763 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n6130)
         );
  OAI21_X1 U7764 ( .B1(n6131), .B2(n6130), .A(n9680), .ZN(n8621) );
  NAND2_X1 U7765 ( .A1(n8622), .A2(n8621), .ZN(n6741) );
  INV_X1 U7766 ( .A(n6139), .ZN(n6132) );
  NAND2_X1 U7767 ( .A1(n6087), .A2(n6749), .ZN(n8094) );
  INV_X1 U7768 ( .A(n6746), .ZN(n6225) );
  AND2_X1 U7769 ( .A1(n9776), .A2(n6225), .ZN(n6134) );
  AND2_X1 U7770 ( .A1(n9681), .A2(n9751), .ZN(n6136) );
  INV_X1 U7771 ( .A(n6087), .ZN(n8089) );
  NAND2_X1 U7772 ( .A1(n6139), .A2(n8089), .ZN(n6135) );
  NAND2_X1 U7773 ( .A1(n8094), .A2(n6746), .ZN(n6137) );
  NAND2_X1 U7774 ( .A1(n6226), .A2(n6137), .ZN(n6199) );
  INV_X1 U7775 ( .A(n9690), .ZN(n9684) );
  NAND3_X1 U7776 ( .A1(n6087), .A2(n6138), .A3(n6082), .ZN(n9755) );
  NAND2_X1 U7777 ( .A1(n6139), .A2(n8620), .ZN(n6201) );
  NAND2_X1 U7778 ( .A1(n6744), .A2(n6201), .ZN(n6357) );
  AOI22_X1 U7779 ( .A1(n9584), .A2(n9703), .B1(n6357), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6152) );
  INV_X1 U7780 ( .A(n8094), .ZN(n6140) );
  INV_X1 U7781 ( .A(n9586), .ZN(n9571) );
  INV_X1 U7782 ( .A(n6142), .ZN(n6143) );
  NAND2_X1 U7783 ( .A1(n6111), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6150) );
  INV_X2 U7784 ( .A(n7448), .ZN(n7489) );
  NAND2_X1 U7785 ( .A1(n7489), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6149) );
  INV_X1 U7786 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6144) );
  INV_X1 U7787 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7788 ( .A1(n6746), .A2(n6142), .ZN(n9613) );
  OAI22_X1 U7789 ( .A1(n6754), .A2(n9611), .B1(n6824), .B2(n9613), .ZN(n9661)
         );
  NAND2_X1 U7790 ( .A1(n9571), .A2(n9661), .ZN(n6151) );
  OAI211_X1 U7791 ( .C1(n6153), .C2(n8250), .A(n6152), .B(n6151), .ZN(P2_U3239) );
  INV_X1 U7792 ( .A(n6462), .ZN(n6155) );
  AND3_X1 U7793 ( .A1(n6156), .A2(n6155), .A3(n6154), .ZN(n7872) );
  INV_X1 U7794 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9380) );
  XOR2_X1 U7795 ( .A(n6159), .B(n6158), .Z(n9399) );
  NAND2_X1 U7796 ( .A1(n9399), .A2(n8849), .ZN(n6161) );
  AOI22_X1 U7797 ( .A1(n8870), .A2(n6605), .B1(n8839), .B2(n5613), .ZN(n6160)
         );
  OAI211_X1 U7798 ( .C1(n7872), .C2(n9380), .A(n6161), .B(n6160), .ZN(P1_U3230) );
  INV_X1 U7799 ( .A(n9483), .ZN(n9408) );
  NOR2_X1 U7800 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6162), .ZN(n7123) );
  INV_X1 U7801 ( .A(n7123), .ZN(n6163) );
  OAI21_X1 U7802 ( .B1(n9408), .B2(n6164), .A(n6163), .ZN(n6176) );
  XNOR2_X1 U7803 ( .A(n9457), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U7804 ( .A1(n6165), .A2(n6062), .ZN(n6168) );
  INV_X1 U7805 ( .A(n6166), .ZN(n6167) );
  AOI21_X1 U7806 ( .B1(n6169), .B2(n6168), .A(n6167), .ZN(n9437) );
  NAND2_X1 U7807 ( .A1(n9441), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7808 ( .B1(n9441), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6170), .ZN(
        n9436) );
  NOR2_X1 U7809 ( .A1(n9437), .A2(n9436), .ZN(n9435) );
  AOI21_X1 U7810 ( .B1(n9441), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9435), .ZN(
        n9450) );
  NAND2_X1 U7811 ( .A1(n9444), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6171) );
  OAI21_X1 U7812 ( .B1(n9444), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6171), .ZN(
        n9449) );
  NAND2_X1 U7813 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6474), .ZN(n6172) );
  OAI21_X1 U7814 ( .B1(n6474), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6172), .ZN(
        n6173) );
  NOR2_X1 U7815 ( .A1(n6174), .A2(n6173), .ZN(n6473) );
  AOI211_X1 U7816 ( .C1(n6174), .C2(n6173), .A(n6473), .B(n9488), .ZN(n6175)
         );
  AOI211_X1 U7817 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n9495), .A(n6176), .B(
        n6175), .ZN(n6187) );
  INV_X1 U7818 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6177) );
  MUX2_X1 U7819 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6177), .S(n6474), .Z(n6184)
         );
  INV_X1 U7820 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U7821 ( .A1(n9444), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n10080), .B2(
        n6178), .ZN(n9447) );
  AOI21_X1 U7822 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6180), .A(n6179), .ZN(
        n9434) );
  NOR2_X1 U7823 ( .A1(n9441), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6181) );
  AOI21_X1 U7824 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9441), .A(n6181), .ZN(
        n9433) );
  NAND2_X1 U7825 ( .A1(n9434), .A2(n9433), .ZN(n9432) );
  OAI21_X1 U7826 ( .B1(n9441), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9432), .ZN(
        n9446) );
  NAND2_X1 U7827 ( .A1(n9447), .A2(n9446), .ZN(n9445) );
  OAI21_X1 U7828 ( .B1(n9444), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9445), .ZN(
        n9460) );
  INV_X1 U7829 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6182) );
  MUX2_X1 U7830 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6182), .S(n9457), .Z(n9459)
         );
  NAND2_X1 U7831 ( .A1(n9460), .A2(n9459), .ZN(n9458) );
  OAI21_X1 U7832 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9457), .A(n9458), .ZN(
        n6183) );
  NAND2_X1 U7833 ( .A1(n6183), .A2(n6184), .ZN(n6468) );
  OAI21_X1 U7834 ( .B1(n6184), .B2(n6183), .A(n6468), .ZN(n6185) );
  NAND2_X1 U7835 ( .A1(n6185), .A2(n9496), .ZN(n6186) );
  NAND2_X1 U7836 ( .A1(n6187), .A2(n6186), .ZN(P1_U3253) );
  NAND2_X1 U7837 ( .A1(n6188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U7838 ( .A(n6189), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8375) );
  INV_X1 U7839 ( .A(n8375), .ZN(n8367) );
  OAI222_X1 U7840 ( .A1(n8727), .A2(n10038), .B1(n7895), .B2(n6190), .C1(n8367), .C2(P2_U3152), .ZN(P2_U3341) );
  NOR2_X1 U7841 ( .A1(n9586), .A2(n9613), .ZN(n8188) );
  INV_X1 U7842 ( .A(n6776), .ZN(n9691) );
  NAND2_X1 U7843 ( .A1(n8281), .A2(n9691), .ZN(n8056) );
  NOR3_X1 U7844 ( .A1(n8250), .A2(n6193), .A3(n8056), .ZN(n6192) );
  AOI21_X1 U7845 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n6357), .A(n6192), .ZN(
        n6196) );
  AOI21_X1 U7846 ( .B1(n8140), .B2(n8281), .A(n8250), .ZN(n6194) );
  OAI21_X1 U7847 ( .B1(n6194), .B2(n9584), .A(n6776), .ZN(n6195) );
  OAI211_X1 U7848 ( .C1(n6754), .C2(n8244), .A(n6196), .B(n6195), .ZN(P2_U3234) );
  INV_X1 U7849 ( .A(n6197), .ZN(n6198) );
  NOR2_X1 U7850 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U7851 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  OR2_X1 U7852 ( .A1(n6583), .A2(n6204), .ZN(n6208) );
  OR2_X1 U7853 ( .A1(n6310), .A2(n6205), .ZN(n6207) );
  OR2_X1 U7854 ( .A1(n6423), .A2(n6294), .ZN(n6206) );
  AND3_X2 U7855 ( .A1(n6208), .A2(n6207), .A3(n6206), .ZN(n9709) );
  XNOR2_X1 U7856 ( .A(n6102), .B(n9709), .ZN(n6306) );
  NAND2_X1 U7857 ( .A1(n8278), .A2(n8140), .ZN(n6305) );
  XNOR2_X1 U7858 ( .A(n6306), .B(n6305), .ZN(n6307) );
  INV_X1 U7859 ( .A(n6209), .ZN(n6211) );
  XOR2_X1 U7860 ( .A(n6307), .B(n6308), .Z(n6214) );
  NAND2_X1 U7861 ( .A1(n6214), .A2(n9589), .ZN(n6224) );
  NAND2_X1 U7862 ( .A1(n7490), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7863 ( .A1(n7459), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6218) );
  NOR2_X1 U7864 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6215) );
  NOR2_X1 U7865 ( .A1(n6320), .A2(n6215), .ZN(n9633) );
  NAND2_X1 U7866 ( .A1(n6145), .A2(n9633), .ZN(n6217) );
  NAND2_X1 U7867 ( .A1(n7488), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7868 ( .A1(n8277), .A2(n8573), .ZN(n6221) );
  NAND2_X1 U7869 ( .A1(n8279), .A2(n8571), .ZN(n6220) );
  NAND2_X1 U7870 ( .A1(n6221), .A2(n6220), .ZN(n9647) );
  NOR2_X1 U7871 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6146), .ZN(n6288) );
  NOR2_X1 U7872 ( .A1(n9573), .A2(n9709), .ZN(n6222) );
  AOI211_X1 U7873 ( .C1(n9571), .C2(n9647), .A(n6288), .B(n6222), .ZN(n6223)
         );
  OAI211_X1 U7874 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9593), .A(n6224), .B(
        n6223), .ZN(P2_U3220) );
  NAND2_X1 U7875 ( .A1(n9681), .A2(n6225), .ZN(n6229) );
  OR2_X1 U7876 ( .A1(n6142), .A2(P2_U3152), .ZN(n7331) );
  OAI21_X1 U7877 ( .B1(n6226), .B2(n7331), .A(n8100), .ZN(n6227) );
  INV_X1 U7878 ( .A(n6227), .ZN(n6228) );
  NAND2_X1 U7879 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  NAND2_X1 U7880 ( .A1(n6230), .A2(n6423), .ZN(n6237) );
  NAND2_X1 U7881 ( .A1(n6237), .A2(n8280), .ZN(n6254) );
  NAND2_X1 U7882 ( .A1(n6254), .A2(n6142), .ZN(n9595) );
  NOR2_X1 U7883 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10027), .ZN(n9582) );
  INV_X1 U7884 ( .A(n6312), .ZN(n6234) );
  INV_X1 U7885 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9603) );
  INV_X1 U7886 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10093) );
  NOR3_X1 U7887 ( .A1(n9603), .A2(n10093), .A3(n9226), .ZN(n9225) );
  AOI21_X1 U7888 ( .B1(n9229), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9225), .ZN(
        n9238) );
  NAND2_X1 U7889 ( .A1(n9240), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7890 ( .B1(n9240), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6231), .ZN(
        n9237) );
  NOR2_X1 U7891 ( .A1(n9238), .A2(n9237), .ZN(n9236) );
  AOI21_X1 U7892 ( .B1(n9240), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9236), .ZN(
        n6286) );
  NAND2_X1 U7893 ( .A1(n6244), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7894 ( .B1(n6244), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6232), .ZN(
        n6285) );
  NOR2_X1 U7895 ( .A1(n6286), .A2(n6285), .ZN(n6284) );
  INV_X1 U7896 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6233) );
  MUX2_X1 U7897 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6233), .S(n6312), .Z(n6260)
         );
  NAND2_X1 U7898 ( .A1(n6241), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7899 ( .B1(n6241), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6235), .ZN(
        n6296) );
  AOI21_X1 U7900 ( .B1(n6241), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6295), .ZN(
        n6239) );
  NAND2_X1 U7901 ( .A1(n6275), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U7902 ( .B1(n6275), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6236), .ZN(
        n6238) );
  INV_X1 U7903 ( .A(n8095), .ZN(n6253) );
  AOI211_X1 U7904 ( .C1(n6239), .C2(n6238), .A(n6270), .B(n9596), .ZN(n6240)
         );
  AOI211_X1 U7905 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9600), .A(n9582), .B(
        n6240), .ZN(n6258) );
  NAND2_X1 U7906 ( .A1(n6241), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6250) );
  INV_X1 U7907 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6242) );
  MUX2_X1 U7908 ( .A(n6242), .B(P2_REG2_REG_5__SCAN_IN), .S(n6241), .Z(n6243)
         );
  INV_X1 U7909 ( .A(n6243), .ZN(n6302) );
  INV_X1 U7910 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U7911 ( .A(n10122), .B(P2_REG2_REG_4__SCAN_IN), .S(n6312), .Z(n6265)
         );
  NAND2_X1 U7912 ( .A1(n6244), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6249) );
  INV_X1 U7913 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6245) );
  MUX2_X1 U7914 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6245), .S(n6244), .Z(n6290)
         );
  NAND2_X1 U7915 ( .A1(n9240), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6248) );
  INV_X1 U7916 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6246) );
  MUX2_X1 U7917 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6246), .S(n9240), .Z(n9244)
         );
  INV_X1 U7918 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10078) );
  XNOR2_X1 U7919 ( .A(n6247), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9231) );
  NAND3_X1 U7920 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9231), .ZN(n9230) );
  OAI21_X1 U7921 ( .B1(n6247), .B2(n10078), .A(n9230), .ZN(n9243) );
  NAND2_X1 U7922 ( .A1(n9244), .A2(n9243), .ZN(n9242) );
  NAND2_X1 U7923 ( .A1(n6248), .A2(n9242), .ZN(n6291) );
  NAND2_X1 U7924 ( .A1(n6290), .A2(n6291), .ZN(n6289) );
  NAND2_X1 U7925 ( .A1(n6249), .A2(n6289), .ZN(n6266) );
  NAND2_X1 U7926 ( .A1(n6265), .A2(n6266), .ZN(n6264) );
  OAI21_X1 U7927 ( .B1(n6312), .B2(n10122), .A(n6264), .ZN(n6301) );
  NAND2_X1 U7928 ( .A1(n6302), .A2(n6301), .ZN(n6300) );
  NAND2_X1 U7929 ( .A1(n6250), .A2(n6300), .ZN(n6256) );
  INV_X1 U7930 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6251) );
  MUX2_X1 U7931 ( .A(n6251), .B(P2_REG2_REG_6__SCAN_IN), .S(n6275), .Z(n6252)
         );
  INV_X1 U7932 ( .A(n6252), .ZN(n6255) );
  NAND2_X1 U7933 ( .A1(n6254), .A2(n6253), .ZN(n8394) );
  NAND2_X1 U7934 ( .A1(n6255), .A2(n6256), .ZN(n6276) );
  OAI211_X1 U7935 ( .C1(n6256), .C2(n6255), .A(n9598), .B(n6276), .ZN(n6257)
         );
  OAI211_X1 U7936 ( .C1(n9595), .C2(n6422), .A(n6258), .B(n6257), .ZN(P2_U3251) );
  INV_X1 U7937 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U7938 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10026), .ZN(n6263) );
  AOI211_X1 U7939 ( .C1(n6261), .C2(n6260), .A(n6259), .B(n9596), .ZN(n6262)
         );
  AOI211_X1 U7940 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9600), .A(n6263), .B(
        n6262), .ZN(n6268) );
  OAI211_X1 U7941 ( .C1(n6266), .C2(n6265), .A(n9598), .B(n6264), .ZN(n6267)
         );
  OAI211_X1 U7942 ( .C1(n9595), .C2(n6312), .A(n6268), .B(n6267), .ZN(P2_U3249) );
  INV_X1 U7943 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6269) );
  NOR2_X1 U7944 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6269), .ZN(n6516) );
  INV_X1 U7945 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6271) );
  MUX2_X1 U7946 ( .A(n6271), .B(P2_REG1_REG_7__SCAN_IN), .S(n6428), .Z(n8289)
         );
  INV_X1 U7947 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6272) );
  MUX2_X1 U7948 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6272), .S(n6389), .Z(n6273)
         );
  NOR2_X1 U7949 ( .A1(n4423), .A2(n6273), .ZN(n6390) );
  AOI211_X1 U7950 ( .C1(n4423), .C2(n6273), .A(n6390), .B(n9596), .ZN(n6274)
         );
  AOI211_X1 U7951 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9600), .A(n6516), .B(
        n6274), .ZN(n6283) );
  INV_X1 U7952 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6278) );
  MUX2_X1 U7953 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6278), .S(n6428), .Z(n8283)
         );
  NAND2_X1 U7954 ( .A1(n6275), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7955 ( .A1(n6277), .A2(n6276), .ZN(n8284) );
  NAND2_X1 U7956 ( .A1(n8283), .A2(n8284), .ZN(n8282) );
  OAI21_X1 U7957 ( .B1(n8286), .B2(n6278), .A(n8282), .ZN(n6281) );
  INV_X1 U7958 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6279) );
  MUX2_X1 U7959 ( .A(n6279), .B(P2_REG2_REG_8__SCAN_IN), .S(n6389), .Z(n6280)
         );
  NAND2_X1 U7960 ( .A1(n6280), .A2(n6281), .ZN(n6384) );
  OAI211_X1 U7961 ( .C1(n6281), .C2(n6280), .A(n9598), .B(n6384), .ZN(n6282)
         );
  OAI211_X1 U7962 ( .C1(n9595), .C2(n6389), .A(n6283), .B(n6282), .ZN(P2_U3253) );
  AOI211_X1 U7963 ( .C1(n6286), .C2(n6285), .A(n6284), .B(n9596), .ZN(n6287)
         );
  AOI211_X1 U7964 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9600), .A(n6288), .B(
        n6287), .ZN(n6293) );
  OAI211_X1 U7965 ( .C1(n6291), .C2(n6290), .A(n9598), .B(n6289), .ZN(n6292)
         );
  OAI211_X1 U7966 ( .C1(n9595), .C2(n6294), .A(n6293), .B(n6292), .ZN(P2_U3248) );
  INV_X1 U7967 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6370) );
  NOR2_X1 U7968 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6370), .ZN(n6299) );
  AOI211_X1 U7969 ( .C1(n6297), .C2(n6296), .A(n6295), .B(n9596), .ZN(n6298)
         );
  AOI211_X1 U7970 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9600), .A(n6299), .B(
        n6298), .ZN(n6304) );
  OAI211_X1 U7971 ( .C1(n6302), .C2(n6301), .A(n9598), .B(n6300), .ZN(n6303)
         );
  OAI211_X1 U7972 ( .C1(n9595), .C2(n6369), .A(n6304), .B(n6303), .ZN(P2_U3250) );
  OR2_X1 U7973 ( .A1(n6583), .A2(n6309), .ZN(n6315) );
  OR2_X1 U7974 ( .A1(n7905), .A2(n6311), .ZN(n6314) );
  OR2_X1 U7975 ( .A1(n6423), .A2(n6312), .ZN(n6313) );
  XNOR2_X1 U7976 ( .A(n8179), .B(n9717), .ZN(n6317) );
  NAND2_X1 U7977 ( .A1(n8277), .A2(n8140), .ZN(n6316) );
  NAND2_X1 U7978 ( .A1(n6317), .A2(n6316), .ZN(n6362) );
  OAI21_X1 U7979 ( .B1(n6317), .B2(n6316), .A(n6362), .ZN(n6318) );
  AOI21_X1 U7980 ( .B1(n6319), .B2(n6318), .A(n6364), .ZN(n6330) );
  NAND2_X1 U7981 ( .A1(n6320), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6371) );
  OAI21_X1 U7982 ( .B1(n6320), .B2(P2_REG3_REG_5__SCAN_IN), .A(n6371), .ZN(
        n9622) );
  OR2_X1 U7983 ( .A1(n7480), .A2(n9622), .ZN(n6324) );
  NAND2_X1 U7984 ( .A1(n7489), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7985 ( .A1(n7488), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7986 ( .A1(n7490), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6321) );
  NAND4_X1 U7987 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(n8276)
         );
  NAND2_X1 U7988 ( .A1(n8276), .A2(n8573), .ZN(n6326) );
  NAND2_X1 U7989 ( .A1(n8278), .A2(n8571), .ZN(n6325) );
  NAND2_X1 U7990 ( .A1(n6326), .A2(n6325), .ZN(n9625) );
  AOI22_X1 U7991 ( .A1(n9571), .A2(n9625), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6327) );
  OAI21_X1 U7992 ( .B1(n9717), .B2(n9573), .A(n6327), .ZN(n6328) );
  AOI21_X1 U7993 ( .B1(n9633), .B2(n8258), .A(n6328), .ZN(n6329) );
  OAI21_X1 U7994 ( .B1(n6330), .B2(n8250), .A(n6329), .ZN(P2_U3232) );
  NAND2_X1 U7995 ( .A1(n6332), .A2(n6331), .ZN(n6334) );
  XOR2_X1 U7996 ( .A(n6334), .B(n6333), .Z(n6339) );
  INV_X1 U7997 ( .A(n5619), .ZN(n6335) );
  OAI22_X1 U7998 ( .A1(n8868), .A2(n7596), .B1(n6335), .B2(n8852), .ZN(n6337)
         );
  INV_X1 U7999 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U8000 ( .A1(n7872), .A2(n9505), .ZN(n6336) );
  AOI211_X1 U8001 ( .C1(n5162), .C2(n8870), .A(n6337), .B(n6336), .ZN(n6338)
         );
  OAI21_X1 U8002 ( .B1(n6339), .B2(n8872), .A(n6338), .ZN(P1_U3220) );
  OR2_X1 U8003 ( .A1(n9534), .A2(n5599), .ZN(n6346) );
  OAI21_X1 U8004 ( .B1(n6342), .B2(P1_D_REG_1__SCAN_IN), .A(n6340), .ZN(n6344)
         );
  OR2_X1 U8005 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  AND2_X1 U8006 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  INV_X1 U8007 ( .A(n6461), .ZN(n6347) );
  NOR2_X1 U8008 ( .A1(n6462), .A2(n6347), .ZN(n6348) );
  INV_X1 U8009 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6353) );
  AND2_X1 U8010 ( .A1(n5619), .A2(n6452), .ZN(n7595) );
  NOR2_X1 U8011 ( .A1(n6455), .A2(n7595), .ZN(n7798) );
  INV_X1 U8012 ( .A(n6349), .ZN(n7836) );
  NOR3_X1 U8013 ( .A1(n7798), .A2(n7836), .A3(n6350), .ZN(n6351) );
  AOI21_X1 U8014 ( .B1(n9251), .B2(n5613), .A(n6351), .ZN(n6608) );
  OAI21_X1 U8015 ( .B1(n6452), .B2(n6603), .A(n6608), .ZN(n9200) );
  NAND2_X1 U8016 ( .A1(n9200), .A2(n9556), .ZN(n6352) );
  OAI21_X1 U8017 ( .B1(n9556), .B2(n6353), .A(n6352), .ZN(P1_U3454) );
  AOI21_X1 U8018 ( .B1(n6356), .B2(n6355), .A(n6354), .ZN(n6361) );
  NOR2_X1 U8019 ( .A1(n9586), .A2(n9611), .ZN(n8187) );
  INV_X1 U8020 ( .A(n6820), .ZN(n6819) );
  AOI22_X1 U8021 ( .A1(n9584), .A2(n4631), .B1(n6357), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U8022 ( .B1(n8244), .B2(n6819), .A(n6358), .ZN(n6359) );
  AOI21_X1 U8023 ( .B1(n8187), .B2(n8281), .A(n6359), .ZN(n6360) );
  OAI21_X1 U8024 ( .B1(n6361), .B2(n8250), .A(n6360), .ZN(P2_U3224) );
  INV_X1 U8025 ( .A(n6362), .ZN(n6363) );
  OR2_X1 U8026 ( .A1(n6583), .A2(n6365), .ZN(n6368) );
  OR2_X1 U8027 ( .A1(n7905), .A2(n6366), .ZN(n6367) );
  XNOR2_X1 U8028 ( .A(n8179), .B(n4395), .ZN(n6414) );
  NAND2_X1 U8029 ( .A1(n8276), .A2(n8140), .ZN(n6413) );
  XNOR2_X1 U8030 ( .A(n6414), .B(n6413), .ZN(n6416) );
  XNOR2_X1 U8031 ( .A(n6417), .B(n6416), .ZN(n6381) );
  INV_X1 U8032 ( .A(n9622), .ZN(n6379) );
  INV_X1 U8033 ( .A(n4395), .ZN(n9725) );
  OAI22_X1 U8034 ( .A1(n9573), .A2(n9725), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6370), .ZN(n6378) );
  INV_X1 U8035 ( .A(n8277), .ZN(n9610) );
  AND2_X1 U8036 ( .A1(n6371), .A2(n10027), .ZN(n6372) );
  OR2_X1 U8037 ( .A1(n6372), .A2(n6432), .ZN(n9592) );
  OR2_X1 U8038 ( .A1(n7480), .A2(n9592), .ZN(n6376) );
  NAND2_X1 U8039 ( .A1(n7459), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6375) );
  INV_X4 U8040 ( .A(n7389), .ZN(n7490) );
  NAND2_X1 U8041 ( .A1(n7490), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8042 ( .A1(n7488), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6373) );
  NAND4_X1 U8043 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n8275)
         );
  INV_X1 U8044 ( .A(n8275), .ZN(n9612) );
  OAI22_X1 U8045 ( .A1(n9610), .A2(n8245), .B1(n8244), .B2(n9612), .ZN(n6377)
         );
  AOI211_X1 U8046 ( .C1(n6379), .C2(n8258), .A(n6378), .B(n6377), .ZN(n6380)
         );
  OAI21_X1 U8047 ( .B1(n6381), .B2(n8250), .A(n6380), .ZN(P2_U3229) );
  NAND2_X1 U8048 ( .A1(n6585), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6386) );
  INV_X1 U8049 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6382) );
  MUX2_X1 U8050 ( .A(n6382), .B(P2_REG2_REG_10__SCAN_IN), .S(n6585), .Z(n6383)
         );
  INV_X1 U8051 ( .A(n6383), .ZN(n8308) );
  NAND2_X1 U8052 ( .A1(n6570), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6385) );
  INV_X1 U8053 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6850) );
  MUX2_X1 U8054 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6850), .S(n6570), .Z(n8297)
         );
  OAI21_X1 U8055 ( .B1(n6389), .B2(n6279), .A(n6384), .ZN(n8296) );
  NAND2_X1 U8056 ( .A1(n8297), .A2(n8296), .ZN(n8295) );
  NAND2_X1 U8057 ( .A1(n6385), .A2(n8295), .ZN(n8309) );
  NAND2_X1 U8058 ( .A1(n8308), .A2(n8309), .ZN(n8307) );
  NAND2_X1 U8059 ( .A1(n6386), .A2(n8307), .ZN(n6388) );
  INV_X1 U8060 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6890) );
  MUX2_X1 U8061 ( .A(n6890), .B(P2_REG2_REG_11__SCAN_IN), .S(n6656), .Z(n6387)
         );
  NOR2_X1 U8062 ( .A1(n6388), .A2(n6387), .ZN(n6483) );
  AOI21_X1 U8063 ( .B1(n6388), .B2(n6387), .A(n6483), .ZN(n6400) );
  INV_X1 U8064 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6659) );
  NOR2_X1 U8065 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6659), .ZN(n6397) );
  INV_X1 U8066 ( .A(n6389), .ZN(n6503) );
  INV_X1 U8067 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6391) );
  MUX2_X1 U8068 ( .A(n6391), .B(P2_REG1_REG_9__SCAN_IN), .S(n6570), .Z(n8301)
         );
  INV_X1 U8069 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6392) );
  MUX2_X1 U8070 ( .A(n6392), .B(P2_REG1_REG_10__SCAN_IN), .S(n6585), .Z(n8314)
         );
  AOI21_X1 U8071 ( .B1(n6585), .B2(P2_REG1_REG_10__SCAN_IN), .A(n8312), .ZN(
        n6395) );
  INV_X1 U8072 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6393) );
  MUX2_X1 U8073 ( .A(n6393), .B(P2_REG1_REG_11__SCAN_IN), .S(n6656), .Z(n6394)
         );
  NOR2_X1 U8074 ( .A1(n6395), .A2(n6394), .ZN(n6488) );
  AOI211_X1 U8075 ( .C1(n6395), .C2(n6394), .A(n6488), .B(n9596), .ZN(n6396)
         );
  AOI211_X1 U8076 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9600), .A(n6397), .B(
        n6396), .ZN(n6399) );
  INV_X1 U8077 ( .A(n9595), .ZN(n9241) );
  NAND2_X1 U8078 ( .A1(n9241), .A2(n6656), .ZN(n6398) );
  OAI211_X1 U8079 ( .C1(n6400), .C2(n8390), .A(n6399), .B(n6398), .ZN(P2_U3256) );
  INV_X1 U8080 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6401) );
  INV_X1 U8081 ( .A(n7368), .ZN(n6403) );
  INV_X1 U8082 ( .A(n9482), .ZN(n7536) );
  OAI222_X1 U8083 ( .A1(n8103), .A2(n6401), .B1(n4396), .B2(n6403), .C1(
        P1_U3084), .C2(n7536), .ZN(P1_U3335) );
  INV_X1 U8084 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6404) );
  XNOR2_X1 U8085 ( .A(n6402), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8385) );
  INV_X1 U8086 ( .A(n8385), .ZN(n8372) );
  OAI222_X1 U8087 ( .A1(n8727), .A2(n6404), .B1(n7895), .B2(n6403), .C1(
        P2_U3152), .C2(n8372), .ZN(P2_U3340) );
  XNOR2_X1 U8088 ( .A(n6406), .B(n6405), .ZN(n6411) );
  AOI22_X1 U8089 ( .A1(n8870), .A2(n5190), .B1(n8886), .B2(n8839), .ZN(n6409)
         );
  AOI21_X1 U8090 ( .B1(n8865), .B2(n5631), .A(n6407), .ZN(n6408) );
  OAI211_X1 U8091 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8812), .A(n6409), .B(
        n6408), .ZN(n6410) );
  AOI21_X1 U8092 ( .B1(n6411), .B2(n8849), .A(n6410), .ZN(n6412) );
  INV_X1 U8093 ( .A(n6412), .ZN(P1_U3216) );
  INV_X1 U8094 ( .A(n6413), .ZN(n6415) );
  AND2_X1 U8095 ( .A1(n8275), .A2(n8140), .ZN(n6425) );
  OR2_X1 U8096 ( .A1(n6583), .A2(n6418), .ZN(n6421) );
  OR2_X1 U8097 ( .A1(n7905), .A2(n6419), .ZN(n6420) );
  XNOR2_X1 U8098 ( .A(n8179), .B(n9583), .ZN(n6424) );
  NOR2_X1 U8099 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  AOI21_X1 U8100 ( .B1(n6425), .B2(n6424), .A(n6426), .ZN(n9581) );
  INV_X1 U8101 ( .A(n6426), .ZN(n6427) );
  AOI22_X1 U8102 ( .A1(n7370), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7369), .B2(
        n6428), .ZN(n6431) );
  OR2_X1 U8103 ( .A1(n6429), .A2(n6583), .ZN(n6430) );
  AND2_X2 U8104 ( .A1(n6431), .A2(n6430), .ZN(n7891) );
  XNOR2_X1 U8105 ( .A(n7891), .B(n8179), .ZN(n6499) );
  NOR2_X1 U8106 ( .A1(n6432), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6433) );
  OR2_X1 U8107 ( .A1(n6438), .A2(n6433), .ZN(n7890) );
  OR2_X1 U8108 ( .A1(n7480), .A2(n7890), .ZN(n6437) );
  NAND2_X1 U8109 ( .A1(n7459), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8110 ( .A1(n7490), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8111 ( .A1(n7488), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6434) );
  NAND4_X1 U8112 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n8274)
         );
  NAND2_X1 U8113 ( .A1(n8274), .A2(n8140), .ZN(n6498) );
  XNOR2_X1 U8114 ( .A(n6499), .B(n6498), .ZN(n6500) );
  XNOR2_X1 U8115 ( .A(n6501), .B(n6500), .ZN(n6448) );
  NOR2_X1 U8116 ( .A1(n6438), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6439) );
  OR2_X1 U8117 ( .A1(n6506), .A2(n6439), .ZN(n7046) );
  OR2_X1 U8118 ( .A1(n7480), .A2(n7046), .ZN(n6443) );
  NAND2_X1 U8119 ( .A1(n7459), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8120 ( .A1(n7488), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8121 ( .A1(n7490), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6440) );
  NAND4_X1 U8122 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n8273)
         );
  INV_X1 U8123 ( .A(n7890), .ZN(n6444) );
  AOI22_X1 U8124 ( .A1(n8188), .A2(n8273), .B1(n8258), .B2(n6444), .ZN(n6447)
         );
  INV_X1 U8125 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U8126 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10123), .ZN(n8285) );
  NOR2_X1 U8127 ( .A1(n9573), .A2(n7891), .ZN(n6445) );
  AOI211_X1 U8128 ( .C1(n8187), .C2(n8275), .A(n8285), .B(n6445), .ZN(n6446)
         );
  OAI211_X1 U8129 ( .C1(n6448), .C2(n8250), .A(n6447), .B(n6446), .ZN(P2_U3215) );
  INV_X1 U8130 ( .A(n9534), .ZN(n9553) );
  OAI21_X1 U8131 ( .B1(n6451), .B2(n6450), .A(n6449), .ZN(n9501) );
  INV_X1 U8132 ( .A(n9501), .ZN(n6460) );
  OAI211_X1 U8133 ( .C1(n6452), .C2(n9507), .A(n9530), .B(n6717), .ZN(n9500)
         );
  OAI21_X1 U8134 ( .B1(n9507), .B2(n9546), .A(n9500), .ZN(n6459) );
  AOI22_X1 U8135 ( .A1(n9251), .A2(n5631), .B1(n5619), .B2(n9254), .ZN(n6458)
         );
  NAND2_X1 U8136 ( .A1(n6456), .A2(n9065), .ZN(n6457) );
  OAI211_X1 U8137 ( .C1(n9501), .C2(n6906), .A(n6458), .B(n6457), .ZN(n9510)
         );
  AOI211_X1 U8138 ( .C1(n9553), .C2(n6460), .A(n6459), .B(n9510), .ZN(n6467)
         );
  NOR2_X1 U8139 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U8140 ( .A1(n9563), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6465) );
  OAI21_X1 U8141 ( .B1(n6467), .B2(n9563), .A(n6465), .ZN(P1_U3524) );
  NAND2_X1 U8142 ( .A1(n9554), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6466) );
  OAI21_X1 U8143 ( .B1(n6467), .B2(n9554), .A(n6466), .ZN(P1_U3457) );
  INV_X1 U8144 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U8145 ( .B1(n6474), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6468), .ZN(
        n6471) );
  INV_X1 U8146 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6469) );
  MUX2_X1 U8147 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6469), .S(n6925), .Z(n6470)
         );
  NAND2_X1 U8148 ( .A1(n6470), .A2(n6471), .ZN(n6924) );
  OAI21_X1 U8149 ( .B1(n6471), .B2(n6470), .A(n6924), .ZN(n6472) );
  NAND2_X1 U8150 ( .A1(n6472), .A2(n9496), .ZN(n6480) );
  AND2_X1 U8151 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7134) );
  MUX2_X1 U8152 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n4560), .S(n6925), .Z(n6475)
         );
  INV_X1 U8153 ( .A(n6475), .ZN(n6476) );
  AOI211_X1 U8154 ( .C1(n6477), .C2(n6476), .A(n6919), .B(n9488), .ZN(n6478)
         );
  AOI211_X1 U8155 ( .C1(n9483), .C2(n6925), .A(n7134), .B(n6478), .ZN(n6479)
         );
  OAI211_X1 U8156 ( .C1(n9481), .C2(n6481), .A(n6480), .B(n6479), .ZN(P1_U3254) );
  INV_X1 U8157 ( .A(n7358), .ZN(n7545) );
  OAI222_X1 U8158 ( .A1(n8727), .A2(n6482), .B1(n7895), .B2(n7545), .C1(
        P2_U3152), .C2(n6749), .ZN(P2_U3339) );
  NOR2_X1 U8159 ( .A1(n6656), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6484) );
  NOR2_X1 U8160 ( .A1(n6484), .A2(n6483), .ZN(n6487) );
  INV_X1 U8161 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6485) );
  MUX2_X1 U8162 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6485), .S(n6953), .Z(n6486)
         );
  NAND2_X1 U8163 ( .A1(n6953), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6610) );
  OAI211_X1 U8164 ( .C1(n6953), .C2(P2_REG2_REG_12__SCAN_IN), .A(n6487), .B(
        n6610), .ZN(n6609) );
  OAI211_X1 U8165 ( .C1(n6487), .C2(n6486), .A(n6609), .B(n9598), .ZN(n6496)
         );
  AOI21_X1 U8166 ( .B1(n6656), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6488), .ZN(
        n6491) );
  INV_X1 U8167 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6489) );
  MUX2_X1 U8168 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6489), .S(n6953), .Z(n6490)
         );
  NAND2_X1 U8169 ( .A1(n6490), .A2(n6491), .ZN(n6613) );
  OAI21_X1 U8170 ( .B1(n6491), .B2(n6490), .A(n6613), .ZN(n6494) );
  AND2_X1 U8171 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n6976) );
  INV_X1 U8172 ( .A(n9600), .ZN(n6619) );
  INV_X1 U8173 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U8174 ( .A1(n6619), .A2(n6492), .ZN(n6493) );
  AOI211_X1 U8175 ( .C1(n9594), .C2(n6494), .A(n6976), .B(n6493), .ZN(n6495)
         );
  OAI211_X1 U8176 ( .C1(n9595), .C2(n6497), .A(n6496), .B(n6495), .ZN(P2_U3257) );
  OR2_X1 U8177 ( .A1(n6502), .A2(n6583), .ZN(n6505) );
  AOI22_X1 U8178 ( .A1(n7370), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7369), .B2(
        n6503), .ZN(n6504) );
  NAND2_X1 U8179 ( .A1(n6505), .A2(n6504), .ZN(n7941) );
  XNOR2_X1 U8180 ( .A(n7941), .B(n8179), .ZN(n6565) );
  NAND2_X1 U8181 ( .A1(n8273), .A2(n8140), .ZN(n6564) );
  XNOR2_X1 U8182 ( .A(n6565), .B(n6564), .ZN(n6567) );
  XNOR2_X1 U8183 ( .A(n6568), .B(n6567), .ZN(n6521) );
  NOR2_X1 U8184 ( .A1(n9593), .A2(n7046), .ZN(n6519) );
  INV_X1 U8185 ( .A(n6506), .ZN(n6508) );
  INV_X1 U8186 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U8187 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  NAND2_X1 U8188 ( .A1(n6577), .A2(n6509), .ZN(n9578) );
  OR2_X1 U8189 ( .A1(n7480), .A2(n9578), .ZN(n6513) );
  NAND2_X1 U8190 ( .A1(n7459), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U8191 ( .A1(n7488), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U8192 ( .A1(n7490), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6510) );
  NAND4_X1 U8193 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n8272)
         );
  NAND2_X1 U8194 ( .A1(n8272), .A2(n8573), .ZN(n6515) );
  NAND2_X1 U8195 ( .A1(n8274), .A2(n8571), .ZN(n6514) );
  AND2_X1 U8196 ( .A1(n6515), .A2(n6514), .ZN(n7043) );
  INV_X1 U8197 ( .A(n6516), .ZN(n6517) );
  OAI21_X1 U8198 ( .B1(n9586), .B2(n7043), .A(n6517), .ZN(n6518) );
  AOI211_X1 U8199 ( .C1(n9584), .C2(n7941), .A(n6519), .B(n6518), .ZN(n6520)
         );
  OAI21_X1 U8200 ( .B1(n6521), .B2(n8250), .A(n6520), .ZN(P2_U3223) );
  INV_X1 U8201 ( .A(n6522), .ZN(n6523) );
  AOI211_X1 U8202 ( .C1(n6525), .C2(n6524), .A(n8872), .B(n6523), .ZN(n6530)
         );
  INV_X1 U8203 ( .A(n6526), .ZN(n6731) );
  AOI22_X1 U8204 ( .A1(n8870), .A2(n6737), .B1(n8885), .B2(n8839), .ZN(n6528)
         );
  AND2_X1 U8205 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9423) );
  AOI21_X1 U8206 ( .B1(n8887), .B2(n8865), .A(n9423), .ZN(n6527) );
  OAI211_X1 U8207 ( .C1(n8812), .C2(n6731), .A(n6528), .B(n6527), .ZN(n6529)
         );
  OR2_X1 U8208 ( .A1(n6530), .A2(n6529), .ZN(P1_U3228) );
  INV_X1 U8209 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U8210 ( .B1(n6532), .B2(n6537), .A(n6531), .ZN(n6692) );
  INV_X1 U8211 ( .A(n6719), .ZN(n6534) );
  INV_X1 U8212 ( .A(n6734), .ZN(n6533) );
  OAI21_X1 U8213 ( .B1(n6535), .B2(n6534), .A(n6533), .ZN(n6688) );
  OAI22_X1 U8214 ( .A1(n6688), .A2(n9548), .B1(n6535), .B2(n9546), .ZN(n6541)
         );
  XNOR2_X1 U8215 ( .A(n6536), .B(n6537), .ZN(n6540) );
  INV_X1 U8216 ( .A(n6906), .ZN(n9259) );
  NAND2_X1 U8217 ( .A1(n6692), .A2(n9259), .ZN(n6539) );
  AOI22_X1 U8218 ( .A1(n8886), .A2(n9251), .B1(n9254), .B2(n5631), .ZN(n6538)
         );
  OAI211_X1 U8219 ( .C1(n9256), .C2(n6540), .A(n6539), .B(n6538), .ZN(n6689)
         );
  AOI211_X1 U8220 ( .C1(n9553), .C2(n6692), .A(n6541), .B(n6689), .ZN(n6544)
         );
  OR2_X1 U8221 ( .A1(n6544), .A2(n9554), .ZN(n6542) );
  OAI21_X1 U8222 ( .B1(n9556), .B2(n6543), .A(n6542), .ZN(P1_U3463) );
  INV_X1 U8223 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6546) );
  OR2_X1 U8224 ( .A1(n6544), .A2(n9563), .ZN(n6545) );
  OAI21_X1 U8225 ( .B1(n9565), .B2(n6546), .A(n6545), .ZN(P1_U3526) );
  INV_X1 U8226 ( .A(n7380), .ZN(n6549) );
  OAI222_X1 U8227 ( .A1(n4396), .A2(n6549), .B1(P1_U3084), .B2(n7825), .C1(
        n6547), .C2(n8108), .ZN(P1_U3332) );
  OAI222_X1 U8228 ( .A1(n8727), .A2(n7381), .B1(n7895), .B2(n6549), .C1(n6548), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8229 ( .A1(n6724), .A2(n6550), .ZN(n6791) );
  INV_X1 U8230 ( .A(n6897), .ZN(n6551) );
  AOI21_X1 U8231 ( .B1(n6902), .B2(n6791), .A(n6551), .ZN(n6865) );
  NAND2_X1 U8232 ( .A1(n6906), .A2(n9534), .ZN(n9537) );
  AOI21_X1 U8233 ( .B1(n6733), .B2(n5247), .A(n9548), .ZN(n6552) );
  NAND2_X1 U8234 ( .A1(n6552), .A2(n6912), .ZN(n6855) );
  OR2_X1 U8235 ( .A1(n7853), .A2(n9104), .ZN(n6856) );
  OAI211_X1 U8236 ( .C1(n6553), .C2(n9546), .A(n6855), .B(n6856), .ZN(n6554)
         );
  AOI21_X1 U8237 ( .B1(n6865), .B2(n9537), .A(n6554), .ZN(n6559) );
  XNOR2_X1 U8238 ( .A(n6555), .B(n6902), .ZN(n6558) );
  NOR2_X1 U8239 ( .A1(n6556), .A2(n5525), .ZN(n6557) );
  AOI21_X1 U8240 ( .B1(n6558), .B2(n9065), .A(n6557), .ZN(n6858) );
  NAND2_X1 U8241 ( .A1(n6559), .A2(n6858), .ZN(n6561) );
  NAND2_X1 U8242 ( .A1(n6561), .A2(n9565), .ZN(n6560) );
  OAI21_X1 U8243 ( .B1(n9565), .B2(n6029), .A(n6560), .ZN(P1_U3528) );
  INV_X1 U8244 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8245 ( .A1(n6561), .A2(n9556), .ZN(n6562) );
  OAI21_X1 U8246 ( .B1(n9556), .B2(n6563), .A(n6562), .ZN(P1_U3469) );
  INV_X1 U8247 ( .A(n6564), .ZN(n6566) );
  AND2_X1 U8248 ( .A1(n8272), .A2(n8140), .ZN(n6574) );
  OR2_X1 U8249 ( .A1(n6569), .A2(n6583), .ZN(n6572) );
  AOI22_X1 U8250 ( .A1(n7370), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7369), .B2(
        n6570), .ZN(n6571) );
  NAND2_X1 U8251 ( .A1(n6572), .A2(n6571), .ZN(n9750) );
  XNOR2_X1 U8252 ( .A(n9750), .B(n8179), .ZN(n6573) );
  NOR2_X1 U8253 ( .A1(n6573), .A2(n6574), .ZN(n6575) );
  AOI21_X1 U8254 ( .B1(n6574), .B2(n6573), .A(n6575), .ZN(n9567) );
  INV_X1 U8255 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U8256 ( .A1(n6577), .A2(n6594), .ZN(n6578) );
  NAND2_X1 U8257 ( .A1(n6661), .A2(n6578), .ZN(n6996) );
  OR2_X1 U8258 ( .A1(n7480), .A2(n6996), .ZN(n6582) );
  NAND2_X1 U8259 ( .A1(n7459), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U8260 ( .A1(n7490), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8261 ( .A1(n7488), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6579) );
  NAND4_X1 U8262 ( .A1(n6582), .A2(n6581), .A3(n6580), .A4(n6579), .ZN(n8271)
         );
  NAND2_X1 U8263 ( .A1(n8271), .A2(n8140), .ZN(n6651) );
  NAND2_X1 U8264 ( .A1(n6584), .A2(n7907), .ZN(n6587) );
  AOI22_X1 U8265 ( .A1(n7370), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7369), .B2(
        n6585), .ZN(n6586) );
  NAND2_X1 U8266 ( .A1(n6587), .A2(n6586), .ZN(n6998) );
  XNOR2_X1 U8267 ( .A(n6998), .B(n8179), .ZN(n6650) );
  XOR2_X1 U8268 ( .A(n6651), .B(n6650), .Z(n6653) );
  XNOR2_X1 U8269 ( .A(n6654), .B(n6653), .ZN(n6599) );
  NOR2_X1 U8270 ( .A1(n9593), .A2(n6996), .ZN(n6597) );
  NAND2_X1 U8271 ( .A1(n7459), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8272 ( .A1(n7488), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6590) );
  XNOR2_X1 U8273 ( .A(n6661), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U8274 ( .A1(n6145), .A2(n6658), .ZN(n6589) );
  NAND2_X1 U8275 ( .A1(n7490), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6588) );
  NAND4_X1 U8276 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n8270)
         );
  NAND2_X1 U8277 ( .A1(n8270), .A2(n8573), .ZN(n6593) );
  NAND2_X1 U8278 ( .A1(n8272), .A2(n8571), .ZN(n6592) );
  AND2_X1 U8279 ( .A1(n6593), .A2(n6592), .ZN(n6992) );
  NOR2_X1 U8280 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6594), .ZN(n8310) );
  INV_X1 U8281 ( .A(n8310), .ZN(n6595) );
  OAI21_X1 U8282 ( .B1(n9586), .B2(n6992), .A(n6595), .ZN(n6596) );
  AOI211_X1 U8283 ( .C1(n9584), .C2(n6998), .A(n6597), .B(n6596), .ZN(n6598)
         );
  OAI21_X1 U8284 ( .B1(n6599), .B2(n8250), .A(n6598), .ZN(P2_U3219) );
  INV_X1 U8285 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6600) );
  OAI22_X1 U8286 ( .A1(n9081), .A2(n6600), .B1(n9380), .B2(n9506), .ZN(n6601)
         );
  INV_X1 U8287 ( .A(n6601), .ZN(n6607) );
  NOR2_X1 U8288 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  OAI21_X1 U8289 ( .B1(n9262), .B2(n9068), .A(n6605), .ZN(n6606) );
  OAI211_X1 U8290 ( .C1(n6608), .C2(n9513), .A(n6607), .B(n6606), .ZN(P1_U3291) );
  NAND2_X1 U8291 ( .A1(n6610), .A2(n6609), .ZN(n6612) );
  INV_X1 U8292 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6628) );
  AOI22_X1 U8293 ( .A1(n7058), .A2(n6628), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6629), .ZN(n6611) );
  NOR2_X1 U8294 ( .A1(n6612), .A2(n6611), .ZN(n6627) );
  AOI21_X1 U8295 ( .B1(n6612), .B2(n6611), .A(n6627), .ZN(n6622) );
  INV_X1 U8296 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6618) );
  INV_X1 U8297 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9331) );
  AOI22_X1 U8298 ( .A1(n7058), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9331), .B2(
        n6629), .ZN(n6615) );
  OAI21_X1 U8299 ( .B1(n6953), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6613), .ZN(
        n6614) );
  NAND2_X1 U8300 ( .A1(n6615), .A2(n6614), .ZN(n6623) );
  OAI21_X1 U8301 ( .B1(n6615), .B2(n6614), .A(n6623), .ZN(n6616) );
  NAND2_X1 U8302 ( .A1(n9594), .A2(n6616), .ZN(n6617) );
  NAND2_X1 U8303 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7068) );
  OAI211_X1 U8304 ( .C1(n6619), .C2(n6618), .A(n6617), .B(n7068), .ZN(n6620)
         );
  AOI21_X1 U8305 ( .B1(n7058), .B2(n9241), .A(n6620), .ZN(n6621) );
  OAI21_X1 U8306 ( .B1(n6622), .B2(n8390), .A(n6621), .ZN(P2_U3258) );
  INV_X1 U8307 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9323) );
  AOI22_X1 U8308 ( .A1(n8322), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9323), .B2(
        n6630), .ZN(n6625) );
  OAI21_X1 U8309 ( .B1(n7058), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6623), .ZN(
        n6624) );
  NAND2_X1 U8310 ( .A1(n6625), .A2(n6624), .ZN(n8320) );
  OAI21_X1 U8311 ( .B1(n6625), .B2(n6624), .A(n8320), .ZN(n6637) );
  AND2_X1 U8312 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7236) );
  AOI21_X1 U8313 ( .B1(n9600), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7236), .ZN(
        n6626) );
  OAI21_X1 U8314 ( .B1(n9595), .B2(n6630), .A(n6626), .ZN(n6636) );
  AOI21_X1 U8315 ( .B1(n6629), .B2(n6628), .A(n6627), .ZN(n6633) );
  INV_X1 U8316 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U8317 ( .A1(n8322), .A2(n6631), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6630), .ZN(n6632) );
  NOR2_X1 U8318 ( .A1(n6633), .A2(n6632), .ZN(n8323) );
  AOI21_X1 U8319 ( .B1(n6633), .B2(n6632), .A(n8323), .ZN(n6634) );
  NOR2_X1 U8320 ( .A1(n6634), .A2(n8390), .ZN(n6635) );
  AOI211_X1 U8321 ( .C1(n6637), .C2(n9594), .A(n6636), .B(n6635), .ZN(n6638)
         );
  INV_X1 U8322 ( .A(n6638), .ZN(P2_U3259) );
  XNOR2_X1 U8323 ( .A(n6640), .B(n6639), .ZN(n6641) );
  XNOR2_X1 U8324 ( .A(n6642), .B(n6641), .ZN(n6649) );
  NAND2_X1 U8325 ( .A1(n8863), .A2(n9260), .ZN(n6645) );
  NOR2_X1 U8326 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6643), .ZN(n9452) );
  AOI21_X1 U8327 ( .B1(n8865), .B2(n9253), .A(n9452), .ZN(n6644) );
  OAI211_X1 U8328 ( .C1(n6646), .C2(n8868), .A(n6645), .B(n6644), .ZN(n6647)
         );
  AOI21_X1 U8329 ( .B1(n9263), .B2(n8870), .A(n6647), .ZN(n6648) );
  OAI21_X1 U8330 ( .B1(n6649), .B2(n8872), .A(n6648), .ZN(P1_U3215) );
  INV_X1 U8331 ( .A(n6650), .ZN(n6652) );
  AOI22_X1 U8332 ( .A1(n7370), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7369), .B2(
        n6656), .ZN(n6657) );
  XNOR2_X1 U8333 ( .A(n7026), .B(n8179), .ZN(n6959) );
  NAND2_X1 U8334 ( .A1(n8270), .A2(n8140), .ZN(n6958) );
  XNOR2_X1 U8335 ( .A(n6959), .B(n6958), .ZN(n6961) );
  XNOR2_X1 U8336 ( .A(n6962), .B(n6961), .ZN(n6672) );
  INV_X1 U8337 ( .A(n6658), .ZN(n6889) );
  OAI22_X1 U8338 ( .A1(n9593), .A2(n6889), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6659), .ZN(n6670) );
  INV_X1 U8339 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U8340 ( .B1(n6661), .B2(n6659), .A(n6660), .ZN(n6664) );
  NAND2_X1 U8341 ( .A1(n6664), .A2(n6968), .ZN(n6966) );
  OR2_X1 U8342 ( .A1(n7480), .A2(n6966), .ZN(n6668) );
  NAND2_X1 U8343 ( .A1(n7489), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8344 ( .A1(n7490), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8345 ( .A1(n7488), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6665) );
  NAND4_X1 U8346 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n8269)
         );
  OAI22_X1 U8347 ( .A1(n6888), .A2(n8245), .B1(n8244), .B2(n7082), .ZN(n6669)
         );
  AOI211_X1 U8348 ( .C1(n9584), .C2(n7026), .A(n6670), .B(n6669), .ZN(n6671)
         );
  OAI21_X1 U8349 ( .B1(n6672), .B2(n8250), .A(n6671), .ZN(P2_U3238) );
  INV_X1 U8350 ( .A(n7391), .ZN(n6674) );
  OAI222_X1 U8351 ( .A1(n8108), .A2(n6673), .B1(n4396), .B2(n6674), .C1(n7755), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U8352 ( .A1(n8727), .A2(n7392), .B1(n7895), .B2(n6674), .C1(
        P2_U3152), .C2(n6082), .ZN(P2_U3336) );
  XNOR2_X1 U8353 ( .A(n6675), .B(n6676), .ZN(n6677) );
  NAND2_X1 U8354 ( .A1(n6677), .A2(n6678), .ZN(n6868) );
  OAI21_X1 U8355 ( .B1(n6678), .B2(n6677), .A(n6868), .ZN(n6684) );
  INV_X1 U8356 ( .A(n6679), .ZN(n6857) );
  AOI22_X1 U8357 ( .A1(n8870), .A2(n5247), .B1(n8884), .B2(n8839), .ZN(n6682)
         );
  AOI21_X1 U8358 ( .B1(n8886), .B2(n8865), .A(n6680), .ZN(n6681) );
  OAI211_X1 U8359 ( .C1(n8812), .C2(n6857), .A(n6682), .B(n6681), .ZN(n6683)
         );
  AOI21_X1 U8360 ( .B1(n6684), .B2(n8849), .A(n6683), .ZN(n6685) );
  INV_X1 U8361 ( .A(n6685), .ZN(P1_U3225) );
  NOR3_X1 U8362 ( .A1(n9513), .A2(n5543), .A3(n5611), .ZN(n9270) );
  INV_X1 U8363 ( .A(n9068), .ZN(n7528) );
  AOI22_X1 U8364 ( .A1(n9262), .A2(n5190), .B1(n9261), .B2(n6686), .ZN(n6687)
         );
  OAI21_X1 U8365 ( .B1(n6688), .B2(n7528), .A(n6687), .ZN(n6691) );
  MUX2_X1 U8366 ( .A(n6689), .B(P1_REG2_REG_3__SCAN_IN), .S(n9513), .Z(n6690)
         );
  AOI211_X1 U8367 ( .C1(n4394), .C2(n6692), .A(n6691), .B(n6690), .ZN(n6693)
         );
  INV_X1 U8368 ( .A(n6693), .ZN(P1_U3288) );
  AND2_X1 U8369 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  OR2_X1 U8370 ( .A1(n6696), .A2(n7801), .ZN(n6698) );
  NAND2_X1 U8371 ( .A1(n6696), .A2(n7801), .ZN(n6697) );
  AND2_X1 U8372 ( .A1(n6698), .A2(n6697), .ZN(n9538) );
  INV_X1 U8373 ( .A(n9538), .ZN(n6708) );
  XNOR2_X1 U8374 ( .A(n6699), .B(n7801), .ZN(n6700) );
  NAND2_X1 U8375 ( .A1(n6700), .A2(n9065), .ZN(n6702) );
  AOI22_X1 U8376 ( .A1(n8883), .A2(n9254), .B1(n9251), .B2(n9253), .ZN(n6701)
         );
  NAND2_X1 U8377 ( .A1(n6702), .A2(n6701), .ZN(n9542) );
  OR2_X1 U8378 ( .A1(n6804), .A2(n9539), .ZN(n6703) );
  NAND2_X1 U8379 ( .A1(n6765), .A2(n6703), .ZN(n9540) );
  AOI22_X1 U8380 ( .A1(n9513), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7012), .B2(
        n9261), .ZN(n6705) );
  NAND2_X1 U8381 ( .A1(n9262), .A2(n7018), .ZN(n6704) );
  OAI211_X1 U8382 ( .C1(n9540), .C2(n7528), .A(n6705), .B(n6704), .ZN(n6706)
         );
  AOI21_X1 U8383 ( .B1(n9542), .B2(n9081), .A(n6706), .ZN(n6707) );
  OAI21_X1 U8384 ( .B1(n6708), .B2(n9114), .A(n6707), .ZN(P1_U3283) );
  INV_X1 U8385 ( .A(n6709), .ZN(n6710) );
  AOI21_X1 U8386 ( .B1(n7795), .B2(n6711), .A(n6710), .ZN(n9516) );
  INV_X1 U8387 ( .A(n9270), .ZN(n6918) );
  OAI21_X1 U8388 ( .B1(n7795), .B2(n7597), .A(n6712), .ZN(n6714) );
  OAI22_X1 U8389 ( .A1(n7866), .A2(n5525), .B1(n7867), .B2(n9104), .ZN(n6713)
         );
  AOI21_X1 U8390 ( .B1(n6714), .B2(n9065), .A(n6713), .ZN(n6715) );
  OAI21_X1 U8391 ( .B1(n9516), .B2(n6906), .A(n6715), .ZN(n9519) );
  NAND2_X1 U8392 ( .A1(n9519), .A2(n9081), .ZN(n6723) );
  INV_X1 U8393 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7873) );
  INV_X1 U8394 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6716) );
  OAI22_X1 U8395 ( .A1(n9506), .A2(n7873), .B1(n6716), .B2(n9081), .ZN(n6721)
         );
  NAND2_X1 U8396 ( .A1(n6717), .A2(n7869), .ZN(n6718) );
  NAND2_X1 U8397 ( .A1(n6719), .A2(n6718), .ZN(n9518) );
  NOR2_X1 U8398 ( .A1(n7528), .A2(n9518), .ZN(n6720) );
  AOI211_X1 U8399 ( .C1(n9262), .C2(n7869), .A(n6721), .B(n6720), .ZN(n6722)
         );
  OAI211_X1 U8400 ( .C1(n9516), .C2(n6918), .A(n6723), .B(n6722), .ZN(P1_U3289) );
  OAI21_X1 U8401 ( .B1(n6725), .B2(n6727), .A(n6724), .ZN(n9527) );
  INV_X1 U8402 ( .A(n9527), .ZN(n6740) );
  XNOR2_X1 U8403 ( .A(n6726), .B(n6727), .ZN(n6730) );
  OAI22_X1 U8404 ( .A1(n7867), .A2(n5525), .B1(n6905), .B2(n9104), .ZN(n6728)
         );
  AOI21_X1 U8405 ( .B1(n9527), .B2(n9259), .A(n6728), .ZN(n6729) );
  OAI21_X1 U8406 ( .B1(n9256), .B2(n6730), .A(n6729), .ZN(n9525) );
  NAND2_X1 U8407 ( .A1(n9525), .A2(n5603), .ZN(n6739) );
  OAI22_X1 U8408 ( .A1(n5603), .A2(n6001), .B1(n6731), .B2(n9506), .ZN(n6736)
         );
  NOR2_X1 U8409 ( .A1(n6732), .A2(n5403), .ZN(n9269) );
  INV_X1 U8410 ( .A(n9269), .ZN(n7301) );
  OAI211_X1 U8411 ( .C1(n6734), .C2(n9524), .A(n6733), .B(n9530), .ZN(n9523)
         );
  NOR2_X1 U8412 ( .A1(n7301), .A2(n9523), .ZN(n6735) );
  AOI211_X1 U8413 ( .C1(n9262), .C2(n6737), .A(n6736), .B(n6735), .ZN(n6738)
         );
  OAI211_X1 U8414 ( .C1(n6740), .C2(n6918), .A(n6739), .B(n6738), .ZN(P1_U3287) );
  OR2_X1 U8415 ( .A1(n8281), .A2(n9691), .ZN(n6772) );
  AND2_X1 U8416 ( .A1(n6772), .A2(n8056), .ZN(n9692) );
  INV_X1 U8417 ( .A(n6741), .ZN(n6742) );
  INV_X1 U8418 ( .A(n8620), .ZN(n6745) );
  NOR2_X1 U8419 ( .A1(n6746), .A2(n6138), .ZN(n6748) );
  NAND2_X1 U8420 ( .A1(n6750), .A2(n6082), .ZN(n6747) );
  NAND2_X1 U8421 ( .A1(n6748), .A2(n6747), .ZN(n9640) );
  OR2_X1 U8422 ( .A1(n6750), .A2(n6749), .ZN(n7078) );
  AND2_X1 U8423 ( .A1(n9640), .A2(n7078), .ZN(n6751) );
  OR2_X1 U8424 ( .A1(n6752), .A2(n6087), .ZN(n9617) );
  NOR2_X2 U8425 ( .A1(n6753), .A2(n8140), .ZN(n9668) );
  OAI21_X1 U8426 ( .B1(n9631), .B2(n9668), .A(n6776), .ZN(n6757) );
  INV_X1 U8427 ( .A(n9666), .ZN(n9632) );
  NAND2_X1 U8428 ( .A1(n8097), .A2(n6138), .ZN(n8086) );
  OR2_X1 U8429 ( .A1(n6087), .A2(n6548), .ZN(n7911) );
  OAI22_X1 U8430 ( .A1(n9692), .A2(n9644), .B1(n6754), .B2(n9613), .ZN(n9694)
         );
  AOI21_X1 U8431 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9632), .A(n9694), .ZN(
        n6755) );
  INV_X1 U8432 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9992) );
  MUX2_X1 U8433 ( .A(n6755), .B(n9992), .S(n9669), .Z(n6756) );
  OAI211_X1 U8434 ( .C1(n9692), .C2(n9676), .A(n6757), .B(n6756), .ZN(P2_U3296) );
  NAND2_X1 U8435 ( .A1(n4787), .A2(n7630), .ZN(n7803) );
  XNOR2_X1 U8436 ( .A(n6758), .B(n7803), .ZN(n6764) );
  XNOR2_X1 U8437 ( .A(n6760), .B(n7803), .ZN(n6762) );
  OAI22_X1 U8438 ( .A1(n6801), .A2(n5525), .B1(n7144), .B2(n9104), .ZN(n6761)
         );
  AOI21_X1 U8439 ( .B1(n6762), .B2(n9065), .A(n6761), .ZN(n6763) );
  OAI21_X1 U8440 ( .B1(n6764), .B2(n6906), .A(n6763), .ZN(n9550) );
  INV_X1 U8441 ( .A(n9550), .ZN(n6771) );
  INV_X1 U8442 ( .A(n6764), .ZN(n9552) );
  NAND2_X1 U8443 ( .A1(n6765), .A2(n6949), .ZN(n6766) );
  NAND2_X1 U8444 ( .A1(n9264), .A2(n6766), .ZN(n9549) );
  AOI22_X1 U8445 ( .A1(n9513), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6945), .B2(
        n9261), .ZN(n6768) );
  NAND2_X1 U8446 ( .A1(n9262), .A2(n6949), .ZN(n6767) );
  OAI211_X1 U8447 ( .C1(n9549), .C2(n7528), .A(n6768), .B(n6767), .ZN(n6769)
         );
  AOI21_X1 U8448 ( .B1(n9552), .B2(n4394), .A(n6769), .ZN(n6770) );
  OAI21_X1 U8449 ( .B1(n6771), .B2(n9513), .A(n6770), .ZN(P1_U3282) );
  OAI211_X1 U8450 ( .C1(n6773), .C2(n6772), .A(n8060), .B(n9662), .ZN(n6775)
         );
  AOI22_X1 U8451 ( .A1(n8571), .A2(n8281), .B1(n8279), .B2(n8573), .ZN(n6774)
         );
  NAND2_X1 U8452 ( .A1(n6775), .A2(n6774), .ZN(n9700) );
  AOI21_X1 U8453 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9632), .A(n9700), .ZN(
        n6781) );
  XNOR2_X1 U8454 ( .A(n6815), .B(n6814), .ZN(n9702) );
  NAND2_X1 U8455 ( .A1(n9691), .A2(n9699), .ZN(n9696) );
  NAND2_X1 U8456 ( .A1(n4631), .A2(n6776), .ZN(n9697) );
  NAND3_X1 U8457 ( .A1(n9668), .A2(n9696), .A3(n9697), .ZN(n6778) );
  NAND2_X1 U8458 ( .A1(n9669), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6777) );
  OAI211_X1 U8459 ( .C1(n9673), .C2(n9699), .A(n6778), .B(n6777), .ZN(n6779)
         );
  AOI21_X1 U8460 ( .B1(n9638), .B2(n9702), .A(n6779), .ZN(n6780) );
  OAI21_X1 U8461 ( .B1(n9669), .B2(n6781), .A(n6780), .ZN(P2_U3295) );
  XNOR2_X1 U8462 ( .A(n6783), .B(n6782), .ZN(n6789) );
  INV_X1 U8463 ( .A(n7150), .ZN(n6786) );
  AND2_X1 U8464 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9456) );
  AOI21_X1 U8465 ( .B1(n8881), .B2(n8865), .A(n9456), .ZN(n6785) );
  NAND2_X1 U8466 ( .A1(n8880), .A2(n8839), .ZN(n6784) );
  OAI211_X1 U8467 ( .C1(n8812), .C2(n6786), .A(n6785), .B(n6784), .ZN(n6787)
         );
  AOI21_X1 U8468 ( .B1(n7151), .B2(n8870), .A(n6787), .ZN(n6788) );
  OAI21_X1 U8469 ( .B1(n6789), .B2(n8872), .A(n6788), .ZN(P1_U3234) );
  OR2_X1 U8470 ( .A1(n6791), .A2(n6790), .ZN(n6794) );
  AND2_X1 U8471 ( .A1(n6794), .A2(n6792), .ZN(n6796) );
  NAND2_X1 U8472 ( .A1(n6794), .A2(n6793), .ZN(n6795) );
  OAI21_X1 U8473 ( .B1(n6796), .B2(n7796), .A(n6795), .ZN(n6797) );
  INV_X1 U8474 ( .A(n6797), .ZN(n6983) );
  NAND2_X1 U8475 ( .A1(n6555), .A2(n7601), .ZN(n6798) );
  NAND2_X1 U8476 ( .A1(n6798), .A2(n7602), .ZN(n6799) );
  XNOR2_X1 U8477 ( .A(n7796), .B(n6799), .ZN(n6800) );
  OAI222_X1 U8478 ( .A1(n9104), .A2(n6801), .B1(n5525), .B2(n7853), .C1(n6800), 
        .C2(n9256), .ZN(n6979) );
  INV_X1 U8479 ( .A(n6979), .ZN(n6802) );
  MUX2_X1 U8480 ( .A(n6803), .B(n6802), .S(n9081), .Z(n6809) );
  INV_X1 U8481 ( .A(n6911), .ZN(n6805) );
  AOI211_X1 U8482 ( .C1(n6981), .C2(n6805), .A(n9548), .B(n6804), .ZN(n6980)
         );
  INV_X1 U8483 ( .A(n7859), .ZN(n6806) );
  OAI22_X1 U8484 ( .A1(n9110), .A2(n7857), .B1(n6806), .B2(n9506), .ZN(n6807)
         );
  AOI21_X1 U8485 ( .B1(n6980), .B2(n9269), .A(n6807), .ZN(n6808) );
  OAI211_X1 U8486 ( .C1(n6983), .C2(n9114), .A(n6809), .B(n6808), .ZN(P1_U3284) );
  NAND2_X1 U8487 ( .A1(n7333), .A2(n7330), .ZN(n6810) );
  OAI211_X1 U8488 ( .C1(n10146), .C2(n8727), .A(n6810), .B(n8100), .ZN(
        P2_U3335) );
  NAND2_X1 U8489 ( .A1(n7333), .A2(n7259), .ZN(n6812) );
  OR2_X1 U8490 ( .A1(n6811), .A2(P1_U3084), .ZN(n7840) );
  OAI211_X1 U8491 ( .C1(n6813), .C2(n8103), .A(n6812), .B(n7840), .ZN(P1_U3330) );
  NAND2_X1 U8492 ( .A1(n6815), .A2(n6814), .ZN(n6817) );
  NAND2_X1 U8493 ( .A1(n6817), .A2(n6816), .ZN(n9674) );
  INV_X1 U8494 ( .A(n6818), .ZN(n9672) );
  NAND2_X1 U8495 ( .A1(n6819), .A2(n6818), .ZN(n7921) );
  NAND2_X1 U8496 ( .A1(n6820), .A2(n9672), .ZN(n7924) );
  NAND2_X1 U8497 ( .A1(n9674), .A2(n9675), .ZN(n6822) );
  OR2_X1 U8498 ( .A1(n8279), .A2(n9703), .ZN(n6821) );
  NAND2_X1 U8499 ( .A1(n6822), .A2(n6821), .ZN(n9641) );
  INV_X1 U8500 ( .A(n9709), .ZN(n6823) );
  NAND2_X1 U8501 ( .A1(n9641), .A2(n9643), .ZN(n6826) );
  NAND2_X1 U8502 ( .A1(n6824), .A2(n9709), .ZN(n6825) );
  NAND2_X1 U8503 ( .A1(n6826), .A2(n6825), .ZN(n9628) );
  NAND2_X1 U8504 ( .A1(n8277), .A2(n9717), .ZN(n9606) );
  NAND2_X1 U8505 ( .A1(n9628), .A2(n9629), .ZN(n6828) );
  INV_X1 U8506 ( .A(n9717), .ZN(n9630) );
  OR2_X1 U8507 ( .A1(n8277), .A2(n9630), .ZN(n6827) );
  NAND2_X1 U8508 ( .A1(n6828), .A2(n6827), .ZN(n9605) );
  INV_X1 U8509 ( .A(n9605), .ZN(n6829) );
  NAND2_X1 U8510 ( .A1(n8276), .A2(n4395), .ZN(n6830) );
  AND2_X1 U8511 ( .A1(n8275), .A2(n9583), .ZN(n6833) );
  INV_X1 U8512 ( .A(n9583), .ZN(n9730) );
  NAND2_X1 U8513 ( .A1(n9612), .A2(n9730), .ZN(n6832) );
  INV_X1 U8514 ( .A(n8274), .ZN(n6834) );
  INV_X1 U8515 ( .A(n7891), .ZN(n9736) );
  NAND2_X1 U8516 ( .A1(n6834), .A2(n9736), .ZN(n7938) );
  NAND2_X1 U8517 ( .A1(n8274), .A2(n7891), .ZN(n7937) );
  NAND2_X1 U8518 ( .A1(n7938), .A2(n7937), .ZN(n8061) );
  INV_X1 U8519 ( .A(n7039), .ZN(n6836) );
  XNOR2_X1 U8520 ( .A(n8273), .B(n7941), .ZN(n8063) );
  INV_X1 U8521 ( .A(n8272), .ZN(n6837) );
  NAND2_X1 U8522 ( .A1(n9750), .A2(n6837), .ZN(n7947) );
  NAND2_X1 U8523 ( .A1(n7948), .A2(n7947), .ZN(n6848) );
  NAND2_X1 U8524 ( .A1(n6838), .A2(n6848), .ZN(n6882) );
  OAI21_X1 U8525 ( .B1(n6838), .B2(n6848), .A(n6882), .ZN(n9760) );
  INV_X1 U8526 ( .A(n9760), .ZN(n9756) );
  NAND2_X1 U8527 ( .A1(n8056), .A2(n6839), .ZN(n7913) );
  NAND2_X1 U8528 ( .A1(n7913), .A2(n6840), .ZN(n7923) );
  INV_X1 U8529 ( .A(n9643), .ZN(n8059) );
  INV_X1 U8530 ( .A(n6841), .ZN(n7916) );
  AOI21_X1 U8531 ( .B1(n9642), .B2(n8059), .A(n7916), .ZN(n9623) );
  INV_X1 U8532 ( .A(n9629), .ZN(n6842) );
  NAND2_X1 U8533 ( .A1(n9623), .A2(n6842), .ZN(n9626) );
  NAND2_X1 U8534 ( .A1(n8276), .A2(n9725), .ZN(n8054) );
  NAND2_X1 U8535 ( .A1(n9626), .A2(n7929), .ZN(n6844) );
  INV_X1 U8536 ( .A(n8276), .ZN(n6843) );
  NAND2_X1 U8537 ( .A1(n6843), .A2(n4395), .ZN(n8055) );
  NAND2_X1 U8538 ( .A1(n6844), .A2(n8055), .ZN(n7875) );
  XNOR2_X1 U8539 ( .A(n8275), .B(n9583), .ZN(n8064) );
  NAND2_X1 U8540 ( .A1(n7875), .A2(n8064), .ZN(n6845) );
  NAND2_X1 U8541 ( .A1(n9612), .A2(n9583), .ZN(n7936) );
  NAND2_X1 U8542 ( .A1(n6845), .A2(n7936), .ZN(n7883) );
  INV_X1 U8543 ( .A(n7883), .ZN(n6847) );
  INV_X1 U8544 ( .A(n8061), .ZN(n6846) );
  INV_X1 U8545 ( .A(n8273), .ZN(n7942) );
  NAND2_X1 U8546 ( .A1(n7942), .A2(n7941), .ZN(n7944) );
  NAND2_X1 U8547 ( .A1(n7040), .A2(n7944), .ZN(n6884) );
  INV_X1 U8548 ( .A(n6848), .ZN(n8065) );
  XNOR2_X1 U8549 ( .A(n6884), .B(n8065), .ZN(n6849) );
  OAI22_X1 U8550 ( .A1(n7942), .A2(n9611), .B1(n6888), .B2(n9613), .ZN(n9570)
         );
  AOI21_X1 U8551 ( .B1(n6849), .B2(n9662), .A(n9570), .ZN(n9757) );
  MUX2_X1 U8552 ( .A(n9757), .B(n6850), .S(n9669), .Z(n6854) );
  NOR2_X1 U8553 ( .A1(n9696), .A2(n9703), .ZN(n9665) );
  NAND2_X1 U8554 ( .A1(n9665), .A2(n9709), .ZN(n9651) );
  INV_X1 U8555 ( .A(n7941), .ZN(n9744) );
  OR2_X1 U8556 ( .A1(n7045), .A2(n9750), .ZN(n6994) );
  INV_X1 U8557 ( .A(n6994), .ZN(n6851) );
  AOI21_X1 U8558 ( .B1(n9750), .B2(n7045), .A(n6851), .ZN(n9753) );
  INV_X1 U8559 ( .A(n9750), .ZN(n9574) );
  OAI22_X1 U8560 ( .A1(n9673), .A2(n9574), .B1(n9666), .B2(n9578), .ZN(n6852)
         );
  AOI21_X1 U8561 ( .B1(n9753), .B2(n9668), .A(n6852), .ZN(n6853) );
  OAI211_X1 U8562 ( .C1(n9676), .C2(n9756), .A(n6854), .B(n6853), .ZN(P2_U3287) );
  INV_X1 U8563 ( .A(n6855), .ZN(n6861) );
  OAI21_X1 U8564 ( .B1(n9506), .B2(n6857), .A(n6856), .ZN(n6860) );
  INV_X1 U8565 ( .A(n6858), .ZN(n6859) );
  AOI211_X1 U8566 ( .C1(n5543), .C2(n6861), .A(n6860), .B(n6859), .ZN(n6862)
         );
  MUX2_X1 U8567 ( .A(n6863), .B(n6862), .S(n9081), .Z(n6867) );
  INV_X1 U8568 ( .A(n9114), .ZN(n6864) );
  AOI22_X1 U8569 ( .A1(n6865), .A2(n6864), .B1(n9262), .B2(n5247), .ZN(n6866)
         );
  NAND2_X1 U8570 ( .A1(n6867), .A2(n6866), .ZN(P1_U3286) );
  OAI21_X1 U8571 ( .B1(n6869), .B2(n6675), .A(n6868), .ZN(n6873) );
  XNOR2_X1 U8572 ( .A(n6871), .B(n6870), .ZN(n6872) );
  XNOR2_X1 U8573 ( .A(n6873), .B(n6872), .ZN(n6879) );
  INV_X1 U8574 ( .A(n6874), .ZN(n6913) );
  AOI22_X1 U8575 ( .A1(n8870), .A2(n5527), .B1(n8883), .B2(n8839), .ZN(n6877)
         );
  AOI21_X1 U8576 ( .B1(n8885), .B2(n8865), .A(n6875), .ZN(n6876) );
  OAI211_X1 U8577 ( .C1(n8812), .C2(n6913), .A(n6877), .B(n6876), .ZN(n6878)
         );
  AOI21_X1 U8578 ( .B1(n6879), .B2(n8849), .A(n6878), .ZN(n6880) );
  INV_X1 U8579 ( .A(n6880), .ZN(P1_U3237) );
  OR2_X1 U8580 ( .A1(n9750), .A2(n8272), .ZN(n6881) );
  OR2_X1 U8581 ( .A1(n6998), .A2(n6888), .ZN(n7951) );
  NAND2_X1 U8582 ( .A1(n6998), .A2(n6888), .ZN(n7952) );
  INV_X1 U8583 ( .A(n6998), .ZN(n9763) );
  INV_X1 U8584 ( .A(n8270), .ZN(n6974) );
  NAND2_X1 U8585 ( .A1(n7026), .A2(n6974), .ZN(n7953) );
  NAND2_X1 U8586 ( .A1(n7961), .A2(n7953), .ZN(n8068) );
  OAI21_X1 U8587 ( .B1(n6883), .B2(n8068), .A(n7028), .ZN(n9769) );
  NAND2_X1 U8588 ( .A1(n6884), .A2(n8065), .ZN(n6885) );
  NAND2_X1 U8589 ( .A1(n7021), .A2(n7951), .ZN(n6886) );
  XOR2_X1 U8590 ( .A(n8068), .B(n6886), .Z(n6887) );
  OAI222_X1 U8591 ( .A1(n9613), .A2(n7082), .B1(n9611), .B2(n6888), .C1(n9644), 
        .C2(n6887), .ZN(n9772) );
  NAND2_X1 U8592 ( .A1(n9772), .A2(n9618), .ZN(n6894) );
  OAI22_X1 U8593 ( .A1(n9618), .A2(n6890), .B1(n6889), .B2(n9666), .ZN(n6892)
         );
  NOR2_X1 U8594 ( .A1(n6994), .A2(n6998), .ZN(n7031) );
  INV_X1 U8595 ( .A(n7026), .ZN(n9770) );
  XNOR2_X1 U8596 ( .A(n7031), .B(n9770), .ZN(n9771) );
  INV_X1 U8597 ( .A(n9668), .ZN(n9636) );
  NOR2_X1 U8598 ( .A1(n9771), .A2(n9636), .ZN(n6891) );
  AOI211_X1 U8599 ( .C1(n9631), .C2(n7026), .A(n6892), .B(n6891), .ZN(n6893)
         );
  OAI211_X1 U8600 ( .C1(n9676), .C2(n9769), .A(n6894), .B(n6893), .ZN(P2_U3285) );
  AND2_X1 U8601 ( .A1(n6897), .A2(n6895), .ZN(n6899) );
  NAND2_X1 U8602 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  OAI21_X1 U8603 ( .B1(n6899), .B2(n6901), .A(n6898), .ZN(n6900) );
  INV_X1 U8604 ( .A(n6900), .ZN(n9535) );
  INV_X1 U8605 ( .A(n6901), .ZN(n7658) );
  NAND2_X1 U8606 ( .A1(n6903), .A2(n7658), .ZN(n7626) );
  OAI21_X1 U8607 ( .B1(n7658), .B2(n6903), .A(n7626), .ZN(n6909) );
  OAI22_X1 U8608 ( .A1(n6905), .A2(n5525), .B1(n6904), .B2(n9104), .ZN(n6908)
         );
  NOR2_X1 U8609 ( .A1(n9535), .A2(n6906), .ZN(n6907) );
  AOI211_X1 U8610 ( .C1(n9065), .C2(n6909), .A(n6908), .B(n6907), .ZN(n9533)
         );
  MUX2_X1 U8611 ( .A(n6910), .B(n9533), .S(n5603), .Z(n6917) );
  AOI21_X1 U8612 ( .B1(n5527), .B2(n6912), .A(n6911), .ZN(n9531) );
  OAI22_X1 U8613 ( .A1(n9110), .A2(n6914), .B1(n6913), .B2(n9506), .ZN(n6915)
         );
  AOI21_X1 U8614 ( .B1(n9531), .B2(n9068), .A(n6915), .ZN(n6916) );
  OAI211_X1 U8615 ( .C1(n9535), .C2(n6918), .A(n6917), .B(n6916), .ZN(P1_U3285) );
  NAND2_X1 U8616 ( .A1(n6920), .A2(n6923), .ZN(n6921) );
  INV_X1 U8617 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U8618 ( .A1(n9472), .A2(n9471), .ZN(n9470) );
  NAND2_X1 U8619 ( .A1(n6921), .A2(n9470), .ZN(n7156) );
  XNOR2_X1 U8620 ( .A(n7156), .B(n7163), .ZN(n6922) );
  INV_X1 U8621 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U8622 ( .A1(n9943), .A2(n6922), .ZN(n7157) );
  AOI211_X1 U8623 ( .C1(n6922), .C2(n9943), .A(n7157), .B(n9488), .ZN(n6934)
         );
  INV_X1 U8624 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9349) );
  AOI22_X1 U8625 ( .A1(n9469), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9349), .B2(
        n6923), .ZN(n9475) );
  OAI21_X1 U8626 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6925), .A(n6924), .ZN(
        n9474) );
  NAND2_X1 U8627 ( .A1(n9475), .A2(n9474), .ZN(n9473) );
  OAI21_X1 U8628 ( .B1(n9469), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9473), .ZN(
        n7162) );
  XNOR2_X1 U8629 ( .A(n7162), .B(n7163), .ZN(n6927) );
  INV_X1 U8630 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U8631 ( .A1(n6926), .A2(n6927), .ZN(n7164) );
  AOI211_X1 U8632 ( .C1(n6927), .C2(n6926), .A(n7164), .B(n9381), .ZN(n6933)
         );
  INV_X1 U8633 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6931) );
  NOR2_X1 U8634 ( .A1(n6928), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8864) );
  AOI21_X1 U8635 ( .B1(n9483), .B2(n6929), .A(n8864), .ZN(n6930) );
  OAI21_X1 U8636 ( .B1(n9481), .B2(n6931), .A(n6930), .ZN(n6932) );
  OR3_X1 U8637 ( .A1(n6934), .A2(n6933), .A3(n6932), .ZN(P1_U3256) );
  NAND2_X1 U8638 ( .A1(n6675), .A2(n6935), .ZN(n7850) );
  NAND2_X1 U8639 ( .A1(n7850), .A2(n6937), .ZN(n6938) );
  AND2_X1 U8640 ( .A1(n6938), .A2(n7847), .ZN(n6941) );
  OR2_X1 U8641 ( .A1(n6941), .A2(n6940), .ZN(n7010) );
  NAND2_X1 U8642 ( .A1(n7010), .A2(n6939), .ZN(n7005) );
  NAND2_X1 U8643 ( .A1(n6941), .A2(n6940), .ZN(n7007) );
  NAND2_X1 U8644 ( .A1(n7005), .A2(n7007), .ZN(n7004) );
  XNOR2_X1 U8645 ( .A(n6943), .B(n6942), .ZN(n6944) );
  XNOR2_X1 U8646 ( .A(n7004), .B(n6944), .ZN(n6951) );
  NAND2_X1 U8647 ( .A1(n8863), .A2(n6945), .ZN(n6947) );
  AND2_X1 U8648 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9439) );
  AOI21_X1 U8649 ( .B1(n8882), .B2(n8865), .A(n9439), .ZN(n6946) );
  OAI211_X1 U8650 ( .C1(n7144), .C2(n8868), .A(n6947), .B(n6946), .ZN(n6948)
         );
  AOI21_X1 U8651 ( .B1(n6949), .B2(n8870), .A(n6948), .ZN(n6950) );
  OAI21_X1 U8652 ( .B1(n6951), .B2(n8872), .A(n6950), .ZN(P1_U3229) );
  NAND2_X1 U8653 ( .A1(n6952), .A2(n7907), .ZN(n6955) );
  AOI22_X1 U8654 ( .A1(n7370), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7369), .B2(
        n6953), .ZN(n6954) );
  NAND2_X1 U8655 ( .A1(n6955), .A2(n6954), .ZN(n7073) );
  INV_X1 U8656 ( .A(n7073), .ZN(n9777) );
  AND2_X1 U8657 ( .A1(n8140), .A2(n8269), .ZN(n6957) );
  XNOR2_X1 U8658 ( .A(n7073), .B(n8179), .ZN(n6956) );
  NOR2_X1 U8659 ( .A1(n6956), .A2(n6957), .ZN(n7054) );
  AOI21_X1 U8660 ( .B1(n6957), .B2(n6956), .A(n7054), .ZN(n6964) );
  INV_X1 U8661 ( .A(n6958), .ZN(n6960) );
  OAI21_X1 U8662 ( .B1(n6964), .B2(n6963), .A(n7056), .ZN(n6965) );
  NAND2_X1 U8663 ( .A1(n6965), .A2(n9589), .ZN(n6978) );
  INV_X1 U8664 ( .A(n6966), .ZN(n7033) );
  INV_X1 U8665 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8666 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  NAND2_X1 U8667 ( .A1(n7062), .A2(n6969), .ZN(n7086) );
  OR2_X1 U8668 ( .A1(n7480), .A2(n7086), .ZN(n6973) );
  NAND2_X1 U8669 ( .A1(n7489), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8670 ( .A1(n7488), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8671 ( .A1(n7490), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6970) );
  NAND4_X1 U8672 ( .A1(n6973), .A2(n6972), .A3(n6971), .A4(n6970), .ZN(n8268)
         );
  INV_X1 U8673 ( .A(n8268), .ZN(n7965) );
  OAI22_X1 U8674 ( .A1(n6974), .A2(n8245), .B1(n8244), .B2(n7965), .ZN(n6975)
         );
  AOI211_X1 U8675 ( .C1(n7033), .C2(n8258), .A(n6976), .B(n6975), .ZN(n6977)
         );
  OAI211_X1 U8676 ( .C1(n9777), .C2(n9573), .A(n6978), .B(n6977), .ZN(P2_U3226) );
  AOI211_X1 U8677 ( .C1(n9529), .C2(n6981), .A(n6980), .B(n6979), .ZN(n6982)
         );
  OAI21_X1 U8678 ( .B1(n9198), .B2(n6983), .A(n6982), .ZN(n6986) );
  NAND2_X1 U8679 ( .A1(n6986), .A2(n9565), .ZN(n6984) );
  OAI21_X1 U8680 ( .B1(n9565), .B2(n6985), .A(n6984), .ZN(P1_U3530) );
  INV_X1 U8681 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U8682 ( .A1(n6986), .A2(n9556), .ZN(n6987) );
  OAI21_X1 U8683 ( .B1(n9556), .B2(n10125), .A(n6987), .ZN(P1_U3475) );
  INV_X1 U8684 ( .A(n7404), .ZN(n7052) );
  OAI222_X1 U8685 ( .A1(n4396), .A2(n7052), .B1(P1_U3084), .B2(n6989), .C1(
        n6988), .C2(n8108), .ZN(P1_U3329) );
  XNOR2_X1 U8686 ( .A(n6990), .B(n8067), .ZN(n9767) );
  INV_X1 U8687 ( .A(n9767), .ZN(n7003) );
  OAI211_X1 U8688 ( .C1(n4477), .C2(n6991), .A(n9662), .B(n7021), .ZN(n6993)
         );
  NAND2_X1 U8689 ( .A1(n6993), .A2(n6992), .ZN(n9765) );
  AND2_X1 U8690 ( .A1(n6994), .A2(n6998), .ZN(n6995) );
  OR2_X1 U8691 ( .A1(n6995), .A2(n7031), .ZN(n9764) );
  NOR2_X1 U8692 ( .A1(n9666), .A2(n6996), .ZN(n6997) );
  AOI21_X1 U8693 ( .B1(n9669), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6997), .ZN(
        n7000) );
  NAND2_X1 U8694 ( .A1(n9631), .A2(n6998), .ZN(n6999) );
  OAI211_X1 U8695 ( .C1(n9764), .C2(n9636), .A(n7000), .B(n6999), .ZN(n7001)
         );
  AOI21_X1 U8696 ( .B1(n9765), .B2(n9618), .A(n7001), .ZN(n7002) );
  OAI21_X1 U8697 ( .B1(n9676), .B2(n7003), .A(n7002), .ZN(P2_U3286) );
  INV_X1 U8698 ( .A(n7004), .ZN(n7011) );
  INV_X1 U8699 ( .A(n7005), .ZN(n7008) );
  AOI21_X1 U8700 ( .B1(n7008), .B2(n7007), .A(n7006), .ZN(n7009) );
  AOI21_X1 U8701 ( .B1(n7011), .B2(n7010), .A(n7009), .ZN(n7020) );
  INV_X1 U8702 ( .A(n7012), .ZN(n7016) );
  AOI21_X1 U8703 ( .B1(n8883), .B2(n8865), .A(n7013), .ZN(n7015) );
  NAND2_X1 U8704 ( .A1(n8839), .A2(n9253), .ZN(n7014) );
  OAI211_X1 U8705 ( .C1(n8812), .C2(n7016), .A(n7015), .B(n7014), .ZN(n7017)
         );
  AOI21_X1 U8706 ( .B1(n7018), .B2(n8870), .A(n7017), .ZN(n7019) );
  OAI21_X1 U8707 ( .B1(n7020), .B2(n8872), .A(n7019), .ZN(P1_U3219) );
  AND2_X1 U8708 ( .A1(n7961), .A2(n7951), .ZN(n7955) );
  NAND2_X1 U8709 ( .A1(n7080), .A2(n7953), .ZN(n7022) );
  OR2_X1 U8710 ( .A1(n7073), .A2(n7082), .ZN(n7957) );
  NAND2_X1 U8711 ( .A1(n7073), .A2(n7082), .ZN(n7963) );
  XNOR2_X1 U8712 ( .A(n7022), .B(n8072), .ZN(n7023) );
  NAND2_X1 U8713 ( .A1(n7023), .A2(n9662), .ZN(n7025) );
  AOI22_X1 U8714 ( .A1(n8571), .A2(n8270), .B1(n8268), .B2(n8573), .ZN(n7024)
         );
  NAND2_X1 U8715 ( .A1(n7025), .A2(n7024), .ZN(n9780) );
  INV_X1 U8716 ( .A(n9780), .ZN(n7038) );
  NAND2_X1 U8717 ( .A1(n7026), .A2(n8270), .ZN(n7027) );
  INV_X1 U8718 ( .A(n8072), .ZN(n7029) );
  OAI21_X1 U8719 ( .B1(n7030), .B2(n7029), .A(n7074), .ZN(n9782) );
  AND2_X1 U8720 ( .A1(n7031), .A2(n9770), .ZN(n7032) );
  NAND2_X1 U8721 ( .A1(n7032), .A2(n9777), .ZN(n7087) );
  OAI21_X1 U8722 ( .B1(n7032), .B2(n9777), .A(n7087), .ZN(n9779) );
  AOI22_X1 U8723 ( .A1(n9669), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7033), .B2(
        n9632), .ZN(n7035) );
  NAND2_X1 U8724 ( .A1(n9631), .A2(n7073), .ZN(n7034) );
  OAI211_X1 U8725 ( .C1(n9779), .C2(n9636), .A(n7035), .B(n7034), .ZN(n7036)
         );
  AOI21_X1 U8726 ( .B1(n9782), .B2(n9638), .A(n7036), .ZN(n7037) );
  OAI21_X1 U8727 ( .B1(n9669), .B2(n7038), .A(n7037), .ZN(P2_U3284) );
  XNOR2_X1 U8728 ( .A(n7039), .B(n6835), .ZN(n9748) );
  INV_X1 U8729 ( .A(n9748), .ZN(n7051) );
  INV_X1 U8730 ( .A(n7040), .ZN(n7041) );
  AOI21_X1 U8731 ( .B1(n6835), .B2(n7042), .A(n7041), .ZN(n7044) );
  OAI21_X1 U8732 ( .B1(n7044), .B2(n9644), .A(n7043), .ZN(n9746) );
  OAI21_X1 U8733 ( .B1(n7888), .B2(n9744), .A(n7045), .ZN(n9745) );
  OAI22_X1 U8734 ( .A1(n9618), .A2(n6279), .B1(n7046), .B2(n9666), .ZN(n7047)
         );
  AOI21_X1 U8735 ( .B1(n9631), .B2(n7941), .A(n7047), .ZN(n7048) );
  OAI21_X1 U8736 ( .B1(n9636), .B2(n9745), .A(n7048), .ZN(n7049) );
  AOI21_X1 U8737 ( .B1(n9746), .B2(n9618), .A(n7049), .ZN(n7050) );
  OAI21_X1 U8738 ( .B1(n9676), .B2(n7051), .A(n7050), .ZN(P2_U3288) );
  OAI222_X1 U8739 ( .A1(n7053), .A2(P2_U3152), .B1(n7895), .B2(n7052), .C1(
        n7405), .C2(n8727), .ZN(P2_U3334) );
  INV_X1 U8740 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U8741 ( .A1(n7057), .A2(n7907), .ZN(n7060) );
  AOI22_X1 U8742 ( .A1(n7370), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7369), .B2(
        n7058), .ZN(n7059) );
  XNOR2_X1 U8743 ( .A(n9325), .B(n8179), .ZN(n7228) );
  NAND2_X1 U8744 ( .A1(n8268), .A2(n8140), .ZN(n7227) );
  XNOR2_X1 U8745 ( .A(n7228), .B(n7227), .ZN(n7230) );
  XNOR2_X1 U8746 ( .A(n7231), .B(n7230), .ZN(n7072) );
  INV_X1 U8747 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8748 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  NAND2_X1 U8749 ( .A1(n7104), .A2(n7063), .ZN(n7112) );
  OR2_X1 U8750 ( .A1(n7480), .A2(n7112), .ZN(n7067) );
  NAND2_X1 U8751 ( .A1(n7459), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8752 ( .A1(n7488), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8753 ( .A1(n7490), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7064) );
  NAND4_X1 U8754 ( .A1(n7067), .A2(n7066), .A3(n7065), .A4(n7064), .ZN(n8267)
         );
  AOI22_X1 U8755 ( .A1(n8187), .A2(n8269), .B1(n8188), .B2(n8267), .ZN(n7069)
         );
  OAI211_X1 U8756 ( .C1(n9593), .C2(n7086), .A(n7069), .B(n7068), .ZN(n7070)
         );
  AOI21_X1 U8757 ( .B1(n9584), .B2(n9325), .A(n7070), .ZN(n7071) );
  OAI21_X1 U8758 ( .B1(n7072), .B2(n8250), .A(n7071), .ZN(P2_U3236) );
  XNOR2_X1 U8759 ( .A(n9325), .B(n8268), .ZN(n8070) );
  NAND2_X1 U8760 ( .A1(n7075), .A2(n8070), .ZN(n7076) );
  NAND2_X1 U8761 ( .A1(n7077), .A2(n7076), .ZN(n9324) );
  OR2_X1 U8762 ( .A1(n9669), .A2(n7078), .ZN(n9648) );
  AND2_X1 U8763 ( .A1(n7963), .A2(n7953), .ZN(n7958) );
  INV_X1 U8764 ( .A(n7957), .ZN(n7079) );
  INV_X1 U8765 ( .A(n8070), .ZN(n7966) );
  NAND2_X1 U8766 ( .A1(n7081), .A2(n8070), .ZN(n7101) );
  OAI21_X1 U8767 ( .B1(n7081), .B2(n8070), .A(n7101), .ZN(n7084) );
  INV_X1 U8768 ( .A(n8267), .ZN(n7244) );
  OAI22_X1 U8769 ( .A1(n7082), .A2(n9611), .B1(n7244), .B2(n9613), .ZN(n7083)
         );
  AOI21_X1 U8770 ( .B1(n7084), .B2(n9662), .A(n7083), .ZN(n7085) );
  OAI21_X1 U8771 ( .B1(n9324), .B2(n9640), .A(n7085), .ZN(n9328) );
  NAND2_X1 U8772 ( .A1(n9328), .A2(n9618), .ZN(n7092) );
  OAI22_X1 U8773 ( .A1(n9618), .A2(n6628), .B1(n7086), .B2(n9666), .ZN(n7090)
         );
  NAND2_X1 U8774 ( .A1(n7087), .A2(n9325), .ZN(n7088) );
  NAND2_X1 U8775 ( .A1(n7198), .A2(n7088), .ZN(n9327) );
  NOR2_X1 U8776 ( .A1(n9327), .A2(n9636), .ZN(n7089) );
  AOI211_X1 U8777 ( .C1(n9631), .C2(n9325), .A(n7090), .B(n7089), .ZN(n7091)
         );
  OAI211_X1 U8778 ( .C1(n9324), .C2(n9648), .A(n7092), .B(n7091), .ZN(P2_U3283) );
  NAND2_X1 U8779 ( .A1(n7094), .A2(n7907), .ZN(n7096) );
  AOI22_X1 U8780 ( .A1(n7370), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7369), .B2(
        n8322), .ZN(n7095) );
  NAND2_X1 U8781 ( .A1(n7222), .A2(n7244), .ZN(n7970) );
  NAND2_X1 U8782 ( .A1(n7971), .A2(n7970), .ZN(n8053) );
  NAND2_X1 U8783 ( .A1(n7097), .A2(n8053), .ZN(n7182) );
  OAI21_X1 U8784 ( .B1(n7097), .B2(n8053), .A(n7182), .ZN(n9322) );
  INV_X1 U8785 ( .A(n9322), .ZN(n7117) );
  AND2_X1 U8786 ( .A1(n9325), .A2(n7965), .ZN(n7959) );
  INV_X1 U8787 ( .A(n7959), .ZN(n7098) );
  NAND2_X1 U8788 ( .A1(n7101), .A2(n7098), .ZN(n7099) );
  NAND2_X1 U8789 ( .A1(n7099), .A2(n8053), .ZN(n7102) );
  NOR2_X1 U8790 ( .A1(n8053), .A2(n7959), .ZN(n7100) );
  NAND3_X1 U8791 ( .A1(n7102), .A2(n7186), .A3(n9662), .ZN(n7111) );
  INV_X1 U8792 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U8793 ( .A1(n7104), .A2(n8327), .ZN(n7105) );
  NAND2_X1 U8794 ( .A1(n7190), .A2(n7105), .ZN(n7243) );
  OR2_X1 U8795 ( .A1(n7480), .A2(n7243), .ZN(n7109) );
  NAND2_X1 U8796 ( .A1(n7490), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8797 ( .A1(n7489), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U8798 ( .A1(n7488), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7106) );
  NAND4_X1 U8799 ( .A1(n7109), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n8266)
         );
  AOI22_X1 U8800 ( .A1(n8571), .A2(n8268), .B1(n8266), .B2(n8573), .ZN(n7110)
         );
  NAND2_X1 U8801 ( .A1(n7111), .A2(n7110), .ZN(n9321) );
  XNOR2_X1 U8802 ( .A(n7198), .B(n7222), .ZN(n9319) );
  INV_X1 U8803 ( .A(n7112), .ZN(n7237) );
  AOI22_X1 U8804 ( .A1(n9669), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7237), .B2(
        n9632), .ZN(n7114) );
  NAND2_X1 U8805 ( .A1(n7222), .A2(n9631), .ZN(n7113) );
  OAI211_X1 U8806 ( .C1(n9319), .C2(n9636), .A(n7114), .B(n7113), .ZN(n7115)
         );
  AOI21_X1 U8807 ( .B1(n9321), .B2(n9618), .A(n7115), .ZN(n7116) );
  OAI21_X1 U8808 ( .B1(n7117), .B2(n9676), .A(n7116), .ZN(P2_U3282) );
  INV_X1 U8809 ( .A(n7120), .ZN(n7121) );
  AOI21_X1 U8810 ( .B1(n7122), .B2(n7119), .A(n7121), .ZN(n7129) );
  NAND2_X1 U8811 ( .A1(n8863), .A2(n7214), .ZN(n7125) );
  AOI21_X1 U8812 ( .B1(n9252), .B2(n8865), .A(n7123), .ZN(n7124) );
  OAI211_X1 U8813 ( .C1(n7126), .C2(n8868), .A(n7125), .B(n7124), .ZN(n7127)
         );
  AOI21_X1 U8814 ( .B1(n7215), .B2(n8870), .A(n7127), .ZN(n7128) );
  OAI21_X1 U8815 ( .B1(n7129), .B2(n8872), .A(n7128), .ZN(P1_U3222) );
  INV_X1 U8816 ( .A(n7130), .ZN(n7132) );
  NOR2_X1 U8817 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  XNOR2_X1 U8818 ( .A(n4472), .B(n7133), .ZN(n7140) );
  INV_X1 U8819 ( .A(n7275), .ZN(n7137) );
  AOI21_X1 U8820 ( .B1(n8880), .B2(n8865), .A(n7134), .ZN(n7136) );
  NAND2_X1 U8821 ( .A1(n8839), .A2(n8878), .ZN(n7135) );
  OAI211_X1 U8822 ( .C1(n8812), .C2(n7137), .A(n7136), .B(n7135), .ZN(n7138)
         );
  AOI21_X1 U8823 ( .B1(n7276), .B2(n8870), .A(n7138), .ZN(n7139) );
  OAI21_X1 U8824 ( .B1(n7140), .B2(n8872), .A(n7139), .ZN(P1_U3232) );
  XNOR2_X1 U8825 ( .A(n7151), .B(n9252), .ZN(n7805) );
  INV_X1 U8826 ( .A(n7805), .ZN(n7643) );
  XNOR2_X1 U8827 ( .A(n7141), .B(n7643), .ZN(n7252) );
  XNOR2_X1 U8828 ( .A(n7142), .B(n7805), .ZN(n7147) );
  OAI22_X1 U8829 ( .A1(n7144), .A2(n5525), .B1(n7143), .B2(n9104), .ZN(n7145)
         );
  INV_X1 U8830 ( .A(n7145), .ZN(n7146) );
  OAI21_X1 U8831 ( .B1(n7147), .B2(n9256), .A(n7146), .ZN(n7148) );
  AOI21_X1 U8832 ( .B1(n7252), .B2(n9259), .A(n7148), .ZN(n7254) );
  NOR2_X1 U8833 ( .A1(n9265), .A2(n7249), .ZN(n7149) );
  OR2_X1 U8834 ( .A1(n7213), .A2(n7149), .ZN(n7250) );
  AOI22_X1 U8835 ( .A1(n9513), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7150), .B2(
        n9261), .ZN(n7153) );
  NAND2_X1 U8836 ( .A1(n9262), .A2(n7151), .ZN(n7152) );
  OAI211_X1 U8837 ( .C1(n7250), .C2(n7528), .A(n7153), .B(n7152), .ZN(n7154)
         );
  AOI21_X1 U8838 ( .B1(n7252), .B2(n4394), .A(n7154), .ZN(n7155) );
  OAI21_X1 U8839 ( .B1(n7254), .B2(n9513), .A(n7155), .ZN(P1_U3280) );
  NOR2_X1 U8840 ( .A1(n7163), .A2(n7156), .ZN(n7158) );
  NAND2_X1 U8841 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7538), .ZN(n7159) );
  OAI21_X1 U8842 ( .B1(n7538), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7159), .ZN(
        n7160) );
  AOI211_X1 U8843 ( .C1(n7161), .C2(n7160), .A(n7530), .B(n9488), .ZN(n7173)
         );
  NOR2_X1 U8844 ( .A1(n7163), .A2(n7162), .ZN(n7165) );
  NOR2_X1 U8845 ( .A1(n7165), .A2(n7164), .ZN(n7167) );
  XNOR2_X1 U8846 ( .A(n7538), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7166) );
  NOR2_X1 U8847 ( .A1(n7167), .A2(n7166), .ZN(n7537) );
  AOI211_X1 U8848 ( .C1(n7167), .C2(n7166), .A(n7537), .B(n9381), .ZN(n7172)
         );
  NAND2_X1 U8849 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7169) );
  NAND2_X1 U8850 ( .A1(n9495), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7168) );
  OAI211_X1 U8851 ( .C1(n9408), .C2(n7170), .A(n7169), .B(n7168), .ZN(n7171)
         );
  OR3_X1 U8852 ( .A1(n7173), .A2(n7172), .A3(n7171), .ZN(P1_U3257) );
  INV_X1 U8853 ( .A(n7415), .ZN(n7177) );
  INV_X1 U8854 ( .A(n7174), .ZN(n7175) );
  OAI222_X1 U8855 ( .A1(n8727), .A2(n7416), .B1(n7895), .B2(n7177), .C1(n7175), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U8856 ( .A1(n8108), .A2(n7178), .B1(n4396), .B2(n7177), .C1(n7176), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U8857 ( .A(n7426), .ZN(n7220) );
  OAI222_X1 U8858 ( .A1(n4396), .A2(n7220), .B1(P1_U3084), .B2(n7180), .C1(
        n7179), .C2(n8103), .ZN(P1_U3327) );
  OR2_X1 U8859 ( .A1(n7222), .A2(n8267), .ZN(n7181) );
  NAND2_X1 U8860 ( .A1(n7182), .A2(n7181), .ZN(n7366) );
  NAND2_X1 U8861 ( .A1(n7183), .A2(n7907), .ZN(n7185) );
  AOI22_X1 U8862 ( .A1(n7370), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7369), .B2(
        n8342), .ZN(n7184) );
  INV_X1 U8863 ( .A(n8266), .ZN(n8599) );
  NAND2_X1 U8864 ( .A1(n7364), .A2(n8599), .ZN(n7976) );
  NAND2_X1 U8865 ( .A1(n7975), .A2(n7976), .ZN(n8075) );
  XNOR2_X1 U8866 ( .A(n7366), .B(n8075), .ZN(n9316) );
  INV_X1 U8867 ( .A(n9316), .ZN(n7206) );
  XNOR2_X1 U8868 ( .A(n7494), .B(n8075), .ZN(n7187) );
  NAND2_X1 U8869 ( .A1(n7187), .A2(n9662), .ZN(n7197) );
  INV_X1 U8870 ( .A(n7190), .ZN(n7188) );
  INV_X1 U8871 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7189) );
  NAND2_X1 U8872 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  NAND2_X1 U8873 ( .A1(n7319), .A2(n7191), .ZN(n8608) );
  OR2_X1 U8874 ( .A1(n7480), .A2(n8608), .ZN(n7195) );
  NAND2_X1 U8875 ( .A1(n7489), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8876 ( .A1(n7490), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8877 ( .A1(n7488), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7192) );
  NAND4_X1 U8878 ( .A1(n7195), .A2(n7194), .A3(n7193), .A4(n7192), .ZN(n8265)
         );
  AOI22_X1 U8879 ( .A1(n8571), .A2(n8267), .B1(n8265), .B2(n8573), .ZN(n7196)
         );
  NAND2_X1 U8880 ( .A1(n7197), .A2(n7196), .ZN(n9315) );
  INV_X1 U8881 ( .A(n7364), .ZN(n9312) );
  OR2_X1 U8882 ( .A1(n7199), .A2(n9312), .ZN(n7200) );
  NAND2_X1 U8883 ( .A1(n8610), .A2(n7200), .ZN(n9313) );
  NAND2_X1 U8884 ( .A1(n9669), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7201) );
  OAI21_X1 U8885 ( .B1(n9666), .B2(n7243), .A(n7201), .ZN(n7202) );
  AOI21_X1 U8886 ( .B1(n7364), .B2(n9631), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8887 ( .B1(n9313), .B2(n9636), .A(n7203), .ZN(n7204) );
  AOI21_X1 U8888 ( .B1(n9315), .B2(n9618), .A(n7204), .ZN(n7205) );
  OAI21_X1 U8889 ( .B1(n7206), .B2(n9676), .A(n7205), .ZN(P2_U3281) );
  INV_X1 U8890 ( .A(n7207), .ZN(n7806) );
  XNOR2_X1 U8891 ( .A(n7208), .B(n7806), .ZN(n9359) );
  XNOR2_X1 U8892 ( .A(n7209), .B(n7806), .ZN(n7211) );
  AOI22_X1 U8893 ( .A1(n9254), .A2(n9252), .B1(n8879), .B2(n9251), .ZN(n7210)
         );
  OAI21_X1 U8894 ( .B1(n7211), .B2(n9256), .A(n7210), .ZN(n7212) );
  AOI21_X1 U8895 ( .B1(n9359), .B2(n9259), .A(n7212), .ZN(n9361) );
  OAI211_X1 U8896 ( .C1(n7213), .C2(n9357), .A(n9530), .B(n7273), .ZN(n9356)
         );
  AOI22_X1 U8897 ( .A1(n9513), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7214), .B2(
        n9261), .ZN(n7217) );
  NAND2_X1 U8898 ( .A1(n9262), .A2(n7215), .ZN(n7216) );
  OAI211_X1 U8899 ( .C1(n9356), .C2(n7301), .A(n7217), .B(n7216), .ZN(n7218)
         );
  AOI21_X1 U8900 ( .B1(n9359), .B2(n4394), .A(n7218), .ZN(n7219) );
  OAI21_X1 U8901 ( .B1(n9361), .B2(n9513), .A(n7219), .ZN(P1_U3279) );
  OAI222_X1 U8902 ( .A1(n7221), .A2(P2_U3152), .B1(n7895), .B2(n7220), .C1(
        n7427), .C2(n8727), .ZN(P2_U3332) );
  INV_X1 U8903 ( .A(n7222), .ZN(n9318) );
  NAND2_X1 U8904 ( .A1(n8267), .A2(n8140), .ZN(n7223) );
  INV_X1 U8905 ( .A(n7223), .ZN(n7226) );
  XNOR2_X1 U8906 ( .A(n7222), .B(n8145), .ZN(n7224) );
  INV_X1 U8907 ( .A(n7224), .ZN(n7225) );
  AOI21_X1 U8908 ( .B1(n7226), .B2(n7225), .A(n7310), .ZN(n7233) );
  INV_X1 U8909 ( .A(n7227), .ZN(n7229) );
  OAI21_X1 U8910 ( .B1(n7233), .B2(n7232), .A(n7316), .ZN(n7234) );
  NAND2_X1 U8911 ( .A1(n7234), .A2(n9589), .ZN(n7239) );
  OAI22_X1 U8912 ( .A1(n7965), .A2(n8245), .B1(n8244), .B2(n8599), .ZN(n7235)
         );
  AOI211_X1 U8913 ( .C1(n7237), .C2(n8258), .A(n7236), .B(n7235), .ZN(n7238)
         );
  OAI211_X1 U8914 ( .C1(n9318), .C2(n9573), .A(n7239), .B(n7238), .ZN(P2_U3217) );
  INV_X1 U8915 ( .A(n7310), .ZN(n7240) );
  NAND2_X1 U8916 ( .A1(n7316), .A2(n7240), .ZN(n7242) );
  XNOR2_X1 U8917 ( .A(n7364), .B(n8145), .ZN(n7311) );
  NAND2_X1 U8918 ( .A1(n8266), .A2(n8140), .ZN(n7312) );
  XNOR2_X1 U8919 ( .A(n7311), .B(n7312), .ZN(n7241) );
  XNOR2_X1 U8920 ( .A(n7242), .B(n7241), .ZN(n7248) );
  OAI22_X1 U8921 ( .A1(n9593), .A2(n7243), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8327), .ZN(n7246) );
  INV_X1 U8922 ( .A(n8265), .ZN(n8592) );
  OAI22_X1 U8923 ( .A1(n7244), .A2(n8245), .B1(n8244), .B2(n8592), .ZN(n7245)
         );
  AOI211_X1 U8924 ( .C1(n9584), .C2(n7364), .A(n7246), .B(n7245), .ZN(n7247)
         );
  OAI21_X1 U8925 ( .B1(n7248), .B2(n8250), .A(n7247), .ZN(P2_U3243) );
  OAI22_X1 U8926 ( .A1(n7250), .A2(n9548), .B1(n7249), .B2(n9546), .ZN(n7251)
         );
  AOI21_X1 U8927 ( .B1(n7252), .B2(n9553), .A(n7251), .ZN(n7253) );
  AND2_X1 U8928 ( .A1(n7254), .A2(n7253), .ZN(n7256) );
  MUX2_X1 U8929 ( .A(n6182), .B(n7256), .S(n9565), .Z(n7255) );
  INV_X1 U8930 ( .A(n7255), .ZN(P1_U3534) );
  INV_X1 U8931 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7257) );
  MUX2_X1 U8932 ( .A(n7257), .B(n7256), .S(n9556), .Z(n7258) );
  INV_X1 U8933 ( .A(n7258), .ZN(P1_U3487) );
  NAND2_X1 U8934 ( .A1(n7440), .A2(n7259), .ZN(n7261) );
  OAI211_X1 U8935 ( .C1(n8103), .C2(n7262), .A(n7261), .B(n7260), .ZN(P1_U3326) );
  INV_X1 U8936 ( .A(n7440), .ZN(n7263) );
  OAI222_X1 U8937 ( .A1(n8727), .A2(n7441), .B1(n7895), .B2(n7263), .C1(n8095), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U8938 ( .A(n7807), .ZN(n7264) );
  XNOR2_X1 U8939 ( .A(n7265), .B(n7264), .ZN(n9353) );
  NAND2_X1 U8940 ( .A1(n7266), .A2(n7635), .ZN(n7268) );
  NAND2_X1 U8941 ( .A1(n7268), .A2(n7807), .ZN(n7267) );
  OAI21_X1 U8942 ( .B1(n7807), .B2(n7268), .A(n7267), .ZN(n7269) );
  NAND2_X1 U8943 ( .A1(n7269), .A2(n9065), .ZN(n7271) );
  AOI22_X1 U8944 ( .A1(n8880), .A2(n9254), .B1(n9251), .B2(n8878), .ZN(n7270)
         );
  NAND2_X1 U8945 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  AOI21_X1 U8946 ( .B1(n9353), .B2(n9259), .A(n7272), .ZN(n9355) );
  NAND2_X1 U8947 ( .A1(n7273), .A2(n7276), .ZN(n7274) );
  NAND2_X1 U8948 ( .A1(n7296), .A2(n7274), .ZN(n9351) );
  AOI22_X1 U8949 ( .A1(n9513), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7275), .B2(
        n9261), .ZN(n7278) );
  NAND2_X1 U8950 ( .A1(n7276), .A2(n9262), .ZN(n7277) );
  OAI211_X1 U8951 ( .C1(n9351), .C2(n7528), .A(n7278), .B(n7277), .ZN(n7279)
         );
  AOI21_X1 U8952 ( .B1(n9353), .B2(n4394), .A(n7279), .ZN(n7280) );
  OAI21_X1 U8953 ( .B1(n9355), .B2(n9513), .A(n7280), .ZN(P1_U3278) );
  INV_X1 U8954 ( .A(n7281), .ZN(n7282) );
  NOR2_X1 U8955 ( .A1(n7283), .A2(n7282), .ZN(n7285) );
  XNOR2_X1 U8956 ( .A(n7285), .B(n7284), .ZN(n7290) );
  NAND2_X1 U8957 ( .A1(n8863), .A2(n7298), .ZN(n7287) );
  NOR2_X1 U8958 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9996), .ZN(n9468) );
  AOI21_X1 U8959 ( .B1(n8865), .B2(n8879), .A(n9468), .ZN(n7286) );
  OAI211_X1 U8960 ( .C1(n9087), .C2(n8868), .A(n7287), .B(n7286), .ZN(n7288)
         );
  AOI21_X1 U8961 ( .B1(n7583), .B2(n8870), .A(n7288), .ZN(n7289) );
  OAI21_X1 U8962 ( .B1(n7290), .B2(n8872), .A(n7289), .ZN(P1_U3213) );
  XOR2_X1 U8963 ( .A(n7809), .B(n7291), .Z(n9348) );
  INV_X1 U8964 ( .A(n9348), .ZN(n7304) );
  XNOR2_X1 U8965 ( .A(n7292), .B(n4810), .ZN(n7293) );
  NAND2_X1 U8966 ( .A1(n7293), .A2(n9065), .ZN(n7295) );
  AOI22_X1 U8967 ( .A1(n9254), .A2(n8879), .B1(n8877), .B2(n9251), .ZN(n7294)
         );
  NAND2_X1 U8968 ( .A1(n7295), .A2(n7294), .ZN(n9347) );
  INV_X1 U8969 ( .A(n7296), .ZN(n7297) );
  OAI211_X1 U8970 ( .C1(n7297), .C2(n9345), .A(n9530), .B(n9106), .ZN(n9344)
         );
  AOI22_X1 U8971 ( .A1(n9513), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7298), .B2(
        n9261), .ZN(n7300) );
  NAND2_X1 U8972 ( .A1(n7583), .A2(n9262), .ZN(n7299) );
  OAI211_X1 U8973 ( .C1(n9344), .C2(n7301), .A(n7300), .B(n7299), .ZN(n7302)
         );
  AOI21_X1 U8974 ( .B1(n9347), .B2(n9081), .A(n7302), .ZN(n7303) );
  OAI21_X1 U8975 ( .B1(n7304), .B2(n9114), .A(n7303), .ZN(P1_U3277) );
  NAND2_X1 U8976 ( .A1(n7305), .A2(n7907), .ZN(n7307) );
  AOI22_X1 U8977 ( .A1(n7370), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7369), .B2(
        n8360), .ZN(n7306) );
  INV_X1 U8978 ( .A(n8695), .ZN(n7329) );
  AND2_X1 U8979 ( .A1(n8265), .A2(n8140), .ZN(n7309) );
  XNOR2_X1 U8980 ( .A(n8695), .B(n8179), .ZN(n7308) );
  NOR2_X1 U8981 ( .A1(n7308), .A2(n7309), .ZN(n8109) );
  AOI21_X1 U8982 ( .B1(n7309), .B2(n7308), .A(n8109), .ZN(n7317) );
  AOI21_X1 U8983 ( .B1(n7311), .B2(n7312), .A(n7310), .ZN(n7315) );
  INV_X1 U8984 ( .A(n7311), .ZN(n7314) );
  INV_X1 U8985 ( .A(n7312), .ZN(n7313) );
  OAI21_X1 U8986 ( .B1(n7317), .B2(n4474), .A(n8110), .ZN(n7318) );
  NAND2_X1 U8987 ( .A1(n7318), .A2(n9589), .ZN(n7328) );
  INV_X1 U8988 ( .A(n8608), .ZN(n7326) );
  AND2_X1 U8989 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8340) );
  INV_X1 U8990 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U8991 ( .A1(n7319), .A2(n8358), .ZN(n7320) );
  NAND2_X1 U8992 ( .A1(n7373), .A2(n7320), .ZN(n8584) );
  OR2_X1 U8993 ( .A1(n7480), .A2(n8584), .ZN(n7324) );
  NAND2_X1 U8994 ( .A1(n7490), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U8995 ( .A1(n7489), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U8996 ( .A1(n7488), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7321) );
  NAND4_X1 U8997 ( .A1(n7324), .A2(n7323), .A3(n7322), .A4(n7321), .ZN(n8572)
         );
  INV_X1 U8998 ( .A(n8572), .ZN(n8598) );
  OAI22_X1 U8999 ( .A1(n8599), .A2(n8245), .B1(n8244), .B2(n8598), .ZN(n7325)
         );
  AOI211_X1 U9000 ( .C1(n8258), .C2(n7326), .A(n8340), .B(n7325), .ZN(n7327)
         );
  OAI211_X1 U9001 ( .C1(n7329), .C2(n9573), .A(n7328), .B(n7327), .ZN(P2_U3228) );
  NAND2_X1 U9002 ( .A1(n8102), .A2(n7330), .ZN(n7332) );
  OAI211_X1 U9003 ( .C1(n8727), .C2(n7453), .A(n7332), .B(n7331), .ZN(P2_U3330) );
  NAND2_X1 U9004 ( .A1(n7333), .A2(n7907), .ZN(n7335) );
  OR2_X1 U9005 ( .A1(n7905), .A2(n10146), .ZN(n7334) );
  INV_X1 U9006 ( .A(n8658), .ZN(n8495) );
  AND2_X1 U9007 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n7336) );
  INV_X1 U9008 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9963) );
  AND2_X1 U9009 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n7338) );
  INV_X1 U9010 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U9011 ( .A1(n7396), .A2(n8160), .ZN(n7340) );
  NAND2_X1 U9012 ( .A1(n7410), .A2(n7340), .ZN(n8492) );
  AOI22_X1 U9013 ( .A1(n7490), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n7459), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U9014 ( .A1(n7488), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7341) );
  OAI211_X1 U9015 ( .C1(n8492), .C2(n7480), .A(n7342), .B(n7341), .ZN(n8263)
         );
  INV_X1 U9016 ( .A(n8263), .ZN(n7403) );
  NAND2_X1 U9017 ( .A1(n7529), .A2(n7907), .ZN(n7344) );
  OR2_X1 U9018 ( .A1(n7905), .A2(n7846), .ZN(n7343) );
  INV_X1 U9019 ( .A(n8675), .ZN(n8546) );
  NAND2_X1 U9020 ( .A1(n7459), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U9021 ( .A1(n7353), .A2(n9963), .ZN(n7345) );
  AND2_X1 U9022 ( .A1(n7395), .A2(n7345), .ZN(n8544) );
  NAND2_X1 U9023 ( .A1(n8544), .A2(n6145), .ZN(n7348) );
  NAND2_X1 U9024 ( .A1(n7488), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U9025 ( .A1(n7490), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7346) );
  NAND4_X1 U9026 ( .A1(n7349), .A2(n7348), .A3(n7347), .A4(n7346), .ZN(n8528)
         );
  INV_X1 U9027 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7351) );
  INV_X1 U9028 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7350) );
  OAI21_X1 U9029 ( .B1(n7373), .B2(n7351), .A(n7350), .ZN(n7352) );
  NAND2_X1 U9030 ( .A1(n7353), .A2(n7352), .ZN(n8170) );
  OR2_X1 U9031 ( .A1(n7480), .A2(n8170), .ZN(n7357) );
  NAND2_X1 U9032 ( .A1(n7489), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U9033 ( .A1(n7488), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U9034 ( .A1(n7490), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7354) );
  NAND4_X1 U9035 ( .A1(n7357), .A2(n7356), .A3(n7355), .A4(n7354), .ZN(n8574)
         );
  INV_X1 U9036 ( .A(n8574), .ZN(n8243) );
  NAND2_X1 U9037 ( .A1(n7358), .A2(n7907), .ZN(n7360) );
  AOI22_X1 U9038 ( .A1(n7370), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6138), .B2(
        n7369), .ZN(n7359) );
  NAND2_X1 U9039 ( .A1(n7361), .A2(n7907), .ZN(n7363) );
  AOI22_X1 U9040 ( .A1(n7370), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7369), .B2(
        n8375), .ZN(n7362) );
  NOR2_X1 U9041 ( .A1(n7364), .A2(n8266), .ZN(n7365) );
  OR2_X1 U9042 ( .A1(n8695), .A2(n8592), .ZN(n7979) );
  NAND2_X1 U9043 ( .A1(n8695), .A2(n8592), .ZN(n8588) );
  NAND2_X1 U9044 ( .A1(n7979), .A2(n8588), .ZN(n8600) );
  AND2_X2 U9045 ( .A1(n8601), .A2(n8600), .ZN(n8603) );
  NAND2_X1 U9046 ( .A1(n8692), .A2(n8598), .ZN(n7985) );
  NAND2_X1 U9047 ( .A1(n7984), .A2(n7985), .ZN(n8589) );
  NAND2_X1 U9048 ( .A1(n7368), .A2(n7907), .ZN(n7372) );
  AOI22_X1 U9049 ( .A1(n7370), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7369), .B2(
        n8385), .ZN(n7371) );
  NAND2_X1 U9050 ( .A1(n7490), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U9051 ( .A1(n7459), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7376) );
  XNOR2_X1 U9052 ( .A(n7373), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U9053 ( .A1(n6145), .A2(n8566), .ZN(n7375) );
  NAND2_X1 U9054 ( .A1(n7488), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7374) );
  NAND4_X1 U9055 ( .A1(n7377), .A2(n7376), .A3(n7375), .A4(n7374), .ZN(n8264)
         );
  NOR2_X1 U9056 ( .A1(n8685), .A2(n8264), .ZN(n7378) );
  INV_X1 U9057 ( .A(n8685), .ZN(n8568) );
  AOI21_X1 U9058 ( .B1(n8682), .B2(n8574), .A(n8550), .ZN(n7379) );
  NAND2_X1 U9059 ( .A1(n8675), .A2(n8555), .ZN(n7999) );
  NAND2_X1 U9060 ( .A1(n8001), .A2(n7999), .ZN(n8539) );
  NAND2_X1 U9061 ( .A1(n8540), .A2(n8539), .ZN(n8673) );
  NAND2_X1 U9062 ( .A1(n7380), .A2(n7907), .ZN(n7383) );
  OR2_X1 U9063 ( .A1(n7905), .A2(n7381), .ZN(n7382) );
  INV_X1 U9064 ( .A(n8668), .ZN(n8525) );
  INV_X1 U9065 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U9066 ( .A1(n7459), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U9067 ( .A1(n7488), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7384) );
  AND2_X1 U9068 ( .A1(n7385), .A2(n7384), .ZN(n7387) );
  XNOR2_X1 U9069 ( .A(n7395), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U9070 ( .A1(n8523), .A2(n6145), .ZN(n7386) );
  OAI211_X1 U9071 ( .C1(n7389), .C2(n7388), .A(n7387), .B(n7386), .ZN(n8537)
         );
  INV_X1 U9072 ( .A(n8537), .ZN(n8227) );
  NAND2_X1 U9073 ( .A1(n8525), .A2(n8227), .ZN(n7390) );
  NAND2_X1 U9074 ( .A1(n7391), .A2(n7907), .ZN(n7394) );
  OR2_X1 U9075 ( .A1(n7905), .A2(n7392), .ZN(n7393) );
  INV_X1 U9076 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7402) );
  INV_X1 U9077 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8193) );
  INV_X1 U9078 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8237) );
  OAI21_X1 U9079 ( .B1(n7395), .B2(n8193), .A(n8237), .ZN(n7397) );
  NAND2_X1 U9080 ( .A1(n7397), .A2(n7396), .ZN(n8236) );
  OR2_X1 U9081 ( .A1(n8236), .A2(n7480), .ZN(n7401) );
  NAND2_X1 U9082 ( .A1(n7490), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U9083 ( .A1(n7489), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7398) );
  AND2_X1 U9084 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  OAI211_X1 U9085 ( .C1(n7477), .C2(n7402), .A(n7401), .B(n7400), .ZN(n8529)
         );
  INV_X1 U9086 ( .A(n8529), .ZN(n8195) );
  NAND2_X1 U9087 ( .A1(n8663), .A2(n8195), .ZN(n8004) );
  NAND2_X1 U9088 ( .A1(n8007), .A2(n8004), .ZN(n8513) );
  INV_X1 U9089 ( .A(n8663), .ZN(n8510) );
  AOI22_X2 U9090 ( .A1(n8506), .A2(n8513), .B1(n8195), .B2(n8510), .ZN(n8489)
         );
  OR2_X1 U9091 ( .A1(n8658), .A2(n7403), .ZN(n8008) );
  NAND2_X1 U9092 ( .A1(n8658), .A2(n7403), .ZN(n8013) );
  NAND2_X1 U9093 ( .A1(n8008), .A2(n8013), .ZN(n8497) );
  NAND2_X1 U9094 ( .A1(n7404), .A2(n7907), .ZN(n7407) );
  OR2_X1 U9095 ( .A1(n7905), .A2(n7405), .ZN(n7406) );
  INV_X1 U9096 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9097 ( .A1(n7410), .A2(n7409), .ZN(n7411) );
  NAND2_X1 U9098 ( .A1(n7419), .A2(n7411), .ZN(n8476) );
  OR2_X1 U9099 ( .A1(n8476), .A2(n7480), .ZN(n7414) );
  AOI22_X1 U9100 ( .A1(n7490), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n7489), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U9101 ( .A1(n7488), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U9102 ( .A1(n8653), .A2(n8161), .ZN(n8014) );
  INV_X1 U9103 ( .A(n8161), .ZN(n8501) );
  NAND2_X1 U9104 ( .A1(n7415), .A2(n7907), .ZN(n7418) );
  OR2_X1 U9105 ( .A1(n7905), .A2(n7416), .ZN(n7417) );
  INV_X1 U9106 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U9107 ( .A1(n7419), .A2(n8204), .ZN(n7420) );
  AND2_X1 U9108 ( .A1(n7431), .A2(n7420), .ZN(n8467) );
  INV_X1 U9109 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9110 ( .A1(n7490), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9111 ( .A1(n7489), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7421) );
  OAI211_X1 U9112 ( .C1(n7423), .C2(n7477), .A(n7422), .B(n7421), .ZN(n7424)
         );
  AOI21_X1 U9113 ( .B1(n8467), .B2(n6145), .A(n7424), .ZN(n8217) );
  XNOR2_X1 U9114 ( .A(n8650), .B(n8217), .ZN(n8459) );
  INV_X1 U9115 ( .A(n8217), .ZN(n8262) );
  NAND2_X1 U9116 ( .A1(n8458), .A2(n7425), .ZN(n8441) );
  NAND2_X1 U9117 ( .A1(n7426), .A2(n7907), .ZN(n7429) );
  OR2_X1 U9118 ( .A1(n7905), .A2(n7427), .ZN(n7428) );
  INV_X1 U9119 ( .A(n7431), .ZN(n7430) );
  NAND2_X1 U9120 ( .A1(n7430), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7444) );
  INV_X1 U9121 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U9122 ( .A1(n7431), .A2(n8256), .ZN(n7432) );
  NAND2_X1 U9123 ( .A1(n7444), .A2(n7432), .ZN(n8255) );
  OR2_X1 U9124 ( .A1(n8255), .A2(n7480), .ZN(n7438) );
  INV_X1 U9125 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9126 ( .A1(n7490), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9127 ( .A1(n7488), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7433) );
  OAI211_X1 U9128 ( .C1(n7448), .C2(n7435), .A(n7434), .B(n7433), .ZN(n7436)
         );
  INV_X1 U9129 ( .A(n7436), .ZN(n7437) );
  NAND2_X1 U9130 ( .A1(n7438), .A2(n7437), .ZN(n8427) );
  INV_X1 U9131 ( .A(n8427), .ZN(n8151) );
  OR2_X1 U9132 ( .A1(n8645), .A2(n8151), .ZN(n8030) );
  NAND2_X1 U9133 ( .A1(n8645), .A2(n8151), .ZN(n8024) );
  NAND2_X1 U9134 ( .A1(n8030), .A2(n8024), .ZN(n8446) );
  NAND2_X1 U9135 ( .A1(n7440), .A2(n7907), .ZN(n7443) );
  OR2_X1 U9136 ( .A1(n7905), .A2(n7441), .ZN(n7442) );
  INV_X1 U9137 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U9138 ( .A1(n7444), .A2(n8150), .ZN(n7445) );
  NAND2_X1 U9139 ( .A1(n7457), .A2(n7445), .ZN(n8434) );
  INV_X1 U9140 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U9141 ( .A1(n7488), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U9142 ( .A1(n7490), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7446) );
  OAI211_X1 U9143 ( .C1(n7448), .C2(n8435), .A(n7447), .B(n7446), .ZN(n7449)
         );
  INV_X1 U9144 ( .A(n7449), .ZN(n7450) );
  NAND2_X1 U9145 ( .A1(n8102), .A2(n7907), .ZN(n7455) );
  OR2_X1 U9146 ( .A1(n7905), .A2(n7453), .ZN(n7454) );
  INV_X1 U9147 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9148 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  NAND2_X1 U9149 ( .A1(n8413), .A2(n6145), .ZN(n7464) );
  INV_X1 U9150 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U9151 ( .A1(n7490), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9152 ( .A1(n7459), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7460) );
  OAI211_X1 U9153 ( .C1(n10001), .C2(n7477), .A(n7461), .B(n7460), .ZN(n7462)
         );
  INV_X1 U9154 ( .A(n7462), .ZN(n7463) );
  NAND2_X1 U9155 ( .A1(n8415), .A2(n8426), .ZN(n8035) );
  INV_X1 U9156 ( .A(SI_28_), .ZN(n7468) );
  NAND2_X1 U9157 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8728) );
  INV_X1 U9159 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7514) );
  MUX2_X1 U9160 ( .A(n8728), .B(n7514), .S(n5868), .Z(n7518) );
  XNOR2_X1 U9161 ( .A(n7518), .B(SI_29_), .ZN(n7472) );
  NOR2_X1 U9162 ( .A1(n7905), .A2(n8728), .ZN(n7473) );
  INV_X1 U9163 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U9164 ( .A1(n7489), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9165 ( .A1(n7490), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7474) );
  OAI211_X1 U9166 ( .C1(n7477), .C2(n7476), .A(n7475), .B(n7474), .ZN(n7478)
         );
  INV_X1 U9167 ( .A(n7478), .ZN(n7479) );
  OAI21_X1 U9168 ( .B1(n7482), .B2(n7480), .A(n7479), .ZN(n8418) );
  NOR2_X1 U9169 ( .A1(n7485), .A2(n8418), .ZN(n8040) );
  INV_X1 U9170 ( .A(n7485), .ZN(n8629) );
  NOR2_X1 U9171 ( .A1(n8582), .A2(n8685), .ZN(n8565) );
  INV_X1 U9172 ( .A(n8645), .ZN(n8455) );
  AOI21_X1 U9173 ( .B1(n8629), .B2(n8411), .A(n8403), .ZN(n8630) );
  INV_X1 U9174 ( .A(n7482), .ZN(n7483) );
  AOI22_X1 U9175 ( .A1(n7483), .A2(n9632), .B1(n9669), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n7484) );
  OAI21_X1 U9176 ( .B1(n7485), .B2(n9673), .A(n7484), .ZN(n7510) );
  INV_X1 U9177 ( .A(P2_B_REG_SCAN_IN), .ZN(n7486) );
  NOR2_X1 U9178 ( .A1(n8095), .A2(n7486), .ZN(n7487) );
  NOR2_X1 U9179 ( .A1(n9613), .A2(n7487), .ZN(n8399) );
  NAND2_X1 U9180 ( .A1(n7488), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U9181 ( .A1(n7489), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9182 ( .A1(n7490), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7491) );
  NAND3_X1 U9183 ( .A1(n7493), .A2(n7492), .A3(n7491), .ZN(n8261) );
  INV_X1 U9184 ( .A(n8261), .ZN(n7508) );
  INV_X1 U9185 ( .A(n8075), .ZN(n7973) );
  INV_X1 U9186 ( .A(n8600), .ZN(n8597) );
  INV_X1 U9187 ( .A(n8588), .ZN(n7981) );
  NOR2_X1 U9188 ( .A1(n8589), .A2(n7981), .ZN(n7495) );
  NAND2_X1 U9189 ( .A1(n8596), .A2(n7495), .ZN(n7496) );
  NAND2_X1 U9190 ( .A1(n7496), .A2(n7984), .ZN(n8570) );
  OR2_X1 U9191 ( .A1(n8685), .A2(n8593), .ZN(n7992) );
  NAND2_X1 U9192 ( .A1(n8685), .A2(n8593), .ZN(n7990) );
  NAND2_X1 U9193 ( .A1(n8570), .A2(n8569), .ZN(n7497) );
  OR2_X1 U9194 ( .A1(n8682), .A2(n8243), .ZN(n7993) );
  NAND2_X1 U9195 ( .A1(n8682), .A2(n8243), .ZN(n8534) );
  NAND2_X1 U9196 ( .A1(n7993), .A2(n8534), .ZN(n8553) );
  INV_X1 U9197 ( .A(n8534), .ZN(n7499) );
  NOR2_X1 U9198 ( .A1(n8539), .A2(n7499), .ZN(n7500) );
  OR2_X1 U9199 ( .A1(n8668), .A2(n8227), .ZN(n8000) );
  NAND2_X1 U9200 ( .A1(n8668), .A2(n8227), .ZN(n8003) );
  NAND2_X1 U9201 ( .A1(n8000), .A2(n8003), .ZN(n8526) );
  INV_X1 U9202 ( .A(n8513), .ZN(n7502) );
  INV_X1 U9203 ( .A(n8007), .ZN(n8498) );
  NOR2_X1 U9204 ( .A1(n8497), .A2(n8498), .ZN(n7503) );
  INV_X1 U9205 ( .A(n8459), .ZN(n8462) );
  OR2_X1 U9206 ( .A1(n8650), .A2(n8217), .ZN(n8019) );
  OR2_X1 U9207 ( .A1(n8638), .A2(n7912), .ZN(n8025) );
  OAI21_X1 U9208 ( .B1(n8425), .B2(n8430), .A(n8025), .ZN(n8417) );
  INV_X1 U9209 ( .A(n8416), .ZN(n8033) );
  INV_X1 U9210 ( .A(n8035), .ZN(n7506) );
  INV_X1 U9211 ( .A(n8037), .ZN(n8081) );
  NOR2_X1 U9212 ( .A1(n4413), .A2(n9669), .ZN(n7509) );
  OAI21_X1 U9213 ( .B1(n8632), .B2(n9676), .A(n7511), .ZN(P2_U3267) );
  INV_X1 U9214 ( .A(n7513), .ZN(n8729) );
  OAI222_X1 U9215 ( .A1(n4396), .A2(n8729), .B1(n7512), .B2(P1_U3084), .C1(
        n7514), .C2(n8108), .ZN(P1_U3324) );
  NAND2_X1 U9216 ( .A1(n7513), .A2(n7560), .ZN(n7516) );
  OR2_X1 U9217 ( .A1(n5185), .A2(n7514), .ZN(n7515) );
  INV_X1 U9218 ( .A(SI_29_), .ZN(n7517) );
  AND2_X1 U9219 ( .A1(n7518), .A2(n7517), .ZN(n7521) );
  INV_X1 U9220 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9221 ( .A1(n7519), .A2(SI_29_), .ZN(n7520) );
  MUX2_X1 U9222 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7555), .Z(n7551) );
  NAND2_X1 U9223 ( .A1(n7898), .A2(n7560), .ZN(n7524) );
  INV_X1 U9224 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10126) );
  OR2_X1 U9225 ( .A1(n5185), .A2(n10126), .ZN(n7523) );
  OAI21_X1 U9226 ( .B1(n8917), .B2(n7619), .A(n4419), .ZN(n9339) );
  INV_X1 U9227 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10077) );
  NOR2_X1 U9228 ( .A1(n9081), .A2(n10077), .ZN(n7526) );
  INV_X1 U9229 ( .A(n9368), .ZN(n9397) );
  AND2_X1 U9230 ( .A1(n9397), .A2(P1_B_REG_SCAN_IN), .ZN(n7525) );
  NOR2_X1 U9231 ( .A1(n9104), .A2(n7525), .ZN(n8914) );
  NAND2_X1 U9232 ( .A1(n8914), .A2(n7740), .ZN(n9338) );
  NOR2_X1 U9233 ( .A1(n9513), .A2(n9338), .ZN(n7842) );
  AOI211_X1 U9234 ( .C1(n9342), .C2(n9262), .A(n7526), .B(n7842), .ZN(n7527)
         );
  OAI21_X1 U9235 ( .B1(n9339), .B2(n7528), .A(n7527), .ZN(P1_U3262) );
  INV_X1 U9236 ( .A(n7529), .ZN(n7845) );
  OAI222_X1 U9237 ( .A1(n4396), .A2(n7845), .B1(P1_U3084), .B2(n5598), .C1(
        n9951), .C2(n8108), .ZN(P1_U3333) );
  NAND2_X1 U9238 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8891), .ZN(n7531) );
  OAI21_X1 U9239 ( .B1(n8891), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7531), .ZN(
        n8889) );
  AOI21_X1 U9240 ( .B1(n8891), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8888), .ZN(
        n9484) );
  OR2_X1 U9241 ( .A1(n9482), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9242 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9482), .ZN(n7532) );
  NAND2_X1 U9243 ( .A1(n7533), .A2(n7532), .ZN(n9485) );
  NOR2_X1 U9244 ( .A1(n9484), .A2(n9485), .ZN(n9487) );
  AOI21_X1 U9245 ( .B1(n9482), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9487), .ZN(
        n7534) );
  XNOR2_X1 U9246 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n7534), .ZN(n7541) );
  INV_X1 U9247 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7535) );
  AOI22_X1 U9248 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9482), .B1(n7536), .B2(
        n7535), .ZN(n9494) );
  AOI21_X1 U9249 ( .B1(n7538), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7537), .ZN(
        n8894) );
  XNOR2_X1 U9250 ( .A(n8891), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8893) );
  NOR2_X1 U9251 ( .A1(n8894), .A2(n8893), .ZN(n8892) );
  AOI21_X1 U9252 ( .B1(n8891), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8892), .ZN(
        n9493) );
  NAND2_X1 U9253 ( .A1(n9494), .A2(n9493), .ZN(n9492) );
  OAI21_X1 U9254 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9482), .A(n9492), .ZN(
        n7539) );
  XNOR2_X1 U9255 ( .A(n7539), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7540) );
  AOI22_X1 U9256 ( .A1(n7541), .A2(n9477), .B1(n7540), .B2(n9496), .ZN(n7543)
         );
  INV_X1 U9257 ( .A(n7540), .ZN(n7542) );
  OAI222_X1 U9258 ( .A1(n7546), .A2(n8103), .B1(n4396), .B2(n7545), .C1(
        P1_U3084), .C2(n5543), .ZN(P1_U3334) );
  NAND2_X1 U9259 ( .A1(n5496), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9260 ( .A1(n5472), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7547) );
  OAI211_X1 U9261 ( .C1(n5296), .C2(n10077), .A(n7548), .B(n7547), .ZN(n8913)
         );
  INV_X1 U9262 ( .A(n8913), .ZN(n7561) );
  INV_X1 U9263 ( .A(n7549), .ZN(n7550) );
  NAND2_X1 U9264 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  NAND2_X1 U9265 ( .A1(n7554), .A2(n7553), .ZN(n7558) );
  MUX2_X1 U9266 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7555), .Z(n7556) );
  XNOR2_X1 U9267 ( .A(n7556), .B(SI_31_), .ZN(n7557) );
  NOR2_X1 U9268 ( .A1(n5185), .A2(n5916), .ZN(n7559) );
  AND2_X1 U9269 ( .A1(n9116), .A2(n7740), .ZN(n7786) );
  INV_X1 U9270 ( .A(n8874), .ZN(n7563) );
  OR2_X1 U9271 ( .A1(n8919), .A2(n7563), .ZN(n7562) );
  AND2_X1 U9272 ( .A1(n7562), .A2(n8907), .ZN(n7565) );
  OAI211_X1 U9273 ( .C1(n4815), .C2(n7789), .A(n7731), .B(n8909), .ZN(n7564)
         );
  AOI22_X1 U9274 ( .A1(n7565), .A2(n7564), .B1(n7563), .B2(n8919), .ZN(n7782)
         );
  INV_X1 U9275 ( .A(n7782), .ZN(n7621) );
  INV_X1 U9276 ( .A(n7565), .ZN(n7785) );
  NAND2_X1 U9277 ( .A1(n7779), .A2(n7772), .ZN(n7713) );
  INV_X1 U9278 ( .A(n7713), .ZN(n7617) );
  NAND2_X1 U9279 ( .A1(n7702), .A2(n4798), .ZN(n7566) );
  NAND2_X1 U9280 ( .A1(n7566), .A2(n7703), .ZN(n7567) );
  NOR2_X1 U9281 ( .A1(n7791), .A2(n7567), .ZN(n7700) );
  INV_X1 U9282 ( .A(n7700), .ZN(n7576) );
  NAND2_X1 U9283 ( .A1(n7690), .A2(n7568), .ZN(n7686) );
  INV_X1 U9284 ( .A(n7686), .ZN(n7573) );
  INV_X1 U9285 ( .A(n7578), .ZN(n7569) );
  NOR2_X1 U9286 ( .A1(n7693), .A2(n7569), .ZN(n7697) );
  INV_X1 U9287 ( .A(n7697), .ZN(n7572) );
  INV_X1 U9288 ( .A(n7692), .ZN(n7570) );
  NAND2_X1 U9289 ( .A1(n9035), .A2(n7570), .ZN(n7696) );
  INV_X1 U9290 ( .A(n7696), .ZN(n7571) );
  OAI211_X1 U9291 ( .C1(n7573), .C2(n7572), .A(n7702), .B(n7571), .ZN(n7574)
         );
  INV_X1 U9292 ( .A(n7574), .ZN(n7575) );
  OAI211_X1 U9293 ( .C1(n7576), .C2(n7575), .A(n8965), .B(n7792), .ZN(n7777)
         );
  NAND2_X1 U9294 ( .A1(n7578), .A2(n7577), .ZN(n7685) );
  INV_X1 U9295 ( .A(n7641), .ZN(n7676) );
  AND2_X1 U9296 ( .A1(n7644), .A2(n7579), .ZN(n7638) );
  INV_X1 U9297 ( .A(n7638), .ZN(n7655) );
  NAND2_X1 U9298 ( .A1(n7667), .A2(n7580), .ZN(n7581) );
  NAND2_X1 U9299 ( .A1(n7581), .A2(n7635), .ZN(n7637) );
  INV_X1 U9300 ( .A(n7637), .ZN(n7582) );
  AND2_X1 U9301 ( .A1(n7582), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U9302 ( .A1(n7583), .A2(n9102), .ZN(n7651) );
  OAI211_X1 U9303 ( .C1(n7655), .C2(n7584), .A(n7677), .B(n7651), .ZN(n7589)
         );
  AND2_X1 U9304 ( .A1(n7651), .A2(n7585), .ZN(n7670) );
  INV_X1 U9305 ( .A(n7670), .ZN(n7646) );
  NAND2_X1 U9306 ( .A1(n7635), .A2(n7586), .ZN(n7642) );
  NOR2_X1 U9307 ( .A1(n7646), .A2(n7642), .ZN(n7608) );
  NAND2_X1 U9308 ( .A1(n7634), .A2(n7630), .ZN(n7587) );
  NAND2_X1 U9309 ( .A1(n7587), .A2(n7632), .ZN(n7664) );
  NAND3_X1 U9310 ( .A1(n4787), .A2(n7632), .A3(n7627), .ZN(n7665) );
  NAND4_X1 U9311 ( .A1(n7608), .A2(n7677), .A3(n7664), .A4(n7665), .ZN(n7588)
         );
  AND4_X1 U9312 ( .A1(n7682), .A2(n7676), .A3(n7589), .A4(n7588), .ZN(n7590)
         );
  OR3_X1 U9313 ( .A1(n7685), .A2(n7610), .A3(n7590), .ZN(n7771) );
  AND2_X1 U9314 ( .A1(n7657), .A2(n7591), .ZN(n7592) );
  AND2_X1 U9315 ( .A1(n7601), .A2(n7592), .ZN(n7799) );
  INV_X1 U9316 ( .A(n7799), .ZN(n7594) );
  INV_X1 U9317 ( .A(n7661), .ZN(n7593) );
  NOR2_X1 U9318 ( .A1(n7594), .A2(n7593), .ZN(n7766) );
  AOI211_X1 U9319 ( .C1(n9507), .C2(n5613), .A(n7825), .B(n7595), .ZN(n7598)
         );
  OAI22_X1 U9320 ( .A1(n7598), .A2(n7597), .B1(n7596), .B2(n7869), .ZN(n7600)
         );
  NAND3_X1 U9321 ( .A1(n7600), .A2(n7757), .A3(n7599), .ZN(n7605) );
  INV_X1 U9322 ( .A(n7601), .ZN(n7603) );
  OAI21_X1 U9323 ( .B1(n7603), .B2(n7758), .A(n7602), .ZN(n7604) );
  AOI22_X1 U9324 ( .A1(n7766), .A2(n7605), .B1(n7604), .B2(n7661), .ZN(n7606)
         );
  INV_X1 U9325 ( .A(n7606), .ZN(n7613) );
  NAND2_X1 U9326 ( .A1(n7629), .A2(n7625), .ZN(n7662) );
  INV_X1 U9327 ( .A(n7662), .ZN(n7607) );
  NAND4_X1 U9328 ( .A1(n7608), .A2(n7607), .A3(n7677), .A4(n7664), .ZN(n7609)
         );
  OR3_X1 U9329 ( .A1(n7685), .A2(n7610), .A3(n7609), .ZN(n7611) );
  AOI21_X1 U9330 ( .B1(n7771), .B2(n7611), .A(n7693), .ZN(n7612) );
  NAND2_X1 U9331 ( .A1(n7700), .A2(n7612), .ZN(n7774) );
  AOI21_X1 U9332 ( .B1(n7771), .B2(n7613), .A(n7774), .ZN(n7615) );
  AND2_X1 U9333 ( .A1(n9156), .A2(n10145), .ZN(n7708) );
  INV_X1 U9334 ( .A(n7708), .ZN(n7614) );
  OAI211_X1 U9335 ( .C1(n7777), .C2(n7615), .A(n7614), .B(n7709), .ZN(n7616)
         );
  AOI21_X1 U9336 ( .B1(n7617), .B2(n7616), .A(n7724), .ZN(n7618) );
  NOR4_X1 U9337 ( .A1(n7785), .A2(n7790), .A3(n7618), .A4(n8926), .ZN(n7620)
         );
  AND2_X1 U9338 ( .A1(n7619), .A2(n8913), .ZN(n7818) );
  INV_X1 U9339 ( .A(n7818), .ZN(n7741) );
  OAI21_X1 U9340 ( .B1(n7621), .B2(n7620), .A(n7741), .ZN(n7624) );
  INV_X1 U9341 ( .A(n9116), .ZN(n7742) );
  INV_X1 U9342 ( .A(n7740), .ZN(n7622) );
  INV_X1 U9343 ( .A(n7819), .ZN(n7623) );
  AOI21_X1 U9344 ( .B1(n7821), .B2(n7624), .A(n7623), .ZN(n7833) );
  NAND3_X1 U9345 ( .A1(n7626), .A2(n7762), .A3(n7625), .ZN(n7628) );
  NAND3_X1 U9346 ( .A1(n7628), .A2(n7627), .A3(n7661), .ZN(n7631) );
  NAND3_X1 U9347 ( .A1(n7631), .A2(n7630), .A3(n7629), .ZN(n7633) );
  NAND3_X1 U9348 ( .A1(n7633), .A2(n7632), .A3(n4787), .ZN(n7636) );
  NAND3_X1 U9349 ( .A1(n7636), .A2(n7635), .A3(n7634), .ZN(n7639) );
  AND2_X1 U9350 ( .A1(n7637), .A2(n7746), .ZN(n7649) );
  NAND3_X1 U9351 ( .A1(n7639), .A2(n7638), .A3(n7649), .ZN(n7675) );
  INV_X1 U9352 ( .A(n7677), .ZN(n7640) );
  NAND2_X1 U9353 ( .A1(n7642), .A2(n7667), .ZN(n7669) );
  INV_X1 U9354 ( .A(n7746), .ZN(n7750) );
  NAND3_X1 U9355 ( .A1(n7669), .A2(n7750), .A3(n7643), .ZN(n7647) );
  NAND3_X1 U9356 ( .A1(n7646), .A2(n7644), .A3(n7746), .ZN(n7645) );
  OAI21_X1 U9357 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7648) );
  NOR2_X1 U9358 ( .A1(n9100), .A2(n7648), .ZN(n7674) );
  INV_X1 U9359 ( .A(n7649), .ZN(n7650) );
  NOR2_X1 U9360 ( .A1(n7650), .A2(n7805), .ZN(n7654) );
  NAND2_X1 U9361 ( .A1(n7651), .A2(n7750), .ZN(n7652) );
  NAND2_X1 U9362 ( .A1(n7655), .A2(n7652), .ZN(n7653) );
  OAI21_X1 U9363 ( .B1(n7655), .B2(n7654), .A(n7653), .ZN(n7673) );
  AND2_X1 U9364 ( .A1(n7657), .A2(n7656), .ZN(n7759) );
  OAI21_X1 U9365 ( .B1(n6726), .B2(n4506), .A(n7759), .ZN(n7659) );
  NAND3_X1 U9366 ( .A1(n7659), .A2(n7658), .A3(n7761), .ZN(n7663) );
  AND2_X1 U9367 ( .A1(n7661), .A2(n7660), .ZN(n7765) );
  AOI21_X1 U9368 ( .B1(n7663), .B2(n7765), .A(n7662), .ZN(n7666) );
  OAI21_X1 U9369 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7668) );
  NAND2_X1 U9370 ( .A1(n7668), .A2(n7667), .ZN(n7671) );
  NAND4_X1 U9371 ( .A1(n7671), .A2(n7750), .A3(n7670), .A4(n7669), .ZN(n7672)
         );
  NAND4_X1 U9372 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n7680)
         );
  MUX2_X1 U9373 ( .A(n7677), .B(n7676), .S(n7746), .Z(n7678) );
  NAND3_X1 U9374 ( .A1(n7680), .A2(n7679), .A3(n7678), .ZN(n7684) );
  MUX2_X1 U9375 ( .A(n7682), .B(n7681), .S(n7746), .Z(n7683) );
  NAND3_X1 U9376 ( .A1(n7684), .A2(n9071), .A3(n7683), .ZN(n7689) );
  MUX2_X1 U9377 ( .A(n7686), .B(n7685), .S(n7750), .Z(n7687) );
  INV_X1 U9378 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U9379 ( .A1(n7689), .A2(n7688), .ZN(n7698) );
  INV_X1 U9380 ( .A(n7690), .ZN(n7691) );
  NOR2_X1 U9381 ( .A1(n7692), .A2(n7691), .ZN(n7695) );
  NAND2_X1 U9382 ( .A1(n7794), .A2(n4801), .ZN(n7694) );
  NAND2_X1 U9383 ( .A1(n7705), .A2(n7702), .ZN(n7701) );
  INV_X1 U9384 ( .A(n7792), .ZN(n7699) );
  AOI21_X1 U9385 ( .B1(n7701), .B2(n7700), .A(n7699), .ZN(n7707) );
  NAND2_X1 U9386 ( .A1(n7702), .A2(n9035), .ZN(n7704) );
  MUX2_X1 U9387 ( .A(n7707), .B(n7706), .S(n7750), .Z(n7716) );
  NAND2_X1 U9388 ( .A1(n8967), .A2(n8980), .ZN(n7715) );
  NAND2_X1 U9389 ( .A1(n7772), .A2(n7708), .ZN(n7710) );
  AND2_X1 U9390 ( .A1(n7710), .A2(n7709), .ZN(n7711) );
  AND2_X1 U9391 ( .A1(n7711), .A2(n7717), .ZN(n7775) );
  INV_X1 U9392 ( .A(n8965), .ZN(n7712) );
  AND2_X1 U9393 ( .A1(n8967), .A2(n7712), .ZN(n7714) );
  NAND2_X1 U9394 ( .A1(n7718), .A2(n8786), .ZN(n7721) );
  AOI21_X1 U9395 ( .B1(n8944), .B2(n4821), .A(n8959), .ZN(n7719) );
  MUX2_X1 U9396 ( .A(n8944), .B(n7719), .S(n7750), .Z(n7720) );
  NAND2_X1 U9397 ( .A1(n7721), .A2(n7720), .ZN(n7730) );
  INV_X1 U9398 ( .A(n7722), .ZN(n7723) );
  NAND2_X1 U9399 ( .A1(n7723), .A2(n8932), .ZN(n7728) );
  OAI21_X1 U9400 ( .B1(n8944), .B2(n4821), .A(n7731), .ZN(n7726) );
  OAI21_X1 U9401 ( .B1(n8786), .B2(n7724), .A(n7781), .ZN(n7725) );
  MUX2_X1 U9402 ( .A(n7726), .B(n7725), .S(n7746), .Z(n7727) );
  NAND2_X1 U9403 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  NAND2_X1 U9404 ( .A1(n7730), .A2(n7729), .ZN(n7734) );
  MUX2_X1 U9405 ( .A(n7731), .B(n7781), .S(n7750), .Z(n7732) );
  AND2_X1 U9406 ( .A1(n7816), .A2(n7732), .ZN(n7733) );
  MUX2_X1 U9407 ( .A(n8909), .B(n8907), .S(n7746), .Z(n7735) );
  NAND2_X1 U9408 ( .A1(n8919), .A2(n7746), .ZN(n7738) );
  NAND2_X1 U9409 ( .A1(n7740), .A2(n8913), .ZN(n7736) );
  NAND2_X1 U9410 ( .A1(n9342), .A2(n7736), .ZN(n7783) );
  INV_X1 U9411 ( .A(n8919), .ZN(n9122) );
  NAND4_X1 U9412 ( .A1(n7783), .A2(n9122), .A3(n7750), .A4(n8874), .ZN(n7737)
         );
  OAI21_X1 U9413 ( .B1(n7749), .B2(n7738), .A(n7737), .ZN(n7745) );
  AOI21_X1 U9414 ( .B1(n8919), .B2(n7750), .A(n8874), .ZN(n7739) );
  NAND2_X1 U9415 ( .A1(n7741), .A2(n7740), .ZN(n7743) );
  NAND2_X1 U9416 ( .A1(n7743), .A2(n7742), .ZN(n7788) );
  OAI21_X1 U9417 ( .B1(n7745), .B2(n7744), .A(n7788), .ZN(n7754) );
  INV_X1 U9418 ( .A(n7783), .ZN(n7747) );
  NAND3_X1 U9419 ( .A1(n7819), .A2(n7747), .A3(n7746), .ZN(n7748) );
  INV_X1 U9420 ( .A(n7786), .ZN(n7756) );
  AND2_X1 U9421 ( .A1(n7748), .A2(n7756), .ZN(n7753) );
  NAND2_X1 U9422 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  AND3_X1 U9423 ( .A1(n7754), .A2(n7753), .A3(n7752), .ZN(n7830) );
  NAND3_X1 U9424 ( .A1(n7756), .A2(n5599), .A3(n7755), .ZN(n7829) );
  INV_X1 U9425 ( .A(n7790), .ZN(n7780) );
  NAND2_X1 U9426 ( .A1(n7758), .A2(n7757), .ZN(n7760) );
  NAND2_X1 U9427 ( .A1(n7760), .A2(n7759), .ZN(n7764) );
  AND2_X1 U9428 ( .A1(n7762), .A2(n7761), .ZN(n7763) );
  NAND2_X1 U9429 ( .A1(n7764), .A2(n7763), .ZN(n7797) );
  INV_X1 U9430 ( .A(n7797), .ZN(n7769) );
  INV_X1 U9431 ( .A(n7765), .ZN(n7768) );
  NAND2_X1 U9432 ( .A1(n6536), .A2(n7766), .ZN(n7767) );
  OAI21_X1 U9433 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n7770) );
  AND2_X1 U9434 ( .A1(n7771), .A2(n7770), .ZN(n7773) );
  OAI21_X1 U9435 ( .B1(n7774), .B2(n7773), .A(n7772), .ZN(n7776) );
  OAI21_X1 U9436 ( .B1(n7777), .B2(n7776), .A(n7775), .ZN(n7778) );
  NAND4_X1 U9437 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n7784)
         );
  OAI211_X1 U9438 ( .C1(n7785), .C2(n7784), .A(n7783), .B(n7782), .ZN(n7787)
         );
  AOI21_X1 U9439 ( .B1(n7788), .B2(n7787), .A(n7786), .ZN(n7822) );
  XNOR2_X1 U9440 ( .A(n8919), .B(n8874), .ZN(n8905) );
  INV_X1 U9441 ( .A(n8905), .ZN(n8911) );
  INV_X1 U9442 ( .A(n8957), .ZN(n7814) );
  INV_X1 U9443 ( .A(n7791), .ZN(n7793) );
  NAND2_X1 U9444 ( .A1(n7793), .A2(n7792), .ZN(n8999) );
  NAND2_X1 U9445 ( .A1(n9035), .A2(n7794), .ZN(n9031) );
  NOR3_X1 U9446 ( .A1(n7797), .A2(n5566), .A3(n7796), .ZN(n7800) );
  INV_X1 U9447 ( .A(n7801), .ZN(n7802) );
  NOR4_X1 U9448 ( .A1(n7804), .A2(n9249), .A3(n7803), .A4(n7802), .ZN(n7808)
         );
  NAND4_X1 U9449 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n7810)
         );
  NOR4_X1 U9450 ( .A1(n9084), .A2(n7810), .A3(n9100), .A4(n7809), .ZN(n7811)
         );
  NAND4_X1 U9451 ( .A1(n9044), .A2(n9071), .A3(n9061), .A4(n7811), .ZN(n7812)
         );
  NOR4_X1 U9452 ( .A1(n8999), .A2(n9006), .A3(n9031), .A4(n7812), .ZN(n7813)
         );
  AND4_X1 U9453 ( .A1(n7814), .A2(n8967), .A3(n7813), .A4(n8980), .ZN(n7815)
         );
  NAND4_X1 U9454 ( .A1(n7816), .A2(n8932), .A3(n8946), .A4(n7815), .ZN(n7817)
         );
  NOR3_X1 U9455 ( .A1(n7818), .A2(n8911), .A3(n7817), .ZN(n7820) );
  NAND3_X1 U9456 ( .A1(n7821), .A2(n7820), .A3(n7819), .ZN(n7826) );
  MUX2_X1 U9457 ( .A(n7822), .B(n7826), .S(n7825), .Z(n7823) );
  NAND4_X1 U9458 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n9397), .ZN(n7837)
         );
  OAI211_X1 U9459 ( .C1(n7838), .C2(n7840), .A(n7837), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7839) );
  OAI21_X1 U9460 ( .B1(n7841), .B2(n7840), .A(n7839), .ZN(P1_U3240) );
  XNOR2_X1 U9461 ( .A(n4419), .B(n9116), .ZN(n9115) );
  NAND2_X1 U9462 ( .A1(n9115), .A2(n9068), .ZN(n7844) );
  AOI21_X1 U9463 ( .B1(n9513), .B2(P1_REG2_REG_31__SCAN_IN), .A(n7842), .ZN(
        n7843) );
  OAI211_X1 U9464 ( .C1(n9116), .C2(n9110), .A(n7844), .B(n7843), .ZN(P1_U3261) );
  OAI222_X1 U9465 ( .A1(n8727), .A2(n7846), .B1(n7895), .B2(n7845), .C1(n6087), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U9466 ( .A1(n7848), .A2(n7847), .ZN(n7852) );
  NAND2_X1 U9467 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  XOR2_X1 U9468 ( .A(n7852), .B(n7851), .Z(n7861) );
  NOR2_X1 U9469 ( .A1(n7853), .A2(n8852), .ZN(n7854) );
  AOI211_X1 U9470 ( .C1(n8839), .C2(n8882), .A(n7855), .B(n7854), .ZN(n7856)
         );
  OAI21_X1 U9471 ( .B1(n7857), .B2(n8859), .A(n7856), .ZN(n7858) );
  AOI21_X1 U9472 ( .B1(n7859), .B2(n8863), .A(n7858), .ZN(n7860) );
  OAI21_X1 U9473 ( .B1(n7861), .B2(n8872), .A(n7860), .ZN(P1_U3211) );
  OAI21_X1 U9474 ( .B1(n7862), .B2(n7864), .A(n7863), .ZN(n7865) );
  NAND2_X1 U9475 ( .A1(n7865), .A2(n8849), .ZN(n7871) );
  OAI22_X1 U9476 ( .A1(n8868), .A2(n7867), .B1(n7866), .B2(n8852), .ZN(n7868)
         );
  AOI21_X1 U9477 ( .B1(n7869), .B2(n8870), .A(n7868), .ZN(n7870) );
  OAI211_X1 U9478 ( .C1(n7873), .C2(n7872), .A(n7871), .B(n7870), .ZN(P1_U3235) );
  XOR2_X1 U9479 ( .A(n8064), .B(n7874), .Z(n9729) );
  XNOR2_X1 U9480 ( .A(n7875), .B(n8064), .ZN(n7877) );
  AOI22_X1 U9481 ( .A1(n8571), .A2(n8276), .B1(n8274), .B2(n8573), .ZN(n9587)
         );
  INV_X1 U9482 ( .A(n9587), .ZN(n7876) );
  AOI21_X1 U9483 ( .B1(n7877), .B2(n9662), .A(n7876), .ZN(n9732) );
  MUX2_X1 U9484 ( .A(n6251), .B(n9732), .S(n9618), .Z(n7881) );
  AND2_X1 U9485 ( .A1(n9615), .A2(n9583), .ZN(n7878) );
  OR2_X1 U9486 ( .A1(n7878), .A2(n7887), .ZN(n9731) );
  OAI22_X1 U9487 ( .A1(n9636), .A2(n9731), .B1(n9592), .B2(n9666), .ZN(n7879)
         );
  AOI21_X1 U9488 ( .B1(n9631), .B2(n9583), .A(n7879), .ZN(n7880) );
  OAI211_X1 U9489 ( .C1(n9729), .C2(n9676), .A(n7881), .B(n7880), .ZN(P2_U3290) );
  XNOR2_X1 U9490 ( .A(n7882), .B(n6846), .ZN(n9741) );
  AOI21_X1 U9491 ( .B1(n7883), .B2(n8061), .A(n9644), .ZN(n7886) );
  OAI22_X1 U9492 ( .A1(n9612), .A2(n9611), .B1(n7942), .B2(n9613), .ZN(n7884)
         );
  AOI21_X1 U9493 ( .B1(n7886), .B2(n7885), .A(n7884), .ZN(n9739) );
  MUX2_X1 U9494 ( .A(n6278), .B(n9739), .S(n9618), .Z(n7894) );
  INV_X1 U9495 ( .A(n7887), .ZN(n7889) );
  AOI21_X1 U9496 ( .B1(n9736), .B2(n7889), .A(n7888), .ZN(n9737) );
  OAI22_X1 U9497 ( .A1(n9673), .A2(n7891), .B1(n9666), .B2(n7890), .ZN(n7892)
         );
  AOI21_X1 U9498 ( .B1(n9737), .B2(n9668), .A(n7892), .ZN(n7893) );
  OAI211_X1 U9499 ( .C1(n9741), .C2(n9676), .A(n7894), .B(n7893), .ZN(P2_U3289) );
  INV_X1 U9500 ( .A(n7898), .ZN(n8107) );
  INV_X1 U9501 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7899) );
  OAI222_X1 U9502 ( .A1(P2_U3152), .A2(n7896), .B1(n7895), .B2(n8107), .C1(
        n7899), .C2(n8727), .ZN(P2_U3328) );
  NAND2_X1 U9503 ( .A1(n7898), .A2(n7907), .ZN(n7901) );
  OR2_X1 U9504 ( .A1(n7905), .A2(n7899), .ZN(n7900) );
  OAI22_X1 U9505 ( .A1(n7902), .A2(n8043), .B1(n6548), .B2(n8398), .ZN(n7903)
         );
  OAI21_X1 U9506 ( .B1(n7904), .B2(n8625), .A(n7903), .ZN(n7910) );
  NOR2_X1 U9507 ( .A1(n7905), .A2(n5963), .ZN(n7906) );
  INV_X1 U9508 ( .A(n8619), .ZN(n7909) );
  INV_X1 U9509 ( .A(n8398), .ZN(n7908) );
  NAND2_X1 U9510 ( .A1(n8625), .A2(n7508), .ZN(n8038) );
  NOR2_X1 U9511 ( .A1(n8619), .A2(n8398), .ZN(n8042) );
  NAND2_X1 U9512 ( .A1(n8638), .A2(n7912), .ZN(n8028) );
  INV_X1 U9513 ( .A(n8046), .ZN(n8029) );
  OR2_X1 U9514 ( .A1(n7913), .A2(n6548), .ZN(n7914) );
  INV_X1 U9515 ( .A(n7921), .ZN(n7915) );
  INV_X1 U9516 ( .A(n7918), .ZN(n7917) );
  AOI211_X1 U9517 ( .C1(n7925), .C2(n8059), .A(n7917), .B(n7916), .ZN(n7920)
         );
  NAND2_X1 U9518 ( .A1(n8055), .A2(n7918), .ZN(n7919) );
  OAI211_X1 U9519 ( .C1(n7920), .C2(n7930), .A(n7936), .B(n8055), .ZN(n7927)
         );
  NAND2_X1 U9520 ( .A1(n8059), .A2(n7921), .ZN(n7922) );
  AOI211_X1 U9521 ( .C1(n7924), .C2(n7923), .A(n7922), .B(n7930), .ZN(n7926)
         );
  AOI22_X1 U9522 ( .A1(n7927), .A2(n8029), .B1(n7926), .B2(n7925), .ZN(n7934)
         );
  AND2_X1 U9523 ( .A1(n8275), .A2(n9730), .ZN(n7933) );
  AOI22_X1 U9524 ( .A1(n7930), .A2(n8054), .B1(n7929), .B2(n7928), .ZN(n7931)
         );
  OAI21_X1 U9525 ( .B1(n7931), .B2(n7933), .A(n8046), .ZN(n7932) );
  OAI21_X1 U9526 ( .B1(n7934), .B2(n7933), .A(n7932), .ZN(n7935) );
  OAI211_X1 U9527 ( .C1(n7936), .C2(n8029), .A(n7935), .B(n6846), .ZN(n7940)
         );
  MUX2_X1 U9528 ( .A(n7938), .B(n7937), .S(n8046), .Z(n7939) );
  OAI21_X1 U9529 ( .B1(n7942), .B2(n7941), .A(n7948), .ZN(n7943) );
  INV_X1 U9530 ( .A(n7943), .ZN(n7945) );
  AND2_X1 U9531 ( .A1(n7952), .A2(n7947), .ZN(n7949) );
  MUX2_X1 U9532 ( .A(n7949), .B(n7948), .S(n8046), .Z(n7950) );
  AND2_X1 U9533 ( .A1(n7953), .A2(n7952), .ZN(n7954) );
  MUX2_X1 U9534 ( .A(n7955), .B(n7954), .S(n8046), .Z(n7956) );
  AOI211_X1 U9535 ( .C1(n7962), .C2(n7958), .A(n7966), .B(n7079), .ZN(n7960)
         );
  OR2_X1 U9536 ( .A1(n7960), .A2(n7959), .ZN(n7969) );
  NAND2_X1 U9537 ( .A1(n7962), .A2(n7961), .ZN(n7964) );
  AOI21_X1 U9538 ( .B1(n7964), .B2(n7963), .A(n7079), .ZN(n7967) );
  OAI22_X1 U9539 ( .A1(n7967), .A2(n7966), .B1(n7965), .B2(n9325), .ZN(n7968)
         );
  MUX2_X1 U9540 ( .A(n7969), .B(n7968), .S(n8046), .Z(n7974) );
  MUX2_X1 U9541 ( .A(n7971), .B(n7970), .S(n8046), .Z(n7972) );
  OAI211_X1 U9542 ( .C1(n7974), .C2(n8053), .A(n7973), .B(n7972), .ZN(n7978)
         );
  MUX2_X1 U9543 ( .A(n7976), .B(n7975), .S(n8046), .Z(n7977) );
  INV_X1 U9544 ( .A(n7979), .ZN(n7980) );
  MUX2_X1 U9545 ( .A(n7981), .B(n7980), .S(n8046), .Z(n7982) );
  NOR3_X1 U9546 ( .A1(n7983), .A2(n7982), .A3(n8589), .ZN(n7989) );
  INV_X1 U9547 ( .A(n7984), .ZN(n7987) );
  NAND2_X1 U9548 ( .A1(n7990), .A2(n7985), .ZN(n7986) );
  MUX2_X1 U9549 ( .A(n7987), .B(n7986), .S(n8046), .Z(n7988) );
  INV_X1 U9550 ( .A(n7990), .ZN(n7991) );
  NAND2_X1 U9551 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  OAI21_X1 U9552 ( .B1(n7995), .B2(n7994), .A(n8534), .ZN(n7996) );
  NAND2_X1 U9553 ( .A1(n7996), .A2(n8001), .ZN(n7997) );
  MUX2_X1 U9554 ( .A(n7998), .B(n7997), .S(n8046), .Z(n8002) );
  NAND3_X1 U9555 ( .A1(n8002), .A2(n8001), .A3(n8000), .ZN(n8005) );
  NAND3_X1 U9556 ( .A1(n8005), .A2(n8004), .A3(n8003), .ZN(n8006) );
  NAND3_X1 U9557 ( .A1(n8010), .A2(n8007), .A3(n8006), .ZN(n8012) );
  NAND2_X1 U9558 ( .A1(n8480), .A2(n8008), .ZN(n8009) );
  OAI21_X1 U9559 ( .B1(n8010), .B2(n8009), .A(n8014), .ZN(n8011) );
  AOI21_X1 U9560 ( .B1(n8029), .B2(n8012), .A(n8011), .ZN(n8016) );
  AOI21_X1 U9561 ( .B1(n8014), .B2(n8013), .A(n8046), .ZN(n8015) );
  NOR2_X1 U9562 ( .A1(n8016), .A2(n8015), .ZN(n8023) );
  OAI21_X1 U9563 ( .B1(n8046), .B2(n8017), .A(n8462), .ZN(n8022) );
  INV_X1 U9564 ( .A(n8024), .ZN(n8018) );
  AOI21_X1 U9565 ( .B1(n8217), .B2(n8650), .A(n8018), .ZN(n8020) );
  MUX2_X1 U9566 ( .A(n8020), .B(n8019), .S(n8046), .Z(n8021) );
  INV_X1 U9567 ( .A(n8430), .ZN(n8424) );
  NAND3_X1 U9568 ( .A1(n8031), .A2(n8424), .A3(n8024), .ZN(n8026) );
  AND2_X1 U9569 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  NAND4_X1 U9570 ( .A1(n8031), .A2(n8424), .A3(n8030), .A4(n8029), .ZN(n8032)
         );
  MUX2_X1 U9571 ( .A(n8035), .B(n8034), .S(n8046), .Z(n8036) );
  MUX2_X1 U9572 ( .A(n8040), .B(n8039), .S(n8046), .Z(n8041) );
  INV_X1 U9573 ( .A(n8042), .ZN(n8047) );
  INV_X1 U9574 ( .A(n8043), .ZN(n8044) );
  NAND2_X1 U9575 ( .A1(n8047), .A2(n8044), .ZN(n8052) );
  INV_X1 U9576 ( .A(n8083), .ZN(n8045) );
  MUX2_X1 U9577 ( .A(n8052), .B(n8045), .S(n8046), .Z(n8050) );
  MUX2_X1 U9578 ( .A(n8048), .B(n8047), .S(n8046), .Z(n8049) );
  INV_X1 U9579 ( .A(n8052), .ZN(n8084) );
  INV_X1 U9580 ( .A(n8539), .ZN(n8535) );
  INV_X1 U9581 ( .A(n8553), .ZN(n8077) );
  INV_X1 U9582 ( .A(n8053), .ZN(n8073) );
  NOR2_X1 U9583 ( .A1(n9629), .A2(n9675), .ZN(n8058) );
  AND2_X1 U9584 ( .A1(n8055), .A2(n8054), .ZN(n9607) );
  AND2_X1 U9585 ( .A1(n8056), .A2(n8089), .ZN(n8057) );
  NAND4_X1 U9586 ( .A1(n8059), .A2(n8058), .A3(n9607), .A4(n8057), .ZN(n8062)
         );
  NOR3_X1 U9587 ( .A1(n8062), .A2(n8061), .A3(n8060), .ZN(n8066) );
  NAND4_X1 U9588 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), .ZN(n8069)
         );
  NOR3_X1 U9589 ( .A1(n8069), .A2(n8068), .A3(n8067), .ZN(n8071) );
  NAND4_X1 U9590 ( .A1(n8073), .A2(n8072), .A3(n8071), .A4(n8070), .ZN(n8074)
         );
  NOR4_X1 U9591 ( .A1(n8589), .A2(n8600), .A3(n8075), .A4(n8074), .ZN(n8076)
         );
  NAND4_X1 U9592 ( .A1(n8535), .A2(n8077), .A3(n8569), .A4(n8076), .ZN(n8078)
         );
  NOR4_X1 U9593 ( .A1(n8497), .A2(n8513), .A3(n8526), .A4(n8078), .ZN(n8079)
         );
  NAND4_X1 U9594 ( .A1(n7505), .A2(n8480), .A3(n8079), .A4(n8462), .ZN(n8080)
         );
  NOR4_X1 U9595 ( .A1(n8081), .A2(n8430), .A3(n8416), .A4(n8080), .ZN(n8082)
         );
  NAND3_X1 U9596 ( .A1(n8084), .A2(n8083), .A3(n8082), .ZN(n8085) );
  XNOR2_X1 U9597 ( .A(n8085), .B(n6138), .ZN(n8087) );
  NOR2_X1 U9598 ( .A1(n8086), .A2(n8089), .ZN(n8091) );
  AOI21_X1 U9599 ( .B1(n8087), .B2(n6548), .A(n8091), .ZN(n8088) );
  OAI21_X1 U9600 ( .B1(n9752), .B2(n8091), .A(n8090), .ZN(n8092) );
  INV_X1 U9601 ( .A(n9681), .ZN(n8096) );
  NOR4_X1 U9602 ( .A1(n8096), .A2(n8095), .A3(n8094), .A4(n9611), .ZN(n8099)
         );
  OAI21_X1 U9603 ( .B1(n8100), .B2(n8097), .A(P2_B_REG_SCAN_IN), .ZN(n8098) );
  OAI22_X1 U9604 ( .A1(n8101), .A2(n8100), .B1(n8099), .B2(n8098), .ZN(
        P2_U3244) );
  INV_X1 U9605 ( .A(n8102), .ZN(n8105) );
  OAI222_X1 U9606 ( .A1(n4396), .A2(n8105), .B1(n5524), .B2(P1_U3084), .C1(
        n8104), .C2(n8103), .ZN(P1_U3325) );
  OAI222_X1 U9607 ( .A1(n8108), .A2(n10126), .B1(n4396), .B2(n8107), .C1(
        P1_U3084), .C2(n8106), .ZN(P1_U3323) );
  XNOR2_X1 U9608 ( .A(n8692), .B(n8145), .ZN(n8112) );
  NAND2_X1 U9609 ( .A1(n8572), .A2(n8140), .ZN(n8111) );
  XNOR2_X1 U9610 ( .A(n8112), .B(n8111), .ZN(n8209) );
  XNOR2_X1 U9611 ( .A(n8685), .B(n8179), .ZN(n8115) );
  NAND2_X1 U9612 ( .A1(n8264), .A2(n8140), .ZN(n8113) );
  XNOR2_X1 U9613 ( .A(n8115), .B(n8113), .ZN(n8241) );
  INV_X1 U9614 ( .A(n8113), .ZN(n8114) );
  AOI21_X2 U9615 ( .B1(n8242), .B2(n8241), .A(n8116), .ZN(n8168) );
  AND2_X1 U9616 ( .A1(n8574), .A2(n8140), .ZN(n8118) );
  XNOR2_X1 U9617 ( .A(n8682), .B(n8179), .ZN(n8117) );
  NOR2_X1 U9618 ( .A1(n8117), .A2(n8118), .ZN(n8119) );
  AOI21_X1 U9619 ( .B1(n8118), .B2(n8117), .A(n8119), .ZN(n8167) );
  INV_X1 U9620 ( .A(n8119), .ZN(n8120) );
  XNOR2_X1 U9621 ( .A(n8675), .B(n8145), .ZN(n8122) );
  NAND2_X1 U9622 ( .A1(n8528), .A2(n8140), .ZN(n8121) );
  XNOR2_X1 U9623 ( .A(n8122), .B(n8121), .ZN(n8224) );
  XNOR2_X1 U9624 ( .A(n8668), .B(n8179), .ZN(n8124) );
  NAND2_X1 U9625 ( .A1(n8537), .A2(n8140), .ZN(n8123) );
  XNOR2_X1 U9626 ( .A(n8124), .B(n8123), .ZN(n8191) );
  INV_X1 U9627 ( .A(n8123), .ZN(n8125) );
  XNOR2_X1 U9628 ( .A(n8663), .B(n8179), .ZN(n8126) );
  XNOR2_X1 U9629 ( .A(n8128), .B(n8126), .ZN(n8234) );
  NAND2_X1 U9630 ( .A1(n8529), .A2(n8140), .ZN(n8233) );
  NAND2_X1 U9631 ( .A1(n8234), .A2(n8233), .ZN(n8232) );
  INV_X1 U9632 ( .A(n8126), .ZN(n8127) );
  NAND2_X1 U9633 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  NAND2_X1 U9634 ( .A1(n8232), .A2(n8129), .ZN(n8159) );
  XNOR2_X1 U9635 ( .A(n8658), .B(n8179), .ZN(n8157) );
  AND2_X1 U9636 ( .A1(n8263), .A2(n8140), .ZN(n8156) );
  NOR2_X1 U9637 ( .A1(n8157), .A2(n8156), .ZN(n8131) );
  NAND2_X1 U9638 ( .A1(n8157), .A2(n8156), .ZN(n8130) );
  XNOR2_X1 U9639 ( .A(n8653), .B(n8145), .ZN(n8132) );
  XNOR2_X1 U9640 ( .A(n8134), .B(n8132), .ZN(n8216) );
  NOR2_X1 U9641 ( .A1(n8161), .A2(n6193), .ZN(n8215) );
  NAND2_X1 U9642 ( .A1(n8216), .A2(n8215), .ZN(n8136) );
  INV_X1 U9643 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U9644 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  XNOR2_X1 U9645 ( .A(n8650), .B(n8179), .ZN(n8201) );
  NOR2_X1 U9646 ( .A1(n8217), .A2(n6193), .ZN(n8202) );
  AOI21_X1 U9647 ( .B1(n8200), .B2(n8201), .A(n8202), .ZN(n8137) );
  INV_X1 U9648 ( .A(n8137), .ZN(n8139) );
  NAND2_X1 U9649 ( .A1(n8139), .A2(n8138), .ZN(n8252) );
  INV_X1 U9650 ( .A(n8252), .ZN(n8144) );
  XNOR2_X1 U9651 ( .A(n8645), .B(n8179), .ZN(n8142) );
  AND2_X1 U9652 ( .A1(n8427), .A2(n8140), .ZN(n8141) );
  NAND2_X1 U9653 ( .A1(n8142), .A2(n8141), .ZN(n8175) );
  OAI21_X1 U9654 ( .B1(n8142), .B2(n8141), .A(n8175), .ZN(n8251) );
  NAND2_X1 U9655 ( .A1(n8253), .A2(n8175), .ZN(n8149) );
  XNOR2_X1 U9656 ( .A(n8638), .B(n8145), .ZN(n8147) );
  NAND2_X1 U9657 ( .A1(n8419), .A2(n8140), .ZN(n8146) );
  NOR2_X1 U9658 ( .A1(n8147), .A2(n8146), .ZN(n8174) );
  AOI21_X1 U9659 ( .B1(n8147), .B2(n8146), .A(n8174), .ZN(n8177) );
  NAND2_X1 U9660 ( .A1(n8149), .A2(n8177), .ZN(n8148) );
  OAI211_X1 U9661 ( .C1(n8149), .C2(n8177), .A(n8148), .B(n9589), .ZN(n8155)
         );
  OAI22_X1 U9662 ( .A1(n8434), .A2(n9593), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8150), .ZN(n8153) );
  OAI22_X1 U9663 ( .A1(n7465), .A2(n8244), .B1(n8245), .B2(n8151), .ZN(n8152)
         );
  AOI211_X1 U9664 ( .C1(n8638), .C2(n9584), .A(n8153), .B(n8152), .ZN(n8154)
         );
  NAND2_X1 U9665 ( .A1(n8155), .A2(n8154), .ZN(P2_U3216) );
  XNOR2_X1 U9666 ( .A(n8157), .B(n8156), .ZN(n8158) );
  XNOR2_X1 U9667 ( .A(n8159), .B(n8158), .ZN(n8165) );
  OAI22_X1 U9668 ( .A1(n9593), .A2(n8492), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8160), .ZN(n8163) );
  OAI22_X1 U9669 ( .A1(n8161), .A2(n8244), .B1(n8245), .B2(n8195), .ZN(n8162)
         );
  AOI211_X1 U9670 ( .C1(n8658), .C2(n9584), .A(n8163), .B(n8162), .ZN(n8164)
         );
  OAI21_X1 U9671 ( .B1(n8165), .B2(n8250), .A(n8164), .ZN(P2_U3218) );
  OAI21_X1 U9672 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8169) );
  NAND2_X1 U9673 ( .A1(n8169), .A2(n9589), .ZN(n8173) );
  INV_X1 U9674 ( .A(n8170), .ZN(n8558) );
  AND2_X1 U9675 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8397) );
  OAI22_X1 U9676 ( .A1(n8593), .A2(n8245), .B1(n8244), .B2(n8555), .ZN(n8171)
         );
  AOI211_X1 U9677 ( .C1(n8258), .C2(n8558), .A(n8397), .B(n8171), .ZN(n8172)
         );
  OAI211_X1 U9678 ( .C1(n8561), .C2(n9573), .A(n8173), .B(n8172), .ZN(P2_U3221) );
  INV_X1 U9679 ( .A(n8174), .ZN(n8176) );
  AND2_X1 U9680 ( .A1(n8175), .A2(n8176), .ZN(n8178) );
  NOR2_X1 U9681 ( .A1(n8415), .A2(n9751), .ZN(n8183) );
  INV_X1 U9682 ( .A(n8183), .ZN(n8181) );
  NAND2_X1 U9683 ( .A1(n8426), .A2(n8140), .ZN(n8180) );
  XNOR2_X1 U9684 ( .A(n8180), .B(n8179), .ZN(n8182) );
  MUX2_X1 U9685 ( .A(n8181), .B(n4621), .S(n8182), .Z(n8186) );
  MUX2_X1 U9686 ( .A(n8415), .B(n8183), .S(n8182), .Z(n8184) );
  OAI21_X1 U9687 ( .B1(n8415), .B2(n9573), .A(n8250), .ZN(n8185) );
  AOI22_X1 U9688 ( .A1(n8413), .A2(n8258), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8190) );
  AOI22_X1 U9689 ( .A1(n8188), .A2(n8418), .B1(n8187), .B2(n8419), .ZN(n8189)
         );
  XNOR2_X1 U9690 ( .A(n8192), .B(n8191), .ZN(n8199) );
  INV_X1 U9691 ( .A(n8523), .ZN(n8194) );
  OAI22_X1 U9692 ( .A1(n9593), .A2(n8194), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8193), .ZN(n8197) );
  OAI22_X1 U9693 ( .A1(n8555), .A2(n8245), .B1(n8244), .B2(n8195), .ZN(n8196)
         );
  AOI211_X1 U9694 ( .C1(n8668), .C2(n9584), .A(n8197), .B(n8196), .ZN(n8198)
         );
  OAI21_X1 U9695 ( .B1(n8199), .B2(n8250), .A(n8198), .ZN(P2_U3225) );
  XOR2_X1 U9696 ( .A(n8202), .B(n8201), .Z(n8203) );
  XNOR2_X1 U9697 ( .A(n8200), .B(n8203), .ZN(n8208) );
  AOI22_X1 U9698 ( .A1(n8427), .A2(n8573), .B1(n8501), .B2(n8571), .ZN(n8464)
         );
  OAI22_X1 U9699 ( .A1(n8464), .A2(n9586), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8204), .ZN(n8205) );
  AOI21_X1 U9700 ( .B1(n8467), .B2(n8258), .A(n8205), .ZN(n8207) );
  NAND2_X1 U9701 ( .A1(n8650), .A2(n9584), .ZN(n8206) );
  OAI211_X1 U9702 ( .C1(n8208), .C2(n8250), .A(n8207), .B(n8206), .ZN(P2_U3227) );
  XNOR2_X1 U9703 ( .A(n8210), .B(n8209), .ZN(n8214) );
  OAI22_X1 U9704 ( .A1(n9593), .A2(n8584), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8358), .ZN(n8212) );
  OAI22_X1 U9705 ( .A1(n8592), .A2(n8245), .B1(n8244), .B2(n8593), .ZN(n8211)
         );
  AOI211_X1 U9706 ( .C1(n8692), .C2(n9584), .A(n8212), .B(n8211), .ZN(n8213)
         );
  OAI21_X1 U9707 ( .B1(n8214), .B2(n8250), .A(n8213), .ZN(P2_U3230) );
  XNOR2_X1 U9708 ( .A(n8216), .B(n8215), .ZN(n8223) );
  OR2_X1 U9709 ( .A1(n8217), .A2(n9613), .ZN(n8219) );
  NAND2_X1 U9710 ( .A1(n8263), .A2(n8571), .ZN(n8218) );
  NAND2_X1 U9711 ( .A1(n8219), .A2(n8218), .ZN(n8482) );
  AOI22_X1 U9712 ( .A1(n8482), .A2(n9571), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8220) );
  OAI21_X1 U9713 ( .B1(n8476), .B2(n9593), .A(n8220), .ZN(n8221) );
  AOI21_X1 U9714 ( .B1(n8653), .B2(n9584), .A(n8221), .ZN(n8222) );
  OAI21_X1 U9715 ( .B1(n8223), .B2(n8250), .A(n8222), .ZN(P2_U3231) );
  XNOR2_X1 U9716 ( .A(n8225), .B(n8224), .ZN(n8231) );
  INV_X1 U9717 ( .A(n8544), .ZN(n8226) );
  OAI22_X1 U9718 ( .A1(n9593), .A2(n8226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9963), .ZN(n8229) );
  OAI22_X1 U9719 ( .A1(n8243), .A2(n8245), .B1(n8244), .B2(n8227), .ZN(n8228)
         );
  AOI211_X1 U9720 ( .C1(n8675), .C2(n9584), .A(n8229), .B(n8228), .ZN(n8230)
         );
  OAI21_X1 U9721 ( .B1(n8231), .B2(n8250), .A(n8230), .ZN(P2_U3235) );
  OAI21_X1 U9722 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8235) );
  NAND2_X1 U9723 ( .A1(n8235), .A2(n9589), .ZN(n8240) );
  INV_X1 U9724 ( .A(n8236), .ZN(n8508) );
  AOI22_X1 U9725 ( .A1(n8263), .A2(n8573), .B1(n8571), .B2(n8537), .ZN(n8514)
         );
  OAI22_X1 U9726 ( .A1(n9586), .A2(n8514), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8237), .ZN(n8238) );
  AOI21_X1 U9727 ( .B1(n8508), .B2(n8258), .A(n8238), .ZN(n8239) );
  OAI211_X1 U9728 ( .C1(n8510), .C2(n9573), .A(n8240), .B(n8239), .ZN(P2_U3237) );
  XNOR2_X1 U9729 ( .A(n8242), .B(n8241), .ZN(n8249) );
  AND2_X1 U9730 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8371) );
  OAI22_X1 U9731 ( .A1(n8598), .A2(n8245), .B1(n8244), .B2(n8243), .ZN(n8246)
         );
  AOI211_X1 U9732 ( .C1(n8258), .C2(n8566), .A(n8371), .B(n8246), .ZN(n8248)
         );
  NAND2_X1 U9733 ( .A1(n8685), .A2(n9584), .ZN(n8247) );
  OAI211_X1 U9734 ( .C1(n8249), .C2(n8250), .A(n8248), .B(n8247), .ZN(P2_U3240) );
  AOI21_X1 U9735 ( .B1(n8252), .B2(n8251), .A(n8250), .ZN(n8254) );
  NAND2_X1 U9736 ( .A1(n8254), .A2(n8253), .ZN(n8260) );
  INV_X1 U9737 ( .A(n8255), .ZN(n8452) );
  AOI22_X1 U9738 ( .A1(n8419), .A2(n8573), .B1(n8262), .B2(n8571), .ZN(n8447)
         );
  OAI22_X1 U9739 ( .A1(n8447), .A2(n9586), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8256), .ZN(n8257) );
  AOI21_X1 U9740 ( .B1(n8452), .B2(n8258), .A(n8257), .ZN(n8259) );
  OAI211_X1 U9741 ( .C1(n8455), .C2(n9573), .A(n8260), .B(n8259), .ZN(P2_U3242) );
  MUX2_X1 U9742 ( .A(n8261), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8280), .Z(
        P2_U3582) );
  MUX2_X1 U9743 ( .A(n8418), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8280), .Z(
        P2_U3581) );
  MUX2_X1 U9744 ( .A(n8426), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8280), .Z(
        P2_U3580) );
  MUX2_X1 U9745 ( .A(n8419), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8280), .Z(
        P2_U3579) );
  MUX2_X1 U9746 ( .A(n8427), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8280), .Z(
        P2_U3578) );
  MUX2_X1 U9747 ( .A(n8262), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8280), .Z(
        P2_U3577) );
  MUX2_X1 U9748 ( .A(n8501), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8280), .Z(
        P2_U3576) );
  MUX2_X1 U9749 ( .A(n8263), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8280), .Z(
        P2_U3575) );
  MUX2_X1 U9750 ( .A(n8529), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8280), .Z(
        P2_U3574) );
  MUX2_X1 U9751 ( .A(n8537), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8280), .Z(
        P2_U3573) );
  MUX2_X1 U9752 ( .A(n8528), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8280), .Z(
        P2_U3572) );
  MUX2_X1 U9753 ( .A(n8574), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8280), .Z(
        P2_U3571) );
  MUX2_X1 U9754 ( .A(n8264), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8280), .Z(
        P2_U3570) );
  MUX2_X1 U9755 ( .A(n8572), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8280), .Z(
        P2_U3569) );
  MUX2_X1 U9756 ( .A(n8265), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8280), .Z(
        P2_U3568) );
  MUX2_X1 U9757 ( .A(n8266), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8280), .Z(
        P2_U3567) );
  MUX2_X1 U9758 ( .A(n8267), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8280), .Z(
        P2_U3566) );
  MUX2_X1 U9759 ( .A(n8268), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8280), .Z(
        P2_U3565) );
  MUX2_X1 U9760 ( .A(n8269), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8280), .Z(
        P2_U3564) );
  MUX2_X1 U9761 ( .A(n8270), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8280), .Z(
        P2_U3563) );
  MUX2_X1 U9762 ( .A(n8271), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8280), .Z(
        P2_U3562) );
  MUX2_X1 U9763 ( .A(n8272), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8280), .Z(
        P2_U3561) );
  MUX2_X1 U9764 ( .A(n8273), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8280), .Z(
        P2_U3560) );
  MUX2_X1 U9765 ( .A(n8274), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8280), .Z(
        P2_U3559) );
  MUX2_X1 U9766 ( .A(n8275), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8280), .Z(
        P2_U3558) );
  MUX2_X1 U9767 ( .A(n8276), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8280), .Z(
        P2_U3557) );
  MUX2_X1 U9768 ( .A(n8277), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8280), .Z(
        P2_U3556) );
  MUX2_X1 U9769 ( .A(n8278), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8280), .Z(
        P2_U3555) );
  MUX2_X1 U9770 ( .A(n8279), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8280), .Z(
        P2_U3554) );
  MUX2_X1 U9771 ( .A(n8281), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8280), .Z(
        P2_U3552) );
  OAI211_X1 U9772 ( .C1(n8284), .C2(n8283), .A(n9598), .B(n8282), .ZN(n8294)
         );
  AOI21_X1 U9773 ( .B1(n9600), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8285), .ZN(
        n8293) );
  OR2_X1 U9774 ( .A1(n9595), .A2(n8286), .ZN(n8292) );
  AOI21_X1 U9775 ( .B1(n8289), .B2(n8288), .A(n8287), .ZN(n8290) );
  NAND2_X1 U9776 ( .A1(n9594), .A2(n8290), .ZN(n8291) );
  NAND4_X1 U9777 ( .A1(n8294), .A2(n8293), .A3(n8292), .A4(n8291), .ZN(
        P2_U3252) );
  OAI211_X1 U9778 ( .C1(n8297), .C2(n8296), .A(n9598), .B(n8295), .ZN(n8306)
         );
  AND2_X1 U9779 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9569) );
  AOI21_X1 U9780 ( .B1(n9600), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9569), .ZN(
        n8305) );
  OR2_X1 U9781 ( .A1(n9595), .A2(n8298), .ZN(n8304) );
  AOI21_X1 U9782 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8302) );
  NAND2_X1 U9783 ( .A1(n9594), .A2(n8302), .ZN(n8303) );
  NAND4_X1 U9784 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(
        P2_U3254) );
  OAI211_X1 U9785 ( .C1(n8309), .C2(n8308), .A(n9598), .B(n8307), .ZN(n8319)
         );
  AOI21_X1 U9786 ( .B1(n9600), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8310), .ZN(
        n8318) );
  OR2_X1 U9787 ( .A1(n9595), .A2(n8311), .ZN(n8317) );
  AOI21_X1 U9788 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(n8315) );
  NAND2_X1 U9789 ( .A1(n9594), .A2(n8315), .ZN(n8316) );
  NAND4_X1 U9790 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(
        P2_U3255) );
  INV_X1 U9791 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9317) );
  AOI211_X1 U9792 ( .C1(n8321), .C2(n9317), .A(n8335), .B(n9596), .ZN(n8332)
         );
  NOR2_X1 U9793 ( .A1(n8322), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8324) );
  NOR2_X1 U9794 ( .A1(n8324), .A2(n8323), .ZN(n8341) );
  XNOR2_X1 U9795 ( .A(n8341), .B(n8342), .ZN(n8325) );
  NOR2_X1 U9796 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8325), .ZN(n8343) );
  AOI21_X1 U9797 ( .B1(n8325), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8343), .ZN(
        n8326) );
  NOR2_X1 U9798 ( .A1(n8326), .A2(n8390), .ZN(n8331) );
  NOR2_X1 U9799 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8327), .ZN(n8328) );
  AOI21_X1 U9800 ( .B1(n9600), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8328), .ZN(
        n8329) );
  OAI21_X1 U9801 ( .B1(n9595), .B2(n8334), .A(n8329), .ZN(n8330) );
  OR3_X1 U9802 ( .A1(n8332), .A2(n8331), .A3(n8330), .ZN(P2_U3260) );
  NOR2_X1 U9803 ( .A1(n8334), .A2(n8333), .ZN(n8336) );
  XOR2_X1 U9804 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8360), .Z(n8337) );
  NAND2_X1 U9805 ( .A1(n8337), .A2(n8338), .ZN(n8359) );
  OAI21_X1 U9806 ( .B1(n8338), .B2(n8337), .A(n8359), .ZN(n8339) );
  NAND2_X1 U9807 ( .A1(n8339), .A2(n9594), .ZN(n8351) );
  AOI21_X1 U9808 ( .B1(n9600), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8340), .ZN(
        n8350) );
  NOR2_X1 U9809 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  NOR2_X1 U9810 ( .A1(n8344), .A2(n8343), .ZN(n8347) );
  INV_X1 U9811 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8345) );
  MUX2_X1 U9812 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8345), .S(n8360), .Z(n8346)
         );
  NAND2_X1 U9813 ( .A1(n8346), .A2(n8347), .ZN(n8352) );
  OAI211_X1 U9814 ( .C1(n8347), .C2(n8346), .A(n9598), .B(n8352), .ZN(n8349)
         );
  NAND2_X1 U9815 ( .A1(n9241), .A2(n8360), .ZN(n8348) );
  NAND4_X1 U9816 ( .A1(n8351), .A2(n8350), .A3(n8349), .A4(n8348), .ZN(
        P2_U3261) );
  NAND2_X1 U9817 ( .A1(n8360), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U9818 ( .A1(n8353), .A2(n8352), .ZN(n8357) );
  INV_X1 U9819 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8354) );
  MUX2_X1 U9820 ( .A(n8354), .B(P2_REG2_REG_17__SCAN_IN), .S(n8375), .Z(n8355)
         );
  INV_X1 U9821 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U9822 ( .A1(n8356), .A2(n8357), .ZN(n8368) );
  OAI211_X1 U9823 ( .C1(n8357), .C2(n8356), .A(n9598), .B(n8368), .ZN(n8366)
         );
  NOR2_X1 U9824 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8358), .ZN(n8364) );
  XNOR2_X1 U9825 ( .A(n8375), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8361) );
  AOI211_X1 U9826 ( .C1(n8362), .C2(n8361), .A(n8374), .B(n9596), .ZN(n8363)
         );
  AOI211_X1 U9827 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9600), .A(n8364), .B(
        n8363), .ZN(n8365) );
  OAI211_X1 U9828 ( .C1(n9595), .C2(n8367), .A(n8366), .B(n8365), .ZN(P2_U3262) );
  NAND2_X1 U9829 ( .A1(n8375), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U9830 ( .A1(n8369), .A2(n8368), .ZN(n8381) );
  XOR2_X1 U9831 ( .A(n8385), .B(n8381), .Z(n8370) );
  NAND2_X1 U9832 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8370), .ZN(n8382) );
  OAI211_X1 U9833 ( .C1(n8370), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9598), .B(
        n8382), .ZN(n8380) );
  AOI21_X1 U9834 ( .B1(n9600), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8371), .ZN(
        n8379) );
  OR2_X1 U9835 ( .A1(n9595), .A2(n8372), .ZN(n8378) );
  INV_X1 U9836 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8373) );
  XNOR2_X1 U9837 ( .A(n8385), .B(n8373), .ZN(n8388) );
  XNOR2_X1 U9838 ( .A(n8388), .B(n8387), .ZN(n8376) );
  NAND2_X1 U9839 ( .A1(n9594), .A2(n8376), .ZN(n8377) );
  NAND4_X1 U9840 ( .A1(n8380), .A2(n8379), .A3(n8378), .A4(n8377), .ZN(
        P2_U3263) );
  NAND2_X1 U9841 ( .A1(n8381), .A2(n8385), .ZN(n8383) );
  NAND2_X1 U9842 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  XOR2_X1 U9843 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8384), .Z(n8395) );
  INV_X1 U9844 ( .A(n8395), .ZN(n8391) );
  NOR2_X1 U9845 ( .A1(n8385), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8386) );
  XNOR2_X1 U9846 ( .A(n8389), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8392) );
  OAI22_X1 U9847 ( .A1(n8391), .A2(n8390), .B1(n9596), .B2(n8392), .ZN(n8396)
         );
  NAND2_X1 U9848 ( .A1(n9594), .A2(n8392), .ZN(n8393) );
  NAND2_X1 U9849 ( .A1(n8404), .A2(n8403), .ZN(n8402) );
  XNOR2_X1 U9850 ( .A(n8619), .B(n8402), .ZN(n8617) );
  NAND2_X1 U9851 ( .A1(n8617), .A2(n9668), .ZN(n8401) );
  NAND2_X1 U9852 ( .A1(n8399), .A2(n8398), .ZN(n8627) );
  NOR2_X1 U9853 ( .A1(n9669), .A2(n8627), .ZN(n8406) );
  AOI21_X1 U9854 ( .B1(n9669), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8406), .ZN(
        n8400) );
  OAI211_X1 U9855 ( .C1(n8619), .C2(n9673), .A(n8401), .B(n8400), .ZN(P2_U3265) );
  OAI21_X1 U9856 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8628) );
  NOR2_X1 U9857 ( .A1(n8404), .A2(n9673), .ZN(n8405) );
  AOI211_X1 U9858 ( .C1(n9669), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8406), .B(
        n8405), .ZN(n8407) );
  OAI21_X1 U9859 ( .B1(n9636), .B2(n8628), .A(n8407), .ZN(P2_U3266) );
  OAI21_X1 U9860 ( .B1(n8409), .B2(n8416), .A(n8408), .ZN(n8410) );
  INV_X1 U9861 ( .A(n8410), .ZN(n8636) );
  INV_X1 U9862 ( .A(n8411), .ZN(n8412) );
  AOI21_X1 U9863 ( .B1(n4621), .B2(n4620), .A(n8412), .ZN(n8633) );
  AOI22_X1 U9864 ( .A1(n8413), .A2(n9632), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9669), .ZN(n8414) );
  OAI21_X1 U9865 ( .B1(n8415), .B2(n9673), .A(n8414), .ZN(n8422) );
  XNOR2_X1 U9866 ( .A(n8417), .B(n8416), .ZN(n8420) );
  AOI222_X1 U9867 ( .A1(n9662), .A2(n8420), .B1(n8419), .B2(n8571), .C1(n8418), 
        .C2(n8573), .ZN(n8635) );
  NOR2_X1 U9868 ( .A1(n8635), .A2(n9669), .ZN(n8421) );
  AOI211_X1 U9869 ( .C1(n8633), .C2(n9668), .A(n8422), .B(n8421), .ZN(n8423)
         );
  OAI21_X1 U9870 ( .B1(n8636), .B2(n9676), .A(n8423), .ZN(P2_U3268) );
  XNOR2_X1 U9871 ( .A(n8425), .B(n8424), .ZN(n8428) );
  AOI222_X1 U9872 ( .A1(n9662), .A2(n8428), .B1(n8427), .B2(n8571), .C1(n8426), 
        .C2(n8573), .ZN(n8641) );
  OAI21_X1 U9873 ( .B1(n8431), .B2(n8430), .A(n8429), .ZN(n8637) );
  NAND2_X1 U9874 ( .A1(n8637), .A2(n9638), .ZN(n8439) );
  AOI21_X1 U9875 ( .B1(n8638), .B2(n8449), .A(n8432), .ZN(n8639) );
  INV_X1 U9876 ( .A(n8638), .ZN(n8433) );
  NOR2_X1 U9877 ( .A1(n8433), .A2(n9673), .ZN(n8437) );
  OAI22_X1 U9878 ( .A1(n9618), .A2(n8435), .B1(n8434), .B2(n9666), .ZN(n8436)
         );
  AOI211_X1 U9879 ( .C1(n8639), .C2(n9668), .A(n8437), .B(n8436), .ZN(n8438)
         );
  OAI211_X1 U9880 ( .C1(n9669), .C2(n8641), .A(n8439), .B(n8438), .ZN(P2_U3269) );
  OAI21_X1 U9881 ( .B1(n8441), .B2(n8446), .A(n8440), .ZN(n8442) );
  INV_X1 U9882 ( .A(n8442), .ZN(n8647) );
  INV_X1 U9883 ( .A(n8443), .ZN(n8444) );
  AOI21_X1 U9884 ( .B1(n8446), .B2(n8445), .A(n8444), .ZN(n8448) );
  OAI21_X1 U9885 ( .B1(n8448), .B2(n9644), .A(n8447), .ZN(n8643) );
  INV_X1 U9886 ( .A(n8449), .ZN(n8450) );
  AOI211_X1 U9887 ( .C1(n8645), .C2(n8451), .A(n9778), .B(n8450), .ZN(n8644)
         );
  NOR2_X1 U9888 ( .A1(n9669), .A2(n6138), .ZN(n8587) );
  NAND2_X1 U9889 ( .A1(n8644), .A2(n8587), .ZN(n8454) );
  AOI22_X1 U9890 ( .A1(n9669), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8452), .B2(
        n9632), .ZN(n8453) );
  OAI211_X1 U9891 ( .C1(n8455), .C2(n9673), .A(n8454), .B(n8453), .ZN(n8456)
         );
  AOI21_X1 U9892 ( .B1(n8643), .B2(n9618), .A(n8456), .ZN(n8457) );
  OAI21_X1 U9893 ( .B1(n8647), .B2(n9676), .A(n8457), .ZN(P2_U3270) );
  OAI21_X1 U9894 ( .B1(n8460), .B2(n8459), .A(n8458), .ZN(n8461) );
  INV_X1 U9895 ( .A(n8461), .ZN(n8652) );
  XNOR2_X1 U9896 ( .A(n8463), .B(n8462), .ZN(n8465) );
  OAI21_X1 U9897 ( .B1(n8465), .B2(n9644), .A(n8464), .ZN(n8648) );
  INV_X1 U9898 ( .A(n8650), .ZN(n8470) );
  AOI211_X1 U9899 ( .C1(n8650), .C2(n8474), .A(n9778), .B(n8466), .ZN(n8649)
         );
  NAND2_X1 U9900 ( .A1(n8649), .A2(n8587), .ZN(n8469) );
  AOI22_X1 U9901 ( .A1(n9669), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8467), .B2(
        n9632), .ZN(n8468) );
  OAI211_X1 U9902 ( .C1(n8470), .C2(n9673), .A(n8469), .B(n8468), .ZN(n8471)
         );
  AOI21_X1 U9903 ( .B1(n8648), .B2(n9618), .A(n8471), .ZN(n8472) );
  OAI21_X1 U9904 ( .B1(n8652), .B2(n9676), .A(n8472), .ZN(P2_U3271) );
  XOR2_X1 U9905 ( .A(n8473), .B(n8480), .Z(n8657) );
  INV_X1 U9906 ( .A(n8474), .ZN(n8475) );
  AOI21_X1 U9907 ( .B1(n8653), .B2(n8490), .A(n8475), .ZN(n8654) );
  INV_X1 U9908 ( .A(n8653), .ZN(n8479) );
  INV_X1 U9909 ( .A(n8476), .ZN(n8477) );
  AOI22_X1 U9910 ( .A1(n9669), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8477), .B2(
        n9632), .ZN(n8478) );
  OAI21_X1 U9911 ( .B1(n8479), .B2(n9673), .A(n8478), .ZN(n8486) );
  INV_X1 U9912 ( .A(n8480), .ZN(n8481) );
  AOI21_X1 U9913 ( .B1(n4432), .B2(n8481), .A(n9644), .ZN(n8484) );
  AOI21_X1 U9914 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8656) );
  NOR2_X1 U9915 ( .A1(n8656), .A2(n9669), .ZN(n8485) );
  AOI211_X1 U9916 ( .C1(n8654), .C2(n9668), .A(n8486), .B(n8485), .ZN(n8487)
         );
  OAI21_X1 U9917 ( .B1(n8657), .B2(n9676), .A(n8487), .ZN(P2_U3272) );
  OAI21_X1 U9918 ( .B1(n8489), .B2(n8497), .A(n8488), .ZN(n8662) );
  INV_X1 U9919 ( .A(n8490), .ZN(n8491) );
  AOI21_X1 U9920 ( .B1(n8658), .B2(n4628), .A(n8491), .ZN(n8659) );
  INV_X1 U9921 ( .A(n8492), .ZN(n8493) );
  AOI22_X1 U9922 ( .A1(n9669), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8493), .B2(
        n9632), .ZN(n8494) );
  OAI21_X1 U9923 ( .B1(n8495), .B2(n9673), .A(n8494), .ZN(n8504) );
  INV_X1 U9924 ( .A(n8496), .ZN(n8511) );
  OAI21_X1 U9925 ( .B1(n8511), .B2(n8498), .A(n8497), .ZN(n8500) );
  NAND2_X1 U9926 ( .A1(n8500), .A2(n8499), .ZN(n8502) );
  AOI222_X1 U9927 ( .A1(n9662), .A2(n8502), .B1(n8529), .B2(n8571), .C1(n8501), 
        .C2(n8573), .ZN(n8661) );
  NOR2_X1 U9928 ( .A1(n8661), .A2(n9669), .ZN(n8503) );
  AOI211_X1 U9929 ( .C1(n8659), .C2(n9668), .A(n8504), .B(n8503), .ZN(n8505)
         );
  OAI21_X1 U9930 ( .B1(n8662), .B2(n9676), .A(n8505), .ZN(P2_U3273) );
  XOR2_X1 U9931 ( .A(n8506), .B(n8513), .Z(n8667) );
  AOI21_X1 U9932 ( .B1(n8663), .B2(n8521), .A(n8507), .ZN(n8664) );
  AOI22_X1 U9933 ( .A1(n9669), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8508), .B2(
        n9632), .ZN(n8509) );
  OAI21_X1 U9934 ( .B1(n8510), .B2(n9673), .A(n8509), .ZN(n8518) );
  AOI211_X1 U9935 ( .C1(n8513), .C2(n8512), .A(n9644), .B(n8511), .ZN(n8516)
         );
  INV_X1 U9936 ( .A(n8514), .ZN(n8515) );
  NOR2_X1 U9937 ( .A1(n8516), .A2(n8515), .ZN(n8666) );
  NOR2_X1 U9938 ( .A1(n8666), .A2(n9669), .ZN(n8517) );
  AOI211_X1 U9939 ( .C1(n8664), .C2(n9668), .A(n8518), .B(n8517), .ZN(n8519)
         );
  OAI21_X1 U9940 ( .B1(n8667), .B2(n9676), .A(n8519), .ZN(P2_U3274) );
  XNOR2_X1 U9941 ( .A(n8520), .B(n8526), .ZN(n8672) );
  INV_X1 U9942 ( .A(n8521), .ZN(n8522) );
  AOI21_X1 U9943 ( .B1(n8668), .B2(n8541), .A(n8522), .ZN(n8669) );
  AOI22_X1 U9944 ( .A1(n9669), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8523), .B2(
        n9632), .ZN(n8524) );
  OAI21_X1 U9945 ( .B1(n8525), .B2(n9673), .A(n8524), .ZN(n8532) );
  XNOR2_X1 U9946 ( .A(n8527), .B(n8526), .ZN(n8530) );
  AOI222_X1 U9947 ( .A1(n9662), .A2(n8530), .B1(n8529), .B2(n8573), .C1(n8528), 
        .C2(n8571), .ZN(n8671) );
  NOR2_X1 U9948 ( .A1(n8671), .A2(n9669), .ZN(n8531) );
  AOI211_X1 U9949 ( .C1(n8669), .C2(n9668), .A(n8532), .B(n8531), .ZN(n8533)
         );
  OAI21_X1 U9950 ( .B1(n8672), .B2(n9676), .A(n8533), .ZN(P2_U3275) );
  NAND2_X1 U9951 ( .A1(n8551), .A2(n8534), .ZN(n8536) );
  XNOR2_X1 U9952 ( .A(n8536), .B(n8535), .ZN(n8538) );
  AOI222_X1 U9953 ( .A1(n9662), .A2(n8538), .B1(n8537), .B2(n8573), .C1(n8574), 
        .C2(n8571), .ZN(n8678) );
  OR2_X1 U9954 ( .A1(n8540), .A2(n8539), .ZN(n8674) );
  NAND3_X1 U9955 ( .A1(n8674), .A2(n8673), .A3(n9638), .ZN(n8549) );
  INV_X1 U9956 ( .A(n8556), .ZN(n8543) );
  INV_X1 U9957 ( .A(n8541), .ZN(n8542) );
  AOI21_X1 U9958 ( .B1(n8675), .B2(n8543), .A(n8542), .ZN(n8676) );
  AOI22_X1 U9959 ( .A1(n9669), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8544), .B2(
        n9632), .ZN(n8545) );
  OAI21_X1 U9960 ( .B1(n8546), .B2(n9673), .A(n8545), .ZN(n8547) );
  AOI21_X1 U9961 ( .B1(n8676), .B2(n9668), .A(n8547), .ZN(n8548) );
  OAI211_X1 U9962 ( .C1(n9669), .C2(n8678), .A(n8549), .B(n8548), .ZN(P2_U3276) );
  XNOR2_X1 U9963 ( .A(n8550), .B(n8553), .ZN(n8684) );
  AOI21_X1 U9964 ( .B1(n8553), .B2(n8552), .A(n7498), .ZN(n8554) );
  OAI222_X1 U9965 ( .A1(n9613), .A2(n8555), .B1(n9611), .B2(n8593), .C1(n9644), 
        .C2(n8554), .ZN(n8680) );
  INV_X1 U9966 ( .A(n8565), .ZN(n8557) );
  AOI211_X1 U9967 ( .C1(n8682), .C2(n8557), .A(n9778), .B(n8556), .ZN(n8681)
         );
  NAND2_X1 U9968 ( .A1(n8681), .A2(n8587), .ZN(n8560) );
  AOI22_X1 U9969 ( .A1(n9669), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8558), .B2(
        n9632), .ZN(n8559) );
  OAI211_X1 U9970 ( .C1(n8561), .C2(n9673), .A(n8560), .B(n8559), .ZN(n8562)
         );
  AOI21_X1 U9971 ( .B1(n8680), .B2(n9618), .A(n8562), .ZN(n8563) );
  OAI21_X1 U9972 ( .B1(n8684), .B2(n9676), .A(n8563), .ZN(P2_U3277) );
  XNOR2_X1 U9973 ( .A(n8564), .B(n8569), .ZN(n8689) );
  AOI21_X1 U9974 ( .B1(n8685), .B2(n8582), .A(n8565), .ZN(n8686) );
  AOI22_X1 U9975 ( .A1(n9669), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8566), .B2(
        n9632), .ZN(n8567) );
  OAI21_X1 U9976 ( .B1(n8568), .B2(n9673), .A(n8567), .ZN(n8577) );
  XOR2_X1 U9977 ( .A(n8570), .B(n8569), .Z(n8575) );
  AOI222_X1 U9978 ( .A1(n9662), .A2(n8575), .B1(n8574), .B2(n8573), .C1(n8572), 
        .C2(n8571), .ZN(n8688) );
  NOR2_X1 U9979 ( .A1(n8688), .A2(n9669), .ZN(n8576) );
  AOI211_X1 U9980 ( .C1(n8686), .C2(n9668), .A(n8577), .B(n8576), .ZN(n8578)
         );
  OAI21_X1 U9981 ( .B1(n8689), .B2(n9676), .A(n8578), .ZN(P2_U3278) );
  OAI21_X1 U9982 ( .B1(n8580), .B2(n8589), .A(n8579), .ZN(n8581) );
  INV_X1 U9983 ( .A(n8581), .ZN(n8694) );
  INV_X1 U9984 ( .A(n8582), .ZN(n8583) );
  AOI211_X1 U9985 ( .C1(n8692), .C2(n8612), .A(n9778), .B(n8583), .ZN(n8691)
         );
  NOR2_X1 U9986 ( .A1(n4615), .A2(n9673), .ZN(n8586) );
  OAI22_X1 U9987 ( .A1(n9618), .A2(n8354), .B1(n8584), .B2(n9666), .ZN(n8585)
         );
  AOI211_X1 U9988 ( .C1(n8691), .C2(n8587), .A(n8586), .B(n8585), .ZN(n8595)
         );
  NAND2_X1 U9989 ( .A1(n8596), .A2(n8588), .ZN(n8590) );
  XNOR2_X1 U9990 ( .A(n8590), .B(n8589), .ZN(n8591) );
  OAI222_X1 U9991 ( .A1(n9613), .A2(n8593), .B1(n9611), .B2(n8592), .C1(n8591), 
        .C2(n9644), .ZN(n8690) );
  NAND2_X1 U9992 ( .A1(n8690), .A2(n9618), .ZN(n8594) );
  OAI211_X1 U9993 ( .C1(n8694), .C2(n9676), .A(n8595), .B(n8594), .ZN(P2_U3279) );
  OAI21_X1 U9994 ( .B1(n8597), .B2(n4473), .A(n8596), .ZN(n8606) );
  OAI22_X1 U9995 ( .A1(n8599), .A2(n9611), .B1(n8598), .B2(n9613), .ZN(n8605)
         );
  NOR2_X1 U9996 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  NOR2_X1 U9997 ( .A1(n8699), .A2(n9640), .ZN(n8604) );
  AOI211_X1 U9998 ( .C1(n9662), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8698)
         );
  NAND2_X1 U9999 ( .A1(n9669), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8607) );
  OAI21_X1 U10000 ( .B1(n9666), .B2(n8608), .A(n8607), .ZN(n8609) );
  AOI21_X1 U10001 ( .B1(n8695), .B2(n9631), .A(n8609), .ZN(n8614) );
  NAND2_X1 U10002 ( .A1(n8610), .A2(n8695), .ZN(n8611) );
  AND2_X1 U10003 ( .A1(n8612), .A2(n8611), .ZN(n8696) );
  NAND2_X1 U10004 ( .A1(n8696), .A2(n9668), .ZN(n8613) );
  OAI211_X1 U10005 ( .C1(n8699), .C2(n9648), .A(n8614), .B(n8613), .ZN(n8615)
         );
  INV_X1 U10006 ( .A(n8615), .ZN(n8616) );
  OAI21_X1 U10007 ( .B1(n8698), .B2(n9669), .A(n8616), .ZN(P2_U3280) );
  NAND2_X1 U10008 ( .A1(n8617), .A2(n9752), .ZN(n8618) );
  OAI211_X1 U10009 ( .C1(n8619), .C2(n9776), .A(n8618), .B(n8627), .ZN(n8705)
         );
  NAND2_X1 U10010 ( .A1(n8621), .A2(n8620), .ZN(n8623) );
  NOR2_X1 U10011 ( .A1(n8702), .A2(n8700), .ZN(n8624) );
  MUX2_X1 U10012 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8705), .S(n9803), .Z(
        P2_U3551) );
  NAND2_X1 U10013 ( .A1(n8625), .A2(n9751), .ZN(n8626) );
  OAI211_X1 U10014 ( .C1(n8628), .C2(n9778), .A(n8627), .B(n8626), .ZN(n8706)
         );
  MUX2_X1 U10015 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8706), .S(n9803), .Z(
        P2_U3550) );
  AOI22_X1 U10016 ( .A1(n8630), .A2(n9752), .B1(n9751), .B2(n8629), .ZN(n8631)
         );
  OAI211_X1 U10017 ( .C1(n8632), .C2(n9740), .A(n4413), .B(n8631), .ZN(n8707)
         );
  MUX2_X1 U10018 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8707), .S(n9803), .Z(
        P2_U3549) );
  AOI22_X1 U10019 ( .A1(n8633), .A2(n9752), .B1(n9751), .B2(n4621), .ZN(n8634)
         );
  OAI211_X1 U10020 ( .C1(n8636), .C2(n9740), .A(n8635), .B(n8634), .ZN(n8708)
         );
  MUX2_X1 U10021 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8708), .S(n9803), .Z(
        P2_U3548) );
  INV_X1 U10022 ( .A(n8637), .ZN(n8642) );
  AOI22_X1 U10023 ( .A1(n8639), .A2(n9752), .B1(n9751), .B2(n8638), .ZN(n8640)
         );
  OAI211_X1 U10024 ( .C1(n8642), .C2(n9740), .A(n8641), .B(n8640), .ZN(n8709)
         );
  MUX2_X1 U10025 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8709), .S(n9803), .Z(
        P2_U3547) );
  AOI211_X1 U10026 ( .C1(n9751), .C2(n8645), .A(n8644), .B(n8643), .ZN(n8646)
         );
  OAI21_X1 U10027 ( .B1(n8647), .B2(n9740), .A(n8646), .ZN(n8710) );
  MUX2_X1 U10028 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8710), .S(n9803), .Z(
        P2_U3546) );
  AOI211_X1 U10029 ( .C1(n9751), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8651)
         );
  OAI21_X1 U10030 ( .B1(n8652), .B2(n9740), .A(n8651), .ZN(n8711) );
  MUX2_X1 U10031 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8711), .S(n9803), .Z(
        P2_U3545) );
  AOI22_X1 U10032 ( .A1(n8654), .A2(n9752), .B1(n9751), .B2(n8653), .ZN(n8655)
         );
  OAI211_X1 U10033 ( .C1(n8657), .C2(n9740), .A(n8656), .B(n8655), .ZN(n8712)
         );
  MUX2_X1 U10034 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8712), .S(n9803), .Z(
        P2_U3544) );
  AOI22_X1 U10035 ( .A1(n8659), .A2(n9752), .B1(n9751), .B2(n8658), .ZN(n8660)
         );
  OAI211_X1 U10036 ( .C1(n8662), .C2(n9740), .A(n8661), .B(n8660), .ZN(n8713)
         );
  MUX2_X1 U10037 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8713), .S(n9803), .Z(
        P2_U3543) );
  AOI22_X1 U10038 ( .A1(n8664), .A2(n9752), .B1(n9751), .B2(n8663), .ZN(n8665)
         );
  OAI211_X1 U10039 ( .C1(n8667), .C2(n9740), .A(n8666), .B(n8665), .ZN(n8714)
         );
  MUX2_X1 U10040 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8714), .S(n9803), .Z(
        P2_U3542) );
  AOI22_X1 U10041 ( .A1(n8669), .A2(n9752), .B1(n9751), .B2(n8668), .ZN(n8670)
         );
  OAI211_X1 U10042 ( .C1(n8672), .C2(n9740), .A(n8671), .B(n8670), .ZN(n8715)
         );
  MUX2_X1 U10043 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8715), .S(n9803), .Z(
        P2_U3541) );
  NAND3_X1 U10044 ( .A1(n8674), .A2(n8673), .A3(n9783), .ZN(n8679) );
  AOI22_X1 U10045 ( .A1(n8676), .A2(n9752), .B1(n9751), .B2(n8675), .ZN(n8677)
         );
  NAND3_X1 U10046 ( .A1(n8679), .A2(n8678), .A3(n8677), .ZN(n8716) );
  MUX2_X1 U10047 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8716), .S(n9803), .Z(
        P2_U3540) );
  AOI211_X1 U10048 ( .C1(n9751), .C2(n8682), .A(n8681), .B(n8680), .ZN(n8683)
         );
  OAI21_X1 U10049 ( .B1(n9740), .B2(n8684), .A(n8683), .ZN(n8717) );
  MUX2_X1 U10050 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8717), .S(n9803), .Z(
        P2_U3539) );
  AOI22_X1 U10051 ( .A1(n8686), .A2(n9752), .B1(n9751), .B2(n8685), .ZN(n8687)
         );
  OAI211_X1 U10052 ( .C1(n8689), .C2(n9740), .A(n8688), .B(n8687), .ZN(n8718)
         );
  MUX2_X1 U10053 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8718), .S(n9803), .Z(
        P2_U3538) );
  AOI211_X1 U10054 ( .C1(n9751), .C2(n8692), .A(n8691), .B(n8690), .ZN(n8693)
         );
  OAI21_X1 U10055 ( .B1(n8694), .B2(n9740), .A(n8693), .ZN(n8719) );
  MUX2_X1 U10056 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8719), .S(n9803), .Z(
        P2_U3537) );
  AOI22_X1 U10057 ( .A1(n8696), .A2(n9752), .B1(n9751), .B2(n8695), .ZN(n8697)
         );
  OAI211_X1 U10058 ( .C1(n9755), .C2(n8699), .A(n8698), .B(n8697), .ZN(n8720)
         );
  MUX2_X1 U10059 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8720), .S(n9803), .Z(
        P2_U3536) );
  INV_X1 U10060 ( .A(n8700), .ZN(n8701) );
  NOR2_X1 U10061 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  MUX2_X1 U10062 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8705), .S(n9785), .Z(
        P2_U3519) );
  MUX2_X1 U10063 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8706), .S(n9785), .Z(
        P2_U3518) );
  MUX2_X1 U10064 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8707), .S(n9785), .Z(
        P2_U3517) );
  MUX2_X1 U10065 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8708), .S(n9785), .Z(
        P2_U3516) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8709), .S(n9785), .Z(
        P2_U3515) );
  MUX2_X1 U10067 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8710), .S(n9785), .Z(
        P2_U3514) );
  MUX2_X1 U10068 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8711), .S(n9785), .Z(
        P2_U3513) );
  MUX2_X1 U10069 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8712), .S(n9785), .Z(
        P2_U3512) );
  MUX2_X1 U10070 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8713), .S(n9785), .Z(
        P2_U3511) );
  MUX2_X1 U10071 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8714), .S(n9785), .Z(
        P2_U3510) );
  MUX2_X1 U10072 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8715), .S(n9785), .Z(
        P2_U3509) );
  MUX2_X1 U10073 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8716), .S(n9785), .Z(
        P2_U3508) );
  MUX2_X1 U10074 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8717), .S(n9785), .Z(
        P2_U3507) );
  MUX2_X1 U10075 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8718), .S(n9785), .Z(
        P2_U3505) );
  MUX2_X1 U10076 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8719), .S(n9785), .Z(
        P2_U3502) );
  MUX2_X1 U10077 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8720), .S(n9785), .Z(
        P2_U3499) );
  INV_X1 U10078 ( .A(n8721), .ZN(n9223) );
  NOR4_X1 U10079 ( .A1(n8723), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8722), .A4(
        P2_U3152), .ZN(n8724) );
  AOI21_X1 U10080 ( .B1(n8725), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8724), .ZN(
        n8726) );
  OAI21_X1 U10081 ( .B1(n9223), .B2(n7895), .A(n8726), .ZN(P2_U3327) );
  OAI222_X1 U10082 ( .A1(n8730), .A2(P2_U3152), .B1(n7895), .B2(n8729), .C1(
        n8728), .C2(n8727), .ZN(P2_U3329) );
  MUX2_X1 U10083 ( .A(n8731), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10084 ( .A(n8732), .ZN(n8733) );
  NAND2_X1 U10085 ( .A1(n8734), .A2(n8733), .ZN(n8736) );
  XNOR2_X1 U10086 ( .A(n8736), .B(n8735), .ZN(n8743) );
  OAI22_X1 U10087 ( .A1(n8984), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8737), .ZN(n8740) );
  NOR2_X1 U10088 ( .A1(n8868), .A2(n8738), .ZN(n8739) );
  AOI211_X1 U10089 ( .C1(n8987), .C2(n8863), .A(n8740), .B(n8739), .ZN(n8742)
         );
  NAND2_X1 U10090 ( .A1(n9156), .A2(n8870), .ZN(n8741) );
  OAI211_X1 U10091 ( .C1(n8743), .C2(n8872), .A(n8742), .B(n8741), .ZN(
        P1_U3214) );
  OAI21_X1 U10092 ( .B1(n8746), .B2(n8745), .A(n8744), .ZN(n8747) );
  NAND2_X1 U10093 ( .A1(n8747), .A2(n8849), .ZN(n8752) );
  OAI22_X1 U10094 ( .A1(n9074), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8748), .ZN(n8750) );
  NOR2_X1 U10095 ( .A1(n8868), .A2(n9046), .ZN(n8749) );
  AOI211_X1 U10096 ( .C1(n9048), .C2(n8863), .A(n8750), .B(n8749), .ZN(n8751)
         );
  OAI211_X1 U10097 ( .C1(n9051), .C2(n8859), .A(n8752), .B(n8751), .ZN(
        P1_U3217) );
  NAND2_X1 U10098 ( .A1(n9130), .A2(n8758), .ZN(n8755) );
  NAND2_X1 U10099 ( .A1(n8934), .A2(n8753), .ZN(n8754) );
  NAND2_X1 U10100 ( .A1(n8755), .A2(n8754), .ZN(n8757) );
  XNOR2_X1 U10101 ( .A(n8757), .B(n8756), .ZN(n8761) );
  AOI22_X1 U10102 ( .A1(n9130), .A2(n8759), .B1(n8758), .B2(n8934), .ZN(n8760)
         );
  XNOR2_X1 U10103 ( .A(n8761), .B(n8760), .ZN(n8768) );
  NAND3_X1 U10104 ( .A1(n8762), .A2(n8849), .A3(n8768), .ZN(n8771) );
  AOI22_X1 U10105 ( .A1(n8874), .A2(n8839), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8763) );
  OAI21_X1 U10106 ( .B1(n8854), .B2(n8852), .A(n8763), .ZN(n8765) );
  NOR2_X1 U10107 ( .A1(n8903), .A2(n8859), .ZN(n8764) );
  AOI211_X1 U10108 ( .C1(n8766), .C2(n8863), .A(n8765), .B(n8764), .ZN(n8770)
         );
  NAND3_X1 U10109 ( .A1(n8768), .A2(n8849), .A3(n8767), .ZN(n8769) );
  NAND4_X1 U10110 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(
        P1_U3218) );
  XOR2_X1 U10111 ( .A(n8773), .B(n8774), .Z(n8779) );
  NAND2_X1 U10112 ( .A1(n8863), .A2(n9010), .ZN(n8776) );
  AOI22_X1 U10113 ( .A1(n9016), .A2(n8865), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8775) );
  OAI211_X1 U10114 ( .C1(n8984), .C2(n8868), .A(n8776), .B(n8775), .ZN(n8777)
         );
  AOI21_X1 U10115 ( .B1(n9165), .B2(n8870), .A(n8777), .ZN(n8778) );
  OAI21_X1 U10116 ( .B1(n8779), .B2(n8872), .A(n8778), .ZN(P1_U3221) );
  INV_X1 U10117 ( .A(n9144), .ZN(n8956) );
  OAI21_X1 U10118 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8783) );
  NAND2_X1 U10119 ( .A1(n8783), .A2(n8849), .ZN(n8789) );
  INV_X1 U10120 ( .A(n8784), .ZN(n8954) );
  AOI22_X1 U10121 ( .A1(n4868), .A2(n8865), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8785) );
  OAI21_X1 U10122 ( .B1(n8786), .B2(n8868), .A(n8785), .ZN(n8787) );
  AOI21_X1 U10123 ( .B1(n8954), .B2(n8863), .A(n8787), .ZN(n8788) );
  OAI211_X1 U10124 ( .C1(n8956), .C2(n8859), .A(n8789), .B(n8788), .ZN(
        P1_U3223) );
  OAI21_X1 U10125 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8793) );
  NAND2_X1 U10126 ( .A1(n8793), .A2(n8849), .ZN(n8797) );
  AOI22_X1 U10127 ( .A1(n8865), .A2(n8877), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8794) );
  OAI21_X1 U10128 ( .B1(n9088), .B2(n8868), .A(n8794), .ZN(n8795) );
  AOI21_X1 U10129 ( .B1(n9092), .B2(n8863), .A(n8795), .ZN(n8796) );
  OAI211_X1 U10130 ( .C1(n9095), .C2(n8859), .A(n8797), .B(n8796), .ZN(
        P1_U3224) );
  OAI21_X1 U10131 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8801) );
  NAND2_X1 U10132 ( .A1(n8801), .A2(n8849), .ZN(n8805) );
  OAI22_X1 U10133 ( .A1(n9103), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10033), .ZN(n8803) );
  NOR2_X1 U10134 ( .A1(n8868), .A2(n9074), .ZN(n8802) );
  AOI211_X1 U10135 ( .C1(n9076), .C2(n8863), .A(n8803), .B(n8802), .ZN(n8804)
         );
  OAI211_X1 U10136 ( .C1(n9079), .C2(n8859), .A(n8805), .B(n8804), .ZN(
        P1_U3226) );
  INV_X1 U10137 ( .A(n8806), .ZN(n8807) );
  AOI21_X1 U10138 ( .B1(n8809), .B2(n8808), .A(n8807), .ZN(n8815) );
  NAND2_X1 U10139 ( .A1(n8969), .A2(n8839), .ZN(n8811) );
  AOI22_X1 U10140 ( .A1(n8865), .A2(n9000), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8810) );
  OAI211_X1 U10141 ( .C1(n8812), .C2(n8974), .A(n8811), .B(n8810), .ZN(n8813)
         );
  AOI21_X1 U10142 ( .B1(n9150), .B2(n8870), .A(n8813), .ZN(n8814) );
  OAI21_X1 U10143 ( .B1(n8815), .B2(n8872), .A(n8814), .ZN(P1_U3227) );
  NAND2_X1 U10144 ( .A1(n4476), .A2(n8816), .ZN(n8817) );
  XNOR2_X1 U10145 ( .A(n8818), .B(n8817), .ZN(n8823) );
  NAND2_X1 U10146 ( .A1(n8863), .A2(n9026), .ZN(n8820) );
  AOI22_X1 U10147 ( .A1(n8865), .A2(n9062), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8819) );
  OAI211_X1 U10148 ( .C1(n9029), .C2(n8868), .A(n8820), .B(n8819), .ZN(n8821)
         );
  AOI21_X1 U10149 ( .B1(n9169), .B2(n8870), .A(n8821), .ZN(n8822) );
  OAI21_X1 U10150 ( .B1(n8823), .B2(n8872), .A(n8822), .ZN(P1_U3231) );
  NOR2_X1 U10151 ( .A1(n8825), .A2(n8824), .ZN(n8827) );
  XNOR2_X1 U10152 ( .A(n8827), .B(n8826), .ZN(n8828) );
  NAND2_X1 U10153 ( .A1(n8828), .A2(n8849), .ZN(n8833) );
  OAI22_X1 U10154 ( .A1(n9029), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8829), .ZN(n8831) );
  NOR2_X1 U10155 ( .A1(n8868), .A2(n10145), .ZN(n8830) );
  AOI211_X1 U10156 ( .C1(n8995), .C2(n8863), .A(n8831), .B(n8830), .ZN(n8832)
         );
  OAI211_X1 U10157 ( .C1(n8997), .C2(n8859), .A(n8833), .B(n8832), .ZN(
        P1_U3233) );
  INV_X1 U10158 ( .A(n8834), .ZN(n8835) );
  NOR2_X1 U10159 ( .A1(n8836), .A2(n8835), .ZN(n8838) );
  XNOR2_X1 U10160 ( .A(n8838), .B(n8837), .ZN(n8844) );
  NAND2_X1 U10161 ( .A1(n8839), .A2(n9062), .ZN(n8840) );
  NAND2_X1 U10162 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9489) );
  OAI211_X1 U10163 ( .C1(n9088), .C2(n8852), .A(n8840), .B(n9489), .ZN(n8842)
         );
  NOR2_X1 U10164 ( .A1(n4573), .A2(n8859), .ZN(n8841) );
  AOI211_X1 U10165 ( .C1(n9057), .C2(n8863), .A(n8842), .B(n8841), .ZN(n8843)
         );
  OAI21_X1 U10166 ( .B1(n8844), .B2(n8872), .A(n8843), .ZN(P1_U3236) );
  INV_X1 U10167 ( .A(n8780), .ZN(n8847) );
  OAI21_X1 U10168 ( .B1(n8847), .B2(n8846), .A(n8845), .ZN(n8850) );
  NAND3_X1 U10169 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n8858) );
  OAI22_X1 U10170 ( .A1(n8853), .A2(n8852), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8851), .ZN(n8856) );
  NOR2_X1 U10171 ( .A1(n8854), .A2(n8868), .ZN(n8855) );
  AOI211_X1 U10172 ( .C1(n8942), .C2(n8863), .A(n8856), .B(n8855), .ZN(n8857)
         );
  OAI211_X1 U10173 ( .C1(n8944), .C2(n8859), .A(n8858), .B(n8857), .ZN(
        P1_U3238) );
  NOR2_X1 U10174 ( .A1(n8860), .A2(n4466), .ZN(n8862) );
  XNOR2_X1 U10175 ( .A(n8862), .B(n8861), .ZN(n8873) );
  NAND2_X1 U10176 ( .A1(n8863), .A2(n9107), .ZN(n8867) );
  AOI21_X1 U10177 ( .B1(n8865), .B2(n8878), .A(n8864), .ZN(n8866) );
  OAI211_X1 U10178 ( .C1(n9103), .C2(n8868), .A(n8867), .B(n8866), .ZN(n8869)
         );
  AOI21_X1 U10179 ( .B1(n9196), .B2(n8870), .A(n8869), .ZN(n8871) );
  OAI21_X1 U10180 ( .B1(n8873), .B2(n8872), .A(n8871), .ZN(P1_U3239) );
  MUX2_X1 U10181 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8913), .S(n10144), .Z(
        P1_U3585) );
  MUX2_X1 U10182 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8874), .S(n10144), .Z(
        P1_U3584) );
  MUX2_X1 U10183 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8934), .S(n10144), .Z(
        P1_U3583) );
  MUX2_X1 U10184 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8947), .S(n10144), .Z(
        P1_U3582) );
  MUX2_X1 U10185 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8959), .S(n10144), .Z(
        P1_U3581) );
  MUX2_X1 U10186 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8969), .S(n10144), .Z(
        P1_U3580) );
  MUX2_X1 U10187 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n4868), .S(n10144), .Z(
        P1_U3579) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9017), .S(n10144), .Z(
        P1_U3577) );
  INV_X1 U10189 ( .A(n9029), .ZN(n9001) );
  MUX2_X1 U10190 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9001), .S(n10144), .Z(
        P1_U3576) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9016), .S(n10144), .Z(
        P1_U3575) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9062), .S(n10144), .Z(
        P1_U3574) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8875), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9063), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8876), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10196 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8877), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10197 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8878), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8879), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10199 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8880), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9252), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8881), .S(n10144), .Z(
        P1_U3565) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9253), .S(n10144), .Z(
        P1_U3564) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8882), .S(n10144), .Z(
        P1_U3563) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8883), .S(n10144), .Z(
        P1_U3562) );
  MUX2_X1 U10205 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8884), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8885), .S(n10144), .Z(
        P1_U3560) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8886), .S(n10144), .Z(
        P1_U3559) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8887), .S(n10144), .Z(
        P1_U3558) );
  MUX2_X1 U10209 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5631), .S(n10144), .Z(
        P1_U3557) );
  MUX2_X1 U10210 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5613), .S(n10144), .Z(
        P1_U3556) );
  AOI211_X1 U10211 ( .C1(n8890), .C2(n8889), .A(n8888), .B(n9488), .ZN(n8900)
         );
  INV_X1 U10212 ( .A(n8891), .ZN(n8898) );
  AOI211_X1 U10213 ( .C1(n8894), .C2(n8893), .A(n8892), .B(n9381), .ZN(n8895)
         );
  INV_X1 U10214 ( .A(n8895), .ZN(n8897) );
  NAND2_X1 U10215 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8896) );
  OAI211_X1 U10216 ( .C1(n9408), .C2(n8898), .A(n8897), .B(n8896), .ZN(n8899)
         );
  AOI211_X1 U10217 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9495), .A(n8900), .B(
        n8899), .ZN(n8901) );
  INV_X1 U10218 ( .A(n8901), .ZN(P1_U3258) );
  XNOR2_X1 U10219 ( .A(n8906), .B(n8905), .ZN(n9120) );
  INV_X1 U10220 ( .A(n9120), .ZN(n8925) );
  INV_X1 U10221 ( .A(n8907), .ZN(n8908) );
  AOI21_X1 U10222 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8912) );
  XNOR2_X1 U10223 ( .A(n8912), .B(n8911), .ZN(n8916) );
  AOI22_X1 U10224 ( .A1(n8934), .A2(n9254), .B1(n8914), .B2(n8913), .ZN(n8915)
         );
  OAI21_X1 U10225 ( .B1(n8916), .B2(n9256), .A(n8915), .ZN(n9123) );
  AOI21_X1 U10226 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n9121) );
  NAND2_X1 U10227 ( .A1(n9121), .A2(n9068), .ZN(n8922) );
  AOI22_X1 U10228 ( .A1(n8920), .A2(n9261), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9513), .ZN(n8921) );
  OAI211_X1 U10229 ( .C1(n9122), .C2(n9110), .A(n8922), .B(n8921), .ZN(n8923)
         );
  AOI21_X1 U10230 ( .B1(n9123), .B2(n9081), .A(n8923), .ZN(n8924) );
  OAI21_X1 U10231 ( .B1(n8925), .B2(n9114), .A(n8924), .ZN(P1_U3355) );
  XNOR2_X1 U10232 ( .A(n8927), .B(n8926), .ZN(n9138) );
  AOI21_X1 U10233 ( .B1(n9134), .B2(n8940), .A(n8928), .ZN(n9135) );
  INV_X1 U10234 ( .A(n8929), .ZN(n8930) );
  AOI22_X1 U10235 ( .A1(n8930), .A2(n9261), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9513), .ZN(n8931) );
  OAI21_X1 U10236 ( .B1(n4743), .B2(n9110), .A(n8931), .ZN(n8937) );
  XNOR2_X1 U10237 ( .A(n8933), .B(n8932), .ZN(n8935) );
  AOI222_X1 U10238 ( .A1(n9065), .A2(n8935), .B1(n8934), .B2(n9251), .C1(n8959), .C2(n9254), .ZN(n9137) );
  NOR2_X1 U10239 ( .A1(n9137), .A2(n9513), .ZN(n8936) );
  AOI211_X1 U10240 ( .C1(n9068), .C2(n9135), .A(n8937), .B(n8936), .ZN(n8938)
         );
  OAI21_X1 U10241 ( .B1(n9138), .B2(n9114), .A(n8938), .ZN(P1_U3264) );
  XOR2_X1 U10242 ( .A(n8946), .B(n8939), .Z(n9143) );
  INV_X1 U10243 ( .A(n8940), .ZN(n8941) );
  AOI21_X1 U10244 ( .B1(n9139), .B2(n8953), .A(n8941), .ZN(n9140) );
  AOI22_X1 U10245 ( .A1(n9513), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n8942), .B2(
        n9261), .ZN(n8943) );
  OAI21_X1 U10246 ( .B1(n8944), .B2(n9110), .A(n8943), .ZN(n8950) );
  XOR2_X1 U10247 ( .A(n8946), .B(n8945), .Z(n8948) );
  AOI222_X1 U10248 ( .A1(n9065), .A2(n8948), .B1(n8947), .B2(n9251), .C1(n8969), .C2(n9254), .ZN(n9142) );
  NOR2_X1 U10249 ( .A1(n9142), .A2(n9513), .ZN(n8949) );
  AOI211_X1 U10250 ( .C1(n9140), .C2(n9068), .A(n8950), .B(n8949), .ZN(n8951)
         );
  OAI21_X1 U10251 ( .B1(n9143), .B2(n9114), .A(n8951), .ZN(P1_U3265) );
  XOR2_X1 U10252 ( .A(n8957), .B(n8952), .Z(n9148) );
  AOI21_X1 U10253 ( .B1(n9144), .B2(n8971), .A(n4584), .ZN(n9145) );
  AOI22_X1 U10254 ( .A1(n9513), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n8954), .B2(
        n9261), .ZN(n8955) );
  OAI21_X1 U10255 ( .B1(n8956), .B2(n9110), .A(n8955), .ZN(n8962) );
  XOR2_X1 U10256 ( .A(n8958), .B(n8957), .Z(n8960) );
  AOI222_X1 U10257 ( .A1(n9065), .A2(n8960), .B1(n8959), .B2(n9251), .C1(n4868), .C2(n9254), .ZN(n9147) );
  NOR2_X1 U10258 ( .A1(n9147), .A2(n9513), .ZN(n8961) );
  AOI211_X1 U10259 ( .C1(n9145), .C2(n9068), .A(n8962), .B(n8961), .ZN(n8963)
         );
  OAI21_X1 U10260 ( .B1(n9148), .B2(n9114), .A(n8963), .ZN(P1_U3266) );
  XOR2_X1 U10261 ( .A(n8967), .B(n8964), .Z(n9153) );
  AOI22_X1 U10262 ( .A1(n9150), .A2(n9262), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9513), .ZN(n8977) );
  AND2_X1 U10263 ( .A1(n8979), .A2(n8965), .ZN(n8968) );
  OAI21_X1 U10264 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(n8970) );
  AOI222_X1 U10265 ( .A1(n9065), .A2(n8970), .B1(n8969), .B2(n9251), .C1(n9000), .C2(n9254), .ZN(n9152) );
  INV_X1 U10266 ( .A(n8985), .ZN(n8972) );
  AOI211_X1 U10267 ( .C1(n9150), .C2(n8972), .A(n9548), .B(n4585), .ZN(n9149)
         );
  NAND2_X1 U10268 ( .A1(n9149), .A2(n5543), .ZN(n8973) );
  OAI211_X1 U10269 ( .C1(n9506), .C2(n8974), .A(n9152), .B(n8973), .ZN(n8975)
         );
  NAND2_X1 U10270 ( .A1(n8975), .A2(n5603), .ZN(n8976) );
  OAI211_X1 U10271 ( .C1(n9153), .C2(n9114), .A(n8977), .B(n8976), .ZN(
        P1_U3267) );
  XNOR2_X1 U10272 ( .A(n8978), .B(n8980), .ZN(n9158) );
  OAI211_X1 U10273 ( .C1(n8981), .C2(n8980), .A(n8979), .B(n9065), .ZN(n8983)
         );
  NAND2_X1 U10274 ( .A1(n4868), .A2(n9251), .ZN(n8982) );
  OAI211_X1 U10275 ( .C1(n8984), .C2(n5525), .A(n8983), .B(n8982), .ZN(n9154)
         );
  INV_X1 U10276 ( .A(n8994), .ZN(n8986) );
  AOI211_X1 U10277 ( .C1(n9156), .C2(n8986), .A(n9548), .B(n8985), .ZN(n9155)
         );
  NAND2_X1 U10278 ( .A1(n9155), .A2(n9269), .ZN(n8989) );
  AOI22_X1 U10279 ( .A1(n9513), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n8987), .B2(
        n9261), .ZN(n8988) );
  OAI211_X1 U10280 ( .C1(n8990), .C2(n9110), .A(n8989), .B(n8988), .ZN(n8991)
         );
  AOI21_X1 U10281 ( .B1(n9154), .B2(n5603), .A(n8991), .ZN(n8992) );
  OAI21_X1 U10282 ( .B1(n9158), .B2(n9114), .A(n8992), .ZN(P1_U3268) );
  XNOR2_X1 U10283 ( .A(n8993), .B(n8999), .ZN(n9163) );
  AOI21_X1 U10284 ( .B1(n9159), .B2(n9008), .A(n8994), .ZN(n9160) );
  AOI22_X1 U10285 ( .A1(n9513), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n8995), .B2(
        n9261), .ZN(n8996) );
  OAI21_X1 U10286 ( .B1(n8997), .B2(n9110), .A(n8996), .ZN(n9004) );
  XOR2_X1 U10287 ( .A(n8999), .B(n8998), .Z(n9002) );
  AOI222_X1 U10288 ( .A1(n9065), .A2(n9002), .B1(n9001), .B2(n9254), .C1(n9000), .C2(n9251), .ZN(n9162) );
  NOR2_X1 U10289 ( .A1(n9162), .A2(n9513), .ZN(n9003) );
  AOI211_X1 U10290 ( .C1(n9160), .C2(n9068), .A(n9004), .B(n9003), .ZN(n9005)
         );
  OAI21_X1 U10291 ( .B1(n9114), .B2(n9163), .A(n9005), .ZN(P1_U3269) );
  XNOR2_X1 U10292 ( .A(n9007), .B(n9006), .ZN(n9168) );
  INV_X1 U10293 ( .A(n9008), .ZN(n9009) );
  AOI211_X1 U10294 ( .C1(n9165), .C2(n9023), .A(n9548), .B(n9009), .ZN(n9164)
         );
  AOI22_X1 U10295 ( .A1(n9513), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9010), .B2(
        n9261), .ZN(n9011) );
  OAI21_X1 U10296 ( .B1(n9012), .B2(n9110), .A(n9011), .ZN(n9020) );
  AND2_X1 U10297 ( .A1(n9030), .A2(n9035), .ZN(n9015) );
  OAI21_X1 U10298 ( .B1(n9015), .B2(n9014), .A(n9013), .ZN(n9018) );
  AOI222_X1 U10299 ( .A1(n9065), .A2(n9018), .B1(n9017), .B2(n9251), .C1(n9016), .C2(n9254), .ZN(n9167) );
  NOR2_X1 U10300 ( .A1(n9167), .A2(n9513), .ZN(n9019) );
  AOI211_X1 U10301 ( .C1(n9269), .C2(n9164), .A(n9020), .B(n9019), .ZN(n9021)
         );
  OAI21_X1 U10302 ( .B1(n9114), .B2(n9168), .A(n9021), .ZN(P1_U3270) );
  XNOR2_X1 U10303 ( .A(n9022), .B(n9031), .ZN(n9173) );
  INV_X1 U10304 ( .A(n9047), .ZN(n9025) );
  INV_X1 U10305 ( .A(n9023), .ZN(n9024) );
  AOI21_X1 U10306 ( .B1(n9169), .B2(n9025), .A(n9024), .ZN(n9170) );
  AOI22_X1 U10307 ( .A1(n9513), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9026), .B2(
        n9261), .ZN(n9027) );
  OAI21_X1 U10308 ( .B1(n9028), .B2(n9110), .A(n9027), .ZN(n9040) );
  NOR2_X1 U10309 ( .A1(n9029), .A2(n9104), .ZN(n9038) );
  INV_X1 U10310 ( .A(n9030), .ZN(n9036) );
  INV_X1 U10311 ( .A(n9031), .ZN(n9032) );
  OAI21_X1 U10312 ( .B1(n9033), .B2(n9032), .A(n9065), .ZN(n9034) );
  AOI21_X1 U10313 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9037) );
  AOI211_X1 U10314 ( .C1(n9254), .C2(n9062), .A(n9038), .B(n9037), .ZN(n9172)
         );
  NOR2_X1 U10315 ( .A1(n9172), .A2(n9513), .ZN(n9039) );
  AOI211_X1 U10316 ( .C1(n9170), .C2(n9068), .A(n9040), .B(n9039), .ZN(n9041)
         );
  OAI21_X1 U10317 ( .B1(n9173), .B2(n9114), .A(n9041), .ZN(P1_U3271) );
  XNOR2_X1 U10318 ( .A(n9042), .B(n9044), .ZN(n9178) );
  XOR2_X1 U10319 ( .A(n9044), .B(n9043), .Z(n9045) );
  OAI222_X1 U10320 ( .A1(n5525), .A2(n9074), .B1(n9104), .B2(n9046), .C1(n9045), .C2(n9256), .ZN(n9174) );
  AOI211_X1 U10321 ( .C1(n9176), .C2(n4575), .A(n9548), .B(n9047), .ZN(n9175)
         );
  NAND2_X1 U10322 ( .A1(n9175), .A2(n9269), .ZN(n9050) );
  AOI22_X1 U10323 ( .A1(n9513), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9048), .B2(
        n9261), .ZN(n9049) );
  OAI211_X1 U10324 ( .C1(n9051), .C2(n9110), .A(n9050), .B(n9049), .ZN(n9052)
         );
  AOI21_X1 U10325 ( .B1(n9174), .B2(n9081), .A(n9052), .ZN(n9053) );
  OAI21_X1 U10326 ( .B1(n9178), .B2(n9114), .A(n9053), .ZN(P1_U3272) );
  XNOR2_X1 U10327 ( .A(n9055), .B(n9054), .ZN(n9183) );
  AOI21_X1 U10328 ( .B1(n9179), .B2(n4981), .A(n9056), .ZN(n9180) );
  AOI22_X1 U10329 ( .A1(n9513), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9057), .B2(
        n9261), .ZN(n9058) );
  OAI21_X1 U10330 ( .B1(n4573), .B2(n9110), .A(n9058), .ZN(n9067) );
  OAI21_X1 U10331 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9064) );
  AOI222_X1 U10332 ( .A1(n9065), .A2(n9064), .B1(n9063), .B2(n9254), .C1(n9062), .C2(n9251), .ZN(n9182) );
  NOR2_X1 U10333 ( .A1(n9182), .A2(n9513), .ZN(n9066) );
  AOI211_X1 U10334 ( .C1(n9180), .C2(n9068), .A(n9067), .B(n9066), .ZN(n9069)
         );
  OAI21_X1 U10335 ( .B1(n9114), .B2(n9183), .A(n9069), .ZN(P1_U3273) );
  XNOR2_X1 U10336 ( .A(n9070), .B(n9071), .ZN(n9188) );
  XNOR2_X1 U10337 ( .A(n9072), .B(n9071), .ZN(n9073) );
  OAI222_X1 U10338 ( .A1(n9104), .A2(n9074), .B1(n5525), .B2(n9103), .C1(n9073), .C2(n9256), .ZN(n9184) );
  INV_X1 U10339 ( .A(n4981), .ZN(n9075) );
  AOI211_X1 U10340 ( .C1(n9186), .C2(n9089), .A(n9548), .B(n9075), .ZN(n9185)
         );
  NAND2_X1 U10341 ( .A1(n9185), .A2(n9269), .ZN(n9078) );
  AOI22_X1 U10342 ( .A1(n9513), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9076), .B2(
        n9261), .ZN(n9077) );
  OAI211_X1 U10343 ( .C1(n9079), .C2(n9110), .A(n9078), .B(n9077), .ZN(n9080)
         );
  AOI21_X1 U10344 ( .B1(n9184), .B2(n9081), .A(n9080), .ZN(n9082) );
  OAI21_X1 U10345 ( .B1(n9188), .B2(n9114), .A(n9082), .ZN(P1_U3274) );
  XNOR2_X1 U10346 ( .A(n9083), .B(n9084), .ZN(n9193) );
  XNOR2_X1 U10347 ( .A(n9085), .B(n9084), .ZN(n9086) );
  OAI222_X1 U10348 ( .A1(n9104), .A2(n9088), .B1(n5525), .B2(n9087), .C1(n9086), .C2(n9256), .ZN(n9189) );
  INV_X1 U10349 ( .A(n9105), .ZN(n9091) );
  INV_X1 U10350 ( .A(n9089), .ZN(n9090) );
  AOI211_X1 U10351 ( .C1(n9191), .C2(n9091), .A(n9548), .B(n9090), .ZN(n9190)
         );
  NAND2_X1 U10352 ( .A1(n9190), .A2(n9269), .ZN(n9094) );
  AOI22_X1 U10353 ( .A1(n9513), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9092), .B2(
        n9261), .ZN(n9093) );
  OAI211_X1 U10354 ( .C1(n9095), .C2(n9110), .A(n9094), .B(n9093), .ZN(n9096)
         );
  AOI21_X1 U10355 ( .B1(n9189), .B2(n5603), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10356 ( .B1(n9193), .B2(n9114), .A(n9097), .ZN(P1_U3275) );
  XNOR2_X1 U10357 ( .A(n9098), .B(n9100), .ZN(n9199) );
  XOR2_X1 U10358 ( .A(n9100), .B(n9099), .Z(n9101) );
  OAI222_X1 U10359 ( .A1(n9104), .A2(n9103), .B1(n5525), .B2(n9102), .C1(n9256), .C2(n9101), .ZN(n9194) );
  AOI211_X1 U10360 ( .C1(n9196), .C2(n9106), .A(n9548), .B(n9105), .ZN(n9195)
         );
  NAND2_X1 U10361 ( .A1(n9195), .A2(n9269), .ZN(n9109) );
  AOI22_X1 U10362 ( .A1(n9513), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9107), .B2(
        n9261), .ZN(n9108) );
  OAI211_X1 U10363 ( .C1(n9111), .C2(n9110), .A(n9109), .B(n9108), .ZN(n9112)
         );
  AOI21_X1 U10364 ( .B1(n9194), .B2(n5603), .A(n9112), .ZN(n9113) );
  OAI21_X1 U10365 ( .B1(n9199), .B2(n9114), .A(n9113), .ZN(P1_U3276) );
  MUX2_X1 U10366 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9201), .S(n9565), .Z(
        P1_U3554) );
  NAND2_X1 U10367 ( .A1(n9120), .A2(n9537), .ZN(n9128) );
  INV_X1 U10368 ( .A(n9121), .ZN(n9125) );
  INV_X1 U10369 ( .A(n9123), .ZN(n9124) );
  OAI211_X1 U10370 ( .C1(n9548), .C2(n9125), .A(n4976), .B(n9124), .ZN(n9126)
         );
  INV_X1 U10371 ( .A(n9126), .ZN(n9127) );
  NAND2_X1 U10372 ( .A1(n9128), .A2(n9127), .ZN(n9202) );
  MUX2_X1 U10373 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9202), .S(n9565), .Z(
        P1_U3552) );
  AOI21_X1 U10374 ( .B1(n9529), .B2(n9130), .A(n9129), .ZN(n9131) );
  OAI211_X1 U10375 ( .C1(n9133), .C2(n9198), .A(n9132), .B(n9131), .ZN(n9203)
         );
  MUX2_X1 U10376 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9203), .S(n9565), .Z(
        P1_U3551) );
  AOI22_X1 U10377 ( .A1(n9135), .A2(n9530), .B1(n9529), .B2(n9134), .ZN(n9136)
         );
  OAI211_X1 U10378 ( .C1(n9138), .C2(n9198), .A(n9137), .B(n9136), .ZN(n9204)
         );
  MUX2_X1 U10379 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9204), .S(n9565), .Z(
        P1_U3550) );
  AOI22_X1 U10380 ( .A1(n9140), .A2(n9530), .B1(n9529), .B2(n9139), .ZN(n9141)
         );
  OAI211_X1 U10381 ( .C1(n9143), .C2(n9198), .A(n9142), .B(n9141), .ZN(n9205)
         );
  MUX2_X1 U10382 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9205), .S(n9565), .Z(
        P1_U3549) );
  AOI22_X1 U10383 ( .A1(n9145), .A2(n9530), .B1(n9529), .B2(n9144), .ZN(n9146)
         );
  OAI211_X1 U10384 ( .C1(n9148), .C2(n9198), .A(n9147), .B(n9146), .ZN(n9206)
         );
  MUX2_X1 U10385 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9206), .S(n9565), .Z(
        P1_U3548) );
  AOI21_X1 U10386 ( .B1(n9529), .B2(n9150), .A(n9149), .ZN(n9151) );
  OAI211_X1 U10387 ( .C1(n9153), .C2(n9198), .A(n9152), .B(n9151), .ZN(n9207)
         );
  MUX2_X1 U10388 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9207), .S(n9565), .Z(
        P1_U3547) );
  AOI211_X1 U10389 ( .C1(n9529), .C2(n9156), .A(n9155), .B(n9154), .ZN(n9157)
         );
  OAI21_X1 U10390 ( .B1(n9158), .B2(n9198), .A(n9157), .ZN(n9208) );
  MUX2_X1 U10391 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9208), .S(n9565), .Z(
        P1_U3546) );
  AOI22_X1 U10392 ( .A1(n9160), .A2(n9530), .B1(n9529), .B2(n9159), .ZN(n9161)
         );
  OAI211_X1 U10393 ( .C1(n9163), .C2(n9198), .A(n9162), .B(n9161), .ZN(n9209)
         );
  MUX2_X1 U10394 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9209), .S(n9565), .Z(
        P1_U3545) );
  AOI21_X1 U10395 ( .B1(n9529), .B2(n9165), .A(n9164), .ZN(n9166) );
  OAI211_X1 U10396 ( .C1(n9168), .C2(n9198), .A(n9167), .B(n9166), .ZN(n9210)
         );
  MUX2_X1 U10397 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9210), .S(n9565), .Z(
        P1_U3544) );
  AOI22_X1 U10398 ( .A1(n9170), .A2(n9530), .B1(n9529), .B2(n9169), .ZN(n9171)
         );
  OAI211_X1 U10399 ( .C1(n9173), .C2(n9198), .A(n9172), .B(n9171), .ZN(n9211)
         );
  MUX2_X1 U10400 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9211), .S(n9565), .Z(
        P1_U3543) );
  AOI211_X1 U10401 ( .C1(n9529), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9177)
         );
  OAI21_X1 U10402 ( .B1(n9178), .B2(n9198), .A(n9177), .ZN(n9212) );
  MUX2_X1 U10403 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9212), .S(n9565), .Z(
        P1_U3542) );
  AOI22_X1 U10404 ( .A1(n9180), .A2(n9530), .B1(n9529), .B2(n9179), .ZN(n9181)
         );
  OAI211_X1 U10405 ( .C1(n9183), .C2(n9198), .A(n9182), .B(n9181), .ZN(n9213)
         );
  MUX2_X1 U10406 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9213), .S(n9565), .Z(
        P1_U3541) );
  AOI211_X1 U10407 ( .C1(n9529), .C2(n9186), .A(n9185), .B(n9184), .ZN(n9187)
         );
  OAI21_X1 U10408 ( .B1(n9188), .B2(n9198), .A(n9187), .ZN(n9214) );
  MUX2_X1 U10409 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9214), .S(n9565), .Z(
        P1_U3540) );
  AOI211_X1 U10410 ( .C1(n9529), .C2(n9191), .A(n9190), .B(n9189), .ZN(n9192)
         );
  OAI21_X1 U10411 ( .B1(n9193), .B2(n9198), .A(n9192), .ZN(n9215) );
  MUX2_X1 U10412 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9215), .S(n9565), .Z(
        P1_U3539) );
  AOI211_X1 U10413 ( .C1(n9529), .C2(n9196), .A(n9195), .B(n9194), .ZN(n9197)
         );
  OAI21_X1 U10414 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9216) );
  MUX2_X1 U10415 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9216), .S(n9565), .Z(
        P1_U3538) );
  MUX2_X1 U10416 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9200), .S(n9565), .Z(
        P1_U3523) );
  MUX2_X1 U10417 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9201), .S(n9556), .Z(
        P1_U3522) );
  MUX2_X1 U10418 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9202), .S(n9556), .Z(
        P1_U3520) );
  MUX2_X1 U10419 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9203), .S(n9556), .Z(
        P1_U3519) );
  MUX2_X1 U10420 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9204), .S(n9556), .Z(
        P1_U3518) );
  MUX2_X1 U10421 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9205), .S(n9556), .Z(
        P1_U3517) );
  MUX2_X1 U10422 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9206), .S(n9556), .Z(
        P1_U3516) );
  MUX2_X1 U10423 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9207), .S(n9556), .Z(
        P1_U3515) );
  MUX2_X1 U10424 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9208), .S(n9556), .Z(
        P1_U3514) );
  MUX2_X1 U10425 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9209), .S(n9556), .Z(
        P1_U3513) );
  MUX2_X1 U10426 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9210), .S(n9556), .Z(
        P1_U3512) );
  MUX2_X1 U10427 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9211), .S(n9556), .Z(
        P1_U3511) );
  MUX2_X1 U10428 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9212), .S(n9556), .Z(
        P1_U3510) );
  MUX2_X1 U10429 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9213), .S(n9556), .Z(
        P1_U3508) );
  MUX2_X1 U10430 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9214), .S(n9556), .Z(
        P1_U3505) );
  MUX2_X1 U10431 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9215), .S(n9556), .Z(
        P1_U3502) );
  MUX2_X1 U10432 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9216), .S(n9556), .Z(
        P1_U3499) );
  MUX2_X1 U10433 ( .A(n9217), .B(P1_D_REG_0__SCAN_IN), .S(n9515), .Z(P1_U3440)
         );
  NOR4_X1 U10434 ( .A1(n9219), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9218), .ZN(n9220) );
  AOI21_X1 U10435 ( .B1(n9221), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9220), .ZN(
        n9222) );
  OAI21_X1 U10436 ( .B1(n9223), .B2(n4396), .A(n9222), .ZN(P1_U3322) );
  MUX2_X1 U10437 ( .A(n9224), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10438 ( .A1(n9600), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9235) );
  NAND2_X1 U10439 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9227) );
  AOI211_X1 U10440 ( .C1(n9227), .C2(n9226), .A(n9225), .B(n9596), .ZN(n9228)
         );
  AOI21_X1 U10441 ( .B1(n9241), .B2(n9229), .A(n9228), .ZN(n9234) );
  NOR2_X1 U10442 ( .A1(n9603), .A2(n9992), .ZN(n9232) );
  OAI211_X1 U10443 ( .C1(n9232), .C2(n9231), .A(n9598), .B(n9230), .ZN(n9233)
         );
  NAND3_X1 U10444 ( .A1(n9235), .A2(n9234), .A3(n9233), .ZN(P2_U3246) );
  AOI22_X1 U10445 ( .A1(n9600), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9247) );
  AOI211_X1 U10446 ( .C1(n9238), .C2(n9237), .A(n9236), .B(n9596), .ZN(n9239)
         );
  AOI21_X1 U10447 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9246) );
  OAI211_X1 U10448 ( .C1(n9244), .C2(n9243), .A(n9598), .B(n9242), .ZN(n9245)
         );
  NAND3_X1 U10449 ( .A1(n9247), .A2(n9246), .A3(n9245), .ZN(P2_U3247) );
  XNOR2_X1 U10450 ( .A(n9248), .B(n9249), .ZN(n9278) );
  XNOR2_X1 U10451 ( .A(n9250), .B(n9249), .ZN(n9257) );
  AOI22_X1 U10452 ( .A1(n9254), .A2(n9253), .B1(n9252), .B2(n9251), .ZN(n9255)
         );
  OAI21_X1 U10453 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9258) );
  AOI21_X1 U10454 ( .B1(n9278), .B2(n9259), .A(n9258), .ZN(n9275) );
  AOI222_X1 U10455 ( .A1(n9263), .A2(n9262), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9513), .C1(n9261), .C2(n9260), .ZN(n9272) );
  INV_X1 U10456 ( .A(n9264), .ZN(n9267) );
  INV_X1 U10457 ( .A(n9265), .ZN(n9266) );
  OAI211_X1 U10458 ( .C1(n9274), .C2(n9267), .A(n9266), .B(n9530), .ZN(n9273)
         );
  INV_X1 U10459 ( .A(n9273), .ZN(n9268) );
  AOI22_X1 U10460 ( .A1(n9278), .A2(n9270), .B1(n9269), .B2(n9268), .ZN(n9271)
         );
  OAI211_X1 U10461 ( .C1(n9513), .C2(n9275), .A(n9272), .B(n9271), .ZN(
        P1_U3281) );
  OAI21_X1 U10462 ( .B1(n9274), .B2(n9546), .A(n9273), .ZN(n9277) );
  INV_X1 U10463 ( .A(n9275), .ZN(n9276) );
  AOI211_X1 U10464 ( .C1(n9553), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9280)
         );
  INV_X1 U10465 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9279) );
  AOI22_X1 U10466 ( .A1(n9556), .A2(n9280), .B1(n9279), .B2(n9554), .ZN(
        P1_U3484) );
  AOI22_X1 U10467 ( .A1(n9565), .A2(n9280), .B1(n10080), .B2(n9563), .ZN(
        P1_U3533) );
  INV_X1 U10468 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10155) );
  NOR2_X1 U10469 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9281) );
  AOI21_X1 U10470 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9281), .ZN(n9811) );
  NOR2_X1 U10471 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9282) );
  AOI21_X1 U10472 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9282), .ZN(n9814) );
  NOR2_X1 U10473 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9283) );
  AOI21_X1 U10474 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9283), .ZN(n9817) );
  NOR2_X1 U10475 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9284) );
  AOI21_X1 U10476 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9284), .ZN(n9820) );
  NOR2_X1 U10477 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9285) );
  AOI21_X1 U10478 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9285), .ZN(n9823) );
  NOR2_X1 U10479 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9292) );
  XNOR2_X1 U10480 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10167) );
  NAND2_X1 U10481 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n9290) );
  XOR2_X1 U10482 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10165) );
  NAND2_X1 U10483 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9288) );
  XOR2_X1 U10484 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10163) );
  AOI21_X1 U10485 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9804) );
  INV_X1 U10486 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9286) );
  NAND3_X1 U10487 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9806) );
  OAI21_X1 U10488 ( .B1(n9804), .B2(n9286), .A(n9806), .ZN(n10162) );
  NAND2_X1 U10489 ( .A1(n10163), .A2(n10162), .ZN(n9287) );
  NAND2_X1 U10490 ( .A1(n9288), .A2(n9287), .ZN(n10164) );
  NAND2_X1 U10491 ( .A1(n10165), .A2(n10164), .ZN(n9289) );
  NAND2_X1 U10492 ( .A1(n9290), .A2(n9289), .ZN(n10166) );
  NOR2_X1 U10493 ( .A1(n10167), .A2(n10166), .ZN(n9291) );
  NOR2_X1 U10494 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  NOR2_X1 U10495 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9293), .ZN(n10150) );
  AND2_X1 U10496 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9293), .ZN(n10151) );
  NOR2_X1 U10497 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10151), .ZN(n9294) );
  NAND2_X1 U10498 ( .A1(n9295), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9297) );
  XOR2_X1 U10499 ( .A(n9295), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10149) );
  NAND2_X1 U10500 ( .A1(n10149), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U10501 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  NAND2_X1 U10502 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9298), .ZN(n9300) );
  XOR2_X1 U10503 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9298), .Z(n10161) );
  NAND2_X1 U10504 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10161), .ZN(n9299) );
  NAND2_X1 U10505 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  NAND2_X1 U10506 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9301), .ZN(n9303) );
  XOR2_X1 U10507 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9301), .Z(n10160) );
  NAND2_X1 U10508 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10160), .ZN(n9302) );
  NAND2_X1 U10509 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  AND2_X1 U10510 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9304), .ZN(n9305) );
  INV_X1 U10511 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10159) );
  XNOR2_X1 U10512 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9304), .ZN(n10158) );
  NAND2_X1 U10513 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9306) );
  OAI21_X1 U10514 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9306), .ZN(n9831) );
  NAND2_X1 U10515 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9307) );
  OAI21_X1 U10516 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9307), .ZN(n9828) );
  NOR2_X1 U10517 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9308) );
  AOI21_X1 U10518 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9308), .ZN(n9825) );
  NAND2_X1 U10519 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  OAI21_X1 U10520 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9824), .ZN(n9822) );
  NAND2_X1 U10521 ( .A1(n9823), .A2(n9822), .ZN(n9821) );
  OAI21_X1 U10522 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9821), .ZN(n9819) );
  NAND2_X1 U10523 ( .A1(n9820), .A2(n9819), .ZN(n9818) );
  OAI21_X1 U10524 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9818), .ZN(n9816) );
  NAND2_X1 U10525 ( .A1(n9817), .A2(n9816), .ZN(n9815) );
  OAI21_X1 U10526 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9815), .ZN(n9813) );
  NAND2_X1 U10527 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  OAI21_X1 U10528 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9812), .ZN(n9810) );
  NAND2_X1 U10529 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  OAI21_X1 U10530 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9809), .ZN(n10154) );
  NOR2_X1 U10531 ( .A1(n10155), .A2(n10154), .ZN(n9309) );
  NAND2_X1 U10532 ( .A1(n10155), .A2(n10154), .ZN(n10153) );
  OAI21_X1 U10533 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9309), .A(n10153), .ZN(
        n9311) );
  XOR2_X1 U10534 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n9310) );
  XNOR2_X1 U10535 ( .A(n9311), .B(n9310), .ZN(ADD_1071_U4) );
  OAI22_X1 U10536 ( .A1(n9313), .A2(n9778), .B1(n9312), .B2(n9776), .ZN(n9314)
         );
  AOI211_X1 U10537 ( .C1(n9316), .C2(n9783), .A(n9315), .B(n9314), .ZN(n9333)
         );
  AOI22_X1 U10538 ( .A1(n9803), .A2(n9333), .B1(n9317), .B2(n9801), .ZN(
        P2_U3535) );
  OAI22_X1 U10539 ( .A1(n9319), .A2(n9778), .B1(n9318), .B2(n9776), .ZN(n9320)
         );
  AOI211_X1 U10540 ( .C1(n9322), .C2(n9783), .A(n9321), .B(n9320), .ZN(n9335)
         );
  AOI22_X1 U10541 ( .A1(n9803), .A2(n9335), .B1(n9323), .B2(n9801), .ZN(
        P2_U3534) );
  INV_X1 U10542 ( .A(n9755), .ZN(n9715) );
  INV_X1 U10543 ( .A(n9324), .ZN(n9330) );
  INV_X1 U10544 ( .A(n9325), .ZN(n9326) );
  OAI22_X1 U10545 ( .A1(n9327), .A2(n9778), .B1(n9326), .B2(n9776), .ZN(n9329)
         );
  AOI211_X1 U10546 ( .C1(n9715), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9337)
         );
  AOI22_X1 U10547 ( .A1(n9803), .A2(n9337), .B1(n9331), .B2(n9801), .ZN(
        P2_U3533) );
  INV_X1 U10548 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9332) );
  AOI22_X1 U10549 ( .A1(n9785), .A2(n9333), .B1(n9332), .B2(n9784), .ZN(
        P2_U3496) );
  INV_X1 U10550 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9334) );
  AOI22_X1 U10551 ( .A1(n9785), .A2(n9335), .B1(n9334), .B2(n9784), .ZN(
        P2_U3493) );
  INV_X1 U10552 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9336) );
  AOI22_X1 U10553 ( .A1(n9785), .A2(n9337), .B1(n9336), .B2(n9784), .ZN(
        P2_U3490) );
  INV_X1 U10554 ( .A(n9338), .ZN(n9341) );
  NOR2_X1 U10555 ( .A1(n9339), .A2(n9548), .ZN(n9340) );
  INV_X1 U10556 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9343) );
  AOI22_X1 U10557 ( .A1(n9565), .A2(n9362), .B1(n9343), .B2(n9563), .ZN(
        P1_U3553) );
  OAI21_X1 U10558 ( .B1(n9345), .B2(n9546), .A(n9344), .ZN(n9346) );
  AOI211_X1 U10559 ( .C1(n9348), .C2(n9537), .A(n9347), .B(n9346), .ZN(n9363)
         );
  AOI22_X1 U10560 ( .A1(n9565), .A2(n9363), .B1(n9349), .B2(n9563), .ZN(
        P1_U3537) );
  OAI22_X1 U10561 ( .A1(n9351), .A2(n9548), .B1(n9350), .B2(n9546), .ZN(n9352)
         );
  AOI21_X1 U10562 ( .B1(n9353), .B2(n9553), .A(n9352), .ZN(n9354) );
  AND2_X1 U10563 ( .A1(n9355), .A2(n9354), .ZN(n9365) );
  AOI22_X1 U10564 ( .A1(n9565), .A2(n9365), .B1(n6469), .B2(n9563), .ZN(
        P1_U3536) );
  OAI21_X1 U10565 ( .B1(n9357), .B2(n9546), .A(n9356), .ZN(n9358) );
  AOI21_X1 U10566 ( .B1(n9359), .B2(n9553), .A(n9358), .ZN(n9360) );
  AND2_X1 U10567 ( .A1(n9361), .A2(n9360), .ZN(n9367) );
  AOI22_X1 U10568 ( .A1(n9565), .A2(n9367), .B1(n6177), .B2(n9563), .ZN(
        P1_U3535) );
  INV_X1 U10569 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U10570 ( .A1(n9556), .A2(n9362), .B1(n10091), .B2(n9554), .ZN(
        P1_U3521) );
  INV_X1 U10571 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U10572 ( .A1(n9556), .A2(n9363), .B1(n10106), .B2(n9554), .ZN(
        P1_U3496) );
  INV_X1 U10573 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9364) );
  AOI22_X1 U10574 ( .A1(n9556), .A2(n9365), .B1(n9364), .B2(n9554), .ZN(
        P1_U3493) );
  INV_X1 U10575 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9366) );
  AOI22_X1 U10576 ( .A1(n9556), .A2(n9367), .B1(n9366), .B2(n9554), .ZN(
        P1_U3490) );
  XNOR2_X1 U10577 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10578 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10579 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9375) );
  AND2_X1 U10580 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9396) );
  OAI22_X1 U10581 ( .A1(n9368), .A2(n9396), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9377), .ZN(n9372) );
  NOR2_X1 U10582 ( .A1(n9368), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9369) );
  OR2_X1 U10583 ( .A1(n5524), .A2(n9369), .ZN(n9371) );
  AOI21_X1 U10584 ( .B1(n9371), .B2(n9370), .A(P1_U3084), .ZN(n9400) );
  OAI211_X1 U10585 ( .C1(n5524), .C2(n9372), .A(n9400), .B(n5168), .ZN(n9373)
         );
  OAI22_X1 U10586 ( .A1(n9481), .A2(n9375), .B1(n9374), .B2(n9373), .ZN(n9376)
         );
  INV_X1 U10587 ( .A(n9376), .ZN(n9379) );
  NAND3_X1 U10588 ( .A1(n9496), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9377), .ZN(
        n9378) );
  OAI211_X1 U10589 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9380), .A(n9379), .B(
        n9378), .ZN(P1_U3241) );
  NAND2_X1 U10590 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9384) );
  AOI211_X1 U10591 ( .C1(n9384), .C2(n9383), .A(n9382), .B(n9381), .ZN(n9385)
         );
  AOI21_X1 U10592 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n9385), 
        .ZN(n9391) );
  AOI22_X1 U10593 ( .A1(n9495), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n9483), .B2(
        n9386), .ZN(n9390) );
  OAI211_X1 U10594 ( .C1(n9396), .C2(n9388), .A(n9477), .B(n9387), .ZN(n9389)
         );
  NAND3_X1 U10595 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(P1_U3242) );
  INV_X1 U10596 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9412) );
  OAI211_X1 U10597 ( .C1(n9394), .C2(n9393), .A(n9496), .B(n9392), .ZN(n9395)
         );
  INV_X1 U10598 ( .A(n9395), .ZN(n9410) );
  INV_X1 U10599 ( .A(n9396), .ZN(n9398) );
  MUX2_X1 U10600 ( .A(n9399), .B(n9398), .S(n9397), .Z(n9402) );
  OAI211_X1 U10601 ( .C1(n9402), .C2(n5524), .A(n9401), .B(n9400), .ZN(n9429)
         );
  XOR2_X1 U10602 ( .A(n9404), .B(n9403), .Z(n9405) );
  NAND2_X1 U10603 ( .A1(n9477), .A2(n9405), .ZN(n9406) );
  OAI211_X1 U10604 ( .C1(n9408), .C2(n9407), .A(n9429), .B(n9406), .ZN(n9409)
         );
  AOI211_X1 U10605 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n9410), 
        .B(n9409), .ZN(n9411) );
  OAI21_X1 U10606 ( .B1(n9481), .B2(n9412), .A(n9411), .ZN(P1_U3243) );
  INV_X1 U10607 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U10608 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  AND2_X1 U10609 ( .A1(n9416), .A2(n9415), .ZN(n9427) );
  INV_X1 U10610 ( .A(n9417), .ZN(n9418) );
  NAND2_X1 U10611 ( .A1(n9483), .A2(n9418), .ZN(n9426) );
  NAND2_X1 U10612 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  NAND2_X1 U10613 ( .A1(n9422), .A2(n9421), .ZN(n9424) );
  AOI21_X1 U10614 ( .B1(n9496), .B2(n9424), .A(n9423), .ZN(n9425) );
  OAI211_X1 U10615 ( .C1(n9488), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9428)
         );
  INV_X1 U10616 ( .A(n9428), .ZN(n9430) );
  OAI211_X1 U10617 ( .C1(n9431), .C2(n9481), .A(n9430), .B(n9429), .ZN(
        P1_U3245) );
  OAI21_X1 U10618 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9440) );
  AOI211_X1 U10619 ( .C1(n9437), .C2(n9436), .A(n9435), .B(n9488), .ZN(n9438)
         );
  AOI211_X1 U10620 ( .C1(n9496), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9443)
         );
  AOI22_X1 U10621 ( .A1(n9495), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9483), .B2(
        n9441), .ZN(n9442) );
  NAND2_X1 U10622 ( .A1(n9443), .A2(n9442), .ZN(P1_U3250) );
  AOI22_X1 U10623 ( .A1(n9495), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9483), .B2(
        n9444), .ZN(n9455) );
  OAI21_X1 U10624 ( .B1(n9447), .B2(n9446), .A(n9445), .ZN(n9453) );
  AOI211_X1 U10625 ( .C1(n9450), .C2(n9449), .A(n9448), .B(n9488), .ZN(n9451)
         );
  AOI211_X1 U10626 ( .C1(n9496), .C2(n9453), .A(n9452), .B(n9451), .ZN(n9454)
         );
  NAND2_X1 U10627 ( .A1(n9455), .A2(n9454), .ZN(P1_U3251) );
  INV_X1 U10628 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9467) );
  AOI21_X1 U10629 ( .B1(n9483), .B2(n9457), .A(n9456), .ZN(n9466) );
  OAI21_X1 U10630 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9464) );
  XNOR2_X1 U10631 ( .A(n9462), .B(n9461), .ZN(n9463) );
  AOI22_X1 U10632 ( .A1(n9464), .A2(n9496), .B1(n9477), .B2(n9463), .ZN(n9465)
         );
  OAI211_X1 U10633 ( .C1(n9481), .C2(n9467), .A(n9466), .B(n9465), .ZN(
        P1_U3252) );
  INV_X1 U10634 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9923) );
  AOI21_X1 U10635 ( .B1(n9483), .B2(n9469), .A(n9468), .ZN(n9480) );
  OAI21_X1 U10636 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9478) );
  OAI21_X1 U10637 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9476) );
  AOI22_X1 U10638 ( .A1(n9478), .A2(n9477), .B1(n9496), .B2(n9476), .ZN(n9479)
         );
  OAI211_X1 U10639 ( .C1(n9481), .C2(n9923), .A(n9480), .B(n9479), .ZN(
        P1_U3255) );
  NAND2_X1 U10640 ( .A1(n9483), .A2(n9482), .ZN(n9491) );
  AND2_X1 U10641 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  OR3_X1 U10642 ( .A1(n9488), .A2(n9487), .A3(n9486), .ZN(n9490) );
  AND3_X1 U10643 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n9499) );
  OAI21_X1 U10644 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9497) );
  AOI22_X1 U10645 ( .A1(n9497), .A2(n9496), .B1(n9495), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U10646 ( .A1(n9499), .A2(n9498), .ZN(P1_U3259) );
  INV_X1 U10647 ( .A(n9500), .ZN(n9503) );
  NOR2_X1 U10648 ( .A1(n9501), .A2(n5611), .ZN(n9502) );
  MUX2_X1 U10649 ( .A(n9503), .B(n9502), .S(n5403), .Z(n9511) );
  INV_X1 U10650 ( .A(n9504), .ZN(n9508) );
  OAI22_X1 U10651 ( .A1(n9508), .A2(n9507), .B1(n9506), .B2(n9505), .ZN(n9509)
         );
  NOR3_X1 U10652 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(n9512) );
  AOI22_X1 U10653 ( .A1(n9513), .A2(n5993), .B1(n9512), .B2(n5603), .ZN(
        P1_U3290) );
  AND2_X1 U10654 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9515), .ZN(P1_U3292) );
  INV_X1 U10655 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U10656 ( .A1(n9514), .A2(n10064), .ZN(P1_U3293) );
  AND2_X1 U10657 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9515), .ZN(P1_U3294) );
  AND2_X1 U10658 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9515), .ZN(P1_U3295) );
  AND2_X1 U10659 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9515), .ZN(P1_U3296) );
  INV_X1 U10660 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U10661 ( .A1(n9514), .A2(n10105), .ZN(P1_U3297) );
  INV_X1 U10662 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U10663 ( .A1(n9514), .A2(n10119), .ZN(P1_U3298) );
  AND2_X1 U10664 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9515), .ZN(P1_U3299) );
  INV_X1 U10665 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U10666 ( .A1(n9514), .A2(n9945), .ZN(P1_U3300) );
  AND2_X1 U10667 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9515), .ZN(P1_U3301) );
  AND2_X1 U10668 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9515), .ZN(P1_U3302) );
  AND2_X1 U10669 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9515), .ZN(P1_U3303) );
  AND2_X1 U10670 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9515), .ZN(P1_U3304) );
  INV_X1 U10671 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U10672 ( .A1(n9514), .A2(n10055), .ZN(P1_U3305) );
  INV_X1 U10673 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U10674 ( .A1(n9514), .A2(n9916), .ZN(P1_U3306) );
  INV_X1 U10675 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U10676 ( .A1(n9514), .A2(n9932), .ZN(P1_U3307) );
  AND2_X1 U10677 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9515), .ZN(P1_U3308) );
  INV_X1 U10678 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U10679 ( .A1(n9514), .A2(n9966), .ZN(P1_U3309) );
  INV_X1 U10680 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10681 ( .A1(n9514), .A2(n10049), .ZN(P1_U3310) );
  INV_X1 U10682 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U10683 ( .A1(n9514), .A2(n10128), .ZN(P1_U3311) );
  INV_X1 U10684 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U10685 ( .A1(n9514), .A2(n9935), .ZN(P1_U3312) );
  AND2_X1 U10686 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9515), .ZN(P1_U3313) );
  AND2_X1 U10687 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9515), .ZN(P1_U3314) );
  AND2_X1 U10688 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9515), .ZN(P1_U3315) );
  AND2_X1 U10689 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9515), .ZN(P1_U3316) );
  AND2_X1 U10690 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9515), .ZN(P1_U3317) );
  AND2_X1 U10691 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9515), .ZN(P1_U3318) );
  INV_X1 U10692 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U10693 ( .A1(n9514), .A2(n10046), .ZN(P1_U3319) );
  AND2_X1 U10694 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9515), .ZN(P1_U3320) );
  AND2_X1 U10695 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9515), .ZN(P1_U3321) );
  INV_X1 U10696 ( .A(n9516), .ZN(n9521) );
  OAI22_X1 U10697 ( .A1(n9518), .A2(n9548), .B1(n9517), .B2(n9546), .ZN(n9520)
         );
  AOI211_X1 U10698 ( .C1(n9553), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9558)
         );
  INV_X1 U10699 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9522) );
  AOI22_X1 U10700 ( .A1(n9556), .A2(n9558), .B1(n9522), .B2(n9554), .ZN(
        P1_U3460) );
  OAI21_X1 U10701 ( .B1(n9524), .B2(n9546), .A(n9523), .ZN(n9526) );
  AOI211_X1 U10702 ( .C1(n9553), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9560)
         );
  INV_X1 U10703 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9528) );
  AOI22_X1 U10704 ( .A1(n9556), .A2(n9560), .B1(n9528), .B2(n9554), .ZN(
        P1_U3466) );
  AOI22_X1 U10705 ( .A1(n9531), .A2(n9530), .B1(n9529), .B2(n5527), .ZN(n9532)
         );
  OAI211_X1 U10706 ( .C1(n9535), .C2(n9534), .A(n9533), .B(n9532), .ZN(n9536)
         );
  INV_X1 U10707 ( .A(n9536), .ZN(n9561) );
  INV_X1 U10708 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U10709 ( .A1(n9556), .A2(n9561), .B1(n10067), .B2(n9554), .ZN(
        P1_U3472) );
  NAND2_X1 U10710 ( .A1(n9538), .A2(n9537), .ZN(n9544) );
  OAI22_X1 U10711 ( .A1(n9540), .A2(n9548), .B1(n9539), .B2(n9546), .ZN(n9541)
         );
  NOR2_X1 U10712 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  INV_X1 U10713 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9545) );
  AOI22_X1 U10714 ( .A1(n9556), .A2(n9562), .B1(n9545), .B2(n9554), .ZN(
        P1_U3478) );
  OAI22_X1 U10715 ( .A1(n9549), .A2(n9548), .B1(n9547), .B2(n9546), .ZN(n9551)
         );
  AOI211_X1 U10716 ( .C1(n9553), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9564)
         );
  INV_X1 U10717 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U10718 ( .A1(n9556), .A2(n9564), .B1(n9555), .B2(n9554), .ZN(
        P1_U3481) );
  INV_X1 U10719 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10720 ( .A1(n9565), .A2(n9558), .B1(n9557), .B2(n9563), .ZN(
        P1_U3525) );
  AOI22_X1 U10721 ( .A1(n9565), .A2(n9560), .B1(n9559), .B2(n9563), .ZN(
        P1_U3527) );
  AOI22_X1 U10722 ( .A1(n9565), .A2(n9561), .B1(n6031), .B2(n9563), .ZN(
        P1_U3529) );
  AOI22_X1 U10723 ( .A1(n9565), .A2(n9562), .B1(n6056), .B2(n9563), .ZN(
        P1_U3531) );
  INV_X1 U10724 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U10725 ( .A1(n9565), .A2(n9564), .B1(n10035), .B2(n9563), .ZN(
        P1_U3532) );
  OAI21_X1 U10726 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9576) );
  AOI21_X1 U10727 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9572) );
  OAI21_X1 U10728 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9575) );
  AOI21_X1 U10729 ( .B1(n9576), .B2(n9589), .A(n9575), .ZN(n9577) );
  OAI21_X1 U10730 ( .B1(n9593), .B2(n9578), .A(n9577), .ZN(P2_U3233) );
  OAI21_X1 U10731 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9590) );
  AOI21_X1 U10732 ( .B1(n9584), .B2(n9583), .A(n9582), .ZN(n9585) );
  OAI21_X1 U10733 ( .B1(n9587), .B2(n9586), .A(n9585), .ZN(n9588) );
  AOI21_X1 U10734 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9591) );
  OAI21_X1 U10735 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(P2_U3241) );
  AOI22_X1 U10736 ( .A1(n9598), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9594), .ZN(n9604) );
  OAI21_X1 U10737 ( .B1(n9596), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9595), .ZN(
        n9597) );
  AOI21_X1 U10738 ( .B1(n9598), .B2(n9992), .A(n9597), .ZN(n9602) );
  AOI22_X1 U10739 ( .A1(n9600), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9601) );
  OAI221_X1 U10740 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9604), .C1(n9603), .C2(
        n9602), .A(n9601), .ZN(P2_U3245) );
  XOR2_X1 U10741 ( .A(n9605), .B(n9607), .Z(n9728) );
  AOI22_X1 U10742 ( .A1(n9728), .A2(n9638), .B1(P2_REG2_REG_5__SCAN_IN), .B2(
        n9669), .ZN(n9621) );
  NAND2_X1 U10743 ( .A1(n9626), .A2(n9606), .ZN(n9608) );
  XNOR2_X1 U10744 ( .A(n9608), .B(n9607), .ZN(n9609) );
  OAI222_X1 U10745 ( .A1(n9613), .A2(n9612), .B1(n9611), .B2(n9610), .C1(n9644), .C2(n9609), .ZN(n9726) );
  OAI21_X1 U10746 ( .B1(n9651), .B2(n9630), .A(n4395), .ZN(n9616) );
  NAND3_X1 U10747 ( .A1(n9616), .A2(n9752), .A3(n9615), .ZN(n9724) );
  OAI22_X1 U10748 ( .A1(n9724), .A2(n6138), .B1(n9725), .B2(n9617), .ZN(n9619)
         );
  OAI21_X1 U10749 ( .B1(n9726), .B2(n9619), .A(n9618), .ZN(n9620) );
  OAI211_X1 U10750 ( .C1(n9666), .C2(n9622), .A(n9621), .B(n9620), .ZN(
        P2_U3291) );
  INV_X1 U10751 ( .A(n9623), .ZN(n9624) );
  AOI21_X1 U10752 ( .B1(n9624), .B2(n9629), .A(n9644), .ZN(n9627) );
  AOI21_X1 U10753 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9719) );
  XNOR2_X1 U10754 ( .A(n9629), .B(n9628), .ZN(n9722) );
  XNOR2_X1 U10755 ( .A(n9651), .B(n9630), .ZN(n9718) );
  NAND2_X1 U10756 ( .A1(n9631), .A2(n9630), .ZN(n9635) );
  AOI22_X1 U10757 ( .A1(n9669), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n9633), .B2(
        n9632), .ZN(n9634) );
  OAI211_X1 U10758 ( .C1(n9718), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9637)
         );
  AOI21_X1 U10759 ( .B1(n9638), .B2(n9722), .A(n9637), .ZN(n9639) );
  OAI21_X1 U10760 ( .B1(n9669), .B2(n9719), .A(n9639), .ZN(P2_U3292) );
  INV_X1 U10761 ( .A(n9640), .ZN(n9761) );
  XNOR2_X1 U10762 ( .A(n9643), .B(n9641), .ZN(n9714) );
  XNOR2_X1 U10763 ( .A(n9643), .B(n9642), .ZN(n9645) );
  NOR2_X1 U10764 ( .A1(n9645), .A2(n9644), .ZN(n9646) );
  AOI211_X1 U10765 ( .C1(n9761), .C2(n9714), .A(n9647), .B(n9646), .ZN(n9711)
         );
  INV_X1 U10766 ( .A(n9648), .ZN(n9649) );
  NAND2_X1 U10767 ( .A1(n9714), .A2(n9649), .ZN(n9657) );
  OR2_X1 U10768 ( .A1(n9665), .A2(n9709), .ZN(n9650) );
  NAND2_X1 U10769 ( .A1(n9651), .A2(n9650), .ZN(n9710) );
  INV_X1 U10770 ( .A(n9710), .ZN(n9652) );
  NAND2_X1 U10771 ( .A1(n9668), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U10772 ( .A1(n9669), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9653) );
  OAI211_X1 U10773 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9666), .A(n9654), .B(
        n9653), .ZN(n9655) );
  INV_X1 U10774 ( .A(n9655), .ZN(n9656) );
  OAI211_X1 U10775 ( .C1(n9709), .C2(n9673), .A(n9657), .B(n9656), .ZN(n9658)
         );
  INV_X1 U10776 ( .A(n9658), .ZN(n9659) );
  OAI21_X1 U10777 ( .B1(n9669), .B2(n9711), .A(n9659), .ZN(P2_U3293) );
  XNOR2_X1 U10778 ( .A(n9675), .B(n9660), .ZN(n9663) );
  AOI21_X1 U10779 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9706) );
  AND2_X1 U10780 ( .A1(n9696), .A2(n9703), .ZN(n9664) );
  NOR2_X1 U10781 ( .A1(n9665), .A2(n9664), .ZN(n9704) );
  INV_X1 U10782 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U10783 ( .A1(n9666), .A2(n10096), .ZN(n9667) );
  AOI21_X1 U10784 ( .B1(n9668), .B2(n9704), .A(n9667), .ZN(n9671) );
  NAND2_X1 U10785 ( .A1(n9669), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9670) );
  OAI211_X1 U10786 ( .C1(n9673), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9678)
         );
  XNOR2_X1 U10787 ( .A(n9674), .B(n4888), .ZN(n9707) );
  NOR2_X1 U10788 ( .A1(n9676), .A2(n9707), .ZN(n9677) );
  NOR2_X1 U10789 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  OAI21_X1 U10790 ( .B1(n9669), .B2(n9706), .A(n9679), .ZN(P2_U3294) );
  INV_X1 U10791 ( .A(n9680), .ZN(n9682) );
  INV_X1 U10792 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U10793 ( .A1(n9685), .A2(n9929), .ZN(P2_U3297) );
  AND2_X1 U10794 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9687), .ZN(P2_U3298) );
  AND2_X1 U10795 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9687), .ZN(P2_U3299) );
  AND2_X1 U10796 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9687), .ZN(P2_U3300) );
  AND2_X1 U10797 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9687), .ZN(P2_U3301) );
  INV_X1 U10798 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U10799 ( .A1(n9685), .A2(n9919), .ZN(P2_U3302) );
  AND2_X1 U10800 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9687), .ZN(P2_U3303) );
  AND2_X1 U10801 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9687), .ZN(P2_U3304) );
  AND2_X1 U10802 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9687), .ZN(P2_U3305) );
  INV_X1 U10803 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U10804 ( .A1(n9685), .A2(n10063), .ZN(P2_U3306) );
  AND2_X1 U10805 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9687), .ZN(P2_U3307) );
  AND2_X1 U10806 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9687), .ZN(P2_U3308) );
  AND2_X1 U10807 ( .A1(n9687), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3309) );
  AND2_X1 U10808 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9687), .ZN(P2_U3310) );
  AND2_X1 U10809 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9687), .ZN(P2_U3311) );
  AND2_X1 U10810 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9687), .ZN(P2_U3312) );
  AND2_X1 U10811 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9687), .ZN(P2_U3313) );
  AND2_X1 U10812 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9687), .ZN(P2_U3314) );
  AND2_X1 U10813 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9687), .ZN(P2_U3315) );
  AND2_X1 U10814 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9687), .ZN(P2_U3316) );
  AND2_X1 U10815 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9687), .ZN(P2_U3317) );
  AND2_X1 U10816 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9687), .ZN(P2_U3318) );
  INV_X1 U10817 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U10818 ( .A1(n9685), .A2(n9974), .ZN(P2_U3319) );
  INV_X1 U10819 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U10820 ( .A1(n9685), .A2(n10112), .ZN(P2_U3320) );
  AND2_X1 U10821 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9687), .ZN(P2_U3321) );
  AND2_X1 U10822 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9687), .ZN(P2_U3322) );
  AND2_X1 U10823 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9687), .ZN(P2_U3323) );
  AND2_X1 U10824 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9687), .ZN(P2_U3324) );
  AND2_X1 U10825 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9687), .ZN(P2_U3325) );
  AND2_X1 U10826 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9687), .ZN(P2_U3326) );
  OAI22_X1 U10827 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9685), .B1(n9684), .B2(
        n9683), .ZN(n9686) );
  INV_X1 U10828 ( .A(n9686), .ZN(P2_U3437) );
  AOI22_X1 U10829 ( .A1(n9690), .A2(n9689), .B1(n9688), .B2(n9687), .ZN(
        P2_U3438) );
  OAI22_X1 U10830 ( .A1(n9692), .A2(n9740), .B1(n6752), .B2(n9691), .ZN(n9693)
         );
  NOR2_X1 U10831 ( .A1(n9694), .A2(n9693), .ZN(n9786) );
  INV_X1 U10832 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10833 ( .A1(n9785), .A2(n9786), .B1(n9695), .B2(n9784), .ZN(
        P2_U3451) );
  NAND3_X1 U10834 ( .A1(n9697), .A2(n9752), .A3(n9696), .ZN(n9698) );
  OAI21_X1 U10835 ( .B1(n9776), .B2(n9699), .A(n9698), .ZN(n9701) );
  AOI211_X1 U10836 ( .C1(n9702), .C2(n9783), .A(n9701), .B(n9700), .ZN(n9787)
         );
  INV_X1 U10837 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U10838 ( .A1(n9785), .A2(n9787), .B1(n10129), .B2(n9784), .ZN(
        P2_U3454) );
  AOI22_X1 U10839 ( .A1(n9704), .A2(n9752), .B1(n9751), .B2(n9703), .ZN(n9705)
         );
  OAI211_X1 U10840 ( .C1(n9740), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9708)
         );
  INV_X1 U10841 ( .A(n9708), .ZN(n9789) );
  INV_X1 U10842 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U10843 ( .A1(n9785), .A2(n9789), .B1(n10113), .B2(n9784), .ZN(
        P2_U3457) );
  OAI22_X1 U10844 ( .A1(n9710), .A2(n9778), .B1(n9709), .B2(n9776), .ZN(n9713)
         );
  INV_X1 U10845 ( .A(n9711), .ZN(n9712) );
  AOI211_X1 U10846 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9790)
         );
  INV_X1 U10847 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U10848 ( .A1(n9785), .A2(n9790), .B1(n9716), .B2(n9784), .ZN(
        P2_U3460) );
  OAI22_X1 U10849 ( .A1(n9718), .A2(n9778), .B1(n9717), .B2(n9776), .ZN(n9721)
         );
  INV_X1 U10850 ( .A(n9719), .ZN(n9720) );
  AOI211_X1 U10851 ( .C1(n9783), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9791)
         );
  INV_X1 U10852 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9723) );
  AOI22_X1 U10853 ( .A1(n9785), .A2(n9791), .B1(n9723), .B2(n9784), .ZN(
        P2_U3463) );
  OAI21_X1 U10854 ( .B1(n9725), .B2(n9776), .A(n9724), .ZN(n9727) );
  AOI211_X1 U10855 ( .C1(n9783), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9793)
         );
  INV_X1 U10856 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U10857 ( .A1(n9785), .A2(n9793), .B1(n9918), .B2(n9784), .ZN(
        P2_U3466) );
  INV_X1 U10858 ( .A(n9729), .ZN(n9735) );
  OAI22_X1 U10859 ( .A1(n9731), .A2(n9778), .B1(n9730), .B2(n9776), .ZN(n9734)
         );
  INV_X1 U10860 ( .A(n9732), .ZN(n9733) );
  AOI211_X1 U10861 ( .C1(n9783), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9795)
         );
  INV_X1 U10862 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U10863 ( .A1(n9785), .A2(n9795), .B1(n10061), .B2(n9784), .ZN(
        P2_U3469) );
  AOI22_X1 U10864 ( .A1(n9737), .A2(n9752), .B1(n9751), .B2(n9736), .ZN(n9738)
         );
  OAI211_X1 U10865 ( .C1(n9741), .C2(n9740), .A(n9739), .B(n9738), .ZN(n9742)
         );
  INV_X1 U10866 ( .A(n9742), .ZN(n9796) );
  INV_X1 U10867 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U10868 ( .A1(n9785), .A2(n9796), .B1(n9743), .B2(n9784), .ZN(
        P2_U3472) );
  OAI22_X1 U10869 ( .A1(n9745), .A2(n9778), .B1(n9744), .B2(n9776), .ZN(n9747)
         );
  AOI211_X1 U10870 ( .C1(n9748), .C2(n9783), .A(n9747), .B(n9746), .ZN(n9797)
         );
  INV_X1 U10871 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9749) );
  AOI22_X1 U10872 ( .A1(n9785), .A2(n9797), .B1(n9749), .B2(n9784), .ZN(
        P2_U3475) );
  AOI22_X1 U10873 ( .A1(n9753), .A2(n9752), .B1(n9751), .B2(n9750), .ZN(n9754)
         );
  OAI21_X1 U10874 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9759) );
  INV_X1 U10875 ( .A(n9757), .ZN(n9758) );
  AOI211_X1 U10876 ( .C1(n9761), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9798)
         );
  INV_X1 U10877 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9762) );
  AOI22_X1 U10878 ( .A1(n9785), .A2(n9798), .B1(n9762), .B2(n9784), .ZN(
        P2_U3478) );
  OAI22_X1 U10879 ( .A1(n9764), .A2(n9778), .B1(n9763), .B2(n9776), .ZN(n9766)
         );
  AOI211_X1 U10880 ( .C1(n9783), .C2(n9767), .A(n9766), .B(n9765), .ZN(n9799)
         );
  INV_X1 U10881 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10882 ( .A1(n9785), .A2(n9799), .B1(n9768), .B2(n9784), .ZN(
        P2_U3481) );
  INV_X1 U10883 ( .A(n9769), .ZN(n9774) );
  OAI22_X1 U10884 ( .A1(n9771), .A2(n9778), .B1(n9770), .B2(n9776), .ZN(n9773)
         );
  AOI211_X1 U10885 ( .C1(n9774), .C2(n9783), .A(n9773), .B(n9772), .ZN(n9800)
         );
  INV_X1 U10886 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9775) );
  AOI22_X1 U10887 ( .A1(n9785), .A2(n9800), .B1(n9775), .B2(n9784), .ZN(
        P2_U3484) );
  OAI22_X1 U10888 ( .A1(n9779), .A2(n9778), .B1(n9777), .B2(n9776), .ZN(n9781)
         );
  AOI211_X1 U10889 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9802)
         );
  INV_X1 U10890 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U10891 ( .A1(n9785), .A2(n9802), .B1(n9949), .B2(n9784), .ZN(
        P2_U3487) );
  AOI22_X1 U10892 ( .A1(n9803), .A2(n9786), .B1(n10093), .B2(n9801), .ZN(
        P2_U3520) );
  AOI22_X1 U10893 ( .A1(n9803), .A2(n9787), .B1(n6071), .B2(n9801), .ZN(
        P2_U3521) );
  INV_X1 U10894 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U10895 ( .A1(n9803), .A2(n9789), .B1(n9788), .B2(n9801), .ZN(
        P2_U3522) );
  AOI22_X1 U10896 ( .A1(n9803), .A2(n9790), .B1(n6144), .B2(n9801), .ZN(
        P2_U3523) );
  AOI22_X1 U10897 ( .A1(n9803), .A2(n9791), .B1(n6233), .B2(n9801), .ZN(
        P2_U3524) );
  INV_X1 U10898 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9792) );
  AOI22_X1 U10899 ( .A1(n9803), .A2(n9793), .B1(n9792), .B2(n9801), .ZN(
        P2_U3525) );
  INV_X1 U10900 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U10901 ( .A1(n9803), .A2(n9795), .B1(n9794), .B2(n9801), .ZN(
        P2_U3526) );
  AOI22_X1 U10902 ( .A1(n9803), .A2(n9796), .B1(n6271), .B2(n9801), .ZN(
        P2_U3527) );
  AOI22_X1 U10903 ( .A1(n9803), .A2(n9797), .B1(n6272), .B2(n9801), .ZN(
        P2_U3528) );
  AOI22_X1 U10904 ( .A1(n9803), .A2(n9798), .B1(n6391), .B2(n9801), .ZN(
        P2_U3529) );
  AOI22_X1 U10905 ( .A1(n9803), .A2(n9799), .B1(n6392), .B2(n9801), .ZN(
        P2_U3530) );
  AOI22_X1 U10906 ( .A1(n9803), .A2(n9800), .B1(n6393), .B2(n9801), .ZN(
        P2_U3531) );
  AOI22_X1 U10907 ( .A1(n9803), .A2(n9802), .B1(n6489), .B2(n9801), .ZN(
        P2_U3532) );
  INV_X1 U10908 ( .A(n9804), .ZN(n9805) );
  NAND2_X1 U10909 ( .A1(n9806), .A2(n9805), .ZN(n9807) );
  XNOR2_X1 U10910 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9807), .ZN(ADD_1071_U5) );
  INV_X1 U10911 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10912 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9808), .B2(n9375), .ZN(ADD_1071_U46) );
  OAI21_X1 U10913 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(ADD_1071_U56) );
  OAI21_X1 U10914 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(ADD_1071_U57) );
  OAI21_X1 U10915 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(ADD_1071_U58) );
  OAI21_X1 U10916 ( .B1(n9820), .B2(n9819), .A(n9818), .ZN(ADD_1071_U59) );
  OAI21_X1 U10917 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(ADD_1071_U60) );
  OAI21_X1 U10918 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(ADD_1071_U61) );
  AOI21_X1 U10919 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(ADD_1071_U62) );
  AOI21_X1 U10920 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(ADD_1071_U63) );
  NAND2_X1 U10921 ( .A1(keyinput15), .A2(keyinput121), .ZN(n9833) );
  NOR3_X1 U10922 ( .A1(keyinput32), .A2(keyinput91), .A3(n9833), .ZN(n9835) );
  INV_X1 U10923 ( .A(keyinput48), .ZN(n9834) );
  NAND4_X1 U10924 ( .A1(keyinput111), .A2(keyinput96), .A3(n9835), .A4(n9834), 
        .ZN(n9847) );
  NOR3_X1 U10925 ( .A1(keyinput79), .A2(keyinput75), .A3(keyinput101), .ZN(
        n9836) );
  NAND2_X1 U10926 ( .A1(keyinput36), .A2(n9836), .ZN(n9846) );
  NAND4_X1 U10927 ( .A1(keyinput122), .A2(keyinput17), .A3(keyinput12), .A4(
        keyinput31), .ZN(n9845) );
  NOR4_X1 U10928 ( .A1(keyinput118), .A2(keyinput7), .A3(keyinput16), .A4(
        keyinput63), .ZN(n9843) );
  NAND3_X1 U10929 ( .A1(keyinput97), .A2(keyinput93), .A3(keyinput20), .ZN(
        n9837) );
  NOR2_X1 U10930 ( .A1(keyinput109), .A2(n9837), .ZN(n9842) );
  INV_X1 U10931 ( .A(keyinput103), .ZN(n9838) );
  NOR4_X1 U10932 ( .A1(keyinput62), .A2(keyinput127), .A3(keyinput43), .A4(
        n9838), .ZN(n9841) );
  NAND2_X1 U10933 ( .A1(keyinput11), .A2(keyinput124), .ZN(n9839) );
  NOR3_X1 U10934 ( .A1(keyinput52), .A2(keyinput50), .A3(n9839), .ZN(n9840) );
  NAND4_X1 U10935 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n9844)
         );
  NOR4_X1 U10936 ( .A1(n9847), .A2(n9846), .A3(n9845), .A4(n9844), .ZN(n9897)
         );
  NAND2_X1 U10937 ( .A1(keyinput125), .A2(keyinput49), .ZN(n9848) );
  NOR3_X1 U10938 ( .A1(keyinput94), .A2(keyinput81), .A3(n9848), .ZN(n9849) );
  NAND3_X1 U10939 ( .A1(keyinput5), .A2(keyinput53), .A3(n9849), .ZN(n9862) );
  INV_X1 U10940 ( .A(keyinput123), .ZN(n9850) );
  NOR4_X1 U10941 ( .A1(keyinput78), .A2(keyinput23), .A3(keyinput120), .A4(
        n9850), .ZN(n9860) );
  NAND2_X1 U10942 ( .A1(keyinput57), .A2(keyinput77), .ZN(n9851) );
  NOR3_X1 U10943 ( .A1(keyinput38), .A2(keyinput39), .A3(n9851), .ZN(n9859) );
  NOR2_X1 U10944 ( .A1(keyinput9), .A2(keyinput89), .ZN(n9852) );
  NAND3_X1 U10945 ( .A1(keyinput85), .A2(keyinput8), .A3(n9852), .ZN(n9857) );
  NAND4_X1 U10946 ( .A1(keyinput99), .A2(keyinput98), .A3(keyinput51), .A4(
        keyinput47), .ZN(n9856) );
  INV_X1 U10947 ( .A(keyinput80), .ZN(n9853) );
  NAND4_X1 U10948 ( .A1(keyinput67), .A2(keyinput68), .A3(keyinput24), .A4(
        n9853), .ZN(n9855) );
  NAND4_X1 U10949 ( .A1(keyinput90), .A2(keyinput110), .A3(keyinput22), .A4(
        keyinput42), .ZN(n9854) );
  NOR4_X1 U10950 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(n9858)
         );
  NAND3_X1 U10951 ( .A1(n9860), .A2(n9859), .A3(n9858), .ZN(n9861) );
  NOR4_X1 U10952 ( .A1(keyinput104), .A2(keyinput34), .A3(n9862), .A4(n9861), 
        .ZN(n9896) );
  NAND2_X1 U10953 ( .A1(keyinput58), .A2(keyinput69), .ZN(n9863) );
  NOR3_X1 U10954 ( .A1(keyinput108), .A2(keyinput61), .A3(n9863), .ZN(n9865)
         );
  INV_X1 U10955 ( .A(keyinput105), .ZN(n9864) );
  NAND3_X1 U10956 ( .A1(keyinput86), .A2(n9865), .A3(n9864), .ZN(n9877) );
  NOR2_X1 U10957 ( .A1(keyinput70), .A2(keyinput54), .ZN(n9866) );
  NAND3_X1 U10958 ( .A1(keyinput25), .A2(keyinput55), .A3(n9866), .ZN(n9867)
         );
  NOR3_X1 U10959 ( .A1(keyinput56), .A2(keyinput2), .A3(n9867), .ZN(n9875) );
  NOR2_X1 U10960 ( .A1(keyinput37), .A2(keyinput87), .ZN(n9868) );
  NAND3_X1 U10961 ( .A1(keyinput107), .A2(keyinput74), .A3(n9868), .ZN(n9873)
         );
  NAND4_X1 U10962 ( .A1(keyinput60), .A2(keyinput64), .A3(keyinput46), .A4(
        keyinput115), .ZN(n9872) );
  NOR2_X1 U10963 ( .A1(keyinput92), .A2(keyinput33), .ZN(n9869) );
  NAND3_X1 U10964 ( .A1(keyinput41), .A2(keyinput0), .A3(n9869), .ZN(n9871) );
  NAND4_X1 U10965 ( .A1(keyinput29), .A2(keyinput106), .A3(keyinput28), .A4(
        keyinput71), .ZN(n9870) );
  NOR4_X1 U10966 ( .A1(n9873), .A2(n9872), .A3(n9871), .A4(n9870), .ZN(n9874)
         );
  NAND4_X1 U10967 ( .A1(keyinput4), .A2(keyinput83), .A3(n9875), .A4(n9874), 
        .ZN(n9876) );
  NOR4_X1 U10968 ( .A1(keyinput6), .A2(keyinput10), .A3(n9877), .A4(n9876), 
        .ZN(n9895) );
  NAND2_X1 U10969 ( .A1(keyinput102), .A2(keyinput1), .ZN(n9878) );
  NOR3_X1 U10970 ( .A1(keyinput113), .A2(keyinput119), .A3(n9878), .ZN(n9879)
         );
  NAND3_X1 U10971 ( .A1(keyinput100), .A2(keyinput35), .A3(n9879), .ZN(n9893)
         );
  INV_X1 U10972 ( .A(keyinput72), .ZN(n9880) );
  NAND4_X1 U10973 ( .A1(keyinput30), .A2(keyinput26), .A3(keyinput45), .A4(
        n9880), .ZN(n9881) );
  NOR3_X1 U10974 ( .A1(keyinput40), .A2(keyinput27), .A3(n9881), .ZN(n9891) );
  INV_X1 U10975 ( .A(keyinput18), .ZN(n9882) );
  NAND4_X1 U10976 ( .A1(keyinput82), .A2(keyinput116), .A3(keyinput73), .A4(
        n9882), .ZN(n9889) );
  NOR2_X1 U10977 ( .A1(keyinput19), .A2(keyinput95), .ZN(n9883) );
  NAND3_X1 U10978 ( .A1(keyinput84), .A2(keyinput88), .A3(n9883), .ZN(n9888)
         );
  NOR2_X1 U10979 ( .A1(keyinput59), .A2(keyinput126), .ZN(n9884) );
  NAND3_X1 U10980 ( .A1(keyinput21), .A2(keyinput66), .A3(n9884), .ZN(n9887)
         );
  NOR2_X1 U10981 ( .A1(keyinput112), .A2(keyinput117), .ZN(n9885) );
  NAND3_X1 U10982 ( .A1(keyinput65), .A2(keyinput3), .A3(n9885), .ZN(n9886) );
  NOR4_X1 U10983 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9890)
         );
  NAND4_X1 U10984 ( .A1(keyinput76), .A2(keyinput44), .A3(n9891), .A4(n9890), 
        .ZN(n9892) );
  NOR4_X1 U10985 ( .A1(keyinput14), .A2(keyinput114), .A3(n9893), .A4(n9892), 
        .ZN(n9894) );
  NAND4_X1 U10986 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9898)
         );
  NAND2_X1 U10987 ( .A1(n9898), .A2(keyinput13), .ZN(n9899) );
  MUX2_X1 U10988 ( .A(keyinput13), .B(n9899), .S(P2_IR_REG_21__SCAN_IN), .Z(
        n10143) );
  INV_X1 U10989 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U10990 ( .A1(n9902), .A2(keyinput43), .B1(n9901), .B2(keyinput94), 
        .ZN(n9900) );
  OAI221_X1 U10991 ( .B1(n9902), .B2(keyinput43), .C1(n9901), .C2(keyinput94), 
        .A(n9900), .ZN(n9913) );
  INV_X1 U10992 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9905) );
  INV_X1 U10993 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10994 ( .A1(n9905), .A2(keyinput50), .B1(n9904), .B2(keyinput62), 
        .ZN(n9903) );
  OAI221_X1 U10995 ( .B1(n9905), .B2(keyinput50), .C1(n9904), .C2(keyinput62), 
        .A(n9903), .ZN(n9912) );
  INV_X1 U10996 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9906) );
  XOR2_X1 U10997 ( .A(n9906), .B(keyinput11), .Z(n9910) );
  XNOR2_X1 U10998 ( .A(keyinput103), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9909)
         );
  XNOR2_X1 U10999 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput124), .ZN(n9908) );
  XNOR2_X1 U11000 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput127), .ZN(n9907) );
  NAND4_X1 U11001 ( .A1(n9910), .A2(n9909), .A3(n9908), .A4(n9907), .ZN(n9911)
         );
  NOR3_X1 U11002 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9960) );
  INV_X1 U11003 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U11004 ( .A1(n9916), .A2(keyinput101), .B1(keyinput75), .B2(n9915), 
        .ZN(n9914) );
  OAI221_X1 U11005 ( .B1(n9916), .B2(keyinput101), .C1(n9915), .C2(keyinput75), 
        .A(n9914), .ZN(n9927) );
  AOI22_X1 U11006 ( .A1(n9919), .A2(keyinput17), .B1(keyinput79), .B2(n9918), 
        .ZN(n9917) );
  OAI221_X1 U11007 ( .B1(n9919), .B2(keyinput17), .C1(n9918), .C2(keyinput79), 
        .A(n9917), .ZN(n9926) );
  AOI22_X1 U11008 ( .A1(n7456), .A2(keyinput31), .B1(n9921), .B2(keyinput52), 
        .ZN(n9920) );
  OAI221_X1 U11009 ( .B1(n7456), .B2(keyinput31), .C1(n9921), .C2(keyinput52), 
        .A(n9920), .ZN(n9925) );
  AOI22_X1 U11010 ( .A1(n5602), .A2(keyinput36), .B1(keyinput12), .B2(n9923), 
        .ZN(n9922) );
  OAI221_X1 U11011 ( .B1(n5602), .B2(keyinput36), .C1(n9923), .C2(keyinput12), 
        .A(n9922), .ZN(n9924) );
  NOR4_X1 U11012 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9959)
         );
  INV_X1 U11013 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U11014 ( .A1(n9930), .A2(keyinput120), .B1(keyinput105), .B2(n9929), 
        .ZN(n9928) );
  OAI221_X1 U11015 ( .B1(n9930), .B2(keyinput120), .C1(n9929), .C2(keyinput105), .A(n9928), .ZN(n9941) );
  AOI22_X1 U11016 ( .A1(n9932), .A2(keyinput38), .B1(keyinput57), .B2(n6890), 
        .ZN(n9931) );
  OAI221_X1 U11017 ( .B1(n9932), .B2(keyinput38), .C1(n6890), .C2(keyinput57), 
        .A(n9931), .ZN(n9940) );
  AOI22_X1 U11018 ( .A1(n9935), .A2(keyinput39), .B1(keyinput78), .B2(n9934), 
        .ZN(n9933) );
  OAI221_X1 U11019 ( .B1(n9935), .B2(keyinput39), .C1(n9934), .C2(keyinput78), 
        .A(n9933), .ZN(n9939) );
  XNOR2_X1 U11020 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput23), .ZN(n9937) );
  XNOR2_X1 U11021 ( .A(SI_12_), .B(keyinput123), .ZN(n9936) );
  NAND2_X1 U11022 ( .A1(n9937), .A2(n9936), .ZN(n9938) );
  NOR4_X1 U11023 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9958)
         );
  AOI22_X1 U11024 ( .A1(n9943), .A2(keyinput42), .B1(keyinput67), .B2(n7435), 
        .ZN(n9942) );
  OAI221_X1 U11025 ( .B1(n9943), .B2(keyinput42), .C1(n7435), .C2(keyinput67), 
        .A(n9942), .ZN(n9956) );
  INV_X1 U11026 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U11027 ( .A1(n9946), .A2(keyinput110), .B1(n9945), .B2(keyinput22), 
        .ZN(n9944) );
  OAI221_X1 U11028 ( .B1(n9946), .B2(keyinput110), .C1(n9945), .C2(keyinput22), 
        .A(n9944), .ZN(n9955) );
  AOI22_X1 U11029 ( .A1(n9949), .A2(keyinput24), .B1(n9948), .B2(keyinput77), 
        .ZN(n9947) );
  OAI221_X1 U11030 ( .B1(n9949), .B2(keyinput24), .C1(n9948), .C2(keyinput77), 
        .A(n9947), .ZN(n9954) );
  AOI22_X1 U11031 ( .A1(n9952), .A2(keyinput80), .B1(n9951), .B2(keyinput68), 
        .ZN(n9950) );
  OAI221_X1 U11032 ( .B1(n9952), .B2(keyinput80), .C1(n9951), .C2(keyinput68), 
        .A(n9950), .ZN(n9953) );
  NOR4_X1 U11033 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(n9957)
         );
  NAND4_X1 U11034 ( .A1(n9960), .A2(n9959), .A3(n9958), .A4(n9957), .ZN(n9990)
         );
  INV_X1 U11035 ( .A(keyinput108), .ZN(n9962) );
  AOI22_X1 U11036 ( .A1(n9963), .A2(keyinput58), .B1(P2_WR_REG_SCAN_IN), .B2(
        n9962), .ZN(n9961) );
  OAI221_X1 U11037 ( .B1(n9963), .B2(keyinput58), .C1(n9962), .C2(
        P2_WR_REG_SCAN_IN), .A(n9961), .ZN(n9969) );
  INV_X1 U11038 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U11039 ( .A1(n6393), .A2(keyinput61), .B1(keyinput6), .B2(n9965), 
        .ZN(n9964) );
  OAI221_X1 U11040 ( .B1(n6393), .B2(keyinput61), .C1(n9965), .C2(keyinput6), 
        .A(n9964), .ZN(n9968) );
  XNOR2_X1 U11041 ( .A(n9966), .B(keyinput65), .ZN(n9967) );
  NOR3_X1 U11042 ( .A1(n9969), .A2(n9968), .A3(n9967), .ZN(n9988) );
  INV_X1 U11043 ( .A(SI_18_), .ZN(n9972) );
  INV_X1 U11044 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9971) );
  OAI22_X1 U11045 ( .A1(n9972), .A2(keyinput81), .B1(n9971), .B2(keyinput99), 
        .ZN(n9970) );
  AOI221_X1 U11046 ( .B1(n9972), .B2(keyinput81), .C1(keyinput99), .C2(n9971), 
        .A(n9970), .ZN(n9987) );
  INV_X1 U11047 ( .A(keyinput45), .ZN(n9973) );
  XNOR2_X1 U11048 ( .A(n9974), .B(n9973), .ZN(n9986) );
  XNOR2_X1 U11049 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput10), .ZN(n9978) );
  XNOR2_X1 U11050 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput117), .ZN(n9977)
         );
  XNOR2_X1 U11051 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput21), .ZN(n9976) );
  XNOR2_X1 U11052 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput3), .ZN(n9975) );
  NAND4_X1 U11053 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n9984)
         );
  XNOR2_X1 U11054 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput40), .ZN(n9982) );
  XNOR2_X1 U11055 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput30), .ZN(n9981) );
  XNOR2_X1 U11056 ( .A(keyinput26), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9980) );
  XNOR2_X1 U11057 ( .A(keyinput69), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9979) );
  NAND4_X1 U11058 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n9983)
         );
  NOR2_X1 U11059 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  NAND4_X1 U11060 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n9989)
         );
  NOR2_X1 U11061 ( .A1(n9990), .A2(n9989), .ZN(n10031) );
  INV_X1 U11062 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11063 ( .A1(n9993), .A2(keyinput66), .B1(keyinput76), .B2(n9992), 
        .ZN(n9991) );
  OAI221_X1 U11064 ( .B1(n9993), .B2(keyinput66), .C1(n9992), .C2(keyinput76), 
        .A(n9991), .ZN(n9999) );
  INV_X1 U11065 ( .A(P1_B_REG_SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11066 ( .A1(n9996), .A2(keyinput27), .B1(n9995), .B2(keyinput113), 
        .ZN(n9994) );
  OAI221_X1 U11067 ( .B1(n9996), .B2(keyinput27), .C1(n9995), .C2(keyinput113), 
        .A(n9994), .ZN(n9998) );
  XOR2_X1 U11068 ( .A(P2_D_REG_19__SCAN_IN), .B(keyinput111), .Z(n9997) );
  NOR3_X1 U11069 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10022) );
  OAI22_X1 U11070 ( .A1(n10002), .A2(keyinput91), .B1(n10001), .B2(keyinput93), 
        .ZN(n10000) );
  AOI221_X1 U11071 ( .B1(n10002), .B2(keyinput91), .C1(keyinput93), .C2(n10001), .A(n10000), .ZN(n10021) );
  INV_X1 U11072 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U11073 ( .A1(n6850), .A2(keyinput44), .B1(n10004), .B2(keyinput72), 
        .ZN(n10003) );
  OAI221_X1 U11074 ( .B1(n6850), .B2(keyinput44), .C1(n10004), .C2(keyinput72), 
        .A(n10003), .ZN(n10008) );
  INV_X1 U11075 ( .A(SI_3_), .ZN(n10006) );
  AOI22_X1 U11076 ( .A1(n6051), .A2(keyinput126), .B1(n10006), .B2(keyinput59), 
        .ZN(n10005) );
  OAI221_X1 U11077 ( .B1(n6051), .B2(keyinput126), .C1(n10006), .C2(keyinput59), .A(n10005), .ZN(n10007) );
  NOR2_X1 U11078 ( .A1(n10008), .A2(n10007), .ZN(n10020) );
  XNOR2_X1 U11079 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput48), .ZN(n10012) );
  XNOR2_X1 U11080 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput49), .ZN(n10011)
         );
  XNOR2_X1 U11081 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput98), .ZN(n10010) );
  XNOR2_X1 U11082 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput32), .ZN(n10009) );
  NAND4_X1 U11083 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10018) );
  XNOR2_X1 U11084 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput85), .ZN(n10016)
         );
  XNOR2_X1 U11085 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput86), .ZN(n10015) );
  XNOR2_X1 U11086 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput5), .ZN(n10014) );
  XNOR2_X1 U11087 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput60), .ZN(n10013)
         );
  NAND4_X1 U11088 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10017) );
  NOR2_X1 U11089 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  AND4_X1 U11090 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10030) );
  INV_X1 U11091 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10024) );
  OAI22_X1 U11092 ( .A1(n10146), .A2(keyinput8), .B1(n10024), .B2(keyinput90), 
        .ZN(n10023) );
  AOI221_X1 U11093 ( .B1(n10146), .B2(keyinput8), .C1(keyinput90), .C2(n10024), 
        .A(n10023), .ZN(n10029) );
  OAI22_X1 U11094 ( .A1(n10027), .A2(keyinput53), .B1(n10026), .B2(keyinput104), .ZN(n10025) );
  AOI221_X1 U11095 ( .B1(n10027), .B2(keyinput53), .C1(keyinput104), .C2(
        n10026), .A(n10025), .ZN(n10028) );
  NAND4_X1 U11096 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10141) );
  OAI22_X1 U11097 ( .A1(n10033), .A2(keyinput34), .B1(n6245), .B2(keyinput125), 
        .ZN(n10032) );
  AOI221_X1 U11098 ( .B1(n10033), .B2(keyinput34), .C1(keyinput125), .C2(n6245), .A(n10032), .ZN(n10044) );
  OAI22_X1 U11099 ( .A1(n6182), .A2(keyinput121), .B1(n10035), .B2(keyinput15), 
        .ZN(n10034) );
  AOI221_X1 U11100 ( .B1(n6182), .B2(keyinput121), .C1(keyinput15), .C2(n10035), .A(n10034), .ZN(n10043) );
  INV_X1 U11101 ( .A(SI_30_), .ZN(n10037) );
  OAI22_X1 U11102 ( .A1(n10038), .A2(keyinput47), .B1(n10037), .B2(keyinput89), 
        .ZN(n10036) );
  AOI221_X1 U11103 ( .B1(n10038), .B2(keyinput47), .C1(keyinput89), .C2(n10037), .A(n10036), .ZN(n10042) );
  OAI22_X1 U11104 ( .A1(n10040), .A2(keyinput9), .B1(n8435), .B2(keyinput51), 
        .ZN(n10039) );
  AOI221_X1 U11105 ( .B1(n10040), .B2(keyinput9), .C1(keyinput51), .C2(n8435), 
        .A(n10039), .ZN(n10041) );
  NAND4_X1 U11106 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10140) );
  AOI22_X1 U11107 ( .A1(n10047), .A2(keyinput106), .B1(n10046), .B2(keyinput28), .ZN(n10045) );
  OAI221_X1 U11108 ( .B1(n10047), .B2(keyinput106), .C1(n10046), .C2(
        keyinput28), .A(n10045), .ZN(n10059) );
  AOI22_X1 U11109 ( .A1(n10050), .A2(keyinput71), .B1(n10049), .B2(keyinput92), 
        .ZN(n10048) );
  OAI221_X1 U11110 ( .B1(n10050), .B2(keyinput71), .C1(n10049), .C2(keyinput92), .A(n10048), .ZN(n10058) );
  INV_X1 U11111 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n10053) );
  INV_X1 U11112 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U11113 ( .A1(n10053), .A2(keyinput41), .B1(n10052), .B2(keyinput33), 
        .ZN(n10051) );
  OAI221_X1 U11114 ( .B1(n10053), .B2(keyinput41), .C1(n10052), .C2(keyinput33), .A(n10051), .ZN(n10057) );
  AOI22_X1 U11115 ( .A1(n6931), .A2(keyinput0), .B1(n10055), .B2(keyinput70), 
        .ZN(n10054) );
  OAI221_X1 U11116 ( .B1(n6931), .B2(keyinput0), .C1(n10055), .C2(keyinput70), 
        .A(n10054), .ZN(n10056) );
  NOR4_X1 U11117 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10075) );
  AOI22_X1 U11118 ( .A1(n10061), .A2(keyinput25), .B1(keyinput4), .B2(n6071), 
        .ZN(n10060) );
  OAI221_X1 U11119 ( .B1(n10061), .B2(keyinput25), .C1(n6071), .C2(keyinput4), 
        .A(n10060), .ZN(n10073) );
  AOI22_X1 U11120 ( .A1(n10064), .A2(keyinput83), .B1(keyinput55), .B2(n10063), 
        .ZN(n10062) );
  OAI221_X1 U11121 ( .B1(n10064), .B2(keyinput83), .C1(n10063), .C2(keyinput55), .A(n10062), .ZN(n10072) );
  AOI22_X1 U11122 ( .A1(n10067), .A2(keyinput54), .B1(n10066), .B2(keyinput56), 
        .ZN(n10065) );
  OAI221_X1 U11123 ( .B1(n10067), .B2(keyinput54), .C1(n10066), .C2(keyinput56), .A(n10065), .ZN(n10071) );
  INV_X1 U11124 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U11125 ( .A1(n10069), .A2(keyinput2), .B1(n5845), .B2(keyinput19), 
        .ZN(n10068) );
  OAI221_X1 U11126 ( .B1(n10069), .B2(keyinput2), .C1(n5845), .C2(keyinput19), 
        .A(n10068), .ZN(n10070) );
  NOR4_X1 U11127 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10074) );
  NAND2_X1 U11128 ( .A1(n10075), .A2(n10074), .ZN(n10139) );
  AOI22_X1 U11129 ( .A1(n10078), .A2(keyinput84), .B1(keyinput88), .B2(n10077), 
        .ZN(n10076) );
  OAI221_X1 U11130 ( .B1(n10078), .B2(keyinput84), .C1(n10077), .C2(keyinput88), .A(n10076), .ZN(n10088) );
  AOI22_X1 U11131 ( .A1(n10080), .A2(keyinput95), .B1(keyinput116), .B2(n9375), 
        .ZN(n10079) );
  OAI221_X1 U11132 ( .B1(n10080), .B2(keyinput95), .C1(n9375), .C2(keyinput116), .A(n10079), .ZN(n10087) );
  INV_X1 U11133 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11134 ( .A1(n10082), .A2(keyinput82), .B1(keyinput73), .B2(
        P2_U3152), .ZN(n10081) );
  OAI221_X1 U11135 ( .B1(n10082), .B2(keyinput82), .C1(P2_U3152), .C2(
        keyinput73), .A(n10081), .ZN(n10086) );
  AOI22_X1 U11136 ( .A1(n10084), .A2(keyinput18), .B1(keyinput112), .B2(n6010), 
        .ZN(n10083) );
  OAI221_X1 U11137 ( .B1(n10084), .B2(keyinput18), .C1(n6010), .C2(keyinput112), .A(n10083), .ZN(n10085) );
  NOR4_X1 U11138 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10137) );
  AOI22_X1 U11139 ( .A1(n10091), .A2(keyinput7), .B1(n10090), .B2(keyinput109), 
        .ZN(n10089) );
  OAI221_X1 U11140 ( .B1(n10091), .B2(keyinput7), .C1(n10090), .C2(keyinput109), .A(n10089), .ZN(n10103) );
  INV_X1 U11141 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11142 ( .A1(n10094), .A2(keyinput20), .B1(n10093), .B2(keyinput118), .ZN(n10092) );
  OAI221_X1 U11143 ( .B1(n10094), .B2(keyinput20), .C1(n10093), .C2(
        keyinput118), .A(n10092), .ZN(n10102) );
  AOI22_X1 U11144 ( .A1(n10155), .A2(keyinput63), .B1(n10096), .B2(keyinput122), .ZN(n10095) );
  OAI221_X1 U11145 ( .B1(n10155), .B2(keyinput63), .C1(n10096), .C2(
        keyinput122), .A(n10095), .ZN(n10101) );
  INV_X1 U11146 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10099) );
  INV_X1 U11147 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U11148 ( .A1(n10099), .A2(keyinput97), .B1(keyinput16), .B2(n10098), 
        .ZN(n10097) );
  OAI221_X1 U11149 ( .B1(n10099), .B2(keyinput97), .C1(n10098), .C2(keyinput16), .A(n10097), .ZN(n10100) );
  NOR4_X1 U11150 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10136) );
  AOI22_X1 U11151 ( .A1(n10106), .A2(keyinput64), .B1(n10105), .B2(keyinput37), 
        .ZN(n10104) );
  OAI221_X1 U11152 ( .B1(n10106), .B2(keyinput64), .C1(n10105), .C2(keyinput37), .A(n10104), .ZN(n10117) );
  AOI22_X1 U11153 ( .A1(n10108), .A2(keyinput107), .B1(keyinput46), .B2(n8345), 
        .ZN(n10107) );
  OAI221_X1 U11154 ( .B1(n10108), .B2(keyinput107), .C1(n8345), .C2(keyinput46), .A(n10107), .ZN(n10116) );
  AOI22_X1 U11155 ( .A1(n10110), .A2(keyinput115), .B1(n6271), .B2(keyinput87), 
        .ZN(n10109) );
  OAI221_X1 U11156 ( .B1(n10110), .B2(keyinput115), .C1(n6271), .C2(keyinput87), .A(n10109), .ZN(n10115) );
  AOI22_X1 U11157 ( .A1(n10113), .A2(keyinput74), .B1(n10112), .B2(keyinput29), 
        .ZN(n10111) );
  OAI221_X1 U11158 ( .B1(n10113), .B2(keyinput74), .C1(n10112), .C2(keyinput29), .A(n10111), .ZN(n10114) );
  NOR4_X1 U11159 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10135) );
  AOI22_X1 U11160 ( .A1(n10120), .A2(keyinput1), .B1(n10119), .B2(keyinput119), 
        .ZN(n10118) );
  OAI221_X1 U11161 ( .B1(n10120), .B2(keyinput1), .C1(n10119), .C2(keyinput119), .A(n10118), .ZN(n10133) );
  AOI22_X1 U11162 ( .A1(n10123), .A2(keyinput102), .B1(keyinput100), .B2(
        n10122), .ZN(n10121) );
  OAI221_X1 U11163 ( .B1(n10123), .B2(keyinput102), .C1(n10122), .C2(
        keyinput100), .A(n10121), .ZN(n10132) );
  AOI22_X1 U11164 ( .A1(n10126), .A2(keyinput35), .B1(n10125), .B2(keyinput14), 
        .ZN(n10124) );
  OAI221_X1 U11165 ( .B1(n10126), .B2(keyinput35), .C1(n10125), .C2(keyinput14), .A(n10124), .ZN(n10131) );
  AOI22_X1 U11166 ( .A1(n10129), .A2(keyinput96), .B1(n10128), .B2(keyinput114), .ZN(n10127) );
  OAI221_X1 U11167 ( .B1(n10129), .B2(keyinput96), .C1(n10128), .C2(
        keyinput114), .A(n10127), .ZN(n10130) );
  NOR4_X1 U11168 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  NAND4_X1 U11169 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  OR4_X1 U11170 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10142) );
  NOR2_X1 U11171 ( .A1(n10143), .A2(n10142), .ZN(n10148) );
  MUX2_X1 U11172 ( .A(n10146), .B(n10145), .S(n10144), .Z(n10147) );
  XNOR2_X1 U11173 ( .A(n10148), .B(n10147), .ZN(P1_U3578) );
  XOR2_X1 U11174 ( .A(n10149), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11175 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  XNOR2_X1 U11176 ( .A(n10152), .B(n6010), .ZN(ADD_1071_U51) );
  OAI21_X1 U11177 ( .B1(n10155), .B2(n10154), .A(n10153), .ZN(n10156) );
  XNOR2_X1 U11178 ( .A(n10156), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11179 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(ADD_1071_U47) );
  XOR2_X1 U11180 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10160), .Z(ADD_1071_U48) );
  XOR2_X1 U11181 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10161), .Z(ADD_1071_U49) );
  XOR2_X1 U11182 ( .A(n10163), .B(n10162), .Z(ADD_1071_U54) );
  XOR2_X1 U11183 ( .A(n10165), .B(n10164), .Z(ADD_1071_U53) );
  XNOR2_X1 U11184 ( .A(n10167), .B(n10166), .ZN(ADD_1071_U52) );
endmodule

