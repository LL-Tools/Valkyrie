

module b14_C_gen_AntiSAT_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4727, n4728;

  OR2_X1 U2284 ( .A1(n3606), .A2(n3831), .ZN(n2213) );
  NAND2_X1 U2286 ( .A1(n2293), .A2(n2292), .ZN(n2377) );
  INV_X1 U2287 ( .A(n3913), .ZN(n2640) );
  INV_X1 U2288 ( .A(n2378), .ZN(n2362) );
  OAI21_X1 U2289 ( .B1(n3609), .B2(n3902), .A(n3241), .ZN(n3336) );
  XNOR2_X1 U2290 ( .A(n2682), .B(IR_REG_24__SCAN_IN), .ZN(n2689) );
  XNOR2_X1 U2291 ( .A(n2368), .B(IR_REG_1__SCAN_IN), .ZN(n4390) );
  NAND3_X2 U2292 ( .A1(n2375), .A2(n2374), .A3(n2373), .ZN(n2815) );
  INV_X2 U2293 ( .A(n3692), .ZN(n2045) );
  OAI21_X1 U2294 ( .B1(n3829), .B2(n3604), .A(n3830), .ZN(n3605) );
  INV_X8 U2295 ( .A(n3273), .ZN(n3693) );
  INV_X4 U2296 ( .A(n2860), .ZN(n3273) );
  NOR2_X2 U2297 ( .A1(n2900), .A2(n2901), .ZN(n2948) );
  INV_X1 U2298 ( .A(n3912), .ZN(n2169) );
  OAI22_X2 U2299 ( .A1(n4043), .A2(n2597), .B1(n3876), .B2(n4236), .ZN(n4024)
         );
  MUX2_X1 U2300 ( .A(n2666), .B(n2665), .S(IR_REG_28__SCAN_IN), .Z(n2042) );
  INV_X1 U2301 ( .A(n2369), .ZN(n2305) );
  NOR2_X2 U2302 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4471), .ZN(n4472) );
  AOI22_X2 U2303 ( .A1(n3336), .A2(n2508), .B1(n4309), .B2(n3891), .ZN(n3571)
         );
  BUF_X2 U2304 ( .A(n2943), .Z(n3694) );
  INV_X2 U2305 ( .A(n2949), .ZN(n2087) );
  NAND2_X1 U2306 ( .A1(n2345), .A2(n2061), .ZN(n3912) );
  INV_X2 U2308 ( .A(n2527), .ZN(n2361) );
  INV_X4 U2309 ( .A(n2527), .ZN(n2337) );
  NAND2_X1 U2310 ( .A1(n2091), .A2(n3162), .ZN(n3165) );
  NOR2_X1 U2311 ( .A1(n3019), .A2(n3109), .ZN(n2093) );
  OR2_X1 U2312 ( .A1(n2220), .A2(n3021), .ZN(n2219) );
  OAI22_X1 U2313 ( .A1(n3979), .A2(n3978), .B1(n4382), .B2(n3977), .ZN(n4396)
         );
  OR2_X1 U2314 ( .A1(n3017), .A2(n3016), .ZN(n2224) );
  CLKBUF_X3 U2315 ( .A(n3692), .Z(n2044) );
  INV_X1 U2316 ( .A(n2879), .ZN(n2916) );
  NAND2_X1 U2317 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  INV_X2 U2318 ( .A(n2377), .ZN(n3404) );
  OR2_X1 U2319 ( .A1(n2826), .A2(n2118), .ZN(n2117) );
  INV_X1 U2320 ( .A(n2292), .ZN(n4378) );
  NAND2_X1 U2321 ( .A1(n2139), .A2(n2137), .ZN(n2292) );
  INV_X1 U2322 ( .A(n4380), .ZN(n3455) );
  XNOR2_X1 U2324 ( .A(n2633), .B(IR_REG_21__SCAN_IN), .ZN(n4380) );
  XNOR2_X1 U2325 ( .A(n2634), .B(IR_REG_19__SCAN_IN), .ZN(n4381) );
  INV_X1 U2326 ( .A(n3584), .ZN(n2706) );
  AND2_X1 U2327 ( .A1(n2686), .A2(n2685), .ZN(n3584) );
  OAI21_X1 U2328 ( .B1(n2550), .B2(IR_REG_19__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2094) );
  NAND2_X1 U2329 ( .A1(n2730), .A2(IR_REG_31__SCAN_IN), .ZN(n2291) );
  AND3_X1 U2330 ( .A1(n2283), .A2(n2402), .A3(n2260), .ZN(n2541) );
  AND2_X1 U2331 ( .A1(n2283), .A2(n2288), .ZN(n2211) );
  INV_X1 U2332 ( .A(n2279), .ZN(n2260) );
  AND4_X1 U2333 ( .A1(n2317), .A2(n2281), .A3(n2282), .A4(n2280), .ZN(n2283)
         );
  AND4_X1 U2334 ( .A1(n2287), .A2(n2286), .A3(n2285), .A4(n2284), .ZN(n2288)
         );
  NAND4_X1 U2335 ( .A1(n2437), .A2(n2401), .A3(n2425), .A4(n2434), .ZN(n2279)
         );
  INV_X1 U2336 ( .A(IR_REG_7__SCAN_IN), .ZN(n2434) );
  INV_X1 U2337 ( .A(IR_REG_6__SCAN_IN), .ZN(n2425) );
  INV_X1 U2338 ( .A(IR_REG_5__SCAN_IN), .ZN(n2401) );
  INV_X1 U2339 ( .A(IR_REG_3__SCAN_IN), .ZN(n2356) );
  NOR2_X1 U2340 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2281)
         );
  NOR2_X1 U2341 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2282)
         );
  NOR2_X1 U2342 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2280)
         );
  NOR2_X1 U2343 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2317)
         );
  OAI21_X2 U2344 ( .B1(n2680), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2690) );
  AND2_X1 U2345 ( .A1(n2890), .A2(n2637), .ZN(n4317) );
  AOI21_X2 U2348 ( .B1(n3774), .B2(n3775), .A(n3777), .ZN(n3872) );
  NAND2_X2 U2349 ( .A1(n2689), .A2(n2688), .ZN(n2811) );
  INV_X1 U2350 ( .A(n2224), .ZN(n2220) );
  NAND2_X1 U2351 ( .A1(n2811), .A2(n2888), .ZN(n2860) );
  OAI22_X1 U2352 ( .A1(n3693), .A2(n2169), .B1(n2167), .B2(n2044), .ZN(n3015)
         );
  OAI22_X1 U2353 ( .A1(n3694), .A2(n2169), .B1(n3693), .B2(n2167), .ZN(n3105)
         );
  NAND2_X1 U2354 ( .A1(n3934), .A2(n2109), .ZN(n2108) );
  NAND2_X1 U2355 ( .A1(n4389), .A2(REG2_REG_2__SCAN_IN), .ZN(n2109) );
  AOI21_X1 U2356 ( .B1(n2187), .B2(n2185), .A(n2063), .ZN(n2184) );
  INV_X1 U2357 ( .A(n2058), .ZN(n2185) );
  INV_X1 U2358 ( .A(n2187), .ZN(n2186) );
  OR2_X1 U2359 ( .A1(n3912), .A2(n2167), .ZN(n3515) );
  NAND2_X1 U2360 ( .A1(n3912), .A2(n2167), .ZN(n3519) );
  OR2_X1 U2361 ( .A1(n2590), .A2(n2588), .ZN(n2600) );
  INV_X1 U2362 ( .A(n2240), .ZN(n2239) );
  OAI21_X1 U2363 ( .B1(n2245), .B2(n2243), .A(n2241), .ZN(n2240) );
  NAND2_X1 U2364 ( .A1(n2242), .A2(n2247), .ZN(n2241) );
  INV_X1 U2365 ( .A(n2244), .ZN(n2242) );
  INV_X1 U2366 ( .A(n2055), .ZN(n3613) );
  NAND2_X1 U2367 ( .A1(n2393), .A2(REG3_REG_5__SCAN_IN), .ZN(n2407) );
  OR2_X1 U2368 ( .A1(n2580), .A2(n4690), .ZN(n2590) );
  AND2_X1 U2369 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2393) );
  OR2_X1 U2370 ( .A1(n2943), .A2(n2949), .ZN(n2089) );
  INV_X1 U2371 ( .A(n3124), .ZN(n2215) );
  NAND2_X1 U2372 ( .A1(n2293), .A2(n4378), .ZN(n2379) );
  NOR2_X1 U2373 ( .A1(n2706), .A2(n2724), .ZN(n2688) );
  XNOR2_X1 U2374 ( .A(n2108), .B(n2765), .ZN(n3946) );
  AOI21_X1 U2375 ( .B1(n3994), .B2(n2112), .A(n3996), .ZN(n2111) );
  NAND2_X1 U2376 ( .A1(n2175), .A2(n2050), .ZN(n2173) );
  NAND2_X1 U2377 ( .A1(n2050), .A2(n2520), .ZN(n2174) );
  OR2_X1 U2378 ( .A1(n3323), .A2(n3284), .ZN(n2193) );
  NAND2_X1 U2379 ( .A1(n2458), .A2(n2194), .ZN(n2192) );
  NOR2_X1 U2380 ( .A1(n2195), .A2(n2469), .ZN(n2194) );
  INV_X1 U2381 ( .A(n2457), .ZN(n2195) );
  AOI22_X1 U2382 ( .A1(n2674), .A2(n4204), .B1(n4007), .B2(n3898), .ZN(n4016)
         );
  NAND2_X1 U2383 ( .A1(n2668), .A2(n2138), .ZN(n2137) );
  NOR2_X1 U2384 ( .A1(n2209), .A2(n2729), .ZN(n2138) );
  INV_X1 U2385 ( .A(n3845), .ZN(n3887) );
  NAND2_X1 U2386 ( .A1(n3962), .A2(n4426), .ZN(n4440) );
  NAND2_X1 U2387 ( .A1(n3851), .A2(n3852), .ZN(n2265) );
  NAND2_X1 U2388 ( .A1(n2661), .A2(n3430), .ZN(n2155) );
  OR2_X1 U2389 ( .A1(n3462), .A2(n3460), .ZN(n2205) );
  NAND2_X1 U2390 ( .A1(n3578), .A2(n2156), .ZN(n4150) );
  AND2_X1 U2391 ( .A1(n2157), .A2(n2051), .ZN(n2156) );
  INV_X1 U2392 ( .A(n3421), .ZN(n2157) );
  NOR2_X1 U2393 ( .A1(n2544), .A2(n4578), .ZN(n2543) );
  AND2_X1 U2394 ( .A1(n2647), .A2(n2146), .ZN(n2145) );
  NAND2_X1 U2395 ( .A1(n2147), .A2(n3496), .ZN(n2146) );
  INV_X1 U2396 ( .A(n3527), .ZN(n2166) );
  AND2_X1 U2397 ( .A1(n2098), .A2(n3813), .ZN(n2097) );
  NOR2_X1 U2398 ( .A1(n2369), .A2(n2561), .ZN(n4153) );
  AND2_X1 U2399 ( .A1(n3724), .A2(n3891), .ZN(n2100) );
  NAND2_X1 U2400 ( .A1(n3178), .A2(n3284), .ZN(n3179) );
  AND2_X1 U2401 ( .A1(n3118), .A2(n3171), .ZN(n2095) );
  INV_X1 U2402 ( .A(IR_REG_27__SCAN_IN), .ZN(n2300) );
  NOR2_X1 U2403 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2284)
         );
  NOR2_X1 U2404 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2285)
         );
  AND2_X1 U2405 ( .A1(n2260), .A2(n2289), .ZN(n2210) );
  INV_X1 U2406 ( .A(IR_REG_25__SCAN_IN), .ZN(n2289) );
  INV_X1 U2407 ( .A(IR_REG_21__SCAN_IN), .ZN(n2628) );
  INV_X1 U2408 ( .A(n3279), .ZN(n3280) );
  XNOR2_X1 U2409 ( .A(n2942), .B(n3695), .ZN(n3017) );
  NAND2_X1 U2410 ( .A1(n3699), .A2(n2244), .ZN(n2243) );
  OR2_X1 U2411 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  INV_X1 U2412 ( .A(n3019), .ZN(n2223) );
  INV_X1 U2413 ( .A(n2219), .ZN(n2218) );
  INV_X1 U2414 ( .A(n3217), .ZN(n2251) );
  NAND2_X1 U2415 ( .A1(n2253), .A2(n2057), .ZN(n2252) );
  INV_X1 U2416 ( .A(n3206), .ZN(n2253) );
  NOR2_X1 U2417 ( .A1(n3842), .A2(n2255), .ZN(n2254) );
  INV_X1 U2418 ( .A(n2257), .ZN(n2255) );
  OR2_X1 U2419 ( .A1(n2564), .A2(n3843), .ZN(n2572) );
  OAI22_X1 U2420 ( .A1(n2928), .A2(n2860), .B1(n2044), .B2(n2859), .ZN(n2863)
         );
  NAND2_X1 U2421 ( .A1(n3785), .A2(n3622), .ZN(n3624) );
  OR2_X1 U2422 ( .A1(n2839), .A2(n4381), .ZN(n2862) );
  AND4_X1 U2423 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n3595)
         );
  AND2_X1 U2424 ( .A1(n2352), .A2(n2351), .ZN(n2353) );
  OR2_X1 U2425 ( .A1(n2377), .A2(n2350), .ZN(n2352) );
  AND2_X1 U2426 ( .A1(n2828), .A2(REG1_REG_4__SCAN_IN), .ZN(n2826) );
  AOI21_X1 U2427 ( .B1(n3946), .B2(REG2_REG_3__SCAN_IN), .A(n2065), .ZN(n2755)
         );
  XNOR2_X1 U2428 ( .A(n2769), .B(n2113), .ZN(n2796) );
  NOR2_X1 U2429 ( .A1(n2780), .A2(n2114), .ZN(n2769) );
  NOR2_X1 U2430 ( .A1(n2787), .A2(n2115), .ZN(n2114) );
  OR2_X1 U2431 ( .A1(n3972), .A2(REG2_REG_13__SCAN_IN), .ZN(n2132) );
  NAND2_X1 U2432 ( .A1(n4462), .A2(n3991), .ZN(n3993) );
  NOR2_X1 U2433 ( .A1(n4457), .A2(n2103), .ZN(n3966) );
  AND2_X1 U2434 ( .A1(n3971), .A2(REG2_REG_15__SCAN_IN), .ZN(n2103) );
  NAND2_X1 U2435 ( .A1(n4476), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2436 ( .A1(n4511), .A2(n2526), .ZN(n2124) );
  AND2_X1 U2437 ( .A1(n3550), .A2(n2153), .ZN(n2152) );
  OR2_X1 U2438 ( .A1(n4075), .A2(n2155), .ZN(n2154) );
  AND2_X1 U2439 ( .A1(n2600), .A2(n2591), .ZN(n4054) );
  NAND2_X1 U2440 ( .A1(n2066), .A2(n2046), .ZN(n2187) );
  NAND2_X1 U2441 ( .A1(n4272), .A2(n2571), .ZN(n4092) );
  OAI21_X1 U2442 ( .B1(n2552), .B2(n2551), .A(n2270), .ZN(n4147) );
  NOR2_X1 U2443 ( .A1(n4202), .A2(n4185), .ZN(n2551) );
  OR2_X1 U2444 ( .A1(n2535), .A2(n2534), .ZN(n2544) );
  NAND2_X1 U2445 ( .A1(n2172), .A2(n2170), .ZN(n4194) );
  AOI21_X1 U2446 ( .B1(n2173), .B2(n2174), .A(n2171), .ZN(n2170) );
  NAND2_X1 U2447 ( .A1(n3571), .A2(n3570), .ZN(n3569) );
  INV_X1 U2448 ( .A(n2177), .ZN(n3243) );
  OAI21_X1 U2449 ( .B1(n3300), .B2(n2179), .A(n2178), .ZN(n2177) );
  AND2_X1 U2450 ( .A1(n3768), .A2(n3835), .ZN(n2179) );
  NAND2_X1 U2451 ( .A1(n3903), .A2(n3295), .ZN(n2178) );
  NOR2_X1 U2452 ( .A1(n3447), .A2(n2191), .ZN(n2190) );
  INV_X1 U2453 ( .A(n2193), .ZN(n2191) );
  NAND2_X1 U2454 ( .A1(n2645), .A2(n3528), .ZN(n3176) );
  OR2_X1 U2455 ( .A1(n3134), .A2(n3133), .ZN(n2645) );
  INV_X1 U2456 ( .A(n4381), .ZN(n4002) );
  OAI21_X1 U2457 ( .B1(n3054), .B2(n3053), .A(n3493), .ZN(n3041) );
  NAND2_X1 U2458 ( .A1(n4066), .A2(n4053), .ZN(n4052) );
  NAND2_X1 U2459 ( .A1(n4122), .A2(n4121), .ZN(n4272) );
  AND4_X1 U2460 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n4302)
         );
  INV_X1 U2461 ( .A(n3767), .ZN(n3596) );
  INV_X1 U2462 ( .A(n3906), .ZN(n3323) );
  INV_X1 U2463 ( .A(n3274), .ZN(n3284) );
  NAND2_X1 U2464 ( .A1(n2664), .A2(n3440), .ZN(n4204) );
  INV_X1 U2465 ( .A(n3127), .ZN(n3100) );
  INV_X1 U2466 ( .A(n4277), .ZN(n4308) );
  NAND2_X1 U2467 ( .A1(n2687), .A2(n3584), .ZN(n2737) );
  NAND2_X1 U2468 ( .A1(n2811), .A2(n2738), .ZN(n2882) );
  AND2_X1 U2469 ( .A1(n2303), .A2(n2300), .ZN(n2299) );
  AND4_X1 U2470 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n4309)
         );
  INV_X1 U2471 ( .A(n4137), .ZN(n4281) );
  AND4_X1 U2472 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n3766)
         );
  NOR2_X1 U2473 ( .A1(n2054), .A2(n3896), .ZN(n2236) );
  NAND2_X1 U2474 ( .A1(n2239), .A2(n2243), .ZN(n2238) );
  OR2_X1 U2475 ( .A1(n2378), .A2(n3925), .ZN(n2382) );
  INV_X1 U2476 ( .A(n4249), .ZN(n3779) );
  NAND2_X1 U2477 ( .A1(n2216), .A2(n2217), .ZN(n3125) );
  AND4_X1 U2478 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), .ZN(n3103)
         );
  OR2_X1 U2479 ( .A1(n2875), .A2(n2854), .ZN(n3845) );
  OR2_X1 U2480 ( .A1(n2875), .A2(n2874), .ZN(n3844) );
  NAND2_X1 U2481 ( .A1(n2954), .A2(n2953), .ZN(n3893) );
  NAND2_X1 U2482 ( .A1(n2606), .A2(n2605), .ZN(n3899) );
  OR2_X1 U2483 ( .A1(n4033), .A2(n2619), .ZN(n2606) );
  INV_X1 U2484 ( .A(n4085), .ZN(n4258) );
  INV_X1 U2485 ( .A(n4302), .ZN(n3900) );
  OR2_X1 U2486 ( .A1(n2619), .A2(n3028), .ZN(n2345) );
  NAND2_X1 U2487 ( .A1(n2754), .A2(n2753), .ZN(n3934) );
  AND2_X1 U2488 ( .A1(n2117), .A2(n2116), .ZN(n2780) );
  INV_X1 U2489 ( .A(n2781), .ZN(n2116) );
  AOI21_X1 U2490 ( .B1(n2129), .B2(n4436), .A(n2082), .ZN(n2127) );
  OR2_X1 U2491 ( .A1(n4440), .A2(n2128), .ZN(n2126) );
  NOR2_X1 U2492 ( .A1(n4459), .A2(n4458), .ZN(n4457) );
  XNOR2_X1 U2493 ( .A(n3966), .B(n3992), .ZN(n4468) );
  NAND2_X1 U2494 ( .A1(n4468), .A2(n2509), .ZN(n4467) );
  NAND2_X1 U2495 ( .A1(n4477), .A2(n4475), .ZN(n4476) );
  NAND2_X1 U2496 ( .A1(n2122), .A2(n4438), .ZN(n2121) );
  NAND2_X1 U2497 ( .A1(n2123), .A2(n4487), .ZN(n2122) );
  AOI21_X1 U2498 ( .B1(n4489), .B2(ADDR_REG_18__SCAN_IN), .A(n4488), .ZN(n2120) );
  NOR2_X1 U2499 ( .A1(n2123), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U2500 ( .A1(n2110), .A2(n2047), .ZN(n4490) );
  AND2_X1 U2501 ( .A1(n2774), .A2(n2759), .ZN(n4491) );
  INV_X1 U2502 ( .A(n3907), .ZN(n3283) );
  AND2_X1 U2503 ( .A1(n4016), .A2(n2158), .ZN(n2718) );
  AOI21_X1 U2504 ( .B1(n4012), .B2(n4531), .A(n2159), .ZN(n2158) );
  NAND2_X1 U2505 ( .A1(n2675), .A2(n2160), .ZN(n2159) );
  NAND2_X1 U2506 ( .A1(n3410), .A2(n4310), .ZN(n2160) );
  INV_X1 U2507 ( .A(n3970), .ZN(n4510) );
  AND2_X1 U2508 ( .A1(n2320), .A2(REG3_REG_15__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U2509 ( .A1(n3914), .A2(n2859), .ZN(n3505) );
  NOR2_X1 U2510 ( .A1(n2332), .A2(n4692), .ZN(n2320) );
  NOR2_X1 U2511 ( .A1(n3863), .A2(n2231), .ZN(n2230) );
  INV_X1 U2512 ( .A(n3630), .ZN(n2231) );
  NAND2_X1 U2513 ( .A1(n3689), .A2(n3688), .ZN(n2244) );
  AND2_X1 U2514 ( .A1(n3741), .A2(n2227), .ZN(n2226) );
  NAND2_X1 U2515 ( .A1(n2228), .A2(n2229), .ZN(n2227) );
  NAND2_X1 U2516 ( .A1(n2045), .A2(n3090), .ZN(n2943) );
  INV_X1 U2517 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2792) );
  INV_X1 U2518 ( .A(n2132), .ZN(n2130) );
  INV_X1 U2519 ( .A(n4480), .ZN(n2112) );
  AND2_X1 U2520 ( .A1(n2275), .A2(REG3_REG_10__SCAN_IN), .ZN(n2460) );
  INV_X1 U2521 ( .A(n2461), .ZN(n2275) );
  NOR2_X1 U2522 ( .A1(n2415), .A2(n2203), .ZN(n2202) );
  INV_X1 U2523 ( .A(n2405), .ZN(n2203) );
  INV_X1 U2524 ( .A(n2199), .ZN(n2197) );
  OAI22_X1 U2525 ( .A1(n2415), .A2(n2200), .B1(n3910), .B2(n3075), .ZN(n2199)
         );
  NAND2_X1 U2526 ( .A1(n2405), .A2(n2201), .ZN(n2200) );
  INV_X1 U2527 ( .A(n2404), .ZN(n2201) );
  NAND2_X1 U2528 ( .A1(n2151), .A2(n2149), .ZN(n3713) );
  AOI21_X1 U2529 ( .B1(n2152), .B2(n2155), .A(n2150), .ZN(n2149) );
  INV_X1 U2530 ( .A(n3412), .ZN(n2150) );
  NOR2_X1 U2531 ( .A1(n2711), .A2(n2099), .ZN(n2098) );
  INV_X1 U2532 ( .A(n4117), .ZN(n2099) );
  OR2_X1 U2533 ( .A1(n2737), .A2(n2703), .ZN(n2837) );
  INV_X1 U2534 ( .A(n2730), .ZN(n2140) );
  NOR2_X1 U2535 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2208)
         );
  NAND2_X1 U2536 ( .A1(n2541), .A2(n2540), .ZN(n2549) );
  INV_X1 U2537 ( .A(IR_REG_17__SCAN_IN), .ZN(n2540) );
  OR3_X1 U2538 ( .A1(n2477), .A2(IR_REG_12__SCAN_IN), .A3(n2318), .ZN(n2327)
         );
  OR2_X1 U2539 ( .A1(n2485), .A2(n2330), .ZN(n2332) );
  AND2_X1 U2540 ( .A1(n3615), .A2(n3614), .ZN(n3719) );
  INV_X1 U2541 ( .A(n2230), .ZN(n2229) );
  AOI21_X1 U2542 ( .B1(n2234), .B2(n2230), .A(n2079), .ZN(n2228) );
  NOR2_X1 U2543 ( .A1(n3690), .A2(n2246), .ZN(n2245) );
  INV_X1 U2544 ( .A(n3874), .ZN(n2246) );
  INV_X1 U2545 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4547) );
  OR2_X1 U2546 ( .A1(n2483), .A2(n4547), .ZN(n2485) );
  NAND2_X1 U2547 ( .A1(n2093), .A2(n2222), .ZN(n2216) );
  NAND2_X1 U2548 ( .A1(n2214), .A2(n2219), .ZN(n2217) );
  INV_X1 U2549 ( .A(n2572), .ZN(n2276) );
  INV_X1 U2550 ( .A(DATAI_0_), .ZN(n2101) );
  INV_X1 U2551 ( .A(n2262), .ZN(n2261) );
  NAND2_X1 U2552 ( .A1(n3278), .A2(n2263), .ZN(n2092) );
  OAI21_X1 U2553 ( .B1(n3280), .B2(n2264), .A(n2071), .ZN(n2262) );
  NAND2_X1 U2554 ( .A1(n3748), .A2(n3654), .ZN(n2257) );
  NAND2_X1 U2555 ( .A1(n3818), .A2(n2258), .ZN(n2256) );
  NAND2_X1 U2556 ( .A1(n2307), .A2(REG3_REG_21__SCAN_IN), .ZN(n2564) );
  AND4_X1 U2557 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n3210)
         );
  AND2_X1 U2558 ( .A1(n2768), .A2(n4387), .ZN(n2118) );
  NOR2_X1 U2559 ( .A1(n2760), .A2(n2406), .ZN(n2105) );
  NOR2_X1 U2560 ( .A1(n2760), .A2(n2113), .ZN(n2104) );
  AND2_X1 U2561 ( .A1(n2107), .A2(n2106), .ZN(n3955) );
  NAND2_X1 U2562 ( .A1(n4384), .A2(REG2_REG_7__SCAN_IN), .ZN(n2106) );
  XNOR2_X1 U2563 ( .A(n3955), .B(n4382), .ZN(n3956) );
  OR2_X1 U2564 ( .A1(n4436), .A2(n3988), .ZN(n2128) );
  NOR2_X1 U2565 ( .A1(n2130), .A2(n2131), .ZN(n2129) );
  AND2_X1 U2566 ( .A1(n2742), .A2(n2741), .ZN(n2774) );
  OAI22_X1 U2567 ( .A1(n4024), .A2(n2608), .B1(n4227), .B2(n4031), .ZN(n3706)
         );
  AOI21_X1 U2568 ( .B1(n2184), .B2(n2186), .A(n2076), .ZN(n2182) );
  OR2_X1 U2569 ( .A1(n4075), .A2(n3485), .ZN(n4060) );
  NAND2_X1 U2570 ( .A1(n2207), .A2(n2206), .ZN(n2204) );
  OAI21_X1 U2571 ( .B1(n4150), .B2(n2655), .A(n3541), .ZN(n4128) );
  NAND2_X1 U2572 ( .A1(n3578), .A2(n2051), .ZN(n4173) );
  AND3_X1 U2573 ( .A1(n2548), .A2(n2547), .A3(n2546), .ZN(n4202) );
  OR2_X1 U2574 ( .A1(n3333), .A2(n3446), .ZN(n3334) );
  NAND2_X1 U2575 ( .A1(n2143), .A2(n2141), .ZN(n3425) );
  AOI21_X1 U2576 ( .B1(n2145), .B2(n2148), .A(n2142), .ZN(n2141) );
  INV_X1 U2577 ( .A(n3496), .ZN(n2148) );
  NAND2_X1 U2578 ( .A1(n3308), .A2(n2062), .ZN(n2180) );
  NAND2_X1 U2579 ( .A1(n2460), .A2(REG3_REG_11__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U2580 ( .A1(n2144), .A2(n3496), .ZN(n3293) );
  NAND2_X1 U2581 ( .A1(n3176), .A2(n3492), .ZN(n2144) );
  NAND2_X1 U2582 ( .A1(n2440), .A2(REG3_REG_9__SCAN_IN), .ZN(n2461) );
  AOI21_X1 U2583 ( .B1(n2165), .B2(n2163), .A(n2162), .ZN(n2161) );
  INV_X1 U2584 ( .A(n2165), .ZN(n2164) );
  INV_X1 U2585 ( .A(n3524), .ZN(n2162) );
  NAND2_X1 U2586 ( .A1(n2197), .A2(n2196), .ZN(n3097) );
  AND2_X1 U2587 ( .A1(n2643), .A2(n3525), .ZN(n3522) );
  INV_X1 U2588 ( .A(n3910), .ZN(n3113) );
  OAI21_X1 U2589 ( .B1(n2981), .B2(n2641), .A(n3519), .ZN(n3054) );
  NAND2_X1 U2590 ( .A1(n2960), .A2(n3514), .ZN(n2981) );
  AND2_X1 U2591 ( .A1(n3514), .A2(n3512), .ZN(n3471) );
  NAND2_X1 U2592 ( .A1(n2911), .A2(n3509), .ZN(n2930) );
  INV_X1 U2593 ( .A(n2639), .ZN(n3472) );
  INV_X1 U2594 ( .A(n4317), .ZN(n3090) );
  OR2_X1 U2595 ( .A1(n2638), .A2(n3504), .ZN(n2911) );
  NAND2_X1 U2596 ( .A1(n2362), .A2(REG3_REG_0__SCAN_IN), .ZN(n2372) );
  AND2_X1 U2597 ( .A1(n2837), .A2(n2836), .ZN(n2886) );
  NOR3_X1 U2598 ( .A1(n4052), .A2(n2102), .A3(n4223), .ZN(n4220) );
  OR2_X1 U2599 ( .A1(n4052), .A2(n4235), .ZN(n4029) );
  AND2_X1 U2600 ( .A1(n2617), .A2(n2616), .ZN(n4238) );
  AND2_X1 U2601 ( .A1(n4133), .A2(n2083), .ZN(n4066) );
  AND2_X1 U2602 ( .A1(n2596), .A2(n2595), .ZN(n4252) );
  NAND2_X1 U2603 ( .A1(n4133), .A2(n2098), .ZN(n4102) );
  NAND2_X1 U2604 ( .A1(n4133), .A2(n4117), .ZN(n4116) );
  AND2_X1 U2605 ( .A1(n4162), .A2(n4142), .ZN(n4133) );
  NOR2_X1 U2606 ( .A1(n4184), .A2(n4153), .ZN(n4162) );
  NAND2_X1 U2607 ( .A1(n4208), .A2(n4207), .ZN(n4206) );
  OR2_X1 U2608 ( .A1(n4206), .A2(n2710), .ZN(n4184) );
  NAND2_X1 U2609 ( .A1(n3302), .A2(n2053), .ZN(n3574) );
  NOR2_X1 U2610 ( .A1(n3574), .A2(n4297), .ZN(n4208) );
  NAND2_X1 U2611 ( .A1(n3302), .A2(n2100), .ZN(n3572) );
  AND4_X1 U2612 ( .A1(n2326), .A2(n2325), .A3(n2324), .A4(n2323), .ZN(n3608)
         );
  NAND2_X1 U2613 ( .A1(n3302), .A2(n3724), .ZN(n3337) );
  INV_X1 U2614 ( .A(n3609), .ZN(n3724) );
  AND2_X1 U2615 ( .A1(n3312), .A2(n3835), .ZN(n3302) );
  NOR2_X1 U2616 ( .A1(n3311), .A2(n3596), .ZN(n3312) );
  INV_X1 U2617 ( .A(n3255), .ZN(n3857) );
  OR2_X1 U2618 ( .A1(n3179), .A2(n3255), .ZN(n3311) );
  AND2_X1 U2619 ( .A1(n3060), .A2(n2077), .ZN(n3178) );
  AND4_X1 U2620 ( .A1(n2433), .A2(n2432), .A3(n2431), .A4(n2430), .ZN(n3196)
         );
  NAND2_X1 U2621 ( .A1(n3060), .A2(n2095), .ZN(n3154) );
  NAND2_X1 U2622 ( .A1(n3060), .A2(n3118), .ZN(n3092) );
  OR2_X1 U2623 ( .A1(n2986), .A2(n2987), .ZN(n3058) );
  NOR2_X1 U2624 ( .A1(n3058), .A2(n3100), .ZN(n3060) );
  NAND2_X1 U2625 ( .A1(n2859), .A2(n2879), .ZN(n2936) );
  INV_X1 U2626 ( .A(n4314), .ZN(n4298) );
  NOR2_X1 U2627 ( .A1(n2299), .A2(n2729), .ZN(n2667) );
  INV_X1 U2628 ( .A(n2299), .ZN(n2302) );
  AND2_X1 U2629 ( .A1(n2685), .A2(n2304), .ZN(n2665) );
  AND2_X1 U2630 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2304)
         );
  NOR2_X1 U2631 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2287)
         );
  NOR2_X1 U2632 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2286)
         );
  XNOR2_X1 U2633 ( .A(n2631), .B(n2630), .ZN(n2839) );
  INV_X1 U2634 ( .A(IR_REG_20__SCAN_IN), .ZN(n2635) );
  AND2_X1 U2635 ( .A1(n2518), .A2(n2507), .ZN(n3971) );
  XNOR2_X1 U2636 ( .A(n3689), .B(n3688), .ZN(n3690) );
  INV_X1 U2637 ( .A(n3278), .ZN(n3281) );
  NAND2_X1 U2638 ( .A1(n2249), .A2(n2252), .ZN(n3218) );
  XNOR2_X1 U2639 ( .A(n2897), .B(n2212), .ZN(n2872) );
  OR2_X1 U2640 ( .A1(n2868), .A2(n3613), .ZN(n2869) );
  NAND2_X1 U2641 ( .A1(n2221), .A2(n2224), .ZN(n3020) );
  NAND2_X1 U2642 ( .A1(n2223), .A2(n2222), .ZN(n2221) );
  AND2_X1 U2643 ( .A1(n2250), .A2(n3219), .ZN(n2248) );
  OR2_X1 U2644 ( .A1(n2252), .A2(n2251), .ZN(n2250) );
  XOR2_X1 U2645 ( .A(n3268), .B(n3269), .Z(n3266) );
  AND4_X2 U2646 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .ZN(n2928)
         );
  OR2_X1 U2647 ( .A1(n2377), .A2(n2363), .ZN(n2364) );
  AND2_X1 U2648 ( .A1(n2555), .A2(n2554), .ZN(n4166) );
  NAND2_X1 U2649 ( .A1(n2256), .A2(n2257), .ZN(n3841) );
  NAND2_X1 U2650 ( .A1(n3628), .A2(n2233), .ZN(n2232) );
  INV_X1 U2651 ( .A(n4252), .ZN(n4236) );
  NAND2_X1 U2652 ( .A1(n2586), .A2(n2585), .ZN(n4249) );
  OR2_X1 U2653 ( .A1(n4080), .A2(n2619), .ZN(n2586) );
  NAND2_X1 U2654 ( .A1(n2570), .A2(n2569), .ZN(n4137) );
  INV_X1 U2655 ( .A(n4202), .ZN(n4154) );
  OAI211_X1 U2656 ( .C1(n3865), .C2(n2619), .A(n2539), .B(n2538), .ZN(n4299)
         );
  INV_X1 U2657 ( .A(n4309), .ZN(n3901) );
  INV_X1 U2658 ( .A(n3608), .ZN(n3902) );
  INV_X1 U2659 ( .A(n3595), .ZN(n3904) );
  INV_X1 U2660 ( .A(n3196), .ZN(n3908) );
  INV_X1 U2661 ( .A(n3210), .ZN(n3909) );
  NAND2_X1 U2662 ( .A1(n2059), .A2(n2355), .ZN(n3913) );
  AOI22_X1 U2663 ( .A1(n2825), .A2(REG2_REG_4__SCAN_IN), .B1(n4387), .B2(n2756), .ZN(n2785) );
  INV_X1 U2664 ( .A(n2117), .ZN(n2782) );
  AOI21_X1 U2665 ( .B1(n4385), .B2(n2770), .A(n2794), .ZN(n2803) );
  AOI21_X1 U2666 ( .B1(n2791), .B2(REG2_REG_6__SCAN_IN), .A(n2084), .ZN(n2761)
         );
  NAND2_X1 U2667 ( .A1(n4453), .A2(n3990), .ZN(n4463) );
  NAND2_X1 U2668 ( .A1(n4463), .A2(n4464), .ZN(n4462) );
  NOR2_X1 U2669 ( .A1(n4449), .A2(n3964), .ZN(n4459) );
  NAND2_X1 U2670 ( .A1(n2133), .A2(n2132), .ZN(n3963) );
  OR2_X1 U2671 ( .A1(n4440), .A2(n4436), .ZN(n2133) );
  XNOR2_X1 U2672 ( .A(n3993), .B(n3992), .ZN(n4471) );
  NAND2_X1 U2673 ( .A1(n4467), .A2(n3967), .ZN(n4475) );
  NOR2_X1 U2674 ( .A1(n4472), .A2(n3994), .ZN(n4481) );
  NOR2_X1 U2675 ( .A1(n4481), .A2(n4480), .ZN(n4482) );
  NAND2_X1 U2676 ( .A1(n2154), .A2(n2152), .ZN(n4028) );
  NAND2_X1 U2677 ( .A1(n2154), .A2(n3550), .ZN(n4026) );
  NAND2_X1 U2678 ( .A1(n2183), .A2(n2187), .ZN(n4063) );
  NAND2_X1 U2679 ( .A1(n4092), .A2(n2058), .ZN(n2183) );
  AND2_X1 U2680 ( .A1(n2188), .A2(n2189), .ZN(n4078) );
  NAND2_X1 U2681 ( .A1(n4092), .A2(n2579), .ZN(n2188) );
  NAND2_X1 U2682 ( .A1(n2298), .A2(n2297), .ZN(n4089) );
  AOI21_X1 U2683 ( .B1(n4147), .B2(n3460), .A(n3462), .ZN(n4130) );
  OAI21_X1 U2684 ( .B1(n3571), .B2(n2174), .A(n2173), .ZN(n4195) );
  NAND2_X1 U2685 ( .A1(n3578), .A2(n3500), .ZN(n3389) );
  NAND2_X1 U2686 ( .A1(n3569), .A2(n2520), .ZN(n3391) );
  NAND2_X1 U2687 ( .A1(n2192), .A2(n2193), .ZN(n3254) );
  NAND4_X1 U2688 ( .A1(n2467), .A2(n2466), .A3(n2465), .A4(n2464), .ZN(n3906)
         );
  NAND2_X1 U2689 ( .A1(n2458), .A2(n2457), .ZN(n3177) );
  OR2_X1 U2690 ( .A1(n2882), .A2(n2849), .ZN(n4496) );
  NAND2_X1 U2691 ( .A1(n2198), .A2(n2405), .ZN(n3040) );
  NAND2_X1 U2692 ( .A1(n3052), .A2(n2404), .ZN(n2198) );
  INV_X1 U2693 ( .A(n2963), .ZN(n3001) );
  OR2_X1 U2694 ( .A1(n4212), .A2(n3090), .ZN(n4187) );
  AND2_X1 U2695 ( .A1(n4191), .A2(n4277), .ZN(n4135) );
  INV_X2 U2696 ( .A(n4543), .ZN(n4545) );
  AND3_X1 U2697 ( .A1(n3352), .A2(n3351), .A3(n3350), .ZN(n3355) );
  NAND2_X1 U2698 ( .A1(n3069), .A2(n2168), .ZN(n3057) );
  AND2_X1 U2699 ( .A1(n3056), .A2(n2085), .ZN(n2168) );
  NAND2_X1 U2700 ( .A1(n2737), .A2(n2736), .ZN(n4507) );
  NAND2_X1 U2701 ( .A1(n2299), .A2(n2266), .ZN(n2730) );
  NOR2_X1 U2702 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2266)
         );
  INV_X1 U2703 ( .A(n2839), .ZN(n4379) );
  NAND2_X1 U2704 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2634) );
  OR2_X1 U2705 ( .A1(n2452), .A2(n2451), .ZN(n4520) );
  NAND2_X1 U2706 ( .A1(n2067), .A2(IR_REG_31__SCAN_IN), .ZN(n2384) );
  CLKBUF_X1 U2707 ( .A(n3915), .Z(U4043) );
  OAI22_X1 U2708 ( .A1(n3844), .A2(n2949), .B1(n2169), .B2(n3845), .ZN(n2956)
         );
  NAND2_X1 U2709 ( .A1(n2238), .A2(n3764), .ZN(n2237) );
  OAI22_X1 U2710 ( .A1(n3844), .A2(n2169), .B1(n3868), .B2(n3127), .ZN(n3128)
         );
  INV_X1 U2711 ( .A(n2119), .ZN(n4494) );
  OAI21_X1 U2712 ( .B1(n4486), .B2(n2121), .A(n2120), .ZN(n2119) );
  OAI211_X1 U2713 ( .C1(n2718), .C2(n4537), .A(n2722), .B(n2080), .ZN(U3515)
         );
  MUX2_X2 U2714 ( .A(n2666), .B(n2665), .S(IR_REG_28__SCAN_IN), .Z(n2369) );
  NAND2_X1 U2715 ( .A1(n3591), .A2(n2265), .ZN(n2264) );
  NAND2_X1 U2716 ( .A1(n3779), .A2(n3813), .ZN(n2046) );
  XNOR2_X1 U2717 ( .A(n2384), .B(IR_REG_2__SCAN_IN), .ZN(n4389) );
  AND2_X1 U2718 ( .A1(n2111), .A2(n4492), .ZN(n2047) );
  INV_X1 U2719 ( .A(IR_REG_28__SCAN_IN), .ZN(n2290) );
  AND2_X1 U2720 ( .A1(n2095), .A2(n3211), .ZN(n2048) );
  AND2_X1 U2721 ( .A1(n2205), .A2(n2074), .ZN(n2049) );
  OR2_X1 U2722 ( .A1(n4315), .A2(n3802), .ZN(n2050) );
  NOR2_X1 U2723 ( .A1(n3388), .A2(n3422), .ZN(n2051) );
  NAND2_X1 U2724 ( .A1(n3281), .A2(n3280), .ZN(n3592) );
  OR2_X1 U2725 ( .A1(n4052), .A2(n2102), .ZN(n2052) );
  AND2_X1 U2726 ( .A1(n2100), .A2(n3791), .ZN(n2053) );
  AND2_X1 U2727 ( .A1(n2239), .A2(n2075), .ZN(n2054) );
  INV_X1 U2728 ( .A(n2234), .ZN(n2233) );
  INV_X2 U2729 ( .A(n4537), .ZN(n4539) );
  AND2_X1 U2730 ( .A1(n2862), .A2(n2861), .ZN(n2055) );
  OR3_X1 U2731 ( .A1(n4052), .A2(n2712), .A3(n4235), .ZN(n2056) );
  NOR2_X1 U2732 ( .A1(n2678), .A2(IR_REG_26__SCAN_IN), .ZN(n2303) );
  NAND2_X1 U2733 ( .A1(n3205), .A2(n3204), .ZN(n2057) );
  AND2_X1 U2734 ( .A1(n2046), .A2(n2579), .ZN(n2058) );
  INV_X1 U2735 ( .A(n3018), .ZN(n2222) );
  INV_X1 U2736 ( .A(n2987), .ZN(n2167) );
  AND2_X1 U2737 ( .A1(n2354), .A2(n2353), .ZN(n2059) );
  OAI21_X1 U2738 ( .B1(n3628), .B2(n2229), .A(n2228), .ZN(n3740) );
  NAND2_X1 U2739 ( .A1(n2232), .A2(n3630), .ZN(n3862) );
  AND2_X1 U2740 ( .A1(n2359), .A2(n2358), .ZN(n4388) );
  AND2_X1 U2741 ( .A1(n4249), .A2(n4257), .ZN(n2060) );
  NAND2_X1 U2742 ( .A1(n2256), .A2(n2254), .ZN(n3731) );
  AND3_X1 U2743 ( .A1(n2346), .A2(n2344), .A3(n2347), .ZN(n2061) );
  OR2_X1 U2744 ( .A1(n3595), .A2(n3767), .ZN(n2062) );
  OAI21_X1 U2745 ( .B1(n3570), .B2(n2176), .A(n2533), .ZN(n2175) );
  NOR2_X1 U2746 ( .A1(n4089), .A2(n4248), .ZN(n2063) );
  AND2_X1 U2747 ( .A1(n3290), .A2(n3292), .ZN(n3447) );
  INV_X1 U2748 ( .A(n2264), .ZN(n2263) );
  INV_X1 U2749 ( .A(IR_REG_31__SCAN_IN), .ZN(n2729) );
  AND2_X1 U2750 ( .A1(n2110), .A2(n2111), .ZN(n2064) );
  AND2_X1 U2751 ( .A1(n2108), .A2(n4388), .ZN(n2065) );
  OR2_X1 U2752 ( .A1(n2268), .A2(n2060), .ZN(n2066) );
  OR2_X1 U2753 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2067) );
  INV_X1 U2754 ( .A(n3032), .ZN(n2935) );
  NOR2_X1 U2755 ( .A1(n3522), .A2(n2455), .ZN(n2068) );
  NAND2_X1 U2756 ( .A1(n3907), .A2(n3220), .ZN(n2069) );
  INV_X1 U2757 ( .A(IR_REG_29__SCAN_IN), .ZN(n2209) );
  INV_X1 U2758 ( .A(n4385), .ZN(n2113) );
  INV_X1 U2759 ( .A(n4025), .ZN(n2153) );
  NOR2_X1 U2760 ( .A1(n2399), .A2(n2279), .ZN(n2315) );
  AND2_X1 U2761 ( .A1(n4133), .A2(n2097), .ZN(n2070) );
  INV_X1 U2762 ( .A(n3535), .ZN(n2142) );
  NAND2_X1 U2763 ( .A1(n3592), .A2(n3591), .ZN(n3850) );
  INV_X1 U2764 ( .A(n3525), .ZN(n2163) );
  OR2_X1 U2765 ( .A1(n3851), .A2(n3852), .ZN(n2071) );
  OR2_X1 U2766 ( .A1(n4299), .A2(n4199), .ZN(n2072) );
  OR2_X1 U2767 ( .A1(n3798), .A2(n3797), .ZN(n2073) );
  INV_X1 U2768 ( .A(n3211), .ZN(n3197) );
  AND2_X1 U2769 ( .A1(n2314), .A2(n2313), .ZN(n4156) );
  INV_X1 U2770 ( .A(n4156), .ZN(n2562) );
  INV_X1 U2771 ( .A(n4315), .ZN(n4200) );
  AND3_X1 U2772 ( .A1(n2530), .A2(n2529), .A3(n2528), .ZN(n4315) );
  NAND2_X1 U2773 ( .A1(n2562), .A2(n4276), .ZN(n2074) );
  INV_X1 U2774 ( .A(n2520), .ZN(n2176) );
  OR2_X1 U2775 ( .A1(n4302), .A2(n3791), .ZN(n2520) );
  NAND2_X1 U2776 ( .A1(n2245), .A2(n2247), .ZN(n2075) );
  NAND2_X1 U2777 ( .A1(n3271), .A2(n3270), .ZN(n3278) );
  NOR2_X1 U2778 ( .A1(n4261), .A2(n4070), .ZN(n2076) );
  INV_X1 U2779 ( .A(n3462), .ZN(n2207) );
  INV_X1 U2780 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2115) );
  AND2_X1 U2781 ( .A1(n2048), .A2(n3227), .ZN(n2077) );
  INV_X1 U2782 ( .A(n2563), .ZN(n2206) );
  NOR2_X1 U2783 ( .A1(n2562), .A2(n4276), .ZN(n2563) );
  NOR2_X1 U2784 ( .A1(n3719), .A2(n3621), .ZN(n2078) );
  INV_X1 U2785 ( .A(n2268), .ZN(n2189) );
  INV_X1 U2786 ( .A(IR_REG_0__SCAN_IN), .ZN(n2136) );
  INV_X1 U2787 ( .A(n3896), .ZN(n3764) );
  NAND2_X1 U2788 ( .A1(n2180), .A2(n2269), .ZN(n3300) );
  NAND2_X1 U2789 ( .A1(n3165), .A2(n2273), .ZN(n3207) );
  INV_X1 U2790 ( .A(n3618), .ZN(n3891) );
  INV_X1 U2791 ( .A(n3492), .ZN(n2147) );
  AND2_X1 U2792 ( .A1(n3636), .A2(n3635), .ZN(n2079) );
  AND2_X1 U2793 ( .A1(n2977), .A2(n2975), .ZN(n2974) );
  OR2_X1 U2794 ( .A1(n4539), .A2(n2719), .ZN(n2080) );
  NAND2_X1 U2795 ( .A1(n3060), .A2(n2048), .ZN(n2096) );
  AND2_X1 U2796 ( .A1(n2218), .A2(n2221), .ZN(n2081) );
  INV_X1 U2797 ( .A(n3988), .ZN(n2131) );
  INV_X1 U2798 ( .A(n4198), .ZN(n2171) );
  AND2_X1 U2799 ( .A1(n2131), .A2(n2130), .ZN(n2082) );
  AND2_X1 U2800 ( .A1(n2097), .A2(n4070), .ZN(n2083) );
  AND2_X1 U2801 ( .A1(n2774), .A2(n3563), .ZN(n4438) );
  AND2_X1 U2802 ( .A1(n2758), .A2(n4385), .ZN(n2084) );
  NAND2_X1 U2803 ( .A1(n2872), .A2(n2871), .ZN(n2899) );
  OR2_X1 U2804 ( .A1(n4308), .A2(n2169), .ZN(n2085) );
  INV_X1 U2805 ( .A(n3995), .ZN(n4511) );
  NAND2_X1 U2806 ( .A1(n3734), .A2(n3665), .ZN(n3668) );
  NAND2_X2 U2807 ( .A1(n3731), .A2(n3660), .ZN(n3734) );
  OAI21_X1 U2808 ( .B1(n2935), .B2(n2044), .A(n2086), .ZN(n2896) );
  NAND2_X1 U2809 ( .A1(n3273), .A2(n2087), .ZN(n2086) );
  NAND2_X1 U2810 ( .A1(n2089), .A2(n2088), .ZN(n2945) );
  NAND2_X1 U2811 ( .A1(n3032), .A2(n3273), .ZN(n2088) );
  NAND2_X1 U2812 ( .A1(n2090), .A2(n2248), .ZN(n3267) );
  NAND4_X1 U2813 ( .A1(n3165), .A2(n2273), .A3(n2057), .A4(n3217), .ZN(n2090)
         );
  OR2_X1 U2814 ( .A1(n3164), .A2(n3161), .ZN(n2273) );
  NAND2_X1 U2815 ( .A1(n3164), .A2(n3161), .ZN(n2091) );
  AOI21_X2 U2816 ( .B1(n3763), .B2(n3759), .A(n3760), .ZN(n3829) );
  NAND2_X2 U2817 ( .A1(n2092), .A2(n2261), .ZN(n3763) );
  AND3_X2 U2818 ( .A1(n2217), .A2(n2215), .A3(n2216), .ZN(n3123) );
  NOR2_X2 U2819 ( .A1(n2948), .A2(n2271), .ZN(n3019) );
  INV_X1 U2820 ( .A(n2096), .ZN(n3153) );
  MUX2_X1 U2821 ( .A(n2136), .B(n2101), .S(n2305), .Z(n2879) );
  NAND3_X1 U2822 ( .A1(n4031), .A2(n4225), .A3(n4014), .ZN(n2102) );
  AOI22_X1 U2823 ( .A1(n2791), .A2(n2105), .B1(n2758), .B2(n2104), .ZN(n2107)
         );
  INV_X1 U2824 ( .A(n2107), .ZN(n2805) );
  NAND2_X1 U2825 ( .A1(n4472), .A2(n2112), .ZN(n2110) );
  NAND2_X1 U2826 ( .A1(n4440), .A2(n2129), .ZN(n2125) );
  NOR2_X1 U2827 ( .A1(n4450), .A2(n2322), .ZN(n4449) );
  NAND3_X1 U2828 ( .A1(n2126), .A2(n2127), .A3(n2125), .ZN(n4450) );
  INV_X1 U2829 ( .A(IR_REG_1__SCAN_IN), .ZN(n2135) );
  INV_X1 U2830 ( .A(IR_REG_2__SCAN_IN), .ZN(n2134) );
  NAND3_X1 U2831 ( .A1(n2136), .A2(n2135), .A3(n2134), .ZN(n2348) );
  NOR2_X1 U2832 ( .A1(n2140), .A2(n2208), .ZN(n2139) );
  NAND2_X1 U2833 ( .A1(n3176), .A2(n2145), .ZN(n2143) );
  NAND2_X1 U2834 ( .A1(n4075), .A2(n2152), .ZN(n2151) );
  NAND2_X1 U2835 ( .A1(n3580), .A2(n3579), .ZN(n3578) );
  OAI21_X1 U2836 ( .B1(n3086), .B2(n2164), .A(n2161), .ZN(n3134) );
  OAI21_X1 U2837 ( .B1(n3086), .B2(n2644), .A(n3525), .ZN(n3146) );
  AOI21_X1 U2838 ( .B1(n2644), .B2(n3525), .A(n2166), .ZN(n2165) );
  AOI21_X1 U2839 ( .B1(n3713), .B2(n3409), .A(n2662), .ZN(n2663) );
  NAND2_X1 U2840 ( .A1(n3509), .A2(n3505), .ZN(n2638) );
  NAND2_X1 U2841 ( .A1(n2642), .A2(n3521), .ZN(n3086) );
  NAND2_X1 U2842 ( .A1(n2929), .A2(n3510), .ZN(n2961) );
  OAI21_X1 U2843 ( .B1(n4128), .B2(n2658), .A(n3431), .ZN(n2659) );
  NAND2_X1 U2844 ( .A1(n3960), .A2(n4418), .ZN(n3961) );
  NAND2_X1 U2845 ( .A1(n3334), .A2(n3498), .ZN(n3580) );
  NAND2_X1 U2846 ( .A1(n2961), .A2(n3471), .ZN(n2960) );
  NAND2_X1 U2847 ( .A1(n2651), .A2(n3417), .ZN(n3333) );
  NAND2_X4 U2848 ( .A1(n4377), .A2(n2292), .ZN(n2527) );
  NAND2_X1 U2849 ( .A1(n3571), .A2(n2173), .ZN(n2172) );
  NAND2_X1 U2850 ( .A1(n4092), .A2(n2184), .ZN(n2181) );
  NAND2_X1 U2851 ( .A1(n2181), .A2(n2182), .ZN(n4043) );
  NAND2_X1 U2852 ( .A1(n2192), .A2(n2190), .ZN(n3252) );
  NAND2_X1 U2853 ( .A1(n2392), .A2(n2202), .ZN(n2196) );
  NAND3_X1 U2854 ( .A1(n2197), .A2(n2196), .A3(n2068), .ZN(n3140) );
  OAI22_X1 U2855 ( .A1(n4147), .A2(n2204), .B1(n2563), .B2(n2049), .ZN(n4122)
         );
  NAND2_X1 U2856 ( .A1(n4377), .A2(n4378), .ZN(n2378) );
  NAND3_X1 U2857 ( .A1(n2402), .A2(n2211), .A3(n2260), .ZN(n2676) );
  NAND3_X1 U2858 ( .A1(n2402), .A2(n2211), .A3(n2210), .ZN(n2678) );
  NAND2_X1 U2859 ( .A1(n2866), .A2(n2212), .ZN(n2898) );
  XNOR2_X1 U2860 ( .A(n2863), .B(n3613), .ZN(n2212) );
  NAND2_X1 U2861 ( .A1(n2213), .A2(n3605), .ZN(n3617) );
  NAND3_X1 U2862 ( .A1(n2213), .A2(n3605), .A3(n2078), .ZN(n3785) );
  INV_X1 U2863 ( .A(n3109), .ZN(n2214) );
  NAND2_X1 U2864 ( .A1(n2225), .A2(n2226), .ZN(n3643) );
  NAND2_X1 U2865 ( .A1(n3628), .A2(n2228), .ZN(n2225) );
  NAND2_X1 U2866 ( .A1(n3628), .A2(n3627), .ZN(n3796) );
  NAND2_X1 U2867 ( .A1(n2073), .A2(n3627), .ZN(n2234) );
  NAND2_X1 U2868 ( .A1(n3681), .A2(n2236), .ZN(n2235) );
  OAI211_X1 U2869 ( .C1(n3681), .C2(n2237), .A(n2235), .B(n3705), .ZN(U3217)
         );
  NAND2_X1 U2870 ( .A1(n3681), .A2(n3874), .ZN(n3691) );
  INV_X1 U2871 ( .A(n3699), .ZN(n2247) );
  NAND3_X1 U2872 ( .A1(n3165), .A2(n2273), .A3(n2057), .ZN(n2249) );
  NAND2_X1 U2873 ( .A1(n3818), .A2(n3822), .ZN(n3750) );
  NOR2_X1 U2874 ( .A1(n3655), .A2(n2259), .ZN(n2258) );
  INV_X1 U2875 ( .A(n3822), .ZN(n2259) );
  NAND2_X1 U2876 ( .A1(n2299), .A2(n2290), .ZN(n2668) );
  OR2_X1 U2877 ( .A1(n2379), .A2(n2360), .ZN(n2367) );
  OR2_X1 U2878 ( .A1(n2377), .A2(n2376), .ZN(n2383) );
  OR2_X1 U2879 ( .A1(n2527), .A2(n2750), .ZN(n2380) );
  AOI21_X2 U2880 ( .B1(n3111), .B2(n3110), .A(n3123), .ZN(n3164) );
  INV_X1 U2881 ( .A(n4377), .ZN(n2293) );
  AND2_X1 U2882 ( .A1(n2356), .A2(n2277), .ZN(n2267) );
  AND2_X1 U2883 ( .A1(n4258), .A2(n2711), .ZN(n2268) );
  OR2_X1 U2884 ( .A1(n3904), .A2(n3596), .ZN(n2269) );
  OR2_X1 U2885 ( .A1(n4154), .A2(n2710), .ZN(n2270) );
  AND2_X1 U2886 ( .A1(n2947), .A2(n2946), .ZN(n2271) );
  AND2_X1 U2887 ( .A1(n3665), .A2(n3666), .ZN(n2272) );
  NAND2_X1 U2888 ( .A1(n3734), .A2(n2272), .ZN(n3808) );
  INV_X1 U2889 ( .A(n4276), .ZN(n4142) );
  NOR2_X1 U2890 ( .A1(n3402), .A2(n2306), .ZN(n4276) );
  NAND2_X1 U2891 ( .A1(n4545), .A2(n4317), .ZN(n4307) );
  INV_X1 U2892 ( .A(n4369), .ZN(n2720) );
  AND2_X1 U2893 ( .A1(n3785), .A2(n3784), .ZN(n2274) );
  INV_X1 U2894 ( .A(IR_REG_4__SCAN_IN), .ZN(n2277) );
  OR2_X1 U2895 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  NAND2_X1 U2896 ( .A1(n2928), .A2(n3011), .ZN(n3509) );
  INV_X1 U2897 ( .A(n3106), .ZN(n3107) );
  NAND2_X1 U2898 ( .A1(n3641), .A2(n3640), .ZN(n3642) );
  AND2_X1 U2899 ( .A1(n2494), .A2(REG3_REG_16__SCAN_IN), .ZN(n2510) );
  OR2_X1 U2900 ( .A1(n4137), .A2(n4117), .ZN(n4096) );
  NAND2_X1 U2901 ( .A1(n3519), .A2(n3515), .ZN(n2977) );
  OR2_X1 U2902 ( .A1(n3615), .A2(n3614), .ZN(n3720) );
  AND2_X1 U2903 ( .A1(n3602), .A2(n3601), .ZN(n3760) );
  NOR2_X1 U2904 ( .A1(n3108), .A2(n3107), .ZN(n3109) );
  AND2_X1 U2905 ( .A1(n2543), .A2(REG3_REG_20__SCAN_IN), .ZN(n2307) );
  INV_X2 U2906 ( .A(n2055), .ZN(n3695) );
  AND2_X1 U2907 ( .A1(n3621), .A2(n3720), .ZN(n3616) );
  NAND2_X1 U2908 ( .A1(n2510), .A2(REG3_REG_17__SCAN_IN), .ZN(n2535) );
  NOR2_X1 U2909 ( .A1(n2407), .A2(n2792), .ZN(n2417) );
  OR2_X1 U2910 ( .A1(n4281), .A2(n4117), .ZN(n2571) );
  INV_X1 U2911 ( .A(n2861), .ZN(n2888) );
  INV_X1 U2912 ( .A(n3802), .ZN(n4297) );
  INV_X1 U2913 ( .A(n4520), .ZN(n3974) );
  INV_X1 U2914 ( .A(n2977), .ZN(n3473) );
  AND2_X1 U2915 ( .A1(n2417), .A2(REG3_REG_7__SCAN_IN), .ZN(n2428) );
  INV_X1 U2916 ( .A(n3220), .ZN(n3227) );
  INV_X1 U2917 ( .A(n3075), .ZN(n3118) );
  INV_X1 U2918 ( .A(n3844), .ZN(n3888) );
  OR2_X1 U2919 ( .A1(n2737), .A2(D_REG_1__SCAN_IN), .ZN(n2883) );
  INV_X1 U2920 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4692) );
  INV_X1 U2921 ( .A(n3899), .ZN(n4227) );
  INV_X1 U2922 ( .A(n4311), .ZN(n3791) );
  OR2_X1 U2923 ( .A1(n2737), .A2(D_REG_0__SCAN_IN), .ZN(n2708) );
  INV_X1 U2924 ( .A(n4248), .ZN(n4070) );
  INV_X1 U2925 ( .A(n4185), .ZN(n2710) );
  INV_X1 U2926 ( .A(n4204), .ZN(n4182) );
  NAND2_X1 U2927 ( .A1(n2276), .A2(REG3_REG_23__SCAN_IN), .ZN(n2580) );
  AND2_X1 U2928 ( .A1(n2428), .A2(REG3_REG_8__SCAN_IN), .ZN(n2440) );
  AND2_X1 U2929 ( .A1(n2578), .A2(n2577), .ZN(n4085) );
  AND4_X1 U2930 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n3768)
         );
  INV_X1 U2931 ( .A(IR_REG_8__SCAN_IN), .ZN(n2437) );
  OR2_X1 U2932 ( .A1(n2670), .A2(n2669), .ZN(n2853) );
  INV_X1 U2933 ( .A(n4226), .ZN(n4310) );
  INV_X1 U2934 ( .A(n4187), .ZN(n4501) );
  INV_X1 U2935 ( .A(n4216), .ZN(n4132) );
  INV_X1 U2936 ( .A(n4141), .ZN(n4082) );
  INV_X1 U2937 ( .A(n4307), .ZN(n2714) );
  NAND2_X1 U2938 ( .A1(n2708), .A2(n2707), .ZN(n2884) );
  INV_X1 U2939 ( .A(n4018), .ZN(n2721) );
  AND2_X1 U2940 ( .A1(n2980), .A2(n2979), .ZN(n4530) );
  INV_X1 U2941 ( .A(n2884), .ZN(n2838) );
  INV_X1 U2942 ( .A(n2637), .ZN(n2726) );
  AND2_X1 U2943 ( .A1(n2481), .A2(n2490), .ZN(n3973) );
  AND2_X1 U2944 ( .A1(n2742), .A2(n2735), .ZN(n4489) );
  INV_X1 U2945 ( .A(n3893), .ZN(n3811) );
  OR2_X1 U2946 ( .A1(n2875), .A2(n2852), .ZN(n3896) );
  INV_X1 U2947 ( .A(n4238), .ZN(n4036) );
  NAND2_X1 U2948 ( .A1(n2560), .A2(n2559), .ZN(n4278) );
  INV_X1 U2949 ( .A(n3768), .ZN(n3903) );
  INV_X1 U2950 ( .A(n4515), .ZN(n4435) );
  INV_X1 U2951 ( .A(n4438), .ZN(n4485) );
  NAND2_X1 U2952 ( .A1(n4191), .A2(n2994), .ZN(n4216) );
  NAND2_X1 U2953 ( .A1(n2721), .A2(n2714), .ZN(n2715) );
  OR2_X1 U2954 ( .A1(n2717), .A2(n2884), .ZN(n4543) );
  NAND2_X1 U2955 ( .A1(n4539), .A2(n4317), .ZN(n4369) );
  AND3_X1 U2956 ( .A1(n4536), .A2(n4535), .A3(n4534), .ZN(n4544) );
  OR2_X1 U2957 ( .A1(n2717), .A2(n2838), .ZN(n4537) );
  INV_X1 U2958 ( .A(n2689), .ZN(n3585) );
  INV_X1 U2959 ( .A(n3972), .ZN(n4514) );
  INV_X1 U2960 ( .A(n2787), .ZN(n4386) );
  INV_X1 U2961 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2709) );
  INV_X1 U2962 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2330) );
  INV_X1 U2963 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2534) );
  INV_X1 U2964 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4578) );
  INV_X1 U2965 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3843) );
  INV_X1 U2966 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4690) );
  XNOR2_X1 U2967 ( .A(n2590), .B(REG3_REG_25__SCAN_IN), .ZN(n4067) );
  INV_X1 U2968 ( .A(n2348), .ZN(n2278) );
  NAND2_X1 U2969 ( .A1(n2278), .A2(n2267), .ZN(n2399) );
  XNOR2_X2 U2970 ( .A(n2291), .B(IR_REG_30__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U2971 ( .A1(n4067), .A2(n2362), .ZN(n2298) );
  INV_X1 U2972 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4255) );
  BUF_X4 U2973 ( .A(n2379), .Z(n3407) );
  NAND2_X1 U2974 ( .A1(n2337), .A2(REG2_REG_25__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2975 ( .A1(n3404), .A2(REG0_REG_25__SCAN_IN), .ZN(n2294) );
  OAI211_X1 U2976 ( .C1(n4255), .C2(n3407), .A(n2295), .B(n2294), .ZN(n2296)
         );
  INV_X1 U2977 ( .A(n2296), .ZN(n2297) );
  INV_X1 U2978 ( .A(n4089), .ZN(n4261) );
  NAND2_X1 U2979 ( .A1(n2300), .A2(n2729), .ZN(n2301) );
  NAND2_X1 U2980 ( .A1(n2302), .A2(n2301), .ZN(n2666) );
  INV_X1 U2981 ( .A(n2303), .ZN(n2685) );
  INV_X1 U2982 ( .A(DATAI_25_), .ZN(n4583) );
  NOR2_X1 U2983 ( .A1(n3402), .A2(n4583), .ZN(n4248) );
  INV_X1 U2984 ( .A(DATAI_21_), .ZN(n2306) );
  INV_X1 U2985 ( .A(n2307), .ZN(n2555) );
  INV_X1 U2986 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2987 ( .A1(n2555), .A2(n2308), .ZN(n2309) );
  NAND2_X1 U2988 ( .A1(n2564), .A2(n2309), .ZN(n3754) );
  OR2_X1 U2989 ( .A1(n3754), .A2(n2619), .ZN(n2314) );
  INV_X1 U2990 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U2991 ( .A1(n3404), .A2(REG0_REG_21__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U2992 ( .A1(n2337), .A2(REG2_REG_21__SCAN_IN), .ZN(n2310) );
  OAI211_X1 U2993 ( .C1(n3407), .C2(n4284), .A(n2311), .B(n2310), .ZN(n2312)
         );
  INV_X1 U2994 ( .A(n2312), .ZN(n2313) );
  INV_X1 U2995 ( .A(IR_REG_9__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2996 ( .A1(n2315), .A2(n2316), .ZN(n2477) );
  INV_X1 U2997 ( .A(n2317), .ZN(n2318) );
  NOR2_X1 U2998 ( .A1(n2327), .A2(IR_REG_13__SCAN_IN), .ZN(n2503) );
  OR2_X1 U2999 ( .A1(n2503), .A2(n2729), .ZN(n2319) );
  XNOR2_X1 U3000 ( .A(n2319), .B(IR_REG_14__SCAN_IN), .ZN(n3988) );
  MUX2_X1 U3001 ( .A(DATAI_14_), .B(n3988), .S(n2369), .Z(n3609) );
  NAND2_X1 U3002 ( .A1(n3404), .A2(REG0_REG_14__SCAN_IN), .ZN(n2326) );
  INV_X1 U3003 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3364) );
  OR2_X1 U3004 ( .A1(n3407), .A2(n3364), .ZN(n2325) );
  INV_X1 U3005 ( .A(n2320), .ZN(n2496) );
  NAND2_X1 U3006 ( .A1(n2332), .A2(n4692), .ZN(n2321) );
  NAND2_X1 U3007 ( .A1(n2496), .A2(n2321), .ZN(n3730) );
  OR2_X1 U3008 ( .A1(n2619), .A2(n3730), .ZN(n2324) );
  INV_X1 U3009 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2322) );
  OR2_X1 U3010 ( .A1(n2527), .A2(n2322), .ZN(n2323) );
  INV_X1 U3011 ( .A(DATAI_13_), .ZN(n2329) );
  NAND2_X1 U3012 ( .A1(n2327), .A2(IR_REG_31__SCAN_IN), .ZN(n2328) );
  XNOR2_X1 U3013 ( .A(n2328), .B(IR_REG_13__SCAN_IN), .ZN(n3972) );
  MUX2_X1 U3014 ( .A(n2329), .B(n4514), .S(n3402), .Z(n3835) );
  INV_X1 U3015 ( .A(n3835), .ZN(n3295) );
  NAND2_X1 U3016 ( .A1(n3404), .A2(REG0_REG_13__SCAN_IN), .ZN(n2336) );
  INV_X1 U3017 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4437) );
  OR2_X1 U3018 ( .A1(n2527), .A2(n4437), .ZN(n2335) );
  NAND2_X1 U3019 ( .A1(n2485), .A2(n2330), .ZN(n2331) );
  NAND2_X1 U3020 ( .A1(n2332), .A2(n2331), .ZN(n3303) );
  OR2_X1 U3021 ( .A1(n2619), .A2(n3303), .ZN(n2334) );
  INV_X1 U3022 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3372) );
  OR2_X1 U3023 ( .A1(n3407), .A2(n3372), .ZN(n2333) );
  NAND2_X1 U3024 ( .A1(n2337), .A2(REG2_REG_4__SCAN_IN), .ZN(n2347) );
  INV_X1 U3025 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2338) );
  OR2_X1 U3026 ( .A1(n2377), .A2(n2338), .ZN(n2346) );
  INV_X1 U3027 ( .A(n2393), .ZN(n2342) );
  INV_X1 U3028 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2340) );
  INV_X1 U3029 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U3030 ( .A1(n2340), .A2(n2339), .ZN(n2341) );
  NAND2_X1 U3031 ( .A1(n2342), .A2(n2341), .ZN(n3028) );
  INV_X1 U3032 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2343) );
  OR2_X1 U3033 ( .A1(n2379), .A2(n2343), .ZN(n2344) );
  NAND2_X1 U3034 ( .A1(n2348), .A2(IR_REG_31__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U3035 ( .A1(n2357), .A2(n2356), .ZN(n2359) );
  NAND2_X1 U3036 ( .A1(n2359), .A2(IR_REG_31__SCAN_IN), .ZN(n2349) );
  XNOR2_X1 U3037 ( .A(n2349), .B(IR_REG_4__SCAN_IN), .ZN(n4387) );
  MUX2_X1 U3038 ( .A(DATAI_4_), .B(n4387), .S(n2369), .Z(n2987) );
  NAND2_X1 U3039 ( .A1(n3912), .A2(n2987), .ZN(n2388) );
  INV_X1 U3040 ( .A(n2388), .ZN(n2391) );
  OR2_X1 U3041 ( .A1(n2378), .A2(REG3_REG_3__SCAN_IN), .ZN(n2354) );
  INV_X1 U3042 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2350) );
  INV_X1 U3043 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3945) );
  OR2_X1 U3044 ( .A1(n2527), .A2(n3945), .ZN(n2351) );
  INV_X1 U3045 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2967) );
  OR2_X1 U3046 ( .A1(n3407), .A2(n2967), .ZN(n2355) );
  OR2_X1 U3047 ( .A1(n2357), .A2(n2356), .ZN(n2358) );
  MUX2_X1 U3048 ( .A(DATAI_3_), .B(n4388), .S(n2369), .Z(n2963) );
  NAND2_X1 U3049 ( .A1(n2640), .A2(n3001), .ZN(n2975) );
  INV_X1 U3050 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U3051 ( .A1(n2361), .A2(REG2_REG_1__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U3052 ( .A1(n2362), .A2(REG3_REG_1__SCAN_IN), .ZN(n2365) );
  INV_X1 U3053 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U3054 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2368)
         );
  MUX2_X1 U3055 ( .A(DATAI_1_), .B(n4390), .S(n2042), .Z(n3011) );
  INV_X1 U3056 ( .A(n2928), .ZN(n3914) );
  INV_X1 U3057 ( .A(n3011), .ZN(n2859) );
  INV_X1 U3058 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2370) );
  OR2_X1 U3059 ( .A1(n2377), .A2(n2370), .ZN(n2371) );
  AND2_X1 U3060 ( .A1(n2372), .A2(n2371), .ZN(n2375) );
  INV_X1 U3061 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2743) );
  OR2_X1 U3062 ( .A1(n2527), .A2(n2743), .ZN(n2374) );
  INV_X1 U3063 ( .A(n2379), .ZN(n2537) );
  NAND2_X1 U3064 ( .A1(n2537), .A2(REG1_REG_0__SCAN_IN), .ZN(n2373) );
  AND2_X1 U3065 ( .A1(n2815), .A2(n2916), .ZN(n2908) );
  NAND2_X1 U3066 ( .A1(n2638), .A2(n2908), .ZN(n2907) );
  INV_X1 U3067 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2376) );
  INV_X1 U3068 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3925) );
  INV_X1 U3069 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2762) );
  OR2_X1 U3070 ( .A1(n2379), .A2(n2762), .ZN(n2381) );
  INV_X1 U3071 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2750) );
  AND4_X2 U3072 ( .A1(n2383), .A2(n2382), .A3(n2381), .A4(n2380), .ZN(n2949)
         );
  MUX2_X1 U3073 ( .A(DATAI_2_), .B(n4389), .S(n2369), .Z(n3032) );
  NAND2_X1 U3074 ( .A1(n2087), .A2(n2935), .ZN(n3503) );
  NAND2_X1 U3075 ( .A1(n2949), .A2(n3032), .ZN(n3510) );
  NAND2_X1 U3076 ( .A1(n3503), .A2(n3510), .ZN(n2639) );
  NAND2_X1 U3077 ( .A1(n3914), .A2(n3011), .ZN(n2923) );
  AND2_X1 U3078 ( .A1(n2639), .A2(n2923), .ZN(n2385) );
  NAND2_X1 U3079 ( .A1(n2907), .A2(n2385), .ZN(n2387) );
  NAND2_X1 U3080 ( .A1(n2949), .A2(n2935), .ZN(n2386) );
  NAND2_X1 U3081 ( .A1(n2387), .A2(n2386), .ZN(n2959) );
  NAND2_X1 U3082 ( .A1(n3913), .A2(n2963), .ZN(n2973) );
  AND2_X1 U3083 ( .A1(n2973), .A2(n2388), .ZN(n2389) );
  NAND2_X1 U3084 ( .A1(n2959), .A2(n2389), .ZN(n2390) );
  OAI21_X1 U3085 ( .B1(n2391), .B2(n2974), .A(n2390), .ZN(n2392) );
  INV_X1 U3086 ( .A(n2392), .ZN(n3052) );
  NAND2_X1 U3087 ( .A1(n3404), .A2(REG0_REG_5__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3088 ( .A1(n3407), .A2(n2115), .ZN(n2397) );
  OAI21_X1 U3089 ( .B1(n2393), .B2(REG3_REG_5__SCAN_IN), .A(n2407), .ZN(n3132)
         );
  OR2_X1 U3090 ( .A1(n2619), .A2(n3132), .ZN(n2396) );
  INV_X1 U3091 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2394) );
  OR2_X1 U3092 ( .A1(n2527), .A2(n2394), .ZN(n2395) );
  INV_X1 U3093 ( .A(DATAI_5_), .ZN(n4704) );
  NAND2_X1 U3094 ( .A1(n2399), .A2(IR_REG_31__SCAN_IN), .ZN(n2400) );
  MUX2_X1 U3095 ( .A(n2400), .B(IR_REG_31__SCAN_IN), .S(n2401), .Z(n2403) );
  INV_X1 U3096 ( .A(n2399), .ZN(n2402) );
  NAND2_X1 U3097 ( .A1(n2402), .A2(n2401), .ZN(n2424) );
  NAND2_X1 U3098 ( .A1(n2403), .A2(n2424), .ZN(n2787) );
  MUX2_X1 U3099 ( .A(n4704), .B(n2787), .S(n2369), .Z(n3127) );
  NAND2_X1 U3100 ( .A1(n3103), .A2(n3127), .ZN(n2404) );
  INV_X1 U3101 ( .A(n3103), .ZN(n3911) );
  NAND2_X1 U3102 ( .A1(n3911), .A2(n3100), .ZN(n2405) );
  NAND2_X1 U3103 ( .A1(n3404), .A2(REG0_REG_6__SCAN_IN), .ZN(n2413) );
  INV_X1 U3104 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3105 ( .A1(n2527), .A2(n2406), .ZN(n2412) );
  AND2_X1 U3106 ( .A1(n2407), .A2(n2792), .ZN(n2408) );
  OR2_X1 U3107 ( .A1(n2408), .A2(n2417), .ZN(n3076) );
  OR2_X1 U3108 ( .A1(n2619), .A2(n3076), .ZN(n2411) );
  INV_X1 U3109 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2409) );
  OR2_X1 U3110 ( .A1(n3407), .A2(n2409), .ZN(n2410) );
  NAND4_X1 U3111 ( .A1(n2413), .A2(n2412), .A3(n2411), .A4(n2410), .ZN(n3910)
         );
  NAND2_X1 U3112 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2414) );
  XNOR2_X1 U3113 ( .A(n2414), .B(IR_REG_6__SCAN_IN), .ZN(n4385) );
  MUX2_X1 U3114 ( .A(DATAI_6_), .B(n4385), .S(n2369), .Z(n3075) );
  AND2_X1 U3115 ( .A1(n3910), .A2(n3075), .ZN(n2415) );
  NAND2_X1 U3116 ( .A1(n3404), .A2(REG0_REG_7__SCAN_IN), .ZN(n2423) );
  INV_X1 U3117 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2416) );
  OR2_X1 U3118 ( .A1(n2527), .A2(n2416), .ZN(n2422) );
  NOR2_X1 U3119 ( .A1(n2417), .A2(REG3_REG_7__SCAN_IN), .ZN(n2418) );
  OR2_X1 U3120 ( .A1(n2428), .A2(n2418), .ZN(n3167) );
  OR2_X1 U3121 ( .A1(n2619), .A2(n3167), .ZN(n2421) );
  INV_X1 U3122 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2419) );
  OR2_X1 U3123 ( .A1(n3407), .A2(n2419), .ZN(n2420) );
  INV_X1 U3124 ( .A(n2424), .ZN(n2426) );
  NAND2_X1 U3125 ( .A1(n2426), .A2(n2425), .ZN(n2427) );
  NAND2_X1 U3126 ( .A1(n2427), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  XNOR2_X1 U3127 ( .A(n2435), .B(IR_REG_7__SCAN_IN), .ZN(n4384) );
  MUX2_X1 U3128 ( .A(DATAI_7_), .B(n4384), .S(n2369), .Z(n3091) );
  NAND2_X1 U3129 ( .A1(n3210), .A2(n3091), .ZN(n2643) );
  INV_X1 U3130 ( .A(n3091), .ZN(n3171) );
  NAND2_X1 U3131 ( .A1(n3909), .A2(n3171), .ZN(n3525) );
  NAND2_X1 U3132 ( .A1(n3404), .A2(REG0_REG_8__SCAN_IN), .ZN(n2433) );
  INV_X1 U3133 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3978) );
  OR2_X1 U3134 ( .A1(n3407), .A2(n3978), .ZN(n2432) );
  NOR2_X1 U3135 ( .A1(n2428), .A2(REG3_REG_8__SCAN_IN), .ZN(n2429) );
  OR2_X1 U3136 ( .A1(n2440), .A2(n2429), .ZN(n4497) );
  OR2_X1 U3137 ( .A1(n2619), .A2(n4497), .ZN(n2431) );
  INV_X1 U3138 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4498) );
  OR2_X1 U3139 ( .A1(n2527), .A2(n4498), .ZN(n2430) );
  INV_X1 U3140 ( .A(DATAI_8_), .ZN(n2439) );
  NAND2_X1 U3141 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3142 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  XNOR2_X1 U3143 ( .A(n2438), .B(n2437), .ZN(n4382) );
  MUX2_X1 U3144 ( .A(n2439), .B(n4382), .S(n2369), .Z(n3211) );
  AND2_X1 U3145 ( .A1(n3196), .A2(n3211), .ZN(n2455) );
  NAND2_X1 U3146 ( .A1(n3404), .A2(REG0_REG_9__SCAN_IN), .ZN(n2449) );
  INV_X1 U3147 ( .A(n2440), .ZN(n2442) );
  INV_X1 U31480 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U31490 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  NAND2_X1 U3150 ( .A1(n2461), .A2(n2443), .ZN(n3224) );
  OR2_X1 U3151 ( .A1(n2619), .A2(n3224), .ZN(n2448) );
  INV_X1 U3152 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2444) );
  OR2_X1 U3153 ( .A1(n3407), .A2(n2444), .ZN(n2447) );
  INV_X1 U3154 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2445) );
  OR2_X1 U3155 ( .A1(n2527), .A2(n2445), .ZN(n2446) );
  NAND4_X1 U3156 ( .A1(n2449), .A2(n2448), .A3(n2447), .A4(n2446), .ZN(n3907)
         );
  NOR2_X1 U3157 ( .A1(n2315), .A2(n2729), .ZN(n2450) );
  MUX2_X1 U3158 ( .A(n2729), .B(n2450), .S(IR_REG_9__SCAN_IN), .Z(n2452) );
  INV_X1 U3159 ( .A(n2477), .ZN(n2451) );
  MUX2_X1 U3160 ( .A(DATAI_9_), .B(n3974), .S(n2369), .Z(n3220) );
  NAND2_X1 U3161 ( .A1(n3909), .A2(n3091), .ZN(n3144) );
  NAND2_X1 U3162 ( .A1(n3908), .A2(n3197), .ZN(n2453) );
  AND2_X1 U3163 ( .A1(n3144), .A2(n2453), .ZN(n2454) );
  OR2_X1 U3164 ( .A1(n2455), .A2(n2454), .ZN(n3139) );
  AND2_X1 U3165 ( .A1(n2069), .A2(n3139), .ZN(n2456) );
  NAND2_X1 U3166 ( .A1(n3140), .A2(n2456), .ZN(n2458) );
  NAND2_X1 U3167 ( .A1(n3283), .A2(n3227), .ZN(n2457) );
  NAND2_X1 U3168 ( .A1(n3404), .A2(REG0_REG_10__SCAN_IN), .ZN(n2467) );
  INV_X1 U3169 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2459) );
  OR2_X1 U3170 ( .A1(n3407), .A2(n2459), .ZN(n2466) );
  INV_X1 U3171 ( .A(n2460), .ZN(n2471) );
  INV_X1 U3172 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U3173 ( .A1(n2461), .A2(n4705), .ZN(n2462) );
  NAND2_X1 U3174 ( .A1(n2471), .A2(n2462), .ZN(n3289) );
  OR2_X1 U3175 ( .A1(n2619), .A2(n3289), .ZN(n2465) );
  INV_X1 U3176 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2463) );
  OR2_X1 U3177 ( .A1(n2527), .A2(n2463), .ZN(n2464) );
  NAND2_X1 U3178 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  XNOR2_X1 U3179 ( .A(n2468), .B(IR_REG_10__SCAN_IN), .ZN(n3981) );
  MUX2_X1 U3180 ( .A(DATAI_10_), .B(n3981), .S(n2369), .Z(n3274) );
  NOR2_X1 U3181 ( .A1(n3906), .A2(n3274), .ZN(n2469) );
  NAND2_X1 U3182 ( .A1(n3404), .A2(REG0_REG_11__SCAN_IN), .ZN(n2476) );
  INV_X1 U3183 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3327) );
  OR2_X1 U3184 ( .A1(n3407), .A2(n3327), .ZN(n2475) );
  INV_X1 U3185 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3186 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U3187 ( .A1(n2483), .A2(n2472), .ZN(n3854) );
  OR2_X1 U3188 ( .A1(n2619), .A2(n3854), .ZN(n2474) );
  INV_X1 U3189 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3259) );
  OR2_X1 U3190 ( .A1(n2527), .A2(n3259), .ZN(n2473) );
  OR2_X1 U3191 ( .A1(n2477), .A2(IR_REG_10__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3192 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  INV_X1 U3193 ( .A(IR_REG_11__SCAN_IN), .ZN(n2479) );
  OR2_X1 U3194 ( .A1(n2480), .A2(n2479), .ZN(n2481) );
  NAND2_X1 U3195 ( .A1(n2480), .A2(n2479), .ZN(n2490) );
  MUX2_X1 U3196 ( .A(DATAI_11_), .B(n3973), .S(n2369), .Z(n3255) );
  NAND2_X1 U3197 ( .A1(n3766), .A2(n3255), .ZN(n3290) );
  INV_X1 U3198 ( .A(n3766), .ZN(n3905) );
  NAND2_X1 U3199 ( .A1(n3905), .A2(n3857), .ZN(n3292) );
  NAND2_X1 U3200 ( .A1(n3766), .A2(n3857), .ZN(n2482) );
  NAND2_X1 U3201 ( .A1(n3252), .A2(n2482), .ZN(n3308) );
  NAND2_X1 U3202 ( .A1(n3404), .A2(REG0_REG_12__SCAN_IN), .ZN(n2489) );
  INV_X1 U3203 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3314) );
  OR2_X1 U3204 ( .A1(n2527), .A2(n3314), .ZN(n2488) );
  NAND2_X1 U3205 ( .A1(n2483), .A2(n4547), .ZN(n2484) );
  NAND2_X1 U3206 ( .A1(n2485), .A2(n2484), .ZN(n3773) );
  OR2_X1 U3207 ( .A1(n2619), .A2(n3773), .ZN(n2487) );
  INV_X1 U3208 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3356) );
  OR2_X1 U3209 ( .A1(n3407), .A2(n3356), .ZN(n2486) );
  INV_X1 U32100 ( .A(DATAI_12_), .ZN(n2492) );
  NAND2_X1 U32110 ( .A1(n2490), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  XNOR2_X1 U32120 ( .A(n2491), .B(IR_REG_12__SCAN_IN), .ZN(n4515) );
  MUX2_X1 U32130 ( .A(n2492), .B(n4435), .S(n2042), .Z(n3767) );
  NAND2_X1 U32140 ( .A1(n3608), .A2(n3609), .ZN(n3417) );
  NAND2_X1 U32150 ( .A1(n3902), .A2(n3724), .ZN(n3499) );
  NAND2_X1 U32160 ( .A1(n3417), .A2(n3499), .ZN(n3242) );
  NAND2_X1 U32170 ( .A1(n3243), .A2(n3242), .ZN(n3241) );
  NAND2_X1 U32180 ( .A1(n3404), .A2(REG0_REG_15__SCAN_IN), .ZN(n2501) );
  INV_X1 U32190 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2493) );
  OR2_X1 U32200 ( .A1(n2527), .A2(n2493), .ZN(n2500) );
  INV_X1 U32210 ( .A(n2494), .ZN(n2511) );
  INV_X1 U32220 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U32230 ( .A1(n2496), .A2(n2495), .ZN(n2497) );
  NAND2_X1 U32240 ( .A1(n2511), .A2(n2497), .ZN(n3339) );
  OR2_X1 U32250 ( .A1(n2619), .A2(n3339), .ZN(n2499) );
  INV_X1 U32260 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3382) );
  OR2_X1 U32270 ( .A1(n3407), .A2(n3382), .ZN(n2498) );
  INV_X1 U32280 ( .A(IR_REG_14__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U32290 ( .A1(n2503), .A2(n2502), .ZN(n2504) );
  NAND2_X1 U32300 ( .A1(n2504), .A2(IR_REG_31__SCAN_IN), .ZN(n2506) );
  INV_X1 U32310 ( .A(IR_REG_15__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32320 ( .A1(n2506), .A2(n2505), .ZN(n2518) );
  OR2_X1 U32330 ( .A1(n2506), .A2(n2505), .ZN(n2507) );
  MUX2_X1 U32340 ( .A(DATAI_15_), .B(n3971), .S(n3402), .Z(n3618) );
  NAND2_X1 U32350 ( .A1(n3901), .A2(n3618), .ZN(n2508) );
  NAND2_X1 U32360 ( .A1(n3404), .A2(REG0_REG_16__SCAN_IN), .ZN(n2517) );
  INV_X1 U32370 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2509) );
  OR2_X1 U32380 ( .A1(n2527), .A2(n2509), .ZN(n2516) );
  INV_X1 U32390 ( .A(n2510), .ZN(n2524) );
  INV_X1 U32400 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U32410 ( .A1(n2511), .A2(n4558), .ZN(n2512) );
  NAND2_X1 U32420 ( .A1(n2524), .A2(n2512), .ZN(n3575) );
  OR2_X1 U32430 ( .A1(n3575), .A2(n2619), .ZN(n2515) );
  INV_X1 U32440 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2513) );
  OR2_X1 U32450 ( .A1(n3407), .A2(n2513), .ZN(n2514) );
  NAND2_X1 U32460 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  XNOR2_X1 U32470 ( .A(n2519), .B(IR_REG_16__SCAN_IN), .ZN(n3992) );
  MUX2_X1 U32480 ( .A(DATAI_16_), .B(n3992), .S(n3402), .Z(n4311) );
  NAND2_X1 U32490 ( .A1(n4302), .A2(n4311), .ZN(n3426) );
  NAND2_X1 U32500 ( .A1(n3900), .A2(n3791), .ZN(n3500) );
  NAND2_X1 U32510 ( .A1(n3426), .A2(n3500), .ZN(n3570) );
  INV_X1 U32520 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4373) );
  OR2_X1 U32530 ( .A1(n2377), .A2(n4373), .ZN(n2522) );
  INV_X1 U32540 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4305) );
  OR2_X1 U32550 ( .A1(n3407), .A2(n4305), .ZN(n2521) );
  AND2_X1 U32560 ( .A1(n2522), .A2(n2521), .ZN(n2530) );
  INV_X1 U32570 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32580 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  NAND2_X1 U32590 ( .A1(n2535), .A2(n2525), .ZN(n3394) );
  OR2_X1 U32600 ( .A1(n3394), .A2(n2619), .ZN(n2529) );
  INV_X1 U32610 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2526) );
  OR2_X1 U32620 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  INV_X1 U32630 ( .A(DATAI_17_), .ZN(n2532) );
  OR2_X1 U32640 ( .A1(n2541), .A2(n2729), .ZN(n2531) );
  XNOR2_X1 U32650 ( .A(n2531), .B(IR_REG_17__SCAN_IN), .ZN(n3995) );
  MUX2_X1 U32660 ( .A(n2532), .B(n4511), .S(n3402), .Z(n3802) );
  NAND2_X1 U32670 ( .A1(n4315), .A2(n3802), .ZN(n2533) );
  NAND2_X1 U32680 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  NAND2_X1 U32690 ( .A1(n2544), .A2(n2536), .ZN(n3865) );
  AOI22_X1 U32700 ( .A1(n2537), .A2(REG1_REG_18__SCAN_IN), .B1(n3404), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32710 ( .A1(n2337), .A2(REG2_REG_18__SCAN_IN), .ZN(n2538) );
  INV_X1 U32720 ( .A(DATAI_18_), .ZN(n4670) );
  NAND2_X1 U32730 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  XNOR2_X1 U32740 ( .A(n2542), .B(IR_REG_18__SCAN_IN), .ZN(n3970) );
  MUX2_X1 U32750 ( .A(n4670), .B(n4510), .S(n3402), .Z(n4207) );
  OR2_X1 U32760 ( .A1(n4299), .A2(n4207), .ZN(n4174) );
  NAND2_X1 U32770 ( .A1(n4299), .A2(n4207), .ZN(n4175) );
  NAND2_X1 U32780 ( .A1(n4174), .A2(n4175), .ZN(n4198) );
  INV_X1 U32790 ( .A(n4207), .ZN(n4199) );
  NAND2_X1 U32800 ( .A1(n4194), .A2(n2072), .ZN(n4171) );
  INV_X1 U32810 ( .A(n4171), .ZN(n2552) );
  INV_X1 U32820 ( .A(n2543), .ZN(n2553) );
  NAND2_X1 U32830 ( .A1(n2544), .A2(n4578), .ZN(n2545) );
  NAND2_X1 U32840 ( .A1(n2553), .A2(n2545), .ZN(n4188) );
  OR2_X1 U32850 ( .A1(n4188), .A2(n2619), .ZN(n2548) );
  AOI22_X1 U32860 ( .A1(n2337), .A2(REG2_REG_19__SCAN_IN), .B1(n3404), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2547) );
  INV_X1 U32870 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4292) );
  OR2_X1 U32880 ( .A1(n3407), .A2(n4292), .ZN(n2546) );
  INV_X1 U32890 ( .A(DATAI_19_), .ZN(n4667) );
  NOR2_X2 U32900 ( .A1(n2549), .A2(IR_REG_18__SCAN_IN), .ZN(n2627) );
  INV_X1 U32910 ( .A(n2627), .ZN(n2550) );
  MUX2_X1 U32920 ( .A(n4667), .B(n4002), .S(n3402), .Z(n4185) );
  INV_X1 U32930 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U32940 ( .A1(n2553), .A2(n4669), .ZN(n2554) );
  NAND2_X1 U32950 ( .A1(n4166), .A2(n2362), .ZN(n2560) );
  INV_X1 U32960 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U32970 ( .A1(n2337), .A2(REG2_REG_20__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U32980 ( .A1(n3404), .A2(REG0_REG_20__SCAN_IN), .ZN(n2556) );
  OAI211_X1 U32990 ( .C1(n4288), .C2(n3407), .A(n2557), .B(n2556), .ZN(n2558)
         );
  INV_X1 U33000 ( .A(n2558), .ZN(n2559) );
  INV_X1 U33010 ( .A(DATAI_20_), .ZN(n2561) );
  NAND2_X1 U33020 ( .A1(n4278), .A2(n4153), .ZN(n3460) );
  NOR2_X1 U33030 ( .A1(n4278), .A2(n4153), .ZN(n3462) );
  NAND2_X1 U33040 ( .A1(n2564), .A2(n3843), .ZN(n2565) );
  AND2_X1 U33050 ( .A1(n2572), .A2(n2565), .ZN(n4118) );
  NAND2_X1 U33060 ( .A1(n4118), .A2(n2362), .ZN(n2570) );
  INV_X1 U33070 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U33080 ( .A1(n3404), .A2(REG0_REG_22__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U33090 ( .A1(n2361), .A2(REG2_REG_22__SCAN_IN), .ZN(n2566) );
  OAI211_X1 U33100 ( .C1(n3407), .C2(n4274), .A(n2567), .B(n2566), .ZN(n2568)
         );
  INV_X1 U33110 ( .A(n2568), .ZN(n2569) );
  NAND2_X1 U33120 ( .A1(n2305), .A2(DATAI_22_), .ZN(n4117) );
  NAND2_X1 U33130 ( .A1(n4137), .A2(n4117), .ZN(n2656) );
  NAND2_X1 U33140 ( .A1(n4096), .A2(n2656), .ZN(n4121) );
  INV_X1 U33150 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U33160 ( .A1(n2572), .A2(n4581), .ZN(n2573) );
  NAND2_X1 U33170 ( .A1(n2580), .A2(n2573), .ZN(n4105) );
  OR2_X1 U33180 ( .A1(n4105), .A2(n2619), .ZN(n2578) );
  INV_X1 U33190 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U33200 ( .A1(n2337), .A2(REG2_REG_23__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U33210 ( .A1(n3404), .A2(REG0_REG_23__SCAN_IN), .ZN(n2574) );
  OAI211_X1 U33220 ( .C1(n4268), .C2(n3407), .A(n2575), .B(n2574), .ZN(n2576)
         );
  INV_X1 U33230 ( .A(n2576), .ZN(n2577) );
  NAND2_X1 U33240 ( .A1(n2305), .A2(DATAI_23_), .ZN(n4103) );
  NAND2_X1 U33250 ( .A1(n4085), .A2(n4103), .ZN(n2579) );
  INV_X1 U33260 ( .A(n4103), .ZN(n2711) );
  NAND2_X1 U33270 ( .A1(n2580), .A2(n4690), .ZN(n2581) );
  NAND2_X1 U33280 ( .A1(n2590), .A2(n2581), .ZN(n4080) );
  INV_X1 U33290 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U33300 ( .A1(n2361), .A2(REG2_REG_24__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33310 ( .A1(n3404), .A2(REG0_REG_24__SCAN_IN), .ZN(n2582) );
  OAI211_X1 U33320 ( .C1(n4264), .C2(n3407), .A(n2583), .B(n2582), .ZN(n2584)
         );
  INV_X1 U33330 ( .A(n2584), .ZN(n2585) );
  INV_X1 U33340 ( .A(DATAI_24_), .ZN(n2587) );
  NOR2_X1 U33350 ( .A1(n3402), .A2(n2587), .ZN(n4257) );
  INV_X1 U33360 ( .A(n4257), .ZN(n3813) );
  NAND2_X1 U33370 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2588) );
  INV_X1 U33380 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4681) );
  INV_X1 U33390 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2589) );
  OAI21_X1 U33400 ( .B1(n2590), .B2(n4681), .A(n2589), .ZN(n2591) );
  NAND2_X1 U33410 ( .A1(n4054), .A2(n2362), .ZN(n2596) );
  INV_X1 U33420 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U33430 ( .A1(n2361), .A2(REG2_REG_26__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U33440 ( .A1(n3404), .A2(REG0_REG_26__SCAN_IN), .ZN(n2592) );
  OAI211_X1 U33450 ( .C1(n4246), .C2(n3407), .A(n2593), .B(n2592), .ZN(n2594)
         );
  INV_X1 U33460 ( .A(n2594), .ZN(n2595) );
  NAND2_X1 U33470 ( .A1(n2305), .A2(DATAI_26_), .ZN(n4053) );
  NOR2_X1 U33480 ( .A1(n4252), .A2(n4053), .ZN(n2597) );
  INV_X1 U33490 ( .A(n4053), .ZN(n3876) );
  INV_X1 U33500 ( .A(n2600), .ZN(n2598) );
  NAND2_X1 U33510 ( .A1(n2598), .A2(REG3_REG_27__SCAN_IN), .ZN(n2610) );
  INV_X1 U33520 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U3353 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  NAND2_X1 U33540 ( .A1(n2610), .A2(n2601), .ZN(n4033) );
  INV_X1 U3355 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U3356 ( .A1(n2337), .A2(REG2_REG_27__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3357 ( .A1(n3404), .A2(REG0_REG_27__SCAN_IN), .ZN(n2602) );
  OAI211_X1 U3358 ( .C1(n4242), .C2(n3407), .A(n2603), .B(n2602), .ZN(n2604)
         );
  INV_X1 U3359 ( .A(n2604), .ZN(n2605) );
  INV_X1 U3360 ( .A(DATAI_27_), .ZN(n2607) );
  NOR2_X1 U3361 ( .A1(n3402), .A2(n2607), .ZN(n4235) );
  NOR2_X1 U3362 ( .A1(n3899), .A2(n4235), .ZN(n2608) );
  INV_X1 U3363 ( .A(n4235), .ZN(n4031) );
  INV_X1 U3364 ( .A(n2610), .ZN(n2609) );
  NAND2_X1 U3365 ( .A1(n2609), .A2(REG3_REG_28__SCAN_IN), .ZN(n4017) );
  INV_X1 U3366 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U3367 ( .A1(n2610), .A2(n3701), .ZN(n2611) );
  NAND2_X1 U3368 ( .A1(n4017), .A2(n2611), .ZN(n3700) );
  OR2_X1 U3369 ( .A1(n3700), .A2(n2619), .ZN(n2617) );
  INV_X1 U3370 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U3371 ( .A1(n2337), .A2(REG2_REG_28__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3372 ( .A1(n3404), .A2(REG0_REG_28__SCAN_IN), .ZN(n2612) );
  OAI211_X1 U3373 ( .C1(n2614), .C2(n3407), .A(n2613), .B(n2612), .ZN(n2615)
         );
  INV_X1 U3374 ( .A(n2615), .ZN(n2616) );
  INV_X1 U3375 ( .A(DATAI_28_), .ZN(n2618) );
  NOR2_X1 U3376 ( .A1(n3402), .A2(n2618), .ZN(n2712) );
  NAND2_X1 U3377 ( .A1(n4238), .A2(n2712), .ZN(n3413) );
  INV_X1 U3378 ( .A(n2712), .ZN(n4225) );
  NAND2_X1 U3379 ( .A1(n4036), .A2(n4225), .ZN(n3409) );
  NAND2_X1 U3380 ( .A1(n3413), .A2(n3409), .ZN(n3711) );
  AOI22_X1 U3381 ( .A1(n3706), .A2(n3711), .B1(n2712), .B2(n4036), .ZN(n2625)
         );
  OR2_X1 U3382 ( .A1(n4017), .A2(n2619), .ZN(n2624) );
  NAND2_X1 U3383 ( .A1(n2361), .A2(REG2_REG_29__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3384 ( .A1(n3404), .A2(REG0_REG_29__SCAN_IN), .ZN(n2620) );
  OAI211_X1 U3385 ( .C1(n2709), .C2(n3407), .A(n2621), .B(n2620), .ZN(n2622)
         );
  INV_X1 U3386 ( .A(n2622), .ZN(n2623) );
  NAND2_X1 U3387 ( .A1(n2624), .A2(n2623), .ZN(n4229) );
  NAND2_X1 U3388 ( .A1(n2305), .A2(DATAI_29_), .ZN(n4014) );
  XNOR2_X1 U3389 ( .A(n4229), .B(n4014), .ZN(n3444) );
  XNOR2_X1 U3390 ( .A(n2625), .B(n3444), .ZN(n4012) );
  NOR2_X1 U3391 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2626)
         );
  NAND2_X1 U3392 ( .A1(n2627), .A2(n2626), .ZN(n2632) );
  INV_X1 U3393 ( .A(n2632), .ZN(n2629) );
  NAND2_X1 U3394 ( .A1(n2629), .A2(n2628), .ZN(n2680) );
  NAND2_X1 U3395 ( .A1(n2680), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  INV_X1 U3396 ( .A(IR_REG_22__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3397 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  OR2_X2 U3398 ( .A1(n3455), .A2(n2726), .ZN(n2861) );
  XNOR2_X1 U3399 ( .A(n4379), .B(n2861), .ZN(n2636) );
  NAND2_X1 U3400 ( .A1(n2636), .A2(n4002), .ZN(n4160) );
  AND2_X1 U3401 ( .A1(n2637), .A2(n4381), .ZN(n2892) );
  NAND2_X1 U3402 ( .A1(n2892), .A2(n2839), .ZN(n4523) );
  NAND2_X1 U3403 ( .A1(n4160), .A2(n4523), .ZN(n4531) );
  NAND2_X1 U3404 ( .A1(n2839), .A2(n3455), .ZN(n2842) );
  OR2_X1 U3405 ( .A1(n2842), .A2(n2637), .ZN(n4226) );
  INV_X1 U3406 ( .A(n2815), .ZN(n2910) );
  NAND2_X1 U3407 ( .A1(n2910), .A2(n2916), .ZN(n3504) );
  NAND2_X1 U3408 ( .A1(n2930), .A2(n3472), .ZN(n2929) );
  NAND2_X1 U3409 ( .A1(n2640), .A2(n2963), .ZN(n3514) );
  NAND2_X1 U3410 ( .A1(n3913), .A2(n3001), .ZN(n3512) );
  INV_X1 U3411 ( .A(n3515), .ZN(n2641) );
  AND2_X1 U3412 ( .A1(n3911), .A2(n3127), .ZN(n3053) );
  NAND2_X1 U3413 ( .A1(n3103), .A2(n3100), .ZN(n3493) );
  NAND2_X1 U3414 ( .A1(n3910), .A2(n3118), .ZN(n3517) );
  NAND2_X1 U3415 ( .A1(n3041), .A2(n3517), .ZN(n2642) );
  NAND2_X1 U3416 ( .A1(n3113), .A2(n3075), .ZN(n3521) );
  INV_X1 U3417 ( .A(n2643), .ZN(n2644) );
  NAND2_X1 U3418 ( .A1(n3196), .A2(n3197), .ZN(n3527) );
  NAND2_X1 U3419 ( .A1(n3908), .A2(n3211), .ZN(n3524) );
  AND2_X1 U3420 ( .A1(n3907), .A2(n3227), .ZN(n3133) );
  NAND2_X1 U3421 ( .A1(n3283), .A2(n3220), .ZN(n3528) );
  NAND2_X1 U3422 ( .A1(n3906), .A2(n3284), .ZN(n3492) );
  NAND2_X1 U3423 ( .A1(n3323), .A2(n3274), .ZN(n3496) );
  NAND2_X1 U3424 ( .A1(n3904), .A2(n3767), .ZN(n3309) );
  NAND2_X1 U3425 ( .A1(n3903), .A2(n3835), .ZN(n2646) );
  NAND2_X1 U3426 ( .A1(n3309), .A2(n2646), .ZN(n3532) );
  INV_X1 U3427 ( .A(n3292), .ZN(n3534) );
  NOR2_X1 U3428 ( .A1(n3532), .A2(n3534), .ZN(n2647) );
  NAND2_X1 U3429 ( .A1(n3595), .A2(n3596), .ZN(n3310) );
  NAND2_X1 U3430 ( .A1(n3290), .A2(n3310), .ZN(n2650) );
  INV_X1 U3431 ( .A(n3532), .ZN(n2649) );
  NOR2_X1 U3432 ( .A1(n3903), .A2(n3835), .ZN(n2648) );
  AOI21_X1 U3433 ( .B1(n2650), .B2(n2649), .A(n2648), .ZN(n3535) );
  INV_X1 U3434 ( .A(n3242), .ZN(n3467) );
  NAND2_X1 U3435 ( .A1(n3425), .A2(n3467), .ZN(n2651) );
  NAND2_X1 U3436 ( .A1(n4309), .A2(n3618), .ZN(n3424) );
  NAND2_X1 U3437 ( .A1(n3901), .A2(n3891), .ZN(n3498) );
  NAND2_X1 U3438 ( .A1(n3424), .A2(n3498), .ZN(n3446) );
  INV_X1 U3439 ( .A(n3570), .ZN(n3579) );
  AND2_X1 U3440 ( .A1(n4200), .A2(n3802), .ZN(n3388) );
  NAND2_X1 U3441 ( .A1(n4154), .A2(n4185), .ZN(n3452) );
  NAND2_X1 U3442 ( .A1(n3452), .A2(n4175), .ZN(n3421) );
  INV_X1 U3443 ( .A(n4153), .ZN(n4164) );
  NAND2_X1 U3444 ( .A1(n4278), .A2(n4164), .ZN(n3419) );
  INV_X1 U3445 ( .A(n3419), .ZN(n2655) );
  NAND2_X1 U3446 ( .A1(n4315), .A2(n4297), .ZN(n4172) );
  AND2_X1 U3447 ( .A1(n4174), .A2(n4172), .ZN(n2652) );
  NAND2_X1 U3448 ( .A1(n4202), .A2(n2710), .ZN(n3453) );
  OAI21_X1 U3449 ( .B1(n3421), .B2(n2652), .A(n3453), .ZN(n4148) );
  NOR2_X1 U3450 ( .A1(n4278), .A2(n4164), .ZN(n2653) );
  OR2_X1 U3451 ( .A1(n4148), .A2(n2653), .ZN(n2654) );
  NAND2_X1 U3452 ( .A1(n2654), .A2(n3419), .ZN(n3541) );
  NAND2_X1 U3453 ( .A1(n4156), .A2(n4276), .ZN(n3445) );
  AND2_X1 U3454 ( .A1(n4096), .A2(n3445), .ZN(n3542) );
  INV_X1 U3455 ( .A(n3542), .ZN(n2658) );
  NAND2_X1 U3456 ( .A1(n4258), .A2(n4103), .ZN(n3450) );
  NAND2_X1 U3457 ( .A1(n3450), .A2(n2656), .ZN(n3491) );
  NOR2_X1 U34580 ( .A1(n4156), .A2(n4276), .ZN(n4093) );
  AND2_X1 U34590 ( .A1(n4096), .A2(n4093), .ZN(n2657) );
  NOR2_X1 U3460 ( .A1(n3491), .A2(n2657), .ZN(n3431) );
  NAND2_X1 U3461 ( .A1(n4085), .A2(n2711), .ZN(n3451) );
  NAND2_X1 U3462 ( .A1(n2659), .A2(n3451), .ZN(n4075) );
  NOR2_X1 U3463 ( .A1(n4249), .A2(n3813), .ZN(n3485) );
  NAND2_X1 U3464 ( .A1(n4252), .A2(n3876), .ZN(n2660) );
  OR2_X1 U3465 ( .A1(n4089), .A2(n4070), .ZN(n4044) );
  AND2_X1 U3466 ( .A1(n2660), .A2(n4044), .ZN(n2661) );
  INV_X1 U34670 ( .A(n2661), .ZN(n3544) );
  NAND2_X1 U3468 ( .A1(n4089), .A2(n4070), .ZN(n3484) );
  NAND2_X1 U34690 ( .A1(n4249), .A2(n3813), .ZN(n4059) );
  NAND2_X1 U3470 ( .A1(n3484), .A2(n4059), .ZN(n4045) );
  AND2_X1 U34710 ( .A1(n4236), .A2(n4053), .ZN(n3411) );
  AOI21_X1 U3472 ( .B1(n2661), .B2(n4045), .A(n3411), .ZN(n3550) );
  XNOR2_X1 U34730 ( .A(n3899), .B(n4031), .ZN(n4025) );
  NAND2_X1 U3474 ( .A1(n4227), .A2(n4235), .ZN(n3412) );
  INV_X1 U34750 ( .A(n3413), .ZN(n2662) );
  XNOR2_X1 U3476 ( .A(n2663), .B(n3444), .ZN(n2674) );
  NAND2_X1 U34770 ( .A1(n4379), .A2(n4381), .ZN(n2664) );
  NAND2_X1 U3478 ( .A1(n4380), .A2(n2726), .ZN(n3440) );
  NOR2_X1 U34790 ( .A1(n2666), .A2(n2665), .ZN(n2822) );
  MUX2_X1 U3480 ( .A(n2729), .B(n2667), .S(IR_REG_28__SCAN_IN), .Z(n2670) );
  INV_X1 U34810 ( .A(n2668), .ZN(n2669) );
  NAND2_X1 U3482 ( .A1(n4379), .A2(n4380), .ZN(n2843) );
  INV_X1 U34830 ( .A(n2843), .ZN(n2734) );
  NAND2_X1 U3484 ( .A1(n2853), .A2(n2734), .ZN(n4314) );
  AOI21_X1 U34850 ( .B1(B_REG_SCAN_IN), .B2(n2822), .A(n4314), .ZN(n4007) );
  INV_X1 U3486 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U34870 ( .A1(n2337), .A2(REG2_REG_30__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3488 ( .A1(n3404), .A2(REG0_REG_30__SCAN_IN), .ZN(n2671) );
  OAI211_X1 U34890 ( .C1(n3407), .C2(n2673), .A(n2672), .B(n2671), .ZN(n3898)
         );
  NOR2_X2 U3490 ( .A1(n2853), .A2(n2843), .ZN(n4277) );
  NAND2_X1 U34910 ( .A1(n4036), .A2(n4277), .ZN(n2675) );
  NAND2_X1 U3492 ( .A1(n2676), .A2(IR_REG_31__SCAN_IN), .ZN(n2677) );
  MUX2_X1 U34930 ( .A(IR_REG_31__SCAN_IN), .B(n2677), .S(IR_REG_25__SCAN_IN), 
        .Z(n2679) );
  NAND2_X1 U3494 ( .A1(n2679), .A2(n2678), .ZN(n2724) );
  NAND2_X1 U34950 ( .A1(n2724), .A2(B_REG_SCAN_IN), .ZN(n2683) );
  INV_X1 U3496 ( .A(IR_REG_23__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U34970 ( .A1(n2690), .A2(n2691), .ZN(n2681) );
  MUX2_X1 U3498 ( .A(n2683), .B(B_REG_SCAN_IN), .S(n2689), .Z(n2687) );
  NAND2_X1 U34990 ( .A1(n2678), .A2(IR_REG_31__SCAN_IN), .ZN(n2684) );
  MUX2_X1 U3500 ( .A(IR_REG_31__SCAN_IN), .B(n2684), .S(IR_REG_26__SCAN_IN), 
        .Z(n2686) );
  NAND2_X1 U35010 ( .A1(n2706), .A2(n2724), .ZN(n2836) );
  NAND2_X1 U3502 ( .A1(n2883), .A2(n2836), .ZN(n2705) );
  XNOR2_X1 U35030 ( .A(n2690), .B(n2691), .ZN(n2733) );
  NAND2_X1 U3504 ( .A1(n2733), .A2(STATE_REG_SCAN_IN), .ZN(n4508) );
  INV_X1 U35050 ( .A(n4508), .ZN(n2738) );
  OR2_X1 U35060 ( .A1(n4523), .A2(n4380), .ZN(n2849) );
  AND2_X1 U35070 ( .A1(n2637), .A2(n4002), .ZN(n2841) );
  OR2_X1 U35080 ( .A1(n2843), .A2(n2841), .ZN(n2880) );
  NAND2_X1 U35090 ( .A1(n2849), .A2(n2880), .ZN(n2692) );
  NOR2_X1 U35100 ( .A1(n2882), .A2(n2692), .ZN(n2704) );
  NOR4_X1 U35110 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2696) );
  NOR4_X1 U35120 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2695) );
  NOR4_X1 U35130 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2694) );
  NOR4_X1 U35140 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2693) );
  NAND4_X1 U35150 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n2702)
         );
  NOR2_X1 U35160 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2700) );
  NOR4_X1 U35170 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2699) );
  NOR4_X1 U35180 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2698) );
  NOR4_X1 U35190 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2697) );
  NAND4_X1 U35200 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .ZN(n2701)
         );
  NOR2_X1 U35210 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND3_X1 U35220 ( .A1(n2705), .A2(n2704), .A3(n2837), .ZN(n2717) );
  NAND2_X1 U35230 ( .A1(n3585), .A2(n2706), .ZN(n2707) );
  MUX2_X1 U35240 ( .A(n2709), .B(n2718), .S(n4545), .Z(n2716) );
  NOR2_X1 U35250 ( .A1(n2936), .A2(n3032), .ZN(n2965) );
  NAND2_X1 U35260 ( .A1(n2965), .A2(n3001), .ZN(n2986) );
  INV_X1 U35270 ( .A(n4014), .ZN(n3410) );
  NAND2_X1 U35280 ( .A1(n2056), .A2(n3410), .ZN(n2713) );
  NAND2_X1 U35290 ( .A1(n2052), .A2(n2713), .ZN(n4018) );
  INV_X1 U35300 ( .A(n2842), .ZN(n2890) );
  NAND2_X1 U35310 ( .A1(n2716), .A2(n2715), .ZN(U3547) );
  INV_X1 U35320 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U35330 ( .A1(n2721), .A2(n2720), .ZN(n2722) );
  INV_X2 U35340 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X2 U35350 ( .A1(n2811), .A2(n4508), .ZN(n3915) );
  NAND2_X1 U35360 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2723) );
  OAI21_X1 U35370 ( .B1(n2724), .B2(U3149), .A(n2723), .ZN(U3327) );
  INV_X1 U35380 ( .A(DATAI_26_), .ZN(n4678) );
  NAND2_X1 U35390 ( .A1(n3584), .A2(STATE_REG_SCAN_IN), .ZN(n2725) );
  OAI21_X1 U35400 ( .B1(STATE_REG_SCAN_IN), .B2(n4678), .A(n2725), .ZN(U3326)
         );
  NAND2_X1 U35410 ( .A1(n2726), .A2(STATE_REG_SCAN_IN), .ZN(n2727) );
  OAI21_X1 U35420 ( .B1(STATE_REG_SCAN_IN), .B2(n2561), .A(n2727), .ZN(U3332)
         );
  NAND2_X1 U35430 ( .A1(n2822), .A2(STATE_REG_SCAN_IN), .ZN(n2728) );
  OAI21_X1 U35440 ( .B1(STATE_REG_SCAN_IN), .B2(n2607), .A(n2728), .ZN(U3325)
         );
  INV_X1 U35450 ( .A(DATAI_31_), .ZN(n4551) );
  OR4_X1 U35460 ( .A1(n2730), .A2(IR_REG_30__SCAN_IN), .A3(n2729), .A4(U3149), 
        .ZN(n2731) );
  OAI21_X1 U35470 ( .B1(STATE_REG_SCAN_IN), .B2(n4551), .A(n2731), .ZN(U3321)
         );
  INV_X1 U35480 ( .A(n2853), .ZN(n2873) );
  NAND2_X1 U35490 ( .A1(n2873), .A2(STATE_REG_SCAN_IN), .ZN(n2732) );
  OAI21_X1 U35500 ( .B1(STATE_REG_SCAN_IN), .B2(n2618), .A(n2732), .ZN(U3324)
         );
  OR2_X1 U35510 ( .A1(n2733), .A2(U3149), .ZN(n3567) );
  NAND2_X1 U35520 ( .A1(n2882), .A2(n3567), .ZN(n2742) );
  AOI21_X1 U35530 ( .B1(n2734), .B2(n2733), .A(n3402), .ZN(n2741) );
  INV_X1 U35540 ( .A(n2741), .ZN(n2735) );
  NOR2_X1 U35550 ( .A1(n4489), .A2(n3915), .ZN(U3148) );
  INV_X1 U35560 ( .A(n2882), .ZN(n2736) );
  INV_X1 U35570 ( .A(D_REG_1__SCAN_IN), .ZN(n2740) );
  INV_X1 U35580 ( .A(n2836), .ZN(n2739) );
  AOI22_X1 U35590 ( .A1(n4507), .A2(n2740), .B1(n2739), .B2(n2738), .ZN(U3459)
         );
  INV_X1 U35600 ( .A(n2774), .ZN(n2746) );
  AOI21_X1 U35610 ( .B1(n2822), .B2(n2743), .A(n2853), .ZN(n2824) );
  OAI21_X1 U35620 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2822), .A(n2824), .ZN(n2744) );
  MUX2_X1 U35630 ( .A(n2744), .B(n2824), .S(IR_REG_0__SCAN_IN), .Z(n2745) );
  INV_X1 U35640 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2858) );
  OAI22_X1 U35650 ( .A1(n2746), .A2(n2745), .B1(STATE_REG_SCAN_IN), .B2(n2858), 
        .ZN(n2747) );
  AOI21_X1 U35660 ( .B1(n4489), .B2(ADDR_REG_0__SCAN_IN), .A(n2747), .ZN(n2749) );
  INV_X1 U35670 ( .A(n2822), .ZN(n2759) );
  INV_X1 U35680 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4540) );
  NAND3_X1 U35690 ( .A1(n4491), .A2(IR_REG_0__SCAN_IN), .A3(n4540), .ZN(n2748)
         );
  NAND2_X1 U35700 ( .A1(n2749), .A2(n2748), .ZN(U3240) );
  INV_X1 U35710 ( .A(n4389), .ZN(n3928) );
  MUX2_X1 U35720 ( .A(REG2_REG_2__SCAN_IN), .B(n2750), .S(n4389), .Z(n2754) );
  INV_X1 U35730 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2751) );
  MUX2_X1 U35740 ( .A(REG2_REG_1__SCAN_IN), .B(n2751), .S(n4390), .Z(n3920) );
  AND2_X1 U35750 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U35760 ( .A1(n3920), .A2(n2752), .ZN(n3931) );
  NAND2_X1 U35770 ( .A1(n4390), .A2(REG2_REG_1__SCAN_IN), .ZN(n3930) );
  NAND2_X1 U35780 ( .A1(n3931), .A2(n3930), .ZN(n2753) );
  XNOR2_X1 U35790 ( .A(n2755), .B(n4387), .ZN(n2825) );
  INV_X1 U35800 ( .A(n2755), .ZN(n2756) );
  MUX2_X1 U35810 ( .A(REG2_REG_5__SCAN_IN), .B(n2394), .S(n2787), .Z(n2784) );
  NOR2_X1 U3582 ( .A1(n2785), .A2(n2784), .ZN(n2783) );
  AOI21_X1 U3583 ( .B1(n4386), .B2(REG2_REG_5__SCAN_IN), .A(n2783), .ZN(n2757)
         );
  XNOR2_X1 U3584 ( .A(n2757), .B(n4385), .ZN(n2791) );
  INV_X1 U3585 ( .A(n2757), .ZN(n2758) );
  MUX2_X1 U3586 ( .A(n2416), .B(REG2_REG_7__SCAN_IN), .S(n4384), .Z(n2760) );
  NOR2_X1 U3587 ( .A1(n2853), .A2(n2759), .ZN(n3563) );
  AOI211_X1 U3588 ( .C1(n2761), .C2(n2760), .A(n4485), .B(n2805), .ZN(n2779)
         );
  XNOR2_X1 U3589 ( .A(n4389), .B(n2762), .ZN(n3937) );
  XNOR2_X1 U3590 ( .A(n4390), .B(n2360), .ZN(n3918) );
  AND2_X1 U3591 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3917)
         );
  NAND2_X1 U3592 ( .A1(n3918), .A2(n3917), .ZN(n3916) );
  NAND2_X1 U3593 ( .A1(n4390), .A2(REG1_REG_1__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U3594 ( .A1(n3916), .A2(n2763), .ZN(n3936) );
  NAND2_X1 U3595 ( .A1(n3937), .A2(n3936), .ZN(n3935) );
  NAND2_X1 U3596 ( .A1(n4389), .A2(REG1_REG_2__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U3597 ( .A1(n3935), .A2(n2764), .ZN(n2766) );
  INV_X1 U3598 ( .A(n4388), .ZN(n2765) );
  XNOR2_X1 U3599 ( .A(n2766), .B(n2765), .ZN(n3944) );
  NAND2_X1 U3600 ( .A1(n3944), .A2(REG1_REG_3__SCAN_IN), .ZN(n3943) );
  NAND2_X1 U3601 ( .A1(n2766), .A2(n4388), .ZN(n2767) );
  NAND2_X1 U3602 ( .A1(n3943), .A2(n2767), .ZN(n2768) );
  INV_X1 U3603 ( .A(n4387), .ZN(n2832) );
  XNOR2_X1 U3604 ( .A(n2768), .B(n2832), .ZN(n2828) );
  XNOR2_X1 U3605 ( .A(n4386), .B(REG1_REG_5__SCAN_IN), .ZN(n2781) );
  INV_X1 U3606 ( .A(n2769), .ZN(n2770) );
  NOR2_X1 U3607 ( .A1(n2796), .A2(n2409), .ZN(n2794) );
  INV_X1 U3608 ( .A(n4384), .ZN(n2776) );
  AND2_X1 U3609 ( .A1(n2776), .A2(n2419), .ZN(n2801) );
  INV_X1 U3610 ( .A(n2801), .ZN(n2771) );
  NAND2_X1 U3611 ( .A1(n4384), .A2(REG1_REG_7__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U3612 ( .A1(n2771), .A2(n2802), .ZN(n2773) );
  OAI21_X1 U3613 ( .B1(n2803), .B2(n2773), .A(n4491), .ZN(n2772) );
  AOI21_X1 U3614 ( .B1(n2803), .B2(n2773), .A(n2772), .ZN(n2778) );
  NAND2_X1 U3615 ( .A1(n2774), .A2(n2853), .ZN(n4495) );
  AND2_X1 U3616 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3168) );
  AOI21_X1 U3617 ( .B1(n4489), .B2(ADDR_REG_7__SCAN_IN), .A(n3168), .ZN(n2775)
         );
  OAI21_X1 U3618 ( .B1(n4495), .B2(n2776), .A(n2775), .ZN(n2777) );
  OR3_X1 U3619 ( .A1(n2779), .A2(n2778), .A3(n2777), .ZN(U3247) );
  INV_X1 U3620 ( .A(n4491), .ZN(n2795) );
  AOI211_X1 U3621 ( .C1(n2782), .C2(n2781), .A(n2780), .B(n2795), .ZN(n2790)
         );
  AOI211_X1 U3622 ( .C1(n2785), .C2(n2784), .A(n2783), .B(n4485), .ZN(n2789)
         );
  INV_X1 U3623 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U3624 ( .A1(STATE_REG_SCAN_IN), .A2(n4665), .ZN(n3129) );
  AOI21_X1 U3625 ( .B1(n4489), .B2(ADDR_REG_5__SCAN_IN), .A(n3129), .ZN(n2786)
         );
  OAI21_X1 U3626 ( .B1(n4495), .B2(n2787), .A(n2786), .ZN(n2788) );
  OR3_X1 U3627 ( .A1(n2790), .A2(n2789), .A3(n2788), .ZN(U3245) );
  XNOR2_X1 U3628 ( .A(n2791), .B(REG2_REG_6__SCAN_IN), .ZN(n2800) );
  INV_X1 U3629 ( .A(n4495), .ZN(n3942) );
  NOR2_X1 U3630 ( .A1(STATE_REG_SCAN_IN), .A2(n2792), .ZN(n3115) );
  AOI21_X1 U3631 ( .B1(n4489), .B2(ADDR_REG_6__SCAN_IN), .A(n3115), .ZN(n2793)
         );
  INV_X1 U3632 ( .A(n2793), .ZN(n2798) );
  AOI211_X1 U3633 ( .C1(n2796), .C2(n2409), .A(n2795), .B(n2794), .ZN(n2797)
         );
  AOI211_X1 U3634 ( .C1(n3942), .C2(n4385), .A(n2798), .B(n2797), .ZN(n2799)
         );
  OAI21_X1 U3635 ( .B1(n2800), .B2(n4485), .A(n2799), .ZN(U3246) );
  AOI21_X1 U3636 ( .B1(n2803), .B2(n2802), .A(n2801), .ZN(n3976) );
  XNOR2_X1 U3637 ( .A(n3976), .B(n4382), .ZN(n3975) );
  XOR2_X1 U3638 ( .A(REG1_REG_8__SCAN_IN), .B(n3975), .Z(n2804) );
  NAND2_X1 U3639 ( .A1(n2804), .A2(n4491), .ZN(n2810) );
  XNOR2_X1 U3640 ( .A(REG2_REG_8__SCAN_IN), .B(n3956), .ZN(n2806) );
  NAND2_X1 U3641 ( .A1(n4438), .A2(n2806), .ZN(n2807) );
  NAND2_X1 U3642 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3212) );
  NAND2_X1 U3643 ( .A1(n2807), .A2(n3212), .ZN(n2808) );
  AOI21_X1 U3644 ( .B1(n4489), .B2(ADDR_REG_8__SCAN_IN), .A(n2808), .ZN(n2809)
         );
  OAI211_X1 U3645 ( .C1(n4495), .C2(n4382), .A(n2810), .B(n2809), .ZN(U3248)
         );
  NAND2_X1 U3646 ( .A1(n2815), .A2(n3273), .ZN(n2813) );
  NAND2_X1 U3647 ( .A1(n2045), .A2(n2916), .ZN(n2812) );
  AND2_X1 U3648 ( .A1(n2813), .A2(n2812), .ZN(n2867) );
  INV_X1 U3649 ( .A(n2811), .ZN(n2950) );
  NAND2_X1 U3650 ( .A1(n2950), .A2(REG1_REG_0__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U3651 ( .A1(n2867), .A2(n2814), .ZN(n2820) );
  INV_X1 U3652 ( .A(n2943), .ZN(n2816) );
  NAND2_X1 U3653 ( .A1(n2816), .A2(n2815), .ZN(n2818) );
  AOI22_X1 U3654 ( .A1(n3273), .A2(n2916), .B1(n2950), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2817) );
  NAND2_X1 U3655 ( .A1(n2818), .A2(n2817), .ZN(n2819) );
  NAND2_X1 U3656 ( .A1(n2820), .A2(n2819), .ZN(n2870) );
  OAI21_X1 U3657 ( .B1(n2820), .B2(n2819), .A(n2870), .ZN(n2855) );
  NAND2_X1 U3658 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3919) );
  AOI21_X1 U3659 ( .B1(n2822), .B2(n3919), .A(n2853), .ZN(n2821) );
  OAI21_X1 U3660 ( .B1(n2855), .B2(n2822), .A(n2821), .ZN(n2823) );
  OAI211_X1 U3661 ( .C1(IR_REG_0__SCAN_IN), .C2(n2824), .A(n2823), .B(n3915), 
        .ZN(n3941) );
  XOR2_X1 U3662 ( .A(REG2_REG_4__SCAN_IN), .B(n2825), .Z(n2834) );
  INV_X1 U3663 ( .A(n2826), .ZN(n2827) );
  OAI211_X1 U3664 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2828), .A(n4491), .B(n2827), 
        .ZN(n2831) );
  NAND2_X1 U3665 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3023) );
  INV_X1 U3666 ( .A(n3023), .ZN(n2829) );
  AOI21_X1 U3667 ( .B1(n4489), .B2(ADDR_REG_4__SCAN_IN), .A(n2829), .ZN(n2830)
         );
  OAI211_X1 U3668 ( .C1(n4495), .C2(n2832), .A(n2831), .B(n2830), .ZN(n2833)
         );
  AOI21_X1 U3669 ( .B1(n4438), .B2(n2834), .A(n2833), .ZN(n2835) );
  NAND2_X1 U3670 ( .A1(n3941), .A2(n2835), .ZN(U3244) );
  NAND3_X1 U3671 ( .A1(n2838), .A2(n2886), .A3(n2883), .ZN(n2875) );
  OR2_X1 U3672 ( .A1(n2862), .A2(n4508), .ZN(n2840) );
  NOR2_X1 U3673 ( .A1(n3693), .A2(n2840), .ZN(n3564) );
  NAND2_X1 U3674 ( .A1(n2875), .A2(n3564), .ZN(n2952) );
  INV_X1 U3675 ( .A(n2952), .ZN(n2847) );
  OR2_X1 U3676 ( .A1(n2842), .A2(n2841), .ZN(n2844) );
  NAND2_X1 U3677 ( .A1(n2844), .A2(n2843), .ZN(n2851) );
  NAND2_X1 U3678 ( .A1(n2851), .A2(n4226), .ZN(n2845) );
  NAND2_X1 U3679 ( .A1(n2875), .A2(n2845), .ZN(n2846) );
  NAND2_X1 U3680 ( .A1(n2846), .A2(n2880), .ZN(n2951) );
  NOR3_X1 U3681 ( .A1(n2847), .A2(n2951), .A3(n2882), .ZN(n2902) );
  OR2_X1 U3682 ( .A1(n2882), .A2(n4226), .ZN(n2848) );
  OR2_X1 U3683 ( .A1(n2875), .A2(n2848), .ZN(n2850) );
  AND2_X2 U3684 ( .A1(n2850), .A2(n4496), .ZN(n3868) );
  INV_X1 U3685 ( .A(n3868), .ZN(n3877) );
  OR2_X1 U3686 ( .A1(n2882), .A2(n2851), .ZN(n2852) );
  NAND2_X1 U3687 ( .A1(n3564), .A2(n2853), .ZN(n2854) );
  OAI22_X1 U3688 ( .A1(n2855), .A2(n3896), .B1(n3845), .B2(n2928), .ZN(n2856)
         );
  AOI21_X1 U3689 ( .B1(n2916), .B2(n3877), .A(n2856), .ZN(n2857) );
  OAI21_X1 U3690 ( .B1(n2902), .B2(n2858), .A(n2857), .ZN(U3229) );
  INV_X1 U3691 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3006) );
  OR2_X1 U3692 ( .A1(n2928), .A2(n2943), .ZN(n2865) );
  NAND2_X1 U3693 ( .A1(n3273), .A2(n3011), .ZN(n2864) );
  NAND2_X1 U3694 ( .A1(n2865), .A2(n2864), .ZN(n2866) );
  INV_X1 U3695 ( .A(n2866), .ZN(n2897) );
  INV_X1 U3696 ( .A(n2867), .ZN(n2868) );
  NAND2_X1 U3697 ( .A1(n2870), .A2(n2869), .ZN(n2871) );
  OAI211_X1 U3698 ( .C1(n2872), .C2(n2871), .A(n2899), .B(n3764), .ZN(n2878)
         );
  NAND2_X1 U3699 ( .A1(n3564), .A2(n2873), .ZN(n2874) );
  OAI22_X1 U3700 ( .A1(n2910), .A2(n3844), .B1(n3845), .B2(n2949), .ZN(n2876)
         );
  AOI21_X1 U3701 ( .B1(n3011), .B2(n3877), .A(n2876), .ZN(n2877) );
  OAI211_X1 U3702 ( .C1(n2902), .C2(n3006), .A(n2878), .B(n2877), .ZN(U3219)
         );
  NAND2_X1 U3703 ( .A1(n2815), .A2(n2879), .ZN(n3506) );
  AND2_X1 U3704 ( .A1(n3504), .A2(n3506), .ZN(n4524) );
  INV_X1 U3705 ( .A(n2880), .ZN(n2881) );
  NOR2_X1 U3706 ( .A1(n2882), .A2(n2881), .ZN(n2885) );
  NAND4_X1 U3707 ( .A1(n2886), .A2(n2885), .A3(n2884), .A4(n2883), .ZN(n2887)
         );
  NAND2_X2 U3708 ( .A1(n2887), .A2(n4496), .ZN(n4191) );
  NAND2_X1 U3709 ( .A1(n2888), .A2(n4381), .ZN(n2993) );
  INV_X1 U3710 ( .A(n2993), .ZN(n2889) );
  AND2_X1 U3711 ( .A1(n4191), .A2(n2889), .ZN(n4502) );
  INV_X1 U3712 ( .A(n4502), .ZN(n3265) );
  NAND2_X1 U3713 ( .A1(n2916), .A2(n2890), .ZN(n4521) );
  AOI21_X1 U3714 ( .B1(n4182), .B2(n4160), .A(n4524), .ZN(n2891) );
  AOI21_X1 U3715 ( .B1(n4298), .B2(n3914), .A(n2891), .ZN(n4522) );
  OAI21_X1 U3716 ( .B1(n2892), .B2(n4521), .A(n4522), .ZN(n2893) );
  INV_X1 U3717 ( .A(n4496), .ZN(n4209) );
  AOI22_X1 U3718 ( .A1(n2893), .A2(n4191), .B1(REG3_REG_0__SCAN_IN), .B2(n4209), .ZN(n2895) );
  NAND2_X1 U3719 ( .A1(n4119), .A2(REG2_REG_0__SCAN_IN), .ZN(n2894) );
  OAI211_X1 U3720 ( .C1(n4524), .C2(n3265), .A(n2895), .B(n2894), .ZN(U3290)
         );
  XNOR2_X1 U3721 ( .A(n2896), .B(n3613), .ZN(n2944) );
  XNOR2_X1 U3722 ( .A(n2944), .B(n2945), .ZN(n2901) );
  NAND2_X1 U3723 ( .A1(n2899), .A2(n2898), .ZN(n2900) );
  AOI21_X1 U3724 ( .B1(n2901), .B2(n2900), .A(n2948), .ZN(n2906) );
  OAI22_X1 U3725 ( .A1(n2640), .A2(n3845), .B1(n3844), .B2(n2928), .ZN(n2904)
         );
  NOR2_X1 U3726 ( .A1(n2902), .A2(n3925), .ZN(n2903) );
  AOI211_X1 U3727 ( .C1(n3032), .C2(n3877), .A(n2904), .B(n2903), .ZN(n2905)
         );
  OAI21_X1 U3728 ( .B1(n2906), .B2(n3896), .A(n2905), .ZN(U3234) );
  INV_X1 U3729 ( .A(n4523), .ZN(n4529) );
  OAI21_X1 U3730 ( .B1(n2638), .B2(n2908), .A(n2907), .ZN(n3007) );
  INV_X1 U3731 ( .A(n3007), .ZN(n2915) );
  AOI22_X1 U3732 ( .A1(n2087), .A2(n4298), .B1(n4310), .B2(n3011), .ZN(n2909)
         );
  OAI21_X1 U3733 ( .B1(n2910), .B2(n4308), .A(n2909), .ZN(n2914) );
  INV_X1 U3734 ( .A(n2911), .ZN(n2912) );
  AOI21_X1 U3735 ( .B1(n2638), .B2(n3504), .A(n2912), .ZN(n2913) );
  OAI22_X1 U3736 ( .A1(n2913), .A2(n4182), .B1(n4160), .B2(n3007), .ZN(n3008)
         );
  AOI211_X1 U3737 ( .C1(n4529), .C2(n2915), .A(n2914), .B(n3008), .ZN(n2922)
         );
  NAND2_X1 U3738 ( .A1(n3011), .A2(n2916), .ZN(n2917) );
  NAND2_X1 U3739 ( .A1(n2936), .A2(n2917), .ZN(n3014) );
  OAI22_X1 U3740 ( .A1(n4307), .A2(n3014), .B1(n4545), .B2(n2360), .ZN(n2918)
         );
  INV_X1 U3741 ( .A(n2918), .ZN(n2919) );
  OAI21_X1 U3742 ( .B1(n2922), .B2(n4543), .A(n2919), .ZN(U3519) );
  OAI22_X1 U3743 ( .A1(n4369), .A2(n3014), .B1(n4539), .B2(n2363), .ZN(n2920)
         );
  INV_X1 U3744 ( .A(n2920), .ZN(n2921) );
  OAI21_X1 U3745 ( .B1(n2922), .B2(n4537), .A(n2921), .ZN(U3469) );
  NAND2_X1 U3746 ( .A1(n2907), .A2(n2923), .ZN(n2924) );
  OR2_X1 U3747 ( .A1(n2924), .A2(n3472), .ZN(n2926) );
  NAND2_X1 U3748 ( .A1(n2924), .A2(n3472), .ZN(n2925) );
  NAND2_X1 U3749 ( .A1(n2926), .A2(n2925), .ZN(n3031) );
  AOI22_X1 U3750 ( .A1(n3913), .A2(n4298), .B1(n3032), .B2(n4310), .ZN(n2927)
         );
  OAI21_X1 U3751 ( .B1(n2928), .B2(n4308), .A(n2927), .ZN(n2934) );
  INV_X1 U3752 ( .A(n4160), .ZN(n3151) );
  NAND2_X1 U3753 ( .A1(n3031), .A2(n3151), .ZN(n2933) );
  OAI21_X1 U3754 ( .B1(n3472), .B2(n2930), .A(n2929), .ZN(n2931) );
  NAND2_X1 U3755 ( .A1(n2931), .A2(n4204), .ZN(n2932) );
  NAND2_X1 U3756 ( .A1(n2933), .A2(n2932), .ZN(n3029) );
  AOI211_X1 U3757 ( .C1(n4529), .C2(n3031), .A(n2934), .B(n3029), .ZN(n2939)
         );
  XNOR2_X1 U3758 ( .A(n2936), .B(n2935), .ZN(n3033) );
  AOI22_X1 U3759 ( .A1(n2720), .A2(n3033), .B1(REG0_REG_2__SCAN_IN), .B2(n4537), .ZN(n2937) );
  OAI21_X1 U3760 ( .B1(n2939), .B2(n4537), .A(n2937), .ZN(U3471) );
  AOI22_X1 U3761 ( .A1(n2714), .A2(n3033), .B1(REG1_REG_2__SCAN_IN), .B2(n4543), .ZN(n2938) );
  OAI21_X1 U3762 ( .B1(n2939), .B2(n4543), .A(n2938), .ZN(U3520) );
  NAND2_X1 U3763 ( .A1(n3913), .A2(n3273), .ZN(n2941) );
  NAND2_X1 U3764 ( .A1(n2045), .A2(n2963), .ZN(n2940) );
  NAND2_X1 U3765 ( .A1(n2941), .A2(n2940), .ZN(n2942) );
  OAI22_X1 U3766 ( .A1(n2640), .A2(n3694), .B1(n3693), .B2(n3001), .ZN(n3016)
         );
  XNOR2_X1 U3767 ( .A(n3017), .B(n3016), .ZN(n3018) );
  INV_X1 U3768 ( .A(n2944), .ZN(n2947) );
  INV_X1 U3769 ( .A(n2945), .ZN(n2946) );
  XOR2_X1 U3770 ( .A(n3018), .B(n3019), .Z(n2958) );
  OAI21_X1 U3771 ( .B1(n2951), .B2(n2950), .A(STATE_REG_SCAN_IN), .ZN(n2954)
         );
  AND2_X1 U3772 ( .A1(n2952), .A2(n3567), .ZN(n2953) );
  MUX2_X1 U3773 ( .A(n3893), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2955) );
  AOI211_X1 U3774 ( .C1(n2963), .C2(n3877), .A(n2956), .B(n2955), .ZN(n2957)
         );
  OAI21_X1 U3775 ( .B1(n2958), .B2(n3896), .A(n2957), .ZN(U3215) );
  INV_X1 U3776 ( .A(n4531), .ZN(n4321) );
  XNOR2_X1 U3777 ( .A(n2959), .B(n3471), .ZN(n3005) );
  OAI21_X1 U3778 ( .B1(n3471), .B2(n2961), .A(n2960), .ZN(n2962) );
  AOI22_X1 U3779 ( .A1(n2962), .A2(n4204), .B1(n4277), .B2(n2087), .ZN(n2995)
         );
  AOI22_X1 U3780 ( .A1(n3912), .A2(n4298), .B1(n4310), .B2(n2963), .ZN(n2964)
         );
  OAI211_X1 U3781 ( .C1(n4321), .C2(n3005), .A(n2995), .B(n2964), .ZN(n2970)
         );
  OR2_X1 U3782 ( .A1(n2965), .A2(n3001), .ZN(n2966) );
  NAND2_X1 U3783 ( .A1(n2966), .A2(n2986), .ZN(n2997) );
  OAI22_X1 U3784 ( .A1(n4307), .A2(n2997), .B1(n4545), .B2(n2967), .ZN(n2968)
         );
  AOI21_X1 U3785 ( .B1(n2970), .B2(n4545), .A(n2968), .ZN(n2969) );
  INV_X1 U3786 ( .A(n2969), .ZN(U3521) );
  NAND2_X1 U3787 ( .A1(n2970), .A2(n4539), .ZN(n2972) );
  NAND2_X1 U3788 ( .A1(n4537), .A2(REG0_REG_3__SCAN_IN), .ZN(n2971) );
  OAI211_X1 U3789 ( .C1(n2997), .C2(n4369), .A(n2972), .B(n2971), .ZN(U3473)
         );
  NAND2_X1 U3790 ( .A1(n2959), .A2(n2973), .ZN(n2976) );
  NAND2_X1 U3791 ( .A1(n2976), .A2(n2974), .ZN(n2980) );
  NAND2_X1 U3792 ( .A1(n2976), .A2(n2975), .ZN(n2978) );
  NAND2_X1 U3793 ( .A1(n2978), .A2(n3473), .ZN(n2979) );
  INV_X1 U3794 ( .A(n4530), .ZN(n2992) );
  XOR2_X1 U3795 ( .A(n3473), .B(n2981), .Z(n2985) );
  AOI22_X1 U3796 ( .A1(n3913), .A2(n4277), .B1(n2987), .B2(n4310), .ZN(n2982)
         );
  OAI21_X1 U3797 ( .B1(n3103), .B2(n4314), .A(n2982), .ZN(n2983) );
  AOI21_X1 U3798 ( .B1(n4530), .B2(n3151), .A(n2983), .ZN(n2984) );
  OAI21_X1 U3799 ( .B1(n2985), .B2(n4182), .A(n2984), .ZN(n4527) );
  INV_X1 U3800 ( .A(n2986), .ZN(n2988) );
  OAI211_X1 U3801 ( .C1(n2988), .C2(n2167), .A(n4317), .B(n3058), .ZN(n4526)
         );
  OAI22_X1 U3802 ( .A1(n4526), .A2(n4381), .B1(n4496), .B2(n3028), .ZN(n2989)
         );
  OAI21_X1 U3803 ( .B1(n4527), .B2(n2989), .A(n4191), .ZN(n2991) );
  NAND2_X1 U3804 ( .A1(n4119), .A2(REG2_REG_4__SCAN_IN), .ZN(n2990) );
  OAI211_X1 U3805 ( .C1(n2992), .C2(n3265), .A(n2991), .B(n2990), .ZN(U3286)
         );
  NAND2_X1 U3806 ( .A1(n4160), .A2(n2993), .ZN(n2994) );
  INV_X1 U3807 ( .A(n2995), .ZN(n3003) );
  NAND2_X1 U3808 ( .A1(n4191), .A2(n4310), .ZN(n4141) );
  AND2_X1 U3809 ( .A1(n4191), .A2(n4298), .ZN(n4136) );
  OAI22_X1 U3810 ( .A1(n4191), .A2(n3945), .B1(REG3_REG_3__SCAN_IN), .B2(n4496), .ZN(n2996) );
  AOI21_X1 U3811 ( .B1(n4136), .B2(n3912), .A(n2996), .ZN(n3000) );
  NAND2_X1 U3812 ( .A1(n4191), .A2(n4002), .ZN(n4212) );
  INV_X1 U3813 ( .A(n2997), .ZN(n2998) );
  NAND2_X1 U3814 ( .A1(n4501), .A2(n2998), .ZN(n2999) );
  OAI211_X1 U3815 ( .C1(n4141), .C2(n3001), .A(n3000), .B(n2999), .ZN(n3002)
         );
  AOI21_X1 U3816 ( .B1(n3003), .B2(n4191), .A(n3002), .ZN(n3004) );
  OAI21_X1 U3817 ( .B1(n4216), .B2(n3005), .A(n3004), .ZN(U3287) );
  OAI22_X1 U3818 ( .A1(n3265), .A2(n3007), .B1(n3006), .B2(n4496), .ZN(n3010)
         );
  MUX2_X1 U3819 ( .A(REG2_REG_1__SCAN_IN), .B(n3008), .S(n4191), .Z(n3009) );
  AOI211_X1 U3820 ( .C1(n4135), .C2(n2815), .A(n3010), .B(n3009), .ZN(n3013)
         );
  AOI22_X1 U3821 ( .A1(n4082), .A2(n3011), .B1(n4136), .B2(n2087), .ZN(n3012)
         );
  OAI211_X1 U3822 ( .C1(n4187), .C2(n3014), .A(n3013), .B(n3012), .ZN(U3289)
         );
  XNOR2_X1 U3823 ( .A(n3015), .B(n3613), .ZN(n3106) );
  XNOR2_X1 U3824 ( .A(n3106), .B(n3105), .ZN(n3021) );
  AOI211_X1 U3825 ( .C1(n3021), .C2(n3020), .A(n3896), .B(n2081), .ZN(n3022)
         );
  INV_X1 U3826 ( .A(n3022), .ZN(n3027) );
  OAI22_X1 U3827 ( .A1(n3868), .A2(n2167), .B1(n2640), .B2(n3844), .ZN(n3025)
         );
  OAI21_X1 U3828 ( .B1(n3845), .B2(n3103), .A(n3023), .ZN(n3024) );
  NOR2_X1 U3829 ( .A1(n3025), .A2(n3024), .ZN(n3026) );
  OAI211_X1 U3830 ( .C1(n3811), .C2(n3028), .A(n3027), .B(n3026), .ZN(U3227)
         );
  MUX2_X1 U3831 ( .A(REG2_REG_2__SCAN_IN), .B(n3029), .S(n4191), .Z(n3039) );
  NOR2_X1 U3832 ( .A1(n4496), .A2(n3925), .ZN(n3030) );
  AOI21_X1 U3833 ( .B1(n3031), .B2(n4502), .A(n3030), .ZN(n3037) );
  AOI22_X1 U3834 ( .A1(n4082), .A2(n3032), .B1(n4136), .B2(n3913), .ZN(n3036)
         );
  NAND2_X1 U3835 ( .A1(n4501), .A2(n3033), .ZN(n3035) );
  NAND2_X1 U3836 ( .A1(n4135), .A2(n3914), .ZN(n3034) );
  NAND4_X1 U3837 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  OR2_X1 U3838 ( .A1(n3039), .A2(n3038), .ZN(U3288) );
  AND2_X1 U3839 ( .A1(n3521), .A2(n3517), .ZN(n3468) );
  XOR2_X1 U3840 ( .A(n3468), .B(n3040), .Z(n3085) );
  XNOR2_X1 U3841 ( .A(n3041), .B(n3468), .ZN(n3082) );
  AOI22_X1 U3842 ( .A1(n3909), .A2(n4298), .B1(n3075), .B2(n4310), .ZN(n3042)
         );
  OAI21_X1 U3843 ( .B1(n3103), .B2(n4308), .A(n3042), .ZN(n3043) );
  AOI21_X1 U3844 ( .B1(n3082), .B2(n4204), .A(n3043), .ZN(n3044) );
  OAI21_X1 U3845 ( .B1(n3085), .B2(n4321), .A(n3044), .ZN(n3050) );
  OR2_X1 U3846 ( .A1(n3060), .A2(n3118), .ZN(n3045) );
  NAND2_X1 U3847 ( .A1(n3092), .A2(n3045), .ZN(n3074) );
  INV_X1 U3848 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3046) );
  OAI22_X1 U3849 ( .A1(n4369), .A2(n3074), .B1(n4539), .B2(n3046), .ZN(n3047)
         );
  AOI21_X1 U3850 ( .B1(n3050), .B2(n4539), .A(n3047), .ZN(n3048) );
  INV_X1 U3851 ( .A(n3048), .ZN(U3479) );
  OAI22_X1 U3852 ( .A1(n4307), .A2(n3074), .B1(n4545), .B2(n2409), .ZN(n3049)
         );
  AOI21_X1 U3853 ( .B1(n3050), .B2(n4545), .A(n3049), .ZN(n3051) );
  INV_X1 U3854 ( .A(n3051), .ZN(U3524) );
  INV_X1 U3855 ( .A(n3053), .ZN(n3518) );
  AND2_X1 U3856 ( .A1(n3518), .A2(n3493), .ZN(n3465) );
  XNOR2_X1 U3857 ( .A(n3052), .B(n3465), .ZN(n3067) );
  XOR2_X1 U3858 ( .A(n3465), .B(n3054), .Z(n3055) );
  NAND2_X1 U3859 ( .A1(n3055), .A2(n4204), .ZN(n3069) );
  AOI22_X1 U3860 ( .A1(n3910), .A2(n4298), .B1(n4310), .B2(n3100), .ZN(n3056)
         );
  AOI21_X1 U3861 ( .B1(n3067), .B2(n4531), .A(n3057), .ZN(n3073) );
  AND2_X1 U3862 ( .A1(n3058), .A2(n3100), .ZN(n3059) );
  NOR2_X1 U3863 ( .A1(n3060), .A2(n3059), .ZN(n3070) );
  AOI22_X1 U3864 ( .A1(n2720), .A2(n3070), .B1(REG0_REG_5__SCAN_IN), .B2(n4537), .ZN(n3061) );
  OAI21_X1 U3865 ( .B1(n3073), .B2(n4537), .A(n3061), .ZN(U3477) );
  INV_X1 U3866 ( .A(n4191), .ZN(n4391) );
  INV_X1 U3867 ( .A(n3070), .ZN(n3065) );
  AOI22_X1 U3868 ( .A1(n4135), .A2(n3912), .B1(n4136), .B2(n3910), .ZN(n3064)
         );
  OAI22_X1 U3869 ( .A1(n4191), .A2(n2394), .B1(n3132), .B2(n4496), .ZN(n3062)
         );
  AOI21_X1 U3870 ( .B1(n3100), .B2(n4082), .A(n3062), .ZN(n3063) );
  OAI211_X1 U3871 ( .C1(n4187), .C2(n3065), .A(n3064), .B(n3063), .ZN(n3066)
         );
  AOI21_X1 U3872 ( .B1(n3067), .B2(n4132), .A(n3066), .ZN(n3068) );
  OAI21_X1 U3873 ( .B1(n3069), .B2(n4391), .A(n3068), .ZN(U3285) );
  NAND2_X1 U3874 ( .A1(n4543), .A2(REG1_REG_5__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3875 ( .A1(n2714), .A2(n3070), .ZN(n3071) );
  OAI211_X1 U3876 ( .C1(n3073), .C2(n4543), .A(n3072), .B(n3071), .ZN(U3523)
         );
  INV_X1 U3877 ( .A(n3074), .ZN(n3080) );
  INV_X1 U3878 ( .A(n4135), .ZN(n4084) );
  AOI22_X1 U3879 ( .A1(n4082), .A2(n3075), .B1(n4136), .B2(n3909), .ZN(n3078)
         );
  INV_X1 U3880 ( .A(n4191), .ZN(n4119) );
  INV_X1 U3881 ( .A(n3076), .ZN(n3120) );
  AOI22_X1 U3882 ( .A1(n4119), .A2(REG2_REG_6__SCAN_IN), .B1(n3120), .B2(n4209), .ZN(n3077) );
  OAI211_X1 U3883 ( .C1(n3103), .C2(n4084), .A(n3078), .B(n3077), .ZN(n3079)
         );
  AOI21_X1 U3884 ( .B1(n4501), .B2(n3080), .A(n3079), .ZN(n3084) );
  NAND2_X1 U3885 ( .A1(n4191), .A2(n4204), .ZN(n3251) );
  INV_X1 U3886 ( .A(n3251), .ZN(n3081) );
  NAND2_X1 U3887 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  OAI211_X1 U3888 ( .C1(n3085), .C2(n4216), .A(n3084), .B(n3083), .ZN(U3284)
         );
  XNOR2_X1 U3889 ( .A(n3086), .B(n3522), .ZN(n3089) );
  AOI22_X1 U3890 ( .A1(n3908), .A2(n4298), .B1(n4310), .B2(n3091), .ZN(n3087)
         );
  OAI21_X1 U3891 ( .B1(n3113), .B2(n4308), .A(n3087), .ZN(n3088) );
  AOI21_X1 U3892 ( .B1(n3089), .B2(n4204), .A(n3088), .ZN(n4536) );
  AOI21_X1 U3893 ( .B1(n3092), .B2(n3091), .A(n3090), .ZN(n3093) );
  NAND2_X1 U3894 ( .A1(n3093), .A2(n3154), .ZN(n4535) );
  INV_X1 U3895 ( .A(n4535), .ZN(n3096) );
  INV_X1 U3896 ( .A(n4212), .ZN(n3095) );
  OAI22_X1 U3897 ( .A1(n4191), .A2(n2416), .B1(n3167), .B2(n4496), .ZN(n3094)
         );
  AOI21_X1 U3898 ( .B1(n3096), .B2(n3095), .A(n3094), .ZN(n3099) );
  OR2_X1 U3899 ( .A1(n3097), .A2(n3522), .ZN(n4533) );
  NAND2_X1 U3900 ( .A1(n3097), .A2(n3522), .ZN(n4532) );
  NAND3_X1 U3901 ( .A1(n4533), .A2(n4532), .A3(n4132), .ZN(n3098) );
  OAI211_X1 U3902 ( .C1(n4536), .C2(n4119), .A(n3099), .B(n3098), .ZN(U3283)
         );
  OR2_X1 U3903 ( .A1(n3103), .A2(n3694), .ZN(n3102) );
  NAND2_X1 U3904 ( .A1(n3273), .A2(n3100), .ZN(n3101) );
  NAND2_X1 U3905 ( .A1(n3102), .A2(n3101), .ZN(n3111) );
  OAI22_X1 U3906 ( .A1(n3103), .A2(n3693), .B1(n2043), .B2(n3127), .ZN(n3104)
         );
  XNOR2_X1 U3907 ( .A(n3104), .B(n3695), .ZN(n3110) );
  INV_X1 U3908 ( .A(n3105), .ZN(n3108) );
  XNOR2_X1 U3909 ( .A(n3110), .B(n3111), .ZN(n3124) );
  OAI22_X1 U3910 ( .A1(n3113), .A2(n3693), .B1(n2044), .B2(n3118), .ZN(n3112)
         );
  XNOR2_X1 U3911 ( .A(n3112), .B(n3695), .ZN(n3162) );
  OAI22_X1 U3912 ( .A1(n3113), .A2(n3694), .B1(n3693), .B2(n3118), .ZN(n3163)
         );
  XNOR2_X1 U3913 ( .A(n3162), .B(n3163), .ZN(n3114) );
  XNOR2_X1 U3914 ( .A(n3164), .B(n3114), .ZN(n3122) );
  AOI21_X1 U3915 ( .B1(n3887), .B2(n3909), .A(n3115), .ZN(n3117) );
  NAND2_X1 U3916 ( .A1(n3888), .A2(n3911), .ZN(n3116) );
  OAI211_X1 U3917 ( .C1(n3868), .C2(n3118), .A(n3117), .B(n3116), .ZN(n3119)
         );
  AOI21_X1 U3918 ( .B1(n3120), .B2(n3893), .A(n3119), .ZN(n3121) );
  OAI21_X1 U3919 ( .B1(n3122), .B2(n3896), .A(n3121), .ZN(U3236) );
  AOI211_X1 U3920 ( .C1(n3125), .C2(n3124), .A(n3896), .B(n3123), .ZN(n3126)
         );
  INV_X1 U3921 ( .A(n3126), .ZN(n3131) );
  AOI211_X1 U3922 ( .C1(n3887), .C2(n3910), .A(n3129), .B(n3128), .ZN(n3130)
         );
  OAI211_X1 U3923 ( .C1(n3811), .C2(n3132), .A(n3131), .B(n3130), .ZN(U3224)
         );
  INV_X1 U3924 ( .A(n3133), .ZN(n3497) );
  AND2_X1 U3925 ( .A1(n3497), .A2(n3528), .ZN(n3470) );
  XOR2_X1 U3926 ( .A(n3470), .B(n3134), .Z(n3135) );
  NAND2_X1 U3927 ( .A1(n3135), .A2(n4204), .ZN(n3188) );
  AOI21_X1 U3928 ( .B1(n3220), .B2(n2096), .A(n3178), .ZN(n3192) );
  AOI22_X1 U3929 ( .A1(n4082), .A2(n3220), .B1(n4136), .B2(n3906), .ZN(n3136)
         );
  OAI21_X1 U3930 ( .B1(n3196), .B2(n4084), .A(n3136), .ZN(n3138) );
  OAI22_X1 U3931 ( .A1(n3224), .A2(n4496), .B1(n2445), .B2(n4191), .ZN(n3137)
         );
  AOI211_X1 U3932 ( .C1(n3192), .C2(n4501), .A(n3138), .B(n3137), .ZN(n3143)
         );
  NAND2_X1 U3933 ( .A1(n3140), .A2(n3139), .ZN(n3141) );
  XNOR2_X1 U3934 ( .A(n3141), .B(n3470), .ZN(n3190) );
  NAND2_X1 U3935 ( .A1(n3190), .A2(n4132), .ZN(n3142) );
  OAI211_X1 U3936 ( .C1(n3188), .C2(n4119), .A(n3143), .B(n3142), .ZN(U3281)
         );
  NAND2_X1 U3937 ( .A1(n4533), .A2(n3144), .ZN(n3145) );
  AND2_X1 U3938 ( .A1(n3527), .A2(n3524), .ZN(n3469) );
  XNOR2_X1 U3939 ( .A(n3145), .B(n3469), .ZN(n4503) );
  INV_X1 U3940 ( .A(n4503), .ZN(n3152) );
  XNOR2_X1 U3941 ( .A(n3146), .B(n3469), .ZN(n3149) );
  OAI22_X1 U3942 ( .A1(n3210), .A2(n4308), .B1(n3211), .B2(n4226), .ZN(n3147)
         );
  AOI21_X1 U3943 ( .B1(n4298), .B2(n3907), .A(n3147), .ZN(n3148) );
  OAI21_X1 U3944 ( .B1(n3149), .B2(n4182), .A(n3148), .ZN(n3150) );
  AOI21_X1 U3945 ( .B1(n3151), .B2(n4503), .A(n3150), .ZN(n4506) );
  OAI21_X1 U3946 ( .B1(n4523), .B2(n3152), .A(n4506), .ZN(n3157) );
  NAND2_X1 U3947 ( .A1(n3157), .A2(n4545), .ZN(n3156) );
  AOI21_X1 U3948 ( .B1(n3197), .B2(n3154), .A(n3153), .ZN(n4500) );
  NAND2_X1 U3949 ( .A1(n4500), .A2(n2714), .ZN(n3155) );
  OAI211_X1 U3950 ( .C1(n4545), .C2(n3978), .A(n3156), .B(n3155), .ZN(U3526)
         );
  INV_X1 U3951 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U3952 ( .A1(n3157), .A2(n4539), .ZN(n3159) );
  NAND2_X1 U3953 ( .A1(n4500), .A2(n2720), .ZN(n3158) );
  OAI211_X1 U3954 ( .C1(n4539), .C2(n3160), .A(n3159), .B(n3158), .ZN(U3483)
         );
  INV_X1 U3955 ( .A(n3163), .ZN(n3161) );
  OAI22_X1 U3956 ( .A1(n3210), .A2(n3694), .B1(n3693), .B2(n3171), .ZN(n3204)
         );
  OAI22_X1 U3957 ( .A1(n3210), .A2(n3693), .B1(n2043), .B2(n3171), .ZN(n3166)
         );
  XNOR2_X1 U3958 ( .A(n3166), .B(n3695), .ZN(n3205) );
  XOR2_X1 U3959 ( .A(n3204), .B(n3205), .Z(n3206) );
  XNOR2_X1 U3960 ( .A(n3207), .B(n3206), .ZN(n3175) );
  INV_X1 U3961 ( .A(n3167), .ZN(n3173) );
  AOI21_X1 U3962 ( .B1(n3887), .B2(n3908), .A(n3168), .ZN(n3170) );
  NAND2_X1 U3963 ( .A1(n3888), .A2(n3910), .ZN(n3169) );
  OAI211_X1 U3964 ( .C1(n3868), .C2(n3171), .A(n3170), .B(n3169), .ZN(n3172)
         );
  AOI21_X1 U3965 ( .B1(n3173), .B2(n3893), .A(n3172), .ZN(n3174) );
  OAI21_X1 U3966 ( .B1(n3175), .B2(n3896), .A(n3174), .ZN(U3210) );
  AND2_X1 U3967 ( .A1(n3496), .A2(n3492), .ZN(n3466) );
  XOR2_X1 U3968 ( .A(n3466), .B(n3176), .Z(n3234) );
  XOR2_X1 U3969 ( .A(n3466), .B(n3177), .Z(n3236) );
  NAND2_X1 U3970 ( .A1(n3236), .A2(n4132), .ZN(n3186) );
  INV_X1 U3971 ( .A(n3178), .ZN(n3180) );
  INV_X1 U3972 ( .A(n3179), .ZN(n3260) );
  AOI21_X1 U3973 ( .B1(n3274), .B2(n3180), .A(n3260), .ZN(n3238) );
  AOI22_X1 U3974 ( .A1(n4082), .A2(n3274), .B1(n4136), .B2(n3905), .ZN(n3183)
         );
  INV_X1 U3975 ( .A(n3289), .ZN(n3181) );
  AOI22_X1 U3976 ( .A1(n4119), .A2(REG2_REG_10__SCAN_IN), .B1(n3181), .B2(
        n4209), .ZN(n3182) );
  OAI211_X1 U3977 ( .C1(n3283), .C2(n4084), .A(n3183), .B(n3182), .ZN(n3184)
         );
  AOI21_X1 U3978 ( .B1(n3238), .B2(n4501), .A(n3184), .ZN(n3185) );
  OAI211_X1 U3979 ( .C1(n3234), .C2(n3251), .A(n3186), .B(n3185), .ZN(U3280)
         );
  AOI22_X1 U3980 ( .A1(n3906), .A2(n4298), .B1(n4310), .B2(n3220), .ZN(n3187)
         );
  OAI211_X1 U3981 ( .C1(n3196), .C2(n4308), .A(n3188), .B(n3187), .ZN(n3189)
         );
  AOI21_X1 U3982 ( .B1(n3190), .B2(n4531), .A(n3189), .ZN(n3194) );
  AOI22_X1 U3983 ( .A1(n3192), .A2(n2714), .B1(REG1_REG_9__SCAN_IN), .B2(n4543), .ZN(n3191) );
  OAI21_X1 U3984 ( .B1(n3194), .B2(n4543), .A(n3191), .ZN(U3527) );
  AOI22_X1 U3985 ( .A1(n3192), .A2(n2720), .B1(REG0_REG_9__SCAN_IN), .B2(n4537), .ZN(n3193) );
  OAI21_X1 U3986 ( .B1(n3194), .B2(n4537), .A(n3193), .ZN(U3485) );
  OAI22_X1 U3987 ( .A1(n3196), .A2(n3693), .B1(n2043), .B2(n3211), .ZN(n3195)
         );
  XNOR2_X1 U3988 ( .A(n3195), .B(n3695), .ZN(n3200) );
  OR2_X1 U3989 ( .A1(n3196), .A2(n3694), .ZN(n3199) );
  NAND2_X1 U3990 ( .A1(n3273), .A2(n3197), .ZN(n3198) );
  NAND2_X1 U3991 ( .A1(n3199), .A2(n3198), .ZN(n3201) );
  NAND2_X1 U3992 ( .A1(n3200), .A2(n3201), .ZN(n3217) );
  INV_X1 U3993 ( .A(n3200), .ZN(n3203) );
  INV_X1 U3994 ( .A(n3201), .ZN(n3202) );
  NAND2_X1 U3995 ( .A1(n3203), .A2(n3202), .ZN(n3219) );
  NAND2_X1 U3996 ( .A1(n3217), .A2(n3219), .ZN(n3208) );
  XOR2_X1 U3997 ( .A(n3208), .B(n3218), .Z(n3209) );
  NAND2_X1 U3998 ( .A1(n3209), .A2(n3764), .ZN(n3216) );
  OAI22_X1 U3999 ( .A1(n3868), .A2(n3211), .B1(n3210), .B2(n3844), .ZN(n3214)
         );
  OAI21_X1 U4000 ( .B1(n3845), .B2(n3283), .A(n3212), .ZN(n3213) );
  NOR2_X1 U4001 ( .A1(n3214), .A2(n3213), .ZN(n3215) );
  OAI211_X1 U4002 ( .C1(n3811), .C2(n4497), .A(n3216), .B(n3215), .ZN(U3218)
         );
  OAI22_X1 U4003 ( .A1(n3283), .A2(n3694), .B1(n3693), .B2(n3227), .ZN(n3268)
         );
  NAND2_X1 U4004 ( .A1(n3907), .A2(n3273), .ZN(n3222) );
  NAND2_X1 U4005 ( .A1(n2045), .A2(n3220), .ZN(n3221) );
  NAND2_X1 U4006 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  XNOR2_X1 U4007 ( .A(n3223), .B(n3695), .ZN(n3269) );
  XOR2_X1 U4008 ( .A(n3267), .B(n3266), .Z(n3231) );
  INV_X1 U4009 ( .A(n3224), .ZN(n3229) );
  AND2_X1 U4010 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4404) );
  AOI21_X1 U4011 ( .B1(n3887), .B2(n3906), .A(n4404), .ZN(n3226) );
  NAND2_X1 U4012 ( .A1(n3888), .A2(n3908), .ZN(n3225) );
  OAI211_X1 U4013 ( .C1(n3868), .C2(n3227), .A(n3226), .B(n3225), .ZN(n3228)
         );
  AOI21_X1 U4014 ( .B1(n3229), .B2(n3893), .A(n3228), .ZN(n3230) );
  OAI21_X1 U4015 ( .B1(n3231), .B2(n3896), .A(n3230), .ZN(U3228) );
  OAI22_X1 U4016 ( .A1(n3766), .A2(n4314), .B1(n4226), .B2(n3284), .ZN(n3232)
         );
  AOI21_X1 U4017 ( .B1(n4277), .B2(n3907), .A(n3232), .ZN(n3233) );
  OAI21_X1 U4018 ( .B1(n3234), .B2(n4182), .A(n3233), .ZN(n3235) );
  AOI21_X1 U4019 ( .B1(n4531), .B2(n3236), .A(n3235), .ZN(n3240) );
  AOI22_X1 U4020 ( .A1(n3238), .A2(n2714), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4543), .ZN(n3237) );
  OAI21_X1 U4021 ( .B1(n3240), .B2(n4543), .A(n3237), .ZN(U3528) );
  AOI22_X1 U4022 ( .A1(n3238), .A2(n2720), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4537), .ZN(n3239) );
  OAI21_X1 U4023 ( .B1(n3240), .B2(n4537), .A(n3239), .ZN(U3487) );
  XNOR2_X1 U4024 ( .A(n3425), .B(n3242), .ZN(n3361) );
  OAI21_X1 U4025 ( .B1(n3243), .B2(n3242), .A(n3241), .ZN(n3363) );
  NAND2_X1 U4026 ( .A1(n3363), .A2(n4132), .ZN(n3250) );
  OAI21_X1 U4027 ( .B1(n3302), .B2(n3724), .A(n3337), .ZN(n3369) );
  INV_X1 U4028 ( .A(n3369), .ZN(n3248) );
  AOI22_X1 U4029 ( .A1(n4082), .A2(n3609), .B1(n4136), .B2(n3901), .ZN(n3246)
         );
  INV_X1 U4030 ( .A(n3730), .ZN(n3244) );
  AOI22_X1 U4031 ( .A1(n4119), .A2(REG2_REG_14__SCAN_IN), .B1(n3244), .B2(
        n4209), .ZN(n3245) );
  OAI211_X1 U4032 ( .C1(n3768), .C2(n4084), .A(n3246), .B(n3245), .ZN(n3247)
         );
  AOI21_X1 U4033 ( .B1(n3248), .B2(n4501), .A(n3247), .ZN(n3249) );
  OAI211_X1 U4034 ( .C1(n3361), .C2(n3251), .A(n3250), .B(n3249), .ZN(U3276)
         );
  INV_X1 U4035 ( .A(n3252), .ZN(n3253) );
  AOI21_X1 U4036 ( .B1(n3447), .B2(n3254), .A(n3253), .ZN(n3324) );
  AOI22_X1 U4037 ( .A1(n3904), .A2(n4298), .B1(n4310), .B2(n3255), .ZN(n3258)
         );
  XNOR2_X1 U4038 ( .A(n3293), .B(n3447), .ZN(n3256) );
  NAND2_X1 U4039 ( .A1(n3256), .A2(n4204), .ZN(n3257) );
  OAI211_X1 U4040 ( .C1(n3324), .C2(n4160), .A(n3258), .B(n3257), .ZN(n3326)
         );
  NAND2_X1 U4041 ( .A1(n3326), .A2(n4191), .ZN(n3264) );
  OAI22_X1 U4042 ( .A1(n4191), .A2(n3259), .B1(n3854), .B2(n4496), .ZN(n3262)
         );
  OAI21_X1 U40430 ( .B1(n3260), .B2(n3857), .A(n3311), .ZN(n3332) );
  NOR2_X1 U4044 ( .A1(n3332), .A2(n4187), .ZN(n3261) );
  AOI211_X1 U4045 ( .C1(n4135), .C2(n3906), .A(n3262), .B(n3261), .ZN(n3263)
         );
  OAI211_X1 U4046 ( .C1(n3324), .C2(n3265), .A(n3264), .B(n3263), .ZN(U3279)
         );
  NAND2_X1 U4047 ( .A1(n3267), .A2(n3266), .ZN(n3271) );
  NOR2_X1 U4048 ( .A1(n3693), .A2(n3284), .ZN(n3272) );
  AOI21_X1 U4049 ( .B1(n2816), .B2(n3906), .A(n3272), .ZN(n3588) );
  NAND2_X1 U4050 ( .A1(n3906), .A2(n3273), .ZN(n3276) );
  NAND2_X1 U4051 ( .A1(n2045), .A2(n3274), .ZN(n3275) );
  NAND2_X1 U4052 ( .A1(n3276), .A2(n3275), .ZN(n3277) );
  XNOR2_X1 U4053 ( .A(n3277), .B(n3695), .ZN(n3590) );
  XOR2_X1 U4054 ( .A(n3588), .B(n3590), .Z(n3279) );
  AOI21_X1 U4055 ( .B1(n3278), .B2(n3279), .A(n3896), .ZN(n3282) );
  NAND2_X1 U4056 ( .A1(n3282), .A2(n3592), .ZN(n3288) );
  OAI22_X1 U4057 ( .A1(n3868), .A2(n3284), .B1(n3283), .B2(n3844), .ZN(n3286)
         );
  NAND2_X1 U4058 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4408) );
  OAI21_X1 U4059 ( .B1(n3845), .B2(n3766), .A(n4408), .ZN(n3285) );
  NOR2_X1 U4060 ( .A1(n3286), .A2(n3285), .ZN(n3287) );
  OAI211_X1 U4061 ( .C1(n3811), .C2(n3289), .A(n3288), .B(n3287), .ZN(U3214)
         );
  INV_X1 U4062 ( .A(n3290), .ZN(n3291) );
  AOI21_X1 U4063 ( .B1(n3293), .B2(n3292), .A(n3291), .ZN(n3318) );
  INV_X1 U4064 ( .A(n3309), .ZN(n3294) );
  AOI21_X1 U4065 ( .B1(n3318), .B2(n3310), .A(n3294), .ZN(n3296) );
  XNOR2_X1 U4066 ( .A(n3768), .B(n3295), .ZN(n3459) );
  XNOR2_X1 U4067 ( .A(n3296), .B(n3459), .ZN(n3299) );
  OAI22_X1 U4068 ( .A1(n3608), .A2(n4314), .B1(n4226), .B2(n3835), .ZN(n3297)
         );
  AOI21_X1 U4069 ( .B1(n4277), .B2(n3904), .A(n3297), .ZN(n3298) );
  OAI21_X1 U4070 ( .B1(n3299), .B2(n4182), .A(n3298), .ZN(n3370) );
  INV_X1 U4071 ( .A(n3370), .ZN(n3307) );
  XNOR2_X1 U4072 ( .A(n3300), .B(n3459), .ZN(n3371) );
  NOR2_X1 U4073 ( .A1(n3312), .A2(n3835), .ZN(n3301) );
  OR2_X1 U4074 ( .A1(n3302), .A2(n3301), .ZN(n3377) );
  INV_X1 U4075 ( .A(n3303), .ZN(n3837) );
  AOI22_X1 U4076 ( .A1(n4119), .A2(REG2_REG_13__SCAN_IN), .B1(n3837), .B2(
        n4209), .ZN(n3304) );
  OAI21_X1 U4077 ( .B1(n3377), .B2(n4187), .A(n3304), .ZN(n3305) );
  AOI21_X1 U4078 ( .B1(n3371), .B2(n4132), .A(n3305), .ZN(n3306) );
  OAI21_X1 U4079 ( .B1(n3307), .B2(n4391), .A(n3306), .ZN(U3277) );
  NAND2_X1 U4080 ( .A1(n3310), .A2(n3309), .ZN(n3463) );
  XNOR2_X1 U4081 ( .A(n3308), .B(n3463), .ZN(n3346) );
  AND2_X1 U4082 ( .A1(n3311), .A2(n3596), .ZN(n3313) );
  OR2_X1 U4083 ( .A1(n3313), .A2(n3312), .ZN(n3358) );
  OAI22_X1 U4084 ( .A1(n4191), .A2(n3314), .B1(n3773), .B2(n4496), .ZN(n3315)
         );
  AOI21_X1 U4085 ( .B1(n3596), .B2(n4082), .A(n3315), .ZN(n3317) );
  AOI22_X1 U4086 ( .A1(n4135), .A2(n3905), .B1(n4136), .B2(n3903), .ZN(n3316)
         );
  OAI211_X1 U4087 ( .C1(n3358), .C2(n4187), .A(n3317), .B(n3316), .ZN(n3321)
         );
  XNOR2_X1 U4088 ( .A(n3318), .B(n3463), .ZN(n3319) );
  NAND2_X1 U4089 ( .A1(n3319), .A2(n4204), .ZN(n3350) );
  NOR2_X1 U4090 ( .A1(n3350), .A2(n4119), .ZN(n3320) );
  AOI211_X1 U4091 ( .C1(n4132), .C2(n3346), .A(n3321), .B(n3320), .ZN(n3322)
         );
  INV_X1 U4092 ( .A(n3322), .ZN(U3278) );
  OAI22_X1 U4093 ( .A1(n3324), .A2(n4523), .B1(n3323), .B2(n4308), .ZN(n3325)
         );
  NOR2_X1 U4094 ( .A1(n3326), .A2(n3325), .ZN(n3329) );
  MUX2_X1 U4095 ( .A(n3327), .B(n3329), .S(n4545), .Z(n3328) );
  OAI21_X1 U4096 ( .B1(n4307), .B2(n3332), .A(n3328), .ZN(U3529) );
  INV_X1 U4097 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3330) );
  MUX2_X1 U4098 ( .A(n3330), .B(n3329), .S(n4539), .Z(n3331) );
  OAI21_X1 U4099 ( .B1(n3332), .B2(n4369), .A(n3331), .ZN(U3489) );
  AOI21_X1 U4100 ( .B1(n3333), .B2(n3446), .A(n4182), .ZN(n3335) );
  NAND2_X1 U4101 ( .A1(n3335), .A2(n3334), .ZN(n3379) );
  XNOR2_X1 U4102 ( .A(n3336), .B(n3446), .ZN(n3381) );
  NAND2_X1 U4103 ( .A1(n3381), .A2(n4132), .ZN(n3345) );
  INV_X1 U4104 ( .A(n3337), .ZN(n3338) );
  OAI21_X1 U4105 ( .B1(n3338), .B2(n3891), .A(n3572), .ZN(n3387) );
  INV_X1 U4106 ( .A(n3387), .ZN(n3343) );
  AOI22_X1 U4107 ( .A1(n4136), .A2(n3900), .B1(n4135), .B2(n3902), .ZN(n3341)
         );
  INV_X1 U4108 ( .A(n3339), .ZN(n3894) );
  AOI22_X1 U4109 ( .A1(n4119), .A2(REG2_REG_15__SCAN_IN), .B1(n3894), .B2(
        n4209), .ZN(n3340) );
  OAI211_X1 U4110 ( .C1(n3891), .C2(n4141), .A(n3341), .B(n3340), .ZN(n3342)
         );
  AOI21_X1 U4111 ( .B1(n3343), .B2(n4501), .A(n3342), .ZN(n3344) );
  OAI211_X1 U4112 ( .C1(n4119), .C2(n3379), .A(n3345), .B(n3344), .ZN(U3275)
         );
  INV_X1 U4113 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4114 ( .A1(n3346), .A2(n4531), .ZN(n3352) );
  OR2_X1 U4115 ( .A1(n3766), .A2(n4308), .ZN(n3348) );
  NAND2_X1 U4116 ( .A1(n3596), .A2(n4310), .ZN(n3347) );
  OAI211_X1 U4117 ( .C1(n3768), .C2(n4314), .A(n3348), .B(n3347), .ZN(n3349)
         );
  INV_X1 U4118 ( .A(n3349), .ZN(n3351) );
  MUX2_X1 U4119 ( .A(n3353), .B(n3355), .S(n4539), .Z(n3354) );
  OAI21_X1 U4120 ( .B1(n3358), .B2(n4369), .A(n3354), .ZN(U3491) );
  MUX2_X1 U4121 ( .A(n3356), .B(n3355), .S(n4545), .Z(n3357) );
  OAI21_X1 U4122 ( .B1(n4307), .B2(n3358), .A(n3357), .ZN(U3530) );
  OAI22_X1 U4123 ( .A1(n4309), .A2(n4314), .B1(n4226), .B2(n3724), .ZN(n3359)
         );
  AOI21_X1 U4124 ( .B1(n4277), .B2(n3903), .A(n3359), .ZN(n3360) );
  OAI21_X1 U4125 ( .B1(n3361), .B2(n4182), .A(n3360), .ZN(n3362) );
  AOI21_X1 U4126 ( .B1(n3363), .B2(n4531), .A(n3362), .ZN(n3366) );
  MUX2_X1 U4127 ( .A(n3364), .B(n3366), .S(n4545), .Z(n3365) );
  OAI21_X1 U4128 ( .B1(n4307), .B2(n3369), .A(n3365), .ZN(U3532) );
  INV_X1 U4129 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3367) );
  MUX2_X1 U4130 ( .A(n3367), .B(n3366), .S(n4539), .Z(n3368) );
  OAI21_X1 U4131 ( .B1(n3369), .B2(n4369), .A(n3368), .ZN(U3495) );
  AOI21_X1 U4132 ( .B1(n4531), .B2(n3371), .A(n3370), .ZN(n3374) );
  MUX2_X1 U4133 ( .A(n3372), .B(n3374), .S(n4545), .Z(n3373) );
  OAI21_X1 U4134 ( .B1(n4307), .B2(n3377), .A(n3373), .ZN(U3531) );
  INV_X1 U4135 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3375) );
  MUX2_X1 U4136 ( .A(n3375), .B(n3374), .S(n4539), .Z(n3376) );
  OAI21_X1 U4137 ( .B1(n3377), .B2(n4369), .A(n3376), .ZN(U3493) );
  AOI22_X1 U4138 ( .A1(n3900), .A2(n4298), .B1(n3618), .B2(n4310), .ZN(n3378)
         );
  OAI211_X1 U4139 ( .C1(n3608), .C2(n4308), .A(n3379), .B(n3378), .ZN(n3380)
         );
  AOI21_X1 U4140 ( .B1(n3381), .B2(n4531), .A(n3380), .ZN(n3384) );
  MUX2_X1 U4141 ( .A(n3382), .B(n3384), .S(n4545), .Z(n3383) );
  OAI21_X1 U4142 ( .B1(n4307), .B2(n3387), .A(n3383), .ZN(U3533) );
  INV_X1 U4143 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3385) );
  MUX2_X1 U4144 ( .A(n3385), .B(n3384), .S(n4539), .Z(n3386) );
  OAI21_X1 U4145 ( .B1(n3387), .B2(n4369), .A(n3386), .ZN(U3497) );
  INV_X1 U4146 ( .A(n3388), .ZN(n3418) );
  NAND2_X1 U4147 ( .A1(n3418), .A2(n4172), .ZN(n3464) );
  XNOR2_X1 U4148 ( .A(n3389), .B(n3464), .ZN(n3390) );
  NAND2_X1 U4149 ( .A1(n3390), .A2(n4204), .ZN(n4301) );
  XOR2_X1 U4150 ( .A(n3464), .B(n3391), .Z(n4304) );
  NAND2_X1 U4151 ( .A1(n4304), .A2(n4132), .ZN(n3400) );
  INV_X1 U4152 ( .A(n3574), .ZN(n3393) );
  INV_X1 U4153 ( .A(n4208), .ZN(n3392) );
  OAI21_X1 U4154 ( .B1(n3393), .B2(n3802), .A(n3392), .ZN(n4375) );
  INV_X1 U4155 ( .A(n4375), .ZN(n3398) );
  AOI22_X1 U4156 ( .A1(n4135), .A2(n3900), .B1(n4136), .B2(n4299), .ZN(n3396)
         );
  INV_X1 U4157 ( .A(n3394), .ZN(n3804) );
  AOI22_X1 U4158 ( .A1(n4119), .A2(REG2_REG_17__SCAN_IN), .B1(n3804), .B2(
        n4209), .ZN(n3395) );
  OAI211_X1 U4159 ( .C1(n3802), .C2(n4141), .A(n3396), .B(n3395), .ZN(n3397)
         );
  AOI21_X1 U4160 ( .B1(n3398), .B2(n4501), .A(n3397), .ZN(n3399) );
  OAI211_X1 U4161 ( .C1(n4119), .C2(n4301), .A(n3400), .B(n3399), .ZN(U3273)
         );
  INV_X1 U4162 ( .A(n3898), .ZN(n3403) );
  INV_X1 U4163 ( .A(DATAI_30_), .ZN(n3401) );
  NOR2_X1 U4164 ( .A1(n3402), .A2(n3401), .ZN(n4223) );
  NOR2_X1 U4165 ( .A1(n3403), .A2(n4223), .ZN(n3554) );
  INV_X1 U4166 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4217) );
  NAND2_X1 U4167 ( .A1(n2361), .A2(REG2_REG_31__SCAN_IN), .ZN(n3406) );
  NAND2_X1 U4168 ( .A1(n3404), .A2(REG0_REG_31__SCAN_IN), .ZN(n3405) );
  OAI211_X1 U4169 ( .C1(n3407), .C2(n4217), .A(n3406), .B(n3405), .ZN(n4008)
         );
  INV_X1 U4170 ( .A(n4008), .ZN(n3408) );
  NOR2_X1 U4171 ( .A1(n3554), .A2(n3408), .ZN(n3443) );
  NAND2_X1 U4172 ( .A1(n2305), .A2(DATAI_31_), .ZN(n4009) );
  INV_X1 U4173 ( .A(n4223), .ZN(n3454) );
  INV_X1 U4174 ( .A(n4229), .ZN(n3702) );
  OAI21_X1 U4175 ( .B1(n3702), .B2(n3410), .A(n3409), .ZN(n3549) );
  NOR3_X1 U4176 ( .A1(n3549), .A2(n4025), .A3(n3411), .ZN(n3438) );
  NAND2_X1 U4177 ( .A1(n3413), .A2(n3412), .ZN(n3434) );
  INV_X1 U4178 ( .A(n3434), .ZN(n3416) );
  NAND2_X1 U4179 ( .A1(n4008), .A2(n4009), .ZN(n3552) );
  OR2_X1 U4180 ( .A1(n3898), .A2(n3454), .ZN(n3414) );
  OAI211_X1 U4181 ( .C1(n4229), .C2(n4014), .A(n3552), .B(n3414), .ZN(n3433)
         );
  INV_X1 U4182 ( .A(n3433), .ZN(n3415) );
  OAI21_X1 U4183 ( .B1(n3416), .B2(n3549), .A(n3415), .ZN(n3556) );
  NAND2_X1 U4184 ( .A1(n3417), .A2(n3424), .ZN(n3537) );
  NAND2_X1 U4185 ( .A1(n3498), .A2(n3499), .ZN(n3423) );
  INV_X1 U4186 ( .A(n3500), .ZN(n3422) );
  NAND2_X1 U4187 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  OR2_X1 U4188 ( .A1(n3421), .A2(n3420), .ZN(n3502) );
  AOI211_X1 U4189 ( .C1(n3424), .C2(n3423), .A(n3422), .B(n3502), .ZN(n3536)
         );
  OAI21_X1 U4190 ( .B1(n3425), .B2(n3537), .A(n3536), .ZN(n3429) );
  INV_X1 U4191 ( .A(n3502), .ZN(n3428) );
  INV_X1 U4192 ( .A(n3426), .ZN(n3427) );
  NAND2_X1 U4193 ( .A1(n3428), .A2(n3427), .ZN(n3540) );
  NAND4_X1 U4194 ( .A1(n3429), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3432)
         );
  INV_X1 U4195 ( .A(n3485), .ZN(n3430) );
  NAND2_X1 U4196 ( .A1(n3430), .A2(n3451), .ZN(n3545) );
  AOI21_X1 U4197 ( .B1(n3432), .B2(n3431), .A(n3545), .ZN(n3436) );
  NOR3_X1 U4198 ( .A1(n3434), .A2(n3544), .A3(n3433), .ZN(n3435) );
  OAI21_X1 U4199 ( .B1(n3436), .B2(n4045), .A(n3435), .ZN(n3437) );
  OAI21_X1 U4200 ( .B1(n3438), .B2(n3556), .A(n3437), .ZN(n3439) );
  OAI21_X1 U4201 ( .B1(n4008), .B2(n3454), .A(n3439), .ZN(n3442) );
  INV_X1 U4202 ( .A(n3440), .ZN(n3441) );
  OAI211_X1 U4203 ( .C1(n3443), .C2(n4009), .A(n3442), .B(n3441), .ZN(n3561)
         );
  XNOR2_X1 U4204 ( .A(n4252), .B(n4053), .ZN(n4042) );
  INV_X1 U4205 ( .A(n4042), .ZN(n4047) );
  NOR2_X1 U4206 ( .A1(n3711), .A2(n4047), .ZN(n3490) );
  INV_X1 U4207 ( .A(n3444), .ZN(n3489) );
  INV_X1 U4208 ( .A(n3445), .ZN(n4094) );
  OR2_X1 U4209 ( .A1(n4093), .A2(n4094), .ZN(n4131) );
  INV_X1 U4210 ( .A(n3446), .ZN(n3448) );
  NAND4_X1 U4211 ( .A1(n3448), .A2(n3447), .A3(n3522), .A4(n4524), .ZN(n3449)
         );
  NOR3_X1 U4212 ( .A1(n4131), .A2(n4121), .A3(n3449), .ZN(n3483) );
  NAND2_X1 U4213 ( .A1(n3451), .A2(n3450), .ZN(n4097) );
  INV_X1 U4214 ( .A(n4097), .ZN(n3482) );
  NAND2_X1 U4215 ( .A1(n3453), .A2(n3452), .ZN(n4178) );
  XNOR2_X1 U4216 ( .A(n3898), .B(n3454), .ZN(n3458) );
  NOR2_X1 U4217 ( .A1(n4008), .A2(n4009), .ZN(n3553) );
  INV_X1 U4218 ( .A(n3553), .ZN(n3456) );
  NAND3_X1 U4219 ( .A1(n3456), .A2(n3552), .A3(n3455), .ZN(n3457) );
  NOR4_X1 U4220 ( .A1(n4178), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n3481)
         );
  INV_X1 U4221 ( .A(n3460), .ZN(n3461) );
  OR2_X1 U4222 ( .A1(n3462), .A2(n3461), .ZN(n4151) );
  NOR2_X1 U4223 ( .A1(n3464), .A2(n3463), .ZN(n3479) );
  AND4_X1 U4224 ( .A1(n2171), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3478)
         );
  NAND4_X1 U4225 ( .A1(n3470), .A2(n3579), .A3(n3469), .A4(n3468), .ZN(n3476)
         );
  INV_X1 U4226 ( .A(n2638), .ZN(n3474) );
  NAND4_X1 U4227 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3475)
         );
  NOR2_X1 U4228 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  AND4_X1 U4229 ( .A1(n4151), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3480)
         );
  NAND4_X1 U4230 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3487)
         );
  NAND2_X1 U4231 ( .A1(n4044), .A2(n3484), .ZN(n4064) );
  INV_X1 U4232 ( .A(n4059), .ZN(n3486) );
  OR2_X1 U4233 ( .A1(n3486), .A2(n3485), .ZN(n4077) );
  NOR3_X1 U4234 ( .A1(n3487), .A2(n4064), .A3(n4077), .ZN(n3488) );
  NAND4_X1 U4235 ( .A1(n3490), .A2(n3489), .A3(n2153), .A4(n3488), .ZN(n3559)
         );
  INV_X1 U4236 ( .A(n3491), .ZN(n3547) );
  NOR2_X1 U4237 ( .A1(n2163), .A2(n3493), .ZN(n3494) );
  NAND4_X1 U4238 ( .A1(n3494), .A2(n3497), .A3(n3524), .A4(n3517), .ZN(n3495)
         );
  NAND2_X1 U4239 ( .A1(n3496), .A2(n3495), .ZN(n3531) );
  NAND4_X1 U4240 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  NOR2_X1 U4241 ( .A1(n3502), .A2(n3501), .ZN(n3530) );
  INV_X1 U4242 ( .A(n3504), .ZN(n3507) );
  OAI211_X1 U4243 ( .C1(n4380), .C2(n3507), .A(n3506), .B(n3505), .ZN(n3508)
         );
  NAND3_X1 U4244 ( .A1(n3510), .A2(n3509), .A3(n3508), .ZN(n3511) );
  NAND3_X1 U4245 ( .A1(n3503), .A2(n3512), .A3(n3511), .ZN(n3513) );
  NAND3_X1 U4246 ( .A1(n3515), .A2(n3514), .A3(n3513), .ZN(n3516) );
  NAND4_X1 U4247 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3520)
         );
  NAND3_X1 U4248 ( .A1(n3522), .A2(n3521), .A3(n3520), .ZN(n3523) );
  NAND3_X1 U4249 ( .A1(n3525), .A2(n3524), .A3(n3523), .ZN(n3526) );
  NAND3_X1 U4250 ( .A1(n3528), .A2(n3527), .A3(n3526), .ZN(n3529) );
  AOI22_X1 U4251 ( .A1(n3536), .A2(n3531), .B1(n3530), .B2(n3529), .ZN(n3533)
         );
  OR4_X1 U4252 ( .A1(n3534), .A2(n2147), .A3(n3533), .A4(n3532), .ZN(n3539) );
  OAI21_X1 U4253 ( .B1(n2142), .B2(n3537), .A(n3536), .ZN(n3538) );
  AND4_X1 U4254 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3543)
         );
  OAI21_X1 U4255 ( .B1(n4093), .B2(n3543), .A(n3542), .ZN(n3546) );
  AOI211_X1 U4256 ( .C1(n3547), .C2(n3546), .A(n3545), .B(n3544), .ZN(n3548)
         );
  AOI211_X1 U4257 ( .C1(n3899), .C2(n4031), .A(n3549), .B(n3548), .ZN(n3551)
         );
  AND2_X1 U4258 ( .A1(n3551), .A2(n3550), .ZN(n3557) );
  OAI21_X1 U4259 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n3555) );
  OAI21_X1 U4260 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3558) );
  MUX2_X1 U4261 ( .A(n3559), .B(n3558), .S(n2637), .Z(n3560) );
  NAND2_X1 U4262 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  XNOR2_X1 U4263 ( .A(n3562), .B(n4381), .ZN(n3568) );
  NAND2_X1 U4264 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  OAI211_X1 U4265 ( .C1(n4379), .C2(n3567), .A(n3565), .B(B_REG_SCAN_IN), .ZN(
        n3566) );
  OAI21_X1 U4266 ( .B1(n3568), .B2(n3567), .A(n3566), .ZN(U3239) );
  OAI21_X1 U4267 ( .B1(n3571), .B2(n3570), .A(n3569), .ZN(n4322) );
  NAND2_X1 U4268 ( .A1(n3572), .A2(n4311), .ZN(n3573) );
  AND2_X1 U4269 ( .A1(n3574), .A2(n3573), .ZN(n4318) );
  AOI22_X1 U4270 ( .A1(n4135), .A2(n3901), .B1(n4136), .B2(n4200), .ZN(n3577)
         );
  INV_X1 U4271 ( .A(n3575), .ZN(n3793) );
  AOI22_X1 U4272 ( .A1(n4391), .A2(REG2_REG_16__SCAN_IN), .B1(n3793), .B2(
        n4209), .ZN(n3576) );
  OAI211_X1 U4273 ( .C1(n3791), .C2(n4141), .A(n3577), .B(n3576), .ZN(n3582)
         );
  OAI211_X1 U4274 ( .C1(n3580), .C2(n3579), .A(n3578), .B(n4204), .ZN(n4319)
         );
  NOR2_X1 U4275 ( .A1(n4319), .A2(n4119), .ZN(n3581) );
  AOI211_X1 U4276 ( .C1(n4318), .C2(n4501), .A(n3582), .B(n3581), .ZN(n3583)
         );
  OAI21_X1 U4277 ( .B1(n4322), .B2(n4216), .A(n3583), .ZN(U3274) );
  INV_X1 U4278 ( .A(D_REG_0__SCAN_IN), .ZN(n3587) );
  NOR2_X1 U4279 ( .A1(n4508), .A2(n3584), .ZN(n3586) );
  AOI22_X1 U4280 ( .A1(n4507), .A2(n3587), .B1(n3586), .B2(n3585), .ZN(U3458)
         );
  INV_X1 U4281 ( .A(n3588), .ZN(n3589) );
  NAND2_X1 U4282 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  OAI22_X1 U4283 ( .A1(n3766), .A2(n3694), .B1(n3693), .B2(n3857), .ZN(n3852)
         );
  OAI22_X1 U4284 ( .A1(n3766), .A2(n3693), .B1(n2043), .B2(n3857), .ZN(n3593)
         );
  XNOR2_X1 U4285 ( .A(n3593), .B(n3695), .ZN(n3851) );
  OAI22_X1 U4286 ( .A1(n3595), .A2(n3693), .B1(n2044), .B2(n3767), .ZN(n3594)
         );
  XNOR2_X1 U4287 ( .A(n3594), .B(n2055), .ZN(n3602) );
  INV_X1 U4288 ( .A(n3602), .ZN(n3599) );
  OR2_X1 U4289 ( .A1(n3595), .A2(n3694), .ZN(n3598) );
  NAND2_X1 U4290 ( .A1(n3273), .A2(n3596), .ZN(n3597) );
  NAND2_X1 U4291 ( .A1(n3598), .A2(n3597), .ZN(n3600) );
  NAND2_X1 U4292 ( .A1(n3599), .A2(n3600), .ZN(n3759) );
  INV_X1 U4293 ( .A(n3600), .ZN(n3601) );
  INV_X1 U4294 ( .A(n3829), .ZN(n3606) );
  OAI22_X1 U4295 ( .A1(n3768), .A2(n3693), .B1(n2044), .B2(n3835), .ZN(n3603)
         );
  XNOR2_X1 U4296 ( .A(n3603), .B(n3695), .ZN(n3604) );
  INV_X1 U4297 ( .A(n3604), .ZN(n3831) );
  OAI22_X1 U4298 ( .A1(n3768), .A2(n3694), .B1(n3693), .B2(n3835), .ZN(n3830)
         );
  OAI22_X1 U4299 ( .A1(n3608), .A2(n3693), .B1(n2043), .B2(n3724), .ZN(n3607)
         );
  XNOR2_X1 U4300 ( .A(n3607), .B(n3695), .ZN(n3615) );
  OR2_X1 U4301 ( .A1(n3608), .A2(n3694), .ZN(n3611) );
  NAND2_X1 U4302 ( .A1(n3273), .A2(n3609), .ZN(n3610) );
  NAND2_X1 U4303 ( .A1(n3611), .A2(n3610), .ZN(n3614) );
  OAI22_X1 U4304 ( .A1(n4309), .A2(n3693), .B1(n2043), .B2(n3891), .ZN(n3612)
         );
  XNOR2_X1 U4305 ( .A(n3613), .B(n3612), .ZN(n3621) );
  OAI21_X2 U4306 ( .B1(n3617), .B2(n3719), .A(n3616), .ZN(n3884) );
  OR2_X1 U4307 ( .A1(n4309), .A2(n3694), .ZN(n3620) );
  NAND2_X1 U4308 ( .A1(n3273), .A2(n3618), .ZN(n3619) );
  NAND2_X1 U4309 ( .A1(n3620), .A2(n3619), .ZN(n3886) );
  OR2_X1 U4310 ( .A1(n3621), .A2(n3720), .ZN(n3784) );
  AND2_X1 U4311 ( .A1(n3886), .A2(n3784), .ZN(n3622) );
  OAI22_X1 U4312 ( .A1(n4302), .A2(n3694), .B1(n3693), .B2(n3791), .ZN(n3625)
         );
  OAI22_X1 U4313 ( .A1(n4302), .A2(n3693), .B1(n2044), .B2(n3791), .ZN(n3623)
         );
  XNOR2_X1 U4314 ( .A(n3623), .B(n3695), .ZN(n3626) );
  XOR2_X1 U4315 ( .A(n3625), .B(n3626), .Z(n3788) );
  NAND3_X1 U4316 ( .A1(n3884), .A2(n3624), .A3(n3788), .ZN(n3628) );
  OAI22_X1 U4317 ( .A1(n4315), .A2(n3693), .B1(n2043), .B2(n3802), .ZN(n3629)
         );
  XNOR2_X1 U4318 ( .A(n3629), .B(n3695), .ZN(n3798) );
  OAI22_X1 U4319 ( .A1(n4315), .A2(n3694), .B1(n3693), .B2(n3802), .ZN(n3797)
         );
  NAND2_X1 U4320 ( .A1(n3798), .A2(n3797), .ZN(n3630) );
  NAND2_X1 U4321 ( .A1(n4299), .A2(n3273), .ZN(n3632) );
  NAND2_X1 U4322 ( .A1(n2045), .A2(n4199), .ZN(n3631) );
  NAND2_X1 U4323 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  XNOR2_X1 U4324 ( .A(n3633), .B(n2055), .ZN(n3636) );
  NOR2_X1 U4325 ( .A1(n3693), .A2(n4207), .ZN(n3634) );
  AOI21_X1 U4326 ( .B1(n4299), .B2(n2816), .A(n3634), .ZN(n3635) );
  NOR2_X1 U4327 ( .A1(n3636), .A2(n3635), .ZN(n3863) );
  OAI22_X1 U4328 ( .A1(n4202), .A2(n3694), .B1(n3693), .B2(n4185), .ZN(n3638)
         );
  OAI22_X1 U4329 ( .A1(n4202), .A2(n3693), .B1(n2044), .B2(n4185), .ZN(n3637)
         );
  XNOR2_X1 U4330 ( .A(n3637), .B(n3695), .ZN(n3639) );
  XOR2_X1 U4331 ( .A(n3638), .B(n3639), .Z(n3741) );
  INV_X1 U4332 ( .A(n3638), .ZN(n3641) );
  INV_X1 U4333 ( .A(n3639), .ZN(n3640) );
  NAND2_X1 U4334 ( .A1(n3643), .A2(n3642), .ZN(n3819) );
  NAND2_X1 U4335 ( .A1(n4278), .A2(n3273), .ZN(n3645) );
  NAND2_X1 U4336 ( .A1(n2045), .A2(n4153), .ZN(n3644) );
  NAND2_X1 U4337 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  XNOR2_X1 U4338 ( .A(n3646), .B(n3695), .ZN(n3649) );
  NAND2_X1 U4339 ( .A1(n4278), .A2(n2816), .ZN(n3648) );
  NAND2_X1 U4340 ( .A1(n3273), .A2(n4153), .ZN(n3647) );
  NAND2_X1 U4341 ( .A1(n3648), .A2(n3647), .ZN(n3650) );
  NAND2_X1 U4342 ( .A1(n3649), .A2(n3650), .ZN(n3820) );
  NAND2_X1 U4343 ( .A1(n3819), .A2(n3820), .ZN(n3818) );
  INV_X1 U4344 ( .A(n3649), .ZN(n3652) );
  INV_X1 U4345 ( .A(n3650), .ZN(n3651) );
  NAND2_X1 U4346 ( .A1(n3652), .A2(n3651), .ZN(n3822) );
  OAI22_X1 U4347 ( .A1(n4156), .A2(n3693), .B1(n2043), .B2(n4142), .ZN(n3653)
         );
  XNOR2_X1 U4348 ( .A(n3653), .B(n3695), .ZN(n3748) );
  OAI22_X1 U4349 ( .A1(n4156), .A2(n3694), .B1(n3693), .B2(n4142), .ZN(n3654)
         );
  NOR2_X1 U4350 ( .A1(n3748), .A2(n3654), .ZN(n3655) );
  INV_X1 U4351 ( .A(n3654), .ZN(n3747) );
  OAI22_X1 U4352 ( .A1(n4281), .A2(n3693), .B1(n2044), .B2(n4117), .ZN(n3656)
         );
  XNOR2_X1 U4353 ( .A(n3656), .B(n3695), .ZN(n3659) );
  OAI22_X1 U4354 ( .A1(n4281), .A2(n3694), .B1(n3693), .B2(n4117), .ZN(n3658)
         );
  XNOR2_X1 U4355 ( .A(n3659), .B(n3658), .ZN(n3842) );
  OAI22_X1 U4356 ( .A1(n4085), .A2(n3693), .B1(n2043), .B2(n4103), .ZN(n3657)
         );
  XNOR2_X1 U4357 ( .A(n3657), .B(n3695), .ZN(n3662) );
  OAI22_X1 U4358 ( .A1(n4085), .A2(n3694), .B1(n3693), .B2(n4103), .ZN(n3661)
         );
  XNOR2_X1 U4359 ( .A(n3662), .B(n3661), .ZN(n3732) );
  NOR2_X1 U4360 ( .A1(n3659), .A2(n3658), .ZN(n3733) );
  NOR2_X1 U4361 ( .A1(n3732), .A2(n3733), .ZN(n3660) );
  NAND2_X1 U4362 ( .A1(n3662), .A2(n3661), .ZN(n3665) );
  NOR2_X1 U4363 ( .A1(n3693), .A2(n3813), .ZN(n3663) );
  AOI21_X1 U4364 ( .B1(n4249), .B2(n2816), .A(n3663), .ZN(n3666) );
  OAI22_X1 U4365 ( .A1(n3779), .A2(n3693), .B1(n2043), .B2(n3813), .ZN(n3664)
         );
  XNOR2_X1 U4366 ( .A(n3664), .B(n3695), .ZN(n3810) );
  NAND2_X1 U4367 ( .A1(n3808), .A2(n3810), .ZN(n3669) );
  INV_X1 U4368 ( .A(n3666), .ZN(n3667) );
  NAND2_X1 U4369 ( .A1(n3668), .A2(n3667), .ZN(n3807) );
  NAND2_X1 U4370 ( .A1(n3669), .A2(n3807), .ZN(n3774) );
  NAND2_X1 U4371 ( .A1(n4089), .A2(n3273), .ZN(n3671) );
  NAND2_X1 U4372 ( .A1(n2045), .A2(n4248), .ZN(n3670) );
  NAND2_X1 U4373 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  XNOR2_X1 U4374 ( .A(n3672), .B(n2055), .ZN(n3675) );
  NOR2_X1 U4375 ( .A1(n3693), .A2(n4070), .ZN(n3673) );
  AOI21_X1 U4376 ( .B1(n4089), .B2(n2816), .A(n3673), .ZN(n3674) );
  NAND2_X1 U4377 ( .A1(n3675), .A2(n3674), .ZN(n3775) );
  NOR2_X1 U4378 ( .A1(n3675), .A2(n3674), .ZN(n3777) );
  OAI22_X1 U4379 ( .A1(n4252), .A2(n3693), .B1(n2043), .B2(n4053), .ZN(n3676)
         );
  XNOR2_X1 U4380 ( .A(n3676), .B(n3695), .ZN(n3677) );
  OAI22_X1 U4381 ( .A1(n4252), .A2(n3694), .B1(n3693), .B2(n4053), .ZN(n3678)
         );
  NAND2_X1 U4382 ( .A1(n3677), .A2(n3678), .ZN(n3873) );
  NAND2_X1 U4383 ( .A1(n3872), .A2(n3873), .ZN(n3681) );
  INV_X1 U4384 ( .A(n3677), .ZN(n3680) );
  INV_X1 U4385 ( .A(n3678), .ZN(n3679) );
  NAND2_X1 U4386 ( .A1(n3680), .A2(n3679), .ZN(n3874) );
  OAI22_X1 U4387 ( .A1(n4227), .A2(n3693), .B1(n4031), .B2(n2044), .ZN(n3682)
         );
  XNOR2_X1 U4388 ( .A(n3682), .B(n3695), .ZN(n3689) );
  OAI22_X1 U4389 ( .A1(n4227), .A2(n3694), .B1(n4031), .B2(n3693), .ZN(n3688)
         );
  XNOR2_X1 U4390 ( .A(n3691), .B(n3690), .ZN(n3687) );
  NOR2_X1 U4391 ( .A1(n4033), .A2(n3811), .ZN(n3685) );
  AOI22_X1 U4392 ( .A1(n4236), .A2(n3888), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3683) );
  OAI21_X1 U4393 ( .B1(n3868), .B2(n4031), .A(n3683), .ZN(n3684) );
  AOI211_X1 U4394 ( .C1(n3887), .C2(n4036), .A(n3685), .B(n3684), .ZN(n3686)
         );
  OAI21_X1 U4395 ( .B1(n3687), .B2(n3896), .A(n3686), .ZN(U3211) );
  OAI22_X1 U4396 ( .A1(n4238), .A2(n3693), .B1(n2044), .B2(n4225), .ZN(n3698)
         );
  OAI22_X1 U4397 ( .A1(n4238), .A2(n3694), .B1(n3693), .B2(n4225), .ZN(n3696)
         );
  XNOR2_X1 U4398 ( .A(n3696), .B(n3695), .ZN(n3697) );
  XOR2_X1 U4399 ( .A(n3698), .B(n3697), .Z(n3699) );
  INV_X1 U4400 ( .A(n3700), .ZN(n3708) );
  OAI22_X1 U4401 ( .A1(n4227), .A2(n3844), .B1(STATE_REG_SCAN_IN), .B2(n3701), 
        .ZN(n3704) );
  OAI22_X1 U4402 ( .A1(n3702), .A2(n3845), .B1(n3868), .B2(n4225), .ZN(n3703)
         );
  AOI211_X1 U4403 ( .C1(n3708), .C2(n3893), .A(n3704), .B(n3703), .ZN(n3705)
         );
  XNOR2_X1 U4404 ( .A(n3706), .B(n3711), .ZN(n4232) );
  INV_X1 U4405 ( .A(n4029), .ZN(n3707) );
  OAI21_X1 U4406 ( .B1(n3707), .B2(n4225), .A(n2056), .ZN(n4333) );
  INV_X1 U4407 ( .A(n4333), .ZN(n3717) );
  AOI22_X1 U4408 ( .A1(n4136), .A2(n4229), .B1(n3899), .B2(n4135), .ZN(n3710)
         );
  AOI22_X1 U4409 ( .A1(n3708), .A2(n4209), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4391), .ZN(n3709) );
  OAI211_X1 U4410 ( .C1(n4225), .C2(n4141), .A(n3710), .B(n3709), .ZN(n3716)
         );
  INV_X1 U4411 ( .A(n3711), .ZN(n3712) );
  XNOR2_X1 U4412 ( .A(n3713), .B(n3712), .ZN(n3714) );
  NAND2_X1 U4413 ( .A1(n3714), .A2(n4204), .ZN(n4230) );
  NOR2_X1 U4414 ( .A1(n4230), .A2(n4391), .ZN(n3715) );
  AOI211_X1 U4415 ( .C1(n4501), .C2(n3717), .A(n3716), .B(n3715), .ZN(n3718)
         );
  OAI21_X1 U4416 ( .B1(n4232), .B2(n4216), .A(n3718), .ZN(U3262) );
  INV_X1 U4417 ( .A(n3719), .ZN(n3721) );
  NAND2_X1 U4418 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  XNOR2_X1 U4419 ( .A(n3617), .B(n3722), .ZN(n3723) );
  NAND2_X1 U4420 ( .A1(n3723), .A2(n3764), .ZN(n3729) );
  OAI22_X1 U4421 ( .A1(n3868), .A2(n3724), .B1(n3768), .B2(n3844), .ZN(n3727)
         );
  NOR2_X1 U4422 ( .A1(n4692), .A2(STATE_REG_SCAN_IN), .ZN(n4452) );
  INV_X1 U4423 ( .A(n4452), .ZN(n3725) );
  OAI21_X1 U4424 ( .B1(n3845), .B2(n4309), .A(n3725), .ZN(n3726) );
  NOR2_X1 U4425 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  OAI211_X1 U4426 ( .C1(n3811), .C2(n3730), .A(n3729), .B(n3728), .ZN(U3212)
         );
  INV_X1 U4427 ( .A(n3731), .ZN(n3840) );
  OAI21_X1 U4428 ( .B1(n3840), .B2(n3733), .A(n3732), .ZN(n3735) );
  NAND3_X1 U4429 ( .A1(n3735), .A2(n3764), .A3(n3734), .ZN(n3739) );
  OAI22_X1 U4430 ( .A1(n3779), .A2(n3845), .B1(n3868), .B2(n4103), .ZN(n3737)
         );
  OAI22_X1 U4431 ( .A1(n4281), .A2(n3844), .B1(STATE_REG_SCAN_IN), .B2(n4581), 
        .ZN(n3736) );
  NOR2_X1 U4432 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  OAI211_X1 U4433 ( .C1(n3811), .C2(n4105), .A(n3739), .B(n3738), .ZN(U3213)
         );
  XNOR2_X1 U4434 ( .A(n3740), .B(n3741), .ZN(n3742) );
  NAND2_X1 U4435 ( .A1(n3742), .A2(n3764), .ZN(n3746) );
  INV_X1 U4436 ( .A(n4299), .ZN(n4179) );
  OAI22_X1 U4437 ( .A1(n3868), .A2(n4185), .B1(n4179), .B2(n3844), .ZN(n3744)
         );
  INV_X1 U4438 ( .A(n4278), .ZN(n3752) );
  NAND2_X1 U4439 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4001) );
  OAI21_X1 U4440 ( .B1(n3845), .B2(n3752), .A(n4001), .ZN(n3743) );
  NOR2_X1 U4441 ( .A1(n3744), .A2(n3743), .ZN(n3745) );
  OAI211_X1 U4442 ( .C1(n3811), .C2(n4188), .A(n3746), .B(n3745), .ZN(U3216)
         );
  XNOR2_X1 U4443 ( .A(n3748), .B(n3747), .ZN(n3749) );
  XNOR2_X1 U4444 ( .A(n3750), .B(n3749), .ZN(n3751) );
  NAND2_X1 U4445 ( .A1(n3751), .A2(n3764), .ZN(n3758) );
  AOI22_X1 U4446 ( .A1(n4137), .A2(n3887), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3757) );
  OAI22_X1 U4447 ( .A1(n3868), .A2(n4142), .B1(n3752), .B2(n3844), .ZN(n3753)
         );
  INV_X1 U4448 ( .A(n3753), .ZN(n3756) );
  INV_X1 U4449 ( .A(n3754), .ZN(n4138) );
  NAND2_X1 U4450 ( .A1(n3893), .A2(n4138), .ZN(n3755) );
  NAND4_X1 U4451 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(U3220)
         );
  INV_X1 U4452 ( .A(n3759), .ZN(n3761) );
  NOR2_X1 U4453 ( .A1(n3761), .A2(n3760), .ZN(n3762) );
  XNOR2_X1 U4454 ( .A(n3763), .B(n3762), .ZN(n3765) );
  NAND2_X1 U4455 ( .A1(n3765), .A2(n3764), .ZN(n3772) );
  OAI22_X1 U4456 ( .A1(n3868), .A2(n3767), .B1(n3766), .B2(n3844), .ZN(n3770)
         );
  NAND2_X1 U4457 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4428) );
  OAI21_X1 U4458 ( .B1(n3845), .B2(n3768), .A(n4428), .ZN(n3769) );
  NOR2_X1 U4459 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  OAI211_X1 U4460 ( .C1(n3811), .C2(n3773), .A(n3772), .B(n3771), .ZN(U3221)
         );
  INV_X1 U4461 ( .A(n3775), .ZN(n3776) );
  NOR2_X1 U4462 ( .A1(n3777), .A2(n3776), .ZN(n3778) );
  XNOR2_X1 U4463 ( .A(n3774), .B(n3778), .ZN(n3783) );
  OAI22_X1 U4464 ( .A1(n3779), .A2(n3844), .B1(STATE_REG_SCAN_IN), .B2(n4681), 
        .ZN(n3781) );
  OAI22_X1 U4465 ( .A1(n4252), .A2(n3845), .B1(n3868), .B2(n4070), .ZN(n3780)
         );
  AOI211_X1 U4466 ( .C1(n4067), .C2(n3893), .A(n3781), .B(n3780), .ZN(n3782)
         );
  OAI21_X1 U4467 ( .B1(n3783), .B2(n3896), .A(n3782), .ZN(U3222) );
  INV_X1 U4468 ( .A(n3884), .ZN(n3786) );
  OAI21_X1 U4469 ( .B1(n3786), .B2(n3886), .A(n2274), .ZN(n3787) );
  XOR2_X1 U4470 ( .A(n3788), .B(n3787), .Z(n3795) );
  AND2_X1 U4471 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4470) );
  AOI21_X1 U4472 ( .B1(n3887), .B2(n4200), .A(n4470), .ZN(n3790) );
  NAND2_X1 U4473 ( .A1(n3888), .A2(n3901), .ZN(n3789) );
  OAI211_X1 U4474 ( .C1(n3868), .C2(n3791), .A(n3790), .B(n3789), .ZN(n3792)
         );
  AOI21_X1 U4475 ( .B1(n3793), .B2(n3893), .A(n3792), .ZN(n3794) );
  OAI21_X1 U4476 ( .B1(n3795), .B2(n3896), .A(n3794), .ZN(U3223) );
  XNOR2_X1 U4477 ( .A(n3798), .B(n3797), .ZN(n3799) );
  XNOR2_X1 U4478 ( .A(n3796), .B(n3799), .ZN(n3806) );
  NOR2_X1 U4479 ( .A1(STATE_REG_SCAN_IN), .A2(n2523), .ZN(n4479) );
  AOI21_X1 U4480 ( .B1(n3887), .B2(n4299), .A(n4479), .ZN(n3801) );
  NAND2_X1 U4481 ( .A1(n3888), .A2(n3900), .ZN(n3800) );
  OAI211_X1 U4482 ( .C1(n3868), .C2(n3802), .A(n3801), .B(n3800), .ZN(n3803)
         );
  AOI21_X1 U4483 ( .B1(n3804), .B2(n3893), .A(n3803), .ZN(n3805) );
  OAI21_X1 U4484 ( .B1(n3806), .B2(n3896), .A(n3805), .ZN(U3225) );
  NAND2_X1 U4485 ( .A1(n3807), .A2(n3808), .ZN(n3809) );
  XOR2_X1 U4486 ( .A(n3810), .B(n3809), .Z(n3817) );
  NOR2_X1 U4487 ( .A1(n3811), .A2(n4080), .ZN(n3815) );
  AOI22_X1 U4488 ( .A1(n4258), .A2(n3888), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3812) );
  OAI21_X1 U4489 ( .B1(n3868), .B2(n3813), .A(n3812), .ZN(n3814) );
  AOI211_X1 U4490 ( .C1(n3887), .C2(n4089), .A(n3815), .B(n3814), .ZN(n3816)
         );
  OAI21_X1 U4491 ( .B1(n3817), .B2(n3896), .A(n3816), .ZN(U3226) );
  INV_X1 U4492 ( .A(n3818), .ZN(n3823) );
  AOI21_X1 U4493 ( .B1(n3822), .B2(n3820), .A(n3819), .ZN(n3821) );
  AOI21_X1 U4494 ( .B1(n3823), .B2(n3822), .A(n3821), .ZN(n3828) );
  OAI22_X1 U4495 ( .A1(n3868), .A2(n4164), .B1(n4202), .B2(n3844), .ZN(n3825)
         );
  OAI22_X1 U4496 ( .A1(n4156), .A2(n3845), .B1(STATE_REG_SCAN_IN), .B2(n4669), 
        .ZN(n3824) );
  NOR2_X1 U4497 ( .A1(n3825), .A2(n3824), .ZN(n3827) );
  NAND2_X1 U4498 ( .A1(n3893), .A2(n4166), .ZN(n3826) );
  OAI211_X1 U4499 ( .C1(n3828), .C2(n3896), .A(n3827), .B(n3826), .ZN(U3230)
         );
  XNOR2_X1 U4500 ( .A(n3831), .B(n3830), .ZN(n3832) );
  XNOR2_X1 U4501 ( .A(n3829), .B(n3832), .ZN(n3839) );
  NOR2_X1 U4502 ( .A1(STATE_REG_SCAN_IN), .A2(n2330), .ZN(n4442) );
  AOI21_X1 U4503 ( .B1(n3887), .B2(n3902), .A(n4442), .ZN(n3834) );
  NAND2_X1 U4504 ( .A1(n3888), .A2(n3904), .ZN(n3833) );
  OAI211_X1 U4505 ( .C1(n3868), .C2(n3835), .A(n3834), .B(n3833), .ZN(n3836)
         );
  AOI21_X1 U4506 ( .B1(n3837), .B2(n3893), .A(n3836), .ZN(n3838) );
  OAI21_X1 U4507 ( .B1(n3839), .B2(n3896), .A(n3838), .ZN(U3231) );
  AOI21_X1 U4508 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3849) );
  OAI22_X1 U4509 ( .A1(n4156), .A2(n3844), .B1(STATE_REG_SCAN_IN), .B2(n3843), 
        .ZN(n3847) );
  OAI22_X1 U4510 ( .A1(n4085), .A2(n3845), .B1(n3868), .B2(n4117), .ZN(n3846)
         );
  AOI211_X1 U4511 ( .C1(n4118), .C2(n3893), .A(n3847), .B(n3846), .ZN(n3848)
         );
  OAI21_X1 U4512 ( .B1(n3849), .B2(n3896), .A(n3848), .ZN(U3232) );
  XOR2_X1 U4513 ( .A(n3852), .B(n3851), .Z(n3853) );
  XNOR2_X1 U4514 ( .A(n3850), .B(n3853), .ZN(n3861) );
  INV_X1 U4515 ( .A(n3854), .ZN(n3859) );
  AND2_X1 U4516 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4424) );
  AOI21_X1 U4517 ( .B1(n3887), .B2(n3904), .A(n4424), .ZN(n3856) );
  NAND2_X1 U4518 ( .A1(n3888), .A2(n3906), .ZN(n3855) );
  OAI211_X1 U4519 ( .C1(n3868), .C2(n3857), .A(n3856), .B(n3855), .ZN(n3858)
         );
  AOI21_X1 U4520 ( .B1(n3859), .B2(n3893), .A(n3858), .ZN(n3860) );
  OAI21_X1 U4521 ( .B1(n3861), .B2(n3896), .A(n3860), .ZN(U3233) );
  NOR2_X1 U4522 ( .A1(n3863), .A2(n2079), .ZN(n3864) );
  XNOR2_X1 U4523 ( .A(n3862), .B(n3864), .ZN(n3871) );
  INV_X1 U4524 ( .A(n3865), .ZN(n4210) );
  AND2_X1 U4525 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4488) );
  AOI21_X1 U4526 ( .B1(n3887), .B2(n4154), .A(n4488), .ZN(n3867) );
  NAND2_X1 U4527 ( .A1(n3888), .A2(n4200), .ZN(n3866) );
  OAI211_X1 U4528 ( .C1(n3868), .C2(n4207), .A(n3867), .B(n3866), .ZN(n3869)
         );
  AOI21_X1 U4529 ( .B1(n4210), .B2(n3893), .A(n3869), .ZN(n3870) );
  OAI21_X1 U4530 ( .B1(n3871), .B2(n3896), .A(n3870), .ZN(U3235) );
  NAND2_X1 U4531 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  XNOR2_X1 U4532 ( .A(n3872), .B(n3875), .ZN(n3883) );
  AOI22_X1 U4533 ( .A1(n3899), .A2(n3887), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3881) );
  NAND2_X1 U4534 ( .A1(n4054), .A2(n3893), .ZN(n3880) );
  NAND2_X1 U4535 ( .A1(n4089), .A2(n3888), .ZN(n3879) );
  NAND2_X1 U4536 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  AND4_X1 U4537 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3882)
         );
  OAI21_X1 U4538 ( .B1(n3883), .B2(n3896), .A(n3882), .ZN(U3237) );
  NAND2_X1 U4539 ( .A1(n3884), .A2(n2274), .ZN(n3885) );
  XOR2_X1 U4540 ( .A(n3886), .B(n3885), .Z(n3897) );
  AND2_X1 U4541 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4461) );
  AOI21_X1 U4542 ( .B1(n3887), .B2(n3900), .A(n4461), .ZN(n3890) );
  NAND2_X1 U4543 ( .A1(n3888), .A2(n3902), .ZN(n3889) );
  OAI211_X1 U4544 ( .C1(n3868), .C2(n3891), .A(n3890), .B(n3889), .ZN(n3892)
         );
  AOI21_X1 U4545 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3895) );
  OAI21_X1 U4546 ( .B1(n3897), .B2(n3896), .A(n3895), .ZN(U3238) );
  MUX2_X1 U4547 ( .A(DATAO_REG_31__SCAN_IN), .B(n4008), .S(n3915), .Z(U3581)
         );
  MUX2_X1 U4548 ( .A(DATAO_REG_30__SCAN_IN), .B(n3898), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4549 ( .A(DATAO_REG_29__SCAN_IN), .B(n4229), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4550 ( .A(DATAO_REG_28__SCAN_IN), .B(n4036), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4551 ( .A(DATAO_REG_27__SCAN_IN), .B(n3899), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4552 ( .A(DATAO_REG_26__SCAN_IN), .B(n4236), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4553 ( .A(DATAO_REG_25__SCAN_IN), .B(n4089), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4554 ( .A(DATAO_REG_24__SCAN_IN), .B(n4249), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4555 ( .A(DATAO_REG_23__SCAN_IN), .B(n4258), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4556 ( .A(DATAO_REG_22__SCAN_IN), .B(n4137), .S(n3915), .Z(U3572)
         );
  MUX2_X1 U4557 ( .A(DATAO_REG_21__SCAN_IN), .B(n2562), .S(n3915), .Z(U3571)
         );
  MUX2_X1 U4558 ( .A(DATAO_REG_20__SCAN_IN), .B(n4278), .S(n3915), .Z(U3570)
         );
  MUX2_X1 U4559 ( .A(DATAO_REG_19__SCAN_IN), .B(n4154), .S(n3915), .Z(U3569)
         );
  MUX2_X1 U4560 ( .A(DATAO_REG_18__SCAN_IN), .B(n4299), .S(n3915), .Z(U3568)
         );
  MUX2_X1 U4561 ( .A(DATAO_REG_17__SCAN_IN), .B(n4200), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4562 ( .A(DATAO_REG_16__SCAN_IN), .B(n3900), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4563 ( .A(DATAO_REG_15__SCAN_IN), .B(n3901), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4564 ( .A(DATAO_REG_14__SCAN_IN), .B(n3902), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4565 ( .A(DATAO_REG_13__SCAN_IN), .B(n3903), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4566 ( .A(DATAO_REG_12__SCAN_IN), .B(n3904), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4567 ( .A(DATAO_REG_11__SCAN_IN), .B(n3905), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4568 ( .A(DATAO_REG_10__SCAN_IN), .B(n3906), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4569 ( .A(DATAO_REG_9__SCAN_IN), .B(n3907), .S(n3915), .Z(U3559) );
  MUX2_X1 U4570 ( .A(DATAO_REG_8__SCAN_IN), .B(n3908), .S(n3915), .Z(U3558) );
  MUX2_X1 U4571 ( .A(DATAO_REG_7__SCAN_IN), .B(n3909), .S(n3915), .Z(U3557) );
  MUX2_X1 U4572 ( .A(DATAO_REG_6__SCAN_IN), .B(n3910), .S(U4043), .Z(U3556) );
  MUX2_X1 U4573 ( .A(DATAO_REG_5__SCAN_IN), .B(n3911), .S(n3915), .Z(U3555) );
  MUX2_X1 U4574 ( .A(DATAO_REG_4__SCAN_IN), .B(n3912), .S(n3915), .Z(U3554) );
  MUX2_X1 U4575 ( .A(DATAO_REG_3__SCAN_IN), .B(n3913), .S(n3915), .Z(U3553) );
  MUX2_X1 U4576 ( .A(DATAO_REG_2__SCAN_IN), .B(n2087), .S(n3915), .Z(U3552) );
  MUX2_X1 U4577 ( .A(DATAO_REG_1__SCAN_IN), .B(n3914), .S(n3915), .Z(U3551) );
  MUX2_X1 U4578 ( .A(DATAO_REG_0__SCAN_IN), .B(n2815), .S(n3915), .Z(U3550) );
  NAND2_X1 U4579 ( .A1(n3942), .A2(n4390), .ZN(n3924) );
  OAI211_X1 U4580 ( .C1(n3918), .C2(n3917), .A(n4491), .B(n3916), .ZN(n3923)
         );
  OAI211_X1 U4581 ( .C1(n2752), .C2(n3920), .A(n4438), .B(n3931), .ZN(n3922)
         );
  AOI22_X1 U4582 ( .A1(n4489), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3921) );
  NAND4_X1 U4583 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(U3241)
         );
  NOR2_X1 U4584 ( .A1(n3925), .A2(STATE_REG_SCAN_IN), .ZN(n3926) );
  AOI21_X1 U4585 ( .B1(n4489), .B2(ADDR_REG_2__SCAN_IN), .A(n3926), .ZN(n3927)
         );
  OAI21_X1 U4586 ( .B1(n4495), .B2(n3928), .A(n3927), .ZN(n3929) );
  INV_X1 U4587 ( .A(n3929), .ZN(n3940) );
  MUX2_X1 U4588 ( .A(n2750), .B(REG2_REG_2__SCAN_IN), .S(n4389), .Z(n3932) );
  NAND3_X1 U4589 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3933) );
  NAND3_X1 U4590 ( .A1(n4438), .A2(n3934), .A3(n3933), .ZN(n3939) );
  OAI211_X1 U4591 ( .C1(n3937), .C2(n3936), .A(n4491), .B(n3935), .ZN(n3938)
         );
  NAND4_X1 U4592 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(U3242)
         );
  NAND2_X1 U4593 ( .A1(n3942), .A2(n4388), .ZN(n3951) );
  OAI211_X1 U4594 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3944), .A(n4491), .B(n3943), 
        .ZN(n3950) );
  AOI22_X1 U4595 ( .A1(n4489), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3949) );
  XNOR2_X1 U4596 ( .A(n3946), .B(n3945), .ZN(n3947) );
  NAND2_X1 U4597 ( .A1(n4438), .A2(n3947), .ZN(n3948) );
  NAND4_X1 U4598 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(U3243)
         );
  INV_X1 U4599 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3952) );
  MUX2_X1 U4600 ( .A(REG2_REG_19__SCAN_IN), .B(n3952), .S(n4381), .Z(n3969) );
  INV_X1 U4601 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4602 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4510), .B1(n3970), .B2(
        n3953), .ZN(n4487) );
  NOR2_X1 U4603 ( .A1(n3995), .A2(REG2_REG_17__SCAN_IN), .ZN(n3954) );
  AOI21_X1 U4604 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3995), .A(n3954), .ZN(n4477) );
  NOR2_X1 U4605 ( .A1(n4437), .A2(n4514), .ZN(n4436) );
  NAND2_X1 U4606 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3973), .ZN(n3960) );
  INV_X1 U4607 ( .A(n3973), .ZN(n4517) );
  AOI22_X1 U4608 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3973), .B1(n4517), .B2(
        n3259), .ZN(n4420) );
  NAND2_X1 U4609 ( .A1(n3974), .A2(REG2_REG_9__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4610 ( .A1(n3974), .A2(REG2_REG_9__SCAN_IN), .B1(n2445), .B2(n4520), .ZN(n4400) );
  OAI22_X1 U4611 ( .A1(n3956), .A2(n4498), .B1(n3955), .B2(n4382), .ZN(n4399)
         );
  NAND2_X1 U4612 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U4613 ( .A1(n3957), .A2(n4398), .ZN(n3958) );
  NAND2_X1 U4614 ( .A1(n3981), .A2(n3958), .ZN(n3959) );
  INV_X1 U4615 ( .A(n3981), .ZN(n4518) );
  XNOR2_X1 U4616 ( .A(n3958), .B(n4518), .ZN(n4407) );
  NAND2_X1 U4617 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4407), .ZN(n4406) );
  NAND2_X1 U4618 ( .A1(n3959), .A2(n4406), .ZN(n4419) );
  NAND2_X1 U4619 ( .A1(n4420), .A2(n4419), .ZN(n4418) );
  NAND2_X1 U4620 ( .A1(n4515), .A2(n3961), .ZN(n3962) );
  XNOR2_X1 U4621 ( .A(n3961), .B(n4435), .ZN(n4427) );
  NAND2_X1 U4622 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4427), .ZN(n4426) );
  NOR2_X1 U4623 ( .A1(n2131), .A2(n3963), .ZN(n3964) );
  NAND2_X1 U4624 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3971), .ZN(n3965) );
  OAI21_X1 U4625 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3971), .A(n3965), .ZN(n4458) );
  INV_X1 U4626 ( .A(n3992), .ZN(n4512) );
  NAND2_X1 U4627 ( .A1(n3966), .A2(n4512), .ZN(n3967) );
  AOI21_X1 U4628 ( .B1(n3970), .B2(REG2_REG_18__SCAN_IN), .A(n4486), .ZN(n3968) );
  XOR2_X1 U4629 ( .A(n3969), .B(n3968), .Z(n4006) );
  INV_X1 U4630 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4631 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3970), .B1(n4510), .B2(
        n3997), .ZN(n4492) );
  NOR2_X1 U4632 ( .A1(n3995), .A2(REG1_REG_17__SCAN_IN), .ZN(n3996) );
  NAND2_X1 U4633 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3971), .ZN(n3991) );
  INV_X1 U4634 ( .A(n3971), .ZN(n4513) );
  AOI22_X1 U4635 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3971), .B1(n4513), .B2(
        n3382), .ZN(n4464) );
  NAND2_X1 U4636 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3972), .ZN(n3987) );
  AOI22_X1 U4637 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3972), .B1(n4514), .B2(
        n3372), .ZN(n4446) );
  NAND2_X1 U4638 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3973), .ZN(n3984) );
  AOI22_X1 U4639 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3973), .B1(n4517), .B2(
        n3327), .ZN(n4417) );
  NAND2_X1 U4640 ( .A1(n3974), .A2(REG1_REG_9__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4641 ( .A1(n3974), .A2(REG1_REG_9__SCAN_IN), .B1(n2444), .B2(n4520), .ZN(n4397) );
  INV_X1 U4642 ( .A(n3975), .ZN(n3979) );
  INV_X1 U4643 ( .A(n3976), .ZN(n3977) );
  NAND2_X1 U4644 ( .A1(n4397), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U4645 ( .A1(n3980), .A2(n4395), .ZN(n3982) );
  NAND2_X1 U4646 ( .A1(n3981), .A2(n3982), .ZN(n3983) );
  XNOR2_X1 U4647 ( .A(n3982), .B(n4518), .ZN(n4412) );
  NAND2_X1 U4648 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U4649 ( .A1(n3983), .A2(n4411), .ZN(n4416) );
  NAND2_X1 U4650 ( .A1(n4417), .A2(n4416), .ZN(n4415) );
  NAND2_X1 U4651 ( .A1(n3984), .A2(n4415), .ZN(n3985) );
  NAND2_X1 U4652 ( .A1(n4515), .A2(n3985), .ZN(n3986) );
  XNOR2_X1 U4653 ( .A(n3985), .B(n4435), .ZN(n4432) );
  NAND2_X1 U4654 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U4655 ( .A1(n3986), .A2(n4431), .ZN(n4445) );
  NAND2_X1 U4656 ( .A1(n4446), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U4657 ( .A1(n3987), .A2(n4444), .ZN(n3989) );
  NAND2_X1 U4658 ( .A1(n3988), .A2(n3989), .ZN(n3990) );
  XNOR2_X1 U4659 ( .A(n3989), .B(n2131), .ZN(n4454) );
  NAND2_X1 U4660 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4454), .ZN(n4453) );
  NOR2_X1 U4661 ( .A1(n3992), .A2(n3993), .ZN(n3994) );
  AOI22_X1 U4662 ( .A1(n3995), .A2(n4305), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4511), .ZN(n4480) );
  OAI21_X1 U4663 ( .B1(n3997), .B2(n4510), .A(n4490), .ZN(n3999) );
  MUX2_X1 U4664 ( .A(n4292), .B(REG1_REG_19__SCAN_IN), .S(n4381), .Z(n3998) );
  XNOR2_X1 U4665 ( .A(n3999), .B(n3998), .ZN(n4004) );
  NAND2_X1 U4666 ( .A1(n4489), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4000) );
  OAI211_X1 U4667 ( .C1(n4495), .C2(n4002), .A(n4001), .B(n4000), .ZN(n4003)
         );
  AOI21_X1 U4668 ( .B1(n4004), .B2(n4491), .A(n4003), .ZN(n4005) );
  OAI21_X1 U4669 ( .B1(n4006), .B2(n4485), .A(n4005), .ZN(U3259) );
  XNOR2_X1 U4670 ( .A(n4220), .B(n4009), .ZN(n4326) );
  NAND2_X1 U4671 ( .A1(n4008), .A2(n4007), .ZN(n4221) );
  OAI21_X1 U4672 ( .B1(n4009), .B2(n4226), .A(n4221), .ZN(n4323) );
  NAND2_X1 U4673 ( .A1(n4191), .A2(n4323), .ZN(n4011) );
  NAND2_X1 U4674 ( .A1(n4119), .A2(REG2_REG_31__SCAN_IN), .ZN(n4010) );
  OAI211_X1 U4675 ( .C1(n4326), .C2(n4187), .A(n4011), .B(n4010), .ZN(U3260)
         );
  INV_X1 U4676 ( .A(n4012), .ZN(n4023) );
  INV_X1 U4677 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4013) );
  OAI22_X1 U4678 ( .A1(n4141), .A2(n4014), .B1(n4013), .B2(n4191), .ZN(n4015)
         );
  AOI21_X1 U4679 ( .B1(n4036), .B2(n4135), .A(n4015), .ZN(n4022) );
  INV_X1 U4680 ( .A(n4016), .ZN(n4020) );
  OAI22_X1 U4681 ( .A1(n4018), .A2(n4187), .B1(n4017), .B2(n4496), .ZN(n4019)
         );
  OAI21_X1 U4682 ( .B1(n4020), .B2(n4019), .A(n4191), .ZN(n4021) );
  OAI211_X1 U4683 ( .C1(n4023), .C2(n4216), .A(n4022), .B(n4021), .ZN(U3354)
         );
  XNOR2_X1 U4684 ( .A(n4024), .B(n4025), .ZN(n4241) );
  INV_X1 U4685 ( .A(n4241), .ZN(n4041) );
  NAND2_X1 U4686 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  AOI21_X1 U4687 ( .B1(n4028), .B2(n4027), .A(n4182), .ZN(n4240) );
  INV_X1 U4688 ( .A(n4052), .ZN(n4030) );
  OAI21_X1 U4689 ( .B1(n4030), .B2(n4031), .A(n4029), .ZN(n4337) );
  NOR2_X1 U4690 ( .A1(n4141), .A2(n4031), .ZN(n4035) );
  INV_X1 U4691 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4032) );
  OAI22_X1 U4692 ( .A1(n4033), .A2(n4496), .B1(n4032), .B2(n4191), .ZN(n4034)
         );
  AOI211_X1 U4693 ( .C1(n4135), .C2(n4236), .A(n4035), .B(n4034), .ZN(n4038)
         );
  NAND2_X1 U4694 ( .A1(n4036), .A2(n4136), .ZN(n4037) );
  OAI211_X1 U4695 ( .C1(n4337), .C2(n4187), .A(n4038), .B(n4037), .ZN(n4039)
         );
  AOI21_X1 U4696 ( .B1(n4240), .B2(n4191), .A(n4039), .ZN(n4040) );
  OAI21_X1 U4697 ( .B1(n4041), .B2(n4216), .A(n4040), .ZN(U3263) );
  XNOR2_X1 U4698 ( .A(n4043), .B(n4042), .ZN(n4245) );
  INV_X1 U4699 ( .A(n4245), .ZN(n4058) );
  INV_X1 U4700 ( .A(n4060), .ZN(n4046) );
  OAI21_X1 U4701 ( .B1(n4046), .B2(n4045), .A(n4044), .ZN(n4048) );
  XNOR2_X1 U4702 ( .A(n4048), .B(n4047), .ZN(n4051) );
  OAI22_X1 U4703 ( .A1(n4227), .A2(n4314), .B1(n4226), .B2(n4053), .ZN(n4049)
         );
  AOI21_X1 U4704 ( .B1(n4277), .B2(n4089), .A(n4049), .ZN(n4050) );
  OAI21_X1 U4705 ( .B1(n4051), .B2(n4182), .A(n4050), .ZN(n4244) );
  OAI21_X1 U4706 ( .B1(n4066), .B2(n4053), .A(n4052), .ZN(n4341) );
  AOI22_X1 U4707 ( .A1(n4054), .A2(n4209), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4391), .ZN(n4055) );
  OAI21_X1 U4708 ( .B1(n4341), .B2(n4187), .A(n4055), .ZN(n4056) );
  AOI21_X1 U4709 ( .B1(n4244), .B2(n4191), .A(n4056), .ZN(n4057) );
  OAI21_X1 U4710 ( .B1(n4058), .B2(n4216), .A(n4057), .ZN(U3264) );
  NAND2_X1 U4711 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  XNOR2_X1 U4712 ( .A(n4061), .B(n4064), .ZN(n4062) );
  NAND2_X1 U4713 ( .A1(n4062), .A2(n4204), .ZN(n4251) );
  XOR2_X1 U4714 ( .A(n4064), .B(n4063), .Z(n4254) );
  NAND2_X1 U4715 ( .A1(n4254), .A2(n4132), .ZN(n4074) );
  NOR2_X1 U4716 ( .A1(n2070), .A2(n4070), .ZN(n4065) );
  OR2_X1 U4717 ( .A1(n4066), .A2(n4065), .ZN(n4345) );
  INV_X1 U4718 ( .A(n4345), .ZN(n4072) );
  AOI22_X1 U4719 ( .A1(n4236), .A2(n4136), .B1(n4135), .B2(n4249), .ZN(n4069)
         );
  AOI22_X1 U4720 ( .A1(n4067), .A2(n4209), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4391), .ZN(n4068) );
  OAI211_X1 U4721 ( .C1(n4070), .C2(n4141), .A(n4069), .B(n4068), .ZN(n4071)
         );
  AOI21_X1 U4722 ( .B1(n4072), .B2(n4501), .A(n4071), .ZN(n4073) );
  OAI211_X1 U4723 ( .C1(n4119), .C2(n4251), .A(n4074), .B(n4073), .ZN(U3265)
         );
  XOR2_X1 U4724 ( .A(n4077), .B(n4075), .Z(n4076) );
  NAND2_X1 U4725 ( .A1(n4076), .A2(n4204), .ZN(n4260) );
  XNOR2_X1 U4726 ( .A(n4078), .B(n4077), .ZN(n4263) );
  NAND2_X1 U4727 ( .A1(n4263), .A2(n4132), .ZN(n4091) );
  INV_X1 U4728 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4079) );
  OAI22_X1 U4729 ( .A1(n4080), .A2(n4496), .B1(n4079), .B2(n4191), .ZN(n4081)
         );
  AOI21_X1 U4730 ( .B1(n4257), .B2(n4082), .A(n4081), .ZN(n4083) );
  OAI21_X1 U4731 ( .B1(n4085), .B2(n4084), .A(n4083), .ZN(n4088) );
  AND2_X1 U4732 ( .A1(n4102), .A2(n4257), .ZN(n4086) );
  OR2_X1 U4733 ( .A1(n4086), .A2(n2070), .ZN(n4349) );
  NOR2_X1 U4734 ( .A1(n4349), .A2(n4187), .ZN(n4087) );
  AOI211_X1 U4735 ( .C1(n4136), .C2(n4089), .A(n4088), .B(n4087), .ZN(n4090)
         );
  OAI211_X1 U4736 ( .C1(n4391), .C2(n4260), .A(n4091), .B(n4090), .ZN(U3266)
         );
  XOR2_X1 U4737 ( .A(n4097), .B(n4092), .Z(n4267) );
  INV_X1 U4738 ( .A(n4267), .ZN(n4110) );
  INV_X1 U4739 ( .A(n4093), .ZN(n4095) );
  AOI21_X1 U4740 ( .B1(n4128), .B2(n4095), .A(n4094), .ZN(n4111) );
  OAI21_X1 U4741 ( .B1(n4111), .B2(n4121), .A(n4096), .ZN(n4098) );
  XNOR2_X1 U4742 ( .A(n4098), .B(n4097), .ZN(n4101) );
  OAI22_X1 U4743 ( .A1(n4281), .A2(n4308), .B1(n4226), .B2(n4103), .ZN(n4099)
         );
  AOI21_X1 U4744 ( .B1(n4298), .B2(n4249), .A(n4099), .ZN(n4100) );
  OAI21_X1 U4745 ( .B1(n4101), .B2(n4182), .A(n4100), .ZN(n4266) );
  INV_X1 U4746 ( .A(n4116), .ZN(n4104) );
  OAI21_X1 U4747 ( .B1(n4104), .B2(n4103), .A(n4102), .ZN(n4353) );
  INV_X1 U4748 ( .A(n4105), .ZN(n4106) );
  AOI22_X1 U4749 ( .A1(n4106), .A2(n4209), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4391), .ZN(n4107) );
  OAI21_X1 U4750 ( .B1(n4353), .B2(n4187), .A(n4107), .ZN(n4108) );
  AOI21_X1 U4751 ( .B1(n4266), .B2(n4191), .A(n4108), .ZN(n4109) );
  OAI21_X1 U4752 ( .B1(n4110), .B2(n4216), .A(n4109), .ZN(U3267) );
  XNOR2_X1 U4753 ( .A(n4111), .B(n4121), .ZN(n4112) );
  NAND2_X1 U4754 ( .A1(n4112), .A2(n4204), .ZN(n4115) );
  OAI22_X1 U4755 ( .A1(n4156), .A2(n4308), .B1(n4117), .B2(n4226), .ZN(n4113)
         );
  AOI21_X1 U4756 ( .B1(n4258), .B2(n4298), .A(n4113), .ZN(n4114) );
  NAND2_X1 U4757 ( .A1(n4115), .A2(n4114), .ZN(n4271) );
  OAI21_X1 U4758 ( .B1(n4133), .B2(n4117), .A(n4116), .ZN(n4357) );
  AOI22_X1 U4759 ( .A1(REG2_REG_22__SCAN_IN), .A2(n4119), .B1(n4118), .B2(
        n4209), .ZN(n4120) );
  OAI21_X1 U4760 ( .B1(n4357), .B2(n4187), .A(n4120), .ZN(n4125) );
  NOR2_X1 U4761 ( .A1(n4122), .A2(n4121), .ZN(n4270) );
  INV_X1 U4762 ( .A(n4272), .ZN(n4123) );
  NOR3_X1 U4763 ( .A1(n4270), .A2(n4123), .A3(n4216), .ZN(n4124) );
  AOI211_X1 U4764 ( .C1(n4191), .C2(n4271), .A(n4125), .B(n4124), .ZN(n4126)
         );
  INV_X1 U4765 ( .A(n4126), .ZN(U3268) );
  INV_X1 U4766 ( .A(n4131), .ZN(n4127) );
  XNOR2_X1 U4767 ( .A(n4128), .B(n4127), .ZN(n4129) );
  NAND2_X1 U4768 ( .A1(n4129), .A2(n4204), .ZN(n4280) );
  XOR2_X1 U4769 ( .A(n4131), .B(n4130), .Z(n4283) );
  NAND2_X1 U4770 ( .A1(n4283), .A2(n4132), .ZN(n4146) );
  INV_X1 U4771 ( .A(n4133), .ZN(n4134) );
  OAI21_X1 U4772 ( .B1(n4162), .B2(n4142), .A(n4134), .ZN(n4361) );
  INV_X1 U4773 ( .A(n4361), .ZN(n4144) );
  AOI22_X1 U4774 ( .A1(n4137), .A2(n4136), .B1(n4135), .B2(n4278), .ZN(n4140)
         );
  AOI22_X1 U4775 ( .A1(n4119), .A2(REG2_REG_21__SCAN_IN), .B1(n4138), .B2(
        n4209), .ZN(n4139) );
  OAI211_X1 U4776 ( .C1(n4142), .C2(n4141), .A(n4140), .B(n4139), .ZN(n4143)
         );
  AOI21_X1 U4777 ( .B1(n4144), .B2(n4501), .A(n4143), .ZN(n4145) );
  OAI211_X1 U4778 ( .C1(n4119), .C2(n4280), .A(n4146), .B(n4145), .ZN(U3269)
         );
  XNOR2_X1 U4779 ( .A(n4147), .B(n4151), .ZN(n4161) );
  INV_X1 U4780 ( .A(n4148), .ZN(n4149) );
  NAND2_X1 U4781 ( .A1(n4150), .A2(n4149), .ZN(n4152) );
  XNOR2_X1 U4782 ( .A(n4152), .B(n4151), .ZN(n4158) );
  AOI22_X1 U4783 ( .A1(n4154), .A2(n4277), .B1(n4153), .B2(n4310), .ZN(n4155)
         );
  OAI21_X1 U4784 ( .B1(n4156), .B2(n4314), .A(n4155), .ZN(n4157) );
  AOI21_X1 U4785 ( .B1(n4158), .B2(n4204), .A(n4157), .ZN(n4159) );
  OAI21_X1 U4786 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4286) );
  INV_X1 U4787 ( .A(n4286), .ZN(n4170) );
  INV_X1 U4788 ( .A(n4161), .ZN(n4287) );
  INV_X1 U4789 ( .A(n4184), .ZN(n4165) );
  INV_X1 U4790 ( .A(n4162), .ZN(n4163) );
  OAI21_X1 U4791 ( .B1(n4165), .B2(n4164), .A(n4163), .ZN(n4365) );
  AOI22_X1 U4792 ( .A1(n4119), .A2(REG2_REG_20__SCAN_IN), .B1(n4166), .B2(
        n4209), .ZN(n4167) );
  OAI21_X1 U4793 ( .B1(n4365), .B2(n4187), .A(n4167), .ZN(n4168) );
  AOI21_X1 U4794 ( .B1(n4287), .B2(n4502), .A(n4168), .ZN(n4169) );
  OAI21_X1 U4795 ( .B1(n4170), .B2(n4391), .A(n4169), .ZN(U3270) );
  XNOR2_X1 U4796 ( .A(n4171), .B(n4178), .ZN(n4291) );
  INV_X1 U4797 ( .A(n4291), .ZN(n4193) );
  NAND2_X1 U4798 ( .A1(n4173), .A2(n4172), .ZN(n4197) );
  INV_X1 U4799 ( .A(n4174), .ZN(n4176) );
  OAI21_X1 U4800 ( .B1(n4197), .B2(n4176), .A(n4175), .ZN(n4177) );
  XOR2_X1 U4801 ( .A(n4178), .B(n4177), .Z(n4183) );
  OAI22_X1 U4802 ( .A1(n4179), .A2(n4308), .B1(n4226), .B2(n4185), .ZN(n4180)
         );
  AOI21_X1 U4803 ( .B1(n4298), .B2(n4278), .A(n4180), .ZN(n4181) );
  OAI21_X1 U4804 ( .B1(n4183), .B2(n4182), .A(n4181), .ZN(n4290) );
  INV_X1 U4805 ( .A(n4206), .ZN(n4186) );
  OAI21_X1 U4806 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4370) );
  NOR2_X1 U4807 ( .A1(n4370), .A2(n4187), .ZN(n4190) );
  OAI22_X1 U4808 ( .A1(n4191), .A2(n3952), .B1(n4188), .B2(n4496), .ZN(n4189)
         );
  AOI211_X1 U4809 ( .C1(n4290), .C2(n4191), .A(n4190), .B(n4189), .ZN(n4192)
         );
  OAI21_X1 U4810 ( .B1(n4193), .B2(n4216), .A(n4192), .ZN(U3271) );
  OAI21_X1 U4811 ( .B1(n4195), .B2(n4198), .A(n4194), .ZN(n4196) );
  INV_X1 U4812 ( .A(n4196), .ZN(n4296) );
  XOR2_X1 U4813 ( .A(n4198), .B(n4197), .Z(n4205) );
  AOI22_X1 U4814 ( .A1(n4200), .A2(n4277), .B1(n4199), .B2(n4310), .ZN(n4201)
         );
  OAI21_X1 U4815 ( .B1(n4202), .B2(n4314), .A(n4201), .ZN(n4203) );
  AOI21_X1 U4816 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n4295) );
  INV_X1 U4817 ( .A(n4295), .ZN(n4214) );
  OAI211_X1 U4818 ( .C1(n4208), .C2(n4207), .A(n4206), .B(n4317), .ZN(n4294)
         );
  AOI22_X1 U4819 ( .A1(n4119), .A2(REG2_REG_18__SCAN_IN), .B1(n4210), .B2(
        n4209), .ZN(n4211) );
  OAI21_X1 U4820 ( .B1(n4294), .B2(n4212), .A(n4211), .ZN(n4213) );
  AOI21_X1 U4821 ( .B1(n4214), .B2(n4191), .A(n4213), .ZN(n4215) );
  OAI21_X1 U4822 ( .B1(n4296), .B2(n4216), .A(n4215), .ZN(U3272) );
  NOR2_X1 U4823 ( .A1(n4545), .A2(n4217), .ZN(n4218) );
  AOI21_X1 U4824 ( .B1(n4545), .B2(n4323), .A(n4218), .ZN(n4219) );
  OAI21_X1 U4825 ( .B1(n4326), .B2(n4307), .A(n4219), .ZN(U3549) );
  AOI21_X1 U4826 ( .B1(n4223), .B2(n2052), .A(n4220), .ZN(n4392) );
  INV_X1 U4827 ( .A(n4392), .ZN(n4329) );
  INV_X1 U4828 ( .A(n4221), .ZN(n4222) );
  AOI21_X1 U4829 ( .B1(n4223), .B2(n4310), .A(n4222), .ZN(n4394) );
  MUX2_X1 U4830 ( .A(n4394), .B(n2673), .S(n4543), .Z(n4224) );
  OAI21_X1 U4831 ( .B1(n4329), .B2(n4307), .A(n4224), .ZN(U3548) );
  OAI22_X1 U4832 ( .A1(n4227), .A2(n4308), .B1(n4226), .B2(n4225), .ZN(n4228)
         );
  AOI21_X1 U4833 ( .B1(n4298), .B2(n4229), .A(n4228), .ZN(n4231) );
  OAI211_X1 U4834 ( .C1(n4232), .C2(n4321), .A(n4231), .B(n4230), .ZN(n4330)
         );
  MUX2_X1 U4835 ( .A(REG1_REG_28__SCAN_IN), .B(n4330), .S(n4545), .Z(n4233) );
  INV_X1 U4836 ( .A(n4233), .ZN(n4234) );
  OAI21_X1 U4837 ( .B1(n4307), .B2(n4333), .A(n4234), .ZN(U3546) );
  AOI22_X1 U4838 ( .A1(n4236), .A2(n4277), .B1(n4235), .B2(n4310), .ZN(n4237)
         );
  OAI21_X1 U4839 ( .B1(n4238), .B2(n4314), .A(n4237), .ZN(n4239) );
  AOI211_X1 U4840 ( .C1(n4241), .C2(n4531), .A(n4240), .B(n4239), .ZN(n4334)
         );
  MUX2_X1 U4841 ( .A(n4242), .B(n4334), .S(n4545), .Z(n4243) );
  OAI21_X1 U4842 ( .B1(n4307), .B2(n4337), .A(n4243), .ZN(U3545) );
  AOI21_X1 U4843 ( .B1(n4245), .B2(n4531), .A(n4244), .ZN(n4338) );
  MUX2_X1 U4844 ( .A(n4246), .B(n4338), .S(n4545), .Z(n4247) );
  OAI21_X1 U4845 ( .B1(n4307), .B2(n4341), .A(n4247), .ZN(U3544) );
  AOI22_X1 U4846 ( .A1(n4249), .A2(n4277), .B1(n4248), .B2(n4310), .ZN(n4250)
         );
  OAI211_X1 U4847 ( .C1(n4252), .C2(n4314), .A(n4251), .B(n4250), .ZN(n4253)
         );
  AOI21_X1 U4848 ( .B1(n4254), .B2(n4531), .A(n4253), .ZN(n4342) );
  MUX2_X1 U4849 ( .A(n4255), .B(n4342), .S(n4545), .Z(n4256) );
  OAI21_X1 U4850 ( .B1(n4307), .B2(n4345), .A(n4256), .ZN(U3543) );
  AOI22_X1 U4851 ( .A1(n4258), .A2(n4277), .B1(n4310), .B2(n4257), .ZN(n4259)
         );
  OAI211_X1 U4852 ( .C1(n4261), .C2(n4314), .A(n4260), .B(n4259), .ZN(n4262)
         );
  AOI21_X1 U4853 ( .B1(n4263), .B2(n4531), .A(n4262), .ZN(n4346) );
  MUX2_X1 U4854 ( .A(n4264), .B(n4346), .S(n4545), .Z(n4265) );
  OAI21_X1 U4855 ( .B1(n4307), .B2(n4349), .A(n4265), .ZN(U3542) );
  AOI21_X1 U4856 ( .B1(n4267), .B2(n4531), .A(n4266), .ZN(n4350) );
  MUX2_X1 U4857 ( .A(n4268), .B(n4350), .S(n4545), .Z(n4269) );
  OAI21_X1 U4858 ( .B1(n4307), .B2(n4353), .A(n4269), .ZN(U3541) );
  NOR2_X1 U4859 ( .A1(n4270), .A2(n4321), .ZN(n4273) );
  AOI21_X1 U4860 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4354) );
  MUX2_X1 U4861 ( .A(n4274), .B(n4354), .S(n4545), .Z(n4275) );
  OAI21_X1 U4862 ( .B1(n4307), .B2(n4357), .A(n4275), .ZN(U3540) );
  AOI22_X1 U4863 ( .A1(n4278), .A2(n4277), .B1(n4276), .B2(n4310), .ZN(n4279)
         );
  OAI211_X1 U4864 ( .C1(n4281), .C2(n4314), .A(n4280), .B(n4279), .ZN(n4282)
         );
  AOI21_X1 U4865 ( .B1(n4283), .B2(n4531), .A(n4282), .ZN(n4358) );
  MUX2_X1 U4866 ( .A(n4284), .B(n4358), .S(n4545), .Z(n4285) );
  OAI21_X1 U4867 ( .B1(n4307), .B2(n4361), .A(n4285), .ZN(U3539) );
  AOI21_X1 U4868 ( .B1(n4529), .B2(n4287), .A(n4286), .ZN(n4362) );
  MUX2_X1 U4869 ( .A(n4288), .B(n4362), .S(n4545), .Z(n4289) );
  OAI21_X1 U4870 ( .B1(n4307), .B2(n4365), .A(n4289), .ZN(U3538) );
  AOI21_X1 U4871 ( .B1(n4291), .B2(n4531), .A(n4290), .ZN(n4366) );
  MUX2_X1 U4872 ( .A(n4292), .B(n4366), .S(n4545), .Z(n4293) );
  OAI21_X1 U4873 ( .B1(n4307), .B2(n4370), .A(n4293), .ZN(U3537) );
  OAI211_X1 U4874 ( .C1(n4296), .C2(n4321), .A(n4295), .B(n4294), .ZN(n4371)
         );
  MUX2_X1 U4875 ( .A(REG1_REG_18__SCAN_IN), .B(n4371), .S(n4545), .Z(U3536) );
  AOI22_X1 U4876 ( .A1(n4299), .A2(n4298), .B1(n4310), .B2(n4297), .ZN(n4300)
         );
  OAI211_X1 U4877 ( .C1(n4302), .C2(n4308), .A(n4301), .B(n4300), .ZN(n4303)
         );
  AOI21_X1 U4878 ( .B1(n4304), .B2(n4531), .A(n4303), .ZN(n4372) );
  MUX2_X1 U4879 ( .A(n4305), .B(n4372), .S(n4545), .Z(n4306) );
  OAI21_X1 U4880 ( .B1(n4307), .B2(n4375), .A(n4306), .ZN(U3535) );
  OR2_X1 U4881 ( .A1(n4309), .A2(n4308), .ZN(n4313) );
  NAND2_X1 U4882 ( .A1(n4311), .A2(n4310), .ZN(n4312) );
  OAI211_X1 U4883 ( .C1(n4315), .C2(n4314), .A(n4313), .B(n4312), .ZN(n4316)
         );
  AOI21_X1 U4884 ( .B1(n4318), .B2(n4317), .A(n4316), .ZN(n4320) );
  OAI211_X1 U4885 ( .C1(n4322), .C2(n4321), .A(n4320), .B(n4319), .ZN(n4376)
         );
  MUX2_X1 U4886 ( .A(REG1_REG_16__SCAN_IN), .B(n4376), .S(n4545), .Z(U3534) );
  NAND2_X1 U4887 ( .A1(n4539), .A2(n4323), .ZN(n4325) );
  NAND2_X1 U4888 ( .A1(n4537), .A2(REG0_REG_31__SCAN_IN), .ZN(n4324) );
  OAI211_X1 U4889 ( .C1(n4326), .C2(n4369), .A(n4325), .B(n4324), .ZN(U3517)
         );
  INV_X1 U4890 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U4891 ( .A(n4394), .B(n4327), .S(n4537), .Z(n4328) );
  OAI21_X1 U4892 ( .B1(n4329), .B2(n4369), .A(n4328), .ZN(U3516) );
  MUX2_X1 U4893 ( .A(REG0_REG_28__SCAN_IN), .B(n4330), .S(n4539), .Z(n4331) );
  INV_X1 U4894 ( .A(n4331), .ZN(n4332) );
  OAI21_X1 U4895 ( .B1(n4333), .B2(n4369), .A(n4332), .ZN(U3514) );
  INV_X1 U4896 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4335) );
  MUX2_X1 U4897 ( .A(n4335), .B(n4334), .S(n4539), .Z(n4336) );
  OAI21_X1 U4898 ( .B1(n4337), .B2(n4369), .A(n4336), .ZN(U3513) );
  INV_X1 U4899 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4339) );
  MUX2_X1 U4900 ( .A(n4339), .B(n4338), .S(n4539), .Z(n4340) );
  OAI21_X1 U4901 ( .B1(n4341), .B2(n4369), .A(n4340), .ZN(U3512) );
  INV_X1 U4902 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4343) );
  MUX2_X1 U4903 ( .A(n4343), .B(n4342), .S(n4539), .Z(n4344) );
  OAI21_X1 U4904 ( .B1(n4345), .B2(n4369), .A(n4344), .ZN(U3511) );
  INV_X1 U4905 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U4906 ( .A(n4347), .B(n4346), .S(n4539), .Z(n4348) );
  OAI21_X1 U4907 ( .B1(n4349), .B2(n4369), .A(n4348), .ZN(U3510) );
  INV_X1 U4908 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U4909 ( .A(n4351), .B(n4350), .S(n4539), .Z(n4352) );
  OAI21_X1 U4910 ( .B1(n4353), .B2(n4369), .A(n4352), .ZN(U3509) );
  INV_X1 U4911 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4355) );
  MUX2_X1 U4912 ( .A(n4355), .B(n4354), .S(n4539), .Z(n4356) );
  OAI21_X1 U4913 ( .B1(n4357), .B2(n4369), .A(n4356), .ZN(U3508) );
  INV_X1 U4914 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U4915 ( .A(n4359), .B(n4358), .S(n4539), .Z(n4360) );
  OAI21_X1 U4916 ( .B1(n4361), .B2(n4369), .A(n4360), .ZN(U3507) );
  INV_X1 U4917 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4918 ( .A(n4363), .B(n4362), .S(n4539), .Z(n4364) );
  OAI21_X1 U4919 ( .B1(n4365), .B2(n4369), .A(n4364), .ZN(U3506) );
  INV_X1 U4920 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4367) );
  MUX2_X1 U4921 ( .A(n4367), .B(n4366), .S(n4539), .Z(n4368) );
  OAI21_X1 U4922 ( .B1(n4370), .B2(n4369), .A(n4368), .ZN(U3505) );
  MUX2_X1 U4923 ( .A(REG0_REG_18__SCAN_IN), .B(n4371), .S(n4539), .Z(U3503) );
  MUX2_X1 U4924 ( .A(n4373), .B(n4372), .S(n4539), .Z(n4374) );
  OAI21_X1 U4925 ( .B1(n4375), .B2(n4369), .A(n4374), .ZN(U3501) );
  MUX2_X1 U4926 ( .A(REG0_REG_16__SCAN_IN), .B(n4376), .S(n4539), .Z(U3499) );
  MUX2_X1 U4927 ( .A(DATAI_30_), .B(n4377), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4928 ( .A(DATAI_29_), .B(n4378), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4929 ( .A(DATAI_24_), .B(n2689), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4930 ( .A(DATAI_22_), .B(n4379), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4931 ( .A(n4380), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4932 ( .A(n4381), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  INV_X1 U4933 ( .A(n4382), .ZN(n4383) );
  MUX2_X1 U4934 ( .A(DATAI_8_), .B(n4383), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4935 ( .A(DATAI_7_), .B(n4384), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4936 ( .A(DATAI_6_), .B(n4385), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U4937 ( .A(n4386), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4938 ( .A(DATAI_4_), .B(n4387), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4939 ( .A(n4388), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4940 ( .A(n4389), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4941 ( .A(n4390), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4942 ( .A1(n4392), .A2(n4501), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4391), .ZN(n4393) );
  OAI21_X1 U4943 ( .B1(n4391), .B2(n4394), .A(n4393), .ZN(U3261) );
  OAI211_X1 U4944 ( .C1(n4397), .C2(n4396), .A(n4491), .B(n4395), .ZN(n4402)
         );
  OAI211_X1 U4945 ( .C1(n4400), .C2(n4399), .A(n4438), .B(n4398), .ZN(n4401)
         );
  OAI211_X1 U4946 ( .C1(n4495), .C2(n4520), .A(n4402), .B(n4401), .ZN(n4403)
         );
  AOI211_X1 U4947 ( .C1(n4489), .C2(ADDR_REG_9__SCAN_IN), .A(n4404), .B(n4403), 
        .ZN(n4405) );
  INV_X1 U4948 ( .A(n4405), .ZN(U3249) );
  OAI211_X1 U4949 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4407), .A(n4438), .B(n4406), .ZN(n4409) );
  NAND2_X1 U4950 ( .A1(n4409), .A2(n4408), .ZN(n4410) );
  AOI21_X1 U4951 ( .B1(n4489), .B2(ADDR_REG_10__SCAN_IN), .A(n4410), .ZN(n4414) );
  OAI211_X1 U4952 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4412), .A(n4491), .B(n4411), .ZN(n4413) );
  OAI211_X1 U4953 ( .C1(n4495), .C2(n4518), .A(n4414), .B(n4413), .ZN(U3250)
         );
  OAI211_X1 U4954 ( .C1(n4417), .C2(n4416), .A(n4491), .B(n4415), .ZN(n4422)
         );
  OAI211_X1 U4955 ( .C1(n4420), .C2(n4419), .A(n4438), .B(n4418), .ZN(n4421)
         );
  OAI211_X1 U4956 ( .C1(n4495), .C2(n4517), .A(n4422), .B(n4421), .ZN(n4423)
         );
  AOI211_X1 U4957 ( .C1(n4489), .C2(ADDR_REG_11__SCAN_IN), .A(n4424), .B(n4423), .ZN(n4425) );
  INV_X1 U4958 ( .A(n4425), .ZN(U3251) );
  OAI211_X1 U4959 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4427), .A(n4438), .B(n4426), .ZN(n4429) );
  NAND2_X1 U4960 ( .A1(n4429), .A2(n4428), .ZN(n4430) );
  AOI21_X1 U4961 ( .B1(n4489), .B2(ADDR_REG_12__SCAN_IN), .A(n4430), .ZN(n4434) );
  OAI211_X1 U4962 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4432), .A(n4491), .B(n4431), .ZN(n4433) );
  OAI211_X1 U4963 ( .C1(n4495), .C2(n4435), .A(n4434), .B(n4433), .ZN(U3252)
         );
  AOI21_X1 U4964 ( .B1(n4437), .B2(n4514), .A(n4436), .ZN(n4441) );
  OAI21_X1 U4965 ( .B1(n4441), .B2(n4440), .A(n4438), .ZN(n4439) );
  AOI21_X1 U4966 ( .B1(n4441), .B2(n4440), .A(n4439), .ZN(n4443) );
  AOI211_X1 U4967 ( .C1(n4489), .C2(ADDR_REG_13__SCAN_IN), .A(n4443), .B(n4442), .ZN(n4448) );
  OAI211_X1 U4968 ( .C1(n4446), .C2(n4445), .A(n4491), .B(n4444), .ZN(n4447)
         );
  OAI211_X1 U4969 ( .C1(n4495), .C2(n4514), .A(n4448), .B(n4447), .ZN(U3253)
         );
  AOI211_X1 U4970 ( .C1(n2322), .C2(n4450), .A(n4449), .B(n4485), .ZN(n4451)
         );
  AOI211_X1 U4971 ( .C1(n4489), .C2(ADDR_REG_14__SCAN_IN), .A(n4452), .B(n4451), .ZN(n4456) );
  OAI211_X1 U4972 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4454), .A(n4491), .B(n4453), .ZN(n4455) );
  OAI211_X1 U4973 ( .C1(n4495), .C2(n2131), .A(n4456), .B(n4455), .ZN(U3254)
         );
  AOI211_X1 U4974 ( .C1(n4459), .C2(n4458), .A(n4457), .B(n4485), .ZN(n4460)
         );
  AOI211_X1 U4975 ( .C1(n4489), .C2(ADDR_REG_15__SCAN_IN), .A(n4461), .B(n4460), .ZN(n4466) );
  OAI211_X1 U4976 ( .C1(n4464), .C2(n4463), .A(n4491), .B(n4462), .ZN(n4465)
         );
  OAI211_X1 U4977 ( .C1(n4495), .C2(n4513), .A(n4466), .B(n4465), .ZN(U3255)
         );
  AOI221_X1 U4978 ( .B1(n4468), .B2(n4467), .C1(n2509), .C2(n4467), .A(n4485), 
        .ZN(n4469) );
  AOI211_X1 U4979 ( .C1(n4489), .C2(ADDR_REG_16__SCAN_IN), .A(n4470), .B(n4469), .ZN(n4474) );
  OAI221_X1 U4980 ( .B1(n4472), .B2(REG1_REG_16__SCAN_IN), .C1(n4472), .C2(
        n4471), .A(n4491), .ZN(n4473) );
  OAI211_X1 U4981 ( .C1(n4495), .C2(n4512), .A(n4474), .B(n4473), .ZN(U3256)
         );
  AOI221_X1 U4982 ( .B1(n4477), .B2(n4476), .C1(n4475), .C2(n4476), .A(n4485), 
        .ZN(n4478) );
  AOI211_X1 U4983 ( .C1(n4489), .C2(ADDR_REG_17__SCAN_IN), .A(n4479), .B(n4478), .ZN(n4484) );
  OAI221_X1 U4984 ( .B1(n4482), .B2(n4481), .C1(n4482), .C2(n4480), .A(n4491), 
        .ZN(n4483) );
  OAI211_X1 U4985 ( .C1(n4495), .C2(n4511), .A(n4484), .B(n4483), .ZN(U3257)
         );
  OAI211_X1 U4986 ( .C1(n4492), .C2(n2064), .A(n4491), .B(n4490), .ZN(n4493)
         );
  OAI211_X1 U4987 ( .C1(n4495), .C2(n4510), .A(n4494), .B(n4493), .ZN(U3258)
         );
  OAI22_X1 U4988 ( .A1(n4191), .A2(n4498), .B1(n4497), .B2(n4496), .ZN(n4499)
         );
  INV_X1 U4989 ( .A(n4499), .ZN(n4505) );
  AOI22_X1 U4990 ( .A1(n4503), .A2(n4502), .B1(n4501), .B2(n4500), .ZN(n4504)
         );
  OAI211_X1 U4991 ( .C1(n4119), .C2(n4506), .A(n4505), .B(n4504), .ZN(U3282)
         );
  AND2_X1 U4992 ( .A1(D_REG_31__SCAN_IN), .A2(n4507), .ZN(U3291) );
  AND2_X1 U4993 ( .A1(D_REG_30__SCAN_IN), .A2(n4507), .ZN(U3292) );
  AND2_X1 U4994 ( .A1(D_REG_29__SCAN_IN), .A2(n4507), .ZN(U3293) );
  AND2_X1 U4995 ( .A1(D_REG_28__SCAN_IN), .A2(n4507), .ZN(U3294) );
  AND2_X1 U4996 ( .A1(D_REG_27__SCAN_IN), .A2(n4507), .ZN(U3295) );
  AND2_X1 U4997 ( .A1(D_REG_26__SCAN_IN), .A2(n4507), .ZN(U3296) );
  AND2_X1 U4998 ( .A1(D_REG_25__SCAN_IN), .A2(n4507), .ZN(U3297) );
  AND2_X1 U4999 ( .A1(D_REG_24__SCAN_IN), .A2(n4507), .ZN(U3298) );
  AND2_X1 U5000 ( .A1(D_REG_23__SCAN_IN), .A2(n4507), .ZN(U3299) );
  AND2_X1 U5001 ( .A1(D_REG_22__SCAN_IN), .A2(n4507), .ZN(U3300) );
  AND2_X1 U5002 ( .A1(D_REG_21__SCAN_IN), .A2(n4507), .ZN(U3301) );
  AND2_X1 U5003 ( .A1(D_REG_20__SCAN_IN), .A2(n4507), .ZN(U3302) );
  AND2_X1 U5004 ( .A1(D_REG_19__SCAN_IN), .A2(n4507), .ZN(U3303) );
  AND2_X1 U5005 ( .A1(D_REG_18__SCAN_IN), .A2(n4507), .ZN(U3304) );
  AND2_X1 U5006 ( .A1(D_REG_17__SCAN_IN), .A2(n4507), .ZN(U3305) );
  AND2_X1 U5007 ( .A1(D_REG_16__SCAN_IN), .A2(n4507), .ZN(U3306) );
  AND2_X1 U5008 ( .A1(D_REG_15__SCAN_IN), .A2(n4507), .ZN(U3307) );
  AND2_X1 U5009 ( .A1(D_REG_14__SCAN_IN), .A2(n4507), .ZN(U3308) );
  AND2_X1 U5010 ( .A1(D_REG_13__SCAN_IN), .A2(n4507), .ZN(U3309) );
  AND2_X1 U5011 ( .A1(D_REG_12__SCAN_IN), .A2(n4507), .ZN(U3310) );
  AND2_X1 U5012 ( .A1(D_REG_11__SCAN_IN), .A2(n4507), .ZN(U3311) );
  AND2_X1 U5013 ( .A1(D_REG_10__SCAN_IN), .A2(n4507), .ZN(U3312) );
  AND2_X1 U5014 ( .A1(D_REG_9__SCAN_IN), .A2(n4507), .ZN(U3313) );
  AND2_X1 U5015 ( .A1(D_REG_8__SCAN_IN), .A2(n4507), .ZN(U3314) );
  AND2_X1 U5016 ( .A1(D_REG_7__SCAN_IN), .A2(n4507), .ZN(U3315) );
  AND2_X1 U5017 ( .A1(D_REG_6__SCAN_IN), .A2(n4507), .ZN(U3316) );
  AND2_X1 U5018 ( .A1(D_REG_5__SCAN_IN), .A2(n4507), .ZN(U3317) );
  AND2_X1 U5019 ( .A1(D_REG_4__SCAN_IN), .A2(n4507), .ZN(U3318) );
  AND2_X1 U5020 ( .A1(D_REG_3__SCAN_IN), .A2(n4507), .ZN(U3319) );
  AND2_X1 U5021 ( .A1(D_REG_2__SCAN_IN), .A2(n4507), .ZN(U3320) );
  OAI21_X1 U5022 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4508), .ZN(
        n4509) );
  INV_X1 U5023 ( .A(n4509), .ZN(U3329) );
  AOI22_X1 U5024 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n4670), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5025 ( .A1(STATE_REG_SCAN_IN), .A2(n4511), .B1(n2532), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5026 ( .A(DATAI_16_), .ZN(n4702) );
  AOI22_X1 U5027 ( .A1(STATE_REG_SCAN_IN), .A2(n4512), .B1(n4702), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5028 ( .A(DATAI_15_), .ZN(n4580) );
  AOI22_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4580), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5030 ( .A(DATAI_14_), .ZN(n4568) );
  AOI22_X1 U5031 ( .A1(STATE_REG_SCAN_IN), .A2(n2131), .B1(n4568), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5032 ( .A1(STATE_REG_SCAN_IN), .A2(n4514), .B1(n2329), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5033 ( .A1(U3149), .A2(n4515), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4516) );
  INV_X1 U5034 ( .A(n4516), .ZN(U3340) );
  INV_X1 U5035 ( .A(DATAI_11_), .ZN(n4679) );
  AOI22_X1 U5036 ( .A1(STATE_REG_SCAN_IN), .A2(n4517), .B1(n4679), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5037 ( .A(DATAI_10_), .ZN(n4720) );
  AOI22_X1 U5038 ( .A1(STATE_REG_SCAN_IN), .A2(n4518), .B1(n4720), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5039 ( .A(DATAI_9_), .ZN(n4519) );
  AOI22_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .B1(n4519), .B2(U3149), 
        .ZN(U3343) );
  OAI211_X1 U5041 ( .C1(n4524), .C2(n4523), .A(n4522), .B(n4521), .ZN(n4525)
         );
  INV_X1 U5042 ( .A(n4525), .ZN(n4541) );
  AOI22_X1 U5043 ( .A1(n4539), .A2(n4541), .B1(n2370), .B2(n4537), .ZN(U3467)
         );
  INV_X1 U5044 ( .A(n4526), .ZN(n4528) );
  AOI211_X1 U5045 ( .C1(n4530), .C2(n4529), .A(n4528), .B(n4527), .ZN(n4542)
         );
  AOI22_X1 U5046 ( .A1(n4539), .A2(n4542), .B1(n2338), .B2(n4537), .ZN(U3475)
         );
  NAND3_X1 U5047 ( .A1(n4533), .A2(n4532), .A3(n4531), .ZN(n4534) );
  INV_X1 U5048 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5049 ( .A1(n4539), .A2(n4544), .B1(n4538), .B2(n4537), .ZN(U3481)
         );
  AOI22_X1 U5050 ( .A1(n4545), .A2(n4541), .B1(n4540), .B2(n4543), .ZN(U3518)
         );
  AOI22_X1 U5051 ( .A1(n4545), .A2(n4542), .B1(n2343), .B2(n4543), .ZN(U3522)
         );
  AOI22_X1 U5052 ( .A1(n4545), .A2(n4544), .B1(n2419), .B2(n4543), .ZN(U3525)
         );
  AOI22_X1 U5053 ( .A1(n4547), .A2(keyinput_g44), .B1(keyinput_g11), .B2(n2561), .ZN(n4546) );
  OAI221_X1 U5054 ( .B1(n4547), .B2(keyinput_g44), .C1(n2561), .C2(
        keyinput_g11), .A(n4546), .ZN(n4556) );
  INV_X1 U5055 ( .A(DATAI_4_), .ZN(n4549) );
  AOI22_X1 U5056 ( .A1(n4549), .A2(keyinput_g27), .B1(n2439), .B2(keyinput_g23), .ZN(n4548) );
  OAI221_X1 U5057 ( .B1(n4549), .B2(keyinput_g27), .C1(n2439), .C2(
        keyinput_g23), .A(n4548), .ZN(n4555) );
  AOI22_X1 U5058 ( .A1(n4551), .A2(keyinput_g0), .B1(n4667), .B2(keyinput_g12), 
        .ZN(n4550) );
  OAI221_X1 U5059 ( .B1(n4551), .B2(keyinput_g0), .C1(n4667), .C2(keyinput_g12), .A(n4550), .ZN(n4554) );
  AOI22_X1 U5060 ( .A1(n4678), .A2(keyinput_g5), .B1(n2308), .B2(keyinput_g43), 
        .ZN(n4552) );
  OAI221_X1 U5061 ( .B1(n4678), .B2(keyinput_g5), .C1(n2308), .C2(keyinput_g43), .A(n4552), .ZN(n4553) );
  NOR4_X1 U5062 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4593)
         );
  AOI22_X1 U5063 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(n4558), .B2(
        keyinput_g46), .ZN(n4557) );
  OAI221_X1 U5064 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(n4558), .C2(
        keyinput_g46), .A(n4557), .ZN(n4566) );
  AOI22_X1 U5065 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput_g49), .ZN(n4559) );
  OAI221_X1 U5066 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4559), .ZN(n4565) );
  AOI22_X1 U5067 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n4560) );
  OAI221_X1 U5068 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_g41), .A(n4560), .ZN(n4564) );
  XNOR2_X1 U5069 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4562) );
  XNOR2_X1 U5070 ( .A(DATAI_7_), .B(keyinput_g24), .ZN(n4561) );
  NAND2_X1 U5071 ( .A1(n4562), .A2(n4561), .ZN(n4563) );
  NOR4_X1 U5072 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4592)
         );
  AOI22_X1 U5073 ( .A1(n4568), .A2(keyinput_g17), .B1(n4692), .B2(keyinput_g35), .ZN(n4567) );
  OAI221_X1 U5074 ( .B1(n4568), .B2(keyinput_g17), .C1(n4692), .C2(
        keyinput_g35), .A(n4567), .ZN(n4576) );
  XNOR2_X1 U5075 ( .A(DATAI_30_), .B(keyinput_g1), .ZN(n4572) );
  XNOR2_X1 U5076 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4571) );
  XNOR2_X1 U5077 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .ZN(n4570) );
  XNOR2_X1 U5078 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4569) );
  NAND4_X1 U5079 ( .A1(n4572), .A2(n4571), .A3(n4570), .A4(n4569), .ZN(n4575)
         );
  XNOR2_X1 U5080 ( .A(keyinput_g40), .B(n3701), .ZN(n4574) );
  XNOR2_X1 U5081 ( .A(keyinput_g18), .B(n2329), .ZN(n4573) );
  NOR4_X1 U5082 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4591)
         );
  AOI22_X1 U5083 ( .A1(n4578), .A2(keyinput_g39), .B1(keyinput_g14), .B2(n2532), .ZN(n4577) );
  OAI221_X1 U5084 ( .B1(n4578), .B2(keyinput_g39), .C1(n2532), .C2(
        keyinput_g14), .A(n4577), .ZN(n4589) );
  AOI22_X1 U5085 ( .A1(n4581), .A2(keyinput_g36), .B1(keyinput_g16), .B2(n4580), .ZN(n4579) );
  OAI221_X1 U5086 ( .B1(n4581), .B2(keyinput_g36), .C1(n4580), .C2(
        keyinput_g16), .A(n4579), .ZN(n4588) );
  AOI22_X1 U5087 ( .A1(U3149), .A2(keyinput_g32), .B1(keyinput_g6), .B2(n4583), 
        .ZN(n4582) );
  OAI221_X1 U5088 ( .B1(U3149), .B2(keyinput_g32), .C1(n4583), .C2(keyinput_g6), .A(n4582), .ZN(n4587) );
  XOR2_X1 U5089 ( .A(n2618), .B(keyinput_g3), .Z(n4585) );
  XNOR2_X1 U5090 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4584) );
  NAND2_X1 U5091 ( .A1(n4585), .A2(n4584), .ZN(n4586) );
  NOR4_X1 U5092 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4590)
         );
  AND4_X1 U5093 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4725)
         );
  OAI22_X1 U5094 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(keyinput_g38), .B2(REG3_REG_3__SCAN_IN), .ZN(n4594) );
  AOI221_X1 U5095 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        REG3_REG_3__SCAN_IN), .C2(keyinput_g38), .A(n4594), .ZN(n4601) );
  OAI22_X1 U5096 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_18_), .B2(
        keyinput_g13), .ZN(n4595) );
  AOI221_X1 U5097 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(keyinput_g13), .C2(
        DATAI_18_), .A(n4595), .ZN(n4600) );
  OAI22_X1 U5098 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(DATAI_12_), .B2(keyinput_g19), .ZN(n4596) );
  AOI221_X1 U5099 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        keyinput_g19), .C2(DATAI_12_), .A(n4596), .ZN(n4599) );
  OAI22_X1 U5100 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(
        keyinput_g33), .B2(REG3_REG_7__SCAN_IN), .ZN(n4597) );
  AOI221_X1 U5101 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_g33), .A(n4597), .ZN(n4598) );
  NAND4_X1 U5102 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4628)
         );
  OAI22_X1 U5103 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_g45), .B1(DATAI_22_), .B2(keyinput_g9), .ZN(n4602) );
  AOI221_X1 U5104 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g9), .C2(DATAI_22_), .A(n4602), .ZN(n4608) );
  OAI22_X1 U5105 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_g53), .B1(DATAI_29_), .B2(keyinput_g2), .ZN(n4603) );
  AOI221_X1 U5106 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_g53), .C1(
        keyinput_g2), .C2(DATAI_29_), .A(n4603), .ZN(n4607) );
  OAI22_X1 U5107 ( .A1(DATAI_27_), .A2(keyinput_g4), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n4604) );
  AOI221_X1 U5108 ( .B1(DATAI_27_), .B2(keyinput_g4), .C1(keyinput_g8), .C2(
        DATAI_23_), .A(n4604), .ZN(n4606) );
  XNOR2_X1 U5109 ( .A(DATAI_1_), .B(keyinput_g30), .ZN(n4605) );
  NAND4_X1 U5110 ( .A1(n4608), .A2(n4607), .A3(n4606), .A4(n4605), .ZN(n4627)
         );
  OAI22_X1 U5111 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(keyinput_g22), .B2(
        DATAI_9_), .ZN(n4609) );
  AOI221_X1 U5112 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(DATAI_9_), .C2(
        keyinput_g22), .A(n4609), .ZN(n4616) );
  OAI22_X1 U5113 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_g62), .B1(keyinput_g47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4610) );
  AOI221_X1 U5114 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_g62), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_g47), .A(n4610), .ZN(n4615) );
  OAI22_X1 U5115 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(DATAI_16_), .B2(keyinput_g15), .ZN(n4611) );
  AOI221_X1 U5116 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g15), .C2(DATAI_16_), .A(n4611), .ZN(n4614) );
  OAI22_X1 U5117 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_g48), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .ZN(n4612) );
  AOI221_X1 U5118 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g37), .C2(REG3_REG_10__SCAN_IN), .A(n4612), .ZN(n4613) );
  NAND4_X1 U5119 ( .A1(n4616), .A2(n4615), .A3(n4614), .A4(n4613), .ZN(n4626)
         );
  OAI22_X1 U5120 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_g57), .B1(keyinput_g31), .B2(DATAI_0_), .ZN(n4617) );
  AOI221_X1 U5121 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_g57), .C1(DATAI_0_), 
        .C2(keyinput_g31), .A(n4617), .ZN(n4624) );
  OAI22_X1 U5122 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(keyinput_g25), .B2(DATAI_6_), .ZN(n4618) );
  AOI221_X1 U5123 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(DATAI_6_), 
        .C2(keyinput_g25), .A(n4618), .ZN(n4623) );
  OAI22_X1 U5124 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_g60), .B1(keyinput_g26), .B2(DATAI_5_), .ZN(n4619) );
  AOI221_X1 U5125 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_g60), .C1(DATAI_5_), 
        .C2(keyinput_g26), .A(n4619), .ZN(n4622) );
  OAI22_X1 U5126 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .ZN(n4620) );
  AOI221_X1 U5127 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g50), .C2(REG3_REG_4__SCAN_IN), .A(n4620), .ZN(n4621) );
  NAND4_X1 U5128 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4625)
         );
  NOR4_X1 U5129 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4724)
         );
  AOI22_X1 U5130 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4629) );
  OAI221_X1 U5131 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4629), .ZN(n4636) );
  AOI22_X1 U5132 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4630) );
  OAI221_X1 U5133 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(REG3_REG_3__SCAN_IN), 
        .C2(keyinput_f38), .A(n4630), .ZN(n4635) );
  AOI22_X1 U5134 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(DATAI_15_), .B2(
        keyinput_f16), .ZN(n4631) );
  OAI221_X1 U5135 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(DATAI_15_), .C2(
        keyinput_f16), .A(n4631), .ZN(n4634) );
  AOI22_X1 U5136 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_f33), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .ZN(n4632) );
  OAI221_X1 U5137 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_f33), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_f51), .A(n4632), .ZN(n4633) );
  NOR4_X1 U5138 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4663)
         );
  AOI22_X1 U5139 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n4637) );
  OAI221_X1 U5140 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4637), .ZN(n4643) );
  AOI22_X1 U5141 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4638) );
  OAI221_X1 U5142 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4638), .ZN(n4642) );
  AOI22_X1 U5143 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n4639) );
  OAI221_X1 U5144 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n4639), .ZN(n4641) );
  XOR2_X1 U5145 ( .A(DATAI_1_), .B(keyinput_f30), .Z(n4640) );
  NOR4_X1 U5146 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4662)
         );
  AOI22_X1 U5147 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(REG3_REG_23__SCAN_IN), 
        .B2(keyinput_f36), .ZN(n4644) );
  OAI221_X1 U5148 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4644), .ZN(n4651) );
  AOI22_X1 U5149 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_f62), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_f63), .ZN(n4645) );
  OAI221_X1 U5150 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_f62), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_f63), .A(n4645), .ZN(n4650) );
  AOI22_X1 U5151 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(U3149), 
        .B2(keyinput_f32), .ZN(n4646) );
  OAI221_X1 U5152 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(U3149), 
        .C2(keyinput_f32), .A(n4646), .ZN(n4649) );
  AOI22_X1 U5153 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_13_), .B2(
        keyinput_f18), .ZN(n4647) );
  OAI221_X1 U5154 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_13_), .C2(
        keyinput_f18), .A(n4647), .ZN(n4648) );
  NOR4_X1 U5155 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n4661)
         );
  AOI22_X1 U5156 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_f56), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n4652) );
  OAI221_X1 U5157 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_f56), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n4652), .ZN(n4659) );
  AOI22_X1 U5158 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4653) );
  OAI221_X1 U5159 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4653), .ZN(n4658) );
  AOI22_X1 U5160 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(DATAI_8_), .B2(
        keyinput_f23), .ZN(n4654) );
  OAI221_X1 U5161 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(DATAI_8_), .C2(
        keyinput_f23), .A(n4654), .ZN(n4657) );
  AOI22_X1 U5162 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(IR_REG_2__SCAN_IN), 
        .B2(keyinput_f57), .ZN(n4655) );
  OAI221_X1 U5163 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_f57), .A(n4655), .ZN(n4656) );
  NOR4_X1 U5164 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4660)
         );
  NAND4_X1 U5165 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4718)
         );
  AOI22_X1 U5166 ( .A1(n4665), .A2(keyinput_f47), .B1(keyinput_f4), .B2(n2607), 
        .ZN(n4664) );
  OAI221_X1 U5167 ( .B1(n4665), .B2(keyinput_f47), .C1(n2607), .C2(keyinput_f4), .A(n4664), .ZN(n4676) );
  AOI22_X1 U5168 ( .A1(n2330), .A2(keyinput_f54), .B1(keyinput_f12), .B2(n4667), .ZN(n4666) );
  OAI221_X1 U5169 ( .B1(n2330), .B2(keyinput_f54), .C1(n4667), .C2(
        keyinput_f12), .A(n4666), .ZN(n4675) );
  AOI22_X1 U5170 ( .A1(n4670), .A2(keyinput_f13), .B1(n4669), .B2(keyinput_f53), .ZN(n4668) );
  OAI221_X1 U5171 ( .B1(n4670), .B2(keyinput_f13), .C1(n4669), .C2(
        keyinput_f53), .A(n4668), .ZN(n4674) );
  XOR2_X1 U5172 ( .A(n2561), .B(keyinput_f11), .Z(n4672) );
  XNOR2_X1 U5173 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4671) );
  NAND2_X1 U5174 ( .A1(n4672), .A2(n4671), .ZN(n4673) );
  NOR4_X1 U5175 ( .A1(n4676), .A2(n4675), .A3(n4674), .A4(n4673), .ZN(n4716)
         );
  AOI22_X1 U5176 ( .A1(n4679), .A2(keyinput_f20), .B1(n4678), .B2(keyinput_f5), 
        .ZN(n4677) );
  OAI221_X1 U5177 ( .B1(n4679), .B2(keyinput_f20), .C1(n4678), .C2(keyinput_f5), .A(n4677), .ZN(n4688) );
  AOI22_X1 U5178 ( .A1(n2618), .A2(keyinput_f3), .B1(n4681), .B2(keyinput_f45), 
        .ZN(n4680) );
  OAI221_X1 U5179 ( .B1(n2618), .B2(keyinput_f3), .C1(n4681), .C2(keyinput_f45), .A(n4680), .ZN(n4687) );
  XOR2_X1 U5180 ( .A(n2308), .B(keyinput_f43), .Z(n4685) );
  XNOR2_X1 U5181 ( .A(keyinput_f25), .B(DATAI_6_), .ZN(n4684) );
  XNOR2_X1 U5182 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n4683) );
  XNOR2_X1 U5183 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4682) );
  NAND4_X1 U5184 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4686)
         );
  NOR3_X1 U5185 ( .A1(n4688), .A2(n4687), .A3(n4686), .ZN(n4715) );
  AOI22_X1 U5186 ( .A1(n2523), .A2(keyinput_f48), .B1(n4690), .B2(keyinput_f49), .ZN(n4689) );
  OAI221_X1 U5187 ( .B1(n2523), .B2(keyinput_f48), .C1(n4690), .C2(
        keyinput_f49), .A(n4689), .ZN(n4700) );
  INV_X1 U5188 ( .A(DATAI_2_), .ZN(n4693) );
  AOI22_X1 U5189 ( .A1(n4693), .A2(keyinput_f29), .B1(n4692), .B2(keyinput_f35), .ZN(n4691) );
  OAI221_X1 U5190 ( .B1(n4693), .B2(keyinput_f29), .C1(n4692), .C2(
        keyinput_f35), .A(n4691), .ZN(n4699) );
  XNOR2_X1 U5191 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_f41), .ZN(n4697) );
  XNOR2_X1 U5192 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_f52), .ZN(n4696) );
  XNOR2_X1 U5193 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4695) );
  XNOR2_X1 U5194 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_f34), .ZN(n4694) );
  NAND4_X1 U5195 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4698)
         );
  NOR3_X1 U5196 ( .A1(n4700), .A2(n4699), .A3(n4698), .ZN(n4714) );
  AOI22_X1 U5197 ( .A1(n4702), .A2(keyinput_f15), .B1(n2532), .B2(keyinput_f14), .ZN(n4701) );
  OAI221_X1 U5198 ( .B1(n4702), .B2(keyinput_f15), .C1(n2532), .C2(
        keyinput_f14), .A(n4701), .ZN(n4712) );
  AOI22_X1 U5199 ( .A1(n4705), .A2(keyinput_f37), .B1(keyinput_f26), .B2(n4704), .ZN(n4703) );
  OAI221_X1 U5200 ( .B1(n4705), .B2(keyinput_f37), .C1(n4704), .C2(
        keyinput_f26), .A(n4703), .ZN(n4711) );
  XNOR2_X1 U5201 ( .A(DATAI_21_), .B(keyinput_f10), .ZN(n4709) );
  XNOR2_X1 U5202 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4708) );
  XNOR2_X1 U5203 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_f39), .ZN(n4707) );
  XNOR2_X1 U5204 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4706) );
  NAND4_X1 U5205 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4710)
         );
  NOR3_X1 U5206 ( .A1(n4712), .A2(n4711), .A3(n4710), .ZN(n4713) );
  NAND4_X1 U5207 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4717)
         );
  OAI22_X1 U5208 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(n4718), .B2(n4717), 
        .ZN(n4722) );
  NAND3_X1 U5209 ( .A1(n4720), .A2(keyinput_g21), .A3(n4722), .ZN(n4719) );
  OAI21_X1 U5210 ( .B1(keyinput_g21), .B2(n4720), .A(n4719), .ZN(n4721) );
  OAI21_X1 U5211 ( .B1(keyinput_f21), .B2(n4722), .A(n4721), .ZN(n4723) );
  AOI21_X1 U5212 ( .B1(n4725), .B2(n4724), .A(n4723), .ZN(n4728) );
  AOI22_X1 U5213 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4727) );
  XNOR2_X1 U5214 ( .A(n4728), .B(n4727), .ZN(U3352) );
  XNOR2_X1 U2346 ( .A(n2094), .B(n2635), .ZN(n2637) );
  BUF_X2 U2285 ( .A(n2378), .Z(n2619) );
  NAND2_X1 U2307 ( .A1(n2811), .A2(n2861), .ZN(n3692) );
  CLKBUF_X1 U2323 ( .A(n3692), .Z(n2043) );
  CLKBUF_X1 U2347 ( .A(n2369), .Z(n3402) );
endmodule

