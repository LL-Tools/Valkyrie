

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10068;

  AOI22_X1 U4777 ( .A1(n6693), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n6698), .B2(
        n6692), .ZN(n9869) );
  AND2_X1 U4778 ( .A1(n7608), .A2(n7609), .ZN(n7507) );
  NAND2_X1 U4779 ( .A1(n8877), .A2(n7181), .ZN(n8822) );
  AND3_X1 U4780 ( .A1(n5018), .A2(n5017), .A3(n5016), .ZN(n7118) );
  CLKBUF_X2 U4781 ( .A(n5037), .Z(n5652) );
  INV_X1 U4782 ( .A(n5019), .ZN(n4732) );
  NAND2_X1 U4783 ( .A1(n6170), .A2(n6167), .ZN(n7483) );
  XNOR2_X1 U4784 ( .A(n4980), .B(n4979), .ZN(n8810) );
  CLKBUF_X2 U4785 ( .A(n5890), .Z(n6020) );
  INV_X1 U4786 ( .A(n4963), .ZN(n9516) );
  OR2_X1 U4787 ( .A1(n7679), .A2(n4510), .ZN(n4509) );
  NOR2_X1 U4788 ( .A1(n4976), .A2(n4968), .ZN(n4981) );
  OAI21_X1 U4789 ( .B1(n8033), .B2(n8341), .A(n8032), .ZN(n8034) );
  AND2_X1 U4790 ( .A1(n4924), .A2(n4816), .ZN(n5776) );
  INV_X1 U4791 ( .A(n8717), .ZN(n5462) );
  INV_X1 U4792 ( .A(n8164), .ZN(n7847) );
  INV_X1 U4793 ( .A(n5817), .ZN(n5818) );
  NOR2_X1 U4794 ( .A1(n9869), .A2(n9870), .ZN(n9868) );
  INV_X1 U4795 ( .A(n7675), .ZN(n7691) );
  CLKBUF_X2 U4796 ( .A(n5825), .Z(n7526) );
  INV_X1 U4797 ( .A(n7526), .ZN(n6102) );
  XNOR2_X1 U4798 ( .A(n5357), .B(n5358), .ZN(n8454) );
  XNOR2_X1 U4799 ( .A(n5195), .B(n5193), .ZN(n7279) );
  INV_X1 U4800 ( .A(n6870), .ZN(n7181) );
  AND3_X2 U4801 ( .A1(n5085), .A2(n5084), .A3(n5083), .ZN(n8819) );
  INV_X1 U4802 ( .A(n6365), .ZN(n8624) );
  AND2_X1 U4803 ( .A1(n5162), .A2(n5161), .ZN(n7133) );
  INV_X1 U4804 ( .A(n6731), .ZN(n9656) );
  NAND4_X2 U4805 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n8126)
         );
  INV_X1 U4806 ( .A(n6924), .ZN(n7167) );
  OR2_X1 U4807 ( .A1(n4967), .A2(n4966), .ZN(n8878) );
  AOI21_X1 U4808 ( .B1(n7089), .B2(n7094), .A(n7956), .ZN(n6120) );
  OAI21_X2 U4809 ( .B1(n7920), .B2(n7923), .A(n7921), .ZN(n7753) );
  NAND2_X2 U4810 ( .A1(n9561), .A2(n9562), .ZN(n9560) );
  AOI21_X2 U4811 ( .B1(n4657), .B2(n9333), .A(n4656), .ZN(n9363) );
  OAI21_X1 U4812 ( .B1(n8282), .B2(n7621), .A(n7498), .ZN(n8262) );
  NAND2_X2 U4813 ( .A1(n7279), .A2(n7280), .ZN(n7278) );
  NAND2_X2 U4814 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  NAND3_X2 U4815 ( .A1(n9045), .A2(n8078), .A3(n4579), .ZN(n4636) );
  XNOR2_X2 U4816 ( .A(n5148), .B(SI_6_), .ZN(n5146) );
  NAND2_X2 U4817 ( .A1(n4540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  NOR2_X2 U4818 ( .A1(n5977), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5989) );
  NOR2_X2 U4819 ( .A1(n9162), .A2(n9379), .ZN(n9136) );
  NAND2_X2 U4820 ( .A1(n4474), .A2(n4718), .ZN(n5357) );
  XNOR2_X2 U4821 ( .A(n5251), .B(n5252), .ZN(n6393) );
  NOR2_X2 U4822 ( .A1(n7100), .A2(n7573), .ZN(n7099) );
  BUF_X1 U4823 ( .A(n5740), .Z(n4271) );
  BUF_X1 U4824 ( .A(n5740), .Z(n4272) );
  NAND2_X1 U4825 ( .A1(n9512), .A2(n4963), .ZN(n5740) );
  NAND2_X1 U4826 ( .A1(n4730), .A2(n6940), .ZN(n4273) );
  NAND2_X1 U4827 ( .A1(n4730), .A2(n6940), .ZN(n4274) );
  CLKBUF_X1 U4828 ( .A(n5629), .Z(n4276) );
  AOI21_X2 U4829 ( .B1(n9772), .B2(n6121), .A(n6120), .ZN(n7240) );
  XNOR2_X2 U4830 ( .A(n5120), .B(SI_5_), .ZN(n5118) );
  OAI21_X2 U4831 ( .B1(n6251), .B2(n4708), .A(n4706), .ZN(n7541) );
  OAI21_X2 U4832 ( .B1(n8123), .B2(n7549), .A(n7496), .ZN(n6251) );
  AOI21_X2 U4833 ( .B1(n7880), .B2(n7876), .A(n7878), .ZN(n7760) );
  OAI22_X2 U4834 ( .A1(n7813), .A2(n7812), .B1(n9547), .B2(n7725), .ZN(n7880)
         );
  CLKBUF_X1 U4835 ( .A(n8096), .Z(n8097) );
  MUX2_X1 U4836 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6208), .S(n4275), .Z(n6198)
         );
  NAND2_X1 U4837 ( .A1(n7456), .A2(n7455), .ZN(n7720) );
  NAND2_X1 U4838 ( .A1(n7136), .A2(n4323), .ZN(n8828) );
  AOI21_X1 U4839 ( .B1(n6115), .B2(n6951), .A(n6114), .ZN(n6808) );
  INV_X1 U4840 ( .A(n7094), .ZN(n9772) );
  XNOR2_X1 U4841 ( .A(n5197), .B(n5196), .ZN(n6359) );
  CLKBUF_X1 U4842 ( .A(n8815), .Z(n4391) );
  CLKBUF_X3 U4843 ( .A(n6267), .Z(n7796) );
  NOR2_X2 U4844 ( .A1(n6581), .A2(n6599), .ZN(n6601) );
  CLKBUF_X1 U4845 ( .A(n5845), .Z(n4418) );
  AND4_X1 U4846 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n7473)
         );
  NAND2_X1 U4847 ( .A1(n5805), .A2(n4457), .ZN(n5825) );
  INV_X2 U4848 ( .A(n5047), .ZN(n5661) );
  INV_X1 U4849 ( .A(n6259), .ZN(n7559) );
  CLKBUF_X2 U4850 ( .A(n6156), .Z(n4398) );
  NAND2_X1 U4851 ( .A1(n6259), .A2(n5782), .ZN(n6805) );
  AND2_X1 U4852 ( .A1(n7532), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5820) );
  AND2_X1 U4853 ( .A1(n4956), .A2(n9507), .ZN(n4959) );
  NAND2_X1 U4854 ( .A1(n4608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5007) );
  INV_X1 U4855 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U4856 ( .A1(n9364), .A2(n9706), .ZN(n4435) );
  MUX2_X1 U4857 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n6208), .S(n9817), .Z(n6209)
         );
  AND2_X1 U4858 ( .A1(n8598), .A2(n5672), .ZN(n7709) );
  AOI21_X1 U4859 ( .B1(n7794), .B2(n7793), .A(n7792), .ZN(n7798) );
  AOI21_X1 U4860 ( .B1(n6158), .B2(n9748), .A(n6157), .ZN(n8113) );
  OR2_X1 U4861 ( .A1(n8809), .A2(n8808), .ZN(n4677) );
  NAND2_X1 U4862 ( .A1(n4512), .A2(n4509), .ZN(n7689) );
  AND2_X1 U4863 ( .A1(n7684), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U4864 ( .A1(n8543), .A2(n5499), .ZN(n8487) );
  NAND2_X1 U4865 ( .A1(n9191), .A2(n9065), .ZN(n9173) );
  NAND2_X1 U4866 ( .A1(n4735), .A2(n4733), .ZN(n8526) );
  NAND2_X1 U4867 ( .A1(n9207), .A2(n4331), .ZN(n9191) );
  INV_X1 U4868 ( .A(n4736), .ZN(n4735) );
  AND2_X1 U4869 ( .A1(n9715), .A2(n4436), .ZN(n8068) );
  NAND2_X1 U4870 ( .A1(n8572), .A2(n4720), .ZN(n4474) );
  NAND2_X1 U4871 ( .A1(n6131), .A2(n6130), .ZN(n8256) );
  NAND2_X1 U4872 ( .A1(n9311), .A2(n4645), .ZN(n9294) );
  OR2_X1 U4873 ( .A1(n8685), .A2(n8722), .ZN(n4663) );
  OR2_X1 U4874 ( .A1(n4830), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U4875 ( .A1(n7278), .A2(n5222), .ZN(n7265) );
  XNOR2_X1 U4876 ( .A(n7720), .B(n7473), .ZN(n7458) );
  NAND2_X1 U4877 ( .A1(n7969), .A2(n7970), .ZN(n7991) );
  NAND2_X1 U4878 ( .A1(n4752), .A2(n5117), .ZN(n6865) );
  INV_X2 U4879 ( .A(n6233), .ZN(n7950) );
  AND2_X1 U4880 ( .A1(n6320), .A2(n6319), .ZN(n7189) );
  AOI21_X1 U4881 ( .B1(n4895), .B2(n4898), .A(n4893), .ZN(n4892) );
  AND2_X1 U4882 ( .A1(n4727), .A2(n4719), .ZN(n4718) );
  OAI21_X1 U4883 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8660) );
  NAND2_X1 U4884 ( .A1(n6279), .A2(n6974), .ZN(n6977) );
  NAND2_X1 U4885 ( .A1(n8812), .A2(n8828), .ZN(n7248) );
  NAND2_X1 U4886 ( .A1(n7054), .A2(n7053), .ZN(n7078) );
  AND2_X1 U4887 ( .A1(n7773), .A2(n6275), .ZN(n7858) );
  NAND2_X1 U4888 ( .A1(n7105), .A2(n7573), .ZN(n7104) );
  NAND2_X1 U4889 ( .A1(n5848), .A2(n7584), .ZN(n7105) );
  AND2_X1 U4890 ( .A1(n6671), .A2(n6272), .ZN(n7775) );
  NAND2_X1 U4891 ( .A1(n4673), .A2(n6662), .ZN(n8630) );
  NAND2_X1 U4892 ( .A1(n5265), .A2(n5264), .ZN(n8581) );
  XNOR2_X1 U4893 ( .A(n5096), .B(n4475), .ZN(n6742) );
  NAND2_X1 U4894 ( .A1(n5920), .A2(n5919), .ZN(n9802) );
  INV_X2 U4895 ( .A(n5832), .ZN(n5833) );
  INV_X2 U4896 ( .A(n9833), .ZN(n4275) );
  NAND2_X1 U4897 ( .A1(n5126), .A2(n5125), .ZN(n6924) );
  XNOR2_X1 U4898 ( .A(n5031), .B(n5658), .ZN(n5035) );
  INV_X2 U4899 ( .A(n5136), .ZN(n5680) );
  AND2_X1 U4900 ( .A1(n5189), .A2(n5188), .ZN(n7153) );
  NAND2_X1 U4901 ( .A1(n4599), .A2(n5172), .ZN(n5197) );
  NAND2_X1 U4902 ( .A1(n5226), .A2(n4937), .ZN(n5228) );
  INV_X2 U4903 ( .A(n4418), .ZN(n7525) );
  INV_X1 U4904 ( .A(n6267), .ZN(n7750) );
  INV_X1 U4905 ( .A(n6982), .ZN(n9746) );
  NAND2_X1 U4906 ( .A1(n4317), .A2(n5840), .ZN(n7957) );
  NOR2_X1 U4907 ( .A1(n6023), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6033) );
  NAND2_X2 U4908 ( .A1(n6261), .A2(n6262), .ZN(n6267) );
  NAND2_X1 U4909 ( .A1(n5805), .A2(n4412), .ZN(n5845) );
  CLKBUF_X1 U4910 ( .A(n5391), .Z(n5645) );
  INV_X1 U4911 ( .A(n4672), .ZN(n8814) );
  INV_X2 U4912 ( .A(n5061), .ZN(n8716) );
  NAND2_X1 U4913 ( .A1(n4637), .A2(n5003), .ZN(n5107) );
  INV_X1 U4914 ( .A(n4959), .ZN(n9512) );
  NAND2_X1 U4915 ( .A1(n6373), .A2(n4457), .ZN(n5061) );
  NAND2_X1 U4916 ( .A1(n4638), .A2(n5000), .ZN(n5077) );
  NAND2_X1 U4917 ( .A1(n5764), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  AND2_X1 U4918 ( .A1(n5711), .A2(n5710), .ZN(n4975) );
  AOI21_X1 U4919 ( .B1(n4652), .B2(n4655), .A(n5169), .ZN(n4651) );
  XNOR2_X1 U4920 ( .A(n6162), .B(n6161), .ZN(n7479) );
  OAI21_X1 U4921 ( .B1(n4958), .B2(n4953), .A(n4952), .ZN(n4956) );
  XNOR2_X1 U4922 ( .A(n5780), .B(n5779), .ZN(n8065) );
  NAND2_X1 U4923 ( .A1(n4985), .A2(n4984), .ZN(n5732) );
  MUX2_X1 U4924 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6169), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6170) );
  XNOR2_X1 U4925 ( .A(n5767), .B(n5766), .ZN(n5782) );
  AOI21_X1 U4926 ( .B1(n6010), .B2(P2_IR_REG_31__SCAN_IN), .A(n4844), .ZN(
        n4843) );
  OR2_X1 U4927 ( .A1(n5796), .A2(n8441), .ZN(n5798) );
  XNOR2_X1 U4928 ( .A(n5714), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8863) );
  XNOR2_X1 U4929 ( .A(n5007), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5711) );
  OAI21_X1 U4930 ( .B1(n6010), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U4931 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U4932 ( .A1(n5005), .A2(n4950), .ZN(n4958) );
  NAND2_X1 U4933 ( .A1(n6165), .A2(n6166), .ZN(n7452) );
  XNOR2_X1 U4934 ( .A(n5858), .B(n5857), .ZN(n6635) );
  AND2_X1 U4936 ( .A1(n4539), .A2(n5789), .ZN(n4538) );
  INV_X1 U4937 ( .A(n4990), .ZN(n4457) );
  AND2_X1 U4938 ( .A1(n4319), .A2(n5797), .ZN(n4539) );
  INV_X1 U4939 ( .A(n6488), .ZN(n6545) );
  AND3_X1 U4940 ( .A1(n4924), .A2(n5775), .A3(n4923), .ZN(n6188) );
  AND2_X1 U4941 ( .A1(n4778), .A2(n4777), .ZN(n6488) );
  AND2_X1 U4942 ( .A1(n4930), .A2(n4910), .ZN(n4909) );
  AND2_X1 U4943 ( .A1(n5758), .A2(n5757), .ZN(n4849) );
  NOR2_X1 U4944 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  OR2_X1 U4945 ( .A1(n5804), .A2(n8441), .ZN(n5826) );
  NAND2_X1 U4946 ( .A1(n4951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U4947 ( .A1(n4938), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4953) );
  CLKBUF_X2 U4948 ( .A(n5803), .Z(n5804) );
  AND2_X1 U4949 ( .A1(n4943), .A2(n4944), .ZN(n4758) );
  NAND2_X1 U4950 ( .A1(n4908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  AND2_X1 U4951 ( .A1(n5081), .A2(n4781), .ZN(n5010) );
  INV_X1 U4952 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5972) );
  NOR2_X1 U4953 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4780) );
  NOR2_X1 U4954 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4943) );
  INV_X1 U4955 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6161) );
  INV_X1 U4956 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6163) );
  INV_X1 U4957 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4977) );
  INV_X1 U4958 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4979) );
  NOR2_X1 U4959 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5772) );
  NOR2_X1 U4960 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4687) );
  NOR2_X1 U4961 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4686) );
  INV_X1 U4962 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4635) );
  INV_X1 U4963 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8078) );
  INV_X4 U4964 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U4965 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4946) );
  NOR2_X2 U4966 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5009) );
  OR2_X1 U4967 ( .A1(n5813), .A2(n8114), .ZN(n6098) );
  INV_X1 U4968 ( .A(n5693), .ZN(n5629) );
  AOI22_X1 U4969 ( .A1(n4899), .A2(n4902), .B1(n4900), .B2(n4905), .ZN(n4897)
         );
  NAND2_X2 U4970 ( .A1(n4730), .A2(n6940), .ZN(n5693) );
  XNOR2_X2 U4971 ( .A(n4988), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U4972 ( .A1(n9258), .A2(n4430), .ZN(n9257) );
  AOI21_X2 U4973 ( .B1(n9273), .B2(n9272), .A(n4396), .ZN(n9258) );
  NAND2_X4 U4974 ( .A1(n8444), .A2(n5792), .ZN(n5817) );
  OAI21_X2 U4975 ( .B1(n7289), .B2(n4887), .A(n4885), .ZN(n7367) );
  AOI21_X2 U4976 ( .B1(n7240), .B2(n7504), .A(n4939), .ZN(n7289) );
  NOR2_X2 U4977 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n4304), .ZN(n6075) );
  INV_X2 U4978 ( .A(n5838), .ZN(n5821) );
  BUF_X4 U4979 ( .A(n5813), .Z(n5838) );
  INV_X2 U4980 ( .A(n5836), .ZN(n5819) );
  INV_X2 U4981 ( .A(n5300), .ZN(n4277) );
  INV_X8 U4982 ( .A(n4277), .ZN(n4278) );
  NAND3_X1 U4983 ( .A1(n5019), .A2(n6570), .A3(n5730), .ZN(n5300) );
  XNOR2_X2 U4984 ( .A(n8111), .B(n7950), .ZN(n7795) );
  AOI21_X1 U4985 ( .B1(n4472), .B2(n4679), .A(n4678), .ZN(n8715) );
  NOR2_X1 U4986 ( .A1(n4854), .A2(n4851), .ZN(n4850) );
  INV_X1 U4987 ( .A(n4801), .ZN(n4799) );
  INV_X1 U4988 ( .A(n7532), .ZN(n6226) );
  NAND2_X1 U4989 ( .A1(n7471), .A2(n7470), .ZN(n5937) );
  NAND2_X1 U4990 ( .A1(n7571), .A2(n7675), .ZN(n4543) );
  AND2_X1 U4991 ( .A1(n8677), .A2(n8676), .ZN(n4683) );
  NAND2_X1 U4992 ( .A1(n7678), .A2(n7677), .ZN(n7683) );
  NAND2_X1 U4993 ( .A1(n7669), .A2(n6250), .ZN(n4709) );
  OR2_X1 U4994 ( .A1(n8101), .A2(n7800), .ZN(n7674) );
  AOI21_X1 U4995 ( .B1(n6384), .B2(n9989), .A(n4305), .ZN(n6798) );
  INV_X1 U4996 ( .A(n4870), .ZN(n4869) );
  OAI21_X1 U4997 ( .B1(n5613), .B2(n4871), .A(n5634), .ZN(n4870) );
  INV_X1 U4998 ( .A(n5434), .ZN(n4449) );
  INV_X1 U4999 ( .A(n5381), .ZN(n5367) );
  NOR2_X1 U5000 ( .A1(n4460), .A2(n4874), .ZN(n4459) );
  INV_X1 U5001 ( .A(n4875), .ZN(n4874) );
  INV_X1 U5002 ( .A(n4461), .ZN(n4460) );
  INV_X1 U5003 ( .A(SI_15_), .ZN(n9943) );
  NAND2_X1 U5004 ( .A1(n4574), .A2(n4572), .ZN(n4770) );
  AOI21_X1 U5005 ( .B1(n4575), .B2(n4576), .A(n4361), .ZN(n4574) );
  NAND2_X1 U5006 ( .A1(n6637), .A2(n4573), .ZN(n4572) );
  INV_X1 U5007 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5757) );
  OR2_X1 U5008 ( .A1(n4284), .A2(n6756), .ZN(n4557) );
  NAND2_X1 U5009 ( .A1(n4550), .A2(n4294), .ZN(n4558) );
  INV_X1 U5010 ( .A(n6756), .ZN(n4768) );
  NOR2_X1 U5011 ( .A1(n6766), .A2(n6765), .ZN(n4559) );
  NOR2_X1 U5012 ( .A1(n4917), .A2(n4913), .ZN(n4912) );
  INV_X1 U5013 ( .A(n4919), .ZN(n4913) );
  NAND2_X1 U5014 ( .A1(n4282), .A2(n4325), .ZN(n4921) );
  NAND2_X1 U5015 ( .A1(n6148), .A2(n4282), .ZN(n4922) );
  AND2_X1 U5016 ( .A1(n6142), .A2(n8178), .ZN(n7662) );
  NAND2_X1 U5017 ( .A1(n8226), .A2(n4906), .ZN(n8200) );
  NOR2_X1 U5018 ( .A1(n8218), .A2(n4907), .ZN(n4906) );
  INV_X1 U5019 ( .A(n6134), .ZN(n4907) );
  INV_X1 U5020 ( .A(n5805), .ZN(n5890) );
  INV_X1 U5021 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5022 ( .A1(n5452), .A2(n8584), .ZN(n4504) );
  AOI21_X1 U5023 ( .B1(n8725), .B2(n8726), .A(n4470), .ZN(n8804) );
  OR2_X1 U5024 ( .A1(n9379), .A2(n9118), .ZN(n8761) );
  OR2_X1 U5025 ( .A1(n9344), .A2(n8625), .ZN(n8767) );
  AND4_X1 U5026 ( .A1(n4970), .A2(n4977), .A3(n4971), .A4(n4947), .ZN(n4929)
         );
  NAND2_X1 U5027 ( .A1(n5596), .A2(n5595), .ZN(n5614) );
  NOR2_X1 U5028 ( .A1(n4762), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U5029 ( .A1(n4882), .A2(n5365), .ZN(n5383) );
  NAND2_X1 U5030 ( .A1(n5363), .A2(n5362), .ZN(n4882) );
  OAI211_X1 U5031 ( .C1(n4651), .C2(n4600), .A(n4596), .B(n5198), .ZN(n5226)
         );
  AND2_X1 U5032 ( .A1(n4652), .A2(n4598), .ZN(n4597) );
  INV_X1 U5033 ( .A(n4600), .ZN(n4598) );
  INV_X1 U5034 ( .A(n7521), .ZN(n4990) );
  AND2_X1 U5035 ( .A1(n7868), .A2(n4835), .ZN(n4833) );
  INV_X1 U5036 ( .A(n7904), .ZN(n4841) );
  AND4_X1 U5037 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n7851)
         );
  CLKBUF_X1 U5038 ( .A(n5836), .Z(n7530) );
  AND4_X1 U5039 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n6263)
         );
  NAND2_X1 U5040 ( .A1(n7717), .A2(n5791), .ZN(n5836) );
  AOI21_X1 U5041 ( .B1(n7604), .B2(n4704), .A(n4703), .ZN(n4702) );
  INV_X1 U5042 ( .A(n7609), .ZN(n4703) );
  AOI21_X1 U5043 ( .B1(n7088), .B2(n4693), .A(n4692), .ZN(n4691) );
  INV_X1 U5044 ( .A(n7575), .ZN(n4693) );
  INV_X1 U5045 ( .A(n7589), .ZN(n4692) );
  NOR2_X1 U5046 ( .A1(n9798), .A2(n6259), .ZN(n6292) );
  INV_X1 U5047 ( .A(n9548), .ZN(n9743) );
  NAND2_X1 U5048 ( .A1(n6150), .A2(n6202), .ZN(n9748) );
  NAND2_X1 U5049 ( .A1(n6164), .A2(n6163), .ZN(n6166) );
  INV_X1 U5050 ( .A(n4925), .ZN(n4816) );
  NOR2_X1 U5051 ( .A1(n4732), .A2(n4731), .ZN(n4730) );
  NOR2_X1 U5052 ( .A1(n6571), .A2(n8863), .ZN(n4731) );
  INV_X1 U5053 ( .A(n4796), .ZN(n4795) );
  OAI21_X1 U5054 ( .B1(n4802), .B2(n4797), .A(n4340), .ZN(n4796) );
  NOR2_X1 U5055 ( .A1(n9097), .A2(n4807), .ZN(n4806) );
  INV_X1 U5056 ( .A(n9094), .ZN(n4807) );
  AND2_X1 U5057 ( .A1(n9263), .A2(n9096), .ZN(n9097) );
  NAND2_X1 U5058 ( .A1(n9270), .A2(n9092), .ZN(n9095) );
  OR2_X1 U5059 ( .A1(n9279), .A2(n9091), .ZN(n9092) );
  NAND2_X1 U5060 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  AND2_X1 U5061 ( .A1(n5571), .A2(n5547), .ZN(n5569) );
  OAI21_X1 U5062 ( .B1(n5502), .B2(n9979), .A(n5501), .ZN(n5504) );
  AND2_X1 U5063 ( .A1(n4560), .A2(n4316), .ZN(n7964) );
  NOR2_X1 U5064 ( .A1(n7964), .A2(n7963), .ZN(n7988) );
  AOI21_X1 U5065 ( .B1(n4395), .B2(n4394), .A(n8631), .ZN(n8637) );
  NOR2_X1 U5066 ( .A1(n8633), .A2(n8629), .ZN(n4394) );
  AND2_X1 U5067 ( .A1(n4528), .A2(n4527), .ZN(n4526) );
  AND2_X1 U5068 ( .A1(n7590), .A2(n7675), .ZN(n4529) );
  INV_X1 U5069 ( .A(n4586), .ZN(n4583) );
  OR2_X1 U5070 ( .A1(n4593), .A2(n4589), .ZN(n4584) );
  NAND2_X1 U5071 ( .A1(n4587), .A2(n4588), .ZN(n4585) );
  INV_X1 U5072 ( .A(n8281), .ZN(n4592) );
  NAND2_X1 U5073 ( .A1(n4681), .A2(n9312), .ZN(n8678) );
  NAND2_X1 U5074 ( .A1(n4684), .A2(n4682), .ZN(n4681) );
  AOI21_X1 U5075 ( .B1(n8675), .B2(n8727), .A(n4683), .ZN(n4682) );
  NAND2_X1 U5076 ( .A1(n7639), .A2(n7636), .ZN(n4532) );
  INV_X1 U5077 ( .A(n4669), .ZN(n4668) );
  INV_X1 U5078 ( .A(n8690), .ZN(n4667) );
  MUX2_X1 U5079 ( .A(n9063), .B(n8742), .S(n8722), .Z(n8690) );
  NOR2_X1 U5080 ( .A1(n8733), .A2(n8727), .ZN(n4468) );
  NAND2_X1 U5081 ( .A1(n7647), .A2(n7648), .ZN(n4595) );
  OR2_X1 U5082 ( .A1(n7652), .A2(n7691), .ZN(n4506) );
  INV_X1 U5083 ( .A(n4537), .ZN(n4536) );
  AOI21_X1 U5084 ( .B1(n7665), .B2(n7675), .A(n8144), .ZN(n4537) );
  AOI21_X1 U5085 ( .B1(n4535), .B2(n7664), .A(n7675), .ZN(n4534) );
  OAI21_X1 U5086 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n4535) );
  INV_X1 U5087 ( .A(n7660), .ZN(n7663) );
  AND2_X1 U5088 ( .A1(n8125), .A2(n7668), .ZN(n4533) );
  OR2_X1 U5089 ( .A1(n8738), .A2(n8761), .ZN(n8704) );
  OAI21_X1 U5090 ( .B1(n8721), .B2(n8720), .A(n8724), .ZN(n4471) );
  OR2_X1 U5091 ( .A1(n9246), .A2(n9100), .ZN(n8689) );
  NAND2_X1 U5092 ( .A1(n8632), .A2(n8628), .ZN(n7132) );
  NOR2_X1 U5093 ( .A1(n9300), .A2(n9321), .ZN(n4632) );
  INV_X1 U5094 ( .A(n5615), .ZN(n4871) );
  INV_X1 U5095 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4970) );
  INV_X1 U5096 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4969) );
  INV_X1 U5097 ( .A(n5410), .ZN(n5411) );
  NOR2_X1 U5098 ( .A1(n4463), .A2(n4462), .ZN(n4461) );
  INV_X1 U5099 ( .A(n5227), .ZN(n4462) );
  INV_X1 U5100 ( .A(n5252), .ZN(n4463) );
  AND2_X1 U5101 ( .A1(n6805), .A2(n6258), .ZN(n6262) );
  NAND3_X1 U5102 ( .A1(n6798), .A2(n7559), .A3(n6260), .ZN(n6261) );
  INV_X1 U5103 ( .A(n7734), .ZN(n4834) );
  NOR2_X1 U5104 ( .A1(n4337), .A2(n4296), .ZN(n4513) );
  AND3_X1 U5105 ( .A1(n4383), .A2(n4766), .A3(n4292), .ZN(n6636) );
  NAND2_X1 U5106 ( .A1(n4555), .A2(n4559), .ZN(n4554) );
  INV_X1 U5107 ( .A(n4559), .ZN(n4556) );
  NAND2_X1 U5108 ( .A1(n7385), .A2(n7384), .ZN(n7965) );
  AOI21_X1 U5109 ( .B1(n4707), .B2(n7670), .A(n4339), .ZN(n4706) );
  OAI21_X1 U5110 ( .B1(n4921), .B2(n4281), .A(n4335), .ZN(n4917) );
  AND2_X1 U5111 ( .A1(n4897), .A2(n4350), .ZN(n4895) );
  AOI21_X1 U5112 ( .B1(n4901), .B2(n7507), .A(n7952), .ZN(n4899) );
  AOI21_X1 U5113 ( .B1(n4904), .B2(n7507), .A(n9808), .ZN(n4900) );
  NAND2_X1 U5114 ( .A1(n4336), .A2(n4280), .ZN(n4887) );
  NAND2_X1 U5115 ( .A1(n9737), .A2(n7600), .ZN(n7364) );
  NAND2_X1 U5116 ( .A1(n4317), .A2(n4523), .ZN(n7584) );
  INV_X1 U5117 ( .A(n5840), .ZN(n4524) );
  NOR2_X1 U5119 ( .A1(n6149), .A2(n4920), .ZN(n4919) );
  INV_X1 U5120 ( .A(n6143), .ZN(n4920) );
  OR2_X1 U5121 ( .A1(n8382), .A2(n7847), .ZN(n7664) );
  OR2_X1 U5122 ( .A1(n8422), .A2(n8242), .ZN(n7629) );
  INV_X1 U5123 ( .A(n7333), .ZN(n7704) );
  INV_X1 U5124 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5797) );
  AND2_X1 U5125 ( .A1(n4849), .A2(n5759), .ZN(n4848) );
  INV_X1 U5126 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5760) );
  INV_X1 U5127 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5986) );
  NOR2_X2 U5128 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5803) );
  OR2_X1 U5129 ( .A1(n5225), .A2(n5224), .ZN(n4935) );
  NAND2_X1 U5130 ( .A1(n8810), .A2(n5732), .ZN(n6571) );
  OR2_X1 U5131 ( .A1(n9373), .A2(n9119), .ZN(n8760) );
  OR2_X1 U5132 ( .A1(n9394), .A2(n9110), .ZN(n9065) );
  OR2_X1 U5133 ( .A1(n9231), .A2(n9106), .ZN(n9204) );
  NOR2_X1 U5134 ( .A1(n9279), .A2(n4631), .ZN(n4630) );
  INV_X1 U5135 ( .A(n4632), .ZN(n4631) );
  OR2_X1 U5136 ( .A1(n9442), .A2(n7434), .ZN(n8670) );
  NOR2_X1 U5137 ( .A1(n4431), .A2(n4787), .ZN(n4786) );
  INV_X1 U5138 ( .A(n7256), .ZN(n4789) );
  NAND2_X1 U5139 ( .A1(n4393), .A2(n4323), .ZN(n8812) );
  INV_X1 U5140 ( .A(n7132), .ZN(n4393) );
  NAND2_X1 U5141 ( .A1(n4647), .A2(n4646), .ZN(n8654) );
  AND2_X1 U5142 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5100) );
  NOR2_X1 U5143 ( .A1(n9231), .A2(n9244), .ZN(n9230) );
  NOR2_X1 U5144 ( .A1(n7157), .A2(n9690), .ZN(n7156) );
  OAI21_X1 U5145 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n7520) );
  XNOR2_X1 U5146 ( .A(n7485), .B(n7484), .ZN(n7488) );
  NAND2_X1 U5147 ( .A1(n5676), .A2(n5675), .ZN(n6215) );
  AND2_X1 U5148 ( .A1(n5636), .A2(n5619), .ZN(n5634) );
  AND2_X1 U5149 ( .A1(n5615), .A2(n5600), .ZN(n5613) );
  AND2_X1 U5150 ( .A1(n4969), .A2(n4970), .ZN(n4765) );
  NOR2_X1 U5151 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4764) );
  INV_X1 U5152 ( .A(n4856), .ZN(n5594) );
  OAI21_X1 U5153 ( .B1(n5522), .B2(n4302), .A(n4376), .ZN(n4856) );
  NOR2_X1 U5154 ( .A1(n5542), .A2(n4863), .ZN(n4862) );
  INV_X1 U5155 ( .A(n5521), .ZN(n4863) );
  INV_X1 U5156 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5157 ( .A1(n4444), .A2(n4442), .ZN(n5480) );
  AND2_X1 U5158 ( .A1(n4443), .A2(n5456), .ZN(n4442) );
  NAND2_X1 U5159 ( .A1(n4978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U5160 ( .A1(n4458), .A2(n4872), .ZN(n5336) );
  AOI21_X1 U5161 ( .B1(n4873), .B2(n4875), .A(n4375), .ZN(n4872) );
  NOR2_X1 U5162 ( .A1(n5282), .A2(n4879), .ZN(n4878) );
  INV_X1 U5163 ( .A(n5255), .ZN(n4879) );
  NAND2_X1 U5164 ( .A1(n5228), .A2(n4461), .ZN(n5256) );
  INV_X1 U5165 ( .A(n4850), .ZN(n4655) );
  INV_X1 U5166 ( .A(n5110), .ZN(n4654) );
  INV_X1 U5167 ( .A(n4852), .ZN(n4653) );
  AOI21_X1 U5168 ( .B1(n5146), .B2(n4853), .A(n4345), .ZN(n4852) );
  NAND2_X1 U5169 ( .A1(n5107), .A2(n5106), .ZN(n5111) );
  NAND2_X1 U5170 ( .A1(n4581), .A2(n4993), .ZN(n4995) );
  NAND2_X1 U5171 ( .A1(n4990), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4581) );
  XNOR2_X1 U5172 ( .A(n4995), .B(n4580), .ZN(n4994) );
  INV_X1 U5173 ( .A(SI_1_), .ZN(n4580) );
  OR2_X1 U5174 ( .A1(n7733), .A2(n8215), .ZN(n7734) );
  NAND2_X1 U5175 ( .A1(n7724), .A2(n7952), .ZN(n4842) );
  AOI21_X1 U5176 ( .B1(n4829), .B2(n4828), .A(n4827), .ZN(n4826) );
  INV_X1 U5177 ( .A(n7888), .ZN(n4828) );
  INV_X1 U5178 ( .A(n7746), .ZN(n4827) );
  NAND2_X1 U5179 ( .A1(n7736), .A2(n8229), .ZN(n4835) );
  NAND2_X1 U5180 ( .A1(n4385), .A2(n7473), .ZN(n7721) );
  NAND2_X1 U5181 ( .A1(n7458), .A2(n7457), .ZN(n7722) );
  NAND2_X1 U5182 ( .A1(n4425), .A2(n6817), .ZN(n6819) );
  NAND2_X1 U5183 ( .A1(n7547), .A2(n7559), .ZN(n4414) );
  OR2_X1 U5184 ( .A1(n5836), .A2(n6436), .ZN(n5812) );
  NAND2_X1 U5185 ( .A1(n6488), .A2(n4776), .ZN(n6489) );
  NAND2_X1 U5186 ( .A1(n6476), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5187 ( .A1(n6495), .A2(n6496), .ZN(n6547) );
  AND2_X1 U5188 ( .A1(n6494), .A2(n6493), .ZN(n6495) );
  AND2_X1 U5189 ( .A1(n4355), .A2(n4406), .ZN(n6637) );
  NAND2_X1 U5190 ( .A1(n6636), .A2(n6644), .ZN(n4406) );
  NAND2_X1 U5191 ( .A1(n6637), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9873) );
  INV_X1 U5192 ( .A(n4770), .ZN(n6752) );
  NAND2_X1 U5193 ( .A1(n4550), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4769) );
  AND2_X1 U5194 ( .A1(n5776), .A2(n5757), .ZN(n5928) );
  NOR2_X1 U5195 ( .A1(n7055), .A2(n4338), .ZN(n7057) );
  INV_X1 U5196 ( .A(n4775), .ZN(n7066) );
  NOR2_X1 U5197 ( .A1(n7056), .A2(n7208), .ZN(n4563) );
  NAND2_X1 U5198 ( .A1(n7067), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4774) );
  XOR2_X1 U5199 ( .A(n7965), .B(n7966), .Z(n7386) );
  NOR2_X1 U5200 ( .A1(n7381), .A2(n4561), .ZN(n7959) );
  AND2_X1 U5201 ( .A1(n7383), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4561) );
  AND4_X1 U5202 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n8243)
         );
  NOR2_X1 U5203 ( .A1(n4899), .A2(n4900), .ZN(n4898) );
  CLKBUF_X1 U5204 ( .A(n7368), .Z(n7369) );
  INV_X1 U5205 ( .A(n7470), .ZN(n7501) );
  INV_X1 U5206 ( .A(n7951), .ZN(n9547) );
  AND2_X1 U5207 ( .A1(n7600), .A2(n7596), .ZN(n9732) );
  NAND2_X1 U5208 ( .A1(n7289), .A2(n7581), .ZN(n7288) );
  AND2_X1 U5209 ( .A1(n7582), .A2(n7590), .ZN(n4713) );
  AND2_X1 U5210 ( .A1(n7575), .A2(n7586), .ZN(n7573) );
  OR2_X1 U5211 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  INV_X1 U5212 ( .A(n8122), .ZN(n8125) );
  OR2_X1 U5213 ( .A1(n7549), .A2(n7548), .ZN(n8122) );
  AND2_X1 U5214 ( .A1(n6064), .A2(n7653), .ZN(n4710) );
  OR2_X1 U5215 ( .A1(n8394), .A2(n7767), .ZN(n7653) );
  NAND2_X1 U5216 ( .A1(n8172), .A2(n8176), .ZN(n4711) );
  OR2_X1 U5217 ( .A1(n7662), .A2(n7497), .ZN(n8162) );
  NAND2_X1 U5218 ( .A1(n8200), .A2(n6135), .ZN(n8203) );
  OR2_X1 U5219 ( .A1(n8330), .A2(n7915), .ZN(n8198) );
  NAND2_X1 U5221 ( .A1(n7691), .A2(n6310), .ZN(n9548) );
  INV_X1 U5222 ( .A(n9745), .ZN(n9550) );
  INV_X1 U5223 ( .A(n9748), .ZN(n9546) );
  AND2_X1 U5224 ( .A1(n7691), .A2(n6231), .ZN(n9745) );
  OR2_X1 U5225 ( .A1(n5845), .A2(n5802), .ZN(n5808) );
  OR2_X1 U5226 ( .A1(n5825), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U5227 ( .A(n6191), .B(n6190), .ZN(n7362) );
  NAND2_X1 U5228 ( .A1(n5776), .A2(n4849), .ZN(n5951) );
  INV_X1 U5229 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10007) );
  INV_X1 U5230 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5754) );
  INV_X1 U5231 ( .A(n4483), .ZN(n4482) );
  NAND2_X1 U5232 ( .A1(n4487), .A2(n4485), .ZN(n4484) );
  INV_X1 U5233 ( .A(n4935), .ZN(n4479) );
  INV_X1 U5234 ( .A(n8534), .ZN(n4744) );
  NOR2_X1 U5235 ( .A1(n4744), .A2(n4741), .ZN(n4740) );
  INV_X1 U5236 ( .A(n4748), .ZN(n4741) );
  AND2_X1 U5237 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  OR2_X1 U5238 ( .A1(n5405), .A2(n8518), .ZN(n5408) );
  INV_X1 U5239 ( .A(n5402), .ZN(n4737) );
  NOR2_X1 U5240 ( .A1(n4737), .A2(n4738), .ZN(n4734) );
  INV_X1 U5241 ( .A(n8455), .ZN(n4738) );
  AOI21_X1 U5242 ( .B1(n4748), .B2(n4306), .A(n4746), .ZN(n4745) );
  INV_X1 U5243 ( .A(n5567), .ZN(n4746) );
  XNOR2_X1 U5244 ( .A(n4476), .B(n4278), .ZN(n5096) );
  NAND2_X1 U5245 ( .A1(n5021), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U5246 ( .A1(n8878), .A2(n5661), .ZN(n4477) );
  NAND2_X1 U5247 ( .A1(n4495), .A2(n4493), .ZN(n8544) );
  AOI21_X1 U5248 ( .B1(n4497), .B2(n4500), .A(n4494), .ZN(n4493) );
  INV_X1 U5249 ( .A(n8481), .ZN(n4494) );
  AND2_X1 U5250 ( .A1(n8495), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U5251 ( .A1(n4724), .A2(n8575), .ZN(n4723) );
  INV_X1 U5252 ( .A(n8573), .ZN(n4724) );
  INV_X1 U5253 ( .A(n8575), .ZN(n4725) );
  NAND2_X1 U5254 ( .A1(n4490), .A2(n4489), .ZN(n6961) );
  INV_X1 U5255 ( .A(n4481), .ZN(n4490) );
  NAND2_X1 U5256 ( .A1(n4487), .A2(n6865), .ZN(n4489) );
  OAI21_X1 U5257 ( .B1(n6963), .B2(n4491), .A(n6962), .ZN(n4481) );
  CLKBUF_X1 U5258 ( .A(n8621), .Z(n4420) );
  AND2_X1 U5259 ( .A1(n5275), .A2(n5274), .ZN(n7301) );
  AND2_X2 U5260 ( .A1(n9516), .A2(n4959), .ZN(n6365) );
  NAND2_X1 U5261 ( .A1(n4959), .A2(n4963), .ZN(n5037) );
  NAND2_X2 U5262 ( .A1(n9512), .A2(n9516), .ZN(n8621) );
  AOI21_X1 U5263 ( .B1(n8926), .B2(P1_REG1_REG_5__SCAN_IN), .A(n8919), .ZN(
        n8935) );
  OR2_X1 U5264 ( .A1(n9531), .A2(n9530), .ZN(n6901) );
  NAND2_X1 U5265 ( .A1(n9579), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4390) );
  INV_X1 U5266 ( .A(n4619), .ZN(n4617) );
  NAND2_X1 U5267 ( .A1(n9136), .A2(n4616), .ZN(n4615) );
  NOR2_X1 U5268 ( .A1(n4617), .A2(n8728), .ZN(n4616) );
  NOR2_X1 U5269 ( .A1(n4620), .A2(n9060), .ZN(n4619) );
  INV_X1 U5270 ( .A(n4621), .ZN(n4620) );
  AOI21_X1 U5271 ( .B1(n4795), .B2(n4792), .A(n4791), .ZN(n4790) );
  NOR2_X1 U5272 ( .A1(n9164), .A2(n9116), .ZN(n4791) );
  OR2_X1 U5273 ( .A1(n9180), .A2(n9114), .ZN(n9155) );
  AND2_X1 U5274 ( .A1(n8762), .A2(n9066), .ZN(n9160) );
  NAND2_X1 U5275 ( .A1(n9230), .A2(n4622), .ZN(n9162) );
  AND2_X1 U5276 ( .A1(n9464), .A2(n4285), .ZN(n4622) );
  NAND2_X1 U5277 ( .A1(n9201), .A2(n9110), .ZN(n4801) );
  NOR2_X1 U5278 ( .A1(n4803), .A2(n9112), .ZN(n4802) );
  INV_X1 U5279 ( .A(n4933), .ZN(n4803) );
  AND2_X1 U5280 ( .A1(n9155), .A2(n8763), .ZN(n9178) );
  OR2_X1 U5281 ( .A1(n9342), .A2(n8810), .ZN(n6562) );
  OAI21_X1 U5282 ( .B1(n9219), .B2(n9107), .A(n9211), .ZN(n9109) );
  AND2_X1 U5283 ( .A1(n9065), .A2(n8734), .ZN(n9189) );
  AND2_X1 U5284 ( .A1(n9102), .A2(n4320), .ZN(n4804) );
  OR2_X1 U5285 ( .A1(n9246), .A2(n9261), .ZN(n9244) );
  INV_X1 U5286 ( .A(n8751), .ZN(n4396) );
  NOR2_X1 U5287 ( .A1(n9300), .A2(n9088), .ZN(n9090) );
  OR2_X1 U5288 ( .A1(n9089), .A2(n9491), .ZN(n4931) );
  NAND2_X1 U5289 ( .A1(n9294), .A2(n8749), .ZN(n9273) );
  AOI21_X1 U5290 ( .B1(n4784), .B2(n4318), .A(n4439), .ZN(n9317) );
  NAND2_X1 U5291 ( .A1(n4349), .A2(n4293), .ZN(n4439) );
  NAND2_X1 U5292 ( .A1(n8747), .A2(n8767), .ZN(n9313) );
  AND2_X1 U5293 ( .A1(n4322), .A2(n9079), .ZN(n4783) );
  OR2_X1 U5294 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  AND2_X1 U5295 ( .A1(n8671), .A2(n9329), .ZN(n8789) );
  AOI21_X1 U5296 ( .B1(n8788), .B2(n4643), .A(n4642), .ZN(n4641) );
  INV_X1 U5297 ( .A(n8833), .ZN(n4643) );
  NAND2_X1 U5298 ( .A1(n4640), .A2(n8788), .ZN(n4639) );
  NAND2_X1 U5299 ( .A1(n4424), .A2(n7337), .ZN(n4423) );
  NAND2_X1 U5300 ( .A1(n7335), .A2(n8830), .ZN(n7336) );
  OR2_X1 U5301 ( .A1(n8581), .A2(n7301), .ZN(n7334) );
  OR2_X1 U5302 ( .A1(n7255), .A2(n8874), .ZN(n7256) );
  NAND2_X1 U5303 ( .A1(n7161), .A2(n7143), .ZN(n7144) );
  OR2_X1 U5304 ( .A1(n9690), .A2(n4646), .ZN(n7143) );
  NAND2_X1 U5305 ( .A1(n7144), .A2(n8768), .ZN(n7257) );
  OR2_X2 U5306 ( .A1(n6576), .A2(n8860), .ZN(n9342) );
  INV_X1 U5307 ( .A(n9333), .ZN(n9240) );
  OR2_X1 U5308 ( .A1(n5730), .A2(n8810), .ZN(n6940) );
  NAND2_X1 U5309 ( .A1(n8803), .A2(n8771), .ZN(n6576) );
  NAND2_X1 U5310 ( .A1(n5641), .A2(n5640), .ZN(n9379) );
  INV_X1 U5311 ( .A(n6373), .ZN(n5461) );
  OAI211_X1 U5312 ( .C1(n6343), .C2(n5061), .A(n4611), .B(n4610), .ZN(n4672)
         );
  NAND2_X1 U5313 ( .A1(n6373), .A2(n4288), .ZN(n4611) );
  OR2_X1 U5314 ( .A1(n6373), .A2(n6414), .ZN(n4610) );
  AND2_X1 U5315 ( .A1(n4814), .A2(n4949), .ZN(n4813) );
  INV_X1 U5316 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4951) );
  XNOR2_X1 U5317 ( .A(n7520), .B(n7519), .ZN(n7718) );
  INV_X1 U5318 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U5319 ( .A(n5635), .B(n5634), .ZN(n7480) );
  NAND2_X1 U5320 ( .A1(n4868), .A2(n5615), .ZN(n5635) );
  NAND2_X1 U5321 ( .A1(n5614), .A2(n5613), .ZN(n4868) );
  XNOR2_X1 U5322 ( .A(n5594), .B(n5593), .ZN(n7431) );
  INV_X1 U5323 ( .A(n4862), .ZN(n4466) );
  XNOR2_X1 U5324 ( .A(n5543), .B(n5542), .ZN(n7330) );
  NAND2_X1 U5325 ( .A1(n4864), .A2(n5521), .ZN(n5543) );
  OAI21_X1 U5326 ( .B1(n5480), .B2(n5481), .A(n5482), .ZN(n5502) );
  NAND2_X1 U5327 ( .A1(n4441), .A2(n4445), .ZN(n5457) );
  OR2_X1 U5328 ( .A1(n5383), .A2(n4448), .ZN(n4441) );
  NAND2_X1 U5329 ( .A1(n4450), .A2(n4452), .ZN(n5435) );
  NAND2_X1 U5330 ( .A1(n5383), .A2(n4455), .ZN(n4450) );
  NAND2_X1 U5331 ( .A1(n4451), .A2(n5368), .ZN(n5414) );
  XNOR2_X1 U5332 ( .A(n4604), .B(n5282), .ZN(n6401) );
  NAND2_X1 U5333 ( .A1(n5256), .A2(n5255), .ZN(n4604) );
  NAND2_X1 U5334 ( .A1(n4457), .A2(n4989), .ZN(n5044) );
  NAND2_X1 U5335 ( .A1(n6187), .A2(n6186), .ZN(n6434) );
  INV_X1 U5337 ( .A(n8178), .ZN(n7766) );
  AND4_X1 U5338 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n7424)
         );
  AND3_X1 U5339 ( .A1(n6037), .A2(n6036), .A3(n6035), .ZN(n8211) );
  INV_X1 U5340 ( .A(n8379), .ZN(n7825) );
  AND4_X1 U5341 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n6982)
         );
  OR2_X1 U5342 ( .A1(n7730), .A2(n8242), .ZN(n4386) );
  AND4_X1 U5343 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n6322)
         );
  INV_X1 U5344 ( .A(n7851), .ZN(n8149) );
  INV_X1 U5345 ( .A(n6322), .ZN(n9729) );
  NAND2_X1 U5346 ( .A1(n4405), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4560) );
  INV_X1 U5347 ( .A(n7382), .ZN(n4405) );
  XNOR2_X1 U5348 ( .A(n7959), .B(n7960), .ZN(n7382) );
  NAND2_X1 U5349 ( .A1(n4545), .A2(n4380), .ZN(n4547) );
  OAI22_X1 U5350 ( .A1(n8068), .A2(n8067), .B1(n8072), .B2(n8335), .ZN(n8069)
         );
  XNOR2_X1 U5351 ( .A(n8066), .B(n4381), .ZN(n4409) );
  AOI21_X1 U5352 ( .B1(n6256), .B2(n9748), .A(n6255), .ZN(n8121) );
  NAND2_X1 U5353 ( .A1(n4884), .A2(n6094), .ZN(n8119) );
  INV_X1 U5354 ( .A(n8372), .ZN(n8131) );
  AND2_X1 U5355 ( .A1(n5950), .A2(n7552), .ZN(n4712) );
  INV_X1 U5356 ( .A(n8362), .ZN(n8298) );
  OAI21_X1 U5357 ( .B1(n6802), .B2(n6292), .A(n6804), .ZN(n6197) );
  NAND2_X1 U5358 ( .A1(n6056), .A2(n6055), .ZN(n8388) );
  AND2_X1 U5359 ( .A1(n6434), .A2(n6387), .ZN(n6385) );
  NAND2_X1 U5360 ( .A1(n4496), .A2(n4501), .ZN(n8478) );
  NAND2_X1 U5361 ( .A1(n8526), .A2(n4502), .ZN(n4496) );
  OR2_X1 U5362 ( .A1(n8526), .A2(n4500), .ZN(n4492) );
  OR2_X1 U5363 ( .A1(n8807), .A2(n9040), .ZN(n4676) );
  INV_X1 U5364 ( .A(n7251), .ZN(n8874) );
  INV_X1 U5365 ( .A(n9076), .ZN(n4656) );
  XNOR2_X1 U5366 ( .A(n4658), .B(n9120), .ZN(n4657) );
  OAI211_X1 U5367 ( .C1(n9370), .C2(n9071), .A(n4811), .B(n4808), .ZN(n9365)
         );
  NAND2_X1 U5368 ( .A1(n9120), .A2(n4360), .ZN(n4811) );
  NAND2_X1 U5369 ( .A1(n9135), .A2(n9134), .ZN(n9370) );
  INV_X1 U5370 ( .A(n8814), .ZN(n4613) );
  NAND2_X1 U5371 ( .A1(n4541), .A2(n7573), .ZN(n7588) );
  NAND2_X1 U5372 ( .A1(n7570), .A2(n7691), .ZN(n4542) );
  NAND2_X1 U5373 ( .A1(n8630), .A2(n8822), .ZN(n4395) );
  NAND2_X1 U5374 ( .A1(n4525), .A2(n7610), .ZN(n4588) );
  NAND2_X1 U5375 ( .A1(n7611), .A2(n4526), .ZN(n4525) );
  AND2_X1 U5376 ( .A1(n7612), .A2(n7620), .ZN(n4587) );
  OAI21_X1 U5377 ( .B1(n7616), .B2(n4589), .A(n7619), .ZN(n4586) );
  AND2_X1 U5378 ( .A1(n8264), .A2(n7624), .ZN(n4590) );
  INV_X1 U5379 ( .A(n8678), .ZN(n8683) );
  OAI21_X1 U5380 ( .B1(n8686), .B2(n8722), .A(n8689), .ZN(n4669) );
  OAI22_X1 U5381 ( .A1(n7642), .A2(n4531), .B1(n7643), .B2(n7691), .ZN(n7649)
         );
  AOI22_X1 U5382 ( .A1(n4532), .A2(n4287), .B1(n7644), .B2(n7675), .ZN(n4531)
         );
  NOR2_X1 U5383 ( .A1(n4665), .A2(n4468), .ZN(n4467) );
  NOR2_X1 U5384 ( .A1(n9224), .A2(n4312), .ZN(n4665) );
  NAND2_X1 U5385 ( .A1(n4505), .A2(n4594), .ZN(n7660) );
  INV_X1 U5386 ( .A(n7657), .ZN(n4594) );
  OAI21_X1 U5387 ( .B1(n4536), .B2(n4534), .A(n4533), .ZN(n7672) );
  INV_X1 U5388 ( .A(n8552), .ZN(n4721) );
  NOR2_X1 U5389 ( .A1(n8705), .A2(n8706), .ZN(n4679) );
  NAND2_X1 U5390 ( .A1(n8702), .A2(n8722), .ZN(n8703) );
  AND2_X1 U5391 ( .A1(n8708), .A2(n8722), .ZN(n4678) );
  AND2_X1 U5392 ( .A1(n7135), .A2(n8645), .ZN(n8640) );
  NOR2_X1 U5393 ( .A1(n7687), .A2(n7680), .ZN(n4605) );
  AND2_X1 U5394 ( .A1(n4514), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U5395 ( .A1(n4347), .A2(n7691), .ZN(n4514) );
  NAND2_X1 U5396 ( .A1(n4297), .A2(n7675), .ZN(n4511) );
  NOR2_X1 U5397 ( .A1(n9872), .A2(n7091), .ZN(n4573) );
  INV_X1 U5398 ( .A(n4355), .ZN(n4575) );
  OAI21_X1 U5399 ( .B1(n8552), .B2(n4729), .A(n5333), .ZN(n4728) );
  OR2_X1 U5400 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  AND2_X1 U5401 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  INV_X1 U5402 ( .A(n5086), .ZN(n5136) );
  NAND2_X1 U5403 ( .A1(n8640), .A2(n8654), .ZN(n8781) );
  INV_X1 U5404 ( .A(n4860), .ZN(n4859) );
  OAI21_X1 U5405 ( .B1(n4862), .B2(n4861), .A(n5569), .ZN(n4860) );
  INV_X1 U5406 ( .A(n5571), .ZN(n4857) );
  INV_X1 U5407 ( .A(n5541), .ZN(n4861) );
  NAND2_X1 U5408 ( .A1(n4364), .A2(n5571), .ZN(n4858) );
  INV_X1 U5409 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5436) );
  INV_X1 U5410 ( .A(SI_17_), .ZN(n5415) );
  NOR2_X1 U5411 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4944) );
  NOR2_X1 U5412 ( .A1(n5308), .A2(n4876), .ZN(n4875) );
  INV_X1 U5413 ( .A(n5283), .ZN(n4876) );
  INV_X1 U5414 ( .A(n4878), .ZN(n4873) );
  NAND2_X1 U5415 ( .A1(n4601), .A2(n5172), .ZN(n4600) );
  INV_X1 U5416 ( .A(n5196), .ZN(n4601) );
  INV_X1 U5417 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5173) );
  INV_X1 U5418 ( .A(n5122), .ZN(n4853) );
  INV_X1 U5419 ( .A(n8444), .ZN(n5791) );
  NOR2_X1 U5420 ( .A1(n6518), .A2(n4577), .ZN(n6494) );
  NOR2_X1 U5421 ( .A1(n6530), .A2(n4578), .ZN(n4577) );
  NAND2_X1 U5422 ( .A1(n7078), .A2(n4411), .ZN(n7224) );
  NAND2_X1 U5423 ( .A1(n7067), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5424 ( .A1(n7991), .A2(n7992), .ZN(n8010) );
  AOI21_X1 U5425 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8036), .A(n8035), .ZN(
        n8037) );
  NOR2_X1 U5426 ( .A1(n4705), .A2(n4701), .ZN(n4700) );
  INV_X1 U5427 ( .A(n7600), .ZN(n4701) );
  INV_X1 U5428 ( .A(n7604), .ZN(n4705) );
  NAND2_X1 U5429 ( .A1(n7024), .A2(n5809), .ZN(n7566) );
  OR2_X1 U5430 ( .A1(n7675), .A2(n7697), .ZN(n6297) );
  OR2_X1 U5431 ( .A1(n7825), .A2(n7851), .ZN(n7667) );
  INV_X1 U5432 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U5433 ( .A1(n4925), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5434 ( .A1(n5756), .A2(n4926), .ZN(n4925) );
  INV_X1 U5435 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5436 ( .A1(n4845), .A2(n5766), .ZN(n4844) );
  NAND2_X1 U5437 ( .A1(n4846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4845) );
  AND3_X1 U5438 ( .A1(n10007), .A2(n5927), .A3(n5938), .ZN(n5758) );
  INV_X1 U5439 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5927) );
  BUF_X1 U5440 ( .A(n4990), .Z(n5815) );
  NOR2_X1 U5441 ( .A1(n4488), .A2(n4491), .ZN(n4485) );
  OAI21_X1 U5442 ( .B1(n6962), .B2(n4488), .A(n7031), .ZN(n4483) );
  NAND2_X1 U5443 ( .A1(n4613), .A2(n5086), .ZN(n5029) );
  AOI22_X1 U5444 ( .A1(n4613), .A2(n5689), .B1(n4391), .B2(n5629), .ZN(n5034)
         );
  INV_X1 U5445 ( .A(n6866), .ZN(n4491) );
  INV_X1 U5446 ( .A(n9258), .ZN(n9255) );
  NOR2_X1 U5447 ( .A1(n9604), .A2(n4388), .ZN(n8991) );
  AND2_X1 U5448 ( .A1(n9608), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4388) );
  NOR2_X1 U5449 ( .A1(n9046), .A2(n9373), .ZN(n4621) );
  INV_X1 U5450 ( .A(n9117), .ZN(n4794) );
  NOR2_X1 U5451 ( .A1(n4798), .A2(n9117), .ZN(n4792) );
  NOR2_X1 U5452 ( .A1(n9219), .A2(n9394), .ZN(n4624) );
  OR2_X1 U5453 ( .A1(n5394), .A2(n5374), .ZN(n5423) );
  NOR2_X1 U5454 ( .A1(n8581), .A2(n8502), .ZN(n4628) );
  INV_X1 U5455 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5456 ( .A1(n6784), .A2(n6924), .ZN(n8628) );
  NAND2_X1 U5457 ( .A1(n6587), .A2(n4613), .ZN(n6613) );
  XNOR2_X1 U5458 ( .A(n8815), .B(n4672), .ZN(n8770) );
  NAND2_X1 U5459 ( .A1(n9230), .A2(n9472), .ZN(n9215) );
  NAND2_X1 U5460 ( .A1(n9341), .A2(n4630), .ZN(n9277) );
  AND2_X1 U5461 ( .A1(n7156), .A2(n9569), .ZN(n7260) );
  NOR2_X1 U5462 ( .A1(n6719), .A2(n9656), .ZN(n6722) );
  NAND2_X1 U5463 ( .A1(n4867), .A2(n4865), .ZN(n5674) );
  AOI21_X1 U5464 ( .B1(n4869), .B2(n4871), .A(n4866), .ZN(n4865) );
  INV_X1 U5465 ( .A(n5636), .ZN(n4866) );
  AND2_X1 U5466 ( .A1(n5675), .A2(n5639), .ZN(n5673) );
  AOI21_X1 U5467 ( .B1(n4309), .B2(n4447), .A(n4446), .ZN(n4445) );
  INV_X1 U5468 ( .A(n5433), .ZN(n4446) );
  INV_X1 U5469 ( .A(n4455), .ZN(n4447) );
  INV_X1 U5470 ( .A(n4309), .ZN(n4448) );
  NOR2_X1 U5471 ( .A1(n5413), .A2(n4456), .ZN(n4455) );
  INV_X1 U5472 ( .A(n5368), .ZN(n4456) );
  INV_X1 U5473 ( .A(n4453), .ZN(n4452) );
  OAI21_X1 U5474 ( .B1(n4454), .B2(n5413), .A(n5412), .ZN(n4453) );
  NAND2_X1 U5475 ( .A1(n5366), .A2(n5368), .ZN(n4454) );
  OR2_X1 U5476 ( .A1(n4421), .A2(n6203), .ZN(n6201) );
  OR2_X1 U5477 ( .A1(n4826), .A2(n4825), .ZN(n4823) );
  INV_X1 U5478 ( .A(n7742), .ZN(n4831) );
  INV_X1 U5479 ( .A(n7821), .ZN(n4825) );
  AND2_X1 U5480 ( .A1(n6311), .A2(n6310), .ZN(n7940) );
  AND2_X1 U5481 ( .A1(n7936), .A2(n4315), .ZN(n4820) );
  NAND2_X1 U5482 ( .A1(n7760), .A2(n7759), .ZN(n4821) );
  NAND2_X1 U5483 ( .A1(n5782), .A2(n8065), .ZN(n6258) );
  INV_X1 U5484 ( .A(n7689), .ZN(n7686) );
  OAI21_X1 U5485 ( .B1(n7692), .B2(n7691), .A(n7690), .ZN(n7693) );
  AND4_X1 U5486 ( .A1(n7536), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n7800)
         );
  AND4_X1 U5487 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n7751)
         );
  AND3_X1 U5488 ( .A1(n6046), .A2(n6045), .A3(n6044), .ZN(n7892) );
  NAND2_X1 U5489 ( .A1(n5819), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5490 ( .A1(n5792), .A2(n4890), .ZN(n4889) );
  AND2_X1 U5491 ( .A1(n8444), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4890) );
  XNOR2_X1 U5492 ( .A(n6530), .B(n4578), .ZN(n6520) );
  NOR2_X1 U5493 ( .A1(n6519), .A2(n6520), .ZN(n6518) );
  NAND2_X1 U5494 ( .A1(n6547), .A2(n4544), .ZN(n4766) );
  AND2_X1 U5495 ( .A1(n4767), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5496 ( .A1(n6547), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6548) );
  AOI21_X1 U5497 ( .B1(n9873), .B2(n4355), .A(n9872), .ZN(n9876) );
  NAND2_X1 U5498 ( .A1(n4558), .A2(n4557), .ZN(n6843) );
  OAI211_X1 U5499 ( .C1(n4558), .C2(n6850), .A(n4552), .B(n4551), .ZN(n6845)
         );
  INV_X1 U5500 ( .A(n4553), .ZN(n4552) );
  OAI21_X1 U5501 ( .B1(n4557), .B2(n6850), .A(n4554), .ZN(n4553) );
  NOR2_X1 U5502 ( .A1(n6845), .A2(n6835), .ZN(n7055) );
  XNOR2_X1 U5503 ( .A(n7224), .B(n7208), .ZN(n7080) );
  NAND2_X1 U5504 ( .A1(n4565), .A2(n4568), .ZN(n4775) );
  NAND3_X1 U5505 ( .A1(n4772), .A2(P2_REG2_REG_17__SCAN_IN), .A3(n4571), .ZN(
        n4569) );
  NAND2_X1 U5506 ( .A1(n8037), .A2(n9714), .ZN(n4571) );
  NAND2_X1 U5507 ( .A1(n4570), .A2(n8039), .ZN(n8064) );
  NAND2_X1 U5508 ( .A1(n4569), .A2(n4772), .ZN(n4570) );
  AOI21_X1 U5509 ( .B1(n6237), .B2(n9786), .A(n6234), .ZN(n6235) );
  NOR2_X1 U5510 ( .A1(n4922), .A2(n4281), .ZN(n4918) );
  AND2_X1 U5511 ( .A1(n8126), .A2(n6094), .ZN(n4883) );
  INV_X1 U5512 ( .A(n4922), .ZN(n4916) );
  OR2_X1 U5513 ( .A1(n7670), .A2(n7669), .ZN(n7551) );
  OR2_X1 U5514 ( .A1(n6050), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U5515 ( .A1(n6042), .A2(n6041), .ZN(n6050) );
  AND2_X1 U5516 ( .A1(n6033), .A2(n6032), .ZN(n6042) );
  NAND2_X1 U5517 ( .A1(n6002), .A2(n6001), .ZN(n6014) );
  OR2_X1 U5518 ( .A1(n6014), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6023) );
  INV_X1 U5519 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7831) );
  AND2_X1 U5520 ( .A1(n5989), .A2(n7831), .ZN(n6002) );
  OR2_X1 U5521 ( .A1(n5966), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5977) );
  INV_X1 U5522 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5955) );
  NOR2_X1 U5523 ( .A1(n5944), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5956) );
  NOR2_X1 U5524 ( .A1(n6123), .A2(n9547), .ZN(n4893) );
  INV_X1 U5525 ( .A(n8266), .ZN(n9549) );
  OR2_X1 U5526 ( .A1(n5931), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5944) );
  OR2_X1 U5527 ( .A1(n5921), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5931) );
  OR2_X1 U5528 ( .A1(n7378), .A2(n7424), .ZN(n7579) );
  NAND2_X1 U5529 ( .A1(n7364), .A2(n7506), .ZN(n7419) );
  AOI21_X1 U5530 ( .B1(n7369), .B2(n7421), .A(n7507), .ZN(n7423) );
  INV_X1 U5531 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5911) );
  INV_X1 U5532 ( .A(n4886), .ZN(n4885) );
  OAI21_X1 U5533 ( .B1(n4887), .B2(n7581), .A(n4888), .ZN(n4886) );
  NAND2_X1 U5534 ( .A1(n5905), .A2(n9732), .ZN(n9737) );
  INV_X1 U5535 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6757) );
  AND2_X1 U5536 ( .A1(n5899), .A2(n6757), .ZN(n5912) );
  NOR2_X1 U5537 ( .A1(n5884), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5899) );
  OR2_X1 U5538 ( .A1(n5873), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5884) );
  INV_X1 U5539 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6638) );
  INV_X1 U5540 ( .A(n7957), .ZN(n7103) );
  XNOR2_X1 U5541 ( .A(n7957), .B(n9751), .ZN(n9749) );
  NAND2_X1 U5542 ( .A1(n4688), .A2(n7565), .ZN(n6806) );
  AND2_X1 U5543 ( .A1(n7667), .A2(n7666), .ZN(n8138) );
  NAND2_X1 U5544 ( .A1(n8140), .A2(n9745), .ZN(n4428) );
  INV_X1 U5545 ( .A(n8138), .ZN(n8144) );
  AND2_X1 U5546 ( .A1(n7664), .A2(n7659), .ZN(n8157) );
  AND2_X1 U5547 ( .A1(n4696), .A2(n7643), .ZN(n4695) );
  NAND2_X1 U5548 ( .A1(n4279), .A2(n7635), .ZN(n4696) );
  AND2_X1 U5549 ( .A1(n7645), .A2(n8184), .ZN(n8201) );
  NAND2_X1 U5550 ( .A1(n8226), .A2(n6134), .ZN(n8213) );
  INV_X1 U5551 ( .A(n8225), .ZN(n6133) );
  AND2_X1 U5552 ( .A1(n7637), .A2(n7640), .ZN(n8225) );
  AND4_X1 U5553 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n8254)
         );
  AND4_X1 U5554 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n8253)
         );
  INV_X1 U5555 ( .A(n8251), .ZN(n6130) );
  INV_X1 U5556 ( .A(n8252), .ZN(n6131) );
  AND2_X1 U5557 ( .A1(n7629), .A2(n7630), .ZN(n8251) );
  INV_X1 U5558 ( .A(n9811), .ZN(n9804) );
  OR3_X1 U5559 ( .A1(n6259), .A2(n5782), .A3(n6202), .ZN(n6300) );
  OR2_X1 U5560 ( .A1(n7675), .A2(n6258), .ZN(n6307) );
  OR2_X1 U5561 ( .A1(n6259), .A2(n7704), .ZN(n9793) );
  NAND2_X1 U5562 ( .A1(n4847), .A2(n5779), .ZN(n4846) );
  INV_X1 U5563 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4847) );
  INV_X1 U5564 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5766) );
  AND4_X1 U5565 ( .A1(n5972), .A2(n5761), .A3(n5986), .A4(n5760), .ZN(n5762)
         );
  INV_X1 U5566 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5761) );
  AND2_X1 U5567 ( .A1(n4924), .A2(n4926), .ZN(n5895) );
  NOR2_X1 U5568 ( .A1(n5804), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U5569 ( .A1(n4346), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4777) );
  NOR2_X1 U5570 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4779) );
  NAND2_X1 U5571 ( .A1(n8454), .A2(n8455), .ZN(n8453) );
  AOI21_X1 U5572 ( .B1(n8487), .B2(n8488), .A(n4306), .ZN(n8466) );
  AND2_X1 U5573 ( .A1(n4504), .A2(n8527), .ZN(n4502) );
  NAND2_X1 U5574 ( .A1(n4298), .A2(n4504), .ZN(n4501) );
  AOI21_X1 U5575 ( .B1(n4499), .B2(n4501), .A(n4498), .ZN(n4497) );
  INV_X1 U5576 ( .A(n8479), .ZN(n4498) );
  INV_X1 U5577 ( .A(n4502), .ZN(n4499) );
  INV_X1 U5578 ( .A(n4501), .ZN(n4500) );
  AND2_X1 U5579 ( .A1(n5096), .A2(n4475), .ZN(n5097) );
  INV_X1 U5580 ( .A(n6742), .ZN(n4751) );
  OR2_X1 U5581 ( .A1(n5486), .A2(n8548), .ZN(n5509) );
  NAND2_X1 U5582 ( .A1(n5465), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5486) );
  INV_X1 U5583 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5319) );
  OR2_X1 U5584 ( .A1(n5320), .A2(n5319), .ZN(n5349) );
  OR2_X1 U5585 ( .A1(n5291), .A2(n6920), .ZN(n5320) );
  XNOR2_X1 U5586 ( .A(n8466), .B(n8464), .ZN(n8562) );
  NAND2_X1 U5587 ( .A1(n8572), .A2(n8573), .ZN(n8571) );
  NOR2_X1 U5588 ( .A1(n5423), .A2(n5422), .ZN(n5443) );
  AND2_X1 U5589 ( .A1(n5443), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5465) );
  NOR2_X1 U5590 ( .A1(n5349), .A2(n8458), .ZN(n5392) );
  INV_X1 U5591 ( .A(n5403), .ZN(n8517) );
  NAND2_X1 U5592 ( .A1(n8453), .A2(n5360), .ZN(n8516) );
  AND2_X1 U5593 ( .A1(n8798), .A2(n8727), .ZN(n4469) );
  OR2_X1 U5594 ( .A1(n8728), .A2(n8756), .ZN(n8855) );
  AND3_X1 U5595 ( .A1(n5688), .A2(n5687), .A3(n5686), .ZN(n9119) );
  AND2_X1 U5596 ( .A1(n5244), .A2(n5243), .ZN(n7251) );
  AND2_X1 U5597 ( .A1(n5105), .A2(n5104), .ZN(n6790) );
  INV_X1 U5598 ( .A(n5037), .ZN(n5685) );
  NAND2_X1 U5599 ( .A1(n8895), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4389) );
  AOI21_X1 U5600 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6895), .A(n6894), .ZN(
        n8921) );
  NOR2_X1 U5601 ( .A1(n8933), .A2(n4362), .ZN(n8949) );
  NOR2_X1 U5602 ( .A1(n8949), .A2(n8948), .ZN(n8947) );
  AND2_X1 U5603 ( .A1(n4780), .A2(n4940), .ZN(n4757) );
  AOI21_X1 U5604 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n8954), .A(n8947), .ZN(
        n8963) );
  AOI21_X1 U5605 ( .B1(n8968), .B2(P1_REG1_REG_8__SCAN_IN), .A(n8961), .ZN(
        n8976) );
  NAND2_X1 U5606 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  NAND2_X1 U5607 ( .A1(n8989), .A2(n8990), .ZN(n9590) );
  AOI21_X1 U5608 ( .B1(n9593), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9589), .ZN(
        n9606) );
  XNOR2_X1 U5609 ( .A(n8991), .B(n9002), .ZN(n9622) );
  NAND2_X1 U5610 ( .A1(n8993), .A2(n8994), .ZN(n9011) );
  AND2_X1 U5611 ( .A1(n6372), .A2(n6426), .ZN(n9074) );
  NOR2_X1 U5612 ( .A1(n9120), .A2(n4360), .ZN(n4810) );
  NAND2_X1 U5613 ( .A1(n9230), .A2(n4624), .ZN(n9196) );
  OR2_X1 U5614 ( .A1(n5551), .A2(n5550), .ZN(n5578) );
  NAND2_X1 U5615 ( .A1(n9341), .A2(n4326), .ZN(n9261) );
  AND2_X1 U5616 ( .A1(n8750), .A2(n8751), .ZN(n9272) );
  AND2_X1 U5617 ( .A1(n9290), .A2(n9289), .ZN(n4645) );
  NAND2_X1 U5618 ( .A1(n9341), .A2(n9495), .ZN(n9318) );
  AND2_X1 U5619 ( .A1(n7443), .A2(n9504), .ZN(n9340) );
  AND2_X1 U5620 ( .A1(n9499), .A2(n9340), .ZN(n9341) );
  AND2_X1 U5621 ( .A1(n7260), .A2(n4626), .ZN(n7443) );
  AND2_X1 U5622 ( .A1(n4283), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U5623 ( .A1(n7260), .A2(n4283), .ZN(n7404) );
  AOI21_X1 U5624 ( .B1(n8784), .B2(n4789), .A(n4343), .ZN(n4788) );
  NAND2_X1 U5625 ( .A1(n7260), .A2(n9699), .ZN(n7304) );
  AND2_X1 U5626 ( .A1(n5235), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5266) );
  OR2_X1 U5627 ( .A1(n5183), .A2(n5182), .ZN(n5211) );
  NOR2_X1 U5628 ( .A1(n5211), .A2(n7270), .ZN(n5235) );
  OR2_X1 U5629 ( .A1(n4649), .A2(n7139), .ZN(n7140) );
  AND2_X1 U5630 ( .A1(n6786), .A2(n7167), .ZN(n6942) );
  NAND2_X1 U5631 ( .A1(n4609), .A2(n7118), .ZN(n6658) );
  NOR2_X1 U5632 ( .A1(n6658), .A2(n6870), .ZN(n6786) );
  NAND2_X1 U5633 ( .A1(n8814), .A2(n6599), .ZN(n6719) );
  INV_X1 U5634 ( .A(n9342), .ZN(n9216) );
  INV_X1 U5635 ( .A(n8770), .ZN(n6602) );
  INV_X1 U5636 ( .A(n9051), .ZN(n8588) );
  NAND2_X1 U5637 ( .A1(n4440), .A2(n5527), .ZN(n9231) );
  NAND2_X1 U5638 ( .A1(n7330), .A2(n8716), .ZN(n4440) );
  OR2_X1 U5639 ( .A1(n8722), .A2(n8860), .ZN(n9700) );
  INV_X1 U5640 ( .A(n9698), .ZN(n9443) );
  AND2_X1 U5641 ( .A1(n6568), .A2(n6936), .ZN(n6595) );
  NAND2_X1 U5642 ( .A1(n6574), .A2(n6573), .ZN(n9333) );
  XNOR2_X1 U5643 ( .A(n5674), .B(n5673), .ZN(n8448) );
  XNOR2_X1 U5644 ( .A(n4974), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5710) );
  AND2_X1 U5645 ( .A1(n4765), .A2(n4764), .ZN(n4763) );
  XNOR2_X1 U5646 ( .A(n5717), .B(n5716), .ZN(n6371) );
  NAND2_X1 U5647 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  INV_X1 U5648 ( .A(SI_20_), .ZN(n9979) );
  NAND2_X1 U5649 ( .A1(n4877), .A2(n5283), .ZN(n5309) );
  NAND2_X1 U5650 ( .A1(n5256), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U5651 ( .A1(n5228), .A2(n5227), .ZN(n5251) );
  OAI21_X1 U5652 ( .B1(n5111), .B2(n4655), .A(n4652), .ZN(n5170) );
  NAND2_X1 U5653 ( .A1(n5111), .A2(n5110), .ZN(n5119) );
  INV_X1 U5654 ( .A(n4994), .ZN(n5026) );
  NAND2_X1 U5655 ( .A1(n7908), .A2(n7734), .ZN(n7782) );
  NAND2_X1 U5656 ( .A1(n6269), .A2(n7560), .ZN(n6817) );
  OR2_X1 U5657 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  AND2_X1 U5658 ( .A1(n4842), .A2(n7457), .ZN(n4839) );
  OAI21_X1 U5659 ( .B1(n7760), .B2(n4819), .A(n4817), .ZN(n7830) );
  AOI21_X1 U5660 ( .B1(n4820), .B2(n4818), .A(n4327), .ZN(n4817) );
  INV_X1 U5661 ( .A(n4820), .ZN(n4819) );
  INV_X1 U5662 ( .A(n7759), .ZN(n4818) );
  NAND2_X1 U5663 ( .A1(n7315), .A2(n6327), .ZN(n6330) );
  AND2_X1 U5664 ( .A1(n4832), .A2(n4835), .ZN(n7869) );
  INV_X1 U5665 ( .A(n4840), .ZN(n4837) );
  INV_X1 U5666 ( .A(n7942), .ZN(n7925) );
  AND3_X1 U5667 ( .A1(n6029), .A2(n6028), .A3(n6027), .ZN(n7915) );
  NAND2_X1 U5668 ( .A1(n6977), .A2(n6281), .ZN(n6289) );
  NAND2_X1 U5669 ( .A1(n6293), .A2(n9540), .ZN(n7930) );
  AND4_X1 U5670 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n8242)
         );
  AND2_X1 U5671 ( .A1(n4821), .A2(n4315), .ZN(n7937) );
  NAND2_X1 U5672 ( .A1(n4821), .A2(n4820), .ZN(n7935) );
  INV_X1 U5673 ( .A(n7932), .ZN(n7934) );
  NAND2_X1 U5674 ( .A1(n7700), .A2(n6260), .ZN(n4520) );
  INV_X1 U5675 ( .A(n6258), .ZN(n7697) );
  NAND2_X1 U5676 ( .A1(n7705), .A2(n7706), .ZN(n4518) );
  INV_X1 U5677 ( .A(n7751), .ZN(n8140) );
  NAND2_X1 U5678 ( .A1(n6063), .A2(n6062), .ZN(n8178) );
  INV_X1 U5679 ( .A(n7915), .ZN(n8229) );
  INV_X1 U5680 ( .A(n8243), .ZN(n8215) );
  INV_X1 U5681 ( .A(n8242), .ZN(n8265) );
  INV_X1 U5682 ( .A(n6263), .ZN(n7955) );
  NAND2_X1 U5683 ( .A1(n4311), .A2(n5814), .ZN(n7958) );
  OR2_X1 U5684 ( .A1(P2_U3150), .A2(n6435), .ZN(n9880) );
  INV_X1 U5685 ( .A(n4924), .ZN(n5891) );
  INV_X1 U5686 ( .A(n4769), .ZN(n6753) );
  OAI211_X1 U5687 ( .C1(n4565), .C2(n4567), .A(n4564), .B(n4562), .ZN(n7068)
         );
  AOI21_X1 U5688 ( .B1(n7056), .B2(n4566), .A(n4374), .ZN(n4564) );
  NOR2_X1 U5689 ( .A1(n7068), .A2(n7070), .ZN(n7209) );
  NOR2_X1 U5690 ( .A1(n7213), .A2(n7212), .ZN(n7381) );
  NAND2_X1 U5691 ( .A1(n4771), .A2(n8016), .ZN(n4548) );
  NOR2_X1 U5692 ( .A1(n8007), .A2(n4366), .ZN(n8009) );
  NOR2_X1 U5693 ( .A1(n8006), .A2(n4332), .ZN(n8007) );
  NOR2_X1 U5694 ( .A1(n8009), .A2(n8008), .ZN(n8035) );
  INV_X1 U5695 ( .A(n4569), .ZN(n9722) );
  AND2_X1 U5696 ( .A1(n6444), .A2(n6443), .ZN(n9882) );
  NAND2_X1 U5697 ( .A1(n8034), .A2(n8038), .ZN(n4436) );
  NAND2_X1 U5698 ( .A1(n6221), .A2(n6220), .ZN(n8101) );
  AND2_X1 U5699 ( .A1(n6108), .A2(n6096), .ZN(n8114) );
  NAND2_X1 U5700 ( .A1(n4698), .A2(n7637), .ZN(n8219) );
  NAND2_X1 U5701 ( .A1(n4416), .A2(n7636), .ZN(n4698) );
  OAI21_X1 U5702 ( .B1(n4416), .B2(n7635), .A(n4279), .ZN(n8197) );
  NAND2_X1 U5703 ( .A1(n6022), .A2(n6021), .ZN(n8330) );
  NAND2_X1 U5704 ( .A1(n6000), .A2(n5999), .ZN(n8339) );
  OR2_X1 U5705 ( .A1(n9793), .A2(n9542), .ZN(n8278) );
  NAND2_X1 U5706 ( .A1(n5937), .A2(n7552), .ZN(n8294) );
  NAND2_X1 U5707 ( .A1(n4896), .A2(n4897), .ZN(n8285) );
  OR2_X1 U5708 ( .A1(n7369), .A2(n4898), .ZN(n4896) );
  NAND2_X1 U5709 ( .A1(n4603), .A2(n5930), .ZN(n9808) );
  NAND2_X1 U5710 ( .A1(n6401), .A2(n7525), .ZN(n4603) );
  OR2_X1 U5711 ( .A1(n7368), .A2(n7507), .ZN(n4903) );
  NAND2_X1 U5712 ( .A1(n7288), .A2(n4280), .ZN(n9728) );
  NAND2_X1 U5713 ( .A1(n5883), .A2(n7590), .ZN(n7292) );
  NAND2_X1 U5714 ( .A1(n7104), .A2(n7575), .ZN(n7087) );
  INV_X1 U5715 ( .A(n6956), .ZN(n7024) );
  NAND2_X1 U5716 ( .A1(n6292), .A2(n6385), .ZN(n9540) );
  INV_X1 U5717 ( .A(n8272), .ZN(n9754) );
  OR2_X1 U5718 ( .A1(n6854), .A2(n8278), .ZN(n8095) );
  INV_X1 U5719 ( .A(n9540), .ZN(n9752) );
  AND2_X1 U5720 ( .A1(n4275), .A2(n9811), .ZN(n8350) );
  AND2_X1 U5721 ( .A1(n7528), .A2(n7527), .ZN(n8362) );
  NAND2_X1 U5722 ( .A1(n7494), .A2(n7493), .ZN(n8363) );
  INV_X1 U5723 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n4403) );
  AND2_X1 U5724 ( .A1(n6085), .A2(n6084), .ZN(n8372) );
  NAND2_X1 U5725 ( .A1(n4914), .A2(n6148), .ZN(n8124) );
  AND2_X1 U5726 ( .A1(n6073), .A2(n6072), .ZN(n8379) );
  AOI21_X1 U5727 ( .B1(n4429), .B2(n9748), .A(n4426), .ZN(n8373) );
  NAND2_X1 U5728 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  XNOR2_X1 U5729 ( .A(n8139), .B(n8138), .ZN(n4429) );
  NAND2_X1 U5730 ( .A1(n8164), .A2(n9743), .ZN(n4427) );
  OR2_X1 U5731 ( .A1(n9819), .A2(n9793), .ZN(n8378) );
  NAND2_X1 U5732 ( .A1(n6066), .A2(n6065), .ZN(n8382) );
  NAND2_X1 U5733 ( .A1(n4711), .A2(n7653), .ZN(n8161) );
  NAND2_X1 U5734 ( .A1(n6049), .A2(n6048), .ZN(n8394) );
  NAND2_X1 U5735 ( .A1(n6040), .A2(n6039), .ZN(n8399) );
  NAND2_X1 U5736 ( .A1(n6031), .A2(n6030), .ZN(n8405) );
  NAND2_X1 U5737 ( .A1(n6013), .A2(n6012), .ZN(n8412) );
  NAND2_X1 U5738 ( .A1(n5988), .A2(n5987), .ZN(n8422) );
  NAND2_X1 U5739 ( .A1(n5965), .A2(n5964), .ZN(n8435) );
  INV_X1 U5740 ( .A(n8425), .ZN(n8437) );
  INV_X1 U5741 ( .A(n8378), .ZN(n8436) );
  AND2_X1 U5742 ( .A1(n7362), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6387) );
  NAND2_X1 U5743 ( .A1(n6386), .A2(n6385), .ZN(n6399) );
  OR2_X1 U5744 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  INV_X1 U5745 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10010) );
  INV_X1 U5746 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10005) );
  AND2_X1 U5747 ( .A1(n4412), .A2(P2_U3151), .ZN(n7360) );
  INV_X1 U5748 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7331) );
  XNOR2_X1 U5749 ( .A(n5778), .B(n5777), .ZN(n7333) );
  INV_X1 U5750 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U5751 ( .A1(n5776), .A2(n5775), .ZN(n5784) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7013) );
  INV_X1 U5753 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6830) );
  INV_X1 U5754 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6715) );
  INV_X1 U5755 ( .A(n8033), .ZN(n8036) );
  XNOR2_X1 U5756 ( .A(n5941), .B(n10007), .ZN(n7383) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6403) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6361) );
  INV_X1 U5759 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6350) );
  INV_X1 U5760 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6348) );
  INV_X1 U5761 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6345) );
  INV_X1 U5762 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6339) );
  INV_X1 U5763 ( .A(n6530), .ZN(n6492) );
  AND2_X1 U5764 ( .A1(n6371), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6246) );
  INV_X1 U5765 ( .A(n7134), .ZN(n9684) );
  NAND2_X1 U5766 ( .A1(n6961), .A2(n5145), .ZN(n7030) );
  INV_X1 U5767 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U5768 ( .A1(n4480), .A2(n4478), .ZN(n5248) );
  NAND2_X1 U5769 ( .A1(n4479), .A2(n5246), .ZN(n4478) );
  NAND2_X1 U5770 ( .A1(n7278), .A2(n4314), .ZN(n4480) );
  AND2_X1 U5771 ( .A1(n5663), .A2(n5662), .ZN(n5721) );
  NAND2_X1 U5772 ( .A1(n5508), .A2(n5507), .ZN(n9246) );
  NAND2_X1 U5773 ( .A1(n8571), .A2(n8575), .ZN(n8496) );
  INV_X1 U5774 ( .A(n4743), .ZN(n4742) );
  OAI21_X1 U5775 ( .B1(n4745), .B2(n4744), .A(n5592), .ZN(n4743) );
  NAND2_X1 U5776 ( .A1(n5373), .A2(n5372), .ZN(n9344) );
  OAI21_X1 U5777 ( .B1(n5360), .B2(n4737), .A(n5409), .ZN(n4736) );
  NAND2_X1 U5778 ( .A1(n8533), .A2(n8534), .ZN(n8532) );
  NAND2_X1 U5779 ( .A1(n4747), .A2(n4745), .ZN(n8533) );
  NAND2_X1 U5780 ( .A1(n8487), .A2(n4748), .ZN(n4747) );
  NOR2_X1 U5781 ( .A1(n4373), .A2(n4726), .ZN(n8553) );
  INV_X1 U5782 ( .A(n4729), .ZN(n4726) );
  OR2_X1 U5783 ( .A1(n8572), .A2(n4725), .ZN(n4717) );
  NAND2_X1 U5784 ( .A1(n4716), .A2(n4715), .ZN(n4714) );
  AND2_X1 U5785 ( .A1(n4503), .A2(n5431), .ZN(n8587) );
  NAND2_X1 U5786 ( .A1(n8526), .A2(n8527), .ZN(n4503) );
  NAND2_X1 U5787 ( .A1(n5442), .A2(n5441), .ZN(n9300) );
  INV_X1 U5788 ( .A(n8601), .ZN(n9566) );
  NOR2_X2 U5789 ( .A1(n5723), .A2(n5720), .ZN(n9571) );
  NAND2_X1 U5790 ( .A1(n5390), .A2(n5389), .ZN(n9078) );
  INV_X1 U5791 ( .A(n9568), .ZN(n8613) );
  INV_X1 U5792 ( .A(n9571), .ZN(n8615) );
  INV_X1 U5793 ( .A(n9119), .ZN(n9075) );
  AND2_X1 U5794 ( .A1(n5655), .A2(n5654), .ZN(n9118) );
  OR2_X1 U5795 ( .A1(n5625), .A2(n5624), .ZN(n9116) );
  OR2_X1 U5796 ( .A1(n5396), .A2(n5395), .ZN(n9077) );
  INV_X1 U5797 ( .A(n6790), .ZN(n8877) );
  NAND2_X1 U5798 ( .A1(n8886), .A2(n8885), .ZN(n8884) );
  NAND2_X1 U5799 ( .A1(n8900), .A2(n8901), .ZN(n8899) );
  AOI21_X1 U5800 ( .B1(n8912), .B2(P1_REG1_REG_3__SCAN_IN), .A(n8906), .ZN(
        n6420) );
  INV_X1 U5801 ( .A(n6901), .ZN(n9529) );
  NAND2_X1 U5802 ( .A1(n9011), .A2(n4387), .ZN(n9024) );
  NAND2_X1 U5803 ( .A1(n9004), .A2(n9999), .ZN(n4387) );
  AND2_X1 U5804 ( .A1(n6418), .A2(n6427), .ZN(n9642) );
  NAND2_X1 U5805 ( .A1(n4617), .A2(n8728), .ZN(n4614) );
  NAND2_X1 U5806 ( .A1(n8719), .A2(n8718), .ZN(n9060) );
  OAI21_X1 U5807 ( .B1(n9109), .B2(n4797), .A(n4795), .ZN(n9161) );
  NAND2_X1 U5808 ( .A1(n4800), .A2(n4801), .ZN(n9177) );
  NAND2_X1 U5809 ( .A1(n9109), .A2(n4802), .ZN(n4800) );
  NAND2_X1 U5810 ( .A1(n9109), .A2(n4933), .ZN(n9188) );
  AND2_X1 U5811 ( .A1(n4805), .A2(n4320), .ZN(n9243) );
  NAND2_X1 U5812 ( .A1(n9095), .A2(n9094), .ZN(n9254) );
  INV_X1 U5813 ( .A(n4782), .ZN(n9338) );
  AOI21_X1 U5814 ( .B1(n4784), .B2(n4783), .A(n4308), .ZN(n4782) );
  AND2_X1 U5815 ( .A1(n4784), .A2(n4322), .ZN(n9080) );
  NAND2_X1 U5816 ( .A1(n4639), .A2(n4641), .ZN(n7410) );
  NAND2_X1 U5817 ( .A1(n7336), .A2(n8833), .ZN(n7408) );
  NAND2_X1 U5818 ( .A1(n7258), .A2(n8784), .ZN(n7302) );
  NAND2_X1 U5819 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  INV_X1 U5820 ( .A(n9302), .ZN(n9673) );
  NAND2_X1 U5821 ( .A1(n6388), .A2(n8716), .ZN(n4648) );
  INV_X1 U5822 ( .A(n9657), .ZN(n9345) );
  INV_X1 U5823 ( .A(n9364), .ZN(n4438) );
  OAI21_X1 U5824 ( .B1(n9364), .B2(n4809), .A(n4812), .ZN(n4660) );
  OR2_X1 U5825 ( .A1(n9707), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U5826 ( .A1(n9707), .A2(n9446), .ZN(n4809) );
  INV_X1 U5827 ( .A(n9365), .ZN(n4434) );
  INV_X1 U5828 ( .A(n9231), .ZN(n9476) );
  INV_X1 U5829 ( .A(n9300), .ZN(n9491) );
  INV_X1 U5830 ( .A(n9344), .ZN(n9499) );
  INV_X1 U5831 ( .A(n9078), .ZN(n9504) );
  NAND2_X1 U5832 ( .A1(n5314), .A2(n5313), .ZN(n8558) );
  INV_X1 U5833 ( .A(n9456), .ZN(n9503) );
  NAND2_X2 U5834 ( .A1(n6565), .A2(n6390), .ZN(n9681) );
  OR2_X1 U5835 ( .A1(n4955), .A2(n4954), .ZN(n9507) );
  CLKBUF_X1 U5836 ( .A(n6378), .Z(n9523) );
  XNOR2_X1 U5837 ( .A(n5570), .B(n5569), .ZN(n7361) );
  NAND2_X1 U5838 ( .A1(n4466), .A2(n5541), .ZN(n4465) );
  INV_X1 U5839 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9936) );
  INV_X1 U5840 ( .A(n8863), .ZN(n8803) );
  NAND2_X1 U5841 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4980) );
  INV_X1 U5842 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10019) );
  INV_X1 U5843 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6829) );
  INV_X1 U5844 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6687) );
  INV_X1 U5845 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9920) );
  INV_X1 U5846 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6352) );
  INV_X1 U5847 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6347) );
  INV_X1 U5848 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6344) );
  INV_X1 U5849 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9992) );
  XNOR2_X1 U5850 ( .A(n5028), .B(n5027), .ZN(n6414) );
  NAND2_X1 U5851 ( .A1(n4457), .A2(SI_0_), .ZN(n5043) );
  INV_X2 U5852 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9045) );
  INV_X1 U5853 ( .A(n4560), .ZN(n7961) );
  INV_X1 U5854 ( .A(n8084), .ZN(n4407) );
  OAI21_X1 U5855 ( .B1(n8304), .B2(n9833), .A(n4399), .ZN(n8305) );
  NAND2_X1 U5856 ( .A1(n9833), .A2(n4400), .ZN(n4399) );
  INV_X1 U5857 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5858 ( .A1(n4404), .A2(n4401), .ZN(P2_U3454) );
  NOR2_X1 U5859 ( .A1(n6257), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U5860 ( .A1(n8304), .A2(n9817), .ZN(n4404) );
  NOR2_X1 U5861 ( .A1(n9817), .A2(n4403), .ZN(n4402) );
  AOI21_X1 U5862 ( .B1(n9367), .B2(n4613), .A(n4612), .ZN(n6653) );
  NOR2_X1 U5863 ( .A1(n9712), .A2(n6413), .ZN(n4612) );
  AND2_X1 U5864 ( .A1(n8218), .A2(n4290), .ZN(n4279) );
  OR2_X1 U5865 ( .A1(n9729), .A2(n7195), .ZN(n4280) );
  NAND2_X1 U5866 ( .A1(n8711), .A2(n8710), .ZN(n9046) );
  INV_X1 U5867 ( .A(n5431), .ZN(n5432) );
  AND2_X1 U5868 ( .A1(n8119), .A2(n8126), .ZN(n4281) );
  INV_X1 U5869 ( .A(n8784), .ZN(n4431) );
  OR2_X1 U5870 ( .A1(n8372), .A2(n7751), .ZN(n4282) );
  AND2_X1 U5871 ( .A1(n4628), .A2(n7344), .ZN(n4283) );
  OR2_X1 U5872 ( .A1(n6752), .A2(n6747), .ZN(n4284) );
  AND2_X1 U5873 ( .A1(n4624), .A2(n4623), .ZN(n4285) );
  AND2_X1 U5874 ( .A1(n4772), .A2(n4571), .ZN(n4286) );
  AND2_X1 U5875 ( .A1(n8218), .A2(n7637), .ZN(n4287) );
  AND2_X1 U5876 ( .A1(n4412), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4288) );
  NAND2_X1 U5877 ( .A1(n4884), .A2(n4883), .ZN(n6250) );
  AND2_X1 U5878 ( .A1(n7579), .A2(n7597), .ZN(n7506) );
  INV_X1 U5879 ( .A(n7506), .ZN(n4704) );
  INV_X1 U5880 ( .A(n7118), .ZN(n6660) );
  AND2_X1 U5881 ( .A1(n7540), .A2(n7539), .ZN(n4289) );
  OR2_X1 U5882 ( .A1(n7636), .A2(n7635), .ZN(n4290) );
  AND2_X1 U5883 ( .A1(n8762), .A2(n8727), .ZN(n4291) );
  NAND2_X1 U5884 ( .A1(n6635), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4292) );
  INV_X1 U5885 ( .A(n7153), .ZN(n4649) );
  INV_X1 U5886 ( .A(n9110), .ZN(n9111) );
  AND2_X1 U5887 ( .A1(n5587), .A2(n5586), .ZN(n9110) );
  NAND2_X1 U5888 ( .A1(n9344), .A2(n9082), .ZN(n4293) );
  AND2_X1 U5889 ( .A1(n4768), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4294) );
  AND2_X1 U5890 ( .A1(n4334), .A2(n4780), .ZN(n4295) );
  NOR2_X1 U5891 ( .A1(n4289), .A2(n7691), .ZN(n4296) );
  AND2_X1 U5892 ( .A1(n7683), .A2(n6233), .ZN(n4297) );
  OR2_X1 U5893 ( .A1(n5432), .A2(n4365), .ZN(n4298) );
  AND2_X1 U5894 ( .A1(n4445), .A2(n5453), .ZN(n4299) );
  AND2_X1 U5895 ( .A1(n4641), .A2(n4644), .ZN(n4300) );
  AND2_X1 U5896 ( .A1(n4823), .A2(n4371), .ZN(n4301) );
  INV_X1 U5898 ( .A(n7620), .ZN(n4589) );
  INV_X1 U5899 ( .A(n7056), .ZN(n4568) );
  AND2_X1 U5900 ( .A1(n5217), .A2(n5216), .ZN(n7142) );
  INV_X1 U5901 ( .A(n7142), .ZN(n4646) );
  NAND2_X1 U5902 ( .A1(n7721), .A2(n7722), .ZN(n7903) );
  AND2_X1 U5903 ( .A1(n5297), .A2(n5296), .ZN(n7337) );
  OR2_X1 U5904 ( .A1(n4858), .A2(n4861), .ZN(n4302) );
  INV_X1 U5905 ( .A(n7208), .ZN(n4773) );
  INV_X1 U5906 ( .A(n7079), .ZN(n7067) );
  NAND2_X1 U5907 ( .A1(n7260), .A2(n4628), .ZN(n4629) );
  AND2_X1 U5908 ( .A1(n4548), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4303) );
  OR2_X1 U5909 ( .A1(n6057), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4304) );
  NAND2_X2 U5910 ( .A1(n5019), .A2(n5020), .ZN(n5047) );
  NAND2_X1 U5911 ( .A1(n8620), .A2(n8619), .ZN(n8728) );
  AND2_X1 U5912 ( .A1(n7483), .A2(n7452), .ZN(n4305) );
  INV_X1 U5913 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U5914 ( .A1(n5519), .A2(n5518), .ZN(n4306) );
  OAI211_X1 U5915 ( .C1(n6443), .C2(n6561), .A(n5847), .B(n5846), .ZN(n9751)
         );
  INV_X1 U5916 ( .A(n9751), .ZN(n4522) );
  NAND2_X1 U5917 ( .A1(n5707), .A2(n4975), .ZN(n5019) );
  AND2_X1 U5918 ( .A1(n9136), .A2(n9047), .ZN(n4307) );
  NOR2_X1 U5919 ( .A1(n9504), .A2(n9081), .ZN(n4308) );
  INV_X1 U5920 ( .A(n9872), .ZN(n4576) );
  AND2_X1 U5921 ( .A1(n4452), .A2(n4449), .ZN(n4309) );
  INV_X1 U5922 ( .A(n5095), .ZN(n4475) );
  OR2_X1 U5923 ( .A1(n6843), .A2(n4559), .ZN(n4310) );
  AND3_X1 U5924 ( .A1(n5812), .A2(n5811), .A3(n5810), .ZN(n4311) );
  OR3_X1 U5925 ( .A1(n9101), .A2(n8727), .A3(n9099), .ZN(n4312) );
  INV_X1 U5926 ( .A(n4830), .ZN(n4829) );
  OR2_X1 U5927 ( .A1(n7747), .A2(n4831), .ZN(n4830) );
  INV_X1 U5928 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4957) );
  INV_X1 U5929 ( .A(n8832), .ZN(n4642) );
  XOR2_X1 U5930 ( .A(n5116), .B(n4278), .Z(n4313) );
  NAND2_X1 U5931 ( .A1(n5602), .A2(n5601), .ZN(n9180) );
  INV_X1 U5932 ( .A(n9180), .ZN(n4623) );
  AND2_X1 U5933 ( .A1(n5222), .A2(n5246), .ZN(n4314) );
  INV_X1 U5934 ( .A(n7088), .ZN(n4694) );
  NAND2_X1 U5935 ( .A1(n7727), .A2(n9549), .ZN(n4315) );
  OR2_X1 U5936 ( .A1(n7960), .A2(n7959), .ZN(n4316) );
  AND3_X1 U5937 ( .A1(n5841), .A2(n5839), .A3(n4521), .ZN(n4317) );
  AND2_X1 U5938 ( .A1(n9337), .A2(n4783), .ZN(n4318) );
  AND2_X1 U5939 ( .A1(n4909), .A2(n4908), .ZN(n4319) );
  NAND2_X1 U5940 ( .A1(n9483), .A2(n9098), .ZN(n4320) );
  AND2_X1 U5941 ( .A1(n8899), .A2(n4389), .ZN(n4321) );
  OR2_X1 U5942 ( .A1(n9442), .A2(n8870), .ZN(n4322) );
  NAND2_X1 U5943 ( .A1(n5485), .A2(n5484), .ZN(n9263) );
  NAND2_X1 U5944 ( .A1(n5834), .A2(n7569), .ZN(n5832) );
  AND2_X1 U5945 ( .A1(n7131), .A2(n8655), .ZN(n4323) );
  OR2_X1 U5946 ( .A1(n8105), .A2(n9798), .ZN(n4324) );
  INV_X1 U5947 ( .A(n9219), .ZN(n9472) );
  NAND2_X1 U5948 ( .A1(n5549), .A2(n5548), .ZN(n9219) );
  AND2_X1 U5949 ( .A1(n8372), .A2(n7751), .ZN(n4325) );
  AND2_X1 U5950 ( .A1(n4630), .A2(n9483), .ZN(n4326) );
  AND2_X1 U5951 ( .A1(n7728), .A2(n7729), .ZN(n4327) );
  AND2_X1 U5952 ( .A1(n9212), .A2(n9204), .ZN(n4328) );
  AND2_X1 U5953 ( .A1(n9576), .A2(n4390), .ZN(n4329) );
  AND2_X1 U5954 ( .A1(n4492), .A2(n4497), .ZN(n4330) );
  INV_X1 U5955 ( .A(n9321), .ZN(n9495) );
  NAND2_X1 U5956 ( .A1(n5421), .A2(n5420), .ZN(n9321) );
  INV_X1 U5957 ( .A(n9279), .ZN(n9487) );
  NAND2_X1 U5958 ( .A1(n5464), .A2(n5463), .ZN(n9279) );
  AND4_X1 U5959 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n6233)
         );
  AND2_X1 U5960 ( .A1(n9189), .A2(n9190), .ZN(n4331) );
  INV_X1 U5961 ( .A(n6498), .ZN(n4767) );
  NAND2_X1 U5962 ( .A1(n5679), .A2(n5678), .ZN(n9373) );
  INV_X1 U5963 ( .A(n6211), .ZN(n8111) );
  AND2_X1 U5964 ( .A1(n6104), .A2(n6103), .ZN(n6211) );
  NOR2_X1 U5965 ( .A1(n7988), .A2(n4771), .ZN(n4332) );
  NAND2_X1 U5966 ( .A1(n9230), .A2(n4285), .ZN(n4625) );
  NAND2_X1 U5967 ( .A1(n4904), .A2(n9808), .ZN(n4902) );
  OR2_X1 U5968 ( .A1(n7696), .A2(n7694), .ZN(n4333) );
  OR2_X1 U5969 ( .A1(n8412), .A2(n8243), .ZN(n7637) );
  INV_X1 U5970 ( .A(n4798), .ZN(n4797) );
  NOR2_X1 U5971 ( .A1(n9115), .A2(n4799), .ZN(n4798) );
  AND3_X1 U5972 ( .A1(n4940), .A2(n4947), .A3(n4945), .ZN(n4334) );
  OR2_X1 U5973 ( .A1(n8119), .A2(n8126), .ZN(n4335) );
  OR2_X1 U5974 ( .A1(n9738), .A2(n7954), .ZN(n4336) );
  NOR2_X1 U5975 ( .A1(n4605), .A2(n7675), .ZN(n4337) );
  AND2_X1 U5976 ( .A1(n4310), .A2(n4555), .ZN(n4338) );
  NOR2_X1 U5977 ( .A1(n8111), .A2(n6233), .ZN(n4339) );
  OR2_X1 U5978 ( .A1(n9114), .A2(n4623), .ZN(n4340) );
  OR2_X1 U5979 ( .A1(n9802), .A2(n7953), .ZN(n4341) );
  OR2_X1 U5980 ( .A1(n5370), .A2(n4948), .ZN(n4342) );
  XNOR2_X1 U5981 ( .A(n6215), .B(n6214), .ZN(n6101) );
  NOR2_X1 U5982 ( .A1(n8581), .A2(n8873), .ZN(n4343) );
  INV_X1 U5983 ( .A(n5809), .ZN(n6264) );
  OR2_X1 U5984 ( .A1(n7686), .A2(n7685), .ZN(n4344) );
  AND4_X1 U5985 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n8287)
         );
  INV_X1 U5986 ( .A(n8287), .ZN(n7952) );
  AND2_X1 U5987 ( .A1(n8752), .A2(n8754), .ZN(n9120) );
  AND2_X1 U5988 ( .A1(n5149), .A2(SI_6_), .ZN(n4345) );
  INV_X1 U5989 ( .A(n9201), .ZN(n9394) );
  AND2_X1 U5990 ( .A1(n5577), .A2(n5576), .ZN(n9201) );
  AND2_X1 U5991 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4346) );
  AND2_X1 U5992 ( .A1(n7683), .A2(n6211), .ZN(n4347) );
  AND2_X1 U5993 ( .A1(n9136), .A2(n4619), .ZN(n4348) );
  INV_X1 U5994 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U5995 ( .A1(n9337), .A2(n4308), .ZN(n4349) );
  OR2_X1 U5996 ( .A1(n9815), .A2(n7951), .ZN(n4350) );
  OR2_X1 U5997 ( .A1(n9744), .A2(n5830), .ZN(n4351) );
  OR2_X1 U5998 ( .A1(n8875), .A2(n7134), .ZN(n4352) );
  AND2_X1 U5999 ( .A1(n7592), .A2(n7691), .ZN(n4353) );
  INV_X1 U6000 ( .A(n5145), .ZN(n4488) );
  OR2_X1 U6001 ( .A1(n4918), .A2(n4917), .ZN(n4354) );
  OR2_X1 U6002 ( .A1(n6636), .A2(n6644), .ZN(n4355) );
  NAND2_X1 U6003 ( .A1(n5621), .A2(n5620), .ZN(n9164) );
  AND2_X1 U6004 ( .A1(n6287), .A2(n6281), .ZN(n4356) );
  AND2_X1 U6005 ( .A1(n4795), .A2(n4794), .ZN(n4357) );
  AND2_X1 U6006 ( .A1(n6328), .A2(n6327), .ZN(n4358) );
  AND2_X1 U6007 ( .A1(n4775), .A2(n4774), .ZN(n4359) );
  OR2_X1 U6008 ( .A1(n8399), .A2(n7892), .ZN(n7650) );
  INV_X1 U6009 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5789) );
  INV_X1 U6010 ( .A(n4772), .ZN(n8040) );
  OR2_X1 U6011 ( .A1(n8037), .A2(n9714), .ZN(n4772) );
  INV_X1 U6012 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5759) );
  INV_X1 U6013 ( .A(n4708), .ZN(n4707) );
  INV_X1 U6014 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4947) );
  INV_X1 U6015 ( .A(n8728), .ZN(n9451) );
  INV_X1 U6016 ( .A(n7409), .ZN(n4644) );
  INV_X1 U6017 ( .A(n6850), .ZN(n4555) );
  NOR2_X1 U6018 ( .A1(n9119), .A2(n9047), .ZN(n4360) );
  AND2_X1 U6019 ( .A1(n9871), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4361) );
  INV_X1 U6020 ( .A(n8768), .ZN(n4787) );
  AND2_X1 U6021 ( .A1(n8940), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U6022 ( .A1(n6128), .A2(n6127), .ZN(n8263) );
  INV_X1 U6023 ( .A(n6766), .ZN(n6844) );
  AND2_X1 U6024 ( .A1(n4903), .A2(n4904), .ZN(n4363) );
  OR2_X1 U6025 ( .A1(n5520), .A2(SI_21_), .ZN(n4364) );
  AND2_X1 U6026 ( .A1(n8585), .A2(n5451), .ZN(n4365) );
  INV_X1 U6027 ( .A(n9256), .ZN(n4430) );
  NOR2_X1 U6028 ( .A1(n5150), .A2(n4762), .ZN(n5384) );
  AND3_X1 U6029 ( .A1(n4547), .A2(n4303), .A3(n4546), .ZN(n4366) );
  OR2_X1 U6030 ( .A1(n6211), .A2(n8313), .ZN(n4367) );
  AND2_X1 U6031 ( .A1(n4556), .A2(n6850), .ZN(n4368) );
  NAND2_X1 U6032 ( .A1(n9341), .A2(n4632), .ZN(n4633) );
  AND2_X1 U6033 ( .A1(n8339), .A2(n8228), .ZN(n4369) );
  OR2_X1 U6034 ( .A1(n6211), .A2(n8378), .ZN(n4370) );
  NAND2_X1 U6035 ( .A1(n7749), .A2(n7851), .ZN(n4371) );
  AND2_X1 U6036 ( .A1(n8198), .A2(n7644), .ZN(n8218) );
  AND2_X1 U6037 ( .A1(n4837), .A2(n7722), .ZN(n4372) );
  AND2_X1 U6038 ( .A1(n4717), .A2(n4722), .ZN(n4373) );
  NOR2_X1 U6039 ( .A1(n4774), .A2(n7208), .ZN(n4374) );
  AND2_X1 U6040 ( .A1(n5307), .A2(SI_12_), .ZN(n4375) );
  OR2_X1 U6041 ( .A1(n4859), .A2(n4857), .ZN(n4376) );
  INV_X1 U6042 ( .A(n4567), .ZN(n4566) );
  NAND2_X1 U6043 ( .A1(n4774), .A2(n7208), .ZN(n4567) );
  NOR2_X1 U6044 ( .A1(n7783), .A2(n4834), .ZN(n4377) );
  INV_X1 U6045 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4926) );
  AND2_X2 U6046 ( .A1(n6595), .A2(n6594), .ZN(n9712) );
  NAND2_X1 U6047 ( .A1(n8803), .A2(n9040), .ZN(n8722) );
  NAND2_X1 U6048 ( .A1(n5346), .A2(n5345), .ZN(n9442) );
  INV_X1 U6049 ( .A(n9442), .ZN(n4627) );
  NOR2_X1 U6050 ( .A1(n6865), .A2(n6866), .ZN(n6864) );
  XNOR2_X1 U6051 ( .A(n4770), .B(n6754), .ZN(n6694) );
  INV_X1 U6052 ( .A(n6694), .ZN(n4550) );
  NAND2_X1 U6053 ( .A1(n6259), .A2(n7704), .ZN(n7675) );
  NAND2_X1 U6054 ( .A1(n4750), .A2(n4751), .ZN(n4755) );
  INV_X2 U6055 ( .A(n9819), .ZN(n9817) );
  AND2_X1 U6056 ( .A1(n6207), .A2(n6206), .ZN(n9819) );
  AND2_X1 U6057 ( .A1(n6854), .A2(n9540), .ZN(n9757) );
  INV_X1 U6058 ( .A(n9757), .ZN(n8268) );
  NAND2_X1 U6059 ( .A1(n5179), .A2(n5178), .ZN(n7139) );
  INV_X1 U6060 ( .A(n7139), .ZN(n4650) );
  NAND2_X1 U6061 ( .A1(n6723), .A2(n9700), .ZN(n9695) );
  INV_X1 U6062 ( .A(n9695), .ZN(n9446) );
  AND3_X1 U6063 ( .A1(n5036), .A2(n5052), .A3(n5051), .ZN(n6459) );
  AND2_X2 U6064 ( .A1(n6595), .A2(n6938), .ZN(n9707) );
  NAND2_X1 U6065 ( .A1(n6197), .A2(n6196), .ZN(n9833) );
  NAND2_X1 U6066 ( .A1(n5287), .A2(n5286), .ZN(n8502) );
  INV_X1 U6067 ( .A(n8502), .ZN(n4424) );
  INV_X1 U6068 ( .A(n7975), .ZN(n7990) );
  NAND2_X1 U6069 ( .A1(n4648), .A2(n5207), .ZN(n9690) );
  INV_X1 U6070 ( .A(n9690), .ZN(n4647) );
  NAND2_X1 U6071 ( .A1(n6722), .A2(n8819), .ZN(n6611) );
  INV_X1 U6072 ( .A(n6611), .ZN(n4609) );
  OR2_X1 U6073 ( .A1(n9817), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4378) );
  AND2_X1 U6074 ( .A1(n4769), .A2(n4284), .ZN(n4379) );
  AND2_X1 U6075 ( .A1(n4549), .A2(n8006), .ZN(n4380) );
  INV_X1 U6076 ( .A(n4771), .ZN(n4549) );
  NOR2_X1 U6077 ( .A1(n7975), .A2(n7974), .ZN(n4771) );
  INV_X1 U6078 ( .A(n8065), .ZN(n8080) );
  XOR2_X1 U6079 ( .A(n8065), .B(P2_REG2_REG_19__SCAN_IN), .Z(n4381) );
  AND2_X1 U6080 ( .A1(n4383), .A2(n4766), .ZN(n4382) );
  OR2_X1 U6081 ( .A1(n6497), .A2(n6498), .ZN(n4383) );
  INV_X1 U6082 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n4397) );
  INV_X1 U6083 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U6084 ( .A1(n6977), .A2(n4356), .ZN(n6320) );
  OAI21_X2 U6085 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7908) );
  NAND2_X1 U6086 ( .A1(n5785), .A2(n4909), .ZN(n6167) );
  OAI21_X1 U6087 ( .B1(n7738), .B2(n8191), .A(n7867), .ZN(n7805) );
  NAND2_X1 U6088 ( .A1(n4384), .A2(n4838), .ZN(n7813) );
  AND3_X2 U6089 ( .A1(n5827), .A2(n5829), .A3(n5828), .ZN(n6807) );
  NAND2_X1 U6090 ( .A1(n5801), .A2(n5800), .ZN(n4689) );
  INV_X1 U6091 ( .A(n7720), .ZN(n4385) );
  NAND2_X2 U6092 ( .A1(n6325), .A2(n7312), .ZN(n7315) );
  NAND2_X1 U6093 ( .A1(n4840), .A2(n4842), .ZN(n4384) );
  NAND2_X1 U6094 ( .A1(n7858), .A2(n7857), .ZN(n6972) );
  NAND2_X1 U6095 ( .A1(n7830), .A2(n7829), .ZN(n7828) );
  NAND2_X1 U6096 ( .A1(n7828), .A2(n4386), .ZN(n7837) );
  NAND2_X1 U6097 ( .A1(n7775), .A2(n7774), .ZN(n7773) );
  XNOR2_X1 U6098 ( .A(n6807), .B(n7750), .ZN(n6271) );
  NAND2_X1 U6099 ( .A1(n4689), .A2(n4690), .ZN(n6156) );
  NOR2_X1 U6100 ( .A1(n7837), .A2(n7838), .ZN(n7911) );
  NAND2_X1 U6101 ( .A1(n7721), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U6102 ( .A1(n6188), .A2(n6190), .ZN(n6160) );
  XNOR2_X1 U6103 ( .A(n6956), .B(n6267), .ZN(n6265) );
  NAND2_X1 U6104 ( .A1(n6819), .A2(n6270), .ZN(n6672) );
  OR2_X2 U6105 ( .A1(n6241), .A2(n9819), .ZN(n6239) );
  NAND2_X1 U6106 ( .A1(n7238), .A2(n7239), .ZN(n5883) );
  NAND2_X1 U6107 ( .A1(n5785), .A2(n4930), .ZN(n6168) );
  NAND2_X1 U6108 ( .A1(n5785), .A2(n4539), .ZN(n5788) );
  NAND2_X1 U6109 ( .A1(n6009), .A2(n6008), .ZN(n8236) );
  OAI21_X1 U6110 ( .B1(n8262), .B2(n5983), .A(n7625), .ZN(n8250) );
  NAND3_X2 U6111 ( .A1(n5823), .A2(n5822), .A3(n5824), .ZN(n9744) );
  NOR2_X1 U6112 ( .A1(n9590), .A2(n9591), .ZN(n9589) );
  NAND2_X1 U6113 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U6114 ( .A1(n6584), .A2(n8772), .ZN(n6608) );
  NAND2_X1 U6115 ( .A1(n7303), .A2(n8786), .ZN(n7342) );
  NAND2_X1 U6116 ( .A1(n6785), .A2(n6789), .ZN(n6926) );
  AOI22_X1 U6117 ( .A1(n9143), .A2(n9144), .B1(n9152), .B2(n9118), .ZN(n9135)
         );
  AOI21_X1 U6118 ( .B1(n9476), .B2(n9106), .A(n9105), .ZN(n9211) );
  NAND2_X1 U6119 ( .A1(n4670), .A2(n4392), .ZN(n8815) );
  AND2_X1 U6120 ( .A1(n5023), .A2(n5024), .ZN(n4392) );
  NAND2_X1 U6121 ( .A1(n6602), .A2(n6598), .ZN(n6597) );
  NAND2_X1 U6122 ( .A1(n7403), .A2(n7402), .ZN(n7436) );
  NAND3_X1 U6123 ( .A1(n4422), .A2(n9712), .A3(n4438), .ZN(n4417) );
  NAND2_X1 U6124 ( .A1(n7343), .A2(n7407), .ZN(n7403) );
  XNOR2_X2 U6125 ( .A(n4958), .B(n4957), .ZN(n4963) );
  INV_X1 U6126 ( .A(n4660), .ZN(n4659) );
  INV_X1 U6127 ( .A(n4905), .ZN(n4904) );
  NAND2_X1 U6128 ( .A1(n8163), .A2(n6141), .ZN(n6144) );
  INV_X1 U6129 ( .A(n4902), .ZN(n4901) );
  INV_X1 U6130 ( .A(n5118), .ZN(n4851) );
  INV_X1 U6131 ( .A(n5146), .ZN(n4854) );
  NAND2_X1 U6132 ( .A1(n8227), .A2(n6133), .ZN(n8226) );
  NAND2_X1 U6133 ( .A1(n4911), .A2(n4354), .ZN(n6213) );
  NAND2_X1 U6134 ( .A1(n4894), .A2(n4892), .ZN(n9544) );
  INV_X2 U6135 ( .A(n6160), .ZN(n5785) );
  NAND2_X1 U6136 ( .A1(n4471), .A2(n8852), .ZN(n4470) );
  NAND2_X1 U6137 ( .A1(n4664), .A2(n4467), .ZN(n8692) );
  AOI21_X1 U6138 ( .B1(n4674), .B2(n8860), .A(n8859), .ZN(n8867) );
  NOR2_X1 U6139 ( .A1(n8804), .A2(n4469), .ZN(n8809) );
  NAND2_X1 U6140 ( .A1(n8674), .A2(n8722), .ZN(n4684) );
  NAND2_X1 U6141 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  NAND2_X2 U6142 ( .A1(n9227), .A2(n4328), .ZN(n9207) );
  OR2_X1 U6143 ( .A1(n5037), .A2(n4397), .ZN(n5024) );
  NAND2_X1 U6144 ( .A1(n4699), .A2(n4702), .ZN(n7471) );
  OAI22_X2 U6145 ( .A1(n9742), .A2(n6118), .B1(n7103), .B2(n4522), .ZN(n7100)
         );
  NOR2_X2 U6146 ( .A1(n7099), .A2(n6119), .ZN(n7089) );
  NAND2_X1 U6147 ( .A1(n7368), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U6148 ( .A1(n4915), .A2(n4921), .ZN(n6252) );
  AND2_X2 U6149 ( .A1(n5785), .A2(n4319), .ZN(n5796) );
  NAND2_X1 U6150 ( .A1(n5890), .A2(n6545), .ZN(n5807) );
  NAND2_X1 U6151 ( .A1(n4914), .A2(n4916), .ZN(n4915) );
  INV_X1 U6152 ( .A(n7057), .ZN(n4565) );
  NAND2_X1 U6153 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  AOI21_X1 U6154 ( .B1(n9104), .B2(n9231), .A(n9223), .ZN(n9105) );
  NAND3_X1 U6155 ( .A1(n4410), .A2(n4408), .A3(n4407), .ZN(P2_U3201) );
  NAND2_X1 U6156 ( .A1(n4409), .A2(n9874), .ZN(n4408) );
  NAND2_X1 U6157 ( .A1(n8085), .A2(n9720), .ZN(n4410) );
  NAND2_X1 U6158 ( .A1(n7080), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7225) );
  AOI22_X2 U6159 ( .A1(n6546), .A2(P2_REG1_REG_3__SCAN_IN), .B1(n6483), .B2(
        n6561), .ZN(n6484) );
  XNOR2_X1 U6160 ( .A(n6482), .B(n6561), .ZN(n6546) );
  NAND2_X1 U6161 ( .A1(n6832), .A2(n6833), .ZN(n7050) );
  NAND2_X1 U6162 ( .A1(n9716), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U6163 ( .A1(n4602), .A2(n4651), .ZN(n4599) );
  OR2_X2 U6164 ( .A1(n8781), .A2(n8631), .ZN(n7136) );
  NAND2_X2 U6165 ( .A1(n5937), .A2(n4712), .ZN(n9812) );
  XNOR2_X1 U6166 ( .A(n4413), .B(n8080), .ZN(n7700) );
  NAND2_X1 U6167 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  NAND2_X1 U6168 ( .A1(n7546), .A2(n6259), .ZN(n4415) );
  NAND2_X1 U6169 ( .A1(n4520), .A2(n7705), .ZN(n4519) );
  NAND2_X1 U6170 ( .A1(n4417), .A2(n4437), .ZN(n9369) );
  NAND2_X1 U6171 ( .A1(n6657), .A2(n8774), .ZN(n6783) );
  NAND2_X1 U6172 ( .A1(n6927), .A2(n8642), .ZN(n6994) );
  NAND2_X1 U6173 ( .A1(n6716), .A2(n6724), .ZN(n6718) );
  AND3_X2 U6174 ( .A1(n5808), .A2(n5807), .A3(n5806), .ZN(n6956) );
  OR2_X1 U6175 ( .A1(n9712), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U6176 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  OAI21_X2 U6179 ( .B1(n9287), .B2(n9090), .A(n4931), .ZN(n9270) );
  NAND2_X1 U6180 ( .A1(n6994), .A2(n4352), .ZN(n6995) );
  NAND2_X1 U6181 ( .A1(n7342), .A2(n4423), .ZN(n7343) );
  NAND2_X1 U6182 ( .A1(n9365), .A2(n9695), .ZN(n4422) );
  NAND2_X1 U6183 ( .A1(n7189), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U6184 ( .A1(n4785), .A2(n4788), .ZN(n7303) );
  NAND2_X1 U6185 ( .A1(n4836), .A2(n4833), .ZN(n7867) );
  NAND2_X1 U6186 ( .A1(n7887), .A2(n7742), .ZN(n7844) );
  XNOR2_X1 U6187 ( .A(n7844), .B(n7845), .ZN(n7846) );
  AOI22_X2 U6188 ( .A1(n7805), .A2(n7806), .B1(n7892), .B2(n7739), .ZN(n7889)
         );
  NAND2_X1 U6189 ( .A1(n6609), .A2(n8775), .ZN(n6656) );
  INV_X1 U6190 ( .A(n6818), .ZN(n4425) );
  NAND2_X1 U6191 ( .A1(n6266), .A2(n6270), .ZN(n6818) );
  AOI21_X2 U6192 ( .B1(n6171), .B2(n7479), .A(n7483), .ZN(n6384) );
  INV_X1 U6193 ( .A(n5796), .ZN(n4690) );
  NAND2_X1 U6194 ( .A1(n8745), .A2(n8789), .ZN(n9330) );
  NAND2_X1 U6195 ( .A1(n4659), .A2(n4433), .ZN(n9458) );
  NAND2_X1 U6196 ( .A1(n9130), .A2(n9131), .ZN(n9129) );
  OAI21_X2 U6197 ( .B1(n7248), .B2(n8768), .A(n8658), .ZN(n7249) );
  OAI21_X2 U6198 ( .B1(n9238), .B2(n9064), .A(n9063), .ZN(n9225) );
  NAND2_X2 U6199 ( .A1(n4432), .A2(n4431), .ZN(n7335) );
  INV_X1 U6200 ( .A(n7249), .ZN(n4432) );
  AND2_X2 U6201 ( .A1(n7437), .A2(n8670), .ZN(n8745) );
  NAND2_X1 U6202 ( .A1(n8011), .A2(n8012), .ZN(n8013) );
  NAND2_X1 U6203 ( .A1(n6751), .A2(n6750), .ZN(n6832) );
  NAND2_X1 U6204 ( .A1(n9317), .A2(n9084), .ZN(n9087) );
  NAND4_X2 U6205 ( .A1(n5074), .A2(n5075), .A3(n5076), .A4(n5073), .ZN(n8879)
         );
  NAND2_X1 U6206 ( .A1(n4639), .A2(n4300), .ZN(n7437) );
  NAND2_X1 U6207 ( .A1(n9129), .A2(n9070), .ZN(n4658) );
  NAND2_X1 U6208 ( .A1(n4793), .A2(n4790), .ZN(n9143) );
  NAND2_X1 U6209 ( .A1(n4815), .A2(n4813), .ZN(n4955) );
  NOR2_X1 U6210 ( .A1(n9620), .A2(n8992), .ZN(n8993) );
  NAND2_X1 U6211 ( .A1(n4519), .A2(n4518), .ZN(n4516) );
  NAND2_X1 U6212 ( .A1(n9812), .A2(n7554), .ZN(n9537) );
  NAND2_X1 U6213 ( .A1(n4697), .A2(n4695), .ZN(n8185) );
  NAND2_X1 U6214 ( .A1(n8250), .A2(n7630), .ZN(n5996) );
  NAND2_X1 U6215 ( .A1(n5383), .A2(n4299), .ZN(n4444) );
  OR2_X1 U6216 ( .A1(n5383), .A2(n5366), .ZN(n4451) );
  NAND3_X1 U6217 ( .A1(n4445), .A2(n4448), .A3(n5453), .ZN(n4443) );
  MUX2_X1 U6218 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n4990), .Z(n5364) );
  MUX2_X1 U6219 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n5815), .Z(n5381) );
  MUX2_X1 U6220 ( .A(n6687), .B(n6715), .S(n4412), .Z(n5410) );
  MUX2_X1 U6221 ( .A(n6829), .B(n6830), .S(n4412), .Z(n5416) );
  MUX2_X1 U6222 ( .A(n6950), .B(n5436), .S(n4412), .Z(n5454) );
  MUX2_X1 U6223 ( .A(n10019), .B(n7013), .S(n4412), .Z(n5458) );
  MUX2_X1 U6224 ( .A(n9936), .B(n7331), .S(n4412), .Z(n5524) );
  MUX2_X1 U6225 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n4412), .Z(n5520) );
  MUX2_X1 U6226 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n4412), .Z(n5500) );
  MUX2_X1 U6227 ( .A(n10025), .B(n10005), .S(n4412), .Z(n5545) );
  MUX2_X1 U6228 ( .A(n7468), .B(n7477), .S(n4412), .Z(n5598) );
  MUX2_X1 U6229 ( .A(n7432), .B(n10010), .S(n4412), .Z(n5573) );
  MUX2_X1 U6230 ( .A(n9998), .B(n10024), .S(n4412), .Z(n5617) );
  MUX2_X1 U6231 ( .A(n9519), .B(n5677), .S(n4412), .Z(n6217) );
  MUX2_X1 U6232 ( .A(n9956), .B(n9982), .S(n4412), .Z(n7484) );
  NAND2_X1 U6233 ( .A1(n5228), .A2(n4459), .ZN(n4458) );
  AND2_X1 U6234 ( .A1(n4464), .A2(n4465), .ZN(n5570) );
  NAND4_X1 U6235 ( .A1(n5504), .A2(n5503), .A3(n5541), .A4(n4364), .ZN(n4464)
         );
  NAND2_X1 U6236 ( .A1(n5504), .A2(n5503), .ZN(n5522) );
  NAND3_X1 U6237 ( .A1(n5504), .A2(n5503), .A3(n4364), .ZN(n4864) );
  NAND3_X1 U6238 ( .A1(n4473), .A2(n4680), .A3(n8707), .ZN(n4472) );
  OAI21_X1 U6239 ( .B1(n8698), .B2(n8735), .A(n4291), .ZN(n4473) );
  NAND2_X2 U6240 ( .A1(n9560), .A2(n5250), .ZN(n8572) );
  NAND2_X1 U6241 ( .A1(n7265), .A2(n4935), .ZN(n5247) );
  INV_X1 U6242 ( .A(n6963), .ZN(n4487) );
  NAND3_X1 U6243 ( .A1(n4486), .A2(n4484), .A3(n4482), .ZN(n7029) );
  NAND3_X1 U6244 ( .A1(n4487), .A2(n6865), .A3(n5145), .ZN(n4486) );
  NAND2_X1 U6245 ( .A1(n8526), .A2(n4497), .ZN(n4495) );
  NAND3_X1 U6246 ( .A1(n4507), .A2(n8176), .A3(n4506), .ZN(n4505) );
  NAND2_X1 U6247 ( .A1(n4508), .A2(n7691), .ZN(n4507) );
  NAND2_X1 U6248 ( .A1(n4595), .A2(n7650), .ZN(n4508) );
  NAND3_X1 U6249 ( .A1(n4880), .A2(n4518), .A3(n4333), .ZN(n4517) );
  NAND3_X1 U6250 ( .A1(n4517), .A2(n4516), .A3(n4515), .ZN(P2_U3296) );
  NAND3_X1 U6251 ( .A1(n7699), .A2(n4518), .A3(n7697), .ZN(n4515) );
  NOR2_X1 U6252 ( .A1(n4524), .A2(n4522), .ZN(n4523) );
  NAND3_X1 U6253 ( .A1(n7594), .A2(n7593), .A3(n4353), .ZN(n4527) );
  NAND3_X1 U6254 ( .A1(n7583), .A2(n7593), .A3(n4529), .ZN(n4528) );
  NAND2_X1 U6255 ( .A1(n4538), .A2(n5785), .ZN(n4540) );
  NAND3_X1 U6256 ( .A1(n4543), .A2(n7572), .A3(n4542), .ZN(n4541) );
  NAND2_X1 U6257 ( .A1(n7988), .A2(n8016), .ZN(n4546) );
  INV_X1 U6258 ( .A(n7988), .ZN(n4545) );
  NAND3_X1 U6259 ( .A1(n4547), .A2(n4548), .A3(n4546), .ZN(n7989) );
  NAND3_X1 U6260 ( .A1(n4557), .A2(n4368), .A3(n4558), .ZN(n4551) );
  NAND2_X1 U6261 ( .A1(n4565), .A2(n4563), .ZN(n4562) );
  INV_X2 U6262 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4579) );
  NAND2_X1 U6263 ( .A1(n4582), .A2(n4592), .ZN(n4591) );
  NAND3_X1 U6264 ( .A1(n4585), .A2(n4584), .A3(n4583), .ZN(n4582) );
  NAND2_X1 U6265 ( .A1(n4591), .A2(n4590), .ZN(n7628) );
  OR2_X1 U6266 ( .A1(n7612), .A2(n7613), .ZN(n4593) );
  NAND2_X1 U6267 ( .A1(n4597), .A2(n5111), .ZN(n4596) );
  NAND2_X1 U6268 ( .A1(n5111), .A2(n4652), .ZN(n4602) );
  NAND3_X1 U6269 ( .A1(n4606), .A2(n4295), .A3(n4759), .ZN(n4976) );
  INV_X1 U6270 ( .A(n4762), .ZN(n4606) );
  NAND2_X1 U6271 ( .A1(n4758), .A2(n4607), .ZN(n4762) );
  AND2_X1 U6272 ( .A1(n4942), .A2(n4941), .ZN(n4607) );
  INV_X1 U6273 ( .A(n4815), .ZN(n5370) );
  NAND2_X1 U6274 ( .A1(n4815), .A2(n4814), .ZN(n4608) );
  AND2_X2 U6275 ( .A1(n4761), .A2(n4760), .ZN(n4815) );
  NAND2_X4 U6276 ( .A1(n6378), .A2(n9520), .ZN(n6373) );
  XNOR2_X2 U6277 ( .A(n5005), .B(n5004), .ZN(n9520) );
  XNOR2_X2 U6278 ( .A(n5008), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6378) );
  NAND2_X2 U6279 ( .A1(n6373), .A2(n4412), .ZN(n8717) );
  OR2_X1 U6280 ( .A1(n9136), .A2(n9451), .ZN(n4618) );
  NAND2_X1 U6281 ( .A1(n9136), .A2(n4621), .ZN(n9123) );
  NAND3_X1 U6282 ( .A1(n4618), .A2(n4615), .A3(n4614), .ZN(n9048) );
  INV_X1 U6283 ( .A(n4625), .ZN(n9179) );
  INV_X1 U6284 ( .A(n4629), .ZN(n7345) );
  INV_X1 U6285 ( .A(n4633), .ZN(n9299) );
  NAND2_X4 U6286 ( .A1(n4636), .A2(n4634), .ZN(n7521) );
  NAND3_X1 U6287 ( .A1(n4635), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U6288 ( .A1(n5077), .A2(n5078), .ZN(n4637) );
  NAND2_X1 U6289 ( .A1(n5059), .A2(n5060), .ZN(n4638) );
  INV_X1 U6290 ( .A(n7336), .ZN(n4640) );
  NAND2_X2 U6291 ( .A1(n9313), .A2(n9312), .ZN(n9311) );
  NAND2_X2 U6292 ( .A1(n4650), .A2(n4649), .ZN(n8645) );
  AOI21_X2 U6293 ( .B1(n4850), .B2(n4654), .A(n4653), .ZN(n4652) );
  OR2_X2 U6294 ( .A1(n9225), .A2(n9224), .ZN(n9227) );
  NAND2_X2 U6295 ( .A1(n9257), .A2(n9062), .ZN(n9238) );
  NAND2_X1 U6296 ( .A1(n4666), .A2(n4661), .ZN(n4664) );
  NAND3_X1 U6297 ( .A1(n4663), .A2(n4668), .A3(n4662), .ZN(n4661) );
  OR2_X1 U6298 ( .A1(n8684), .A2(n8727), .ZN(n4662) );
  NOR2_X1 U6299 ( .A1(n4667), .A2(n9224), .ZN(n4666) );
  OAI22_X1 U6300 ( .A1(n5740), .A2(n6413), .B1(n8621), .B2(n5022), .ZN(n4671)
         );
  INV_X1 U6301 ( .A(n4671), .ZN(n4670) );
  OAI21_X2 U6302 ( .B1(n8630), .B2(n8629), .A(n8822), .ZN(n8632) );
  NAND2_X1 U6303 ( .A1(n6659), .A2(n8821), .ZN(n4673) );
  NAND3_X1 U6304 ( .A1(n4677), .A2(n4676), .A3(n4675), .ZN(n4674) );
  NAND3_X1 U6305 ( .A1(n8806), .A2(n9040), .A3(n8805), .ZN(n4675) );
  NAND3_X1 U6306 ( .A1(n8701), .A2(n8722), .A3(n9066), .ZN(n4680) );
  NAND2_X1 U6307 ( .A1(n4685), .A2(n9749), .ZN(n5848) );
  XNOR2_X1 U6308 ( .A(n4685), .B(n9749), .ZN(n9764) );
  NAND2_X1 U6309 ( .A1(n5835), .A2(n5834), .ZN(n4685) );
  NAND3_X1 U6310 ( .A1(n5803), .A2(n4687), .A3(n4686), .ZN(n5879) );
  NAND2_X1 U6311 ( .A1(n4688), .A2(n6955), .ZN(n7026) );
  OR2_X1 U6312 ( .A1(n6115), .A2(n7560), .ZN(n4688) );
  NAND2_X2 U6313 ( .A1(n6156), .A2(n6155), .ZN(n5805) );
  OAI21_X2 U6314 ( .B1(n7104), .B2(n4694), .A(n4691), .ZN(n7238) );
  NAND2_X1 U6315 ( .A1(n8236), .A2(n4279), .ZN(n4697) );
  NAND2_X1 U6316 ( .A1(n9737), .A2(n4700), .ZN(n4699) );
  OAI21_X1 U6317 ( .B1(n6251), .B2(n7669), .A(n6250), .ZN(n6224) );
  NAND2_X1 U6318 ( .A1(n7795), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U6319 ( .A1(n4711), .A2(n4710), .ZN(n8156) );
  NAND2_X1 U6320 ( .A1(n5883), .A2(n4713), .ZN(n9735) );
  NAND2_X1 U6321 ( .A1(n9735), .A2(n9734), .ZN(n5905) );
  NAND2_X1 U6322 ( .A1(n6083), .A2(n7667), .ZN(n8123) );
  OAI21_X1 U6323 ( .B1(n7545), .B2(n7544), .A(n7543), .ZN(n7546) );
  NAND2_X2 U6324 ( .A1(n7566), .A2(n7565), .ZN(n6115) );
  NAND2_X1 U6325 ( .A1(n6071), .A2(n7664), .ZN(n8145) );
  NAND2_X1 U6326 ( .A1(n5962), .A2(n7618), .ZN(n8282) );
  AOI211_X1 U6327 ( .C1(n8669), .C2(n8668), .A(n8667), .B(n4642), .ZN(n8673)
         );
  OAI21_X1 U6328 ( .B1(n8695), .B2(n8694), .A(n8693), .ZN(n8700) );
  INV_X1 U6329 ( .A(n5150), .ZN(n4761) );
  NAND2_X1 U6330 ( .A1(n5119), .A2(n5118), .ZN(n4855) );
  NAND2_X1 U6331 ( .A1(n4855), .A2(n5122), .ZN(n5147) );
  NAND2_X1 U6332 ( .A1(n8648), .A2(n8647), .ZN(n8657) );
  AOI21_X1 U6333 ( .B1(n8660), .B2(n8826), .A(n8829), .ZN(n8662) );
  XNOR2_X2 U6334 ( .A(n8879), .B(n8819), .ZN(n8772) );
  NAND2_X1 U6335 ( .A1(n6047), .A2(n7650), .ZN(n8172) );
  INV_X2 U6336 ( .A(n7717), .ZN(n5792) );
  OAI21_X2 U6337 ( .B1(n6459), .B2(n6461), .A(n6460), .ZN(n6458) );
  INV_X1 U6338 ( .A(n5051), .ZN(n6506) );
  NAND2_X1 U6339 ( .A1(n5036), .A2(n5052), .ZN(n6505) );
  NAND2_X1 U6340 ( .A1(n6458), .A2(n5070), .ZN(n6680) );
  AND2_X1 U6341 ( .A1(n5070), .A2(n4714), .ZN(n6460) );
  INV_X1 U6342 ( .A(n5068), .ZN(n4715) );
  INV_X1 U6343 ( .A(n5069), .ZN(n4716) );
  NAND3_X1 U6344 ( .A1(n4722), .A2(n4721), .A3(n4725), .ZN(n4719) );
  INV_X1 U6345 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U6346 ( .A1(n5304), .A2(n5303), .ZN(n4729) );
  NAND2_X2 U6347 ( .A1(n4278), .A2(n4273), .ZN(n5086) );
  NAND2_X1 U6348 ( .A1(n8454), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6349 ( .A1(n8487), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U6350 ( .A1(n4739), .A2(n4742), .ZN(n8506) );
  NOR2_X1 U6351 ( .A1(n5568), .A2(n4749), .ZN(n4748) );
  NOR2_X1 U6352 ( .A1(n8488), .A2(n4306), .ZN(n4749) );
  NAND2_X1 U6353 ( .A1(n4755), .A2(n4753), .ZN(n4756) );
  INV_X1 U6354 ( .A(n6741), .ZN(n4750) );
  INV_X1 U6355 ( .A(n4755), .ZN(n6740) );
  NAND2_X1 U6356 ( .A1(n4755), .A2(n4754), .ZN(n5117) );
  NAND2_X1 U6357 ( .A1(n4756), .A2(n4313), .ZN(n4752) );
  INV_X1 U6358 ( .A(n5097), .ZN(n4753) );
  NOR2_X1 U6359 ( .A1(n5097), .A2(n4313), .ZN(n4754) );
  AND2_X2 U6360 ( .A1(n5010), .A2(n5009), .ZN(n4759) );
  NAND2_X2 U6361 ( .A1(n4759), .A2(n4757), .ZN(n5150) );
  NAND2_X1 U6362 ( .A1(n4981), .A2(n4765), .ZN(n4986) );
  NAND2_X1 U6363 ( .A1(n4981), .A2(n4763), .ZN(n4972) );
  AND2_X1 U6364 ( .A1(n4981), .A2(n4969), .ZN(n4987) );
  NAND3_X1 U6365 ( .A1(n5010), .A2(n5009), .A3(n4780), .ZN(n5123) );
  INV_X2 U6366 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U6367 ( .A1(n7436), .A2(n7435), .ZN(n4784) );
  NAND2_X1 U6368 ( .A1(n7144), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U6369 ( .A1(n9109), .A2(n4357), .ZN(n4793) );
  NAND2_X1 U6370 ( .A1(n4805), .A2(n4804), .ZN(n9103) );
  NAND2_X1 U6371 ( .A1(n9095), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U6372 ( .A1(n9370), .A2(n4810), .ZN(n4808) );
  NOR2_X2 U6373 ( .A1(n4948), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4814) );
  AND2_X2 U6374 ( .A1(n5755), .A2(n5754), .ZN(n4924) );
  NAND2_X1 U6375 ( .A1(n7889), .A2(n7888), .ZN(n7887) );
  OAI21_X1 U6376 ( .B1(n7889), .B2(n4830), .A(n4826), .ZN(n7820) );
  INV_X1 U6377 ( .A(n4822), .ZN(n7920) );
  OAI21_X1 U6378 ( .B1(n7889), .B2(n4824), .A(n4301), .ZN(n4822) );
  NAND2_X1 U6379 ( .A1(n7908), .A2(n4377), .ZN(n4836) );
  CLKBUF_X1 U6380 ( .A(n4836), .Z(n4832) );
  INV_X1 U6381 ( .A(n4832), .ZN(n7781) );
  NAND2_X1 U6382 ( .A1(n7458), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U6383 ( .A1(n7315), .A2(n4358), .ZN(n7456) );
  OAI21_X1 U6384 ( .B1(n6010), .B2(n4846), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5767) );
  INV_X1 U6385 ( .A(n4843), .ZN(n5764) );
  NAND2_X1 U6386 ( .A1(n5776), .A2(n4848), .ZN(n5963) );
  NAND2_X1 U6387 ( .A1(n5614), .A2(n4869), .ZN(n4867) );
  AOI21_X1 U6388 ( .B1(n7693), .B2(n7695), .A(n7698), .ZN(n4880) );
  INV_X1 U6389 ( .A(n7693), .ZN(n4881) );
  AOI21_X1 U6390 ( .B1(n7696), .B2(n4881), .A(n7694), .ZN(n7699) );
  INV_X1 U6391 ( .A(n6250), .ZN(n7670) );
  NAND2_X1 U6392 ( .A1(n8448), .A2(n7525), .ZN(n4884) );
  INV_X1 U6393 ( .A(n7367), .ZN(n6122) );
  OR2_X1 U6394 ( .A1(n7371), .A2(n9789), .ZN(n4888) );
  NAND3_X1 U6395 ( .A1(n5795), .A2(n5793), .A3(n4891), .ZN(n5809) );
  AND2_X1 U6396 ( .A1(n5794), .A2(n4889), .ZN(n4891) );
  OAI21_X2 U6397 ( .B1(n7507), .B2(n7421), .A(n4341), .ZN(n4905) );
  NAND2_X1 U6398 ( .A1(n6144), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U6399 ( .A1(n6144), .A2(n4919), .ZN(n4914) );
  NAND2_X1 U6400 ( .A1(n6144), .A2(n6143), .ZN(n8148) );
  OAI21_X2 U6401 ( .B1(n8263), .B2(n8264), .A(n6129), .ZN(n8252) );
  NAND2_X1 U6402 ( .A1(n4976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6403 ( .A1(n4986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5714) );
  OR2_X1 U6404 ( .A1(n4987), .A2(n5386), .ZN(n4988) );
  INV_X1 U6405 ( .A(n9287), .ZN(n9288) );
  INV_X1 U6406 ( .A(n9373), .ZN(n9047) );
  CLKBUF_X1 U6407 ( .A(n9270), .Z(n9271) );
  NAND2_X1 U6408 ( .A1(n5357), .A2(n5359), .ZN(n5360) );
  XNOR2_X1 U6409 ( .A(n7488), .B(SI_29_), .ZN(n8709) );
  AND2_X1 U6410 ( .A1(n7521), .A2(P2_U3151), .ZN(n8446) );
  NAND2_X1 U6411 ( .A1(n7521), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6412 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  AND2_X1 U6413 ( .A1(n6246), .A2(n5019), .ZN(n6565) );
  OR2_X2 U6414 ( .A1(n6241), .A2(n9833), .ZN(n6244) );
  AND2_X1 U6415 ( .A1(n7419), .A2(n7365), .ZN(n7373) );
  NAND2_X1 U6416 ( .A1(n6122), .A2(n4704), .ZN(n7368) );
  NAND2_X1 U6417 ( .A1(n6265), .A2(n6264), .ZN(n6270) );
  OR2_X1 U6418 ( .A1(n6499), .A2(n4398), .ZN(n8086) );
  AND2_X1 U6419 ( .A1(n6475), .A2(n4398), .ZN(n9720) );
  OR2_X1 U6420 ( .A1(n9101), .A2(n9100), .ZN(n4927) );
  INV_X1 U6421 ( .A(n8253), .ZN(n7729) );
  OR2_X1 U6422 ( .A1(n5353), .A2(n5352), .ZN(n8870) );
  OR2_X1 U6423 ( .A1(n7676), .A2(n8378), .ZN(n4928) );
  AND2_X1 U6424 ( .A1(n6163), .A2(n6161), .ZN(n4930) );
  AND2_X1 U6425 ( .A1(n5819), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4932) );
  OR2_X1 U6426 ( .A1(n9472), .A2(n9108), .ZN(n4933) );
  OR2_X1 U6427 ( .A1(n7676), .A2(n8313), .ZN(n4934) );
  INV_X1 U6428 ( .A(n9060), .ZN(n8720) );
  AND2_X1 U6429 ( .A1(n5227), .A2(n5202), .ZN(n4937) );
  INV_X1 U6430 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6431 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4938) );
  INV_X2 U6432 ( .A(n9678), .ZN(n9304) );
  NAND2_X2 U6433 ( .A1(n6939), .A2(n9673), .ZN(n9678) );
  INV_X1 U6434 ( .A(n9744), .ZN(n5831) );
  INV_X1 U6435 ( .A(n9246), .ZN(n9101) );
  AND2_X1 U6436 ( .A1(n7955), .A2(n7245), .ZN(n4939) );
  INV_X1 U6437 ( .A(n8558), .ZN(n7344) );
  INV_X1 U6438 ( .A(n8435), .ZN(n6125) );
  NAND2_X1 U6439 ( .A1(n6125), .A2(n9549), .ZN(n6126) );
  NOR2_X1 U6440 ( .A1(n8363), .A2(n7495), .ZN(n7687) );
  OAI211_X1 U6441 ( .C1(n9060), .C2(n8722), .A(n8728), .B(n9073), .ZN(n8723)
         );
  INV_X1 U6442 ( .A(n7694), .ZN(n7695) );
  INV_X1 U6443 ( .A(n5358), .ZN(n5359) );
  INV_X1 U6444 ( .A(n8723), .ZN(n8724) );
  INV_X1 U6445 ( .A(n9099), .ZN(n9100) );
  NAND2_X1 U6446 ( .A1(n10068), .A2(n4929), .ZN(n4948) );
  INV_X1 U6447 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4940) );
  INV_X1 U6448 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6001) );
  INV_X1 U6449 ( .A(n7662), .ZN(n6064) );
  NAND2_X1 U6450 ( .A1(n9495), .A2(n9085), .ZN(n9086) );
  INV_X1 U6451 ( .A(SI_27_), .ZN(n9931) );
  INV_X1 U6452 ( .A(SI_25_), .ZN(n5597) );
  INV_X1 U6453 ( .A(SI_22_), .ZN(n5523) );
  INV_X1 U6454 ( .A(SI_19_), .ZN(n9934) );
  INV_X1 U6455 ( .A(SI_9_), .ZN(n9937) );
  INV_X1 U6456 ( .A(n6290), .ZN(n6287) );
  OR2_X1 U6457 ( .A1(n5836), .A2(n6959), .ZN(n5795) );
  NOR2_X1 U6458 ( .A1(n6201), .A2(n6799), .ZN(n6302) );
  INV_X1 U6459 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U6460 ( .A1(n5578), .A2(n8538), .ZN(n5603) );
  OR2_X1 U6461 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  INV_X1 U6462 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5422) );
  INV_X1 U6463 ( .A(n6365), .ZN(n5391) );
  OR2_X1 U6464 ( .A1(n9638), .A2(n9639), .ZN(n9641) );
  NAND2_X1 U6465 ( .A1(n9279), .A2(n9091), .ZN(n9094) );
  AND2_X1 U6466 ( .A1(n6372), .A2(n6571), .ZN(n6566) );
  NOR2_X1 U6467 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4949) );
  INV_X1 U6468 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5437) );
  INV_X1 U6469 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4945) );
  INV_X1 U6470 ( .A(n7958), .ZN(n6822) );
  INV_X1 U6471 ( .A(n6155), .ZN(n7701) );
  AND2_X1 U6472 ( .A1(n6441), .A2(n8445), .ZN(n6475) );
  AND2_X1 U6473 ( .A1(n8087), .A2(n6109), .ZN(n8106) );
  AND2_X1 U6474 ( .A1(n7589), .A2(n7585), .ZN(n7088) );
  INV_X1 U6475 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6242) );
  INV_X1 U6476 ( .A(n6204), .ZN(n6195) );
  AND2_X1 U6477 ( .A1(n7625), .A2(n7626), .ZN(n8264) );
  INV_X1 U6478 ( .A(n8275), .ZN(n8288) );
  OR2_X1 U6479 ( .A1(n7698), .A2(n7704), .ZN(n9798) );
  AND2_X1 U6480 ( .A1(n6294), .A2(n6385), .ZN(n6291) );
  INV_X1 U6481 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8538) );
  AND2_X1 U6482 ( .A1(n7267), .A2(n7266), .ZN(n5222) );
  OR2_X1 U6483 ( .A1(n5737), .A2(n5736), .ZN(n8601) );
  INV_X1 U6484 ( .A(n6571), .ZN(n8858) );
  NOR2_X1 U6485 ( .A1(n5509), .A2(n8490), .ZN(n5528) );
  INV_X1 U6486 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7270) );
  INV_X1 U6487 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6920) );
  INV_X1 U6488 ( .A(n9136), .ZN(n9148) );
  AND2_X1 U6489 ( .A1(n8764), .A2(n9190), .ZN(n9212) );
  AND2_X1 U6490 ( .A1(n8748), .A2(n8749), .ZN(n9290) );
  OR2_X1 U6491 ( .A1(n8558), .A2(n8871), .ZN(n7402) );
  OR2_X1 U6492 ( .A1(n8759), .A2(n6426), .ZN(n9051) );
  INV_X1 U6493 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5712) );
  OR2_X1 U6494 ( .A1(n6576), .A2(n8858), .ZN(n9698) );
  AOI21_X1 U6495 ( .B1(n9681), .B2(n6567), .A(n6566), .ZN(n6936) );
  AND2_X1 U6496 ( .A1(n5595), .A2(n5575), .ZN(n5593) );
  NOR2_X1 U6497 ( .A1(n7483), .A2(n7452), .ZN(n6187) );
  OR2_X1 U6498 ( .A1(n6309), .A2(n6310), .ZN(n7942) );
  INV_X1 U6499 ( .A(n7928), .ZN(n7944) );
  OR2_X1 U6500 ( .A1(n5838), .A2(n8087), .ZN(n7536) );
  NOR2_X1 U6501 ( .A1(n7210), .A2(n7209), .ZN(n7213) );
  INV_X1 U6502 ( .A(n8082), .ZN(n9887) );
  INV_X1 U6503 ( .A(n9880), .ZN(n9713) );
  NAND2_X1 U6504 ( .A1(n6254), .A2(n6253), .ZN(n6255) );
  INV_X1 U6505 ( .A(n8095), .ZN(n9750) );
  INV_X1 U6506 ( .A(n9757), .ZN(n8291) );
  NAND2_X1 U6507 ( .A1(n9833), .A2(n6242), .ZN(n6243) );
  INV_X1 U6508 ( .A(n8313), .ZN(n8349) );
  NOR2_X1 U6509 ( .A1(n6801), .A2(n6195), .ZN(n6196) );
  INV_X1 U6510 ( .A(n9793), .ZN(n9816) );
  AND2_X1 U6511 ( .A1(n5783), .A2(n6307), .ZN(n9786) );
  OR2_X1 U6512 ( .A1(n9786), .A2(n8354), .ZN(n9811) );
  AND2_X1 U6513 ( .A1(n6175), .A2(n6174), .ZN(n6799) );
  INV_X1 U6514 ( .A(n9575), .ZN(n8568) );
  AND2_X1 U6515 ( .A1(n6565), .A2(n5724), .ZN(n9302) );
  INV_X1 U6516 ( .A(n5732), .ZN(n8860) );
  OR2_X1 U6517 ( .A1(n9182), .A2(n5652), .ZN(n5609) );
  AND2_X1 U6518 ( .A1(n5326), .A2(n5325), .ZN(n7411) );
  AND2_X1 U6519 ( .A1(n6418), .A2(n9520), .ZN(n9630) );
  INV_X1 U6520 ( .A(n9619), .ZN(n9634) );
  OR2_X1 U6521 ( .A1(n6565), .A2(n6370), .ZN(n6377) );
  AND2_X1 U6522 ( .A1(n9678), .A2(n6943), .ZN(n9657) );
  INV_X1 U6523 ( .A(n9660), .ZN(n9350) );
  AOI21_X1 U6524 ( .B1(n5713), .B2(n5712), .A(n6392), .ZN(n6594) );
  AND2_X1 U6525 ( .A1(n9712), .A2(n9443), .ZN(n9367) );
  AND2_X1 U6526 ( .A1(n9707), .A2(n9443), .ZN(n9456) );
  INV_X1 U6527 ( .A(n6387), .ZN(n6247) );
  INV_X1 U6528 ( .A(n9738), .ZN(n9789) );
  AND2_X1 U6529 ( .A1(n6306), .A2(n6305), .ZN(n7928) );
  INV_X1 U6530 ( .A(n8394), .ZN(n7898) );
  AND2_X1 U6531 ( .A1(n6286), .A2(n6285), .ZN(n7932) );
  AND4_X1 U6532 ( .A1(n7536), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n7495)
         );
  NAND4_X1 U6533 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n8164)
         );
  INV_X1 U6534 ( .A(n8254), .ZN(n8228) );
  INV_X1 U6535 ( .A(n7424), .ZN(n9730) );
  INV_X1 U6536 ( .A(n9882), .ZN(n8050) );
  INV_X1 U6537 ( .A(n9720), .ZN(n9891) );
  NAND2_X1 U6538 ( .A1(n8291), .A2(n9552), .ZN(n8272) );
  NAND2_X1 U6539 ( .A1(n4275), .A2(n9816), .ZN(n8313) );
  INV_X1 U6540 ( .A(n8350), .ZN(n8344) );
  OR2_X1 U6541 ( .A1(n9819), .A2(n9804), .ZN(n8425) );
  AND3_X1 U6542 ( .A1(n8357), .A2(n8356), .A3(n8355), .ZN(n9760) );
  INV_X1 U6543 ( .A(n6399), .ZN(n6400) );
  INV_X1 U6544 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6358) );
  INV_X1 U6545 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8450) );
  INV_X1 U6546 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6450) );
  AND2_X1 U6547 ( .A1(n5735), .A2(n5734), .ZN(n9575) );
  OR2_X1 U6548 ( .A1(n5742), .A2(n5741), .ZN(n8868) );
  OAI21_X1 U6549 ( .B1(n9248), .B2(n5652), .A(n5514), .ZN(n9099) );
  OR2_X1 U6550 ( .A1(n5377), .A2(n5376), .ZN(n9082) );
  NAND2_X1 U6551 ( .A1(n6418), .A2(n9523), .ZN(n9619) );
  NAND2_X1 U6552 ( .A1(n6377), .A2(n6375), .ZN(n9650) );
  AND2_X1 U6553 ( .A1(n6935), .A2(n6934), .ZN(n9689) );
  INV_X1 U6554 ( .A(n9367), .ZN(n9440) );
  INV_X1 U6555 ( .A(n9712), .ZN(n9710) );
  INV_X1 U6556 ( .A(n9164), .ZN(n9464) );
  INV_X1 U6557 ( .A(n9263), .ZN(n9483) );
  AND2_X1 U6558 ( .A1(n9689), .A2(n9688), .ZN(n9708) );
  INV_X1 U6559 ( .A(n9707), .ZN(n9706) );
  AND2_X1 U6560 ( .A1(n7433), .A2(n7481), .ZN(n6392) );
  INV_X1 U6561 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10025) );
  INV_X1 U6562 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6950) );
  INV_X1 U6563 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6449) );
  NOR2_X2 U6564 ( .A1(n6434), .A2(n6247), .ZN(P2_U3893) );
  AND2_X2 U6565 ( .A1(n6246), .A2(n4732), .ZN(P1_U3973) );
  NOR2_X1 U6566 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4942) );
  NOR2_X1 U6567 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4941) );
  NAND2_X2 U6568 ( .A1(n4955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6569 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4950) );
  NAND3_X1 U6570 ( .A1(n4957), .A2(n5004), .A3(n4951), .ZN(n4954) );
  INV_X1 U6571 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6907) );
  INV_X1 U6572 ( .A(n5100), .ZN(n4962) );
  INV_X1 U6573 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5071) );
  INV_X1 U6574 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U6575 ( .A1(n5071), .A2(n4960), .ZN(n4961) );
  NAND2_X1 U6576 ( .A1(n4962), .A2(n4961), .ZN(n6736) );
  OAI22_X1 U6577 ( .A1(n8624), .A2(n6907), .B1(n5652), .B2(n6736), .ZN(n4967)
         );
  INV_X1 U6578 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n4965) );
  INV_X1 U6579 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n4964) );
  OAI22_X1 U6580 ( .A1(n4271), .A2(n4965), .B1(n8621), .B2(n4964), .ZN(n4966)
         );
  NAND3_X1 U6581 ( .A1(n5437), .A2(n4977), .A3(n4979), .ZN(n4968) );
  INV_X1 U6582 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6583 ( .A1(n4972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4973) );
  XNOR2_X1 U6584 ( .A(n4973), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6585 ( .A1(n4342), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6586 ( .A1(n5419), .A2(n4977), .ZN(n4978) );
  NAND2_X1 U6587 ( .A1(n5438), .A2(n5437), .ZN(n5440) );
  INV_X1 U6588 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6589 ( .A1(n4982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4983) );
  MUX2_X1 U6590 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4983), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n4985) );
  INV_X1 U6591 ( .A(n4987), .ZN(n4984) );
  NAND2_X1 U6592 ( .A1(n5719), .A2(n5732), .ZN(n5730) );
  AND2_X1 U6593 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4989) );
  NAND3_X1 U6594 ( .A1(n5815), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4991) );
  NAND2_X1 U6595 ( .A1(n5044), .A2(n4991), .ZN(n5025) );
  NAND2_X1 U6596 ( .A1(n5025), .A2(n4994), .ZN(n4997) );
  NAND2_X1 U6597 ( .A1(n4995), .A2(SI_1_), .ZN(n4996) );
  NAND2_X1 U6598 ( .A1(n4997), .A2(n4996), .ZN(n5059) );
  INV_X1 U6599 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6342) );
  INV_X1 U6600 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6338) );
  MUX2_X1 U6601 ( .A(n6342), .B(n6338), .S(n7521), .Z(n4998) );
  XNOR2_X1 U6602 ( .A(n4998), .B(SI_2_), .ZN(n5060) );
  INV_X1 U6603 ( .A(n4998), .ZN(n4999) );
  NAND2_X1 U6604 ( .A1(n4999), .A2(SI_2_), .ZN(n5000) );
  MUX2_X1 U6605 ( .A(n6339), .B(n9992), .S(n7521), .Z(n5001) );
  XNOR2_X1 U6606 ( .A(n5001), .B(SI_3_), .ZN(n5078) );
  INV_X1 U6607 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6608 ( .A1(n5002), .A2(SI_3_), .ZN(n5003) );
  MUX2_X1 U6609 ( .A(n6345), .B(n6344), .S(n7521), .Z(n5108) );
  XNOR2_X1 U6610 ( .A(n5108), .B(SI_4_), .ZN(n5106) );
  XNOR2_X1 U6611 ( .A(n5107), .B(n5106), .ZN(n6346) );
  NAND2_X1 U6612 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5006) );
  NAND2_X1 U6613 ( .A1(n5007), .A2(n5006), .ZN(n5008) );
  OR2_X1 U6614 ( .A1(n6346), .A2(n5061), .ZN(n5018) );
  OR2_X1 U6615 ( .A1(n5009), .A2(n5386), .ZN(n5079) );
  OR2_X1 U6616 ( .A1(n5010), .A2(n5386), .ZN(n5011) );
  AND2_X1 U6617 ( .A1(n5079), .A2(n5011), .ZN(n5013) );
  INV_X1 U6618 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6619 ( .A1(n5013), .A2(n5012), .ZN(n5112) );
  INV_X1 U6620 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6621 ( .A1(n5014), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6622 ( .A1(n5112), .A2(n5015), .ZN(n6906) );
  OR2_X1 U6623 ( .A1(n6373), .A2(n6906), .ZN(n5017) );
  OR2_X1 U6624 ( .A1(n8717), .A2(n6344), .ZN(n5016) );
  INV_X1 U6625 ( .A(n5730), .ZN(n5020) );
  INV_X2 U6626 ( .A(n5047), .ZN(n5689) );
  AOI22_X1 U6627 ( .A1(n8878), .A2(n4276), .B1(n6660), .B2(n5689), .ZN(n5095)
         );
  NAND2_X1 U6628 ( .A1(n8863), .A2(n8810), .ZN(n6570) );
  NAND2_X1 U6629 ( .A1(n6660), .A2(n5680), .ZN(n5021) );
  NAND2_X1 U6630 ( .A1(n6365), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5023) );
  INV_X1 U6631 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6413) );
  INV_X1 U6632 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6633 ( .A1(n4391), .A2(n5661), .ZN(n5030) );
  XNOR2_X1 U6634 ( .A(n5025), .B(n5026), .ZN(n5802) );
  INV_X1 U6635 ( .A(n5802), .ZN(n6343) );
  INV_X1 U6636 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6337) );
  INV_X1 U6637 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6638 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5027) );
  NAND2_X1 U6639 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  INV_X2 U6640 ( .A(n4278), .ZN(n5658) );
  INV_X1 U6641 ( .A(n5035), .ZN(n5033) );
  INV_X1 U6642 ( .A(n5034), .ZN(n5032) );
  NAND2_X1 U6643 ( .A1(n5033), .A2(n5032), .ZN(n5036) );
  NAND2_X1 U6644 ( .A1(n5035), .A2(n5034), .ZN(n5052) );
  INV_X1 U6645 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6379) );
  INV_X1 U6646 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9672) );
  OAI22_X1 U6647 ( .A1(n5037), .A2(n9672), .B1(n5740), .B2(n6379), .ZN(n5041)
         );
  INV_X1 U6648 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5039) );
  INV_X1 U6649 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5038) );
  OAI22_X1 U6650 ( .A1(n5391), .A2(n5039), .B1(n8621), .B2(n5038), .ZN(n5040)
         );
  OR2_X2 U6651 ( .A1(n5041), .A2(n5040), .ZN(n6581) );
  NAND2_X1 U6652 ( .A1(n6581), .A2(n5661), .ZN(n5046) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6654 ( .A1(n5043), .A2(n5042), .ZN(n5045) );
  AND2_X1 U6655 ( .A1(n5045), .A2(n5044), .ZN(n9525) );
  MUX2_X1 U6656 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9525), .S(n6373), .Z(n6585) );
  NAND2_X1 U6657 ( .A1(n5086), .A2(n6585), .ZN(n5050) );
  OAI211_X1 U6658 ( .C1(n6379), .C2(n5019), .A(n5046), .B(n5050), .ZN(n6424)
         );
  NAND2_X1 U6659 ( .A1(n6581), .A2(n5629), .ZN(n5049) );
  AOI22_X1 U6660 ( .A1(n5661), .A2(n6585), .B1(n4732), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6661 ( .A1(n5049), .A2(n5048), .ZN(n6423) );
  AOI22_X1 U6662 ( .A1(n6424), .A2(n6423), .B1(n5658), .B2(n5050), .ZN(n5051)
         );
  INV_X1 U6663 ( .A(n5052), .ZN(n6461) );
  NAND2_X1 U6664 ( .A1(n5685), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6665 ( .A1(n6365), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5057) );
  INV_X1 U6666 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5053) );
  OR2_X1 U6667 ( .A1(n5740), .A2(n5053), .ZN(n5056) );
  INV_X1 U6668 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6669 ( .A1(n8621), .A2(n5054), .ZN(n5055) );
  NAND4_X2 U6670 ( .A1(n5058), .A2(n5057), .A3(n5056), .A4(n5055), .ZN(n8880)
         );
  NAND2_X1 U6671 ( .A1(n8880), .A2(n5661), .ZN(n5066) );
  XNOR2_X1 U6672 ( .A(n5059), .B(n5060), .ZN(n6341) );
  OR2_X1 U6673 ( .A1(n5061), .A2(n6341), .ZN(n5064) );
  OR2_X1 U6674 ( .A1(n8717), .A2(n6338), .ZN(n5063) );
  XNOR2_X1 U6675 ( .A(n5079), .B(n4781), .ZN(n6415) );
  OR2_X1 U6676 ( .A1(n6373), .A2(n6415), .ZN(n5062) );
  AND3_X2 U6677 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n6731) );
  NAND2_X1 U6678 ( .A1(n9656), .A2(n5086), .ZN(n5065) );
  NAND2_X1 U6679 ( .A1(n5066), .A2(n5065), .ZN(n5067) );
  XNOR2_X1 U6680 ( .A(n5067), .B(n5658), .ZN(n5069) );
  AOI22_X1 U6681 ( .A1(n8880), .A2(n5629), .B1(n9656), .B2(n5689), .ZN(n5068)
         );
  NAND2_X1 U6682 ( .A1(n5069), .A2(n5068), .ZN(n5070) );
  NAND2_X1 U6683 ( .A1(n5685), .A2(n5071), .ZN(n5076) );
  NAND2_X1 U6684 ( .A1(n6365), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5075) );
  INV_X1 U6685 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6417) );
  OR2_X1 U6686 ( .A1(n5740), .A2(n6417), .ZN(n5074) );
  INV_X1 U6687 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5072) );
  OR2_X1 U6688 ( .A1(n8621), .A2(n5072), .ZN(n5073) );
  INV_X1 U6689 ( .A(n8879), .ZN(n6617) );
  XNOR2_X1 U6690 ( .A(n5077), .B(n5078), .ZN(n6340) );
  OR2_X1 U6691 ( .A1(n5061), .A2(n6340), .ZN(n5085) );
  OR2_X1 U6692 ( .A1(n8717), .A2(n9992), .ZN(n5084) );
  NAND2_X1 U6693 ( .A1(n5079), .A2(n4781), .ZN(n5080) );
  NAND2_X1 U6694 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  INV_X1 U6695 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U6696 ( .A(n5082), .B(n5081), .ZN(n6416) );
  OR2_X1 U6697 ( .A1(n6373), .A2(n6416), .ZN(n5083) );
  OAI22_X1 U6698 ( .A1(n6617), .A2(n4274), .B1(n8819), .B2(n5047), .ZN(n5091)
         );
  NAND2_X1 U6699 ( .A1(n8879), .A2(n5661), .ZN(n5088) );
  INV_X1 U6700 ( .A(n8819), .ZN(n6650) );
  NAND2_X1 U6701 ( .A1(n6650), .A2(n5086), .ZN(n5087) );
  NAND2_X1 U6702 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XNOR2_X1 U6703 ( .A(n5089), .B(n4278), .ZN(n5090) );
  XOR2_X1 U6704 ( .A(n5091), .B(n5090), .Z(n6681) );
  NAND2_X1 U6705 ( .A1(n6680), .A2(n6681), .ZN(n6679) );
  INV_X1 U6706 ( .A(n5090), .ZN(n5093) );
  INV_X1 U6707 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6708 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  NAND2_X1 U6709 ( .A1(n6679), .A2(n5094), .ZN(n6741) );
  INV_X1 U6710 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7179) );
  INV_X1 U6711 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6896) );
  OR2_X1 U6712 ( .A1(n4272), .A2(n6896), .ZN(n5098) );
  OAI21_X1 U6713 ( .B1(n8624), .B2(n7179), .A(n5098), .ZN(n5099) );
  INV_X1 U6714 ( .A(n5099), .ZN(n5105) );
  NAND2_X1 U6715 ( .A1(n5100), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5128) );
  OAI21_X1 U6716 ( .B1(n5100), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5128), .ZN(
        n7180) );
  INV_X1 U6717 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6718 ( .A1(n8621), .A2(n5101), .ZN(n5102) );
  OAI21_X1 U6719 ( .B1(n5652), .B2(n7180), .A(n5102), .ZN(n5103) );
  INV_X1 U6720 ( .A(n5103), .ZN(n5104) );
  INV_X1 U6721 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6722 ( .A1(n5109), .A2(SI_4_), .ZN(n5110) );
  MUX2_X1 U6723 ( .A(n6348), .B(n6347), .S(n7521), .Z(n5120) );
  XNOR2_X1 U6724 ( .A(n5119), .B(n5118), .ZN(n6349) );
  OR2_X1 U6725 ( .A1(n6349), .A2(n5061), .ZN(n5115) );
  NAND2_X1 U6726 ( .A1(n5112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U6727 ( .A(n5113), .B(P1_IR_REG_5__SCAN_IN), .ZN(n8926) );
  AOI22_X1 U6728 ( .A1(n5462), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5461), .B2(
        n8926), .ZN(n5114) );
  NAND2_X1 U6729 ( .A1(n5115), .A2(n5114), .ZN(n6870) );
  AOI22_X1 U6730 ( .A1(n8877), .A2(n5689), .B1(n6870), .B2(n5680), .ZN(n5116)
         );
  OAI22_X1 U6731 ( .A1(n6790), .A2(n5693), .B1(n7181), .B2(n5047), .ZN(n6866)
         );
  INV_X1 U6732 ( .A(n5117), .ZN(n6963) );
  INV_X1 U6733 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6734 ( .A1(n5121), .A2(SI_5_), .ZN(n5122) );
  MUX2_X1 U6735 ( .A(n6350), .B(n6352), .S(n7521), .Z(n5148) );
  XNOR2_X1 U6736 ( .A(n5147), .B(n5146), .ZN(n6351) );
  OR2_X1 U6737 ( .A1(n6351), .A2(n5061), .ZN(n5126) );
  NAND2_X1 U6738 ( .A1(n5123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U6739 ( .A(n5124), .B(P1_IR_REG_6__SCAN_IN), .ZN(n8940) );
  AOI22_X1 U6740 ( .A1(n5462), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5461), .B2(
        n8940), .ZN(n5125) );
  NAND2_X1 U6741 ( .A1(n6365), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5134) );
  INV_X1 U6742 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5127) );
  NOR2_X1 U6743 ( .A1(n5128), .A2(n5127), .ZN(n5156) );
  AND2_X1 U6744 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  NOR2_X1 U6745 ( .A1(n5156), .A2(n5129), .ZN(n6966) );
  NAND2_X1 U6746 ( .A1(n5685), .A2(n6966), .ZN(n5133) );
  INV_X1 U6747 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6897) );
  OR2_X1 U6748 ( .A1(n4272), .A2(n6897), .ZN(n5132) );
  INV_X1 U6749 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5130) );
  OR2_X1 U6750 ( .A1(n8621), .A2(n5130), .ZN(n5131) );
  NAND4_X1 U6751 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n8876)
         );
  NAND2_X1 U6752 ( .A1(n8876), .A2(n5661), .ZN(n5135) );
  OAI21_X1 U6753 ( .B1(n7167), .B2(n5136), .A(n5135), .ZN(n5137) );
  XNOR2_X1 U6754 ( .A(n5137), .B(n5658), .ZN(n5141) );
  OR2_X1 U6755 ( .A1(n7167), .A2(n5047), .ZN(n5139) );
  NAND2_X1 U6756 ( .A1(n8876), .A2(n4276), .ZN(n5138) );
  NAND2_X1 U6757 ( .A1(n5139), .A2(n5138), .ZN(n5142) );
  INV_X1 U6758 ( .A(n5142), .ZN(n5140) );
  NAND2_X1 U6759 ( .A1(n5141), .A2(n5140), .ZN(n5145) );
  INV_X1 U6760 ( .A(n5141), .ZN(n5143) );
  NAND2_X1 U6761 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  AND2_X1 U6762 ( .A1(n5145), .A2(n5144), .ZN(n6962) );
  INV_X1 U6763 ( .A(n5148), .ZN(n5149) );
  MUX2_X1 U6764 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7521), .Z(n5171) );
  XNOR2_X1 U6765 ( .A(n5171), .B(SI_7_), .ZN(n5169) );
  XNOR2_X1 U6766 ( .A(n5170), .B(n5169), .ZN(n6353) );
  NAND2_X1 U6767 ( .A1(n6353), .A2(n8716), .ZN(n5153) );
  NAND2_X1 U6768 ( .A1(n5150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5151) );
  XNOR2_X1 U6769 ( .A(n5151), .B(P1_IR_REG_7__SCAN_IN), .ZN(n8954) );
  AOI22_X1 U6770 ( .A1(n5462), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5461), .B2(
        n8954), .ZN(n5152) );
  NAND2_X1 U6771 ( .A1(n5153), .A2(n5152), .ZN(n7134) );
  INV_X1 U6772 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6944) );
  INV_X1 U6773 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6898) );
  OR2_X1 U6774 ( .A1(n4271), .A2(n6898), .ZN(n5154) );
  OAI21_X1 U6775 ( .B1(n8624), .B2(n6944), .A(n5154), .ZN(n5155) );
  INV_X1 U6776 ( .A(n5155), .ZN(n5162) );
  NAND2_X1 U6777 ( .A1(n5156), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5183) );
  OR2_X1 U6778 ( .A1(n5156), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6779 ( .A1(n5183), .A2(n5157), .ZN(n7033) );
  INV_X1 U6780 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5158) );
  OR2_X1 U6781 ( .A1(n8621), .A2(n5158), .ZN(n5159) );
  OAI21_X1 U6782 ( .B1(n5652), .B2(n7033), .A(n5159), .ZN(n5160) );
  INV_X1 U6783 ( .A(n5160), .ZN(n5161) );
  OAI22_X1 U6784 ( .A1(n9684), .A2(n5047), .B1(n7133), .B2(n5693), .ZN(n5166)
         );
  NAND2_X1 U6785 ( .A1(n7134), .A2(n5680), .ZN(n5164) );
  OR2_X1 U6786 ( .A1(n7133), .A2(n5047), .ZN(n5163) );
  NAND2_X1 U6787 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  XNOR2_X1 U6788 ( .A(n5165), .B(n4278), .ZN(n5167) );
  XOR2_X1 U6789 ( .A(n5166), .B(n5167), .Z(n7031) );
  NAND2_X1 U6790 ( .A1(n7029), .A2(n5168), .ZN(n5195) );
  NAND2_X1 U6791 ( .A1(n5171), .A2(SI_7_), .ZN(n5172) );
  MUX2_X1 U6792 ( .A(n6361), .B(n5173), .S(n7521), .Z(n5175) );
  INV_X1 U6793 ( .A(SI_8_), .ZN(n5174) );
  NAND2_X1 U6794 ( .A1(n5175), .A2(n5174), .ZN(n5198) );
  INV_X1 U6795 ( .A(n5175), .ZN(n5176) );
  NAND2_X1 U6796 ( .A1(n5176), .A2(SI_8_), .ZN(n5177) );
  NAND2_X1 U6797 ( .A1(n5198), .A2(n5177), .ZN(n5196) );
  NAND2_X1 U6798 ( .A1(n6359), .A2(n8716), .ZN(n5179) );
  NOR2_X1 U6799 ( .A1(n5150), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5231) );
  OR2_X1 U6800 ( .A1(n5231), .A2(n5386), .ZN(n5204) );
  XNOR2_X1 U6801 ( .A(n5204), .B(P1_IR_REG_8__SCAN_IN), .ZN(n8968) );
  AOI22_X1 U6802 ( .A1(n5462), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5461), .B2(
        n8968), .ZN(n5178) );
  NAND2_X1 U6803 ( .A1(n7139), .A2(n5680), .ZN(n5191) );
  INV_X1 U6804 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7006) );
  INV_X1 U6805 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6899) );
  OR2_X1 U6806 ( .A1(n4271), .A2(n6899), .ZN(n5180) );
  OAI21_X1 U6807 ( .B1(n8624), .B2(n7006), .A(n5180), .ZN(n5181) );
  INV_X1 U6808 ( .A(n5181), .ZN(n5189) );
  NAND2_X1 U6809 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  NAND2_X1 U6810 ( .A1(n5211), .A2(n5184), .ZN(n7282) );
  INV_X1 U6811 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5185) );
  OR2_X1 U6812 ( .A1(n8621), .A2(n5185), .ZN(n5186) );
  OAI21_X1 U6813 ( .B1(n5652), .B2(n7282), .A(n5186), .ZN(n5187) );
  INV_X1 U6814 ( .A(n5187), .ZN(n5188) );
  OR2_X1 U6815 ( .A1(n7153), .A2(n5047), .ZN(n5190) );
  NAND2_X1 U6816 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  XNOR2_X1 U6817 ( .A(n5192), .B(n4278), .ZN(n5193) );
  AOI22_X1 U6818 ( .A1(n7139), .A2(n5661), .B1(n4276), .B2(n4649), .ZN(n7280)
         );
  INV_X1 U6819 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6820 ( .A1(n5195), .A2(n5194), .ZN(n7267) );
  INV_X1 U6821 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6395) );
  INV_X1 U6822 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5199) );
  MUX2_X1 U6823 ( .A(n6395), .B(n5199), .S(n7521), .Z(n5200) );
  NAND2_X1 U6824 ( .A1(n5200), .A2(n9937), .ZN(n5227) );
  INV_X1 U6825 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6826 ( .A1(n5201), .A2(SI_9_), .ZN(n5202) );
  XNOR2_X1 U6827 ( .A(n5226), .B(n4937), .ZN(n6388) );
  INV_X1 U6828 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6829 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U6830 ( .A1(n5205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6831 ( .A(n5206), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8984) );
  AOI22_X1 U6832 ( .A1(n5462), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5461), .B2(
        n8984), .ZN(n5207) );
  NAND2_X1 U6833 ( .A1(n9690), .A2(n5680), .ZN(n5219) );
  INV_X1 U6834 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7155) );
  INV_X1 U6835 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6836 ( .A1(n4271), .A2(n5208), .ZN(n5209) );
  OAI21_X1 U6837 ( .B1(n8624), .B2(n7155), .A(n5209), .ZN(n5210) );
  INV_X1 U6838 ( .A(n5210), .ZN(n5217) );
  AND2_X1 U6839 ( .A1(n5211), .A2(n7270), .ZN(n5212) );
  OR2_X1 U6840 ( .A1(n5212), .A2(n5235), .ZN(n7273) );
  INV_X1 U6841 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6842 ( .A1(n8621), .A2(n5213), .ZN(n5214) );
  OAI21_X1 U6843 ( .B1(n5652), .B2(n7273), .A(n5214), .ZN(n5215) );
  INV_X1 U6844 ( .A(n5215), .ZN(n5216) );
  OR2_X1 U6845 ( .A1(n7142), .A2(n5047), .ZN(n5218) );
  NAND2_X1 U6846 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  XNOR2_X1 U6847 ( .A(n5220), .B(n4278), .ZN(n5223) );
  NOR2_X1 U6848 ( .A1(n7142), .A2(n5693), .ZN(n5221) );
  AOI21_X1 U6849 ( .B1(n9690), .B2(n5689), .A(n5221), .ZN(n5224) );
  XNOR2_X1 U6850 ( .A(n5223), .B(n5224), .ZN(n7266) );
  INV_X1 U6851 ( .A(n5223), .ZN(n5225) );
  INV_X1 U6852 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6397) );
  INV_X1 U6853 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6854 ( .A(n6397), .B(n5229), .S(n7521), .Z(n5253) );
  XNOR2_X1 U6855 ( .A(n5253), .B(SI_10_), .ZN(n5252) );
  NAND2_X1 U6856 ( .A1(n6393), .A2(n8716), .ZN(n5234) );
  NOR2_X1 U6857 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5230) );
  AND2_X1 U6858 ( .A1(n5231), .A2(n5230), .ZN(n5262) );
  OR2_X1 U6859 ( .A1(n5262), .A2(n5386), .ZN(n5232) );
  XNOR2_X1 U6860 ( .A(n5232), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9534) );
  AOI22_X1 U6861 ( .A1(n5462), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5461), .B2(
        n9534), .ZN(n5233) );
  NAND2_X1 U6862 ( .A1(n5234), .A2(n5233), .ZN(n7255) );
  NOR2_X1 U6863 ( .A1(n5235), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5236) );
  OR2_X1 U6864 ( .A1(n5266), .A2(n5236), .ZN(n9574) );
  INV_X1 U6865 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6866 ( .A1(n4271), .A2(n5237), .ZN(n5238) );
  OAI21_X1 U6867 ( .B1(n5652), .B2(n9574), .A(n5238), .ZN(n5239) );
  INV_X1 U6868 ( .A(n5239), .ZN(n5244) );
  INV_X1 U6869 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7145) );
  INV_X1 U6870 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6871 ( .A1(n4420), .A2(n5240), .ZN(n5241) );
  OAI21_X1 U6872 ( .B1(n8624), .B2(n7145), .A(n5241), .ZN(n5242) );
  INV_X1 U6873 ( .A(n5242), .ZN(n5243) );
  AOI22_X1 U6874 ( .A1(n7255), .A2(n5680), .B1(n5689), .B2(n8874), .ZN(n5245)
         );
  XOR2_X1 U6875 ( .A(n4278), .B(n5245), .Z(n5246) );
  NOR2_X2 U6876 ( .A1(n5247), .A2(n5246), .ZN(n5249) );
  NOR2_X1 U6877 ( .A1(n5249), .A2(n5248), .ZN(n9561) );
  AOI22_X1 U6878 ( .A1(n7255), .A2(n5689), .B1(n4276), .B2(n8874), .ZN(n9562)
         );
  INV_X1 U6879 ( .A(n5249), .ZN(n5250) );
  INV_X1 U6880 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6881 ( .A1(n5254), .A2(SI_10_), .ZN(n5255) );
  MUX2_X1 U6882 ( .A(n6403), .B(n9920), .S(n7521), .Z(n5258) );
  INV_X1 U6883 ( .A(SI_11_), .ZN(n5257) );
  NAND2_X1 U6884 ( .A1(n5258), .A2(n5257), .ZN(n5283) );
  INV_X1 U6885 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6886 ( .A1(n5259), .A2(SI_11_), .ZN(n5260) );
  NAND2_X1 U6887 ( .A1(n5283), .A2(n5260), .ZN(n5282) );
  NAND2_X1 U6888 ( .A1(n6401), .A2(n8716), .ZN(n5265) );
  INV_X1 U6889 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5261) );
  AND2_X1 U6890 ( .A1(n5262), .A2(n5261), .ZN(n5285) );
  INV_X1 U6891 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6892 ( .A1(n5285), .A2(n5386), .ZN(n5263) );
  XNOR2_X1 U6893 ( .A(n5263), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9579) );
  AOI22_X1 U6894 ( .A1(n5462), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5461), .B2(
        n9579), .ZN(n5264) );
  NAND2_X1 U6895 ( .A1(n8581), .A2(n5680), .ZN(n5277) );
  NAND2_X1 U6896 ( .A1(n5266), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5291) );
  OR2_X1 U6897 ( .A1(n5266), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6898 ( .A1(n5291), .A2(n5267), .ZN(n8579) );
  INV_X1 U6899 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6900 ( .A1(n4271), .A2(n5268), .ZN(n5269) );
  OAI21_X1 U6901 ( .B1(n5652), .B2(n8579), .A(n5269), .ZN(n5270) );
  INV_X1 U6902 ( .A(n5270), .ZN(n5275) );
  INV_X1 U6903 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7259) );
  INV_X1 U6904 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5271) );
  OR2_X1 U6905 ( .A1(n4420), .A2(n5271), .ZN(n5272) );
  OAI21_X1 U6906 ( .B1(n8624), .B2(n7259), .A(n5272), .ZN(n5273) );
  INV_X1 U6907 ( .A(n5273), .ZN(n5274) );
  OR2_X1 U6908 ( .A1(n7301), .A2(n5047), .ZN(n5276) );
  NAND2_X1 U6909 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  XNOR2_X1 U6910 ( .A(n5278), .B(n5658), .ZN(n5281) );
  NOR2_X1 U6911 ( .A1(n7301), .A2(n5693), .ZN(n5279) );
  AOI21_X1 U6912 ( .B1(n8581), .B2(n5689), .A(n5279), .ZN(n5280) );
  OR2_X1 U6913 ( .A1(n5281), .A2(n5280), .ZN(n8573) );
  NAND2_X1 U6914 ( .A1(n5281), .A2(n5280), .ZN(n8575) );
  MUX2_X1 U6915 ( .A(n6450), .B(n6449), .S(n7521), .Z(n5306) );
  XNOR2_X1 U6916 ( .A(n5306), .B(SI_12_), .ZN(n5305) );
  XNOR2_X1 U6917 ( .A(n5309), .B(n5305), .ZN(n6448) );
  NAND2_X1 U6918 ( .A1(n6448), .A2(n8716), .ZN(n5287) );
  INV_X1 U6919 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6920 ( .A1(n5285), .A2(n5284), .ZN(n5343) );
  NAND2_X1 U6921 ( .A1(n5343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U6922 ( .A(n5310), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8999) );
  AOI22_X1 U6923 ( .A1(n5462), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5461), .B2(
        n8999), .ZN(n5286) );
  NAND2_X1 U6924 ( .A1(n8502), .A2(n5680), .ZN(n5299) );
  INV_X1 U6925 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7305) );
  INV_X1 U6926 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5288) );
  OR2_X1 U6927 ( .A1(n4272), .A2(n5288), .ZN(n5289) );
  OAI21_X1 U6928 ( .B1(n8624), .B2(n7305), .A(n5289), .ZN(n5290) );
  INV_X1 U6929 ( .A(n5290), .ZN(n5297) );
  NAND2_X1 U6930 ( .A1(n5291), .A2(n6920), .ZN(n5292) );
  NAND2_X1 U6931 ( .A1(n5320), .A2(n5292), .ZN(n8500) );
  INV_X1 U6932 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5293) );
  OR2_X1 U6933 ( .A1(n4420), .A2(n5293), .ZN(n5294) );
  OAI21_X1 U6934 ( .B1(n5652), .B2(n8500), .A(n5294), .ZN(n5295) );
  INV_X1 U6935 ( .A(n5295), .ZN(n5296) );
  OR2_X1 U6936 ( .A1(n7337), .A2(n5047), .ZN(n5298) );
  NAND2_X1 U6937 ( .A1(n5299), .A2(n5298), .ZN(n5301) );
  XNOR2_X1 U6938 ( .A(n5301), .B(n4278), .ZN(n5302) );
  INV_X1 U6939 ( .A(n7337), .ZN(n8872) );
  AOI22_X1 U6940 ( .A1(n8502), .A2(n5661), .B1(n4276), .B2(n8872), .ZN(n5303)
         );
  XNOR2_X1 U6941 ( .A(n5302), .B(n5303), .ZN(n8495) );
  INV_X1 U6942 ( .A(n5302), .ZN(n5304) );
  INV_X1 U6943 ( .A(n5305), .ZN(n5308) );
  INV_X1 U6944 ( .A(n5306), .ZN(n5307) );
  MUX2_X1 U6945 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7521), .Z(n5337) );
  XNOR2_X1 U6946 ( .A(n5337), .B(SI_13_), .ZN(n5334) );
  XNOR2_X1 U6947 ( .A(n5336), .B(n5334), .ZN(n6455) );
  NAND2_X1 U6948 ( .A1(n6455), .A2(n8716), .ZN(n5314) );
  INV_X1 U6949 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6950 ( .A1(n5310), .A2(n5341), .ZN(n5311) );
  NAND2_X1 U6951 ( .A1(n5311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6952 ( .A(n5312), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U6953 ( .A1(n5462), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5461), .B2(
        n9593), .ZN(n5313) );
  INV_X1 U6954 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5317) );
  INV_X1 U6955 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5315) );
  OR2_X1 U6956 ( .A1(n4272), .A2(n5315), .ZN(n5316) );
  OAI21_X1 U6957 ( .B1(n8624), .B2(n5317), .A(n5316), .ZN(n5318) );
  INV_X1 U6958 ( .A(n5318), .ZN(n5326) );
  NAND2_X1 U6959 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U6960 ( .A1(n5349), .A2(n5321), .ZN(n8556) );
  INV_X1 U6961 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5322) );
  OR2_X1 U6962 ( .A1(n4420), .A2(n5322), .ZN(n5323) );
  OAI21_X1 U6963 ( .B1(n5652), .B2(n8556), .A(n5323), .ZN(n5324) );
  INV_X1 U6964 ( .A(n5324), .ZN(n5325) );
  INV_X1 U6965 ( .A(n7411), .ZN(n8871) );
  AOI22_X1 U6966 ( .A1(n8558), .A2(n5689), .B1(n4276), .B2(n8871), .ZN(n5330)
         );
  NAND2_X1 U6967 ( .A1(n8558), .A2(n5680), .ZN(n5328) );
  OR2_X1 U6968 ( .A1(n7411), .A2(n5047), .ZN(n5327) );
  NAND2_X1 U6969 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  XNOR2_X1 U6970 ( .A(n5329), .B(n4278), .ZN(n5332) );
  XOR2_X1 U6971 ( .A(n5330), .B(n5332), .Z(n8552) );
  INV_X1 U6972 ( .A(n5330), .ZN(n5331) );
  INV_X1 U6973 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6974 ( .A1(n5336), .A2(n5335), .ZN(n5339) );
  NAND2_X1 U6975 ( .A1(n5337), .A2(SI_13_), .ZN(n5338) );
  NAND2_X1 U6976 ( .A1(n5339), .A2(n5338), .ZN(n5363) );
  XNOR2_X1 U6977 ( .A(n5364), .B(SI_14_), .ZN(n5361) );
  XNOR2_X1 U6978 ( .A(n5363), .B(n5361), .ZN(n6512) );
  NAND2_X1 U6979 ( .A1(n6512), .A2(n8716), .ZN(n5346) );
  INV_X1 U6980 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6981 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  OAI21_X1 U6982 ( .B1(n5343), .B2(n5342), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5344) );
  XNOR2_X1 U6983 ( .A(n5344), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9608) );
  AOI22_X1 U6984 ( .A1(n5462), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5461), .B2(
        n9608), .ZN(n5345) );
  NAND2_X1 U6985 ( .A1(n9442), .A2(n5680), .ZN(n5355) );
  INV_X1 U6986 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5348) );
  INV_X1 U6987 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5347) );
  OAI22_X1 U6988 ( .A1(n8624), .A2(n5348), .B1(n4272), .B2(n5347), .ZN(n5353)
         );
  AND2_X1 U6989 ( .A1(n5349), .A2(n8458), .ZN(n5350) );
  OR2_X1 U6990 ( .A1(n5350), .A2(n5392), .ZN(n7405) );
  INV_X1 U6991 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5351) );
  OAI22_X1 U6992 ( .A1(n5652), .A2(n7405), .B1(n4420), .B2(n5351), .ZN(n5352)
         );
  NAND2_X1 U6993 ( .A1(n8870), .A2(n5689), .ZN(n5354) );
  NAND2_X1 U6994 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  XNOR2_X1 U6995 ( .A(n5356), .B(n4278), .ZN(n5358) );
  AOI22_X1 U6996 ( .A1(n9442), .A2(n5689), .B1(n4276), .B2(n8870), .ZN(n8455)
         );
  INV_X1 U6997 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6998 ( .A1(n5364), .A2(SI_14_), .ZN(n5365) );
  NOR2_X1 U6999 ( .A1(n5367), .A2(n9943), .ZN(n5366) );
  NAND2_X1 U7000 ( .A1(n5367), .A2(n9943), .ZN(n5368) );
  XNOR2_X1 U7001 ( .A(n5410), .B(SI_16_), .ZN(n5369) );
  XNOR2_X1 U7002 ( .A(n5414), .B(n5369), .ZN(n6686) );
  NAND2_X1 U7003 ( .A1(n6686), .A2(n8716), .ZN(n5373) );
  NAND2_X1 U7004 ( .A1(n5370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U7005 ( .A(n5371), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9013) );
  AOI22_X1 U7006 ( .A1(n5462), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5461), .B2(
        n9013), .ZN(n5372) );
  NAND2_X1 U7007 ( .A1(n9344), .A2(n5680), .ZN(n5379) );
  NAND2_X1 U7008 ( .A1(n5392), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5394) );
  INV_X1 U7009 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U7010 ( .A1(n5394), .A2(n5374), .ZN(n5375) );
  NAND2_X1 U7011 ( .A1(n5423), .A2(n5375), .ZN(n9346) );
  INV_X1 U7012 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9497) );
  OAI22_X1 U7013 ( .A1(n9346), .A2(n5652), .B1(n4420), .B2(n9497), .ZN(n5377)
         );
  INV_X1 U7014 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9347) );
  INV_X1 U7015 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9999) );
  OAI22_X1 U7016 ( .A1(n8624), .A2(n9347), .B1(n4272), .B2(n9999), .ZN(n5376)
         );
  NAND2_X1 U7017 ( .A1(n9082), .A2(n5689), .ZN(n5378) );
  NAND2_X1 U7018 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  XNOR2_X1 U7019 ( .A(n5380), .B(n4278), .ZN(n8518) );
  INV_X1 U7020 ( .A(n9082), .ZN(n8625) );
  OAI22_X1 U7021 ( .A1(n9499), .A2(n5047), .B1(n8625), .B2(n5693), .ZN(n5404)
         );
  XNOR2_X1 U7022 ( .A(n5381), .B(SI_15_), .ZN(n5382) );
  XNOR2_X1 U7023 ( .A(n5383), .B(n5382), .ZN(n6626) );
  NAND2_X1 U7024 ( .A1(n6626), .A2(n8716), .ZN(n5390) );
  NOR2_X1 U7025 ( .A1(n5384), .A2(n5386), .ZN(n5385) );
  MUX2_X1 U7026 ( .A(n5386), .B(n5385), .S(P1_IR_REG_15__SCAN_IN), .Z(n5387)
         );
  INV_X1 U7027 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U7028 ( .A1(n5388), .A2(n5370), .ZN(n9002) );
  INV_X1 U7029 ( .A(n9002), .ZN(n9629) );
  AOI22_X1 U7030 ( .A1(n5462), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5461), .B2(
        n9629), .ZN(n5389) );
  NAND2_X1 U7031 ( .A1(n9078), .A2(n5689), .ZN(n5398) );
  INV_X1 U7032 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9625) );
  INV_X1 U7033 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9621) );
  OAI22_X1 U7034 ( .A1(n5645), .A2(n9625), .B1(n4271), .B2(n9621), .ZN(n5396)
         );
  OR2_X1 U7035 ( .A1(n5392), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U7036 ( .A1(n5394), .A2(n5393), .ZN(n8611) );
  INV_X1 U7037 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9501) );
  OAI22_X1 U7038 ( .A1(n5652), .A2(n8611), .B1(n4420), .B2(n9501), .ZN(n5395)
         );
  NAND2_X1 U7039 ( .A1(n9077), .A2(n4276), .ZN(n5397) );
  NAND2_X1 U7040 ( .A1(n5398), .A2(n5397), .ZN(n8607) );
  NAND2_X1 U7041 ( .A1(n9078), .A2(n5680), .ZN(n5400) );
  NAND2_X1 U7042 ( .A1(n9077), .A2(n5689), .ZN(n5399) );
  NAND2_X1 U7043 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  XNOR2_X1 U7044 ( .A(n5401), .B(n4278), .ZN(n5403) );
  AOI22_X1 U7045 ( .A1(n8518), .A2(n5404), .B1(n8607), .B2(n5403), .ZN(n5402)
         );
  INV_X1 U7046 ( .A(n8607), .ZN(n5406) );
  INV_X1 U7047 ( .A(n5404), .ZN(n8519) );
  AOI21_X1 U7048 ( .B1(n8517), .B2(n5406), .A(n8519), .ZN(n5405) );
  NAND3_X1 U7049 ( .A1(n8519), .A2(n5406), .A3(n8517), .ZN(n5407) );
  NOR2_X1 U7050 ( .A1(n5411), .A2(SI_16_), .ZN(n5413) );
  NAND2_X1 U7051 ( .A1(n5411), .A2(SI_16_), .ZN(n5412) );
  NAND2_X1 U7052 ( .A1(n5416), .A2(n5415), .ZN(n5433) );
  INV_X1 U7053 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U7054 ( .A1(n5417), .A2(SI_17_), .ZN(n5418) );
  NAND2_X1 U7055 ( .A1(n5433), .A2(n5418), .ZN(n5434) );
  XNOR2_X1 U7056 ( .A(n5435), .B(n5434), .ZN(n6828) );
  NAND2_X1 U7057 ( .A1(n6828), .A2(n8716), .ZN(n5421) );
  XNOR2_X1 U7058 ( .A(n5419), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9031) );
  AOI22_X1 U7059 ( .A1(n5462), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5461), .B2(
        n9031), .ZN(n5420) );
  AND2_X1 U7060 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  OR2_X1 U7061 ( .A1(n5424), .A2(n5443), .ZN(n9322) );
  INV_X1 U7062 ( .A(n4272), .ZN(n5468) );
  INV_X1 U7063 ( .A(n4420), .ZN(n5467) );
  AOI22_X1 U7064 ( .A1(n5468), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5467), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7065 ( .A1(n6365), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5425) );
  OAI211_X1 U7066 ( .C1(n9322), .C2(n5652), .A(n5426), .B(n5425), .ZN(n9083)
         );
  AND2_X1 U7067 ( .A1(n9083), .A2(n4276), .ZN(n5427) );
  AOI21_X1 U7068 ( .B1(n9321), .B2(n5689), .A(n5427), .ZN(n5429) );
  AOI22_X1 U7069 ( .A1(n9321), .A2(n5680), .B1(n5689), .B2(n9083), .ZN(n5428)
         );
  XNOR2_X1 U7070 ( .A(n5428), .B(n4278), .ZN(n5430) );
  XOR2_X1 U7071 ( .A(n5429), .B(n5430), .Z(n8527) );
  NAND2_X1 U7072 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  XNOR2_X1 U7073 ( .A(n5454), .B(SI_18_), .ZN(n5453) );
  XNOR2_X1 U7074 ( .A(n5457), .B(n5453), .ZN(n6862) );
  NAND2_X1 U7075 ( .A1(n6862), .A2(n8716), .ZN(n5442) );
  OR2_X1 U7076 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  AND2_X1 U7077 ( .A1(n5440), .A2(n5439), .ZN(n9028) );
  AOI22_X1 U7078 ( .A1(n5462), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5461), .B2(
        n9028), .ZN(n5441) );
  NAND2_X1 U7079 ( .A1(n9300), .A2(n5680), .ZN(n5448) );
  NOR2_X1 U7080 ( .A1(n5443), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5444) );
  OR2_X1 U7081 ( .A1(n5465), .A2(n5444), .ZN(n9301) );
  AOI22_X1 U7082 ( .A1(n6365), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5468), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5446) );
  INV_X1 U7083 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9489) );
  OR2_X1 U7084 ( .A1(n4420), .A2(n9489), .ZN(n5445) );
  OAI211_X1 U7085 ( .C1(n9301), .C2(n5652), .A(n5446), .B(n5445), .ZN(n9088)
         );
  NAND2_X1 U7086 ( .A1(n9088), .A2(n5661), .ZN(n5447) );
  NAND2_X1 U7087 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  XNOR2_X1 U7088 ( .A(n5449), .B(n5658), .ZN(n8585) );
  AND2_X1 U7089 ( .A1(n9088), .A2(n4276), .ZN(n5450) );
  AOI21_X1 U7090 ( .B1(n9300), .B2(n5689), .A(n5450), .ZN(n5451) );
  INV_X1 U7091 ( .A(n8585), .ZN(n5452) );
  INV_X1 U7092 ( .A(n5451), .ZN(n8584) );
  INV_X1 U7093 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U7094 ( .A1(n5455), .A2(SI_18_), .ZN(n5456) );
  NAND2_X1 U7095 ( .A1(n5458), .A2(n9934), .ZN(n5482) );
  INV_X1 U7096 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U7097 ( .A1(n5459), .A2(SI_19_), .ZN(n5460) );
  NAND2_X1 U7098 ( .A1(n5482), .A2(n5460), .ZN(n5481) );
  XNOR2_X1 U7099 ( .A(n5480), .B(n5481), .ZN(n7012) );
  NAND2_X1 U7100 ( .A1(n7012), .A2(n8716), .ZN(n5464) );
  INV_X1 U7101 ( .A(n8810), .ZN(n9040) );
  AOI22_X1 U7102 ( .A1(n5462), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9040), .B2(
        n5461), .ZN(n5463) );
  NAND2_X1 U7103 ( .A1(n9279), .A2(n5680), .ZN(n5472) );
  OR2_X1 U7104 ( .A1(n5465), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7105 ( .A1(n5486), .A2(n5466), .ZN(n9280) );
  AOI22_X1 U7106 ( .A1(n5468), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5467), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7107 ( .A1(n6365), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5469) );
  OAI211_X1 U7108 ( .C1(n9280), .C2(n5652), .A(n5470), .B(n5469), .ZN(n9091)
         );
  NAND2_X1 U7109 ( .A1(n9091), .A2(n5689), .ZN(n5471) );
  NAND2_X1 U7110 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  XNOR2_X1 U7111 ( .A(n5473), .B(n4278), .ZN(n5476) );
  NAND2_X1 U7112 ( .A1(n9279), .A2(n5661), .ZN(n5475) );
  NAND2_X1 U7113 ( .A1(n9091), .A2(n4276), .ZN(n5474) );
  NAND2_X1 U7114 ( .A1(n5475), .A2(n5474), .ZN(n5477) );
  NAND2_X1 U7115 ( .A1(n5476), .A2(n5477), .ZN(n8479) );
  INV_X1 U7116 ( .A(n5476), .ZN(n5479) );
  INV_X1 U7117 ( .A(n5477), .ZN(n5478) );
  NAND2_X1 U7118 ( .A1(n5479), .A2(n5478), .ZN(n8481) );
  XNOR2_X1 U7119 ( .A(n5500), .B(n9979), .ZN(n5483) );
  XNOR2_X1 U7120 ( .A(n5502), .B(n5483), .ZN(n7110) );
  NAND2_X1 U7121 ( .A1(n7110), .A2(n8716), .ZN(n5485) );
  INV_X1 U7122 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10004) );
  OR2_X1 U7123 ( .A1(n8717), .A2(n10004), .ZN(n5484) );
  INV_X1 U7124 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U7125 ( .A1(n5486), .A2(n8548), .ZN(n5487) );
  AND2_X1 U7126 ( .A1(n5509), .A2(n5487), .ZN(n9264) );
  NAND2_X1 U7127 ( .A1(n9264), .A2(n5685), .ZN(n5493) );
  INV_X1 U7128 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5490) );
  INV_X1 U7129 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9481) );
  OR2_X1 U7130 ( .A1(n4420), .A2(n9481), .ZN(n5489) );
  INV_X1 U7131 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9415) );
  OR2_X1 U7132 ( .A1(n4272), .A2(n9415), .ZN(n5488) );
  OAI211_X1 U7133 ( .C1(n8624), .C2(n5490), .A(n5489), .B(n5488), .ZN(n5491)
         );
  INV_X1 U7134 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U7135 ( .A1(n5493), .A2(n5492), .ZN(n9096) );
  INV_X1 U7136 ( .A(n9096), .ZN(n9098) );
  OAI22_X1 U7137 ( .A1(n9483), .A2(n5047), .B1(n9098), .B2(n5693), .ZN(n5497)
         );
  NAND2_X1 U7138 ( .A1(n9263), .A2(n5680), .ZN(n5495) );
  NAND2_X1 U7139 ( .A1(n9096), .A2(n5661), .ZN(n5494) );
  NAND2_X1 U7140 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  XNOR2_X1 U7141 ( .A(n5496), .B(n4278), .ZN(n5498) );
  XOR2_X1 U7142 ( .A(n5497), .B(n5498), .Z(n8545) );
  NAND2_X1 U7143 ( .A1(n8544), .A2(n8545), .ZN(n8543) );
  OR2_X1 U7144 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  INV_X1 U7145 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U7146 ( .A1(n5502), .A2(n9979), .ZN(n5503) );
  INV_X1 U7147 ( .A(SI_21_), .ZN(n5505) );
  XNOR2_X1 U7148 ( .A(n5520), .B(n5505), .ZN(n5506) );
  XNOR2_X1 U7149 ( .A(n5522), .B(n5506), .ZN(n6038) );
  NAND2_X1 U7150 ( .A1(n6038), .A2(n8716), .ZN(n5508) );
  INV_X1 U7151 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7204) );
  OR2_X1 U7152 ( .A1(n8717), .A2(n7204), .ZN(n5507) );
  INV_X1 U7153 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8490) );
  AND2_X1 U7154 ( .A1(n5509), .A2(n8490), .ZN(n5510) );
  OR2_X1 U7155 ( .A1(n5510), .A2(n5528), .ZN(n9248) );
  INV_X1 U7156 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9247) );
  INV_X1 U7157 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9478) );
  OR2_X1 U7158 ( .A1(n4420), .A2(n9478), .ZN(n5512) );
  INV_X1 U7159 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9410) );
  OR2_X1 U7160 ( .A1(n4271), .A2(n9410), .ZN(n5511) );
  OAI211_X1 U7161 ( .C1(n5645), .C2(n9247), .A(n5512), .B(n5511), .ZN(n5513)
         );
  INV_X1 U7162 ( .A(n5513), .ZN(n5514) );
  OAI22_X1 U7163 ( .A1(n9101), .A2(n5047), .B1(n9100), .B2(n5693), .ZN(n5518)
         );
  NAND2_X1 U7164 ( .A1(n9246), .A2(n5680), .ZN(n5516) );
  NAND2_X1 U7165 ( .A1(n9099), .A2(n5689), .ZN(n5515) );
  NAND2_X1 U7166 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  XNOR2_X1 U7167 ( .A(n5517), .B(n4278), .ZN(n5519) );
  XOR2_X1 U7168 ( .A(n5518), .B(n5519), .Z(n8488) );
  NAND2_X1 U7169 ( .A1(n5520), .A2(SI_21_), .ZN(n5521) );
  NAND2_X1 U7170 ( .A1(n5524), .A2(n5523), .ZN(n5541) );
  INV_X1 U7171 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U7172 ( .A1(n5525), .A2(SI_22_), .ZN(n5526) );
  NAND2_X1 U7173 ( .A1(n5541), .A2(n5526), .ZN(n5542) );
  OR2_X1 U7174 ( .A1(n8717), .A2(n9936), .ZN(n5527) );
  NAND2_X1 U7175 ( .A1(n9231), .A2(n5661), .ZN(n5537) );
  NAND2_X1 U7176 ( .A1(n5528), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5551) );
  OR2_X1 U7177 ( .A1(n5528), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7178 ( .A1(n5551), .A2(n5529), .ZN(n8565) );
  OR2_X1 U7179 ( .A1(n8565), .A2(n5652), .ZN(n5535) );
  INV_X1 U7180 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5532) );
  INV_X1 U7181 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9474) );
  OR2_X1 U7182 ( .A1(n4420), .A2(n9474), .ZN(n5531) );
  INV_X1 U7183 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9945) );
  OR2_X1 U7184 ( .A1(n4272), .A2(n9945), .ZN(n5530) );
  OAI211_X1 U7185 ( .C1(n5645), .C2(n5532), .A(n5531), .B(n5530), .ZN(n5533)
         );
  INV_X1 U7186 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7187 ( .A1(n5535), .A2(n5534), .ZN(n9104) );
  NAND2_X1 U7188 ( .A1(n9104), .A2(n4276), .ZN(n5536) );
  NAND2_X1 U7189 ( .A1(n5537), .A2(n5536), .ZN(n5563) );
  INV_X1 U7190 ( .A(n5563), .ZN(n8563) );
  NAND2_X1 U7191 ( .A1(n9231), .A2(n5680), .ZN(n5539) );
  NAND2_X1 U7192 ( .A1(n9104), .A2(n5689), .ZN(n5538) );
  NAND2_X1 U7193 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  XNOR2_X1 U7194 ( .A(n5540), .B(n4278), .ZN(n8465) );
  INV_X1 U7195 ( .A(n8465), .ZN(n8464) );
  INV_X1 U7196 ( .A(SI_23_), .ZN(n5544) );
  NAND2_X1 U7197 ( .A1(n5545), .A2(n5544), .ZN(n5571) );
  INV_X1 U7198 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7199 ( .A1(n5546), .A2(SI_23_), .ZN(n5547) );
  NAND2_X1 U7200 ( .A1(n7361), .A2(n8716), .ZN(n5549) );
  OR2_X1 U7201 ( .A1(n8717), .A2(n10025), .ZN(n5548) );
  NAND2_X1 U7202 ( .A1(n9219), .A2(n5680), .ZN(n5559) );
  INV_X1 U7203 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7204 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  NAND2_X1 U7205 ( .A1(n5578), .A2(n5552), .ZN(n9214) );
  OR2_X1 U7206 ( .A1(n9214), .A2(n5652), .ZN(n5557) );
  INV_X1 U7207 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9213) );
  INV_X1 U7208 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9470) );
  OR2_X1 U7209 ( .A1(n4420), .A2(n9470), .ZN(n5554) );
  INV_X1 U7210 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9401) );
  OR2_X1 U7211 ( .A1(n4271), .A2(n9401), .ZN(n5553) );
  OAI211_X1 U7212 ( .C1(n8624), .C2(n9213), .A(n5554), .B(n5553), .ZN(n5555)
         );
  INV_X1 U7213 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7214 ( .A1(n5557), .A2(n5556), .ZN(n9107) );
  NAND2_X1 U7215 ( .A1(n9107), .A2(n5689), .ZN(n5558) );
  NAND2_X1 U7216 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  XNOR2_X1 U7217 ( .A(n5560), .B(n5658), .ZN(n5566) );
  INV_X1 U7218 ( .A(n5566), .ZN(n8469) );
  NAND2_X1 U7219 ( .A1(n9219), .A2(n5689), .ZN(n5562) );
  NAND2_X1 U7220 ( .A1(n9107), .A2(n4276), .ZN(n5561) );
  NAND2_X1 U7221 ( .A1(n5562), .A2(n5561), .ZN(n8468) );
  NAND2_X1 U7222 ( .A1(n8469), .A2(n8468), .ZN(n8467) );
  OAI21_X1 U7223 ( .B1(n8563), .B2(n8464), .A(n8467), .ZN(n5568) );
  OAI21_X1 U7224 ( .B1(n8465), .B2(n5563), .A(n8468), .ZN(n5565) );
  NOR3_X1 U7225 ( .A1(n8465), .A2(n8468), .A3(n5563), .ZN(n5564) );
  AOI21_X1 U7226 ( .B1(n5566), .B2(n5565), .A(n5564), .ZN(n5567) );
  INV_X1 U7227 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7432) );
  INV_X1 U7228 ( .A(SI_24_), .ZN(n5572) );
  NAND2_X1 U7229 ( .A1(n5573), .A2(n5572), .ZN(n5595) );
  INV_X1 U7230 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7231 ( .A1(n5574), .A2(SI_24_), .ZN(n5575) );
  NAND2_X1 U7232 ( .A1(n7431), .A2(n8716), .ZN(n5577) );
  OR2_X1 U7233 ( .A1(n8717), .A2(n7432), .ZN(n5576) );
  AND2_X1 U7234 ( .A1(n5578), .A2(n8538), .ZN(n5579) );
  OR2_X1 U7235 ( .A1(n5603), .A2(n5579), .ZN(n8539) );
  INV_X1 U7236 ( .A(n8539), .ZN(n9198) );
  NAND2_X1 U7237 ( .A1(n9198), .A2(n5685), .ZN(n5587) );
  INV_X1 U7238 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5584) );
  INV_X1 U7239 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5580) );
  OR2_X1 U7240 ( .A1(n4420), .A2(n5580), .ZN(n5583) );
  INV_X1 U7241 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5581) );
  OR2_X1 U7242 ( .A1(n4272), .A2(n5581), .ZN(n5582) );
  OAI211_X1 U7243 ( .C1(n8624), .C2(n5584), .A(n5583), .B(n5582), .ZN(n5585)
         );
  INV_X1 U7244 ( .A(n5585), .ZN(n5586) );
  AOI22_X1 U7245 ( .A1(n9394), .A2(n5680), .B1(n5661), .B2(n9111), .ZN(n5588)
         );
  XOR2_X1 U7246 ( .A(n4278), .B(n5588), .Z(n5590) );
  OAI22_X1 U7247 ( .A1(n9201), .A2(n5047), .B1(n9110), .B2(n5693), .ZN(n5589)
         );
  NOR2_X1 U7248 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  AOI21_X1 U7249 ( .B1(n5590), .B2(n5589), .A(n5591), .ZN(n8534) );
  INV_X1 U7250 ( .A(n5591), .ZN(n5592) );
  NAND2_X1 U7251 ( .A1(n5594), .A2(n5593), .ZN(n5596) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7477) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U7254 ( .A1(n5598), .A2(n5597), .ZN(n5615) );
  INV_X1 U7255 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U7256 ( .A1(n5599), .A2(SI_25_), .ZN(n5600) );
  XNOR2_X1 U7257 ( .A(n5614), .B(n5613), .ZN(n7467) );
  NAND2_X1 U7258 ( .A1(n7467), .A2(n8716), .ZN(n5602) );
  OR2_X1 U7259 ( .A1(n8717), .A2(n7468), .ZN(n5601) );
  OR2_X1 U7260 ( .A1(n5603), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7261 ( .A1(n5603), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7262 ( .A1(n5604), .A2(n5622), .ZN(n9182) );
  INV_X1 U7263 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9181) );
  INV_X1 U7264 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9466) );
  OR2_X1 U7265 ( .A1(n4420), .A2(n9466), .ZN(n5606) );
  INV_X1 U7266 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9390) );
  OR2_X1 U7267 ( .A1(n4271), .A2(n9390), .ZN(n5605) );
  OAI211_X1 U7268 ( .C1(n5645), .C2(n9181), .A(n5606), .B(n5605), .ZN(n5607)
         );
  INV_X1 U7269 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7270 ( .A1(n5609), .A2(n5608), .ZN(n9113) );
  INV_X1 U7271 ( .A(n9113), .ZN(n9114) );
  OAI22_X1 U7272 ( .A1(n4623), .A2(n5047), .B1(n9114), .B2(n5693), .ZN(n5631)
         );
  NAND2_X1 U7273 ( .A1(n9180), .A2(n5680), .ZN(n5611) );
  NAND2_X1 U7274 ( .A1(n9113), .A2(n5689), .ZN(n5610) );
  NAND2_X1 U7275 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  XNOR2_X1 U7276 ( .A(n5612), .B(n4278), .ZN(n5632) );
  XOR2_X1 U7277 ( .A(n5631), .B(n5632), .Z(n8507) );
  NAND2_X1 U7278 ( .A1(n8506), .A2(n8507), .ZN(n8505) );
  INV_X1 U7279 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10024) );
  INV_X1 U7280 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9998) );
  INV_X1 U7281 ( .A(SI_26_), .ZN(n5616) );
  NAND2_X1 U7282 ( .A1(n5617), .A2(n5616), .ZN(n5636) );
  INV_X1 U7283 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7284 ( .A1(n5618), .A2(SI_26_), .ZN(n5619) );
  NAND2_X1 U7285 ( .A1(n7480), .A2(n8716), .ZN(n5621) );
  OR2_X1 U7286 ( .A1(n8717), .A2(n9998), .ZN(n5620) );
  NAND2_X1 U7287 ( .A1(n9164), .A2(n5680), .ZN(n5627) );
  INV_X1 U7288 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9166) );
  INV_X1 U7289 ( .A(n5622), .ZN(n5623) );
  NAND2_X1 U7290 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n5623), .ZN(n5648) );
  OAI21_X1 U7291 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5623), .A(n5648), .ZN(
        n9165) );
  OAI22_X1 U7292 ( .A1(n8624), .A2(n9166), .B1(n5652), .B2(n9165), .ZN(n5625)
         );
  INV_X1 U7293 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9385) );
  INV_X1 U7294 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9462) );
  OAI22_X1 U7295 ( .A1(n4272), .A2(n9385), .B1(n4420), .B2(n9462), .ZN(n5624)
         );
  NAND2_X1 U7296 ( .A1(n9116), .A2(n5689), .ZN(n5626) );
  NAND2_X1 U7297 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  XNOR2_X1 U7298 ( .A(n5628), .B(n5658), .ZN(n5666) );
  AND2_X1 U7299 ( .A1(n9116), .A2(n4276), .ZN(n5630) );
  AOI21_X1 U7300 ( .B1(n9164), .B2(n5661), .A(n5630), .ZN(n5667) );
  XNOR2_X1 U7301 ( .A(n5666), .B(n5667), .ZN(n8595) );
  NOR2_X1 U7302 ( .A1(n5632), .A2(n5631), .ZN(n8596) );
  NOR2_X1 U7303 ( .A1(n8595), .A2(n8596), .ZN(n5633) );
  NAND2_X1 U7304 ( .A1(n8505), .A2(n5633), .ZN(n8598) );
  INV_X1 U7305 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U7306 ( .A(n8450), .B(n9933), .S(n7521), .Z(n5637) );
  NAND2_X1 U7307 ( .A1(n5637), .A2(n9931), .ZN(n5675) );
  INV_X1 U7308 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7309 ( .A1(n5638), .A2(SI_27_), .ZN(n5639) );
  NAND2_X1 U7310 ( .A1(n8448), .A2(n8716), .ZN(n5641) );
  OR2_X1 U7311 ( .A1(n8717), .A2(n9933), .ZN(n5640) );
  NAND2_X1 U7312 ( .A1(n9379), .A2(n5680), .ZN(n5657) );
  INV_X1 U7313 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5644) );
  INV_X1 U7314 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5642) );
  OR2_X1 U7315 ( .A1(n4272), .A2(n5642), .ZN(n5643) );
  OAI21_X1 U7316 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5646) );
  INV_X1 U7317 ( .A(n5646), .ZN(n5655) );
  INV_X1 U7318 ( .A(n5648), .ZN(n5647) );
  NAND2_X1 U7319 ( .A1(n5647), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5738) );
  INV_X1 U7320 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U7321 ( .A1(n5648), .A2(n7712), .ZN(n5649) );
  NAND2_X1 U7322 ( .A1(n5738), .A2(n5649), .ZN(n7711) );
  INV_X1 U7323 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5650) );
  OR2_X1 U7324 ( .A1(n4420), .A2(n5650), .ZN(n5651) );
  OAI21_X1 U7325 ( .B1(n5652), .B2(n7711), .A(n5651), .ZN(n5653) );
  INV_X1 U7326 ( .A(n5653), .ZN(n5654) );
  OR2_X1 U7327 ( .A1(n9118), .A2(n5047), .ZN(n5656) );
  NAND2_X1 U7328 ( .A1(n5657), .A2(n5656), .ZN(n5659) );
  XNOR2_X1 U7329 ( .A(n5659), .B(n5658), .ZN(n5663) );
  INV_X1 U7330 ( .A(n5663), .ZN(n5665) );
  NOR2_X1 U7331 ( .A1(n9118), .A2(n5693), .ZN(n5660) );
  AOI21_X1 U7332 ( .B1(n9379), .B2(n5661), .A(n5660), .ZN(n5662) );
  INV_X1 U7333 ( .A(n5662), .ZN(n5664) );
  AOI21_X1 U7334 ( .B1(n5665), .B2(n5664), .A(n5721), .ZN(n7707) );
  INV_X1 U7335 ( .A(n7707), .ZN(n5671) );
  INV_X1 U7336 ( .A(n5666), .ZN(n5669) );
  INV_X1 U7337 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U7338 ( .A1(n5669), .A2(n5668), .ZN(n7708) );
  INV_X1 U7339 ( .A(n7708), .ZN(n5670) );
  NOR2_X1 U7340 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U7341 ( .A1(n5674), .A2(n5673), .ZN(n5676) );
  INV_X1 U7342 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5677) );
  INV_X1 U7343 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U7344 ( .A(n6217), .B(SI_28_), .ZN(n6214) );
  NAND2_X1 U7345 ( .A1(n6101), .A2(n8716), .ZN(n5679) );
  OR2_X1 U7346 ( .A1(n8717), .A2(n9519), .ZN(n5678) );
  NAND2_X1 U7347 ( .A1(n9373), .A2(n5680), .ZN(n5691) );
  INV_X1 U7348 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5681) );
  OR2_X1 U7349 ( .A1(n4271), .A2(n5681), .ZN(n5684) );
  INV_X1 U7350 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5682) );
  OR2_X1 U7351 ( .A1(n4420), .A2(n5682), .ZN(n5683) );
  AND2_X1 U7352 ( .A1(n5684), .A2(n5683), .ZN(n5688) );
  XNOR2_X1 U7353 ( .A(n5738), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U7354 ( .A1(n5685), .A2(n9137), .ZN(n5687) );
  NAND2_X1 U7355 ( .A1(n6365), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7356 ( .A1(n9075), .A2(n5689), .ZN(n5690) );
  NAND2_X1 U7357 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  XNOR2_X1 U7358 ( .A(n5692), .B(n4278), .ZN(n5696) );
  NOR2_X1 U7359 ( .A1(n9119), .A2(n5693), .ZN(n5694) );
  AOI21_X1 U7360 ( .B1(n9373), .B2(n5689), .A(n5694), .ZN(n5695) );
  XNOR2_X1 U7361 ( .A(n5696), .B(n5695), .ZN(n5722) );
  NOR2_X1 U7362 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n5700) );
  NOR4_X1 U7363 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5699) );
  NOR4_X1 U7364 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5698) );
  NOR4_X1 U7365 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5697) );
  NAND4_X1 U7366 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n5706)
         );
  NOR4_X1 U7367 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5704) );
  NOR4_X1 U7368 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5703) );
  NOR4_X1 U7369 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5702) );
  NOR4_X1 U7370 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5701) );
  NAND4_X1 U7371 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), .ZN(n5705)
         );
  NOR2_X1 U7372 ( .A1(n5706), .A2(n5705), .ZN(n6564) );
  INV_X1 U7373 ( .A(n5710), .ZN(n7469) );
  NAND2_X1 U7374 ( .A1(n7469), .A2(P1_B_REG_SCAN_IN), .ZN(n5708) );
  MUX2_X1 U7375 ( .A(n5708), .B(P1_B_REG_SCAN_IN), .S(n5707), .Z(n5709) );
  NAND2_X1 U7376 ( .A1(n5709), .A2(n5711), .ZN(n6390) );
  OR2_X1 U7377 ( .A1(n5711), .A2(n5710), .ZN(n9506) );
  OAI21_X1 U7378 ( .B1(n6390), .B2(P1_D_REG_1__SCAN_IN), .A(n9506), .ZN(n6563)
         );
  INV_X1 U7379 ( .A(n6563), .ZN(n6937) );
  INV_X1 U7380 ( .A(n6390), .ZN(n5713) );
  INV_X1 U7381 ( .A(n5707), .ZN(n7433) );
  INV_X1 U7382 ( .A(n5711), .ZN(n7481) );
  OAI211_X1 U7383 ( .C1(n6564), .C2(n6390), .A(n6937), .B(n6594), .ZN(n5737)
         );
  NAND2_X1 U7384 ( .A1(n5714), .A2(n4971), .ZN(n5715) );
  INV_X1 U7385 ( .A(n6565), .ZN(n5718) );
  OR2_X1 U7386 ( .A1(n5737), .A2(n5718), .ZN(n5723) );
  AND2_X1 U7387 ( .A1(n8863), .A2(n5719), .ZN(n6372) );
  INV_X1 U7388 ( .A(n6372), .ZN(n8759) );
  INV_X1 U7389 ( .A(n5719), .ZN(n8771) );
  AND2_X1 U7390 ( .A1(n8759), .A2(n9698), .ZN(n5726) );
  INV_X1 U7391 ( .A(n5726), .ZN(n5720) );
  OR4_X2 U7392 ( .A1(n7709), .A2(n5721), .A3(n5722), .A4(n8615), .ZN(n5753) );
  AND2_X1 U7393 ( .A1(n5722), .A2(n9571), .ZN(n5751) );
  NAND3_X1 U7394 ( .A1(n5722), .A2(n9571), .A3(n5721), .ZN(n5749) );
  INV_X1 U7395 ( .A(n5723), .ZN(n5725) );
  NOR2_X1 U7396 ( .A1(n6576), .A2(n5732), .ZN(n6943) );
  INV_X1 U7397 ( .A(n6562), .ZN(n5724) );
  AOI21_X2 U7398 ( .B1(n5725), .B2(n6943), .A(n9302), .ZN(n9568) );
  NAND2_X1 U7399 ( .A1(n5737), .A2(n5726), .ZN(n5728) );
  INV_X1 U7400 ( .A(n6566), .ZN(n5727) );
  NAND4_X1 U7401 ( .A1(n5728), .A2(n5019), .A3(n6371), .A4(n5727), .ZN(n5729)
         );
  NAND2_X1 U7402 ( .A1(n5729), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5735) );
  OR2_X1 U7403 ( .A1(n6570), .A2(n5730), .ZN(n6569) );
  INV_X1 U7404 ( .A(n6569), .ZN(n5731) );
  NAND2_X1 U7405 ( .A1(n6565), .A2(n5731), .ZN(n8862) );
  OR2_X1 U7406 ( .A1(n5732), .A2(P1_U3086), .ZN(n7097) );
  NAND2_X1 U7407 ( .A1(n8862), .A2(n7097), .ZN(n5733) );
  NAND2_X1 U7408 ( .A1(n5737), .A2(n5733), .ZN(n5734) );
  INV_X1 U7409 ( .A(n9137), .ZN(n5746) );
  NAND2_X1 U7410 ( .A1(n6565), .A2(n8858), .ZN(n5736) );
  INV_X1 U7411 ( .A(n9520), .ZN(n6426) );
  INV_X1 U7412 ( .A(n9074), .ZN(n8508) );
  OR2_X1 U7413 ( .A1(n9118), .A2(n8508), .ZN(n5744) );
  INV_X1 U7414 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9122) );
  INV_X1 U7415 ( .A(n5738), .ZN(n5739) );
  NAND2_X1 U7416 ( .A1(n5739), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9121) );
  OAI22_X1 U7417 ( .A1(n8624), .A2(n9122), .B1(n5652), .B2(n9121), .ZN(n5742)
         );
  INV_X1 U7418 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9366) );
  INV_X1 U7419 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9455) );
  OAI22_X1 U7420 ( .A1(n4271), .A2(n9366), .B1(n4420), .B2(n9455), .ZN(n5741)
         );
  NAND2_X1 U7421 ( .A1(n8868), .A2(n8588), .ZN(n5743) );
  NAND2_X1 U7422 ( .A1(n5744), .A2(n5743), .ZN(n9132) );
  AOI22_X1 U7423 ( .A1(n9566), .A2(n9132), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5745) );
  OAI21_X1 U7424 ( .B1(n9575), .B2(n5746), .A(n5745), .ZN(n5747) );
  AOI21_X1 U7425 ( .B1(n9373), .B2(n8613), .A(n5747), .ZN(n5748) );
  NAND2_X1 U7426 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  AOI21_X1 U7427 ( .B1(n7709), .B2(n5751), .A(n5750), .ZN(n5752) );
  NAND2_X1 U7428 ( .A1(n5753), .A2(n5752), .ZN(P1_U3220) );
  INV_X1 U7429 ( .A(n5879), .ZN(n5755) );
  INV_X1 U7430 ( .A(n5963), .ZN(n5763) );
  NAND2_X1 U7431 ( .A1(n5763), .A2(n5762), .ZN(n6010) );
  XNOR2_X2 U7432 ( .A(n5765), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6259) );
  NOR2_X1 U7433 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5771) );
  NOR2_X1 U7434 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5770) );
  NOR2_X1 U7435 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5769) );
  NOR2_X1 U7436 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5768) );
  NAND4_X1 U7437 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n5774)
         );
  NAND4_X1 U7438 ( .A1(n5772), .A2(n5759), .A3(n5779), .A4(n5972), .ZN(n5773)
         );
  NAND2_X1 U7439 ( .A1(n5784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7440 ( .A1(n6805), .A2(n7333), .ZN(n5781) );
  NAND2_X1 U7441 ( .A1(n5781), .A2(n8065), .ZN(n6159) );
  INV_X1 U7442 ( .A(n6159), .ZN(n5783) );
  NAND2_X1 U7443 ( .A1(n5782), .A2(n8080), .ZN(n7698) );
  INV_X1 U7444 ( .A(n9798), .ZN(n8354) );
  INV_X1 U7445 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5786) );
  XNOR2_X2 U7446 ( .A(n5787), .B(n5786), .ZN(n7717) );
  XNOR2_X2 U7447 ( .A(n5790), .B(n5789), .ZN(n8444) );
  INV_X1 U7448 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6959) );
  AND2_X2 U7449 ( .A1(n7717), .A2(n8444), .ZN(n5837) );
  NAND2_X1 U7450 ( .A1(n5837), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7451 ( .A1(n5792), .A2(n5791), .ZN(n5813) );
  INV_X1 U7452 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7023) );
  OR2_X1 U7453 ( .A1(n5813), .A2(n7023), .ZN(n5793) );
  INV_X1 U7454 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7021) );
  XNOR2_X2 U7455 ( .A(n5798), .B(n5797), .ZN(n6155) );
  NAND2_X1 U7456 ( .A1(n6167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7457 ( .A1(n5799), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5801) );
  NAND2_X2 U7458 ( .A1(n6264), .A2(n6956), .ZN(n7565) );
  INV_X1 U7459 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U7460 ( .A1(n5837), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5811) );
  INV_X1 U7461 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6859) );
  OR2_X1 U7462 ( .A1(n5817), .A2(n6859), .ZN(n5810) );
  INV_X1 U7463 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6649) );
  OR2_X1 U7464 ( .A1(n5838), .A2(n6649), .ZN(n5814) );
  NAND2_X1 U7465 ( .A1(n4412), .A2(SI_0_), .ZN(n5816) );
  XNOR2_X1 U7466 ( .A(n5816), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8452) );
  MUX2_X1 U7467 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8452), .S(n6443), .Z(n6268) );
  NAND2_X1 U7468 ( .A1(n6822), .A2(n6268), .ZN(n7560) );
  NAND2_X1 U7469 ( .A1(n5818), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5824) );
  NOR2_X1 U7470 ( .A1(n4932), .A2(n5820), .ZN(n5823) );
  NAND2_X1 U7471 ( .A1(n5821), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5822) );
  OR2_X1 U7472 ( .A1(n7526), .A2(n6342), .ZN(n5829) );
  OR2_X1 U7473 ( .A1(n5845), .A2(n6341), .ZN(n5828) );
  XNOR2_X2 U7474 ( .A(n5826), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U7475 ( .A1(n6020), .A2(n6530), .ZN(n5827) );
  INV_X1 U7476 ( .A(n6807), .ZN(n5830) );
  NAND2_X1 U7477 ( .A1(n5831), .A2(n5830), .ZN(n5834) );
  NAND2_X1 U7478 ( .A1(n9744), .A2(n6807), .ZN(n7569) );
  NAND2_X1 U7479 ( .A1(n6806), .A2(n5833), .ZN(n5835) );
  BUF_X4 U7480 ( .A(n5837), .Z(n7532) );
  NAND2_X1 U7481 ( .A1(n7532), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5841) );
  OR2_X1 U7482 ( .A1(n5838), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7483 ( .A1(n5818), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7484 ( .A1(n5804), .A2(n5842), .ZN(n5856) );
  NAND2_X1 U7485 ( .A1(n5856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5844) );
  INV_X1 U7486 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U7487 ( .A(n5844), .B(n5843), .ZN(n6561) );
  OR2_X1 U7488 ( .A1(n4418), .A2(n6340), .ZN(n5847) );
  OR2_X1 U7489 ( .A1(n7526), .A2(n6339), .ZN(n5846) );
  NAND2_X1 U7490 ( .A1(n5819), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5855) );
  INV_X1 U7491 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7492 ( .A1(n6226), .A2(n5849), .ZN(n5854) );
  NOR2_X1 U7493 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5861) );
  AND2_X1 U7494 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5850) );
  NOR2_X1 U7495 ( .A1(n5861), .A2(n5850), .ZN(n7862) );
  OR2_X1 U7496 ( .A1(n5838), .A2(n7862), .ZN(n5853) );
  INV_X1 U7497 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7498 ( .A1(n5817), .A2(n5851), .ZN(n5852) );
  OR2_X1 U7499 ( .A1(n5856), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7500 ( .A1(n5867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  INV_X1 U7501 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7502 ( .A1(n4418), .A2(n6346), .ZN(n5860) );
  OR2_X1 U7503 ( .A1(n7526), .A2(n6345), .ZN(n5859) );
  OAI211_X1 U7504 ( .C1(n6443), .C2(n6635), .A(n5860), .B(n5859), .ZN(n7861)
         );
  NAND2_X1 U7505 ( .A1(n6982), .A2(n7861), .ZN(n7575) );
  INV_X1 U7506 ( .A(n7861), .ZN(n9766) );
  NAND2_X1 U7507 ( .A1(n9746), .A2(n9766), .ZN(n7586) );
  NAND2_X1 U7508 ( .A1(n7532), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5866) );
  INV_X1 U7509 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7091) );
  OR2_X1 U7510 ( .A1(n5817), .A2(n7091), .ZN(n5865) );
  NAND2_X1 U7511 ( .A1(n5861), .A2(n6638), .ZN(n5873) );
  OR2_X1 U7512 ( .A1(n5861), .A2(n6638), .ZN(n5862) );
  AND2_X1 U7513 ( .A1(n5873), .A2(n5862), .ZN(n7092) );
  OR2_X1 U7514 ( .A1(n5838), .A2(n7092), .ZN(n5864) );
  NAND2_X1 U7515 ( .A1(n5819), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5863) );
  NAND4_X1 U7516 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n7956)
         );
  INV_X1 U7517 ( .A(n7956), .ZN(n7102) );
  OAI21_X1 U7518 ( .B1(n5867), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5869) );
  INV_X1 U7519 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5868) );
  XNOR2_X1 U7520 ( .A(n5869), .B(n5868), .ZN(n6698) );
  OR2_X1 U7521 ( .A1(n4418), .A2(n6349), .ZN(n5871) );
  OR2_X1 U7522 ( .A1(n7526), .A2(n6348), .ZN(n5870) );
  OAI211_X1 U7523 ( .C1(n6443), .C2(n6698), .A(n5871), .B(n5870), .ZN(n7094)
         );
  NAND2_X1 U7524 ( .A1(n7102), .A2(n7094), .ZN(n7589) );
  NAND2_X1 U7525 ( .A1(n7956), .A2(n9772), .ZN(n7585) );
  NAND2_X1 U7526 ( .A1(n5819), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5878) );
  INV_X1 U7527 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7528 ( .A1(n6226), .A2(n5872), .ZN(n5877) );
  NAND2_X1 U7529 ( .A1(n5873), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5874) );
  AND2_X1 U7530 ( .A1(n5884), .A2(n5874), .ZN(n7243) );
  OR2_X1 U7531 ( .A1(n5838), .A2(n7243), .ZN(n5876) );
  INV_X1 U7532 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7242) );
  OR2_X1 U7533 ( .A1(n5817), .A2(n7242), .ZN(n5875) );
  NAND2_X1 U7534 ( .A1(n5879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7535 ( .A(n5880), .B(n5754), .ZN(n9871) );
  OR2_X1 U7536 ( .A1(n4418), .A2(n6351), .ZN(n5882) );
  OR2_X1 U7537 ( .A1(n7526), .A2(n6350), .ZN(n5881) );
  OAI211_X1 U7538 ( .C1(n6443), .C2(n9871), .A(n5882), .B(n5881), .ZN(n7245)
         );
  NAND2_X1 U7539 ( .A1(n6263), .A2(n7245), .ZN(n7590) );
  INV_X1 U7540 ( .A(n7245), .ZN(n9776) );
  NAND2_X1 U7541 ( .A1(n7955), .A2(n9776), .ZN(n7592) );
  NAND2_X1 U7542 ( .A1(n7590), .A2(n7592), .ZN(n7504) );
  INV_X1 U7543 ( .A(n7504), .ZN(n7239) );
  NAND2_X1 U7544 ( .A1(n7532), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5889) );
  INV_X1 U7545 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6748) );
  OR2_X1 U7546 ( .A1(n7530), .A2(n6748), .ZN(n5888) );
  AND2_X1 U7547 ( .A1(n5884), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5885) );
  NOR2_X1 U7548 ( .A1(n5899), .A2(n5885), .ZN(n7293) );
  OR2_X1 U7549 ( .A1(n5838), .A2(n7293), .ZN(n5887) );
  INV_X1 U7550 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6704) );
  OR2_X1 U7551 ( .A1(n5817), .A2(n6704), .ZN(n5886) );
  NAND2_X1 U7552 ( .A1(n5891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U7553 ( .A(n5892), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7554 ( .A1(n6102), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6020), .B2(
        n6747), .ZN(n5894) );
  NAND2_X1 U7555 ( .A1(n6353), .A2(n7525), .ZN(n5893) );
  NAND2_X1 U7556 ( .A1(n5894), .A2(n5893), .ZN(n7195) );
  NAND2_X1 U7557 ( .A1(n6322), .A2(n7195), .ZN(n7595) );
  INV_X1 U7558 ( .A(n7195), .ZN(n9780) );
  NAND2_X1 U7559 ( .A1(n9729), .A2(n9780), .ZN(n9734) );
  NAND2_X1 U7560 ( .A1(n7595), .A2(n9734), .ZN(n7581) );
  NAND2_X1 U7561 ( .A1(n6359), .A2(n7525), .ZN(n5898) );
  OR2_X1 U7562 ( .A1(n5895), .A2(n8441), .ZN(n5896) );
  XNOR2_X1 U7563 ( .A(n5896), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7564 ( .A1(n6102), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6020), .B2(
        n6766), .ZN(n5897) );
  NAND2_X1 U7565 ( .A1(n5898), .A2(n5897), .ZN(n9738) );
  NAND2_X1 U7566 ( .A1(n7532), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7567 ( .A1(n5818), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5903) );
  INV_X1 U7568 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6764) );
  OR2_X1 U7569 ( .A1(n7530), .A2(n6764), .ZN(n5902) );
  NOR2_X1 U7570 ( .A1(n5899), .A2(n6757), .ZN(n5900) );
  OR2_X1 U7571 ( .A1(n5912), .A2(n5900), .ZN(n9740) );
  NAND2_X1 U7572 ( .A1(n5821), .A2(n9740), .ZN(n5901) );
  NAND4_X1 U7573 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n7954)
         );
  NAND2_X1 U7574 ( .A1(n9789), .A2(n7954), .ZN(n7600) );
  INV_X1 U7575 ( .A(n7954), .ZN(n7371) );
  NAND2_X1 U7576 ( .A1(n7371), .A2(n9738), .ZN(n7596) );
  NAND2_X1 U7577 ( .A1(n6388), .A2(n7525), .ZN(n5909) );
  INV_X1 U7578 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8441) );
  NOR2_X1 U7579 ( .A1(n5776), .A2(n8441), .ZN(n5906) );
  MUX2_X1 U7580 ( .A(n8441), .B(n5906), .S(P2_IR_REG_9__SCAN_IN), .Z(n5907) );
  NOR2_X1 U7581 ( .A1(n5907), .A2(n5928), .ZN(n6850) );
  AOI22_X1 U7582 ( .A1(n6102), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6020), .B2(
        n6850), .ZN(n5908) );
  NAND2_X1 U7583 ( .A1(n5909), .A2(n5908), .ZN(n7378) );
  NAND2_X1 U7584 ( .A1(n5819), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5917) );
  INV_X1 U7585 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7586 ( .A1(n6226), .A2(n5910), .ZN(n5916) );
  NAND2_X1 U7587 ( .A1(n5912), .A2(n5911), .ZN(n5921) );
  OR2_X1 U7588 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  AND2_X1 U7589 ( .A1(n5921), .A2(n5913), .ZN(n7376) );
  OR2_X1 U7590 ( .A1(n5838), .A2(n7376), .ZN(n5915) );
  INV_X1 U7591 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6835) );
  OR2_X1 U7592 ( .A1(n5817), .A2(n6835), .ZN(n5914) );
  NAND2_X1 U7593 ( .A1(n7378), .A2(n7424), .ZN(n7597) );
  NAND2_X1 U7594 ( .A1(n6393), .A2(n7525), .ZN(n5920) );
  OR2_X1 U7595 ( .A1(n5928), .A2(n8441), .ZN(n5918) );
  XNOR2_X1 U7596 ( .A(n5918), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7079) );
  AOI22_X1 U7597 ( .A1(n6102), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6020), .B2(
        n7079), .ZN(n5919) );
  NAND2_X1 U7598 ( .A1(n7532), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5926) );
  INV_X1 U7599 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7040) );
  OR2_X1 U7600 ( .A1(n7530), .A2(n7040), .ZN(n5925) );
  NAND2_X1 U7601 ( .A1(n5921), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5922) );
  AND2_X1 U7602 ( .A1(n5931), .A2(n5922), .ZN(n7460) );
  OR2_X1 U7603 ( .A1(n5838), .A2(n7460), .ZN(n5924) );
  INV_X1 U7604 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7041) );
  OR2_X1 U7605 ( .A1(n5817), .A2(n7041), .ZN(n5923) );
  OR2_X1 U7606 ( .A1(n9802), .A2(n7473), .ZN(n7608) );
  AND2_X1 U7607 ( .A1(n7608), .A2(n7579), .ZN(n7604) );
  NAND2_X1 U7608 ( .A1(n9802), .A2(n7473), .ZN(n7609) );
  NAND2_X1 U7609 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7610 ( .A1(n5929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5939) );
  XNOR2_X1 U7611 ( .A(n5939), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7208) );
  AOI22_X1 U7612 ( .A1(n6102), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6020), .B2(
        n7208), .ZN(n5930) );
  NAND2_X1 U7613 ( .A1(n7532), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5936) );
  INV_X1 U7614 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7069) );
  OR2_X1 U7615 ( .A1(n7530), .A2(n7069), .ZN(n5935) );
  NAND2_X1 U7616 ( .A1(n5931), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5932) );
  AND2_X1 U7617 ( .A1(n5944), .A2(n5932), .ZN(n7902) );
  OR2_X1 U7618 ( .A1(n5838), .A2(n7902), .ZN(n5934) );
  INV_X1 U7619 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7070) );
  OR2_X1 U7620 ( .A1(n5817), .A2(n7070), .ZN(n5933) );
  XNOR2_X1 U7621 ( .A(n9808), .B(n7952), .ZN(n7470) );
  NAND2_X1 U7622 ( .A1(n9808), .A2(n8287), .ZN(n7552) );
  NAND2_X1 U7623 ( .A1(n6448), .A2(n7525), .ZN(n5943) );
  NAND2_X1 U7624 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U7625 ( .A1(n5940), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5941) );
  INV_X1 U7626 ( .A(n7383), .ZN(n7215) );
  AOI22_X1 U7627 ( .A1(n6102), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6020), .B2(
        n7215), .ZN(n5942) );
  NAND2_X1 U7628 ( .A1(n5943), .A2(n5942), .ZN(n9815) );
  INV_X1 U7629 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7227) );
  OR2_X1 U7630 ( .A1(n7530), .A2(n7227), .ZN(n5949) );
  AND2_X1 U7631 ( .A1(n5944), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U7632 ( .A1(n5956), .A2(n5945), .ZN(n8289) );
  OR2_X1 U7633 ( .A1(n5838), .A2(n8289), .ZN(n5948) );
  INV_X1 U7634 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8290) );
  OR2_X1 U7635 ( .A1(n5817), .A2(n8290), .ZN(n5947) );
  NAND2_X1 U7636 ( .A1(n7532), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5946) );
  NAND4_X1 U7637 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n7951)
         );
  OR2_X1 U7638 ( .A1(n9815), .A2(n9547), .ZN(n7554) );
  NAND2_X1 U7639 ( .A1(n9815), .A2(n9547), .ZN(n7555) );
  NAND2_X1 U7640 ( .A1(n7554), .A2(n7555), .ZN(n8293) );
  INV_X1 U7641 ( .A(n8293), .ZN(n5950) );
  NAND2_X1 U7642 ( .A1(n6455), .A2(n7525), .ZN(n5954) );
  NAND2_X1 U7643 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7644 ( .A(n5952), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7960) );
  AOI22_X1 U7645 ( .A1(n6102), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6020), .B2(
        n7960), .ZN(n5953) );
  NAND2_X1 U7646 ( .A1(n5954), .A2(n5953), .ZN(n9538) );
  NAND2_X1 U7647 ( .A1(n7532), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5961) );
  OR2_X1 U7648 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7649 ( .A1(n5956), .A2(n5955), .ZN(n5966) );
  AND2_X1 U7650 ( .A1(n5957), .A2(n5966), .ZN(n9541) );
  OR2_X1 U7651 ( .A1(n5838), .A2(n9541), .ZN(n5960) );
  INV_X1 U7652 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7388) );
  OR2_X1 U7653 ( .A1(n7530), .A2(n7388), .ZN(n5959) );
  NAND2_X1 U7654 ( .A1(n5818), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5958) );
  NAND4_X1 U7655 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n8275)
         );
  NAND2_X1 U7656 ( .A1(n9538), .A2(n8288), .ZN(n7617) );
  NAND2_X1 U7657 ( .A1(n9537), .A2(n7617), .ZN(n5962) );
  OR2_X1 U7658 ( .A1(n9538), .A2(n8288), .ZN(n7618) );
  NAND2_X1 U7659 ( .A1(n6512), .A2(n7525), .ZN(n5965) );
  NAND2_X1 U7660 ( .A1(n5963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7661 ( .A(n5985), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7975) );
  AOI22_X1 U7662 ( .A1(n6102), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6020), .B2(
        n7975), .ZN(n5964) );
  INV_X1 U7663 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8348) );
  OR2_X1 U7664 ( .A1(n7530), .A2(n8348), .ZN(n5971) );
  NAND2_X1 U7665 ( .A1(n5966), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5967) );
  AND2_X1 U7666 ( .A1(n5977), .A2(n5967), .ZN(n8277) );
  OR2_X1 U7667 ( .A1(n5838), .A2(n8277), .ZN(n5970) );
  INV_X1 U7668 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7974) );
  OR2_X1 U7669 ( .A1(n5817), .A2(n7974), .ZN(n5969) );
  NAND2_X1 U7670 ( .A1(n7532), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5968) );
  NAND4_X1 U7671 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n8266)
         );
  NOR2_X1 U7672 ( .A1(n8435), .A2(n9549), .ZN(n7621) );
  NAND2_X1 U7673 ( .A1(n8435), .A2(n9549), .ZN(n7498) );
  NAND2_X1 U7674 ( .A1(n6626), .A2(n7525), .ZN(n5976) );
  NAND2_X1 U7675 ( .A1(n5985), .A2(n5972), .ZN(n5973) );
  NAND2_X1 U7676 ( .A1(n5973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7677 ( .A(n5974), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8006) );
  AOI22_X1 U7678 ( .A1(n6102), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6020), .B2(
        n8006), .ZN(n5975) );
  NAND2_X1 U7679 ( .A1(n5976), .A2(n5975), .ZN(n8429) );
  NAND2_X1 U7680 ( .A1(n7532), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5982) );
  INV_X1 U7681 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8345) );
  OR2_X1 U7682 ( .A1(n7530), .A2(n8345), .ZN(n5981) );
  AND2_X1 U7683 ( .A1(n5977), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U7684 ( .A1(n5989), .A2(n5978), .ZN(n7938) );
  OR2_X1 U7685 ( .A1(n5813), .A2(n7938), .ZN(n5980) );
  INV_X1 U7686 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10021) );
  OR2_X1 U7687 ( .A1(n5817), .A2(n10021), .ZN(n5979) );
  NAND2_X1 U7688 ( .A1(n8429), .A2(n8253), .ZN(n7626) );
  INV_X1 U7689 ( .A(n7626), .ZN(n5983) );
  OR2_X1 U7690 ( .A1(n8429), .A2(n8253), .ZN(n7625) );
  NAND2_X1 U7691 ( .A1(n6686), .A2(n7525), .ZN(n5988) );
  OAI21_X1 U7692 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7693 ( .A1(n5985), .A2(n5984), .ZN(n5997) );
  XNOR2_X1 U7694 ( .A(n5997), .B(n5986), .ZN(n8033) );
  AOI22_X1 U7695 ( .A1(n6102), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6020), .B2(
        n8033), .ZN(n5987) );
  NAND2_X1 U7696 ( .A1(n7532), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5995) );
  INV_X1 U7697 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8341) );
  OR2_X1 U7698 ( .A1(n7530), .A2(n8341), .ZN(n5994) );
  NOR2_X1 U7699 ( .A1(n5989), .A2(n7831), .ZN(n5990) );
  OR2_X1 U7700 ( .A1(n6002), .A2(n5990), .ZN(n8259) );
  INV_X1 U7701 ( .A(n8259), .ZN(n5991) );
  OR2_X1 U7702 ( .A1(n5838), .A2(n5991), .ZN(n5993) );
  INV_X1 U7703 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8258) );
  OR2_X1 U7704 ( .A1(n5817), .A2(n8258), .ZN(n5992) );
  NAND2_X1 U7705 ( .A1(n8422), .A2(n8242), .ZN(n7630) );
  NAND2_X1 U7706 ( .A1(n5996), .A2(n7629), .ZN(n8238) );
  INV_X1 U7707 ( .A(n8238), .ZN(n6009) );
  NAND2_X1 U7708 ( .A1(n6828), .A2(n7525), .ZN(n6000) );
  OAI21_X1 U7709 ( .B1(n5997), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7710 ( .A(n5998), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U7711 ( .A1(n6102), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6020), .B2(
        n9714), .ZN(n5999) );
  OR2_X1 U7712 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  NAND2_X1 U7713 ( .A1(n6014), .A2(n6003), .ZN(n8244) );
  NAND2_X1 U7714 ( .A1(n5821), .A2(n8244), .ZN(n6007) );
  INV_X1 U7715 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9930) );
  OR2_X1 U7716 ( .A1(n7530), .A2(n9930), .ZN(n6006) );
  INV_X1 U7717 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8417) );
  OR2_X1 U7718 ( .A1(n6226), .A2(n8417), .ZN(n6005) );
  INV_X1 U7719 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8246) );
  OR2_X1 U7720 ( .A1(n5817), .A2(n8246), .ZN(n6004) );
  OR2_X1 U7721 ( .A1(n8339), .A2(n8254), .ZN(n7638) );
  NAND2_X1 U7722 ( .A1(n8339), .A2(n8254), .ZN(n8223) );
  NAND2_X1 U7723 ( .A1(n7638), .A2(n8223), .ZN(n8239) );
  INV_X1 U7724 ( .A(n8239), .ZN(n6008) );
  NAND2_X1 U7725 ( .A1(n6862), .A2(n7525), .ZN(n6013) );
  NAND2_X1 U7726 ( .A1(n6010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U7727 ( .A(n6011), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8072) );
  AOI22_X1 U7728 ( .A1(n6102), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6020), .B2(
        n8072), .ZN(n6012) );
  NAND2_X1 U7729 ( .A1(n6014), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7730 ( .A1(n6023), .A2(n6015), .ZN(n8232) );
  NAND2_X1 U7731 ( .A1(n5821), .A2(n8232), .ZN(n6019) );
  INV_X1 U7732 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8335) );
  OR2_X1 U7733 ( .A1(n7530), .A2(n8335), .ZN(n6018) );
  INV_X1 U7734 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8411) );
  OR2_X1 U7735 ( .A1(n6226), .A2(n8411), .ZN(n6017) );
  INV_X1 U7736 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8231) );
  OR2_X1 U7737 ( .A1(n5817), .A2(n8231), .ZN(n6016) );
  NAND2_X1 U7738 ( .A1(n8412), .A2(n8243), .ZN(n7640) );
  AND2_X1 U7739 ( .A1(n7640), .A2(n8223), .ZN(n7636) );
  NAND2_X1 U7740 ( .A1(n7012), .A2(n7525), .ZN(n6022) );
  AOI22_X1 U7741 ( .A1(n6102), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8080), .B2(
        n6020), .ZN(n6021) );
  AND2_X1 U7742 ( .A1(n6023), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6024) );
  OR2_X1 U7743 ( .A1(n6024), .A2(n6033), .ZN(n8217) );
  NAND2_X1 U7744 ( .A1(n8217), .A2(n5821), .ZN(n6029) );
  NAND2_X1 U7745 ( .A1(n5819), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7746 ( .A1(n7532), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6025) );
  AND2_X1 U7747 ( .A1(n6026), .A2(n6025), .ZN(n6028) );
  NAND2_X1 U7748 ( .A1(n5818), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7749 ( .A1(n8330), .A2(n7915), .ZN(n7644) );
  NAND2_X1 U7750 ( .A1(n7110), .A2(n7525), .ZN(n6031) );
  NAND2_X1 U7751 ( .A1(n6102), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6030) );
  INV_X1 U7752 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6032) );
  NOR2_X1 U7753 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  OR2_X1 U7754 ( .A1(n6042), .A2(n6034), .ZN(n8208) );
  NAND2_X1 U7755 ( .A1(n8208), .A2(n5821), .ZN(n6037) );
  AOI22_X1 U7756 ( .A1(n5819), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7532), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7757 ( .A1(n5818), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6035) );
  OR2_X1 U7758 ( .A1(n8405), .A2(n8211), .ZN(n7645) );
  AND2_X1 U7759 ( .A1(n7645), .A2(n8198), .ZN(n7643) );
  NAND2_X1 U7760 ( .A1(n6038), .A2(n7525), .ZN(n6040) );
  NAND2_X1 U7761 ( .A1(n6102), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6039) );
  INV_X1 U7762 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6041) );
  OR2_X1 U7763 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND2_X1 U7764 ( .A1(n6050), .A2(n6043), .ZN(n8194) );
  NAND2_X1 U7765 ( .A1(n8194), .A2(n5821), .ZN(n6046) );
  AOI22_X1 U7766 ( .A1(n7532), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5818), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7767 ( .A1(n5819), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7768 ( .A1(n8399), .A2(n7892), .ZN(n6136) );
  NAND2_X1 U7769 ( .A1(n8405), .A2(n8211), .ZN(n8184) );
  AND2_X1 U7770 ( .A1(n6136), .A2(n8184), .ZN(n7648) );
  NAND2_X1 U7771 ( .A1(n8185), .A2(n7648), .ZN(n6047) );
  NAND2_X1 U7772 ( .A1(n7330), .A2(n7525), .ZN(n6049) );
  NAND2_X1 U7773 ( .A1(n6102), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7774 ( .A1(n6050), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7775 ( .A1(n6057), .A2(n6051), .ZN(n8180) );
  INV_X1 U7776 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U7777 ( .A1(n5819), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7778 ( .A1(n7532), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6052) );
  OAI211_X1 U7779 ( .C1(n9960), .C2(n5817), .A(n6053), .B(n6052), .ZN(n6054)
         );
  AOI21_X1 U7780 ( .B1(n8180), .B2(n5821), .A(n6054), .ZN(n7767) );
  NAND2_X1 U7781 ( .A1(n8394), .A2(n7767), .ZN(n7654) );
  NAND2_X1 U7782 ( .A1(n7653), .A2(n7654), .ZN(n8171) );
  INV_X1 U7783 ( .A(n8171), .ZN(n8176) );
  NAND2_X1 U7784 ( .A1(n7361), .A2(n7525), .ZN(n6056) );
  OR2_X1 U7785 ( .A1(n7526), .A2(n10005), .ZN(n6055) );
  INV_X1 U7786 ( .A(n8388), .ZN(n6142) );
  NAND2_X1 U7787 ( .A1(n6057), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7788 ( .A1(n6058), .A2(n4304), .ZN(n8167) );
  NAND2_X1 U7789 ( .A1(n8167), .A2(n5821), .ZN(n6063) );
  INV_X1 U7790 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U7791 ( .A1(n5818), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7792 ( .A1(n7532), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7793 ( .C1(n7530), .C2(n8317), .A(n6060), .B(n6059), .ZN(n6061)
         );
  INV_X1 U7794 ( .A(n6061), .ZN(n6062) );
  NAND2_X1 U7795 ( .A1(n7431), .A2(n7525), .ZN(n6066) );
  OR2_X1 U7796 ( .A1(n7526), .A2(n10010), .ZN(n6065) );
  NAND2_X1 U7797 ( .A1(n7532), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7798 ( .A1(n5818), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6069) );
  AOI21_X1 U7799 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n4304), .A(n6075), .ZN(
        n8151) );
  OR2_X1 U7800 ( .A1(n5838), .A2(n8151), .ZN(n6068) );
  NAND2_X1 U7801 ( .A1(n5819), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7802 ( .A1(n8382), .A2(n7847), .ZN(n7659) );
  NAND2_X1 U7803 ( .A1(n8388), .A2(n7766), .ZN(n8155) );
  AND2_X1 U7804 ( .A1(n7659), .A2(n8155), .ZN(n7661) );
  NAND2_X1 U7805 ( .A1(n8156), .A2(n7661), .ZN(n6071) );
  NAND2_X1 U7806 ( .A1(n7467), .A2(n7525), .ZN(n6073) );
  NAND2_X1 U7807 ( .A1(n6102), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7808 ( .A1(n5819), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6082) );
  INV_X1 U7809 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8374) );
  OR2_X1 U7810 ( .A1(n6226), .A2(n8374), .ZN(n6081) );
  INV_X1 U7811 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7812 ( .A1(n6074), .A2(n6075), .ZN(n6088) );
  INV_X1 U7813 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7814 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n6076), .ZN(n6077) );
  AND2_X1 U7815 ( .A1(n6088), .A2(n6077), .ZN(n8141) );
  OR2_X1 U7816 ( .A1(n5838), .A2(n8141), .ZN(n6080) );
  INV_X1 U7817 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7818 ( .A1(n5817), .A2(n6078), .ZN(n6079) );
  NAND2_X1 U7819 ( .A1(n7825), .A2(n7851), .ZN(n7666) );
  NAND2_X1 U7820 ( .A1(n8145), .A2(n8138), .ZN(n6083) );
  NAND2_X1 U7821 ( .A1(n7480), .A2(n7525), .ZN(n6085) );
  OR2_X1 U7822 ( .A1(n7526), .A2(n10024), .ZN(n6084) );
  NAND2_X1 U7823 ( .A1(n7532), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6093) );
  INV_X1 U7824 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8128) );
  OR2_X1 U7825 ( .A1(n5817), .A2(n8128), .ZN(n6092) );
  INV_X1 U7826 ( .A(n6088), .ZN(n6087) );
  INV_X1 U7827 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7828 ( .A1(n6087), .A2(n6086), .ZN(n6095) );
  NAND2_X1 U7829 ( .A1(n6088), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6089) );
  AND2_X1 U7830 ( .A1(n6095), .A2(n6089), .ZN(n8129) );
  OR2_X1 U7831 ( .A1(n5813), .A2(n8129), .ZN(n6091) );
  INV_X1 U7832 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8307) );
  OR2_X1 U7833 ( .A1(n7530), .A2(n8307), .ZN(n6090) );
  NOR2_X1 U7834 ( .A1(n8131), .A2(n7751), .ZN(n7549) );
  NAND2_X1 U7835 ( .A1(n8131), .A2(n7751), .ZN(n7496) );
  NAND2_X1 U7836 ( .A1(n6102), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7837 ( .A1(n5819), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7838 ( .A1(n7532), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6099) );
  OR2_X2 U7839 ( .A1(n6095), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7840 ( .A1(n6095), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7841 ( .A1(n5818), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6097) );
  INV_X1 U7842 ( .A(n8126), .ZN(n7790) );
  AND2_X1 U7843 ( .A1(n8119), .A2(n7790), .ZN(n7669) );
  NAND2_X1 U7844 ( .A1(n6101), .A2(n7525), .ZN(n6104) );
  NAND2_X1 U7845 ( .A1(n6102), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7846 ( .A1(n5819), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6113) );
  INV_X1 U7847 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6105) );
  OR2_X1 U7848 ( .A1(n6226), .A2(n6105), .ZN(n6112) );
  INV_X1 U7849 ( .A(n6108), .ZN(n6107) );
  INV_X1 U7850 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7851 ( .A1(n6107), .A2(n6106), .ZN(n8087) );
  NAND2_X1 U7852 ( .A1(n6108), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7853 ( .A1(n5813), .A2(n8106), .ZN(n6111) );
  INV_X1 U7854 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8107) );
  OR2_X1 U7855 ( .A1(n5817), .A2(n8107), .ZN(n6110) );
  XNOR2_X1 U7856 ( .A(n6224), .B(n7795), .ZN(n8108) );
  NAND2_X1 U7857 ( .A1(n7958), .A2(n6268), .ZN(n6951) );
  NOR2_X1 U7858 ( .A1(n5809), .A2(n6956), .ZN(n6114) );
  INV_X1 U7859 ( .A(n6808), .ZN(n6116) );
  NAND2_X1 U7860 ( .A1(n6116), .A2(n5832), .ZN(n6117) );
  NAND2_X1 U7861 ( .A1(n6117), .A2(n4351), .ZN(n9742) );
  NOR2_X1 U7862 ( .A1(n7957), .A2(n9751), .ZN(n6118) );
  AND2_X1 U7863 ( .A1(n6982), .A2(n9766), .ZN(n6119) );
  INV_X1 U7864 ( .A(n7089), .ZN(n6121) );
  INV_X1 U7865 ( .A(n7378), .ZN(n9794) );
  NAND2_X1 U7866 ( .A1(n9794), .A2(n7424), .ZN(n7421) );
  INV_X1 U7867 ( .A(n7473), .ZN(n7953) );
  INV_X1 U7868 ( .A(n9815), .ZN(n6123) );
  OR2_X1 U7869 ( .A1(n9538), .A2(n8275), .ZN(n7500) );
  NAND2_X1 U7870 ( .A1(n9544), .A2(n7500), .ZN(n6124) );
  NAND2_X1 U7871 ( .A1(n9538), .A2(n8275), .ZN(n7499) );
  NAND2_X1 U7872 ( .A1(n6124), .A2(n7499), .ZN(n8274) );
  NAND2_X1 U7873 ( .A1(n8274), .A2(n6126), .ZN(n6128) );
  NAND2_X1 U7874 ( .A1(n8435), .A2(n8266), .ZN(n6127) );
  INV_X1 U7875 ( .A(n8429), .ZN(n7948) );
  NAND2_X1 U7876 ( .A1(n7948), .A2(n8253), .ZN(n6129) );
  NAND2_X1 U7877 ( .A1(n8422), .A2(n8265), .ZN(n6132) );
  NAND2_X1 U7878 ( .A1(n8256), .A2(n6132), .ZN(n8240) );
  AOI21_X1 U7879 ( .B1(n8240), .B2(n8239), .A(n4369), .ZN(n8227) );
  INV_X1 U7880 ( .A(n8412), .ZN(n7919) );
  NAND2_X1 U7881 ( .A1(n7919), .A2(n8243), .ZN(n6134) );
  AND2_X1 U7882 ( .A1(n8330), .A2(n8229), .ZN(n8202) );
  NOR2_X1 U7883 ( .A1(n8201), .A2(n8202), .ZN(n6135) );
  INV_X1 U7884 ( .A(n8405), .ZN(n7875) );
  NAND2_X1 U7885 ( .A1(n7875), .A2(n8211), .ZN(n8188) );
  NAND2_X1 U7886 ( .A1(n8203), .A2(n8188), .ZN(n6137) );
  NAND2_X1 U7887 ( .A1(n7650), .A2(n6136), .ZN(n8187) );
  NAND2_X1 U7888 ( .A1(n6137), .A2(n8187), .ZN(n8174) );
  INV_X1 U7889 ( .A(n8399), .ZN(n6138) );
  NAND2_X1 U7890 ( .A1(n6138), .A2(n7892), .ZN(n8175) );
  NAND2_X1 U7891 ( .A1(n8174), .A2(n8175), .ZN(n6139) );
  NAND2_X1 U7892 ( .A1(n6139), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U7893 ( .A1(n7898), .A2(n7767), .ZN(n6140) );
  NAND2_X1 U7894 ( .A1(n8173), .A2(n6140), .ZN(n8163) );
  NAND2_X1 U7895 ( .A1(n8388), .A2(n8178), .ZN(n6141) );
  NAND2_X1 U7896 ( .A1(n6142), .A2(n7766), .ZN(n6143) );
  NOR2_X1 U7897 ( .A1(n8382), .A2(n8164), .ZN(n8135) );
  AND2_X1 U7898 ( .A1(n8379), .A2(n7851), .ZN(n6147) );
  OR2_X1 U7899 ( .A1(n8135), .A2(n6147), .ZN(n6149) );
  OR2_X1 U7900 ( .A1(n8379), .A2(n7851), .ZN(n6145) );
  NAND2_X1 U7901 ( .A1(n8382), .A2(n8164), .ZN(n8136) );
  AND2_X1 U7902 ( .A1(n6145), .A2(n8136), .ZN(n6146) );
  XNOR2_X1 U7903 ( .A(n6213), .B(n7795), .ZN(n6158) );
  INV_X1 U7904 ( .A(n5782), .ZN(n6260) );
  NAND2_X1 U7905 ( .A1(n6259), .A2(n6260), .ZN(n6150) );
  NAND2_X1 U7906 ( .A1(n8080), .A2(n7704), .ZN(n6202) );
  INV_X1 U7907 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6151) );
  OR2_X1 U7908 ( .A1(n6226), .A2(n6151), .ZN(n6154) );
  INV_X1 U7909 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8099) );
  OR2_X1 U7910 ( .A1(n5817), .A2(n8099), .ZN(n6153) );
  OR2_X1 U7911 ( .A1(n7530), .A2(n6242), .ZN(n6152) );
  INV_X1 U7912 ( .A(n7800), .ZN(n7949) );
  NAND2_X1 U7913 ( .A1(n7949), .A2(n7691), .ZN(n7677) );
  INV_X1 U7914 ( .A(n4398), .ZN(n8073) );
  XNOR2_X1 U7915 ( .A(n7701), .B(n8073), .ZN(n6231) );
  INV_X1 U7916 ( .A(n6231), .ZN(n6310) );
  OAI22_X1 U7917 ( .A1(n7677), .A2(n6310), .B1(n7790), .B2(n9548), .ZN(n6157)
         );
  OAI21_X1 U7918 ( .B1(n9804), .B2(n8108), .A(n8113), .ZN(n6208) );
  OR2_X1 U7919 ( .A1(n6159), .A2(n5782), .ZN(n6173) );
  NAND2_X1 U7920 ( .A1(n6160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6164) );
  XNOR2_X1 U7921 ( .A(n7452), .B(P2_B_REG_SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7922 ( .A1(n6168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6169) );
  INV_X1 U7923 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9989) );
  AND2_X1 U7924 ( .A1(n7675), .A2(n4421), .ZN(n6172) );
  NAND2_X1 U7925 ( .A1(n6173), .A2(n6172), .ZN(n6802) );
  NAND2_X1 U7926 ( .A1(n6173), .A2(n7675), .ZN(n6176) );
  NAND2_X1 U7927 ( .A1(n6384), .A2(n6358), .ZN(n6175) );
  NAND2_X1 U7928 ( .A1(n7483), .A2(n7479), .ZN(n6174) );
  NAND2_X1 U7929 ( .A1(n6176), .A2(n6799), .ZN(n6804) );
  NOR2_X1 U7930 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .ZN(
        n9905) );
  NOR4_X1 U7931 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6179) );
  NOR4_X1 U7932 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6178) );
  NOR4_X1 U7933 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7934 ( .A1(n9905), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n6185)
         );
  NOR4_X1 U7935 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6183) );
  NOR4_X1 U7936 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6182) );
  NOR4_X1 U7937 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6181) );
  NOR4_X1 U7938 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6180) );
  NAND4_X1 U7939 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n6184)
         );
  OAI21_X1 U7940 ( .B1(n6185), .B2(n6184), .A(n6384), .ZN(n6200) );
  INV_X1 U7941 ( .A(n7479), .ZN(n6186) );
  INV_X1 U7942 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7943 ( .A1(n6189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6191) );
  AND2_X1 U7944 ( .A1(n6200), .A2(n6385), .ZN(n6192) );
  NAND2_X1 U7945 ( .A1(n6297), .A2(n6192), .ZN(n6801) );
  INV_X1 U7946 ( .A(n6799), .ZN(n6194) );
  INV_X1 U7947 ( .A(n4421), .ZN(n6193) );
  OR2_X1 U7948 ( .A1(n6194), .A2(n6193), .ZN(n6204) );
  INV_X1 U7949 ( .A(n6198), .ZN(n6199) );
  NAND2_X1 U7950 ( .A1(n6199), .A2(n4367), .ZN(P2_U3487) );
  INV_X1 U7951 ( .A(n6200), .ZN(n6203) );
  AND2_X1 U7952 ( .A1(n6302), .A2(n6385), .ZN(n6308) );
  NAND3_X1 U7953 ( .A1(n9793), .A2(n6300), .A3(n7675), .ZN(n6283) );
  INV_X1 U7954 ( .A(n7698), .ZN(n9542) );
  NAND2_X1 U7955 ( .A1(n6283), .A2(n8278), .ZN(n6295) );
  NAND2_X1 U7956 ( .A1(n6308), .A2(n6295), .ZN(n6207) );
  NOR2_X1 U7957 ( .A1(n6204), .A2(n6203), .ZN(n6294) );
  NAND2_X1 U7958 ( .A1(n6307), .A2(n6300), .ZN(n6205) );
  NAND2_X1 U7959 ( .A1(n6291), .A2(n6205), .ZN(n6206) );
  INV_X1 U7960 ( .A(n6209), .ZN(n6210) );
  NAND2_X1 U7961 ( .A1(n6210), .A2(n4370), .ZN(P2_U3455) );
  NAND2_X1 U7962 ( .A1(n6211), .A2(n6233), .ZN(n6212) );
  AOI22_X1 U7963 ( .A1(n6213), .A2(n6212), .B1(n7950), .B2(n8111), .ZN(n6222)
         );
  NAND2_X1 U7964 ( .A1(n6215), .A2(n6214), .ZN(n6219) );
  INV_X1 U7965 ( .A(SI_28_), .ZN(n6216) );
  NAND2_X1 U7966 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  NAND2_X1 U7967 ( .A1(n6219), .A2(n6218), .ZN(n7485) );
  INV_X1 U7968 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9982) );
  INV_X1 U7969 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U7970 ( .A1(n8709), .A2(n7525), .ZN(n6221) );
  OR2_X1 U7971 ( .A1(n7526), .A2(n9982), .ZN(n6220) );
  NAND2_X1 U7972 ( .A1(n8101), .A2(n7800), .ZN(n7539) );
  NAND2_X1 U7973 ( .A1(n7674), .A2(n7539), .ZN(n7517) );
  XNOR2_X1 U7974 ( .A(n6222), .B(n7517), .ZN(n6223) );
  NAND2_X1 U7975 ( .A1(n6223), .A2(n9748), .ZN(n6236) );
  XNOR2_X1 U7976 ( .A(n7541), .B(n7517), .ZN(n6237) );
  INV_X1 U7977 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9948) );
  OR2_X1 U7978 ( .A1(n7530), .A2(n9948), .ZN(n6230) );
  INV_X1 U7979 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7980 ( .A1(n6226), .A2(n6225), .ZN(n6229) );
  INV_X1 U7981 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6227) );
  OR2_X1 U7982 ( .A1(n5817), .A2(n6227), .ZN(n6228) );
  NAND2_X1 U7983 ( .A1(n6443), .A2(P2_B_REG_SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7984 ( .A1(n9745), .A2(n6232), .ZN(n8089) );
  OAI22_X1 U7985 ( .A1(n6233), .A2(n9548), .B1(n7495), .B2(n8089), .ZN(n6234)
         );
  NAND2_X1 U7986 ( .A1(n6236), .A2(n6235), .ZN(n8096) );
  INV_X1 U7987 ( .A(n8096), .ZN(n6238) );
  INV_X1 U7988 ( .A(n6237), .ZN(n8105) );
  NAND2_X1 U7989 ( .A1(n6238), .A2(n4324), .ZN(n6241) );
  NAND2_X1 U7990 ( .A1(n6239), .A2(n4378), .ZN(n6240) );
  INV_X1 U7991 ( .A(n8101), .ZN(n7676) );
  NAND2_X1 U7992 ( .A1(n6240), .A2(n4928), .ZN(P2_U3456) );
  NAND2_X1 U7993 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  NAND2_X1 U7994 ( .A1(n6245), .A2(n4934), .ZN(P2_U3488) );
  INV_X4 U7995 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U7996 ( .A1(n7675), .A2(n6434), .ZN(n6248) );
  NAND2_X1 U7997 ( .A1(n6248), .A2(n7362), .ZN(n6441) );
  NAND2_X1 U7998 ( .A1(n6441), .A2(n6443), .ZN(n6249) );
  NAND2_X1 U7999 ( .A1(n6249), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U8000 ( .A(n6251), .B(n7551), .ZN(n8116) );
  XNOR2_X1 U8001 ( .A(n6252), .B(n7551), .ZN(n6256) );
  NAND2_X1 U8002 ( .A1(n7950), .A2(n9745), .ZN(n6254) );
  NAND2_X1 U8003 ( .A1(n8140), .A2(n9743), .ZN(n6253) );
  OAI21_X1 U8004 ( .B1(n9804), .B2(n8116), .A(n8121), .ZN(n8304) );
  INV_X1 U8005 ( .A(n8119), .ZN(n8306) );
  NOR2_X1 U8006 ( .A1(n8306), .A2(n8378), .ZN(n6257) );
  XNOR2_X1 U8007 ( .A(n7796), .B(n7245), .ZN(n6317) );
  XNOR2_X1 U8008 ( .A(n6317), .B(n6263), .ZN(n6290) );
  INV_X1 U8009 ( .A(n6268), .ZN(n6861) );
  NAND2_X1 U8010 ( .A1(n7750), .A2(n6861), .ZN(n6269) );
  XNOR2_X1 U8011 ( .A(n6271), .B(n9744), .ZN(n6673) );
  NAND2_X1 U8012 ( .A1(n6672), .A2(n6673), .ZN(n6671) );
  NAND2_X1 U8013 ( .A1(n6271), .A2(n5831), .ZN(n6272) );
  XNOR2_X1 U8014 ( .A(n7796), .B(n9751), .ZN(n6273) );
  XNOR2_X1 U8015 ( .A(n6273), .B(n7957), .ZN(n7774) );
  INV_X1 U8016 ( .A(n6273), .ZN(n6274) );
  NAND2_X1 U8017 ( .A1(n6274), .A2(n7957), .ZN(n6275) );
  XNOR2_X1 U8018 ( .A(n9766), .B(n7796), .ZN(n6276) );
  NAND2_X1 U8019 ( .A1(n9746), .A2(n6276), .ZN(n6278) );
  INV_X1 U8020 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U8021 ( .A1(n6982), .A2(n6277), .ZN(n6973) );
  AND2_X1 U8022 ( .A1(n6278), .A2(n6973), .ZN(n7857) );
  NAND2_X1 U8023 ( .A1(n6972), .A2(n6973), .ZN(n6279) );
  XNOR2_X1 U8024 ( .A(n7796), .B(n7094), .ZN(n6280) );
  XNOR2_X1 U8025 ( .A(n6280), .B(n7956), .ZN(n6974) );
  NAND2_X1 U8026 ( .A1(n7102), .A2(n6280), .ZN(n6281) );
  INV_X1 U8027 ( .A(n6300), .ZN(n6282) );
  NAND2_X1 U8028 ( .A1(n6308), .A2(n6282), .ZN(n6286) );
  INV_X1 U8029 ( .A(n6283), .ZN(n6284) );
  NAND2_X1 U8030 ( .A1(n6291), .A2(n6284), .ZN(n6285) );
  INV_X1 U8031 ( .A(n6320), .ZN(n6288) );
  AOI211_X1 U8032 ( .C1(n6290), .C2(n6289), .A(n7932), .B(n6288), .ZN(n6316)
         );
  NAND2_X1 U8033 ( .A1(n6291), .A2(n9816), .ZN(n6293) );
  INV_X1 U8034 ( .A(n7930), .ZN(n7947) );
  NOR2_X1 U8035 ( .A1(n7947), .A2(n9776), .ZN(n6315) );
  INV_X1 U8036 ( .A(n6294), .ZN(n6296) );
  NAND2_X1 U8037 ( .A1(n6296), .A2(n6295), .ZN(n6299) );
  AND3_X1 U8038 ( .A1(n6297), .A2(n6434), .A3(n7362), .ZN(n6298) );
  OAI211_X1 U8039 ( .C1(n6302), .C2(n6300), .A(n6299), .B(n6298), .ZN(n6301)
         );
  NAND2_X1 U8040 ( .A1(n6301), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6306) );
  INV_X1 U8041 ( .A(n6302), .ZN(n6304) );
  INV_X1 U8042 ( .A(n6385), .ZN(n6303) );
  NOR2_X1 U8043 ( .A1(n6307), .A2(n6303), .ZN(n7702) );
  NAND2_X1 U8044 ( .A1(n6304), .A2(n7702), .ZN(n6305) );
  NOR2_X1 U8045 ( .A1(n7928), .A2(n7243), .ZN(n6314) );
  INV_X1 U8046 ( .A(n6307), .ZN(n6855) );
  AND2_X1 U8047 ( .A1(n6308), .A2(n6855), .ZN(n6311) );
  INV_X1 U8048 ( .A(n6311), .ZN(n6309) );
  NAND2_X1 U8049 ( .A1(n7940), .A2(n7956), .ZN(n6312) );
  NAND2_X1 U8050 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9877) );
  OAI211_X1 U8051 ( .C1(n6322), .C2(n7942), .A(n6312), .B(n9877), .ZN(n6313)
         );
  OR4_X1 U8052 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(P2_U3179)
         );
  XNOR2_X1 U8053 ( .A(n7378), .B(n7796), .ZN(n7453) );
  XNOR2_X1 U8054 ( .A(n7453), .B(n7424), .ZN(n6331) );
  INV_X1 U8055 ( .A(n6317), .ZN(n6318) );
  NAND2_X1 U8056 ( .A1(n7955), .A2(n6318), .ZN(n6319) );
  XNOR2_X1 U8057 ( .A(n7750), .B(n7195), .ZN(n6321) );
  NAND2_X1 U8058 ( .A1(n9729), .A2(n6321), .ZN(n6324) );
  INV_X1 U8059 ( .A(n6321), .ZN(n6323) );
  NAND2_X1 U8060 ( .A1(n6323), .A2(n6322), .ZN(n7311) );
  AND2_X1 U8061 ( .A1(n6324), .A2(n7311), .ZN(n7188) );
  NAND2_X1 U8062 ( .A1(n7187), .A2(n7311), .ZN(n6325) );
  XNOR2_X1 U8063 ( .A(n9738), .B(n7796), .ZN(n6326) );
  XNOR2_X1 U8064 ( .A(n6326), .B(n7954), .ZN(n7312) );
  NAND2_X1 U8065 ( .A1(n6326), .A2(n7371), .ZN(n6327) );
  INV_X1 U8066 ( .A(n6331), .ZN(n6328) );
  INV_X1 U8067 ( .A(n7456), .ZN(n6329) );
  AOI211_X1 U8068 ( .C1(n6331), .C2(n6330), .A(n7932), .B(n6329), .ZN(n6336)
         );
  NOR2_X1 U8069 ( .A1(n9794), .A2(n7947), .ZN(n6335) );
  NOR2_X1 U8070 ( .A1(n7928), .A2(n7376), .ZN(n6334) );
  NAND2_X1 U8071 ( .A1(n7940), .A2(n7954), .ZN(n6332) );
  NAND2_X1 U8072 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6846) );
  OAI211_X1 U8073 ( .C1(n7473), .C2(n7942), .A(n6332), .B(n6846), .ZN(n6333)
         );
  OR4_X1 U8074 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(P2_U3171)
         );
  NOR2_X1 U8075 ( .A1(n7521), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9509) );
  INV_X2 U8076 ( .A(n9509), .ZN(n9522) );
  AND2_X1 U8077 ( .A1(n7521), .A2(P1_U3086), .ZN(n7358) );
  INV_X2 U8078 ( .A(n7358), .ZN(n9514) );
  OAI222_X1 U8079 ( .A1(n9522), .A2(n6337), .B1(n9514), .B2(n6343), .C1(
        P1_U3086), .C2(n6414), .ZN(P1_U3354) );
  OAI222_X1 U8080 ( .A1(n9522), .A2(n6338), .B1(n9514), .B2(n6341), .C1(
        P1_U3086), .C2(n6415), .ZN(P1_U3353) );
  OAI222_X1 U8081 ( .A1(n9522), .A2(n9992), .B1(n9514), .B2(n6340), .C1(
        P1_U3086), .C2(n6416), .ZN(P1_U3352) );
  INV_X2 U8082 ( .A(n7360), .ZN(n8451) );
  INV_X2 U8083 ( .A(n8446), .ZN(n8449) );
  OAI222_X1 U8084 ( .A1(n6561), .A2(P2_U3151), .B1(n8451), .B2(n6340), .C1(
        n6339), .C2(n8449), .ZN(P2_U3292) );
  OAI222_X1 U8085 ( .A1(n8449), .A2(n6342), .B1(n8451), .B2(n6341), .C1(n6492), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8086 ( .A1(n6545), .A2(P2_U3151), .B1(n8451), .B2(n6343), .C1(
        n8449), .C2(n4992), .ZN(P2_U3294) );
  OAI222_X1 U8087 ( .A1(n9522), .A2(n6344), .B1(n9514), .B2(n6346), .C1(
        P1_U3086), .C2(n6906), .ZN(P1_U3351) );
  OAI222_X1 U8088 ( .A1(n6635), .A2(P2_U3151), .B1(n8451), .B2(n6346), .C1(
        n6345), .C2(n8449), .ZN(P2_U3291) );
  INV_X1 U8089 ( .A(n8926), .ZN(n6908) );
  OAI222_X1 U8090 ( .A1(n9522), .A2(n6347), .B1(n9514), .B2(n6349), .C1(
        P1_U3086), .C2(n6908), .ZN(P1_U3350) );
  OAI222_X1 U8091 ( .A1(n6698), .A2(P2_U3151), .B1(n8451), .B2(n6349), .C1(
        n6348), .C2(n8449), .ZN(P2_U3290) );
  OAI222_X1 U8092 ( .A1(n9871), .A2(P2_U3151), .B1(n8451), .B2(n6351), .C1(
        n6350), .C2(n8449), .ZN(P2_U3289) );
  INV_X1 U8093 ( .A(n8940), .ZN(n6910) );
  OAI222_X1 U8094 ( .A1(n9522), .A2(n6352), .B1(n9514), .B2(n6351), .C1(
        P1_U3086), .C2(n6910), .ZN(P1_U3349) );
  INV_X1 U8095 ( .A(n6747), .ZN(n6754) );
  INV_X1 U8096 ( .A(n6353), .ZN(n6355) );
  INV_X1 U8097 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6354) );
  OAI222_X1 U8098 ( .A1(n6754), .A2(P2_U3151), .B1(n8451), .B2(n6355), .C1(
        n6354), .C2(n8449), .ZN(P2_U3288) );
  INV_X1 U8099 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6356) );
  INV_X1 U8100 ( .A(n8954), .ZN(n6911) );
  OAI222_X1 U8101 ( .A1(n9522), .A2(n6356), .B1(n9514), .B2(n6355), .C1(
        P1_U3086), .C2(n6911), .ZN(P1_U3348) );
  NAND2_X1 U8102 ( .A1(n6799), .A2(n6385), .ZN(n6357) );
  OAI21_X1 U8103 ( .B1(n6385), .B2(n6358), .A(n6357), .ZN(P2_U3377) );
  INV_X1 U8104 ( .A(n6359), .ZN(n6362) );
  AOI22_X1 U8105 ( .A1(n8968), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9509), .ZN(n6360) );
  OAI21_X1 U8106 ( .B1(n6362), .B2(n9514), .A(n6360), .ZN(P1_U3347) );
  OAI222_X1 U8107 ( .A1(n6844), .A2(P2_U3151), .B1(n8451), .B2(n6362), .C1(
        n6361), .C2(n8449), .ZN(P2_U3287) );
  NAND2_X1 U8108 ( .A1(n4391), .A2(P1_U3973), .ZN(n6363) );
  OAI21_X1 U8109 ( .B1(P1_U3973), .B2(n4992), .A(n6363), .ZN(P1_U3555) );
  INV_X1 U8110 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U8111 ( .A1(n6581), .A2(P1_U3973), .ZN(n6364) );
  OAI21_X1 U8112 ( .B1(P1_U3973), .B2(n9946), .A(n6364), .ZN(P1_U3554) );
  INV_X1 U8113 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6369) );
  INV_X1 U8114 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U8115 ( .A1(n6365), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6367) );
  INV_X1 U8116 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9449) );
  OR2_X1 U8117 ( .A1(n4420), .A2(n9449), .ZN(n6366) );
  OAI211_X1 U8118 ( .C1(n9356), .C2(n4272), .A(n6367), .B(n6366), .ZN(n9052)
         );
  NAND2_X1 U8119 ( .A1(n9052), .A2(P1_U3973), .ZN(n6368) );
  OAI21_X1 U8120 ( .B1(P1_U3973), .B2(n6369), .A(n6368), .ZN(P1_U3585) );
  OR2_X1 U8121 ( .A1(n6371), .A2(P1_U3086), .ZN(n8866) );
  INV_X1 U8122 ( .A(n8866), .ZN(n6370) );
  NAND2_X1 U8123 ( .A1(n6372), .A2(n6371), .ZN(n6374) );
  NAND2_X1 U8124 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  INV_X1 U8125 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6383) );
  INV_X1 U8126 ( .A(n6375), .ZN(n6376) );
  AND2_X1 U8127 ( .A1(n6377), .A2(n6376), .ZN(n6418) );
  OAI21_X1 U8128 ( .B1(n9523), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6426), .ZN(
        n6428) );
  AOI21_X1 U8129 ( .B1(n9523), .B2(n6379), .A(n6428), .ZN(n6380) );
  INV_X1 U8130 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U8131 ( .A(n6380), .B(n6429), .ZN(n6381) );
  AOI22_X1 U8132 ( .A1(n6418), .A2(n6381), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6382) );
  OAI21_X1 U8133 ( .B1(n9650), .B2(n6383), .A(n6382), .ZN(P1_U3243) );
  INV_X1 U8134 ( .A(n9650), .ZN(n9014) );
  NOR2_X1 U8135 ( .A1(n9014), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8136 ( .A(n6384), .ZN(n6386) );
  AOI22_X1 U8137 ( .A1(n6399), .A2(n9989), .B1(n6387), .B2(n4305), .ZN(
        P2_U3376) );
  INV_X1 U8138 ( .A(n6388), .ZN(n6396) );
  AOI22_X1 U8139 ( .A1(n8984), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9509), .ZN(n6389) );
  OAI21_X1 U8140 ( .B1(n6396), .B2(n9514), .A(n6389), .ZN(P1_U3346) );
  NAND2_X1 U8141 ( .A1(n9681), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6391) );
  OAI21_X1 U8142 ( .B1(n9681), .B2(n6392), .A(n6391), .ZN(P1_U3439) );
  INV_X1 U8143 ( .A(n6393), .ZN(n6398) );
  AOI22_X1 U8144 ( .A1(n9534), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9509), .ZN(n6394) );
  OAI21_X1 U8145 ( .B1(n6398), .B2(n9514), .A(n6394), .ZN(P1_U3345) );
  AND2_X1 U8146 ( .A1(n6399), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8147 ( .A1(n6399), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8148 ( .A1(n6399), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8149 ( .A1(n6399), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8150 ( .A1(n6399), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8151 ( .A1(n6399), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8152 ( .A1(n6399), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8153 ( .A1(n6399), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8154 ( .A1(n6399), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8155 ( .A1(n6399), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8156 ( .A1(n6399), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8157 ( .A1(n6399), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8158 ( .A1(n6399), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8159 ( .A1(n6399), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8160 ( .A1(n6399), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8161 ( .A1(n6399), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8162 ( .A1(n6399), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8163 ( .A1(n6399), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8164 ( .A1(n6399), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8165 ( .A1(n6399), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8166 ( .A1(n6399), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8167 ( .A1(n6399), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8168 ( .A1(n6399), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8169 ( .A1(n6399), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8170 ( .A1(n6399), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  OAI222_X1 U8171 ( .A1(P2_U3151), .A2(n4555), .B1(n8451), .B2(n6396), .C1(
        n6395), .C2(n8449), .ZN(P2_U3286) );
  OAI222_X1 U8172 ( .A1(P2_U3151), .A2(n7067), .B1(n8451), .B2(n6398), .C1(
        n6397), .C2(n8449), .ZN(P2_U3285) );
  INV_X1 U8173 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U8174 ( .A1(n6400), .A2(n9957), .ZN(P2_U3253) );
  INV_X1 U8175 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9963) );
  NOR2_X1 U8176 ( .A1(n6400), .A2(n9963), .ZN(P2_U3261) );
  INV_X1 U8177 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9978) );
  NOR2_X1 U8178 ( .A1(n6400), .A2(n9978), .ZN(P2_U3251) );
  INV_X1 U8179 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U8180 ( .A1(n6400), .A2(n9928), .ZN(P2_U3249) );
  INV_X1 U8181 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U8182 ( .A1(n6400), .A2(n10008), .ZN(P2_U3260) );
  INV_X1 U8183 ( .A(n6401), .ZN(n6404) );
  INV_X1 U8184 ( .A(n9579), .ZN(n6402) );
  OAI222_X1 U8185 ( .A1(n9522), .A2(n9920), .B1(n9514), .B2(n6404), .C1(
        P1_U3086), .C2(n6402), .ZN(P1_U3344) );
  OAI222_X1 U8186 ( .A1(n4773), .A2(P2_U3151), .B1(n8451), .B2(n6404), .C1(
        n6403), .C2(n8449), .ZN(P2_U3284) );
  INV_X1 U8187 ( .A(n6906), .ZN(n6895) );
  INV_X1 U8188 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6412) );
  XNOR2_X1 U8189 ( .A(n6906), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6410) );
  INV_X1 U8190 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9654) );
  MUX2_X1 U8191 ( .A(n9654), .B(P1_REG2_REG_2__SCAN_IN), .S(n6415), .Z(n8898)
         );
  INV_X1 U8192 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6405) );
  MUX2_X1 U8193 ( .A(n6405), .B(P1_REG2_REG_1__SCAN_IN), .S(n6414), .Z(n8889)
         );
  AND2_X1 U8194 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8888) );
  NAND2_X1 U8195 ( .A1(n8889), .A2(n8888), .ZN(n8887) );
  INV_X1 U8196 ( .A(n6414), .ZN(n8883) );
  NAND2_X1 U8197 ( .A1(n8883), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8198 ( .A1(n8887), .A2(n6406), .ZN(n8897) );
  NAND2_X1 U8199 ( .A1(n8898), .A2(n8897), .ZN(n8896) );
  INV_X1 U8200 ( .A(n6415), .ZN(n8895) );
  NAND2_X1 U8201 ( .A1(n8895), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8202 ( .A1(n8896), .A2(n6407), .ZN(n8914) );
  INV_X1 U8203 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9975) );
  MUX2_X1 U8204 ( .A(n9975), .B(P1_REG2_REG_3__SCAN_IN), .S(n6416), .Z(n8915)
         );
  NAND2_X1 U8205 ( .A1(n8914), .A2(n8915), .ZN(n8913) );
  INV_X1 U8206 ( .A(n6416), .ZN(n8912) );
  NAND2_X1 U8207 ( .A1(n8912), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8208 ( .A1(n8913), .A2(n6408), .ZN(n6409) );
  OR2_X1 U8209 ( .A1(n9520), .A2(n9523), .ZN(n8861) );
  INV_X1 U8210 ( .A(n8861), .ZN(n6427) );
  NAND2_X1 U8211 ( .A1(n6409), .A2(n6410), .ZN(n6905) );
  OAI211_X1 U8212 ( .C1(n6410), .C2(n6409), .A(n9642), .B(n6905), .ZN(n6411)
         );
  NAND2_X1 U8213 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n6739) );
  OAI211_X1 U8214 ( .C1(n9650), .C2(n6412), .A(n6411), .B(n6739), .ZN(n6422)
         );
  MUX2_X1 U8215 ( .A(n6413), .B(P1_REG1_REG_1__SCAN_IN), .S(n6414), .Z(n8886)
         );
  OAI21_X1 U8216 ( .B1(n6414), .B2(n6413), .A(n8884), .ZN(n8900) );
  MUX2_X1 U8217 ( .A(n5053), .B(P1_REG1_REG_2__SCAN_IN), .S(n6415), .Z(n8901)
         );
  MUX2_X1 U8218 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6417), .S(n6416), .Z(n8907)
         );
  NOR2_X1 U8219 ( .A1(n4321), .A2(n8907), .ZN(n8906) );
  XOR2_X1 U8220 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6906), .Z(n6419) );
  NOR2_X1 U8221 ( .A1(n6420), .A2(n6419), .ZN(n6894) );
  AOI211_X1 U8222 ( .C1(n6420), .C2(n6419), .A(n6894), .B(n9619), .ZN(n6421)
         );
  AOI211_X1 U8223 ( .C1(n9630), .C2(n6895), .A(n6422), .B(n6421), .ZN(n6432)
         );
  INV_X1 U8224 ( .A(n6423), .ZN(n6425) );
  XNOR2_X1 U8225 ( .A(n6425), .B(n6424), .ZN(n6452) );
  NAND2_X1 U8226 ( .A1(n6426), .A2(n9523), .ZN(n6431) );
  AOI22_X1 U8227 ( .A1(n6429), .A2(n6428), .B1(n6427), .B2(n8888), .ZN(n6430)
         );
  OAI211_X1 U8228 ( .C1(n6452), .C2(n6431), .A(P1_U3973), .B(n6430), .ZN(n8905) );
  NAND2_X1 U8229 ( .A1(n6432), .A2(n8905), .ZN(P1_U3247) );
  INV_X1 U8230 ( .A(n7362), .ZN(n6433) );
  NOR2_X1 U8231 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  INV_X1 U8232 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6447) );
  NOR2_X1 U8233 ( .A1(n6155), .A2(P2_U3151), .ZN(n8445) );
  INV_X1 U8234 ( .A(n6475), .ZN(n6499) );
  NAND2_X1 U8235 ( .A1(P2_U3893), .A2(n6155), .ZN(n8082) );
  INV_X1 U8236 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6476) );
  MUX2_X1 U8237 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n4398), .Z(n6438) );
  MUX2_X1 U8238 ( .A(n6859), .B(n6436), .S(n4398), .Z(n6437) );
  NAND2_X1 U8239 ( .A1(n6437), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6533) );
  INV_X1 U8240 ( .A(n6533), .ZN(n6468) );
  AOI21_X1 U8241 ( .B1(n6476), .B2(n6438), .A(n6468), .ZN(n6439) );
  AOI21_X1 U8242 ( .B1(n6499), .B2(n8082), .A(n6439), .ZN(n6440) );
  AOI21_X1 U8243 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6440), .ZN(
        n6446) );
  AND2_X1 U8244 ( .A1(n6441), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6442) );
  MUX2_X1 U8245 ( .A(P2_U3893), .B(n6442), .S(n6155), .Z(n6444) );
  NAND2_X1 U8246 ( .A1(n9882), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6445) );
  OAI211_X1 U8247 ( .C1(n9880), .C2(n6447), .A(n6446), .B(n6445), .ZN(P2_U3182) );
  INV_X1 U8248 ( .A(n6448), .ZN(n6451) );
  INV_X1 U8249 ( .A(n8999), .ZN(n6923) );
  OAI222_X1 U8250 ( .A1(n9514), .A2(n6451), .B1(n6923), .B2(P1_U3086), .C1(
        n6449), .C2(n9522), .ZN(P1_U3343) );
  OAI222_X1 U8251 ( .A1(P2_U3151), .A2(n7383), .B1(n8451), .B2(n6451), .C1(
        n6450), .C2(n8449), .ZN(P2_U3283) );
  NOR2_X1 U8252 ( .A1(n8568), .A2(P1_U3086), .ZN(n6507) );
  AND2_X1 U8253 ( .A1(n4391), .A2(n8588), .ZN(n9675) );
  AOI22_X1 U8254 ( .A1(n9571), .A2(n6452), .B1(n9566), .B2(n9675), .ZN(n6454)
         );
  NAND2_X1 U8255 ( .A1(n8613), .A2(n6585), .ZN(n6453) );
  OAI211_X1 U8256 ( .C1(n6507), .C2(n9672), .A(n6454), .B(n6453), .ZN(P1_U3232) );
  INV_X1 U8257 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9959) );
  INV_X1 U8258 ( .A(n6455), .ZN(n6457) );
  INV_X1 U8259 ( .A(n9593), .ZN(n8997) );
  OAI222_X1 U8260 ( .A1(n9522), .A2(n9959), .B1(n9514), .B2(n6457), .C1(
        P1_U3086), .C2(n8997), .ZN(P1_U3342) );
  INV_X1 U8261 ( .A(n7960), .ZN(n7966) );
  INV_X1 U8262 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6456) );
  OAI222_X1 U8263 ( .A1(n7966), .A2(P2_U3151), .B1(n8451), .B2(n6457), .C1(
        n6456), .C2(n8449), .ZN(P2_U3282) );
  INV_X1 U8264 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9653) );
  INV_X1 U8265 ( .A(n6458), .ZN(n6463) );
  NOR3_X1 U8266 ( .A1(n6459), .A2(n6461), .A3(n6460), .ZN(n6462) );
  OAI21_X1 U8267 ( .B1(n6463), .B2(n6462), .A(n9571), .ZN(n6465) );
  INV_X1 U8268 ( .A(n8815), .ZN(n6587) );
  OAI22_X1 U8269 ( .A1(n6587), .A2(n8508), .B1(n6617), .B2(n9051), .ZN(n6728)
         );
  AOI22_X1 U8270 ( .A1(n8613), .A2(n9656), .B1(n9566), .B2(n6728), .ZN(n6464)
         );
  OAI211_X1 U8271 ( .C1(n6507), .C2(n9653), .A(n6465), .B(n6464), .ZN(P1_U3237) );
  MUX2_X1 U8272 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n4398), .Z(n6466) );
  XNOR2_X1 U8273 ( .A(n6466), .B(n6545), .ZN(n6534) );
  INV_X1 U8274 ( .A(n6466), .ZN(n6467) );
  OAI22_X1 U8275 ( .A1(n6534), .A2(n6468), .B1(n6488), .B2(n6467), .ZN(n6517)
         );
  MUX2_X1 U8276 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4398), .Z(n6469) );
  XNOR2_X1 U8277 ( .A(n6469), .B(n6530), .ZN(n6516) );
  AOI22_X1 U8278 ( .A1(n6517), .A2(n6516), .B1(n6469), .B2(n6492), .ZN(n6557)
         );
  MUX2_X1 U8279 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4398), .Z(n6470) );
  XOR2_X1 U8280 ( .A(n6561), .B(n6470), .Z(n6556) );
  NAND2_X1 U8281 ( .A1(n6557), .A2(n6556), .ZN(n6555) );
  INV_X1 U8282 ( .A(n6470), .ZN(n6471) );
  INV_X1 U8283 ( .A(n6561), .ZN(n6493) );
  NAND2_X1 U8284 ( .A1(n6471), .A2(n6493), .ZN(n6472) );
  AND2_X1 U8285 ( .A1(n6555), .A2(n6472), .ZN(n6474) );
  MUX2_X1 U8286 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4398), .Z(n6630) );
  XOR2_X1 U8287 ( .A(n6635), .B(n6630), .Z(n6473) );
  NAND3_X1 U8288 ( .A1(n6555), .A2(n6472), .A3(n6473), .ZN(n6631) );
  OAI211_X1 U8289 ( .C1(n6474), .C2(n6473), .A(n9887), .B(n6631), .ZN(n6504)
         );
  INV_X1 U8290 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9822) );
  MUX2_X1 U8291 ( .A(n9822), .B(P2_REG1_REG_4__SCAN_IN), .S(n6635), .Z(n6485)
         );
  XNOR2_X1 U8292 ( .A(n6530), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8293 ( .A1(n5804), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8294 ( .A1(n6545), .A2(n6480), .ZN(n6479) );
  NAND2_X1 U8295 ( .A1(n6476), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6477) );
  OR2_X1 U8296 ( .A1(n6477), .A2(n5804), .ZN(n6478) );
  NAND2_X1 U8297 ( .A1(n6479), .A2(n6478), .ZN(n6538) );
  NAND2_X1 U8298 ( .A1(n6538), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8299 ( .A1(n6481), .A2(n6480), .ZN(n6523) );
  AOI22_X1 U8300 ( .A1(n6524), .A2(n6523), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n6492), .ZN(n6482) );
  INV_X1 U8301 ( .A(n6482), .ZN(n6483) );
  NOR2_X1 U8302 ( .A1(n6484), .A2(n6485), .ZN(n6634) );
  AOI21_X1 U8303 ( .B1(n6485), .B2(n6484), .A(n6634), .ZN(n6487) );
  INV_X1 U8304 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6486) );
  OAI22_X1 U8305 ( .A1(n9891), .A2(n6487), .B1(n9880), .B2(n6486), .ZN(n6502)
         );
  AND2_X1 U8306 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U8307 ( .A1(n5804), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8308 ( .A1(n6489), .A2(n6490), .ZN(n6536) );
  NOR2_X1 U8309 ( .A1(n6536), .A2(n7021), .ZN(n6535) );
  INV_X1 U8310 ( .A(n6490), .ZN(n6491) );
  NOR2_X1 U8311 ( .A1(n6535), .A2(n6491), .ZN(n6519) );
  NOR2_X1 U8312 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  INV_X1 U8313 ( .A(n6496), .ZN(n6497) );
  XNOR2_X1 U8314 ( .A(n6635), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6498) );
  NAND3_X1 U8315 ( .A1(n6548), .A2(n6498), .A3(n6497), .ZN(n6500) );
  AOI21_X1 U8316 ( .B1(n4382), .B2(n6500), .A(n8086), .ZN(n6501) );
  NOR3_X1 U8317 ( .A1(n6502), .A2(n7860), .A3(n6501), .ZN(n6503) );
  OAI211_X1 U8318 ( .C1(n8050), .C2(n6635), .A(n6504), .B(n6503), .ZN(P2_U3186) );
  AOI21_X1 U8319 ( .B1(n6506), .B2(n6505), .A(n6459), .ZN(n6511) );
  INV_X1 U8320 ( .A(n6507), .ZN(n6509) );
  AOI22_X1 U8321 ( .A1(n8588), .A2(n8880), .B1(n6581), .B2(n9074), .ZN(n6603)
         );
  OAI22_X1 U8322 ( .A1(n9568), .A2(n8814), .B1(n6603), .B2(n8601), .ZN(n6508)
         );
  AOI21_X1 U8323 ( .B1(n6509), .B2(P1_REG3_REG_1__SCAN_IN), .A(n6508), .ZN(
        n6510) );
  OAI21_X1 U8324 ( .B1(n6511), .B2(n8615), .A(n6510), .ZN(P1_U3222) );
  INV_X1 U8325 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6513) );
  INV_X1 U8326 ( .A(n6512), .ZN(n6515) );
  INV_X1 U8327 ( .A(n9608), .ZN(n9000) );
  OAI222_X1 U8328 ( .A1(n9522), .A2(n6513), .B1(n9514), .B2(n6515), .C1(
        P1_U3086), .C2(n9000), .ZN(P1_U3341) );
  INV_X1 U8329 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6514) );
  OAI222_X1 U8330 ( .A1(n7990), .A2(P2_U3151), .B1(n8451), .B2(n6515), .C1(
        n6514), .C2(n8449), .ZN(P2_U3281) );
  XNOR2_X1 U8331 ( .A(n6517), .B(n6516), .ZN(n6532) );
  AOI21_X1 U8332 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6522) );
  INV_X1 U8333 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6521) );
  OAI22_X1 U8334 ( .A1(n8086), .A2(n6522), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6521), .ZN(n6529) );
  INV_X1 U8335 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6527) );
  XNOR2_X1 U8336 ( .A(n6524), .B(n6523), .ZN(n6525) );
  NAND2_X1 U8337 ( .A1(n9720), .A2(n6525), .ZN(n6526) );
  OAI21_X1 U8338 ( .B1(n6527), .B2(n9880), .A(n6526), .ZN(n6528) );
  AOI211_X1 U8339 ( .C1(n6530), .C2(n9882), .A(n6529), .B(n6528), .ZN(n6531)
         );
  OAI21_X1 U8340 ( .B1(n8082), .B2(n6532), .A(n6531), .ZN(P2_U3184) );
  XNOR2_X1 U8341 ( .A(n6534), .B(n6533), .ZN(n6543) );
  INV_X1 U8342 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9839) );
  AOI21_X1 U8343 ( .B1(n7021), .B2(n6536), .A(n6535), .ZN(n6537) );
  OAI22_X1 U8344 ( .A1(n9880), .A2(n9839), .B1(n8086), .B2(n6537), .ZN(n6542)
         );
  XNOR2_X1 U8345 ( .A(n6538), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8346 ( .A1(n9720), .A2(n6539), .ZN(n6540) );
  OAI21_X1 U8347 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7023), .A(n6540), .ZN(n6541) );
  AOI211_X1 U8348 ( .C1(n9887), .C2(n6543), .A(n6542), .B(n6541), .ZN(n6544)
         );
  OAI21_X1 U8349 ( .B1(n6545), .B2(n8050), .A(n6544), .ZN(P2_U3183) );
  XNOR2_X1 U8350 ( .A(n6546), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6554) );
  AND2_X1 U8351 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7776) );
  INV_X1 U8352 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6552) );
  INV_X1 U8353 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9756) );
  INV_X1 U8354 ( .A(n6547), .ZN(n6550) );
  INV_X1 U8355 ( .A(n6548), .ZN(n6549) );
  AOI21_X1 U8356 ( .B1(n9756), .B2(n6550), .A(n6549), .ZN(n6551) );
  OAI22_X1 U8357 ( .A1(n9880), .A2(n6552), .B1(n6551), .B2(n8086), .ZN(n6553)
         );
  AOI211_X1 U8358 ( .C1(n9720), .C2(n6554), .A(n7776), .B(n6553), .ZN(n6560)
         );
  OAI21_X1 U8359 ( .B1(n6557), .B2(n6556), .A(n6555), .ZN(n6558) );
  NAND2_X1 U8360 ( .A1(n6558), .A2(n9887), .ZN(n6559) );
  OAI211_X1 U8361 ( .C1(n8050), .C2(n6561), .A(n6560), .B(n6559), .ZN(P2_U3185) );
  AND2_X1 U8362 ( .A1(n6563), .A2(n6562), .ZN(n6568) );
  NAND2_X1 U8363 ( .A1(n6565), .A2(n6564), .ZN(n6567) );
  INV_X1 U8364 ( .A(n6585), .ZN(n6599) );
  AND2_X1 U8365 ( .A1(n6581), .A2(n6599), .ZN(n8813) );
  NOR2_X1 U8366 ( .A1(n6601), .A2(n8813), .ZN(n9667) );
  NAND2_X1 U8367 ( .A1(n6569), .A2(n6576), .ZN(n9668) );
  AND2_X1 U8368 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  OR2_X1 U8369 ( .A1(n9668), .A2(n6572), .ZN(n6723) );
  NAND2_X1 U8370 ( .A1(n8863), .A2(n9040), .ZN(n6574) );
  NAND2_X1 U8371 ( .A1(n5719), .A2(n8860), .ZN(n6573) );
  NOR2_X1 U8372 ( .A1(n9695), .A2(n9333), .ZN(n6575) );
  OR2_X1 U8373 ( .A1(n9667), .A2(n6575), .ZN(n6579) );
  INV_X1 U8374 ( .A(n6576), .ZN(n6577) );
  AND2_X1 U8375 ( .A1(n6585), .A2(n6577), .ZN(n9669) );
  NOR2_X1 U8376 ( .A1(n9675), .A2(n9669), .ZN(n6578) );
  AND2_X1 U8377 ( .A1(n6579), .A2(n6578), .ZN(n9682) );
  NAND2_X1 U8378 ( .A1(n9710), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U8379 ( .B1(n9710), .B2(n9682), .A(n6580), .ZN(P1_U3522) );
  NAND2_X1 U8380 ( .A1(n6581), .A2(n6585), .ZN(n6598) );
  NAND2_X1 U8381 ( .A1(n6587), .A2(n8814), .ZN(n6582) );
  NAND2_X1 U8382 ( .A1(n6597), .A2(n6582), .ZN(n6716) );
  XNOR2_X1 U8383 ( .A(n8880), .B(n6731), .ZN(n6724) );
  INV_X1 U8384 ( .A(n8880), .ZN(n6588) );
  NAND2_X1 U8385 ( .A1(n6588), .A2(n6731), .ZN(n6583) );
  NAND2_X1 U8386 ( .A1(n6718), .A2(n6583), .ZN(n6584) );
  OAI21_X1 U8387 ( .B1(n6584), .B2(n8772), .A(n6608), .ZN(n7128) );
  INV_X1 U8388 ( .A(n6722), .ZN(n6586) );
  AOI211_X1 U8389 ( .C1(n6650), .C2(n6586), .A(n9342), .B(n4609), .ZN(n7124)
         );
  NAND2_X1 U8390 ( .A1(n8770), .A2(n6601), .ZN(n6614) );
  AND2_X1 U8391 ( .A1(n6614), .A2(n6613), .ZN(n6725) );
  NAND2_X1 U8392 ( .A1(n6588), .A2(n9656), .ZN(n6612) );
  OAI21_X1 U8393 ( .B1(n6725), .B2(n6724), .A(n6612), .ZN(n6589) );
  XNOR2_X1 U8394 ( .A(n6589), .B(n8772), .ZN(n6593) );
  NAND2_X1 U8395 ( .A1(n8878), .A2(n8588), .ZN(n6591) );
  NAND2_X1 U8396 ( .A1(n8880), .A2(n9074), .ZN(n6590) );
  NAND2_X1 U8397 ( .A1(n6591), .A2(n6590), .ZN(n6677) );
  INV_X1 U8398 ( .A(n6677), .ZN(n6592) );
  OAI21_X1 U8399 ( .B1(n6593), .B2(n9240), .A(n6592), .ZN(n7123) );
  AOI211_X1 U8400 ( .C1(n9695), .C2(n7128), .A(n7124), .B(n7123), .ZN(n6652)
         );
  INV_X1 U8401 ( .A(n6594), .ZN(n6938) );
  AOI22_X1 U8402 ( .A1(n9456), .A2(n6650), .B1(n9706), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n6596) );
  OAI21_X1 U8403 ( .B1(n6652), .B2(n9706), .A(n6596), .ZN(P1_U3462) );
  OAI21_X1 U8404 ( .B1(n6602), .B2(n6598), .A(n6597), .ZN(n6986) );
  OR2_X1 U8405 ( .A1(n8814), .A2(n6599), .ZN(n6600) );
  AND3_X1 U8406 ( .A1(n6600), .A2(n9216), .A3(n6719), .ZN(n6988) );
  XNOR2_X1 U8407 ( .A(n6602), .B(n6601), .ZN(n6604) );
  OAI21_X1 U8408 ( .B1(n6604), .B2(n9240), .A(n6603), .ZN(n6989) );
  AOI211_X1 U8409 ( .C1(n9695), .C2(n6986), .A(n6988), .B(n6989), .ZN(n6654)
         );
  OAI22_X1 U8410 ( .A1(n9503), .A2(n8814), .B1(n9707), .B2(n5022), .ZN(n6605)
         );
  INV_X1 U8411 ( .A(n6605), .ZN(n6606) );
  OAI21_X1 U8412 ( .B1(n6654), .B2(n9706), .A(n6606), .ZN(P1_U3456) );
  NAND2_X1 U8413 ( .A1(n6617), .A2(n8819), .ZN(n6607) );
  XNOR2_X1 U8414 ( .A(n8878), .B(n7118), .ZN(n8775) );
  OAI21_X1 U8415 ( .B1(n6609), .B2(n8775), .A(n6656), .ZN(n7120) );
  INV_X1 U8416 ( .A(n6658), .ZN(n6610) );
  AOI211_X1 U8417 ( .C1(n6660), .C2(n6611), .A(n9342), .B(n6610), .ZN(n7114)
         );
  NAND3_X1 U8418 ( .A1(n6614), .A2(n6613), .A3(n6612), .ZN(n6616) );
  INV_X1 U8419 ( .A(n8772), .ZN(n6615) );
  NAND2_X1 U8420 ( .A1(n8880), .A2(n6731), .ZN(n8817) );
  NAND3_X1 U8421 ( .A1(n6616), .A2(n6615), .A3(n8817), .ZN(n6619) );
  NAND2_X1 U8422 ( .A1(n6617), .A2(n6650), .ZN(n6618) );
  NAND2_X1 U8423 ( .A1(n6619), .A2(n6618), .ZN(n6659) );
  XNOR2_X1 U8424 ( .A(n6659), .B(n8775), .ZN(n6623) );
  OR2_X1 U8425 ( .A1(n6790), .A2(n9051), .ZN(n6621) );
  NAND2_X1 U8426 ( .A1(n8879), .A2(n9074), .ZN(n6620) );
  NAND2_X1 U8427 ( .A1(n6621), .A2(n6620), .ZN(n6737) );
  INV_X1 U8428 ( .A(n6737), .ZN(n6622) );
  OAI21_X1 U8429 ( .B1(n6623), .B2(n9240), .A(n6622), .ZN(n7113) );
  AOI211_X1 U8430 ( .C1(n9695), .C2(n7120), .A(n7114), .B(n7113), .ZN(n6690)
         );
  OAI22_X1 U8431 ( .A1(n9503), .A2(n7118), .B1(n9707), .B2(n4964), .ZN(n6624)
         );
  INV_X1 U8432 ( .A(n6624), .ZN(n6625) );
  OAI21_X1 U8433 ( .B1(n6690), .B2(n9706), .A(n6625), .ZN(P1_U3465) );
  INV_X1 U8434 ( .A(n8006), .ZN(n8016) );
  INV_X1 U8435 ( .A(n6626), .ZN(n6628) );
  INV_X1 U8436 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6627) );
  OAI222_X1 U8437 ( .A1(n8016), .A2(P2_U3151), .B1(n8451), .B2(n6628), .C1(
        n6627), .C2(n8449), .ZN(P2_U3280) );
  INV_X1 U8438 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6629) );
  OAI222_X1 U8439 ( .A1(n9522), .A2(n6629), .B1(n9514), .B2(n6628), .C1(
        P1_U3086), .C2(n9002), .ZN(P1_U3340) );
  INV_X1 U8440 ( .A(n6635), .ZN(n6633) );
  INV_X1 U8441 ( .A(n6630), .ZN(n6632) );
  OAI21_X1 U8442 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(n6701) );
  MUX2_X1 U8443 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4398), .Z(n6699) );
  XOR2_X1 U8444 ( .A(n6698), .B(n6699), .Z(n6700) );
  XNOR2_X1 U8445 ( .A(n6701), .B(n6700), .ZN(n6646) );
  INV_X1 U8446 ( .A(n6698), .ZN(n6644) );
  AOI21_X1 U8447 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6635), .A(n6634), .ZN(
        n6691) );
  XNOR2_X1 U8448 ( .A(n6691), .B(n6698), .ZN(n6693) );
  XOR2_X1 U8449 ( .A(n6693), .B(P2_REG1_REG_5__SCAN_IN), .Z(n6642) );
  OAI21_X1 U8450 ( .B1(n6637), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9873), .ZN(
        n6639) );
  INV_X1 U8451 ( .A(n8086), .ZN(n9874) );
  NOR2_X1 U8452 ( .A1(n6638), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6980) );
  AOI21_X1 U8453 ( .B1(n6639), .B2(n9874), .A(n6980), .ZN(n6641) );
  NAND2_X1 U8454 ( .A1(n9713), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6640) );
  OAI211_X1 U8455 ( .C1(n6642), .C2(n9891), .A(n6641), .B(n6640), .ZN(n6643)
         );
  AOI21_X1 U8456 ( .B1(n6644), .B2(n9882), .A(n6643), .ZN(n6645) );
  OAI21_X1 U8457 ( .B1(n8082), .B2(n6646), .A(n6645), .ZN(P2_U3187) );
  NOR2_X1 U8458 ( .A1(n7944), .A2(P2_U3151), .ZN(n6823) );
  AND2_X1 U8459 ( .A1(n7958), .A2(n6861), .ZN(n7558) );
  INV_X1 U8460 ( .A(n7558), .ZN(n7561) );
  AND2_X1 U8461 ( .A1(n7560), .A2(n7561), .ZN(n7502) );
  INV_X1 U8462 ( .A(n7502), .ZN(n6777) );
  OAI22_X1 U8463 ( .A1(n6264), .A2(n7942), .B1(n7947), .B2(n6861), .ZN(n6647)
         );
  AOI21_X1 U8464 ( .B1(n6777), .B2(n7934), .A(n6647), .ZN(n6648) );
  OAI21_X1 U8465 ( .B1(n6823), .B2(n6649), .A(n6648), .ZN(P2_U3172) );
  AOI22_X1 U8466 ( .A1(n9367), .A2(n6650), .B1(n9710), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6651) );
  OAI21_X1 U8467 ( .B1(n6652), .B2(n9710), .A(n6651), .ZN(P1_U3525) );
  OAI21_X1 U8468 ( .B1(n6654), .B2(n9710), .A(n6653), .ZN(P1_U3523) );
  INV_X1 U8469 ( .A(n8878), .ZN(n6661) );
  NAND2_X1 U8470 ( .A1(n6661), .A2(n7118), .ZN(n6655) );
  NAND2_X1 U8471 ( .A1(n6790), .A2(n6870), .ZN(n6788) );
  NAND2_X1 U8472 ( .A1(n6788), .A2(n8822), .ZN(n8774) );
  OAI21_X1 U8473 ( .B1(n6657), .B2(n8774), .A(n6783), .ZN(n7176) );
  AOI211_X1 U8474 ( .C1(n6870), .C2(n6658), .A(n9342), .B(n6786), .ZN(n7183)
         );
  NAND2_X1 U8475 ( .A1(n8878), .A2(n7118), .ZN(n8821) );
  NAND2_X1 U8476 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  XNOR2_X1 U8477 ( .A(n8630), .B(n8774), .ZN(n6665) );
  NAND2_X1 U8478 ( .A1(n8878), .A2(n9074), .ZN(n6664) );
  NAND2_X1 U8479 ( .A1(n8876), .A2(n8588), .ZN(n6663) );
  AND2_X1 U8480 ( .A1(n6664), .A2(n6663), .ZN(n6867) );
  OAI21_X1 U8481 ( .B1(n6665), .B2(n9240), .A(n6867), .ZN(n7177) );
  AOI211_X1 U8482 ( .C1(n9695), .C2(n7176), .A(n7183), .B(n7177), .ZN(n6669)
         );
  OAI22_X1 U8483 ( .A1(n9503), .A2(n7181), .B1(n9707), .B2(n5101), .ZN(n6666)
         );
  INV_X1 U8484 ( .A(n6666), .ZN(n6667) );
  OAI21_X1 U8485 ( .B1(n6669), .B2(n9706), .A(n6667), .ZN(P1_U3468) );
  AOI22_X1 U8486 ( .A1(n9367), .A2(n6870), .B1(n9710), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6668) );
  OAI21_X1 U8487 ( .B1(n6669), .B2(n9710), .A(n6668), .ZN(P1_U3527) );
  INV_X1 U8488 ( .A(n7940), .ZN(n7893) );
  OAI22_X1 U8489 ( .A1(n7893), .A2(n6264), .B1(n6807), .B2(n7947), .ZN(n6670)
         );
  AOI21_X1 U8490 ( .B1(n7925), .B2(n7957), .A(n6670), .ZN(n6676) );
  OAI21_X1 U8491 ( .B1(n6673), .B2(n6672), .A(n6671), .ZN(n6674) );
  NAND2_X1 U8492 ( .A1(n6674), .A2(n7934), .ZN(n6675) );
  OAI211_X1 U8493 ( .C1(n6823), .C2(n6521), .A(n6676), .B(n6675), .ZN(P2_U3177) );
  AOI22_X1 U8494 ( .A1(n9566), .A2(n6677), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n6678) );
  OAI21_X1 U8495 ( .B1(n9568), .B2(n8819), .A(n6678), .ZN(n6684) );
  OAI21_X1 U8496 ( .B1(n6681), .B2(n6680), .A(n6679), .ZN(n6682) );
  AND2_X1 U8497 ( .A1(n6682), .A2(n9571), .ZN(n6683) );
  AOI211_X1 U8498 ( .C1(n5071), .C2(n8568), .A(n6684), .B(n6683), .ZN(n6685)
         );
  INV_X1 U8499 ( .A(n6685), .ZN(P1_U3218) );
  INV_X1 U8500 ( .A(n6686), .ZN(n6714) );
  INV_X1 U8501 ( .A(n9013), .ZN(n9004) );
  OAI222_X1 U8502 ( .A1(n9514), .A2(n6714), .B1(n9004), .B2(P1_U3086), .C1(
        n6687), .C2(n9522), .ZN(P1_U3339) );
  OAI22_X1 U8503 ( .A1(n9440), .A2(n7118), .B1(n9712), .B2(n4965), .ZN(n6688)
         );
  INV_X1 U8504 ( .A(n6688), .ZN(n6689) );
  OAI21_X1 U8505 ( .B1(n6690), .B2(n9710), .A(n6689), .ZN(P1_U3526) );
  INV_X1 U8506 ( .A(n6691), .ZN(n6692) );
  INV_X1 U8507 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9826) );
  MUX2_X1 U8508 ( .A(n9826), .B(P2_REG1_REG_6__SCAN_IN), .S(n9871), .Z(n9870)
         );
  AOI21_X1 U8509 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n9871), .A(n9868), .ZN(
        n6746) );
  XNOR2_X1 U8510 ( .A(n6746), .B(n6747), .ZN(n6749) );
  XNOR2_X1 U8511 ( .A(n6749), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n6713) );
  INV_X1 U8512 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U8513 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7191) );
  OAI21_X1 U8514 ( .B1(n9880), .B2(n9916), .A(n7191), .ZN(n6697) );
  XNOR2_X1 U8515 ( .A(n9871), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n9872) );
  AOI21_X1 U8516 ( .B1(n6704), .B2(n6694), .A(n6753), .ZN(n6695) );
  NOR2_X1 U8517 ( .A1(n6695), .A2(n8086), .ZN(n6696) );
  AOI211_X1 U8518 ( .C1(n9882), .C2(n6747), .A(n6697), .B(n6696), .ZN(n6712)
         );
  AOI22_X1 U8519 ( .A1(n6701), .A2(n6700), .B1(n6699), .B2(n6698), .ZN(n9886)
         );
  MUX2_X1 U8520 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4398), .Z(n6702) );
  NOR2_X1 U8521 ( .A1(n6702), .A2(n9871), .ZN(n6703) );
  AOI21_X1 U8522 ( .B1(n6702), .B2(n9871), .A(n6703), .ZN(n9885) );
  NAND2_X1 U8523 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  INV_X1 U8524 ( .A(n6703), .ZN(n6709) );
  MUX2_X1 U8525 ( .A(n6704), .B(n6748), .S(n4398), .Z(n6705) );
  NAND2_X1 U8526 ( .A1(n6705), .A2(n6747), .ZN(n6763) );
  INV_X1 U8527 ( .A(n6705), .ZN(n6706) );
  NAND2_X1 U8528 ( .A1(n6706), .A2(n6754), .ZN(n6707) );
  NAND2_X1 U8529 ( .A1(n6763), .A2(n6707), .ZN(n6708) );
  AOI21_X1 U8530 ( .B1(n9884), .B2(n6709), .A(n6708), .ZN(n6772) );
  AND3_X1 U8531 ( .A1(n9884), .A2(n6709), .A3(n6708), .ZN(n6710) );
  OAI21_X1 U8532 ( .B1(n6772), .B2(n6710), .A(n9887), .ZN(n6711) );
  OAI211_X1 U8533 ( .C1(n6713), .C2(n9891), .A(n6712), .B(n6711), .ZN(P2_U3189) );
  OAI222_X1 U8534 ( .A1(n8449), .A2(n6715), .B1(P2_U3151), .B2(n8036), .C1(
        n6714), .C2(n8451), .ZN(P2_U3279) );
  INV_X1 U8535 ( .A(n9700), .ZN(n9686) );
  OR2_X1 U8536 ( .A1(n6716), .A2(n6724), .ZN(n6717) );
  NAND2_X1 U8537 ( .A1(n6718), .A2(n6717), .ZN(n9652) );
  NAND2_X1 U8538 ( .A1(n9656), .A2(n6719), .ZN(n6720) );
  NAND2_X1 U8539 ( .A1(n6720), .A2(n9216), .ZN(n6721) );
  NOR2_X1 U8540 ( .A1(n6722), .A2(n6721), .ZN(n9658) );
  INV_X1 U8541 ( .A(n6723), .ZN(n9705) );
  INV_X1 U8542 ( .A(n6724), .ZN(n8769) );
  XNOR2_X1 U8543 ( .A(n6725), .B(n8769), .ZN(n6726) );
  NOR2_X1 U8544 ( .A1(n6726), .A2(n9240), .ZN(n6727) );
  AOI211_X1 U8545 ( .C1(n9705), .C2(n9652), .A(n6728), .B(n6727), .ZN(n9666)
         );
  INV_X1 U8546 ( .A(n9666), .ZN(n6729) );
  AOI211_X1 U8547 ( .C1(n9686), .C2(n9652), .A(n9658), .B(n6729), .ZN(n6734)
         );
  AOI22_X1 U8548 ( .A1(n9367), .A2(n9656), .B1(n9710), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U8549 ( .B1(n6734), .B2(n9710), .A(n6730), .ZN(P1_U3524) );
  OAI22_X1 U8550 ( .A1(n9503), .A2(n6731), .B1(n9707), .B2(n5054), .ZN(n6732)
         );
  INV_X1 U8551 ( .A(n6732), .ZN(n6733) );
  OAI21_X1 U8552 ( .B1(n6734), .B2(n9706), .A(n6733), .ZN(P1_U3459) );
  INV_X1 U8553 ( .A(P1_U3973), .ZN(n8869) );
  NAND2_X1 U8554 ( .A1(n8869), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6735) );
  OAI21_X1 U8555 ( .B1(n9118), .B2(n8869), .A(n6735), .ZN(P1_U3581) );
  INV_X1 U8556 ( .A(n6736), .ZN(n7115) );
  NAND2_X1 U8557 ( .A1(n9566), .A2(n6737), .ZN(n6738) );
  OAI211_X1 U8558 ( .C1(n9568), .C2(n7118), .A(n6739), .B(n6738), .ZN(n6744)
         );
  AOI211_X1 U8559 ( .C1(n6742), .C2(n6741), .A(n8615), .B(n6740), .ZN(n6743)
         );
  AOI211_X1 U8560 ( .C1(n7115), .C2(n8568), .A(n6744), .B(n6743), .ZN(n6745)
         );
  INV_X1 U8561 ( .A(n6745), .ZN(P1_U3230) );
  OAI22_X1 U8562 ( .A1(n6749), .A2(n6748), .B1(n6747), .B2(n6746), .ZN(n6751)
         );
  AOI22_X1 U8563 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6844), .B1(n6766), .B2(
        n6764), .ZN(n6750) );
  OAI21_X1 U8564 ( .B1(n6751), .B2(n6750), .A(n6832), .ZN(n6762) );
  NAND2_X1 U8565 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6844), .ZN(n6755) );
  OAI21_X1 U8566 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6844), .A(n6755), .ZN(
        n6756) );
  AOI21_X1 U8567 ( .B1(n4379), .B2(n6756), .A(n6843), .ZN(n6760) );
  NOR2_X1 U8568 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6757), .ZN(n7318) );
  NOR2_X1 U8569 ( .A1(n8050), .A2(n6844), .ZN(n6758) );
  AOI211_X1 U8570 ( .C1(n9713), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7318), .B(
        n6758), .ZN(n6759) );
  OAI21_X1 U8571 ( .B1(n6760), .B2(n8086), .A(n6759), .ZN(n6761) );
  AOI21_X1 U8572 ( .B1(n9720), .B2(n6762), .A(n6761), .ZN(n6776) );
  INV_X1 U8573 ( .A(n6763), .ZN(n6771) );
  INV_X1 U8574 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6765) );
  MUX2_X1 U8575 ( .A(n6765), .B(n6764), .S(n4398), .Z(n6767) );
  NAND2_X1 U8576 ( .A1(n6767), .A2(n6766), .ZN(n6840) );
  INV_X1 U8577 ( .A(n6767), .ZN(n6768) );
  NAND2_X1 U8578 ( .A1(n6768), .A2(n6844), .ZN(n6769) );
  AND2_X1 U8579 ( .A1(n6840), .A2(n6769), .ZN(n6770) );
  OAI21_X1 U8580 ( .B1(n6772), .B2(n6771), .A(n6770), .ZN(n6841) );
  INV_X1 U8581 ( .A(n6841), .ZN(n6774) );
  NOR3_X1 U8582 ( .A1(n6772), .A2(n6771), .A3(n6770), .ZN(n6773) );
  OAI21_X1 U8583 ( .B1(n6774), .B2(n6773), .A(n9887), .ZN(n6775) );
  NAND2_X1 U8584 ( .A1(n6776), .A2(n6775), .ZN(P2_U3190) );
  INV_X1 U8585 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6781) );
  OAI21_X1 U8586 ( .B1(n9748), .B2(n9811), .A(n6777), .ZN(n6779) );
  NOR2_X1 U8587 ( .A1(n6264), .A2(n9550), .ZN(n6857) );
  INV_X1 U8588 ( .A(n6857), .ZN(n6778) );
  OAI211_X1 U8589 ( .C1(n9793), .C2(n6861), .A(n6779), .B(n6778), .ZN(n8359)
         );
  NAND2_X1 U8590 ( .A1(n8359), .A2(n9817), .ZN(n6780) );
  OAI21_X1 U8591 ( .B1(n6781), .B2(n9817), .A(n6780), .ZN(P2_U3390) );
  NAND2_X1 U8592 ( .A1(n6790), .A2(n7181), .ZN(n6782) );
  NAND2_X1 U8593 ( .A1(n6783), .A2(n6782), .ZN(n6785) );
  NAND2_X1 U8594 ( .A1(n7167), .A2(n8876), .ZN(n8634) );
  INV_X1 U8595 ( .A(n8876), .ZN(n6784) );
  NAND2_X1 U8596 ( .A1(n8634), .A2(n8628), .ZN(n6789) );
  OAI21_X1 U8597 ( .B1(n6785), .B2(n6789), .A(n6926), .ZN(n7172) );
  INV_X1 U8598 ( .A(n6786), .ZN(n6787) );
  AOI211_X1 U8599 ( .C1(n6924), .C2(n6787), .A(n9342), .B(n6942), .ZN(n7171)
         );
  INV_X1 U8600 ( .A(n6788), .ZN(n8629) );
  INV_X1 U8601 ( .A(n6789), .ZN(n8778) );
  XNOR2_X1 U8602 ( .A(n8632), .B(n8778), .ZN(n6793) );
  OR2_X1 U8603 ( .A1(n6790), .A2(n8508), .ZN(n6791) );
  OAI21_X1 U8604 ( .B1(n7133), .B2(n9051), .A(n6791), .ZN(n6969) );
  INV_X1 U8605 ( .A(n6969), .ZN(n6792) );
  OAI21_X1 U8606 ( .B1(n6793), .B2(n9240), .A(n6792), .ZN(n7166) );
  AOI211_X1 U8607 ( .C1(n9695), .C2(n7172), .A(n7171), .B(n7166), .ZN(n6797)
         );
  OAI22_X1 U8608 ( .A1(n9503), .A2(n7167), .B1(n9707), .B2(n5130), .ZN(n6794)
         );
  INV_X1 U8609 ( .A(n6794), .ZN(n6795) );
  OAI21_X1 U8610 ( .B1(n6797), .B2(n9706), .A(n6795), .ZN(P1_U3471) );
  AOI22_X1 U8611 ( .A1(n9367), .A2(n6924), .B1(n9710), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6796) );
  OAI21_X1 U8612 ( .B1(n6797), .B2(n9710), .A(n6796), .ZN(P1_U3528) );
  NOR2_X1 U8613 ( .A1(n6799), .A2(n4421), .ZN(n6800) );
  NOR2_X1 U8614 ( .A1(n6801), .A2(n6800), .ZN(n6803) );
  NAND3_X1 U8615 ( .A1(n6804), .A2(n6803), .A3(n6802), .ZN(n6854) );
  NOR2_X1 U8616 ( .A1(n6805), .A2(n8065), .ZN(n7366) );
  OR2_X1 U8617 ( .A1(n9786), .A2(n7366), .ZN(n9552) );
  XNOR2_X1 U8618 ( .A(n6806), .B(n5833), .ZN(n8353) );
  INV_X1 U8619 ( .A(n8353), .ZN(n6816) );
  NOR2_X1 U8620 ( .A1(n6807), .A2(n8278), .ZN(n6813) );
  XNOR2_X1 U8621 ( .A(n6808), .B(n5833), .ZN(n6811) );
  NAND2_X1 U8622 ( .A1(n7957), .A2(n9745), .ZN(n6809) );
  OAI21_X1 U8623 ( .B1(n6264), .B2(n9548), .A(n6809), .ZN(n6810) );
  AOI21_X1 U8624 ( .B1(n6811), .B2(n9748), .A(n6810), .ZN(n8357) );
  INV_X1 U8625 ( .A(n8357), .ZN(n6812) );
  AOI211_X1 U8626 ( .C1(n9752), .C2(P2_REG3_REG_2__SCAN_IN), .A(n6813), .B(
        n6812), .ZN(n6814) );
  MUX2_X1 U8627 ( .A(n4578), .B(n6814), .S(n8268), .Z(n6815) );
  OAI21_X1 U8628 ( .B1(n8272), .B2(n6816), .A(n6815), .ZN(P2_U3231) );
  INV_X1 U8629 ( .A(n6817), .ZN(n6821) );
  INV_X1 U8630 ( .A(n6819), .ZN(n6820) );
  AOI21_X1 U8631 ( .B1(n6821), .B2(n6818), .A(n6820), .ZN(n6827) );
  OAI22_X1 U8632 ( .A1(n7893), .A2(n6822), .B1(n7947), .B2(n7024), .ZN(n6825)
         );
  NOR2_X1 U8633 ( .A1(n6823), .A2(n7023), .ZN(n6824) );
  AOI211_X1 U8634 ( .C1(n7925), .C2(n9744), .A(n6825), .B(n6824), .ZN(n6826)
         );
  OAI21_X1 U8635 ( .B1(n7932), .B2(n6827), .A(n6826), .ZN(P2_U3162) );
  INV_X1 U8636 ( .A(n6828), .ZN(n6831) );
  INV_X1 U8637 ( .A(n9031), .ZN(n9017) );
  OAI222_X1 U8638 ( .A1(n9522), .A2(n6829), .B1(n9514), .B2(n6831), .C1(
        P1_U3086), .C2(n9017), .ZN(P1_U3338) );
  INV_X1 U8639 ( .A(n9714), .ZN(n8038) );
  OAI222_X1 U8640 ( .A1(n8038), .A2(P2_U3151), .B1(n8451), .B2(n6831), .C1(
        n6830), .C2(n8449), .ZN(P2_U3278) );
  NAND2_X1 U8641 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6844), .ZN(n6833) );
  XNOR2_X1 U8642 ( .A(n7050), .B(n6850), .ZN(n7051) );
  INV_X1 U8643 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U8644 ( .A(n7051), .B(n6834), .ZN(n6853) );
  MUX2_X1 U8645 ( .A(n6835), .B(n6834), .S(n4398), .Z(n6836) );
  NAND2_X1 U8646 ( .A1(n6836), .A2(n6850), .ZN(n7039) );
  INV_X1 U8647 ( .A(n6836), .ZN(n6837) );
  NAND2_X1 U8648 ( .A1(n6837), .A2(n4555), .ZN(n6838) );
  NAND2_X1 U8649 ( .A1(n7039), .A2(n6838), .ZN(n6839) );
  AOI21_X1 U8650 ( .B1(n6841), .B2(n6840), .A(n6839), .ZN(n7047) );
  AND3_X1 U8651 ( .A1(n6841), .A2(n6840), .A3(n6839), .ZN(n6842) );
  OAI21_X1 U8652 ( .B1(n7047), .B2(n6842), .A(n9887), .ZN(n6852) );
  AOI21_X1 U8653 ( .B1(n6835), .B2(n6845), .A(n7055), .ZN(n6847) );
  OAI21_X1 U8654 ( .B1(n8086), .B2(n6847), .A(n6846), .ZN(n6849) );
  INV_X1 U8655 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9991) );
  NOR2_X1 U8656 ( .A1(n9880), .A2(n9991), .ZN(n6848) );
  AOI211_X1 U8657 ( .C1(n9882), .C2(n6850), .A(n6849), .B(n6848), .ZN(n6851)
         );
  OAI211_X1 U8658 ( .C1(n9891), .C2(n6853), .A(n6852), .B(n6851), .ZN(P2_U3191) );
  NOR3_X1 U8659 ( .A1(n7502), .A2(n6855), .A3(n9816), .ZN(n6856) );
  AOI211_X1 U8660 ( .C1(n9752), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6857), .B(
        n6856), .ZN(n6858) );
  MUX2_X1 U8661 ( .A(n6859), .B(n6858), .S(n8268), .Z(n6860) );
  OAI21_X1 U8662 ( .B1(n8095), .B2(n6861), .A(n6860), .ZN(P2_U3233) );
  INV_X1 U8663 ( .A(n6862), .ZN(n6949) );
  AOI22_X1 U8664 ( .A1(n8072), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8446), .ZN(n6863) );
  OAI21_X1 U8665 ( .B1(n6949), .B2(n8451), .A(n6863), .ZN(P2_U3277) );
  AOI21_X1 U8666 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n6872) );
  NAND2_X1 U8667 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n8923) );
  OAI21_X1 U8668 ( .B1(n8601), .B2(n6867), .A(n8923), .ZN(n6869) );
  NOR2_X1 U8669 ( .A1(n9575), .A2(n7180), .ZN(n6868) );
  AOI211_X1 U8670 ( .C1(n6870), .C2(n8613), .A(n6869), .B(n6868), .ZN(n6871)
         );
  OAI21_X1 U8671 ( .B1(n6872), .B2(n8615), .A(n6871), .ZN(P1_U3227) );
  INV_X2 U8672 ( .A(P2_U3893), .ZN(n8051) );
  NAND2_X1 U8673 ( .A1(n8051), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6873) );
  OAI21_X1 U8674 ( .B1(n7495), .B2(n8051), .A(n6873), .ZN(P2_U3521) );
  INV_X1 U8675 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9841) );
  NOR2_X1 U8676 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6874) );
  AOI21_X1 U8677 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6874), .ZN(n9846) );
  NOR2_X1 U8678 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6875) );
  AOI21_X1 U8679 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6875), .ZN(n9849) );
  NOR2_X1 U8680 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6876) );
  AOI21_X1 U8681 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6876), .ZN(n9852) );
  NOR2_X1 U8682 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6877) );
  AOI21_X1 U8683 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6877), .ZN(n9855) );
  NOR2_X1 U8684 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6878) );
  AOI21_X1 U8685 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6878), .ZN(n9858) );
  NOR2_X1 U8686 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6879) );
  AOI21_X1 U8687 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6879), .ZN(n9861) );
  NOR2_X1 U8688 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6880) );
  AOI21_X1 U8689 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6880), .ZN(n9864) );
  NOR2_X1 U8690 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6881) );
  AOI21_X1 U8691 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6881), .ZN(n9867) );
  NOR2_X1 U8692 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6882) );
  AOI21_X1 U8693 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6882), .ZN(n10050) );
  NOR2_X1 U8694 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6883) );
  AOI21_X1 U8695 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6883), .ZN(n10056) );
  NOR2_X1 U8696 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6884) );
  AOI21_X1 U8697 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6884), .ZN(n10053) );
  NOR2_X1 U8698 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6885) );
  AOI21_X1 U8699 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6885), .ZN(n10044) );
  NOR2_X1 U8700 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6886) );
  AOI21_X1 U8701 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6886), .ZN(n10047) );
  AND2_X1 U8702 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6887) );
  NOR2_X1 U8703 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6887), .ZN(n9836) );
  INV_X1 U8704 ( .A(n9836), .ZN(n9837) );
  NAND3_X1 U8705 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U8706 ( .A1(n9839), .A2(n9838), .ZN(n9835) );
  NAND2_X1 U8707 ( .A1(n9837), .A2(n9835), .ZN(n10059) );
  NAND2_X1 U8708 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6888) );
  OAI21_X1 U8709 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6888), .ZN(n10058) );
  NOR2_X1 U8710 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  AOI21_X1 U8711 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10057), .ZN(n10062) );
  NAND2_X1 U8712 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6889) );
  OAI21_X1 U8713 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6889), .ZN(n10061) );
  NOR2_X1 U8714 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  AOI21_X1 U8715 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10060), .ZN(n10065) );
  NOR2_X1 U8716 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6890) );
  AOI21_X1 U8717 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6890), .ZN(n10064) );
  NAND2_X1 U8718 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  OAI21_X1 U8719 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10063), .ZN(n10046) );
  NAND2_X1 U8720 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  OAI21_X1 U8721 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10045), .ZN(n10043) );
  NAND2_X1 U8722 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  OAI21_X1 U8723 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10042), .ZN(n10052) );
  NAND2_X1 U8724 ( .A1(n10053), .A2(n10052), .ZN(n10051) );
  OAI21_X1 U8725 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10051), .ZN(n10055) );
  NAND2_X1 U8726 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  OAI21_X1 U8727 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10054), .ZN(n10049) );
  NAND2_X1 U8728 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  OAI21_X1 U8729 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10048), .ZN(n9866) );
  NAND2_X1 U8730 ( .A1(n9867), .A2(n9866), .ZN(n9865) );
  OAI21_X1 U8731 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9865), .ZN(n9863) );
  NAND2_X1 U8732 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  OAI21_X1 U8733 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9862), .ZN(n9860) );
  NAND2_X1 U8734 ( .A1(n9861), .A2(n9860), .ZN(n9859) );
  OAI21_X1 U8735 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9859), .ZN(n9857) );
  NAND2_X1 U8736 ( .A1(n9858), .A2(n9857), .ZN(n9856) );
  OAI21_X1 U8737 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9856), .ZN(n9854) );
  NAND2_X1 U8738 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  OAI21_X1 U8739 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9853), .ZN(n9851) );
  NAND2_X1 U8740 ( .A1(n9852), .A2(n9851), .ZN(n9850) );
  OAI21_X1 U8741 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9850), .ZN(n9848) );
  NAND2_X1 U8742 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  OAI21_X1 U8743 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9847), .ZN(n9845) );
  NAND2_X1 U8744 ( .A1(n9846), .A2(n9845), .ZN(n9844) );
  OAI21_X1 U8745 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9844), .ZN(n9842) );
  NAND2_X1 U8746 ( .A1(n9841), .A2(n9842), .ZN(n6891) );
  NOR2_X1 U8747 ( .A1(n9841), .A2(n9842), .ZN(n9840) );
  AOI21_X1 U8748 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6891), .A(n9840), .ZN(
        n6893) );
  XNOR2_X1 U8749 ( .A(n9045), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n6892) );
  XNOR2_X1 U8750 ( .A(n6893), .B(n6892), .ZN(ADD_1068_U4) );
  INV_X1 U8751 ( .A(n9630), .ZN(n9646) );
  MUX2_X1 U8752 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n5268), .S(n9579), .Z(n9578)
         );
  NAND2_X1 U8753 ( .A1(n9534), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6902) );
  OAI21_X1 U8754 ( .B1(n9534), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6902), .ZN(
        n9530) );
  MUX2_X1 U8755 ( .A(n6896), .B(P1_REG1_REG_5__SCAN_IN), .S(n8926), .Z(n8920)
         );
  NOR2_X1 U8756 ( .A1(n8921), .A2(n8920), .ZN(n8919) );
  MUX2_X1 U8757 ( .A(n6897), .B(P1_REG1_REG_6__SCAN_IN), .S(n8940), .Z(n8934)
         );
  NOR2_X1 U8758 ( .A1(n8935), .A2(n8934), .ZN(n8933) );
  MUX2_X1 U8759 ( .A(n6898), .B(P1_REG1_REG_7__SCAN_IN), .S(n8954), .Z(n8948)
         );
  MUX2_X1 U8760 ( .A(n6899), .B(P1_REG1_REG_8__SCAN_IN), .S(n8968), .Z(n8962)
         );
  NOR2_X1 U8761 ( .A1(n8963), .A2(n8962), .ZN(n8961) );
  NOR2_X1 U8762 ( .A1(n8984), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6900) );
  AOI21_X1 U8763 ( .B1(n8984), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6900), .ZN(
        n8977) );
  NAND2_X1 U8764 ( .A1(n8976), .A2(n8977), .ZN(n8975) );
  OAI21_X1 U8765 ( .B1(n8984), .B2(P1_REG1_REG_9__SCAN_IN), .A(n8975), .ZN(
        n9531) );
  NAND2_X1 U8766 ( .A1(n6902), .A2(n6901), .ZN(n9577) );
  AOI22_X1 U8767 ( .A1(n8999), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5288), .B2(
        n6923), .ZN(n6903) );
  NAND2_X1 U8768 ( .A1(n4329), .A2(n6903), .ZN(n8989) );
  OAI21_X1 U8769 ( .B1(n4329), .B2(n6903), .A(n8989), .ZN(n6919) );
  AOI22_X1 U8770 ( .A1(n8999), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7305), .B2(
        n6923), .ZN(n6917) );
  MUX2_X1 U8771 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7259), .S(n9579), .Z(n9582)
         );
  NAND2_X1 U8772 ( .A1(n9534), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6904) );
  OAI21_X1 U8773 ( .B1(n9534), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6904), .ZN(
        n9527) );
  INV_X1 U8774 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6909) );
  OAI21_X1 U8775 ( .B1(n6907), .B2(n6906), .A(n6905), .ZN(n8928) );
  MUX2_X1 U8776 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7179), .S(n8926), .Z(n8929)
         );
  NAND2_X1 U8777 ( .A1(n8928), .A2(n8929), .ZN(n8927) );
  OAI21_X1 U8778 ( .B1(n6908), .B2(n7179), .A(n8927), .ZN(n8942) );
  MUX2_X1 U8779 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6909), .S(n8940), .Z(n8943)
         );
  NAND2_X1 U8780 ( .A1(n8942), .A2(n8943), .ZN(n8941) );
  OAI21_X1 U8781 ( .B1(n6910), .B2(n6909), .A(n8941), .ZN(n8956) );
  MUX2_X1 U8782 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6944), .S(n8954), .Z(n8957)
         );
  NAND2_X1 U8783 ( .A1(n8956), .A2(n8957), .ZN(n8955) );
  OAI21_X1 U8784 ( .B1(n6944), .B2(n6911), .A(n8955), .ZN(n8970) );
  MUX2_X1 U8785 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7006), .S(n8968), .Z(n8971)
         );
  NAND2_X1 U8786 ( .A1(n8970), .A2(n8971), .ZN(n8969) );
  INV_X1 U8787 ( .A(n8969), .ZN(n6912) );
  AOI21_X1 U8788 ( .B1(n8968), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6912), .ZN(
        n8981) );
  NOR2_X1 U8789 ( .A1(n8984), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6913) );
  AOI21_X1 U8790 ( .B1(n8984), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6913), .ZN(
        n8982) );
  NAND2_X1 U8791 ( .A1(n8981), .A2(n8982), .ZN(n8980) );
  OAI21_X1 U8792 ( .B1(n8984), .B2(P1_REG2_REG_9__SCAN_IN), .A(n8980), .ZN(
        n9528) );
  NOR2_X1 U8793 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  AOI21_X1 U8794 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9534), .A(n9526), .ZN(
        n6914) );
  INV_X1 U8795 ( .A(n6914), .ZN(n9581) );
  NAND2_X1 U8796 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  NAND2_X1 U8797 ( .A1(n9579), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6915) );
  AND2_X1 U8798 ( .A1(n9580), .A2(n6915), .ZN(n6916) );
  NAND2_X1 U8799 ( .A1(n6917), .A2(n6916), .ZN(n8998) );
  OAI21_X1 U8800 ( .B1(n6917), .B2(n6916), .A(n8998), .ZN(n6918) );
  AOI22_X1 U8801 ( .A1(n9634), .A2(n6919), .B1(n9642), .B2(n6918), .ZN(n6922)
         );
  NOR2_X1 U8802 ( .A1(n6920), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8497) );
  AOI21_X1 U8803 ( .B1(n9014), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8497), .ZN(
        n6921) );
  OAI211_X1 U8804 ( .C1(n6923), .C2(n9646), .A(n6922), .B(n6921), .ZN(P1_U3255) );
  OR2_X1 U8805 ( .A1(n8876), .A2(n6924), .ZN(n6925) );
  NAND2_X1 U8806 ( .A1(n6926), .A2(n6925), .ZN(n6927) );
  XNOR2_X1 U8807 ( .A(n7134), .B(n7133), .ZN(n8642) );
  OR2_X1 U8808 ( .A1(n6927), .A2(n8642), .ZN(n6928) );
  NAND2_X1 U8809 ( .A1(n6994), .A2(n6928), .ZN(n9687) );
  NAND2_X1 U8810 ( .A1(n9687), .A2(n9705), .ZN(n6935) );
  NAND2_X1 U8811 ( .A1(n7132), .A2(n8634), .ZN(n6929) );
  NOR2_X1 U8812 ( .A1(n6929), .A2(n8642), .ZN(n7151) );
  AND2_X1 U8813 ( .A1(n6929), .A2(n8642), .ZN(n6930) );
  OR2_X1 U8814 ( .A1(n7151), .A2(n6930), .ZN(n6933) );
  OR2_X1 U8815 ( .A1(n7153), .A2(n9051), .ZN(n6932) );
  NAND2_X1 U8816 ( .A1(n8876), .A2(n9074), .ZN(n6931) );
  NAND2_X1 U8817 ( .A1(n6932), .A2(n6931), .ZN(n7036) );
  AOI21_X1 U8818 ( .B1(n6933), .B2(n9333), .A(n7036), .ZN(n6934) );
  NAND3_X1 U8819 ( .A1(n6938), .A2(n6937), .A3(n6936), .ZN(n6939) );
  INV_X1 U8820 ( .A(n6940), .ZN(n6941) );
  AND2_X1 U8821 ( .A1(n9678), .A2(n6941), .ZN(n9651) );
  NAND2_X1 U8822 ( .A1(n6942), .A2(n9684), .ZN(n7005) );
  OAI211_X1 U8823 ( .C1(n6942), .C2(n9684), .A(n9216), .B(n7005), .ZN(n9683)
         );
  NAND2_X1 U8824 ( .A1(n9678), .A2(n8810), .ZN(n9660) );
  OAI22_X1 U8825 ( .A1(n9678), .A2(n6944), .B1(n7033), .B2(n9673), .ZN(n6945)
         );
  AOI21_X1 U8826 ( .B1(n9657), .B2(n7134), .A(n6945), .ZN(n6946) );
  OAI21_X1 U8827 ( .B1(n9683), .B2(n9660), .A(n6946), .ZN(n6947) );
  AOI21_X1 U8828 ( .B1(n9687), .B2(n9651), .A(n6947), .ZN(n6948) );
  OAI21_X1 U8829 ( .B1(n9689), .B2(n9304), .A(n6948), .ZN(P1_U3286) );
  INV_X1 U8830 ( .A(n9028), .ZN(n9645) );
  OAI222_X1 U8831 ( .A1(n9522), .A2(n6950), .B1(n9645), .B2(P1_U3086), .C1(
        n9514), .C2(n6949), .ZN(P1_U3337) );
  XNOR2_X1 U8832 ( .A(n6115), .B(n6951), .ZN(n6952) );
  NAND2_X1 U8833 ( .A1(n6952), .A2(n9748), .ZN(n6954) );
  AOI22_X1 U8834 ( .A1(n9743), .A2(n7958), .B1(n9744), .B2(n9745), .ZN(n6953)
         );
  AND2_X1 U8835 ( .A1(n6954), .A2(n6953), .ZN(n7022) );
  NAND2_X1 U8836 ( .A1(n6115), .A2(n7560), .ZN(n6955) );
  AOI22_X1 U8837 ( .A1(n7026), .A2(n8354), .B1(n6956), .B2(n9816), .ZN(n6958)
         );
  NAND2_X1 U8838 ( .A1(n7026), .A2(n9786), .ZN(n6957) );
  AND3_X1 U8839 ( .A1(n7022), .A2(n6958), .A3(n6957), .ZN(n9758) );
  MUX2_X1 U8840 ( .A(n6959), .B(n9758), .S(n4275), .Z(n6960) );
  INV_X1 U8841 ( .A(n6960), .ZN(P2_U3460) );
  INV_X1 U8842 ( .A(n6961), .ZN(n6965) );
  NOR3_X1 U8843 ( .A1(n6864), .A2(n6963), .A3(n6962), .ZN(n6964) );
  OAI21_X1 U8844 ( .B1(n6965), .B2(n6964), .A(n9571), .ZN(n6971) );
  NAND2_X1 U8845 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8937) );
  INV_X1 U8846 ( .A(n8937), .ZN(n6968) );
  INV_X1 U8847 ( .A(n6966), .ZN(n7168) );
  NOR2_X1 U8848 ( .A1(n9575), .A2(n7168), .ZN(n6967) );
  AOI211_X1 U8849 ( .C1(n9566), .C2(n6969), .A(n6968), .B(n6967), .ZN(n6970)
         );
  OAI211_X1 U8850 ( .C1(n7167), .C2(n9568), .A(n6971), .B(n6970), .ZN(P1_U3239) );
  INV_X1 U8851 ( .A(n6972), .ZN(n6976) );
  INV_X1 U8852 ( .A(n6973), .ZN(n6975) );
  NOR3_X1 U8853 ( .A1(n6976), .A2(n6975), .A3(n6974), .ZN(n6979) );
  INV_X1 U8854 ( .A(n6977), .ZN(n6978) );
  OAI21_X1 U8855 ( .B1(n6979), .B2(n6978), .A(n7934), .ZN(n6985) );
  AOI21_X1 U8856 ( .B1(n7925), .B2(n7955), .A(n6980), .ZN(n6981) );
  OAI21_X1 U8857 ( .B1(n6982), .B2(n7893), .A(n6981), .ZN(n6983) );
  AOI21_X1 U8858 ( .B1(n7094), .B2(n7930), .A(n6983), .ZN(n6984) );
  OAI211_X1 U8859 ( .C1(n7092), .C2(n7928), .A(n6985), .B(n6984), .ZN(P2_U3167) );
  AOI21_X1 U8860 ( .B1(n9705), .B2(n9678), .A(n9651), .ZN(n7418) );
  INV_X1 U8861 ( .A(n6986), .ZN(n6993) );
  OAI22_X1 U8862 ( .A1(n9345), .A2(n8814), .B1(n4397), .B2(n9673), .ZN(n6987)
         );
  AOI21_X1 U8863 ( .B1(n9350), .B2(n6988), .A(n6987), .ZN(n6992) );
  INV_X1 U8864 ( .A(n6989), .ZN(n6990) );
  MUX2_X1 U8865 ( .A(n6405), .B(n6990), .S(n9678), .Z(n6991) );
  OAI211_X1 U8866 ( .C1(n7418), .C2(n6993), .A(n6992), .B(n6991), .ZN(P1_U3292) );
  INV_X1 U8867 ( .A(n7133), .ZN(n8875) );
  NAND2_X1 U8868 ( .A1(n7139), .A2(n7153), .ZN(n8644) );
  NAND2_X1 U8869 ( .A1(n8645), .A2(n8644), .ZN(n7001) );
  NAND2_X1 U8870 ( .A1(n6995), .A2(n7001), .ZN(n7141) );
  OAI21_X1 U8871 ( .B1(n6995), .B2(n7001), .A(n7141), .ZN(n7016) );
  INV_X1 U8872 ( .A(n7016), .ZN(n7011) );
  INV_X1 U8873 ( .A(n7151), .ZN(n6996) );
  NAND2_X1 U8874 ( .A1(n7134), .A2(n7133), .ZN(n6997) );
  NAND2_X1 U8875 ( .A1(n6996), .A2(n6997), .ZN(n7000) );
  INV_X1 U8876 ( .A(n8645), .ZN(n6998) );
  NAND2_X1 U8877 ( .A1(n8644), .A2(n6997), .ZN(n8638) );
  NOR3_X1 U8878 ( .A1(n7151), .A2(n6998), .A3(n8638), .ZN(n6999) );
  AOI211_X1 U8879 ( .C1(n7001), .C2(n7000), .A(n9240), .B(n6999), .ZN(n7003)
         );
  OR2_X1 U8880 ( .A1(n7133), .A2(n8508), .ZN(n7002) );
  OAI21_X1 U8881 ( .B1(n7142), .B2(n9051), .A(n7002), .ZN(n7285) );
  OR2_X1 U8882 ( .A1(n7003), .A2(n7285), .ZN(n7014) );
  NAND2_X1 U8883 ( .A1(n7014), .A2(n9678), .ZN(n7010) );
  OR2_X1 U8884 ( .A1(n7005), .A2(n7139), .ZN(n7157) );
  INV_X1 U8885 ( .A(n7157), .ZN(n7004) );
  AOI211_X1 U8886 ( .C1(n7139), .C2(n7005), .A(n9342), .B(n7004), .ZN(n7015)
         );
  NOR2_X1 U8887 ( .A1(n9345), .A2(n4650), .ZN(n7008) );
  OAI22_X1 U8888 ( .A1(n9678), .A2(n7006), .B1(n7282), .B2(n9673), .ZN(n7007)
         );
  AOI211_X1 U8889 ( .C1(n7015), .C2(n9350), .A(n7008), .B(n7007), .ZN(n7009)
         );
  OAI211_X1 U8890 ( .C1(n7418), .C2(n7011), .A(n7010), .B(n7009), .ZN(P1_U3285) );
  INV_X1 U8891 ( .A(n7012), .ZN(n7716) );
  OAI222_X1 U8892 ( .A1(P2_U3151), .A2(n8065), .B1(n8451), .B2(n7716), .C1(
        n7013), .C2(n8449), .ZN(P2_U3276) );
  AOI211_X1 U8893 ( .C1(n9695), .C2(n7016), .A(n7015), .B(n7014), .ZN(n7020)
         );
  AOI22_X1 U8894 ( .A1(n9367), .A2(n7139), .B1(n9710), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7017) );
  OAI21_X1 U8895 ( .B1(n7020), .B2(n9710), .A(n7017), .ZN(P1_U3530) );
  OAI22_X1 U8896 ( .A1(n9503), .A2(n4650), .B1(n9707), .B2(n5185), .ZN(n7018)
         );
  INV_X1 U8897 ( .A(n7018), .ZN(n7019) );
  OAI21_X1 U8898 ( .B1(n7020), .B2(n9706), .A(n7019), .ZN(P1_U3477) );
  MUX2_X1 U8899 ( .A(n7022), .B(n7021), .S(n9757), .Z(n7028) );
  OAI22_X1 U8900 ( .A1(n8095), .A2(n7024), .B1(n7023), .B2(n9540), .ZN(n7025)
         );
  AOI21_X1 U8901 ( .B1(n9754), .B2(n7026), .A(n7025), .ZN(n7027) );
  NAND2_X1 U8902 ( .A1(n7028), .A2(n7027), .ZN(P2_U3232) );
  OAI21_X1 U8903 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7032) );
  NAND2_X1 U8904 ( .A1(n7032), .A2(n9571), .ZN(n7038) );
  NAND2_X1 U8905 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n8951) );
  INV_X1 U8906 ( .A(n8951), .ZN(n7035) );
  NOR2_X1 U8907 ( .A1(n9575), .A2(n7033), .ZN(n7034) );
  AOI211_X1 U8908 ( .C1(n9566), .C2(n7036), .A(n7035), .B(n7034), .ZN(n7037)
         );
  OAI211_X1 U8909 ( .C1(n9684), .C2(n9568), .A(n7038), .B(n7037), .ZN(P1_U3213) );
  INV_X1 U8910 ( .A(n7039), .ZN(n7046) );
  MUX2_X1 U8911 ( .A(n7041), .B(n7040), .S(n4398), .Z(n7042) );
  NAND2_X1 U8912 ( .A1(n7042), .A2(n7079), .ZN(n7075) );
  INV_X1 U8913 ( .A(n7042), .ZN(n7043) );
  NAND2_X1 U8914 ( .A1(n7043), .A2(n7067), .ZN(n7044) );
  AND2_X1 U8915 ( .A1(n7075), .A2(n7044), .ZN(n7045) );
  OAI21_X1 U8916 ( .B1(n7047), .B2(n7046), .A(n7045), .ZN(n7076) );
  INV_X1 U8917 ( .A(n7076), .ZN(n7049) );
  NOR3_X1 U8918 ( .A1(n7047), .A2(n7046), .A3(n7045), .ZN(n7048) );
  OAI21_X1 U8919 ( .B1(n7049), .B2(n7048), .A(n9887), .ZN(n7065) );
  AOI22_X1 U8920 ( .A1(n7051), .A2(P2_REG1_REG_9__SCAN_IN), .B1(n7050), .B2(
        n4555), .ZN(n7052) );
  INV_X1 U8921 ( .A(n7052), .ZN(n7054) );
  AOI22_X1 U8922 ( .A1(n7079), .A2(n7040), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7067), .ZN(n7053) );
  OAI21_X1 U8923 ( .B1(n7054), .B2(n7053), .A(n7078), .ZN(n7063) );
  AOI22_X1 U8924 ( .A1(n7079), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7041), .B2(
        n7067), .ZN(n7056) );
  AOI21_X1 U8925 ( .B1(n7057), .B2(n7056), .A(n7066), .ZN(n7059) );
  INV_X1 U8926 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7058) );
  OR2_X1 U8927 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7058), .ZN(n7461) );
  OAI21_X1 U8928 ( .B1(n8086), .B2(n7059), .A(n7461), .ZN(n7060) );
  AOI21_X1 U8929 ( .B1(n9713), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7060), .ZN(
        n7061) );
  OAI21_X1 U8930 ( .B1(n8050), .B2(n7067), .A(n7061), .ZN(n7062) );
  AOI21_X1 U8931 ( .B1(n7063), .B2(n9720), .A(n7062), .ZN(n7064) );
  NAND2_X1 U8932 ( .A1(n7065), .A2(n7064), .ZN(P2_U3192) );
  AOI21_X1 U8933 ( .B1(n7070), .B2(n7068), .A(n7209), .ZN(n7086) );
  MUX2_X1 U8934 ( .A(n7070), .B(n7069), .S(n4398), .Z(n7071) );
  NAND2_X1 U8935 ( .A1(n7071), .A2(n7208), .ZN(n7214) );
  INV_X1 U8936 ( .A(n7071), .ZN(n7072) );
  NAND2_X1 U8937 ( .A1(n7072), .A2(n4773), .ZN(n7073) );
  NAND2_X1 U8938 ( .A1(n7214), .A2(n7073), .ZN(n7074) );
  AOI21_X1 U8939 ( .B1(n7076), .B2(n7075), .A(n7074), .ZN(n7221) );
  AND3_X1 U8940 ( .A1(n7076), .A2(n7075), .A3(n7074), .ZN(n7077) );
  OAI21_X1 U8941 ( .B1(n7221), .B2(n7077), .A(n9887), .ZN(n7085) );
  OAI21_X1 U8942 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7080), .A(n7225), .ZN(
        n7083) );
  AND2_X1 U8943 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7900) );
  AOI21_X1 U8944 ( .B1(n9713), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7900), .ZN(
        n7081) );
  OAI21_X1 U8945 ( .B1(n8050), .B2(n4773), .A(n7081), .ZN(n7082) );
  AOI21_X1 U8946 ( .B1(n7083), .B2(n9720), .A(n7082), .ZN(n7084) );
  OAI211_X1 U8947 ( .C1(n7086), .C2(n8086), .A(n7085), .B(n7084), .ZN(P2_U3193) );
  XNOR2_X1 U8948 ( .A(n7087), .B(n4694), .ZN(n9770) );
  XNOR2_X1 U8949 ( .A(n7089), .B(n7088), .ZN(n7090) );
  AOI222_X1 U8950 ( .A1(n9748), .A2(n7090), .B1(n7955), .B2(n9745), .C1(n9746), 
        .C2(n9743), .ZN(n9771) );
  MUX2_X1 U8951 ( .A(n7091), .B(n9771), .S(n8268), .Z(n7096) );
  INV_X1 U8952 ( .A(n7092), .ZN(n7093) );
  AOI22_X1 U8953 ( .A1(n9750), .A2(n7094), .B1(n9752), .B2(n7093), .ZN(n7095)
         );
  OAI211_X1 U8954 ( .C1(n8272), .C2(n9770), .A(n7096), .B(n7095), .ZN(P2_U3228) );
  NAND2_X1 U8955 ( .A1(n7110), .A2(n7358), .ZN(n7098) );
  OAI211_X1 U8956 ( .C1(n10004), .C2(n9522), .A(n7098), .B(n7097), .ZN(
        P1_U3335) );
  AOI21_X1 U8957 ( .B1(n7573), .B2(n7100), .A(n7099), .ZN(n7101) );
  OAI222_X1 U8958 ( .A1(n9548), .A2(n7103), .B1(n9550), .B2(n7102), .C1(n9546), 
        .C2(n7101), .ZN(n9767) );
  INV_X1 U8959 ( .A(n9767), .ZN(n7109) );
  OAI21_X1 U8960 ( .B1(n7105), .B2(n7573), .A(n7104), .ZN(n9769) );
  NOR2_X1 U8961 ( .A1(n8268), .A2(n5851), .ZN(n7107) );
  OAI22_X1 U8962 ( .A1(n8095), .A2(n9766), .B1(n7862), .B2(n9540), .ZN(n7106)
         );
  AOI211_X1 U8963 ( .C1(n9769), .C2(n9754), .A(n7107), .B(n7106), .ZN(n7108)
         );
  OAI21_X1 U8964 ( .B1(n7109), .B2(n9757), .A(n7108), .ZN(P2_U3229) );
  INV_X1 U8965 ( .A(n7110), .ZN(n7112) );
  INV_X1 U8966 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7111) );
  OAI222_X1 U8967 ( .A1(n5782), .A2(P2_U3151), .B1(n8451), .B2(n7112), .C1(
        n7111), .C2(n8449), .ZN(P2_U3275) );
  INV_X1 U8968 ( .A(n7113), .ZN(n7122) );
  INV_X1 U8969 ( .A(n7418), .ZN(n9339) );
  NAND2_X1 U8970 ( .A1(n7114), .A2(n9350), .ZN(n7117) );
  AOI22_X1 U8971 ( .A1(n9304), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7115), .B2(
        n9302), .ZN(n7116) );
  OAI211_X1 U8972 ( .C1(n7118), .C2(n9345), .A(n7117), .B(n7116), .ZN(n7119)
         );
  AOI21_X1 U8973 ( .B1(n9339), .B2(n7120), .A(n7119), .ZN(n7121) );
  OAI21_X1 U8974 ( .B1(n9304), .B2(n7122), .A(n7121), .ZN(P1_U3289) );
  INV_X1 U8975 ( .A(n7123), .ZN(n7130) );
  NAND2_X1 U8976 ( .A1(n7124), .A2(n9350), .ZN(n7126) );
  AOI22_X1 U8977 ( .A1(n9304), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9302), .B2(
        n5071), .ZN(n7125) );
  OAI211_X1 U8978 ( .C1(n8819), .C2(n9345), .A(n7126), .B(n7125), .ZN(n7127)
         );
  AOI21_X1 U8979 ( .B1(n9339), .B2(n7128), .A(n7127), .ZN(n7129) );
  OAI21_X1 U8980 ( .B1(n7130), .B2(n9304), .A(n7129), .ZN(P1_U3290) );
  NAND3_X1 U8981 ( .A1(n8654), .A2(n8638), .A3(n8645), .ZN(n7131) );
  NAND2_X1 U8982 ( .A1(n9690), .A2(n7142), .ZN(n8655) );
  OR2_X1 U8983 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  INV_X1 U8984 ( .A(n8634), .ZN(n8631) );
  OR2_X1 U8985 ( .A1(n7255), .A2(n7251), .ZN(n8826) );
  NAND2_X1 U8986 ( .A1(n7255), .A2(n7251), .ZN(n8658) );
  NAND2_X1 U8987 ( .A1(n8826), .A2(n8658), .ZN(n8768) );
  XNOR2_X1 U8988 ( .A(n7248), .B(n8768), .ZN(n7138) );
  OR2_X1 U8989 ( .A1(n7142), .A2(n8508), .ZN(n7137) );
  OAI21_X1 U8990 ( .B1(n7301), .B2(n9051), .A(n7137), .ZN(n9565) );
  AOI21_X1 U8991 ( .B1(n7138), .B2(n9333), .A(n9565), .ZN(n7200) );
  NAND2_X1 U8992 ( .A1(n7141), .A2(n7140), .ZN(n7163) );
  NAND2_X1 U8993 ( .A1(n8654), .A2(n8655), .ZN(n7162) );
  OAI21_X1 U8994 ( .B1(n7144), .B2(n8768), .A(n7257), .ZN(n7198) );
  NAND2_X1 U8995 ( .A1(n7198), .A2(n9339), .ZN(n7150) );
  OAI22_X1 U8996 ( .A1(n9678), .A2(n7145), .B1(n9574), .B2(n9673), .ZN(n7148)
         );
  INV_X1 U8997 ( .A(n7255), .ZN(n9569) );
  INV_X1 U8998 ( .A(n7260), .ZN(n7146) );
  OAI211_X1 U8999 ( .C1(n9569), .C2(n7156), .A(n7146), .B(n9216), .ZN(n7199)
         );
  NOR2_X1 U9000 ( .A1(n7199), .A2(n9660), .ZN(n7147) );
  AOI211_X1 U9001 ( .C1(n9657), .C2(n7255), .A(n7148), .B(n7147), .ZN(n7149)
         );
  OAI211_X1 U9002 ( .C1(n9304), .C2(n7200), .A(n7150), .B(n7149), .ZN(P1_U3283) );
  OAI21_X1 U9003 ( .B1(n7151), .B2(n8638), .A(n8645), .ZN(n7152) );
  XNOR2_X1 U9004 ( .A(n7152), .B(n7162), .ZN(n7154) );
  NOR2_X1 U9005 ( .A1(n7153), .A2(n8508), .ZN(n7268) );
  AOI21_X1 U9006 ( .B1(n7154), .B2(n9333), .A(n7268), .ZN(n9692) );
  OAI22_X1 U9007 ( .A1(n9678), .A2(n7155), .B1(n7273), .B2(n9673), .ZN(n7160)
         );
  AOI211_X1 U9008 ( .C1(n9690), .C2(n7157), .A(n9342), .B(n7156), .ZN(n7158)
         );
  NOR2_X1 U9009 ( .A1(n7251), .A2(n9051), .ZN(n7269) );
  NOR2_X1 U9010 ( .A1(n7158), .A2(n7269), .ZN(n9691) );
  NOR2_X1 U9011 ( .A1(n9691), .A2(n9660), .ZN(n7159) );
  AOI211_X1 U9012 ( .C1(n9657), .C2(n9690), .A(n7160), .B(n7159), .ZN(n7165)
         );
  OAI21_X1 U9013 ( .B1(n7163), .B2(n7162), .A(n7161), .ZN(n9694) );
  NAND2_X1 U9014 ( .A1(n9694), .A2(n9339), .ZN(n7164) );
  OAI211_X1 U9015 ( .C1(n9304), .C2(n9692), .A(n7165), .B(n7164), .ZN(P1_U3284) );
  INV_X1 U9016 ( .A(n7166), .ZN(n7175) );
  NOR2_X1 U9017 ( .A1(n9345), .A2(n7167), .ZN(n7170) );
  OAI22_X1 U9018 ( .A1(n9678), .A2(n6909), .B1(n7168), .B2(n9673), .ZN(n7169)
         );
  AOI211_X1 U9019 ( .C1(n7171), .C2(n9350), .A(n7170), .B(n7169), .ZN(n7174)
         );
  NAND2_X1 U9020 ( .A1(n7172), .A2(n9339), .ZN(n7173) );
  OAI211_X1 U9021 ( .C1(n7175), .C2(n9304), .A(n7174), .B(n7173), .ZN(P1_U3287) );
  INV_X1 U9022 ( .A(n7176), .ZN(n7186) );
  INV_X1 U9023 ( .A(n9339), .ZN(n9309) );
  INV_X1 U9024 ( .A(n7177), .ZN(n7178) );
  MUX2_X1 U9025 ( .A(n7179), .B(n7178), .S(n9678), .Z(n7185) );
  OAI22_X1 U9026 ( .A1(n9345), .A2(n7181), .B1(n7180), .B2(n9673), .ZN(n7182)
         );
  AOI21_X1 U9027 ( .B1(n7183), .B2(n9350), .A(n7182), .ZN(n7184) );
  OAI211_X1 U9028 ( .C1(n7186), .C2(n9309), .A(n7185), .B(n7184), .ZN(P1_U3288) );
  OAI21_X1 U9029 ( .B1(n7189), .B2(n7188), .A(n7187), .ZN(n7190) );
  NAND2_X1 U9030 ( .A1(n7190), .A2(n7934), .ZN(n7197) );
  NOR2_X1 U9031 ( .A1(n7928), .A2(n7293), .ZN(n7194) );
  NAND2_X1 U9032 ( .A1(n7940), .A2(n7955), .ZN(n7192) );
  OAI211_X1 U9033 ( .C1(n7371), .C2(n7942), .A(n7192), .B(n7191), .ZN(n7193)
         );
  AOI211_X1 U9034 ( .C1(n7195), .C2(n7930), .A(n7194), .B(n7193), .ZN(n7196)
         );
  NAND2_X1 U9035 ( .A1(n7197), .A2(n7196), .ZN(P2_U3153) );
  INV_X1 U9036 ( .A(n7198), .ZN(n7201) );
  OAI211_X1 U9037 ( .C1(n7201), .C2(n9446), .A(n7200), .B(n7199), .ZN(n7206)
         );
  INV_X1 U9038 ( .A(n7206), .ZN(n7203) );
  AOI22_X1 U9039 ( .A1(n7255), .A2(n9456), .B1(n9706), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7202) );
  OAI21_X1 U9040 ( .B1(n7203), .B2(n9706), .A(n7202), .ZN(P1_U3483) );
  INV_X1 U9041 ( .A(n6038), .ZN(n7237) );
  OAI222_X1 U9042 ( .A1(n9514), .A2(n7237), .B1(n8771), .B2(P1_U3086), .C1(
        n7204), .C2(n9522), .ZN(P1_U3334) );
  OAI22_X1 U9043 ( .A1(n9569), .A2(n9440), .B1(n9712), .B2(n5237), .ZN(n7205)
         );
  AOI21_X1 U9044 ( .B1(n7206), .B2(n9712), .A(n7205), .ZN(n7207) );
  INV_X1 U9045 ( .A(n7207), .ZN(P1_U3532) );
  NOR2_X1 U9046 ( .A1(n7208), .A2(n4359), .ZN(n7210) );
  NAND2_X1 U9047 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7383), .ZN(n7211) );
  OAI21_X1 U9048 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7383), .A(n7211), .ZN(
        n7212) );
  AOI21_X1 U9049 ( .B1(n7213), .B2(n7212), .A(n7381), .ZN(n7235) );
  INV_X1 U9050 ( .A(n7214), .ZN(n7220) );
  MUX2_X1 U9051 ( .A(n8290), .B(n7227), .S(n4398), .Z(n7216) );
  NAND2_X1 U9052 ( .A1(n7216), .A2(n7215), .ZN(n7393) );
  INV_X1 U9053 ( .A(n7216), .ZN(n7217) );
  NAND2_X1 U9054 ( .A1(n7217), .A2(n7383), .ZN(n7218) );
  AND2_X1 U9055 ( .A1(n7393), .A2(n7218), .ZN(n7219) );
  OAI21_X1 U9056 ( .B1(n7221), .B2(n7220), .A(n7219), .ZN(n7394) );
  INV_X1 U9057 ( .A(n7394), .ZN(n7223) );
  NOR3_X1 U9058 ( .A1(n7221), .A2(n7220), .A3(n7219), .ZN(n7222) );
  OAI21_X1 U9059 ( .B1(n7223), .B2(n7222), .A(n9887), .ZN(n7234) );
  NAND2_X1 U9060 ( .A1(n4773), .A2(n7224), .ZN(n7226) );
  NAND2_X1 U9061 ( .A1(n7226), .A2(n7225), .ZN(n7229) );
  MUX2_X1 U9062 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7227), .S(n7383), .Z(n7228)
         );
  NAND2_X1 U9063 ( .A1(n7228), .A2(n7229), .ZN(n7384) );
  OAI21_X1 U9064 ( .B1(n7229), .B2(n7228), .A(n7384), .ZN(n7232) );
  NAND2_X1 U9065 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n7814) );
  NAND2_X1 U9066 ( .A1(n9713), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7230) );
  OAI211_X1 U9067 ( .C1(n8050), .C2(n7383), .A(n7814), .B(n7230), .ZN(n7231)
         );
  AOI21_X1 U9068 ( .B1(n7232), .B2(n9720), .A(n7231), .ZN(n7233) );
  OAI211_X1 U9069 ( .C1(n7235), .C2(n8086), .A(n7234), .B(n7233), .ZN(P2_U3194) );
  INV_X1 U9070 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7236) );
  OAI222_X1 U9071 ( .A1(n7559), .A2(P2_U3151), .B1(n8451), .B2(n7237), .C1(
        n7236), .C2(n8449), .ZN(P2_U3274) );
  XNOR2_X1 U9072 ( .A(n7238), .B(n7504), .ZN(n9777) );
  XNOR2_X1 U9073 ( .A(n7240), .B(n7239), .ZN(n7241) );
  AOI222_X1 U9074 ( .A1(n9748), .A2(n7241), .B1(n9729), .B2(n9745), .C1(n7956), 
        .C2(n9743), .ZN(n9775) );
  MUX2_X1 U9075 ( .A(n7242), .B(n9775), .S(n8268), .Z(n7247) );
  INV_X1 U9076 ( .A(n7243), .ZN(n7244) );
  AOI22_X1 U9077 ( .A1(n9750), .A2(n7245), .B1(n9752), .B2(n7244), .ZN(n7246)
         );
  OAI211_X1 U9078 ( .C1(n8272), .C2(n9777), .A(n7247), .B(n7246), .ZN(P2_U3227) );
  NAND2_X1 U9079 ( .A1(n8581), .A2(n7301), .ZN(n8659) );
  NAND2_X1 U9080 ( .A1(n7334), .A2(n8659), .ZN(n8784) );
  NAND2_X1 U9081 ( .A1(n7249), .A2(n8784), .ZN(n7250) );
  NAND3_X1 U9082 ( .A1(n7335), .A2(n9333), .A3(n7250), .ZN(n7254) );
  OR2_X1 U9083 ( .A1(n7251), .A2(n8508), .ZN(n7252) );
  OAI21_X1 U9084 ( .B1(n7337), .B2(n9051), .A(n7252), .ZN(n8577) );
  INV_X1 U9085 ( .A(n8577), .ZN(n7253) );
  AND2_X1 U9086 ( .A1(n7254), .A2(n7253), .ZN(n9697) );
  OAI21_X1 U9087 ( .B1(n7258), .B2(n8784), .A(n7302), .ZN(n9704) );
  NAND2_X1 U9088 ( .A1(n9704), .A2(n9339), .ZN(n7264) );
  OAI22_X1 U9089 ( .A1(n9678), .A2(n7259), .B1(n8579), .B2(n9673), .ZN(n7262)
         );
  INV_X1 U9090 ( .A(n8581), .ZN(n9699) );
  OAI211_X1 U9091 ( .C1(n7260), .C2(n9699), .A(n9216), .B(n7304), .ZN(n9696)
         );
  NOR2_X1 U9092 ( .A1(n9696), .A2(n9660), .ZN(n7261) );
  AOI211_X1 U9093 ( .C1(n9657), .C2(n8581), .A(n7262), .B(n7261), .ZN(n7263)
         );
  OAI211_X1 U9094 ( .C1(n9304), .C2(n9697), .A(n7264), .B(n7263), .ZN(P1_U3282) );
  NAND2_X1 U9095 ( .A1(n7265), .A2(n9571), .ZN(n7277) );
  AOI21_X1 U9096 ( .B1(n7278), .B2(n7267), .A(n7266), .ZN(n7276) );
  OAI21_X1 U9097 ( .B1(n7269), .B2(n7268), .A(n9566), .ZN(n7272) );
  NOR2_X1 U9098 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7270), .ZN(n8979) );
  INV_X1 U9099 ( .A(n8979), .ZN(n7271) );
  OAI211_X1 U9100 ( .C1(n9575), .C2(n7273), .A(n7272), .B(n7271), .ZN(n7274)
         );
  AOI21_X1 U9101 ( .B1(n9690), .B2(n8613), .A(n7274), .ZN(n7275) );
  OAI21_X1 U9102 ( .B1(n7277), .B2(n7276), .A(n7275), .ZN(P1_U3231) );
  OAI21_X1 U9103 ( .B1(n7280), .B2(n7279), .A(n7278), .ZN(n7281) );
  NAND2_X1 U9104 ( .A1(n7281), .A2(n9571), .ZN(n7287) );
  NAND2_X1 U9105 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8965) );
  INV_X1 U9106 ( .A(n8965), .ZN(n7284) );
  NOR2_X1 U9107 ( .A1(n9575), .A2(n7282), .ZN(n7283) );
  AOI211_X1 U9108 ( .C1(n9566), .C2(n7285), .A(n7284), .B(n7283), .ZN(n7286)
         );
  OAI211_X1 U9109 ( .C1(n4650), .C2(n9568), .A(n7287), .B(n7286), .ZN(P1_U3221) );
  OAI21_X1 U9110 ( .B1(n7289), .B2(n7581), .A(n7288), .ZN(n7290) );
  AOI222_X1 U9111 ( .A1(n9748), .A2(n7290), .B1(n7954), .B2(n9745), .C1(n7955), 
        .C2(n9743), .ZN(n9782) );
  INV_X1 U9112 ( .A(n9735), .ZN(n7291) );
  AOI21_X1 U9113 ( .B1(n7581), .B2(n7292), .A(n7291), .ZN(n9785) );
  NOR2_X1 U9114 ( .A1(n8095), .A2(n9780), .ZN(n7295) );
  OAI22_X1 U9115 ( .A1(n8291), .A2(n6704), .B1(n7293), .B2(n9540), .ZN(n7294)
         );
  AOI211_X1 U9116 ( .C1(n9785), .C2(n9754), .A(n7295), .B(n7294), .ZN(n7296)
         );
  OAI21_X1 U9117 ( .B1(n9782), .B2(n9757), .A(n7296), .ZN(P2_U3226) );
  OR2_X1 U9118 ( .A1(n8502), .A2(n7337), .ZN(n8652) );
  NAND2_X1 U9119 ( .A1(n8502), .A2(n7337), .ZN(n8833) );
  NAND2_X1 U9120 ( .A1(n8652), .A2(n8833), .ZN(n8786) );
  NAND2_X1 U9121 ( .A1(n7335), .A2(n7334), .ZN(n7297) );
  XOR2_X1 U9122 ( .A(n8786), .B(n7297), .Z(n7300) );
  OR2_X1 U9123 ( .A1(n7301), .A2(n8508), .ZN(n7298) );
  OAI21_X1 U9124 ( .B1(n7411), .B2(n9051), .A(n7298), .ZN(n8498) );
  INV_X1 U9125 ( .A(n8498), .ZN(n7299) );
  OAI21_X1 U9126 ( .B1(n7300), .B2(n9240), .A(n7299), .ZN(n7323) );
  INV_X1 U9127 ( .A(n7323), .ZN(n7310) );
  INV_X1 U9128 ( .A(n7301), .ZN(n8873) );
  OAI21_X1 U9129 ( .B1(n7303), .B2(n8786), .A(n7342), .ZN(n7325) );
  NAND2_X1 U9130 ( .A1(n7325), .A2(n9339), .ZN(n7309) );
  AOI211_X1 U9131 ( .C1(n8502), .C2(n7304), .A(n9342), .B(n7345), .ZN(n7324)
         );
  NOR2_X1 U9132 ( .A1(n4424), .A2(n9345), .ZN(n7307) );
  OAI22_X1 U9133 ( .A1(n9678), .A2(n7305), .B1(n8500), .B2(n9673), .ZN(n7306)
         );
  AOI211_X1 U9134 ( .C1(n7324), .C2(n9350), .A(n7307), .B(n7306), .ZN(n7308)
         );
  OAI211_X1 U9135 ( .C1(n9304), .C2(n7310), .A(n7309), .B(n7308), .ZN(P1_U3281) );
  INV_X1 U9136 ( .A(n7187), .ZN(n7314) );
  INV_X1 U9137 ( .A(n7311), .ZN(n7313) );
  NOR3_X1 U9138 ( .A1(n7314), .A2(n7313), .A3(n7312), .ZN(n7317) );
  INV_X1 U9139 ( .A(n7315), .ZN(n7316) );
  OAI21_X1 U9140 ( .B1(n7317), .B2(n7316), .A(n7934), .ZN(n7322) );
  AOI21_X1 U9141 ( .B1(n7940), .B2(n9729), .A(n7318), .ZN(n7319) );
  OAI21_X1 U9142 ( .B1(n7424), .B2(n7942), .A(n7319), .ZN(n7320) );
  AOI21_X1 U9143 ( .B1(n9740), .B2(n7944), .A(n7320), .ZN(n7321) );
  OAI211_X1 U9144 ( .C1(n9789), .C2(n7947), .A(n7322), .B(n7321), .ZN(P2_U3161) );
  AOI211_X1 U9145 ( .C1(n7325), .C2(n9695), .A(n7324), .B(n7323), .ZN(n7329)
         );
  AOI22_X1 U9146 ( .A1(n8502), .A2(n9367), .B1(n9710), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7326) );
  OAI21_X1 U9147 ( .B1(n7329), .B2(n9710), .A(n7326), .ZN(P1_U3534) );
  NOR2_X1 U9148 ( .A1(n9707), .A2(n5293), .ZN(n7327) );
  AOI21_X1 U9149 ( .B1(n8502), .B2(n9456), .A(n7327), .ZN(n7328) );
  OAI21_X1 U9150 ( .B1(n7329), .B2(n9706), .A(n7328), .ZN(P1_U3489) );
  INV_X1 U9151 ( .A(n7330), .ZN(n7332) );
  OAI222_X1 U9152 ( .A1(n9522), .A2(n9936), .B1(n9514), .B2(n7332), .C1(
        P1_U3086), .C2(n8803), .ZN(P1_U3333) );
  OAI222_X1 U9153 ( .A1(P2_U3151), .A2(n7333), .B1(n8451), .B2(n7332), .C1(
        n7331), .C2(n8449), .ZN(P2_U3273) );
  AND2_X1 U9154 ( .A1(n8652), .A2(n7334), .ZN(n8830) );
  OR2_X1 U9155 ( .A1(n8558), .A2(n7411), .ZN(n8668) );
  NAND2_X1 U9156 ( .A1(n8558), .A2(n7411), .ZN(n8832) );
  NAND2_X1 U9157 ( .A1(n8668), .A2(n8832), .ZN(n7407) );
  XNOR2_X1 U9158 ( .A(n7408), .B(n7407), .ZN(n7341) );
  OR2_X1 U9159 ( .A1(n7337), .A2(n8508), .ZN(n7339) );
  NAND2_X1 U9160 ( .A1(n8870), .A2(n8588), .ZN(n7338) );
  NAND2_X1 U9161 ( .A1(n7339), .A2(n7338), .ZN(n8554) );
  INV_X1 U9162 ( .A(n8554), .ZN(n7340) );
  OAI21_X1 U9163 ( .B1(n7341), .B2(n9240), .A(n7340), .ZN(n7352) );
  INV_X1 U9164 ( .A(n7352), .ZN(n7351) );
  OAI21_X1 U9165 ( .B1(n7343), .B2(n7407), .A(n7403), .ZN(n7354) );
  NAND2_X1 U9166 ( .A1(n7354), .A2(n9339), .ZN(n7350) );
  INV_X1 U9167 ( .A(n7404), .ZN(n7346) );
  AOI211_X1 U9168 ( .C1(n8558), .C2(n4629), .A(n9342), .B(n7346), .ZN(n7353)
         );
  NOR2_X1 U9169 ( .A1(n7344), .A2(n9345), .ZN(n7348) );
  OAI22_X1 U9170 ( .A1(n9678), .A2(n5317), .B1(n8556), .B2(n9673), .ZN(n7347)
         );
  AOI211_X1 U9171 ( .C1(n7353), .C2(n9350), .A(n7348), .B(n7347), .ZN(n7349)
         );
  OAI211_X1 U9172 ( .C1(n9304), .C2(n7351), .A(n7350), .B(n7349), .ZN(P1_U3280) );
  AOI211_X1 U9173 ( .C1(n7354), .C2(n9695), .A(n7353), .B(n7352), .ZN(n7357)
         );
  AOI22_X1 U9174 ( .A1(n8558), .A2(n9456), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9706), .ZN(n7355) );
  OAI21_X1 U9175 ( .B1(n7357), .B2(n9706), .A(n7355), .ZN(P1_U3492) );
  AOI22_X1 U9176 ( .A1(n8558), .A2(n9367), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9710), .ZN(n7356) );
  OAI21_X1 U9177 ( .B1(n7357), .B2(n9710), .A(n7356), .ZN(P1_U3535) );
  NAND2_X1 U9178 ( .A1(n7361), .A2(n7358), .ZN(n7359) );
  OAI211_X1 U9179 ( .C1(n10025), .C2(n9522), .A(n7359), .B(n8866), .ZN(
        P1_U3332) );
  NAND2_X1 U9180 ( .A1(n7361), .A2(n7360), .ZN(n7363) );
  OR2_X1 U9181 ( .A1(n7362), .A2(P2_U3151), .ZN(n7706) );
  OAI211_X1 U9182 ( .C1(n10005), .C2(n8449), .A(n7363), .B(n7706), .ZN(
        P2_U3272) );
  OR2_X1 U9183 ( .A1(n7364), .A2(n7506), .ZN(n7365) );
  INV_X1 U9184 ( .A(n7373), .ZN(n9795) );
  NAND2_X1 U9185 ( .A1(n8291), .A2(n7366), .ZN(n8104) );
  INV_X1 U9186 ( .A(n7369), .ZN(n7370) );
  AOI21_X1 U9187 ( .B1(n7506), .B2(n7367), .A(n7370), .ZN(n7375) );
  OAI22_X1 U9188 ( .A1(n7371), .A2(n9548), .B1(n7473), .B2(n9550), .ZN(n7372)
         );
  AOI21_X1 U9189 ( .B1(n7373), .B2(n9786), .A(n7372), .ZN(n7374) );
  OAI21_X1 U9190 ( .B1(n7375), .B2(n9546), .A(n7374), .ZN(n9797) );
  NAND2_X1 U9191 ( .A1(n9797), .A2(n8268), .ZN(n7380) );
  OAI22_X1 U9192 ( .A1(n8291), .A2(n6835), .B1(n7376), .B2(n9540), .ZN(n7377)
         );
  AOI21_X1 U9193 ( .B1(n9750), .B2(n7378), .A(n7377), .ZN(n7379) );
  OAI211_X1 U9194 ( .C1(n9795), .C2(n8104), .A(n7380), .B(n7379), .ZN(P2_U3224) );
  INV_X1 U9195 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9554) );
  AOI21_X1 U9196 ( .B1(n9554), .B2(n7382), .A(n7961), .ZN(n7401) );
  NAND2_X1 U9197 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7383), .ZN(n7385) );
  NAND2_X1 U9198 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7386), .ZN(n7967) );
  OAI21_X1 U9199 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7386), .A(n7967), .ZN(
        n7399) );
  AND2_X1 U9200 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7882) );
  AOI21_X1 U9201 ( .B1(n9713), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7882), .ZN(
        n7387) );
  OAI21_X1 U9202 ( .B1(n8050), .B2(n7966), .A(n7387), .ZN(n7398) );
  MUX2_X1 U9203 ( .A(n9554), .B(n7388), .S(n4398), .Z(n7389) );
  NAND2_X1 U9204 ( .A1(n7389), .A2(n7960), .ZN(n7973) );
  INV_X1 U9205 ( .A(n7389), .ZN(n7390) );
  NAND2_X1 U9206 ( .A1(n7390), .A2(n7966), .ZN(n7391) );
  NAND2_X1 U9207 ( .A1(n7973), .A2(n7391), .ZN(n7392) );
  AOI21_X1 U9208 ( .B1(n7394), .B2(n7393), .A(n7392), .ZN(n7981) );
  INV_X1 U9209 ( .A(n7981), .ZN(n7396) );
  NAND3_X1 U9210 ( .A1(n7394), .A2(n7393), .A3(n7392), .ZN(n7395) );
  AOI21_X1 U9211 ( .B1(n7396), .B2(n7395), .A(n8082), .ZN(n7397) );
  AOI211_X1 U9212 ( .C1(n9720), .C2(n7399), .A(n7398), .B(n7397), .ZN(n7400)
         );
  OAI21_X1 U9213 ( .B1(n7401), .B2(n8086), .A(n7400), .ZN(P2_U3195) );
  INV_X1 U9214 ( .A(n8870), .ZN(n7434) );
  NAND2_X1 U9215 ( .A1(n9442), .A2(n7434), .ZN(n8835) );
  NAND2_X1 U9216 ( .A1(n8670), .A2(n8835), .ZN(n7409) );
  XNOR2_X1 U9217 ( .A(n7436), .B(n4644), .ZN(n9447) );
  AOI211_X1 U9218 ( .C1(n9442), .C2(n7404), .A(n9342), .B(n7443), .ZN(n9441)
         );
  INV_X1 U9219 ( .A(n7405), .ZN(n8461) );
  AOI22_X1 U9220 ( .A1(n9304), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8461), .B2(
        n9302), .ZN(n7406) );
  OAI21_X1 U9221 ( .B1(n4627), .B2(n9345), .A(n7406), .ZN(n7416) );
  INV_X1 U9222 ( .A(n7407), .ZN(n8788) );
  AOI21_X1 U9223 ( .B1(n7410), .B2(n7409), .A(n9240), .ZN(n7414) );
  OR2_X1 U9224 ( .A1(n7411), .A2(n8508), .ZN(n7413) );
  NAND2_X1 U9225 ( .A1(n9077), .A2(n8588), .ZN(n7412) );
  NAND2_X1 U9226 ( .A1(n7413), .A2(n7412), .ZN(n8457) );
  AOI21_X1 U9227 ( .B1(n7414), .B2(n7437), .A(n8457), .ZN(n9445) );
  NOR2_X1 U9228 ( .A1(n9445), .A2(n9304), .ZN(n7415) );
  AOI211_X1 U9229 ( .C1(n9441), .C2(n9350), .A(n7416), .B(n7415), .ZN(n7417)
         );
  OAI21_X1 U9230 ( .B1(n9447), .B2(n7418), .A(n7417), .ZN(P1_U3279) );
  NAND2_X1 U9231 ( .A1(n7419), .A2(n7579), .ZN(n7420) );
  XNOR2_X1 U9232 ( .A(n7420), .B(n7507), .ZN(n9799) );
  INV_X1 U9233 ( .A(n9786), .ZN(n7427) );
  AND3_X1 U9234 ( .A1(n7369), .A2(n7507), .A3(n7421), .ZN(n7422) );
  OAI21_X1 U9235 ( .B1(n7423), .B2(n7422), .A(n9748), .ZN(n7426) );
  AOI22_X1 U9236 ( .A1(n9743), .A2(n9730), .B1(n7952), .B2(n9745), .ZN(n7425)
         );
  OAI211_X1 U9237 ( .C1(n9799), .C2(n7427), .A(n7426), .B(n7425), .ZN(n9800)
         );
  NAND2_X1 U9238 ( .A1(n9800), .A2(n8268), .ZN(n7430) );
  OAI22_X1 U9239 ( .A1(n8268), .A2(n7041), .B1(n7460), .B2(n9540), .ZN(n7428)
         );
  AOI21_X1 U9240 ( .B1(n9750), .B2(n9802), .A(n7428), .ZN(n7429) );
  OAI211_X1 U9241 ( .C1(n9799), .C2(n8104), .A(n7430), .B(n7429), .ZN(P2_U3223) );
  INV_X1 U9242 ( .A(n7431), .ZN(n7451) );
  OAI222_X1 U9243 ( .A1(n9514), .A2(n7451), .B1(P1_U3086), .B2(n7433), .C1(
        n7432), .C2(n9522), .ZN(P1_U3331) );
  NAND2_X1 U9244 ( .A1(n9442), .A2(n8870), .ZN(n7435) );
  INV_X1 U9245 ( .A(n9077), .ZN(n9081) );
  OR2_X1 U9246 ( .A1(n9078), .A2(n9081), .ZN(n8671) );
  NAND2_X1 U9247 ( .A1(n9078), .A2(n9081), .ZN(n9329) );
  XNOR2_X1 U9248 ( .A(n9080), .B(n8789), .ZN(n9438) );
  INV_X1 U9249 ( .A(n9438), .ZN(n7450) );
  XNOR2_X1 U9250 ( .A(n8745), .B(n8789), .ZN(n7438) );
  NAND2_X1 U9251 ( .A1(n7438), .A2(n9333), .ZN(n7442) );
  NAND2_X1 U9252 ( .A1(n8870), .A2(n9074), .ZN(n7440) );
  NAND2_X1 U9253 ( .A1(n9082), .A2(n8588), .ZN(n7439) );
  NAND2_X1 U9254 ( .A1(n7440), .A2(n7439), .ZN(n8609) );
  INV_X1 U9255 ( .A(n8609), .ZN(n7441) );
  NAND2_X1 U9256 ( .A1(n7442), .A2(n7441), .ZN(n9436) );
  INV_X1 U9257 ( .A(n7443), .ZN(n7444) );
  AOI211_X1 U9258 ( .C1(n9078), .C2(n7444), .A(n9342), .B(n9340), .ZN(n9437)
         );
  NAND2_X1 U9259 ( .A1(n9437), .A2(n9350), .ZN(n7447) );
  INV_X1 U9260 ( .A(n8611), .ZN(n7445) );
  AOI22_X1 U9261 ( .A1(n9304), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7445), .B2(
        n9302), .ZN(n7446) );
  OAI211_X1 U9262 ( .C1(n9504), .C2(n9345), .A(n7447), .B(n7446), .ZN(n7448)
         );
  AOI21_X1 U9263 ( .B1(n9678), .B2(n9436), .A(n7448), .ZN(n7449) );
  OAI21_X1 U9264 ( .B1(n7450), .B2(n9309), .A(n7449), .ZN(P1_U3278) );
  OAI222_X1 U9265 ( .A1(n7452), .A2(P2_U3151), .B1(n8451), .B2(n7451), .C1(
        n10010), .C2(n8449), .ZN(P2_U3271) );
  INV_X1 U9266 ( .A(n7453), .ZN(n7454) );
  NAND2_X1 U9267 ( .A1(n7454), .A2(n9730), .ZN(n7455) );
  XNOR2_X1 U9268 ( .A(n9802), .B(n7796), .ZN(n7457) );
  OAI21_X1 U9269 ( .B1(n7458), .B2(n7457), .A(n7722), .ZN(n7459) );
  NAND2_X1 U9270 ( .A1(n7459), .A2(n7934), .ZN(n7466) );
  NOR2_X1 U9271 ( .A1(n7928), .A2(n7460), .ZN(n7464) );
  NAND2_X1 U9272 ( .A1(n7940), .A2(n9730), .ZN(n7462) );
  OAI211_X1 U9273 ( .C1(n8287), .C2(n7942), .A(n7462), .B(n7461), .ZN(n7463)
         );
  AOI211_X1 U9274 ( .C1(n9802), .C2(n7930), .A(n7464), .B(n7463), .ZN(n7465)
         );
  NAND2_X1 U9275 ( .A1(n7466), .A2(n7465), .ZN(P2_U3157) );
  INV_X1 U9276 ( .A(n7467), .ZN(n7478) );
  OAI222_X1 U9277 ( .A1(n9514), .A2(n7478), .B1(P1_U3086), .B2(n7469), .C1(
        n7468), .C2(n9522), .ZN(P1_U3330) );
  XNOR2_X1 U9278 ( .A(n7471), .B(n7501), .ZN(n9805) );
  XNOR2_X1 U9279 ( .A(n4363), .B(n7501), .ZN(n7472) );
  OAI222_X1 U9280 ( .A1(n9550), .A2(n9547), .B1(n9548), .B2(n7473), .C1(n7472), 
        .C2(n9546), .ZN(n9806) );
  NAND2_X1 U9281 ( .A1(n9806), .A2(n8268), .ZN(n7476) );
  OAI22_X1 U9282 ( .A1(n8291), .A2(n7070), .B1(n7902), .B2(n9540), .ZN(n7474)
         );
  AOI21_X1 U9283 ( .B1(n9808), .B2(n9750), .A(n7474), .ZN(n7475) );
  OAI211_X1 U9284 ( .C1(n9805), .C2(n8272), .A(n7476), .B(n7475), .ZN(P2_U3222) );
  OAI222_X1 U9285 ( .A1(n7479), .A2(P2_U3151), .B1(n8451), .B2(n7478), .C1(
        n7477), .C2(n8449), .ZN(P2_U3270) );
  INV_X1 U9286 ( .A(n7480), .ZN(n7482) );
  OAI222_X1 U9287 ( .A1(n9514), .A2(n7482), .B1(P1_U3086), .B2(n7481), .C1(
        n9998), .C2(n9522), .ZN(P1_U3329) );
  OAI222_X1 U9288 ( .A1(n7483), .A2(P2_U3151), .B1(n8451), .B2(n7482), .C1(
        n10024), .C2(n8449), .ZN(P2_U3269) );
  INV_X1 U9289 ( .A(SI_29_), .ZN(n7487) );
  OR2_X1 U9290 ( .A1(n7485), .A2(n7484), .ZN(n7486) );
  INV_X1 U9291 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7719) );
  INV_X1 U9292 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9515) );
  MUX2_X1 U9293 ( .A(n7719), .B(n9515), .S(n7521), .Z(n7490) );
  INV_X1 U9294 ( .A(SI_30_), .ZN(n7489) );
  NAND2_X1 U9295 ( .A1(n7490), .A2(n7489), .ZN(n7518) );
  INV_X1 U9296 ( .A(n7490), .ZN(n7491) );
  NAND2_X1 U9297 ( .A1(n7491), .A2(SI_30_), .ZN(n7492) );
  NAND2_X1 U9298 ( .A1(n7518), .A2(n7492), .ZN(n7519) );
  NAND2_X1 U9299 ( .A1(n7718), .A2(n7525), .ZN(n7494) );
  OR2_X1 U9300 ( .A1(n7526), .A2(n7719), .ZN(n7493) );
  NAND2_X1 U9301 ( .A1(n8363), .A2(n7495), .ZN(n7540) );
  INV_X1 U9302 ( .A(n7540), .ZN(n7685) );
  NOR2_X1 U9303 ( .A1(n7685), .A2(n7687), .ZN(n7538) );
  INV_X1 U9304 ( .A(n7795), .ZN(n7516) );
  INV_X1 U9305 ( .A(n7496), .ZN(n7548) );
  INV_X1 U9306 ( .A(n8155), .ZN(n7497) );
  INV_X1 U9307 ( .A(n7498), .ZN(n7622) );
  OR2_X1 U9308 ( .A1(n7621), .A2(n7622), .ZN(n8281) );
  NAND2_X1 U9309 ( .A1(n7500), .A2(n7499), .ZN(n7620) );
  NOR2_X1 U9310 ( .A1(n8293), .A2(n7501), .ZN(n7612) );
  INV_X1 U9311 ( .A(n7612), .ZN(n7510) );
  NOR2_X1 U9312 ( .A1(n5832), .A2(n6115), .ZN(n7503) );
  NAND4_X1 U9313 ( .A1(n7503), .A2(n7573), .A3(n7502), .A4(n9749), .ZN(n7505)
         );
  NOR4_X1 U9314 ( .A1(n7505), .A2(n4694), .A3(n7581), .A4(n7504), .ZN(n7508)
         );
  NAND4_X1 U9315 ( .A1(n7508), .A2(n7507), .A3(n7506), .A4(n9732), .ZN(n7509)
         );
  NOR4_X1 U9316 ( .A1(n8281), .A2(n4589), .A3(n7510), .A4(n7509), .ZN(n7511)
         );
  AND4_X1 U9317 ( .A1(n6008), .A2(n8264), .A3(n8251), .A4(n7511), .ZN(n7512)
         );
  NAND4_X1 U9318 ( .A1(n8201), .A2(n8218), .A3(n8225), .A4(n7512), .ZN(n7513)
         );
  NOR4_X1 U9319 ( .A1(n8162), .A2(n8171), .A3(n8187), .A4(n7513), .ZN(n7514)
         );
  NAND4_X1 U9320 ( .A1(n8125), .A2(n8138), .A3(n8157), .A4(n7514), .ZN(n7515)
         );
  NOR4_X1 U9321 ( .A1(n7517), .A2(n7516), .A3(n7551), .A4(n7515), .ZN(n7537)
         );
  OAI21_X1 U9322 ( .B1(n7520), .B2(n7519), .A(n7518), .ZN(n7524) );
  INV_X1 U9323 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8618) );
  MUX2_X1 U9324 ( .A(n6369), .B(n8618), .S(n7521), .Z(n7522) );
  XNOR2_X1 U9325 ( .A(n7522), .B(SI_31_), .ZN(n7523) );
  XNOR2_X1 U9326 ( .A(n7524), .B(n7523), .ZN(n8617) );
  NAND2_X1 U9327 ( .A1(n8617), .A2(n7525), .ZN(n7528) );
  OR2_X1 U9328 ( .A1(n7526), .A2(n6369), .ZN(n7527) );
  INV_X1 U9329 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7529) );
  OR2_X1 U9330 ( .A1(n7530), .A2(n7529), .ZN(n7535) );
  INV_X1 U9331 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7531) );
  OR2_X1 U9332 ( .A1(n5817), .A2(n7531), .ZN(n7534) );
  NAND2_X1 U9333 ( .A1(n7532), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7533) );
  NAND4_X1 U9334 ( .A1(n7536), .A2(n7535), .A3(n7534), .A4(n7533), .ZN(n8091)
         );
  INV_X1 U9335 ( .A(n8091), .ZN(n7542) );
  AND2_X1 U9336 ( .A1(n8298), .A2(n7542), .ZN(n7694) );
  NAND2_X1 U9337 ( .A1(n8362), .A2(n8091), .ZN(n7690) );
  NAND4_X1 U9338 ( .A1(n7538), .A2(n7537), .A3(n7695), .A4(n7690), .ZN(n7547)
         );
  INV_X1 U9339 ( .A(n7674), .ZN(n7680) );
  OAI21_X1 U9340 ( .B1(n7541), .B2(n7680), .A(n4289), .ZN(n7545) );
  INV_X1 U9341 ( .A(n8363), .ZN(n8303) );
  OAI21_X1 U9342 ( .B1(n8303), .B2(n8298), .A(n7690), .ZN(n7544) );
  OAI21_X1 U9343 ( .B1(n7687), .B2(n7542), .A(n8298), .ZN(n7543) );
  MUX2_X1 U9344 ( .A(n7549), .B(n7548), .S(n7675), .Z(n7550) );
  NOR2_X1 U9345 ( .A1(n7551), .A2(n7550), .ZN(n7673) );
  INV_X1 U9346 ( .A(n7552), .ZN(n7553) );
  NAND2_X1 U9347 ( .A1(n7554), .A2(n7553), .ZN(n7556) );
  AND2_X1 U9348 ( .A1(n7556), .A2(n7555), .ZN(n7614) );
  NAND2_X1 U9349 ( .A1(n7614), .A2(n7691), .ZN(n7613) );
  NAND2_X1 U9350 ( .A1(n7565), .A2(n7675), .ZN(n7557) );
  OAI21_X1 U9351 ( .B1(n6115), .B2(n7558), .A(n7557), .ZN(n7564) );
  NAND2_X1 U9352 ( .A1(n7560), .A2(n7559), .ZN(n7562) );
  NAND3_X1 U9353 ( .A1(n7562), .A2(n7675), .A3(n7561), .ZN(n7563) );
  NAND2_X1 U9354 ( .A1(n7564), .A2(n7563), .ZN(n7568) );
  MUX2_X1 U9355 ( .A(n7566), .B(n7565), .S(n7691), .Z(n7567) );
  NAND3_X1 U9356 ( .A1(n7568), .A2(n5833), .A3(n7567), .ZN(n7572) );
  NAND2_X1 U9357 ( .A1(n7584), .A2(n5834), .ZN(n7571) );
  NAND2_X1 U9358 ( .A1(n7957), .A2(n4522), .ZN(n7574) );
  NAND2_X1 U9359 ( .A1(n7574), .A2(n7569), .ZN(n7570) );
  INV_X1 U9360 ( .A(n7574), .ZN(n7576) );
  OAI211_X1 U9361 ( .C1(n7588), .C2(n7576), .A(n7589), .B(n7575), .ZN(n7577)
         );
  NAND3_X1 U9362 ( .A1(n7577), .A2(n7585), .A3(n7592), .ZN(n7583) );
  AND2_X1 U9363 ( .A1(n7600), .A2(n7691), .ZN(n7578) );
  NAND2_X1 U9364 ( .A1(n7579), .A2(n7578), .ZN(n7599) );
  NAND3_X1 U9365 ( .A1(n7597), .A2(n7675), .A3(n7596), .ZN(n7580) );
  NAND2_X1 U9366 ( .A1(n7599), .A2(n7580), .ZN(n7602) );
  INV_X1 U9367 ( .A(n7581), .ZN(n7582) );
  AND2_X1 U9368 ( .A1(n7602), .A2(n7582), .ZN(n7593) );
  INV_X1 U9369 ( .A(n7584), .ZN(n7587) );
  OAI211_X1 U9370 ( .C1(n7588), .C2(n7587), .A(n7586), .B(n7585), .ZN(n7591)
         );
  NAND3_X1 U9371 ( .A1(n7591), .A2(n7590), .A3(n7589), .ZN(n7594) );
  AND2_X1 U9372 ( .A1(n7596), .A2(n7595), .ZN(n7598) );
  OAI211_X1 U9373 ( .C1(n7599), .C2(n7598), .A(n7597), .B(n7609), .ZN(n7606)
         );
  NAND2_X1 U9374 ( .A1(n7600), .A2(n9734), .ZN(n7601) );
  NAND2_X1 U9375 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  NAND2_X1 U9376 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  MUX2_X1 U9377 ( .A(n7606), .B(n7605), .S(n7675), .Z(n7607) );
  INV_X1 U9378 ( .A(n7607), .ZN(n7611) );
  MUX2_X1 U9379 ( .A(n7609), .B(n7608), .S(n7691), .Z(n7610) );
  INV_X1 U9380 ( .A(n7614), .ZN(n7615) );
  NAND2_X1 U9381 ( .A1(n7615), .A2(n7675), .ZN(n7616) );
  MUX2_X1 U9382 ( .A(n7618), .B(n7617), .S(n7675), .Z(n7619) );
  MUX2_X1 U9383 ( .A(n7622), .B(n7621), .S(n7691), .Z(n7623) );
  INV_X1 U9384 ( .A(n7623), .ZN(n7624) );
  MUX2_X1 U9385 ( .A(n7626), .B(n7625), .S(n7675), .Z(n7627) );
  NAND3_X1 U9386 ( .A1(n7628), .A2(n8251), .A3(n7627), .ZN(n7634) );
  MUX2_X1 U9387 ( .A(n7630), .B(n7629), .S(n7691), .Z(n7631) );
  INV_X1 U9388 ( .A(n7631), .ZN(n7632) );
  NOR2_X1 U9389 ( .A1(n8239), .A2(n7632), .ZN(n7633) );
  NAND2_X1 U9390 ( .A1(n7634), .A2(n7633), .ZN(n7639) );
  INV_X1 U9391 ( .A(n7637), .ZN(n7635) );
  NAND3_X1 U9392 ( .A1(n7639), .A2(n7638), .A3(n7637), .ZN(n7641) );
  AOI21_X1 U9393 ( .B1(n7641), .B2(n7640), .A(n7691), .ZN(n7642) );
  INV_X1 U9394 ( .A(n7644), .ZN(n7646) );
  OAI21_X1 U9395 ( .B1(n7649), .B2(n7646), .A(n7645), .ZN(n7647) );
  NAND2_X1 U9396 ( .A1(n7649), .A2(n7648), .ZN(n7651) );
  NAND2_X1 U9397 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  INV_X1 U9398 ( .A(n7653), .ZN(n7656) );
  INV_X1 U9399 ( .A(n7654), .ZN(n7655) );
  MUX2_X1 U9400 ( .A(n7656), .B(n7655), .S(n7691), .Z(n7657) );
  NAND2_X1 U9401 ( .A1(n6064), .A2(n7664), .ZN(n7658) );
  AOI22_X1 U9402 ( .A1(n7660), .A2(n7661), .B1(n7659), .B2(n7658), .ZN(n7665)
         );
  MUX2_X1 U9403 ( .A(n7667), .B(n7666), .S(n7691), .Z(n7668) );
  MUX2_X1 U9404 ( .A(n7670), .B(n7669), .S(n7691), .Z(n7671) );
  AOI21_X1 U9405 ( .B1(n7673), .B2(n7672), .A(n7671), .ZN(n7682) );
  MUX2_X1 U9406 ( .A(n7950), .B(n8111), .S(n7675), .Z(n7681) );
  NOR2_X1 U9407 ( .A1(n7682), .A2(n7681), .ZN(n7679) );
  OAI21_X1 U9408 ( .B1(n7676), .B2(n7675), .A(n7674), .ZN(n7678) );
  NAND3_X1 U9409 ( .A1(n7683), .A2(n7682), .A3(n7681), .ZN(n7684) );
  NAND2_X1 U9410 ( .A1(n4344), .A2(n7691), .ZN(n7696) );
  INV_X1 U9411 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U9412 ( .A1(n7689), .A2(n7688), .ZN(n7692) );
  NAND3_X1 U9413 ( .A1(n7702), .A2(n7701), .A3(n4398), .ZN(n7703) );
  OAI211_X1 U9414 ( .C1(n7704), .C2(n7706), .A(n7703), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7705) );
  INV_X1 U9415 ( .A(n9379), .ZN(n9152) );
  AOI21_X1 U9416 ( .B1(n8598), .B2(n7708), .A(n7707), .ZN(n7710) );
  OAI21_X1 U9417 ( .B1(n7710), .B2(n7709), .A(n9571), .ZN(n7715) );
  INV_X1 U9418 ( .A(n7711), .ZN(n9149) );
  AOI22_X1 U9419 ( .A1(n9075), .A2(n8588), .B1(n9074), .B2(n9116), .ZN(n9146)
         );
  OAI22_X1 U9420 ( .A1(n8601), .A2(n9146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7712), .ZN(n7713) );
  AOI21_X1 U9421 ( .B1(n8568), .B2(n9149), .A(n7713), .ZN(n7714) );
  OAI211_X1 U9422 ( .C1(n9152), .C2(n9568), .A(n7715), .B(n7714), .ZN(P1_U3214) );
  OAI222_X1 U9423 ( .A1(n9522), .A2(n10019), .B1(n9514), .B2(n7716), .C1(
        P1_U3086), .C2(n8810), .ZN(P1_U3336) );
  INV_X1 U9424 ( .A(n7718), .ZN(n9513) );
  OAI222_X1 U9425 ( .A1(n7717), .A2(P2_U3151), .B1(n8451), .B2(n9513), .C1(
        n7719), .C2(n8449), .ZN(P2_U3265) );
  XNOR2_X1 U9426 ( .A(n8405), .B(n7796), .ZN(n7737) );
  INV_X1 U9427 ( .A(n7737), .ZN(n7738) );
  INV_X1 U9428 ( .A(n8211), .ZN(n8191) );
  XNOR2_X1 U9429 ( .A(n8330), .B(n7796), .ZN(n7735) );
  INV_X1 U9430 ( .A(n7735), .ZN(n7736) );
  XNOR2_X1 U9431 ( .A(n8422), .B(n7796), .ZN(n7730) );
  XNOR2_X1 U9432 ( .A(n9808), .B(n7796), .ZN(n7723) );
  INV_X1 U9433 ( .A(n7723), .ZN(n7724) );
  XNOR2_X1 U9434 ( .A(n7723), .B(n8287), .ZN(n7904) );
  XNOR2_X1 U9435 ( .A(n9815), .B(n7796), .ZN(n7725) );
  XNOR2_X1 U9436 ( .A(n7725), .B(n9547), .ZN(n7812) );
  XNOR2_X1 U9437 ( .A(n9538), .B(n7796), .ZN(n7726) );
  NAND2_X1 U9438 ( .A1(n7726), .A2(n8288), .ZN(n7876) );
  NOR2_X1 U9439 ( .A1(n7726), .A2(n8288), .ZN(n7878) );
  XNOR2_X1 U9440 ( .A(n8435), .B(n7796), .ZN(n7727) );
  XNOR2_X1 U9441 ( .A(n7727), .B(n8266), .ZN(n7759) );
  XNOR2_X1 U9442 ( .A(n7948), .B(n7796), .ZN(n7728) );
  XNOR2_X1 U9443 ( .A(n7728), .B(n8253), .ZN(n7936) );
  XNOR2_X1 U9444 ( .A(n7730), .B(n8265), .ZN(n7829) );
  XNOR2_X1 U9445 ( .A(n8339), .B(n7796), .ZN(n7731) );
  XNOR2_X1 U9446 ( .A(n7731), .B(n8254), .ZN(n7838) );
  INV_X1 U9447 ( .A(n7731), .ZN(n7732) );
  NOR2_X1 U9448 ( .A1(n7732), .A2(n8228), .ZN(n7910) );
  XNOR2_X1 U9449 ( .A(n8412), .B(n7750), .ZN(n7733) );
  XNOR2_X1 U9450 ( .A(n7733), .B(n8243), .ZN(n7909) );
  XNOR2_X1 U9451 ( .A(n7735), .B(n7915), .ZN(n7783) );
  XOR2_X1 U9452 ( .A(n8211), .B(n7737), .Z(n7868) );
  XNOR2_X1 U9453 ( .A(n8399), .B(n7796), .ZN(n7739) );
  XOR2_X1 U9454 ( .A(n7892), .B(n7739), .Z(n7806) );
  XNOR2_X1 U9455 ( .A(n7898), .B(n7796), .ZN(n7740) );
  XNOR2_X1 U9456 ( .A(n7740), .B(n7767), .ZN(n7888) );
  INV_X1 U9457 ( .A(n7767), .ZN(n7741) );
  NAND2_X1 U9458 ( .A1(n7740), .A2(n7741), .ZN(n7742) );
  XNOR2_X1 U9459 ( .A(n8382), .B(n7796), .ZN(n7848) );
  XNOR2_X1 U9460 ( .A(n8388), .B(n7750), .ZN(n7845) );
  INV_X1 U9461 ( .A(n7845), .ZN(n7743) );
  OAI22_X1 U9462 ( .A1(n7848), .A2(n7847), .B1(n7766), .B2(n7743), .ZN(n7747)
         );
  OAI21_X1 U9463 ( .B1(n7845), .B2(n8178), .A(n8164), .ZN(n7745) );
  NOR2_X1 U9464 ( .A1(n8178), .A2(n8164), .ZN(n7744) );
  AOI22_X1 U9465 ( .A1(n7745), .A2(n7848), .B1(n7744), .B2(n7743), .ZN(n7746)
         );
  XNOR2_X1 U9466 ( .A(n8379), .B(n7796), .ZN(n7748) );
  XNOR2_X1 U9467 ( .A(n7748), .B(n7851), .ZN(n7821) );
  INV_X1 U9468 ( .A(n7748), .ZN(n7749) );
  XNOR2_X1 U9469 ( .A(n8372), .B(n7750), .ZN(n7752) );
  NOR2_X1 U9470 ( .A1(n7752), .A2(n7751), .ZN(n7923) );
  NAND2_X1 U9471 ( .A1(n7752), .A2(n7751), .ZN(n7921) );
  INV_X1 U9472 ( .A(n7753), .ZN(n7794) );
  XNOR2_X1 U9473 ( .A(n8119), .B(n7796), .ZN(n7791) );
  XNOR2_X1 U9474 ( .A(n7791), .B(n8126), .ZN(n7793) );
  XNOR2_X1 U9475 ( .A(n7794), .B(n7793), .ZN(n7758) );
  AOI22_X1 U9476 ( .A1(n7925), .A2(n7950), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7755) );
  NAND2_X1 U9477 ( .A1(n7940), .A2(n8140), .ZN(n7754) );
  OAI211_X1 U9478 ( .C1(n8114), .C2(n7928), .A(n7755), .B(n7754), .ZN(n7756)
         );
  AOI21_X1 U9479 ( .B1(n8119), .B2(n7930), .A(n7756), .ZN(n7757) );
  OAI21_X1 U9480 ( .B1(n7758), .B2(n7932), .A(n7757), .ZN(P2_U3154) );
  XOR2_X1 U9481 ( .A(n7760), .B(n7759), .Z(n7765) );
  NAND2_X1 U9482 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7972) );
  OAI21_X1 U9483 ( .B1(n7893), .B2(n8288), .A(n7972), .ZN(n7761) );
  AOI21_X1 U9484 ( .B1(n7925), .B2(n7729), .A(n7761), .ZN(n7762) );
  OAI21_X1 U9485 ( .B1(n8277), .B2(n7928), .A(n7762), .ZN(n7763) );
  AOI21_X1 U9486 ( .B1(n8435), .B2(n7930), .A(n7763), .ZN(n7764) );
  OAI21_X1 U9487 ( .B1(n7765), .B2(n7932), .A(n7764), .ZN(P2_U3155) );
  XNOR2_X1 U9488 ( .A(n7846), .B(n7766), .ZN(n7772) );
  AOI22_X1 U9489 ( .A1(n7741), .A2(n7940), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7769) );
  NAND2_X1 U9490 ( .A1(n7944), .A2(n8167), .ZN(n7768) );
  OAI211_X1 U9491 ( .C1(n7847), .C2(n7942), .A(n7769), .B(n7768), .ZN(n7770)
         );
  AOI21_X1 U9492 ( .B1(n8388), .B2(n7930), .A(n7770), .ZN(n7771) );
  OAI21_X1 U9493 ( .B1(n7772), .B2(n7932), .A(n7771), .ZN(P2_U3156) );
  OAI211_X1 U9494 ( .C1(n7775), .C2(n7774), .A(n7773), .B(n7934), .ZN(n7780)
         );
  AOI21_X1 U9495 ( .B1(n7930), .B2(n9751), .A(n7776), .ZN(n7779) );
  AOI22_X1 U9496 ( .A1(n7940), .A2(n9744), .B1(n7925), .B2(n9746), .ZN(n7778)
         );
  OR2_X1 U9497 ( .A1(n7928), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7777) );
  NAND4_X1 U9498 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(
        P2_U3158) );
  INV_X1 U9499 ( .A(n8330), .ZN(n7789) );
  AOI211_X1 U9500 ( .C1(n7783), .C2(n7782), .A(n7932), .B(n7781), .ZN(n7784)
         );
  INV_X1 U9501 ( .A(n7784), .ZN(n7788) );
  NAND2_X1 U9502 ( .A1(n7940), .A2(n8215), .ZN(n7785) );
  NAND2_X1 U9503 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8077) );
  OAI211_X1 U9504 ( .C1(n8211), .C2(n7942), .A(n7785), .B(n8077), .ZN(n7786)
         );
  AOI21_X1 U9505 ( .B1(n8217), .B2(n7944), .A(n7786), .ZN(n7787) );
  OAI211_X1 U9506 ( .C1(n7789), .C2(n7947), .A(n7788), .B(n7787), .ZN(P2_U3159) );
  NOR2_X1 U9507 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  XOR2_X1 U9508 ( .A(n7796), .B(n7795), .Z(n7797) );
  XNOR2_X1 U9509 ( .A(n7798), .B(n7797), .ZN(n7804) );
  NOR2_X1 U9510 ( .A1(n7928), .A2(n8106), .ZN(n7802) );
  AOI22_X1 U9511 ( .A1(n7940), .A2(n8126), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7799) );
  OAI21_X1 U9512 ( .B1(n7800), .B2(n7942), .A(n7799), .ZN(n7801) );
  AOI211_X1 U9513 ( .C1(n8111), .C2(n7930), .A(n7802), .B(n7801), .ZN(n7803)
         );
  OAI21_X1 U9514 ( .B1(n7804), .B2(n7932), .A(n7803), .ZN(P2_U3160) );
  XOR2_X1 U9515 ( .A(n7806), .B(n7805), .Z(n7811) );
  AOI22_X1 U9516 ( .A1(n7741), .A2(n7925), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7808) );
  NAND2_X1 U9517 ( .A1(n7944), .A2(n8194), .ZN(n7807) );
  OAI211_X1 U9518 ( .C1(n8211), .C2(n7893), .A(n7808), .B(n7807), .ZN(n7809)
         );
  AOI21_X1 U9519 ( .B1(n8399), .B2(n7930), .A(n7809), .ZN(n7810) );
  OAI21_X1 U9520 ( .B1(n7811), .B2(n7932), .A(n7810), .ZN(P2_U3163) );
  XNOR2_X1 U9521 ( .A(n7813), .B(n7812), .ZN(n7819) );
  OAI21_X1 U9522 ( .B1(n7893), .B2(n8287), .A(n7814), .ZN(n7815) );
  AOI21_X1 U9523 ( .B1(n7925), .B2(n8275), .A(n7815), .ZN(n7816) );
  OAI21_X1 U9524 ( .B1(n8289), .B2(n7928), .A(n7816), .ZN(n7817) );
  AOI21_X1 U9525 ( .B1(n9815), .B2(n7930), .A(n7817), .ZN(n7818) );
  OAI21_X1 U9526 ( .B1(n7819), .B2(n7932), .A(n7818), .ZN(P2_U3164) );
  XOR2_X1 U9527 ( .A(n7821), .B(n7820), .Z(n7827) );
  AOI22_X1 U9528 ( .A1(n7925), .A2(n8140), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7823) );
  NAND2_X1 U9529 ( .A1(n7940), .A2(n8164), .ZN(n7822) );
  OAI211_X1 U9530 ( .C1(n8141), .C2(n7928), .A(n7823), .B(n7822), .ZN(n7824)
         );
  AOI21_X1 U9531 ( .B1(n7825), .B2(n7930), .A(n7824), .ZN(n7826) );
  OAI21_X1 U9532 ( .B1(n7827), .B2(n7932), .A(n7826), .ZN(P2_U3165) );
  INV_X1 U9533 ( .A(n8422), .ZN(n7836) );
  OAI211_X1 U9534 ( .C1(n7830), .C2(n7829), .A(n7828), .B(n7934), .ZN(n7835)
         );
  NOR2_X1 U9535 ( .A1(n7831), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8025) );
  AOI21_X1 U9536 ( .B1(n7925), .B2(n8228), .A(n8025), .ZN(n7832) );
  OAI21_X1 U9537 ( .B1(n7893), .B2(n8253), .A(n7832), .ZN(n7833) );
  AOI21_X1 U9538 ( .B1(n8259), .B2(n7944), .A(n7833), .ZN(n7834) );
  OAI211_X1 U9539 ( .C1(n7836), .C2(n7947), .A(n7835), .B(n7834), .ZN(P2_U3166) );
  AOI21_X1 U9540 ( .B1(n7838), .B2(n7837), .A(n7911), .ZN(n7843) );
  AOI22_X1 U9541 ( .A1(n7925), .A2(n8215), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7840) );
  NAND2_X1 U9542 ( .A1(n7944), .A2(n8244), .ZN(n7839) );
  OAI211_X1 U9543 ( .C1(n7893), .C2(n8242), .A(n7840), .B(n7839), .ZN(n7841)
         );
  AOI21_X1 U9544 ( .B1(n8339), .B2(n7930), .A(n7841), .ZN(n7842) );
  OAI21_X1 U9545 ( .B1(n7843), .B2(n7932), .A(n7842), .ZN(P2_U3168) );
  OAI22_X1 U9546 ( .A1(n7846), .A2(n8178), .B1(n7845), .B2(n7844), .ZN(n7850)
         );
  XNOR2_X1 U9547 ( .A(n7848), .B(n7847), .ZN(n7849) );
  XNOR2_X1 U9548 ( .A(n7850), .B(n7849), .ZN(n7856) );
  NAND2_X1 U9549 ( .A1(n8178), .A2(n7940), .ZN(n7853) );
  AOI22_X1 U9550 ( .A1(n7925), .A2(n8149), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7852) );
  OAI211_X1 U9551 ( .C1(n8151), .C2(n7928), .A(n7853), .B(n7852), .ZN(n7854)
         );
  AOI21_X1 U9552 ( .B1(n8382), .B2(n7930), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9553 ( .B1(n7856), .B2(n7932), .A(n7855), .ZN(P2_U3169) );
  OAI21_X1 U9554 ( .B1(n7858), .B2(n7857), .A(n6972), .ZN(n7859) );
  NAND2_X1 U9555 ( .A1(n7859), .A2(n7934), .ZN(n7866) );
  AOI21_X1 U9556 ( .B1(n7930), .B2(n7861), .A(n7860), .ZN(n7865) );
  AOI22_X1 U9557 ( .A1(n7925), .A2(n7956), .B1(n7940), .B2(n7957), .ZN(n7864)
         );
  OR2_X1 U9558 ( .A1(n7928), .A2(n7862), .ZN(n7863) );
  NAND4_X1 U9559 ( .A1(n7866), .A2(n7865), .A3(n7864), .A4(n7863), .ZN(
        P2_U3170) );
  OAI21_X1 U9560 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7870) );
  NAND2_X1 U9561 ( .A1(n7870), .A2(n7934), .ZN(n7874) );
  INV_X1 U9562 ( .A(n7892), .ZN(n8205) );
  AOI22_X1 U9563 ( .A1(n8205), .A2(n7925), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7871) );
  OAI21_X1 U9564 ( .B1(n7915), .B2(n7893), .A(n7871), .ZN(n7872) );
  AOI21_X1 U9565 ( .B1(n8208), .B2(n7944), .A(n7872), .ZN(n7873) );
  OAI211_X1 U9566 ( .C1(n7875), .C2(n7947), .A(n7874), .B(n7873), .ZN(P2_U3173) );
  INV_X1 U9567 ( .A(n7876), .ZN(n7877) );
  NOR2_X1 U9568 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  XNOR2_X1 U9569 ( .A(n7880), .B(n7879), .ZN(n7886) );
  NOR2_X1 U9570 ( .A1(n7942), .A2(n9549), .ZN(n7881) );
  AOI211_X1 U9571 ( .C1(n7940), .C2(n7951), .A(n7882), .B(n7881), .ZN(n7883)
         );
  OAI21_X1 U9572 ( .B1(n9541), .B2(n7928), .A(n7883), .ZN(n7884) );
  AOI21_X1 U9573 ( .B1(n9538), .B2(n7930), .A(n7884), .ZN(n7885) );
  OAI21_X1 U9574 ( .B1(n7886), .B2(n7932), .A(n7885), .ZN(P2_U3174) );
  OAI211_X1 U9575 ( .C1(n7889), .C2(n7888), .A(n7887), .B(n7934), .ZN(n7897)
         );
  INV_X1 U9576 ( .A(n8180), .ZN(n7890) );
  NOR2_X1 U9577 ( .A1(n7928), .A2(n7890), .ZN(n7895) );
  INV_X1 U9578 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7891) );
  OAI22_X1 U9579 ( .A1(n7893), .A2(n7892), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7891), .ZN(n7894) );
  AOI211_X1 U9580 ( .C1(n7925), .C2(n8178), .A(n7895), .B(n7894), .ZN(n7896)
         );
  OAI211_X1 U9581 ( .C1(n7898), .C2(n7947), .A(n7897), .B(n7896), .ZN(P2_U3175) );
  NOR2_X1 U9582 ( .A1(n7942), .A2(n9547), .ZN(n7899) );
  AOI211_X1 U9583 ( .C1(n7940), .C2(n7953), .A(n7900), .B(n7899), .ZN(n7901)
         );
  OAI21_X1 U9584 ( .B1(n7902), .B2(n7928), .A(n7901), .ZN(n7906) );
  AOI211_X1 U9585 ( .C1(n7904), .C2(n7903), .A(n7932), .B(n4372), .ZN(n7905)
         );
  AOI211_X1 U9586 ( .C1(n9808), .C2(n7930), .A(n7906), .B(n7905), .ZN(n7907)
         );
  INV_X1 U9587 ( .A(n7907), .ZN(P2_U3176) );
  INV_X1 U9588 ( .A(n7908), .ZN(n7913) );
  NOR3_X1 U9589 ( .A1(n7911), .A2(n7910), .A3(n7909), .ZN(n7912) );
  OAI21_X1 U9590 ( .B1(n7913), .B2(n7912), .A(n7934), .ZN(n7918) );
  NAND2_X1 U9591 ( .A1(n7940), .A2(n8228), .ZN(n7914) );
  NAND2_X1 U9592 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8053) );
  OAI211_X1 U9593 ( .C1(n7915), .C2(n7942), .A(n7914), .B(n8053), .ZN(n7916)
         );
  AOI21_X1 U9594 ( .B1(n8232), .B2(n7944), .A(n7916), .ZN(n7917) );
  OAI211_X1 U9595 ( .C1(n7919), .C2(n7947), .A(n7918), .B(n7917), .ZN(P2_U3178) );
  INV_X1 U9596 ( .A(n7921), .ZN(n7922) );
  NOR2_X1 U9597 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  XNOR2_X1 U9598 ( .A(n7920), .B(n7924), .ZN(n7933) );
  AOI22_X1 U9599 ( .A1(n7940), .A2(n8149), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7927) );
  NAND2_X1 U9600 ( .A1(n7925), .A2(n8126), .ZN(n7926) );
  OAI211_X1 U9601 ( .C1(n8129), .C2(n7928), .A(n7927), .B(n7926), .ZN(n7929)
         );
  AOI21_X1 U9602 ( .B1(n8131), .B2(n7930), .A(n7929), .ZN(n7931) );
  OAI21_X1 U9603 ( .B1(n7933), .B2(n7932), .A(n7931), .ZN(P2_U3180) );
  OAI211_X1 U9604 ( .C1(n7937), .C2(n7936), .A(n7935), .B(n7934), .ZN(n7946)
         );
  INV_X1 U9605 ( .A(n7938), .ZN(n8269) );
  AND2_X1 U9606 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7999) );
  AOI21_X1 U9607 ( .B1(n7940), .B2(n8266), .A(n7999), .ZN(n7941) );
  OAI21_X1 U9608 ( .B1(n8242), .B2(n7942), .A(n7941), .ZN(n7943) );
  AOI21_X1 U9609 ( .B1(n8269), .B2(n7944), .A(n7943), .ZN(n7945) );
  OAI211_X1 U9610 ( .C1(n7948), .C2(n7947), .A(n7946), .B(n7945), .ZN(P2_U3181) );
  MUX2_X1 U9611 ( .A(n8091), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8051), .Z(
        P2_U3522) );
  MUX2_X1 U9612 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n7949), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9613 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n7950), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9614 ( .A(n8126), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8051), .Z(
        P2_U3518) );
  MUX2_X1 U9615 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8140), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9616 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8149), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9617 ( .A(n8164), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8051), .Z(
        P2_U3515) );
  MUX2_X1 U9618 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8178), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9619 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n7741), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9620 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8205), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9621 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8191), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9622 ( .A(n8229), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8051), .Z(
        P2_U3510) );
  MUX2_X1 U9623 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8215), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9624 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8228), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9625 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8265), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9626 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7729), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9627 ( .A(n8266), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8051), .Z(
        P2_U3505) );
  MUX2_X1 U9628 ( .A(n8275), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8051), .Z(
        P2_U3504) );
  MUX2_X1 U9629 ( .A(n7951), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8051), .Z(
        P2_U3503) );
  MUX2_X1 U9630 ( .A(n7952), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8051), .Z(
        P2_U3502) );
  MUX2_X1 U9631 ( .A(n7953), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8051), .Z(
        P2_U3501) );
  MUX2_X1 U9632 ( .A(n9730), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8051), .Z(
        P2_U3500) );
  MUX2_X1 U9633 ( .A(n7954), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8051), .Z(
        P2_U3499) );
  MUX2_X1 U9634 ( .A(n9729), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8051), .Z(
        P2_U3498) );
  MUX2_X1 U9635 ( .A(n7955), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8051), .Z(
        P2_U3497) );
  MUX2_X1 U9636 ( .A(n7956), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8051), .Z(
        P2_U3496) );
  MUX2_X1 U9637 ( .A(n9746), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8051), .Z(
        P2_U3495) );
  MUX2_X1 U9638 ( .A(n7957), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8051), .Z(
        P2_U3494) );
  MUX2_X1 U9639 ( .A(n9744), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8051), .Z(
        P2_U3493) );
  MUX2_X1 U9640 ( .A(n5809), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8051), .Z(
        P2_U3492) );
  MUX2_X1 U9641 ( .A(n7958), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8051), .Z(
        P2_U3491) );
  NAND2_X1 U9642 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7990), .ZN(n7962) );
  OAI21_X1 U9643 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7990), .A(n7962), .ZN(
        n7963) );
  AOI21_X1 U9644 ( .B1(n7964), .B2(n7963), .A(n7988), .ZN(n7987) );
  AOI22_X1 U9645 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7990), .B1(n7975), .B2(
        n8348), .ZN(n7970) );
  NAND2_X1 U9646 ( .A1(n7966), .A2(n7965), .ZN(n7968) );
  NAND2_X1 U9647 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  OAI21_X1 U9648 ( .B1(n7970), .B2(n7969), .A(n7991), .ZN(n7985) );
  NAND2_X1 U9649 ( .A1(n9713), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7971) );
  OAI211_X1 U9650 ( .C1(n8050), .C2(n7990), .A(n7972), .B(n7971), .ZN(n7984)
         );
  INV_X1 U9651 ( .A(n7973), .ZN(n7980) );
  MUX2_X1 U9652 ( .A(n7974), .B(n8348), .S(n4398), .Z(n7976) );
  NAND2_X1 U9653 ( .A1(n7976), .A2(n7975), .ZN(n7994) );
  INV_X1 U9654 ( .A(n7976), .ZN(n7977) );
  NAND2_X1 U9655 ( .A1(n7977), .A2(n7990), .ZN(n7978) );
  AND2_X1 U9656 ( .A1(n7994), .A2(n7978), .ZN(n7979) );
  OAI21_X1 U9657 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(n7995) );
  OR3_X1 U9658 ( .A1(n7981), .A2(n7980), .A3(n7979), .ZN(n7982) );
  AOI21_X1 U9659 ( .B1(n7995), .B2(n7982), .A(n8082), .ZN(n7983) );
  AOI211_X1 U9660 ( .C1(n7985), .C2(n9720), .A(n7984), .B(n7983), .ZN(n7986)
         );
  OAI21_X1 U9661 ( .B1(n7987), .B2(n8086), .A(n7986), .ZN(P2_U3196) );
  AOI21_X1 U9662 ( .B1(n10021), .B2(n7989), .A(n4366), .ZN(n8005) );
  NAND2_X1 U9663 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7990), .ZN(n7992) );
  XNOR2_X1 U9664 ( .A(n8006), .B(n8010), .ZN(n7993) );
  NAND2_X1 U9665 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7993), .ZN(n8011) );
  OAI21_X1 U9666 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n7993), .A(n8011), .ZN(
        n8003) );
  NAND2_X1 U9667 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  MUX2_X1 U9668 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4398), .Z(n8017) );
  XNOR2_X1 U9669 ( .A(n8017), .B(n8006), .ZN(n7996) );
  NAND2_X1 U9670 ( .A1(n7997), .A2(n7996), .ZN(n8015) );
  OAI21_X1 U9671 ( .B1(n7997), .B2(n7996), .A(n8015), .ZN(n7998) );
  NAND2_X1 U9672 ( .A1(n7998), .A2(n9887), .ZN(n8001) );
  AOI21_X1 U9673 ( .B1(n9713), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7999), .ZN(
        n8000) );
  OAI211_X1 U9674 ( .C1(n8050), .C2(n8016), .A(n8001), .B(n8000), .ZN(n8002)
         );
  AOI21_X1 U9675 ( .B1(n9720), .B2(n8003), .A(n8002), .ZN(n8004) );
  OAI21_X1 U9676 ( .B1(n8005), .B2(n8086), .A(n8004), .ZN(P2_U3197) );
  AOI22_X1 U9677 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8033), .B1(n8036), .B2(
        n8258), .ZN(n8008) );
  AOI21_X1 U9678 ( .B1(n8009), .B2(n8008), .A(n8035), .ZN(n8031) );
  AOI22_X1 U9679 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8036), .B1(n8033), .B2(
        n8341), .ZN(n8014) );
  NAND2_X1 U9680 ( .A1(n8016), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U9681 ( .A1(n8014), .A2(n8013), .ZN(n8032) );
  OAI21_X1 U9682 ( .B1(n8014), .B2(n8013), .A(n8032), .ZN(n8029) );
  OAI21_X1 U9683 ( .B1(n8017), .B2(n8016), .A(n8015), .ZN(n8021) );
  MUX2_X1 U9684 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4398), .Z(n8018) );
  NAND2_X1 U9685 ( .A1(n8018), .A2(n8036), .ZN(n8022) );
  NAND2_X1 U9686 ( .A1(n8021), .A2(n8022), .ZN(n8044) );
  INV_X1 U9687 ( .A(n8018), .ZN(n8019) );
  NAND2_X1 U9688 ( .A1(n8019), .A2(n8033), .ZN(n8043) );
  INV_X1 U9689 ( .A(n8043), .ZN(n8020) );
  NOR2_X1 U9690 ( .A1(n8044), .A2(n8020), .ZN(n8024) );
  AOI21_X1 U9691 ( .B1(n8022), .B2(n8043), .A(n8021), .ZN(n8023) );
  OAI21_X1 U9692 ( .B1(n8024), .B2(n8023), .A(n9887), .ZN(n8027) );
  AOI21_X1 U9693 ( .B1(n9713), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8025), .ZN(
        n8026) );
  OAI211_X1 U9694 ( .C1(n8036), .C2(n8050), .A(n8027), .B(n8026), .ZN(n8028)
         );
  AOI21_X1 U9695 ( .B1(n9720), .B2(n8029), .A(n8028), .ZN(n8030) );
  OAI21_X1 U9696 ( .B1(n8031), .B2(n8086), .A(n8030), .ZN(P2_U3198) );
  XOR2_X1 U9697 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8072), .Z(n8067) );
  XNOR2_X1 U9698 ( .A(n9714), .B(n8034), .ZN(n9716) );
  XOR2_X1 U9699 ( .A(n8067), .B(n8068), .Z(n8061) );
  NOR2_X1 U9700 ( .A1(n8072), .A2(n8231), .ZN(n8062) );
  AOI21_X1 U9701 ( .B1(n8072), .B2(n8231), .A(n8062), .ZN(n8039) );
  INV_X1 U9702 ( .A(n8064), .ZN(n8042) );
  NOR3_X1 U9703 ( .A1(n8040), .A2(n9722), .A3(n8039), .ZN(n8041) );
  OAI21_X1 U9704 ( .B1(n8042), .B2(n8041), .A(n9874), .ZN(n8060) );
  NAND2_X1 U9705 ( .A1(n8044), .A2(n8043), .ZN(n9718) );
  MUX2_X1 U9706 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4398), .Z(n8045) );
  XNOR2_X1 U9707 ( .A(n8045), .B(n9714), .ZN(n9717) );
  INV_X1 U9708 ( .A(n8045), .ZN(n8046) );
  AOI22_X1 U9709 ( .A1(n9718), .A2(n9717), .B1(n9714), .B2(n8046), .ZN(n8048)
         );
  MUX2_X1 U9710 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4398), .Z(n8047) );
  NOR2_X1 U9711 ( .A1(n8048), .A2(n8047), .ZN(n8070) );
  NAND2_X1 U9712 ( .A1(n8048), .A2(n8047), .ZN(n8071) );
  INV_X1 U9713 ( .A(n8071), .ZN(n8049) );
  NOR2_X1 U9714 ( .A1(n8070), .A2(n8049), .ZN(n8055) );
  INV_X1 U9715 ( .A(n8055), .ZN(n8052) );
  OAI21_X1 U9716 ( .B1(n8052), .B2(n8051), .A(n8050), .ZN(n8058) );
  INV_X1 U9717 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8054) );
  OAI21_X1 U9718 ( .B1(n9880), .B2(n8054), .A(n8053), .ZN(n8057) );
  NOR3_X1 U9719 ( .A1(n8055), .A2(n8072), .A3(n8082), .ZN(n8056) );
  AOI211_X1 U9720 ( .C1(n8072), .C2(n8058), .A(n8057), .B(n8056), .ZN(n8059)
         );
  OAI211_X1 U9721 ( .C1(n8061), .C2(n9891), .A(n8060), .B(n8059), .ZN(P2_U3200) );
  INV_X1 U9722 ( .A(n8062), .ZN(n8063) );
  NAND2_X1 U9723 ( .A1(n8064), .A2(n8063), .ZN(n8066) );
  XNOR2_X1 U9724 ( .A(n8080), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8074) );
  XNOR2_X1 U9725 ( .A(n8069), .B(n8074), .ZN(n8085) );
  AOI21_X1 U9726 ( .B1(n8072), .B2(n8071), .A(n8070), .ZN(n8076) );
  MUX2_X1 U9727 ( .A(n8074), .B(n4381), .S(n8073), .Z(n8075) );
  XNOR2_X1 U9728 ( .A(n8076), .B(n8075), .ZN(n8083) );
  OAI21_X1 U9729 ( .B1(n9880), .B2(n8078), .A(n8077), .ZN(n8079) );
  AOI21_X1 U9730 ( .B1(n8080), .B2(n9882), .A(n8079), .ZN(n8081) );
  OAI21_X1 U9731 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8084) );
  INV_X1 U9732 ( .A(n8087), .ZN(n8088) );
  NAND2_X1 U9733 ( .A1(n9752), .A2(n8088), .ZN(n8098) );
  INV_X1 U9734 ( .A(n8089), .ZN(n8090) );
  NAND2_X1 U9735 ( .A1(n8091), .A2(n8090), .ZN(n8360) );
  AOI21_X1 U9736 ( .B1(n8098), .B2(n8360), .A(n9757), .ZN(n8093) );
  AOI21_X1 U9737 ( .B1(n9757), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8093), .ZN(
        n8092) );
  OAI21_X1 U9738 ( .B1(n8362), .B2(n8095), .A(n8092), .ZN(P2_U3202) );
  AOI21_X1 U9739 ( .B1(n9757), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8093), .ZN(
        n8094) );
  OAI21_X1 U9740 ( .B1(n8303), .B2(n8095), .A(n8094), .ZN(P2_U3203) );
  NAND2_X1 U9741 ( .A1(n8097), .A2(n8268), .ZN(n8103) );
  OAI21_X1 U9742 ( .B1(n8268), .B2(n8099), .A(n8098), .ZN(n8100) );
  AOI21_X1 U9743 ( .B1(n8101), .B2(n9750), .A(n8100), .ZN(n8102) );
  OAI211_X1 U9744 ( .C1(n8105), .C2(n8104), .A(n8103), .B(n8102), .ZN(P2_U3204) );
  OAI22_X1 U9745 ( .A1(n8291), .A2(n8107), .B1(n8106), .B2(n9540), .ZN(n8110)
         );
  NOR2_X1 U9746 ( .A1(n8108), .A2(n8272), .ZN(n8109) );
  AOI211_X1 U9747 ( .C1(n9750), .C2(n8111), .A(n8110), .B(n8109), .ZN(n8112)
         );
  OAI21_X1 U9748 ( .B1(n8113), .B2(n9757), .A(n8112), .ZN(P2_U3205) );
  INV_X1 U9749 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8115) );
  OAI22_X1 U9750 ( .A1(n8291), .A2(n8115), .B1(n8114), .B2(n9540), .ZN(n8118)
         );
  NOR2_X1 U9751 ( .A1(n8116), .A2(n8272), .ZN(n8117) );
  AOI211_X1 U9752 ( .C1(n9750), .C2(n8119), .A(n8118), .B(n8117), .ZN(n8120)
         );
  OAI21_X1 U9753 ( .B1(n8121), .B2(n9757), .A(n8120), .ZN(P2_U3206) );
  XNOR2_X1 U9754 ( .A(n8123), .B(n8122), .ZN(n8369) );
  INV_X1 U9755 ( .A(n8369), .ZN(n8134) );
  XNOR2_X1 U9756 ( .A(n8124), .B(n8125), .ZN(n8127) );
  AOI222_X1 U9757 ( .A1(n9748), .A2(n8127), .B1(n8149), .B2(n9743), .C1(n8126), 
        .C2(n9745), .ZN(n8367) );
  MUX2_X1 U9758 ( .A(n8128), .B(n8367), .S(n8268), .Z(n8133) );
  INV_X1 U9759 ( .A(n8129), .ZN(n8130) );
  AOI22_X1 U9760 ( .A1(n8131), .A2(n9750), .B1(n9752), .B2(n8130), .ZN(n8132)
         );
  OAI211_X1 U9761 ( .C1(n8134), .C2(n8272), .A(n8133), .B(n8132), .ZN(P2_U3207) );
  OR2_X1 U9762 ( .A1(n8148), .A2(n8135), .ZN(n8137) );
  NAND2_X1 U9763 ( .A1(n8137), .A2(n8136), .ZN(n8139) );
  INV_X1 U9764 ( .A(n8373), .ZN(n8143) );
  OAI22_X1 U9765 ( .A1(n8379), .A2(n8278), .B1(n8141), .B2(n9540), .ZN(n8142)
         );
  OAI21_X1 U9766 ( .B1(n8143), .B2(n8142), .A(n8291), .ZN(n8147) );
  XNOR2_X1 U9767 ( .A(n8145), .B(n8144), .ZN(n8375) );
  AOI22_X1 U9768 ( .A1(n8375), .A2(n9754), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9757), .ZN(n8146) );
  NAND2_X1 U9769 ( .A1(n8147), .A2(n8146), .ZN(P2_U3208) );
  XOR2_X1 U9770 ( .A(n8157), .B(n8148), .Z(n8150) );
  AOI222_X1 U9771 ( .A1(n9748), .A2(n8150), .B1(n8149), .B2(n9745), .C1(n8178), 
        .C2(n9743), .ZN(n8380) );
  INV_X1 U9772 ( .A(n8380), .ZN(n8154) );
  INV_X1 U9773 ( .A(n8382), .ZN(n8152) );
  OAI22_X1 U9774 ( .A1(n8152), .A2(n8278), .B1(n8151), .B2(n9540), .ZN(n8153)
         );
  OAI21_X1 U9775 ( .B1(n8154), .B2(n8153), .A(n8291), .ZN(n8160) );
  NAND2_X1 U9776 ( .A1(n8156), .A2(n8155), .ZN(n8158) );
  XNOR2_X1 U9777 ( .A(n8158), .B(n8157), .ZN(n8383) );
  AOI22_X1 U9778 ( .A1(n8383), .A2(n9754), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9757), .ZN(n8159) );
  NAND2_X1 U9779 ( .A1(n8160), .A2(n8159), .ZN(P2_U3209) );
  XNOR2_X1 U9780 ( .A(n8161), .B(n8162), .ZN(n8389) );
  INV_X1 U9781 ( .A(n8389), .ZN(n8170) );
  INV_X1 U9782 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8166) );
  XNOR2_X1 U9783 ( .A(n8163), .B(n8162), .ZN(n8165) );
  AOI222_X1 U9784 ( .A1(n9748), .A2(n8165), .B1(n8164), .B2(n9745), .C1(n7741), 
        .C2(n9743), .ZN(n8386) );
  MUX2_X1 U9785 ( .A(n8166), .B(n8386), .S(n8268), .Z(n8169) );
  AOI22_X1 U9786 ( .A1(n8388), .A2(n9750), .B1(n9752), .B2(n8167), .ZN(n8168)
         );
  OAI211_X1 U9787 ( .C1(n8170), .C2(n8272), .A(n8169), .B(n8168), .ZN(P2_U3210) );
  XNOR2_X1 U9788 ( .A(n8172), .B(n8171), .ZN(n8395) );
  INV_X1 U9789 ( .A(n8395), .ZN(n8183) );
  NAND3_X1 U9790 ( .A1(n8174), .A2(n8176), .A3(n8175), .ZN(n8177) );
  NAND2_X1 U9791 ( .A1(n8173), .A2(n8177), .ZN(n8179) );
  AOI222_X1 U9792 ( .A1(n9748), .A2(n8179), .B1(n8178), .B2(n9745), .C1(n8205), 
        .C2(n9743), .ZN(n8392) );
  MUX2_X1 U9793 ( .A(n9960), .B(n8392), .S(n8268), .Z(n8182) );
  AOI22_X1 U9794 ( .A1(n8394), .A2(n9750), .B1(n9752), .B2(n8180), .ZN(n8181)
         );
  OAI211_X1 U9795 ( .C1(n8183), .C2(n8272), .A(n8182), .B(n8181), .ZN(P2_U3211) );
  NAND2_X1 U9796 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  XNOR2_X1 U9797 ( .A(n8186), .B(n8187), .ZN(n8402) );
  INV_X1 U9798 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8193) );
  INV_X1 U9799 ( .A(n8187), .ZN(n8189) );
  NAND3_X1 U9800 ( .A1(n8203), .A2(n8189), .A3(n8188), .ZN(n8190) );
  NAND2_X1 U9801 ( .A1(n8174), .A2(n8190), .ZN(n8192) );
  AOI222_X1 U9802 ( .A1(n9748), .A2(n8192), .B1(n7741), .B2(n9745), .C1(n8191), 
        .C2(n9743), .ZN(n8398) );
  MUX2_X1 U9803 ( .A(n8193), .B(n8398), .S(n8268), .Z(n8196) );
  AOI22_X1 U9804 ( .A1(n8399), .A2(n9750), .B1(n9752), .B2(n8194), .ZN(n8195)
         );
  OAI211_X1 U9805 ( .C1(n8402), .C2(n8272), .A(n8196), .B(n8195), .ZN(P2_U3212) );
  NAND2_X1 U9806 ( .A1(n8197), .A2(n8198), .ZN(n8199) );
  XNOR2_X1 U9807 ( .A(n8199), .B(n8201), .ZN(n8408) );
  INV_X1 U9808 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8207) );
  INV_X1 U9809 ( .A(n8200), .ZN(n8212) );
  OAI21_X1 U9810 ( .B1(n8212), .B2(n8202), .A(n8201), .ZN(n8204) );
  NAND2_X1 U9811 ( .A1(n8204), .A2(n8203), .ZN(n8206) );
  AOI222_X1 U9812 ( .A1(n9748), .A2(n8206), .B1(n8205), .B2(n9745), .C1(n8229), 
        .C2(n9743), .ZN(n8403) );
  MUX2_X1 U9813 ( .A(n8207), .B(n8403), .S(n8268), .Z(n8210) );
  AOI22_X1 U9814 ( .A1(n8405), .A2(n9750), .B1(n9752), .B2(n8208), .ZN(n8209)
         );
  OAI211_X1 U9815 ( .C1(n8408), .C2(n8272), .A(n8210), .B(n8209), .ZN(P2_U3213) );
  NOR2_X1 U9816 ( .A1(n8211), .A2(n9550), .ZN(n8329) );
  AOI211_X1 U9817 ( .C1(n8218), .C2(n8213), .A(n9546), .B(n8212), .ZN(n8214)
         );
  AOI21_X1 U9818 ( .B1(n9743), .B2(n8215), .A(n8214), .ZN(n8334) );
  INV_X1 U9819 ( .A(n8334), .ZN(n8216) );
  AOI211_X1 U9820 ( .C1(n9752), .C2(n8217), .A(n8329), .B(n8216), .ZN(n8222)
         );
  AOI22_X1 U9821 ( .A1(n8330), .A2(n9750), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9757), .ZN(n8221) );
  OR2_X1 U9822 ( .A1(n8219), .A2(n8218), .ZN(n8331) );
  NAND3_X1 U9823 ( .A1(n8331), .A2(n9754), .A3(n8197), .ZN(n8220) );
  OAI211_X1 U9824 ( .C1(n8222), .C2(n9757), .A(n8221), .B(n8220), .ZN(P2_U3214) );
  NAND2_X1 U9825 ( .A1(n4416), .A2(n8223), .ZN(n8224) );
  XNOR2_X1 U9826 ( .A(n8224), .B(n8225), .ZN(n8413) );
  INV_X1 U9827 ( .A(n8413), .ZN(n8235) );
  OAI21_X1 U9828 ( .B1(n8227), .B2(n6133), .A(n8226), .ZN(n8230) );
  AOI222_X1 U9829 ( .A1(n9748), .A2(n8230), .B1(n8229), .B2(n9745), .C1(n8228), 
        .C2(n9743), .ZN(n8410) );
  MUX2_X1 U9830 ( .A(n8231), .B(n8410), .S(n8268), .Z(n8234) );
  AOI22_X1 U9831 ( .A1(n8412), .A2(n9750), .B1(n9752), .B2(n8232), .ZN(n8233)
         );
  OAI211_X1 U9832 ( .C1(n8235), .C2(n8272), .A(n8234), .B(n8233), .ZN(P2_U3215) );
  INV_X1 U9833 ( .A(n4416), .ZN(n8237) );
  AOI21_X1 U9834 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8419) );
  XNOR2_X1 U9835 ( .A(n8240), .B(n8239), .ZN(n8241) );
  OAI222_X1 U9836 ( .A1(n9550), .A2(n8243), .B1(n9548), .B2(n8242), .C1(n8241), 
        .C2(n9546), .ZN(n8338) );
  NAND2_X1 U9837 ( .A1(n8338), .A2(n8268), .ZN(n8249) );
  INV_X1 U9838 ( .A(n8244), .ZN(n8245) );
  OAI22_X1 U9839 ( .A1(n8291), .A2(n8246), .B1(n8245), .B2(n9540), .ZN(n8247)
         );
  AOI21_X1 U9840 ( .B1(n8339), .B2(n9750), .A(n8247), .ZN(n8248) );
  OAI211_X1 U9841 ( .C1(n8419), .C2(n8272), .A(n8249), .B(n8248), .ZN(P2_U3216) );
  XNOR2_X1 U9842 ( .A(n8250), .B(n8251), .ZN(n8426) );
  AOI21_X1 U9843 ( .B1(n8252), .B2(n8251), .A(n9546), .ZN(n8257) );
  OAI22_X1 U9844 ( .A1(n8254), .A2(n9550), .B1(n8253), .B2(n9548), .ZN(n8255)
         );
  AOI21_X1 U9845 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(n8420) );
  MUX2_X1 U9846 ( .A(n8258), .B(n8420), .S(n8268), .Z(n8261) );
  AOI22_X1 U9847 ( .A1(n8422), .A2(n9750), .B1(n9752), .B2(n8259), .ZN(n8260)
         );
  OAI211_X1 U9848 ( .C1(n8426), .C2(n8272), .A(n8261), .B(n8260), .ZN(P2_U3217) );
  XNOR2_X1 U9849 ( .A(n8262), .B(n8264), .ZN(n8430) );
  INV_X1 U9850 ( .A(n8430), .ZN(n8273) );
  XNOR2_X1 U9851 ( .A(n8263), .B(n8264), .ZN(n8267) );
  AOI222_X1 U9852 ( .A1(n9748), .A2(n8267), .B1(n8266), .B2(n9743), .C1(n8265), 
        .C2(n9745), .ZN(n8427) );
  MUX2_X1 U9853 ( .A(n10021), .B(n8427), .S(n8268), .Z(n8271) );
  AOI22_X1 U9854 ( .A1(n8429), .A2(n9750), .B1(n9752), .B2(n8269), .ZN(n8270)
         );
  OAI211_X1 U9855 ( .C1(n8273), .C2(n8272), .A(n8271), .B(n8270), .ZN(P2_U3218) );
  XOR2_X1 U9856 ( .A(n8274), .B(n8281), .Z(n8276) );
  AOI222_X1 U9857 ( .A1(n9748), .A2(n8276), .B1(n8275), .B2(n9743), .C1(n7729), 
        .C2(n9745), .ZN(n8433) );
  INV_X1 U9858 ( .A(n8433), .ZN(n8280) );
  OAI22_X1 U9859 ( .A1(n6125), .A2(n8278), .B1(n8277), .B2(n9540), .ZN(n8279)
         );
  OAI21_X1 U9860 ( .B1(n8280), .B2(n8279), .A(n8291), .ZN(n8284) );
  XNOR2_X1 U9861 ( .A(n8282), .B(n8281), .ZN(n8438) );
  AOI22_X1 U9862 ( .A1(n8438), .A2(n9754), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9757), .ZN(n8283) );
  NAND2_X1 U9863 ( .A1(n8284), .A2(n8283), .ZN(P2_U3219) );
  XOR2_X1 U9864 ( .A(n8293), .B(n8285), .Z(n8286) );
  OAI222_X1 U9865 ( .A1(n9550), .A2(n8288), .B1(n9548), .B2(n8287), .C1(n9546), 
        .C2(n8286), .ZN(n9813) );
  INV_X1 U9866 ( .A(n9813), .ZN(n8297) );
  OAI22_X1 U9867 ( .A1(n8291), .A2(n8290), .B1(n8289), .B2(n9540), .ZN(n8292)
         );
  AOI21_X1 U9868 ( .B1(n9815), .B2(n9750), .A(n8292), .ZN(n8296) );
  NAND2_X1 U9869 ( .A1(n8294), .A2(n8293), .ZN(n9810) );
  NAND3_X1 U9870 ( .A1(n9812), .A2(n9810), .A3(n9754), .ZN(n8295) );
  OAI211_X1 U9871 ( .C1(n8297), .C2(n9757), .A(n8296), .B(n8295), .ZN(P2_U3221) );
  NAND2_X1 U9872 ( .A1(n8298), .A2(n8349), .ZN(n8300) );
  INV_X1 U9873 ( .A(n8360), .ZN(n8299) );
  NAND2_X1 U9874 ( .A1(n4275), .A2(n8299), .ZN(n8301) );
  OAI211_X1 U9875 ( .C1(n4275), .C2(n7529), .A(n8300), .B(n8301), .ZN(P2_U3490) );
  NAND2_X1 U9876 ( .A1(n9833), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8302) );
  OAI211_X1 U9877 ( .C1(n8303), .C2(n8313), .A(n8302), .B(n8301), .ZN(P2_U3489) );
  OAI21_X1 U9878 ( .B1(n8306), .B2(n8313), .A(n8305), .ZN(P2_U3486) );
  MUX2_X1 U9879 ( .A(n8307), .B(n8367), .S(n4275), .Z(n8309) );
  NAND2_X1 U9880 ( .A1(n8369), .A2(n8350), .ZN(n8308) );
  OAI211_X1 U9881 ( .C1(n8372), .C2(n8313), .A(n8309), .B(n8308), .ZN(P2_U3485) );
  INV_X1 U9882 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8310) );
  MUX2_X1 U9883 ( .A(n8310), .B(n8373), .S(n4275), .Z(n8312) );
  NAND2_X1 U9884 ( .A1(n8375), .A2(n8350), .ZN(n8311) );
  OAI211_X1 U9885 ( .C1(n8379), .C2(n8313), .A(n8312), .B(n8311), .ZN(P2_U3484) );
  INV_X1 U9886 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8314) );
  MUX2_X1 U9887 ( .A(n8314), .B(n8380), .S(n4275), .Z(n8316) );
  AOI22_X1 U9888 ( .A1(n8383), .A2(n8350), .B1(n8349), .B2(n8382), .ZN(n8315)
         );
  NAND2_X1 U9889 ( .A1(n8316), .A2(n8315), .ZN(P2_U3483) );
  MUX2_X1 U9890 ( .A(n8317), .B(n8386), .S(n4275), .Z(n8319) );
  AOI22_X1 U9891 ( .A1(n8389), .A2(n8350), .B1(n8349), .B2(n8388), .ZN(n8318)
         );
  NAND2_X1 U9892 ( .A1(n8319), .A2(n8318), .ZN(P2_U3482) );
  INV_X1 U9893 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8320) );
  MUX2_X1 U9894 ( .A(n8320), .B(n8392), .S(n4275), .Z(n8322) );
  AOI22_X1 U9895 ( .A1(n8395), .A2(n8350), .B1(n8349), .B2(n8394), .ZN(n8321)
         );
  NAND2_X1 U9896 ( .A1(n8322), .A2(n8321), .ZN(P2_U3481) );
  INV_X1 U9897 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8323) );
  MUX2_X1 U9898 ( .A(n8323), .B(n8398), .S(n4275), .Z(n8325) );
  NAND2_X1 U9899 ( .A1(n8399), .A2(n8349), .ZN(n8324) );
  OAI211_X1 U9900 ( .C1(n8344), .C2(n8402), .A(n8325), .B(n8324), .ZN(P2_U3480) );
  INV_X1 U9901 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8326) );
  MUX2_X1 U9902 ( .A(n8326), .B(n8403), .S(n4275), .Z(n8328) );
  NAND2_X1 U9903 ( .A1(n8405), .A2(n8349), .ZN(n8327) );
  OAI211_X1 U9904 ( .C1(n8408), .C2(n8344), .A(n8328), .B(n8327), .ZN(P2_U3479) );
  AOI21_X1 U9905 ( .B1(n8330), .B2(n9816), .A(n8329), .ZN(n8333) );
  NAND3_X1 U9906 ( .A1(n8331), .A2(n8197), .A3(n9811), .ZN(n8332) );
  NAND3_X1 U9907 ( .A1(n8334), .A2(n8333), .A3(n8332), .ZN(n8409) );
  MUX2_X1 U9908 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8409), .S(n4275), .Z(
        P2_U3478) );
  MUX2_X1 U9909 ( .A(n8335), .B(n8410), .S(n4275), .Z(n8337) );
  AOI22_X1 U9910 ( .A1(n8413), .A2(n8350), .B1(n8349), .B2(n8412), .ZN(n8336)
         );
  NAND2_X1 U9911 ( .A1(n8337), .A2(n8336), .ZN(P2_U3477) );
  AOI21_X1 U9912 ( .B1(n9816), .B2(n8339), .A(n8338), .ZN(n8416) );
  MUX2_X1 U9913 ( .A(n9930), .B(n8416), .S(n4275), .Z(n8340) );
  OAI21_X1 U9914 ( .B1(n8419), .B2(n8344), .A(n8340), .ZN(P2_U3476) );
  MUX2_X1 U9915 ( .A(n8341), .B(n8420), .S(n4275), .Z(n8343) );
  NAND2_X1 U9916 ( .A1(n8422), .A2(n8349), .ZN(n8342) );
  OAI211_X1 U9917 ( .C1(n8426), .C2(n8344), .A(n8343), .B(n8342), .ZN(P2_U3475) );
  MUX2_X1 U9918 ( .A(n8345), .B(n8427), .S(n4275), .Z(n8347) );
  AOI22_X1 U9919 ( .A1(n8430), .A2(n8350), .B1(n8349), .B2(n8429), .ZN(n8346)
         );
  NAND2_X1 U9920 ( .A1(n8347), .A2(n8346), .ZN(P2_U3474) );
  MUX2_X1 U9921 ( .A(n8348), .B(n8433), .S(n4275), .Z(n8352) );
  AOI22_X1 U9922 ( .A1(n8438), .A2(n8350), .B1(n8349), .B2(n8435), .ZN(n8351)
         );
  NAND2_X1 U9923 ( .A1(n8352), .A2(n8351), .ZN(P2_U3473) );
  OAI21_X1 U9924 ( .B1(n8354), .B2(n9786), .A(n8353), .ZN(n8356) );
  NAND2_X1 U9925 ( .A1(n5830), .A2(n9816), .ZN(n8355) );
  INV_X1 U9926 ( .A(n9760), .ZN(n8358) );
  MUX2_X1 U9927 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8358), .S(n4275), .Z(
        P2_U3461) );
  MUX2_X1 U9928 ( .A(n8359), .B(P2_REG1_REG_0__SCAN_IN), .S(n9833), .Z(
        P2_U3459) );
  NOR2_X1 U9929 ( .A1(n9819), .A2(n8360), .ZN(n8364) );
  AOI21_X1 U9930 ( .B1(n9819), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8364), .ZN(
        n8361) );
  OAI21_X1 U9931 ( .B1(n8362), .B2(n8378), .A(n8361), .ZN(P2_U3458) );
  NAND2_X1 U9932 ( .A1(n8363), .A2(n8436), .ZN(n8366) );
  INV_X1 U9933 ( .A(n8364), .ZN(n8365) );
  OAI211_X1 U9934 ( .C1(n6225), .C2(n9817), .A(n8366), .B(n8365), .ZN(P2_U3457) );
  INV_X1 U9935 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8368) );
  MUX2_X1 U9936 ( .A(n8368), .B(n8367), .S(n9817), .Z(n8371) );
  NAND2_X1 U9937 ( .A1(n8369), .A2(n8437), .ZN(n8370) );
  OAI211_X1 U9938 ( .C1(n8372), .C2(n8378), .A(n8371), .B(n8370), .ZN(P2_U3453) );
  MUX2_X1 U9939 ( .A(n8374), .B(n8373), .S(n9817), .Z(n8377) );
  NAND2_X1 U9940 ( .A1(n8375), .A2(n8437), .ZN(n8376) );
  OAI211_X1 U9941 ( .C1(n8379), .C2(n8378), .A(n8377), .B(n8376), .ZN(P2_U3452) );
  INV_X1 U9942 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8381) );
  MUX2_X1 U9943 ( .A(n8381), .B(n8380), .S(n9817), .Z(n8385) );
  AOI22_X1 U9944 ( .A1(n8383), .A2(n8437), .B1(n8436), .B2(n8382), .ZN(n8384)
         );
  NAND2_X1 U9945 ( .A1(n8385), .A2(n8384), .ZN(P2_U3451) );
  INV_X1 U9946 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8387) );
  MUX2_X1 U9947 ( .A(n8387), .B(n8386), .S(n9817), .Z(n8391) );
  AOI22_X1 U9948 ( .A1(n8389), .A2(n8437), .B1(n8436), .B2(n8388), .ZN(n8390)
         );
  NAND2_X1 U9949 ( .A1(n8391), .A2(n8390), .ZN(P2_U3450) );
  INV_X1 U9950 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8393) );
  MUX2_X1 U9951 ( .A(n8393), .B(n8392), .S(n9817), .Z(n8397) );
  AOI22_X1 U9952 ( .A1(n8395), .A2(n8437), .B1(n8436), .B2(n8394), .ZN(n8396)
         );
  NAND2_X1 U9953 ( .A1(n8397), .A2(n8396), .ZN(P2_U3449) );
  INV_X1 U9954 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U9955 ( .A(n9965), .B(n8398), .S(n9817), .Z(n8401) );
  NAND2_X1 U9956 ( .A1(n8399), .A2(n8436), .ZN(n8400) );
  OAI211_X1 U9957 ( .C1(n8402), .C2(n8425), .A(n8401), .B(n8400), .ZN(P2_U3448) );
  INV_X1 U9958 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8404) );
  MUX2_X1 U9959 ( .A(n8404), .B(n8403), .S(n9817), .Z(n8407) );
  NAND2_X1 U9960 ( .A1(n8405), .A2(n8436), .ZN(n8406) );
  OAI211_X1 U9961 ( .C1(n8408), .C2(n8425), .A(n8407), .B(n8406), .ZN(P2_U3447) );
  MUX2_X1 U9962 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8409), .S(n9817), .Z(
        P2_U3446) );
  MUX2_X1 U9963 ( .A(n8411), .B(n8410), .S(n9817), .Z(n8415) );
  AOI22_X1 U9964 ( .A1(n8413), .A2(n8437), .B1(n8436), .B2(n8412), .ZN(n8414)
         );
  NAND2_X1 U9965 ( .A1(n8415), .A2(n8414), .ZN(P2_U3444) );
  MUX2_X1 U9966 ( .A(n8417), .B(n8416), .S(n9817), .Z(n8418) );
  OAI21_X1 U9967 ( .B1(n8419), .B2(n8425), .A(n8418), .ZN(P2_U3441) );
  INV_X1 U9968 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8421) );
  MUX2_X1 U9969 ( .A(n8421), .B(n8420), .S(n9817), .Z(n8424) );
  NAND2_X1 U9970 ( .A1(n8422), .A2(n8436), .ZN(n8423) );
  OAI211_X1 U9971 ( .C1(n8426), .C2(n8425), .A(n8424), .B(n8423), .ZN(P2_U3438) );
  INV_X1 U9972 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8428) );
  MUX2_X1 U9973 ( .A(n8428), .B(n8427), .S(n9817), .Z(n8432) );
  AOI22_X1 U9974 ( .A1(n8430), .A2(n8437), .B1(n8436), .B2(n8429), .ZN(n8431)
         );
  NAND2_X1 U9975 ( .A1(n8432), .A2(n8431), .ZN(P2_U3435) );
  INV_X1 U9976 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8434) );
  MUX2_X1 U9977 ( .A(n8434), .B(n8433), .S(n9817), .Z(n8440) );
  AOI22_X1 U9978 ( .A1(n8438), .A2(n8437), .B1(n8436), .B2(n8435), .ZN(n8439)
         );
  NAND2_X1 U9979 ( .A1(n8440), .A2(n8439), .ZN(P2_U3432) );
  INV_X1 U9980 ( .A(n8617), .ZN(n9511) );
  NOR4_X1 U9981 ( .A1(n4540), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8441), .ZN(n8442) );
  AOI21_X1 U9982 ( .B1(n8446), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8442), .ZN(
        n8443) );
  OAI21_X1 U9983 ( .B1(n9511), .B2(n8451), .A(n8443), .ZN(P2_U3264) );
  INV_X1 U9984 ( .A(n8709), .ZN(n9518) );
  OAI222_X1 U9985 ( .A1(P2_U3151), .A2(n8444), .B1(n8451), .B2(n9518), .C1(
        n9982), .C2(n8449), .ZN(P2_U3266) );
  INV_X1 U9986 ( .A(n6101), .ZN(n9521) );
  AOI21_X1 U9987 ( .B1(n8446), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8445), .ZN(
        n8447) );
  OAI21_X1 U9988 ( .B1(n9521), .B2(n8451), .A(n8447), .ZN(P2_U3267) );
  INV_X1 U9989 ( .A(n8448), .ZN(n9524) );
  OAI222_X1 U9990 ( .A1(P2_U3151), .A2(n4398), .B1(n8451), .B2(n9524), .C1(
        n8450), .C2(n8449), .ZN(P2_U3268) );
  MUX2_X1 U9991 ( .A(n8452), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U9992 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8456) );
  NAND2_X1 U9993 ( .A1(n8456), .A2(n9571), .ZN(n8463) );
  INV_X1 U9994 ( .A(n8457), .ZN(n8459) );
  OAI22_X1 U9995 ( .A1(n8601), .A2(n8459), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8458), .ZN(n8460) );
  AOI21_X1 U9996 ( .B1(n8568), .B2(n8461), .A(n8460), .ZN(n8462) );
  OAI211_X1 U9997 ( .C1(n4627), .C2(n9568), .A(n8463), .B(n8462), .ZN(P1_U3215) );
  NAND2_X1 U9998 ( .A1(n8562), .A2(n8563), .ZN(n8561) );
  OAI21_X1 U9999 ( .B1(n8466), .B2(n8465), .A(n8561), .ZN(n8471) );
  OAI21_X1 U10000 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8470) );
  XNOR2_X1 U10001 ( .A(n8471), .B(n8470), .ZN(n8477) );
  OR2_X1 U10002 ( .A1(n9110), .A2(n9051), .ZN(n8473) );
  NAND2_X1 U10003 ( .A1(n9104), .A2(n9074), .ZN(n8472) );
  NAND2_X1 U10004 ( .A1(n8473), .A2(n8472), .ZN(n9209) );
  AOI22_X1 U10005 ( .A1(n9209), .A2(n9566), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8474) );
  OAI21_X1 U10006 ( .B1(n9575), .B2(n9214), .A(n8474), .ZN(n8475) );
  AOI21_X1 U10007 ( .B1(n9219), .B2(n8613), .A(n8475), .ZN(n8476) );
  OAI21_X1 U10008 ( .B1(n8477), .B2(n8615), .A(n8476), .ZN(P1_U3216) );
  AOI21_X1 U10009 ( .B1(n8479), .B2(n8481), .A(n8478), .ZN(n8480) );
  AOI21_X1 U10010 ( .B1(n4330), .B2(n8481), .A(n8480), .ZN(n8486) );
  NOR2_X1 U10011 ( .A1(n9575), .A2(n9280), .ZN(n8484) );
  AOI22_X1 U10012 ( .A1(n9096), .A2(n8588), .B1(n9074), .B2(n9088), .ZN(n9275)
         );
  INV_X1 U10013 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8482) );
  OAI22_X1 U10014 ( .A1(n9275), .A2(n8601), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8482), .ZN(n8483) );
  AOI211_X1 U10015 ( .C1(n9279), .C2(n8613), .A(n8484), .B(n8483), .ZN(n8485)
         );
  OAI21_X1 U10016 ( .B1(n8486), .B2(n8615), .A(n8485), .ZN(P1_U3219) );
  XOR2_X1 U10017 ( .A(n8488), .B(n8487), .Z(n8494) );
  NOR2_X1 U10018 ( .A1(n9575), .A2(n9248), .ZN(n8492) );
  AND2_X1 U10019 ( .A1(n9096), .A2(n9074), .ZN(n8489) );
  AOI21_X1 U10020 ( .B1(n9104), .B2(n8588), .A(n8489), .ZN(n9239) );
  OAI22_X1 U10021 ( .A1(n9239), .A2(n8601), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8490), .ZN(n8491) );
  AOI211_X1 U10022 ( .C1(n9246), .C2(n8613), .A(n8492), .B(n8491), .ZN(n8493)
         );
  OAI21_X1 U10023 ( .B1(n8494), .B2(n8615), .A(n8493), .ZN(P1_U3223) );
  XOR2_X1 U10024 ( .A(n8496), .B(n8495), .Z(n8504) );
  AOI21_X1 U10025 ( .B1(n9566), .B2(n8498), .A(n8497), .ZN(n8499) );
  OAI21_X1 U10026 ( .B1(n9575), .B2(n8500), .A(n8499), .ZN(n8501) );
  AOI21_X1 U10027 ( .B1(n8502), .B2(n8613), .A(n8501), .ZN(n8503) );
  OAI21_X1 U10028 ( .B1(n8504), .B2(n8615), .A(n8503), .ZN(P1_U3224) );
  OAI21_X1 U10029 ( .B1(n8507), .B2(n8506), .A(n8505), .ZN(n8514) );
  NAND2_X1 U10030 ( .A1(n9180), .A2(n8613), .ZN(n8512) );
  OR2_X1 U10031 ( .A1(n9110), .A2(n8508), .ZN(n8510) );
  NAND2_X1 U10032 ( .A1(n9116), .A2(n8588), .ZN(n8509) );
  NAND2_X1 U10033 ( .A1(n8510), .A2(n8509), .ZN(n9174) );
  AOI22_X1 U10034 ( .A1(n9174), .A2(n9566), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8511) );
  OAI211_X1 U10035 ( .C1(n9575), .C2(n9182), .A(n8512), .B(n8511), .ZN(n8513)
         );
  AOI21_X1 U10036 ( .B1(n8514), .B2(n9571), .A(n8513), .ZN(n8515) );
  INV_X1 U10037 ( .A(n8515), .ZN(P1_U3225) );
  XNOR2_X1 U10038 ( .A(n8516), .B(n8517), .ZN(n8608) );
  NOR2_X1 U10039 ( .A1(n8608), .A2(n8607), .ZN(n8606) );
  AOI21_X1 U10040 ( .B1(n8517), .B2(n8516), .A(n8606), .ZN(n8521) );
  XNOR2_X1 U10041 ( .A(n8519), .B(n8518), .ZN(n8520) );
  XNOR2_X1 U10042 ( .A(n8521), .B(n8520), .ZN(n8525) );
  NOR2_X1 U10043 ( .A1(n9575), .A2(n9346), .ZN(n8523) );
  AOI22_X1 U10044 ( .A1(n9083), .A2(n8588), .B1(n9074), .B2(n9077), .ZN(n9335)
         );
  NAND2_X1 U10045 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8996) );
  OAI21_X1 U10046 ( .B1(n8601), .B2(n9335), .A(n8996), .ZN(n8522) );
  AOI211_X1 U10047 ( .C1(n9344), .C2(n8613), .A(n8523), .B(n8522), .ZN(n8524)
         );
  OAI21_X1 U10048 ( .B1(n8525), .B2(n8615), .A(n8524), .ZN(P1_U3226) );
  XOR2_X1 U10049 ( .A(n8527), .B(n8526), .Z(n8531) );
  NOR2_X1 U10050 ( .A1(n9575), .A2(n9322), .ZN(n8529) );
  AOI22_X1 U10051 ( .A1(n9088), .A2(n8588), .B1(n9074), .B2(n9082), .ZN(n9314)
         );
  NAND2_X1 U10052 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9016) );
  OAI21_X1 U10053 ( .B1(n9314), .B2(n8601), .A(n9016), .ZN(n8528) );
  AOI211_X1 U10054 ( .C1(n9321), .C2(n8613), .A(n8529), .B(n8528), .ZN(n8530)
         );
  OAI21_X1 U10055 ( .B1(n8531), .B2(n8615), .A(n8530), .ZN(P1_U3228) );
  OAI21_X1 U10056 ( .B1(n8534), .B2(n8533), .A(n8532), .ZN(n8535) );
  NAND2_X1 U10057 ( .A1(n8535), .A2(n9571), .ZN(n8542) );
  NAND2_X1 U10058 ( .A1(n9113), .A2(n8588), .ZN(n8537) );
  NAND2_X1 U10059 ( .A1(n9107), .A2(n9074), .ZN(n8536) );
  NAND2_X1 U10060 ( .A1(n8537), .A2(n8536), .ZN(n9192) );
  OAI22_X1 U10061 ( .A1(n8539), .A2(n9575), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8538), .ZN(n8540) );
  AOI21_X1 U10062 ( .B1(n9192), .B2(n9566), .A(n8540), .ZN(n8541) );
  OAI211_X1 U10063 ( .C1(n9201), .C2(n9568), .A(n8542), .B(n8541), .ZN(
        P1_U3229) );
  OAI21_X1 U10064 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8546) );
  NAND2_X1 U10065 ( .A1(n8546), .A2(n9571), .ZN(n8551) );
  AND2_X1 U10066 ( .A1(n9091), .A2(n9074), .ZN(n8547) );
  AOI21_X1 U10067 ( .B1(n9099), .B2(n8588), .A(n8547), .ZN(n9259) );
  OAI22_X1 U10068 ( .A1(n9259), .A2(n8601), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8548), .ZN(n8549) );
  AOI21_X1 U10069 ( .B1(n9264), .B2(n8568), .A(n8549), .ZN(n8550) );
  OAI211_X1 U10070 ( .C1(n9483), .C2(n9568), .A(n8551), .B(n8550), .ZN(
        P1_U3233) );
  XOR2_X1 U10071 ( .A(n8553), .B(n8552), .Z(n8560) );
  AOI22_X1 U10072 ( .A1(n9566), .A2(n8554), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8555) );
  OAI21_X1 U10073 ( .B1(n9575), .B2(n8556), .A(n8555), .ZN(n8557) );
  AOI21_X1 U10074 ( .B1(n8558), .B2(n8613), .A(n8557), .ZN(n8559) );
  OAI21_X1 U10075 ( .B1(n8560), .B2(n8615), .A(n8559), .ZN(P1_U3234) );
  OAI21_X1 U10076 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8564) );
  NAND2_X1 U10077 ( .A1(n8564), .A2(n9571), .ZN(n8570) );
  INV_X1 U10078 ( .A(n8565), .ZN(n9232) );
  AOI22_X1 U10079 ( .A1(n9107), .A2(n8588), .B1(n9074), .B2(n9099), .ZN(n9228)
         );
  INV_X1 U10080 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8566) );
  OAI22_X1 U10081 ( .A1(n9228), .A2(n8601), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8566), .ZN(n8567) );
  AOI21_X1 U10082 ( .B1(n9232), .B2(n8568), .A(n8567), .ZN(n8569) );
  OAI211_X1 U10083 ( .C1(n9476), .C2(n9568), .A(n8570), .B(n8569), .ZN(
        P1_U3235) );
  INV_X1 U10084 ( .A(n8571), .ZN(n8576) );
  AOI21_X1 U10085 ( .B1(n8573), .B2(n8575), .A(n8572), .ZN(n8574) );
  AOI21_X1 U10086 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n8583) );
  AOI22_X1 U10087 ( .A1(n9566), .A2(n8577), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8578) );
  OAI21_X1 U10088 ( .B1(n9575), .B2(n8579), .A(n8578), .ZN(n8580) );
  AOI21_X1 U10089 ( .B1(n8581), .B2(n8613), .A(n8580), .ZN(n8582) );
  OAI21_X1 U10090 ( .B1(n8583), .B2(n8615), .A(n8582), .ZN(P1_U3236) );
  XNOR2_X1 U10091 ( .A(n8585), .B(n8584), .ZN(n8586) );
  XNOR2_X1 U10092 ( .A(n8587), .B(n8586), .ZN(n8594) );
  NAND2_X1 U10093 ( .A1(n9091), .A2(n8588), .ZN(n8590) );
  NAND2_X1 U10094 ( .A1(n9083), .A2(n9074), .ZN(n8589) );
  NAND2_X1 U10095 ( .A1(n8590), .A2(n8589), .ZN(n9296) );
  AOI22_X1 U10096 ( .A1(n9296), .A2(n9566), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8591) );
  OAI21_X1 U10097 ( .B1(n9575), .B2(n9301), .A(n8591), .ZN(n8592) );
  AOI21_X1 U10098 ( .B1(n9300), .B2(n8613), .A(n8592), .ZN(n8593) );
  OAI21_X1 U10099 ( .B1(n8594), .B2(n8615), .A(n8593), .ZN(P1_U3238) );
  INV_X1 U10100 ( .A(n8505), .ZN(n8597) );
  OAI21_X1 U10101 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8599) );
  NAND3_X1 U10102 ( .A1(n8599), .A2(n9571), .A3(n8598), .ZN(n8605) );
  NOR2_X1 U10103 ( .A1(n9575), .A2(n9165), .ZN(n8603) );
  NOR2_X1 U10104 ( .A1(n9118), .A2(n9051), .ZN(n8600) );
  AOI21_X1 U10105 ( .B1(n9113), .B2(n9074), .A(n8600), .ZN(n9158) );
  NOR2_X1 U10106 ( .A1(n9158), .A2(n8601), .ZN(n8602) );
  AOI211_X1 U10107 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n8603), 
        .B(n8602), .ZN(n8604) );
  OAI211_X1 U10108 ( .C1(n9464), .C2(n9568), .A(n8605), .B(n8604), .ZN(
        P1_U3240) );
  AOI21_X1 U10109 ( .B1(n8608), .B2(n8607), .A(n8606), .ZN(n8616) );
  AOI22_X1 U10110 ( .A1(n9566), .A2(n8609), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8610) );
  OAI21_X1 U10111 ( .B1(n9575), .B2(n8611), .A(n8610), .ZN(n8612) );
  AOI21_X1 U10112 ( .B1(n9078), .B2(n8613), .A(n8612), .ZN(n8614) );
  OAI21_X1 U10113 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(P1_U3241) );
  NAND2_X1 U10114 ( .A1(n8617), .A2(n8716), .ZN(n8620) );
  OR2_X1 U10115 ( .A1(n8717), .A2(n8618), .ZN(n8619) );
  INV_X1 U10116 ( .A(n9052), .ZN(n8756) );
  AND2_X1 U10117 ( .A1(n8728), .A2(n8756), .ZN(n8798) );
  INV_X1 U10118 ( .A(n8722), .ZN(n8727) );
  INV_X1 U10119 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9057) );
  INV_X1 U10120 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9360) );
  OR2_X1 U10121 ( .A1(n4271), .A2(n9360), .ZN(n8623) );
  INV_X1 U10122 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9452) );
  OR2_X1 U10123 ( .A1(n4420), .A2(n9452), .ZN(n8622) );
  OAI211_X1 U10124 ( .C1(n8624), .C2(n9057), .A(n8623), .B(n8622), .ZN(n9073)
         );
  OAI21_X1 U10125 ( .B1(n9451), .B2(n9073), .A(n9052), .ZN(n8726) );
  NAND2_X1 U10126 ( .A1(n8760), .A2(n8761), .ZN(n8708) );
  OR2_X1 U10127 ( .A1(n9263), .A2(n9098), .ZN(n9062) );
  INV_X1 U10128 ( .A(n9091), .ZN(n9093) );
  OR2_X1 U10129 ( .A1(n9279), .A2(n9093), .ZN(n8750) );
  AND2_X1 U10130 ( .A1(n9062), .A2(n8750), .ZN(n8686) );
  NAND2_X1 U10131 ( .A1(n9344), .A2(n8625), .ZN(n8843) );
  AND2_X1 U10132 ( .A1(n8843), .A2(n9329), .ZN(n8746) );
  INV_X1 U10133 ( .A(n8767), .ZN(n8626) );
  OAI22_X1 U10134 ( .A1(n8746), .A2(n8626), .B1(n8722), .B2(n9078), .ZN(n8677)
         );
  INV_X1 U10135 ( .A(n8843), .ZN(n8627) );
  OAI21_X1 U10136 ( .B1(n8627), .B2(n9081), .A(n8727), .ZN(n8676) );
  INV_X1 U10137 ( .A(n8628), .ZN(n8633) );
  INV_X1 U10138 ( .A(n8632), .ZN(n8635) );
  AOI21_X1 U10139 ( .B1(n8635), .B2(n8634), .A(n8633), .ZN(n8636) );
  MUX2_X1 U10140 ( .A(n8637), .B(n8636), .S(n8722), .Z(n8643) );
  INV_X1 U10141 ( .A(n8638), .ZN(n8639) );
  MUX2_X1 U10142 ( .A(n8640), .B(n8639), .S(n8722), .Z(n8641) );
  OAI21_X1 U10143 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8648) );
  AND2_X1 U10144 ( .A1(n8655), .A2(n8644), .ZN(n8646) );
  MUX2_X1 U10145 ( .A(n8646), .B(n8645), .S(n8722), .Z(n8647) );
  INV_X1 U10146 ( .A(n8657), .ZN(n8650) );
  NAND2_X1 U10147 ( .A1(n8826), .A2(n8654), .ZN(n8649) );
  OAI21_X1 U10148 ( .B1(n8650), .B2(n8649), .A(n8658), .ZN(n8653) );
  NAND2_X1 U10149 ( .A1(n8833), .A2(n8659), .ZN(n8651) );
  AOI22_X1 U10150 ( .A1(n8653), .A2(n8830), .B1(n8652), .B2(n8651), .ZN(n8664)
         );
  INV_X1 U10151 ( .A(n8654), .ZN(n8656) );
  NAND2_X1 U10152 ( .A1(n8659), .A2(n8658), .ZN(n8829) );
  INV_X1 U10153 ( .A(n8830), .ZN(n8661) );
  OAI21_X1 U10154 ( .B1(n8662), .B2(n8661), .A(n8833), .ZN(n8663) );
  MUX2_X1 U10155 ( .A(n8664), .B(n8663), .S(n8722), .Z(n8669) );
  NAND2_X1 U10156 ( .A1(n8670), .A2(n8668), .ZN(n8837) );
  AOI21_X1 U10157 ( .B1(n8669), .B2(n8832), .A(n8837), .ZN(n8666) );
  NAND2_X1 U10158 ( .A1(n8746), .A2(n8835), .ZN(n8665) );
  OAI21_X1 U10159 ( .B1(n8666), .B2(n8665), .A(n8767), .ZN(n8675) );
  INV_X1 U10160 ( .A(n8835), .ZN(n8667) );
  INV_X1 U10161 ( .A(n8670), .ZN(n8672) );
  NAND2_X1 U10162 ( .A1(n8767), .A2(n8671), .ZN(n8811) );
  NOR3_X1 U10163 ( .A1(n8673), .A2(n8672), .A3(n8811), .ZN(n8674) );
  XNOR2_X1 U10164 ( .A(n9321), .B(n9083), .ZN(n9312) );
  INV_X1 U10165 ( .A(n9312), .ZN(n9316) );
  INV_X1 U10166 ( .A(n9088), .ZN(n9089) );
  OR2_X1 U10167 ( .A1(n9300), .A2(n9089), .ZN(n8748) );
  INV_X1 U10168 ( .A(n9083), .ZN(n9085) );
  OR2_X1 U10169 ( .A1(n9321), .A2(n9085), .ZN(n9289) );
  NAND3_X1 U10170 ( .A1(n8678), .A2(n8748), .A3(n9289), .ZN(n8679) );
  NAND2_X1 U10171 ( .A1(n9279), .A2(n9093), .ZN(n8751) );
  NAND2_X1 U10172 ( .A1(n9300), .A2(n9089), .ZN(n8749) );
  NAND3_X1 U10173 ( .A1(n8679), .A2(n8751), .A3(n8749), .ZN(n8685) );
  NAND2_X1 U10174 ( .A1(n8750), .A2(n8748), .ZN(n8840) );
  INV_X1 U10175 ( .A(n8840), .ZN(n8682) );
  AND2_X1 U10176 ( .A1(n9263), .A2(n9098), .ZN(n8765) );
  INV_X1 U10177 ( .A(n8749), .ZN(n8680) );
  AOI21_X1 U10178 ( .B1(n9085), .B2(n9321), .A(n8680), .ZN(n8681) );
  OAI21_X1 U10179 ( .B1(n8681), .B2(n8840), .A(n8751), .ZN(n8846) );
  AOI211_X1 U10180 ( .C1(n8683), .C2(n8682), .A(n8765), .B(n8846), .ZN(n8684)
         );
  NAND2_X1 U10181 ( .A1(n8689), .A2(n8765), .ZN(n8688) );
  NAND2_X1 U10182 ( .A1(n9246), .A2(n9100), .ZN(n8687) );
  AND2_X1 U10183 ( .A1(n8688), .A2(n8687), .ZN(n9063) );
  AND2_X1 U10184 ( .A1(n8689), .A2(n9062), .ZN(n8742) );
  INV_X1 U10185 ( .A(n9104), .ZN(n9106) );
  NAND2_X1 U10186 ( .A1(n9231), .A2(n9106), .ZN(n8691) );
  NAND2_X1 U10187 ( .A1(n9204), .A2(n8691), .ZN(n9224) );
  INV_X1 U10188 ( .A(n9107), .ZN(n9108) );
  NAND2_X1 U10189 ( .A1(n9219), .A2(n9108), .ZN(n9190) );
  AND2_X1 U10190 ( .A1(n9190), .A2(n8691), .ZN(n8733) );
  OR2_X1 U10191 ( .A1(n9219), .A2(n9108), .ZN(n8764) );
  NAND2_X1 U10192 ( .A1(n8764), .A2(n9204), .ZN(n8729) );
  AOI22_X1 U10193 ( .A1(n8692), .A2(n8764), .B1(n8727), .B2(n8729), .ZN(n8695)
         );
  NAND2_X1 U10194 ( .A1(n9394), .A2(n9110), .ZN(n8734) );
  OAI21_X1 U10195 ( .B1(n8722), .B2(n9190), .A(n9189), .ZN(n8694) );
  MUX2_X1 U10196 ( .A(n9065), .B(n8734), .S(n8722), .Z(n8693) );
  INV_X1 U10197 ( .A(n9155), .ZN(n8696) );
  NOR2_X1 U10198 ( .A1(n8700), .A2(n8696), .ZN(n8698) );
  INV_X1 U10199 ( .A(n9116), .ZN(n8697) );
  NAND2_X1 U10200 ( .A1(n9164), .A2(n8697), .ZN(n9066) );
  NAND2_X1 U10201 ( .A1(n9180), .A2(n9114), .ZN(n8763) );
  NAND2_X1 U10202 ( .A1(n9066), .A2(n8763), .ZN(n8735) );
  OR2_X1 U10203 ( .A1(n9164), .A2(n8697), .ZN(n8762) );
  INV_X1 U10204 ( .A(n8763), .ZN(n8699) );
  OAI211_X1 U10205 ( .C1(n8700), .C2(n8699), .A(n8762), .B(n9155), .ZN(n8701)
         );
  NAND2_X1 U10206 ( .A1(n9373), .A2(n9119), .ZN(n9070) );
  NAND2_X1 U10207 ( .A1(n9379), .A2(n9118), .ZN(n9068) );
  NAND2_X1 U10208 ( .A1(n9070), .A2(n9068), .ZN(n8738) );
  INV_X1 U10209 ( .A(n8738), .ZN(n8707) );
  INV_X1 U10210 ( .A(n8760), .ZN(n8706) );
  INV_X1 U10211 ( .A(n9068), .ZN(n8702) );
  NAND2_X1 U10212 ( .A1(n8709), .A2(n8716), .ZN(n8711) );
  OR2_X1 U10213 ( .A1(n8717), .A2(n9956), .ZN(n8710) );
  INV_X1 U10214 ( .A(n8868), .ZN(n8712) );
  OR2_X1 U10215 ( .A1(n9046), .A2(n8712), .ZN(n8752) );
  NAND2_X1 U10216 ( .A1(n9046), .A2(n8712), .ZN(n8754) );
  OAI21_X1 U10217 ( .B1(n8727), .B2(n9070), .A(n9120), .ZN(n8714) );
  MUX2_X1 U10218 ( .A(n8754), .B(n8752), .S(n8722), .Z(n8713) );
  OAI21_X1 U10219 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8721) );
  NAND2_X1 U10220 ( .A1(n7718), .A2(n8716), .ZN(n8719) );
  OR2_X1 U10221 ( .A1(n8717), .A2(n9515), .ZN(n8718) );
  MUX2_X1 U10222 ( .A(n8721), .B(n8727), .S(n9060), .Z(n8725) );
  OAI211_X1 U10223 ( .C1(n8855), .C2(n8810), .A(n5719), .B(n8803), .ZN(n8808)
         );
  NAND2_X1 U10224 ( .A1(n8729), .A2(n9190), .ZN(n8730) );
  NAND2_X1 U10225 ( .A1(n9065), .A2(n8730), .ZN(n8731) );
  NAND2_X1 U10226 ( .A1(n8731), .A2(n8734), .ZN(n8732) );
  AND2_X1 U10227 ( .A1(n9155), .A2(n8732), .ZN(n8741) );
  NAND3_X1 U10228 ( .A1(n8734), .A2(n8733), .A3(n9063), .ZN(n8736) );
  AOI21_X1 U10229 ( .B1(n8741), .B2(n8736), .A(n8735), .ZN(n8737) );
  NAND2_X1 U10230 ( .A1(n8761), .A2(n8762), .ZN(n8740) );
  NOR2_X1 U10231 ( .A1(n8737), .A2(n8740), .ZN(n8739) );
  NOR2_X1 U10232 ( .A1(n8739), .A2(n8738), .ZN(n8850) );
  INV_X1 U10233 ( .A(n8740), .ZN(n8845) );
  INV_X1 U10234 ( .A(n8741), .ZN(n8744) );
  INV_X1 U10235 ( .A(n8742), .ZN(n8743) );
  NOR2_X1 U10236 ( .A1(n8744), .A2(n8743), .ZN(n8844) );
  NAND2_X1 U10237 ( .A1(n9330), .A2(n8746), .ZN(n8747) );
  NAND3_X1 U10238 ( .A1(n8845), .A2(n8844), .A3(n9255), .ZN(n8753) );
  NAND2_X1 U10239 ( .A1(n8752), .A2(n8760), .ZN(n8848) );
  AOI21_X1 U10240 ( .B1(n8850), .B2(n8753), .A(n8848), .ZN(n8757) );
  INV_X1 U10241 ( .A(n9073), .ZN(n8755) );
  NAND2_X1 U10242 ( .A1(n9060), .A2(n8755), .ZN(n8796) );
  NAND2_X1 U10243 ( .A1(n8796), .A2(n8754), .ZN(n8853) );
  OR2_X1 U10244 ( .A1(n9060), .A2(n8755), .ZN(n8851) );
  OAI22_X1 U10245 ( .A1(n8757), .A2(n8853), .B1(n8756), .B2(n8851), .ZN(n8758)
         );
  OAI211_X1 U10246 ( .C1(n8720), .C2(n9052), .A(n8758), .B(n8855), .ZN(n8802)
         );
  NOR2_X1 U10247 ( .A1(n8798), .A2(n8759), .ZN(n8801) );
  NAND2_X1 U10248 ( .A1(n8760), .A2(n9070), .ZN(n9134) );
  NAND2_X1 U10249 ( .A1(n8761), .A2(n9068), .ZN(n9144) );
  INV_X1 U10250 ( .A(n9224), .ZN(n9222) );
  INV_X1 U10251 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U10252 ( .A1(n9062), .A2(n8766), .ZN(n9256) );
  NAND2_X1 U10253 ( .A1(n8767), .A2(n8843), .ZN(n9337) );
  NAND4_X1 U10254 ( .A1(n8770), .A2(n8771), .A3(n9667), .A4(n8769), .ZN(n8773)
         );
  NOR2_X1 U10255 ( .A1(n8773), .A2(n8772), .ZN(n8779) );
  INV_X1 U10256 ( .A(n8774), .ZN(n8777) );
  INV_X1 U10257 ( .A(n8775), .ZN(n8776) );
  NAND4_X1 U10258 ( .A1(n8779), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n8780)
         );
  NOR2_X1 U10259 ( .A1(n8781), .A2(n8780), .ZN(n8782) );
  NAND3_X1 U10260 ( .A1(n4787), .A2(n4323), .A3(n8782), .ZN(n8783) );
  OR2_X1 U10261 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  NOR2_X1 U10262 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  NAND4_X1 U10263 ( .A1(n8789), .A2(n4644), .A3(n8788), .A4(n8787), .ZN(n8790)
         );
  NOR2_X1 U10264 ( .A1(n9337), .A2(n8790), .ZN(n8791) );
  NAND4_X1 U10265 ( .A1(n9272), .A2(n9290), .A3(n8791), .A4(n9312), .ZN(n8792)
         );
  NOR2_X1 U10266 ( .A1(n9256), .A2(n8792), .ZN(n8793) );
  XNOR2_X1 U10267 ( .A(n9246), .B(n9100), .ZN(n9064) );
  INV_X1 U10268 ( .A(n9064), .ZN(n9242) );
  AND4_X1 U10269 ( .A1(n9212), .A2(n9222), .A3(n8793), .A4(n9242), .ZN(n8794)
         );
  NAND4_X1 U10270 ( .A1(n9160), .A2(n9189), .A3(n9178), .A4(n8794), .ZN(n8795)
         );
  NOR3_X1 U10271 ( .A1(n9134), .A2(n9144), .A3(n8795), .ZN(n8797) );
  AND4_X1 U10272 ( .A1(n9120), .A2(n8851), .A3(n8797), .A4(n8796), .ZN(n8799)
         );
  INV_X1 U10273 ( .A(n8798), .ZN(n8852) );
  NAND3_X1 U10274 ( .A1(n8855), .A2(n8799), .A3(n8852), .ZN(n8805) );
  INV_X1 U10275 ( .A(n8805), .ZN(n8800) );
  AOI21_X1 U10276 ( .B1(n8802), .B2(n8801), .A(n8800), .ZN(n8807) );
  OAI21_X1 U10277 ( .B1(n8804), .B2(n8803), .A(n5719), .ZN(n8806) );
  NOR2_X1 U10278 ( .A1(n8810), .A2(n8860), .ZN(n9671) );
  INV_X1 U10279 ( .A(n8811), .ZN(n8839) );
  INV_X1 U10280 ( .A(n8812), .ZN(n8825) );
  INV_X1 U10281 ( .A(n8813), .ZN(n8818) );
  NAND2_X1 U10282 ( .A1(n4391), .A2(n8814), .ZN(n8816) );
  AND4_X1 U10283 ( .A1(n8818), .A2(n8817), .A3(n5719), .A4(n8816), .ZN(n8823)
         );
  NAND2_X1 U10284 ( .A1(n8879), .A2(n8819), .ZN(n8820) );
  NAND4_X1 U10285 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n8824)
         );
  NAND2_X1 U10286 ( .A1(n8825), .A2(n8824), .ZN(n8827) );
  NAND4_X1 U10287 ( .A1(n8830), .A2(n8828), .A3(n8827), .A4(n8826), .ZN(n8834)
         );
  NAND2_X1 U10288 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  AND4_X1 U10289 ( .A1(n8834), .A2(n8833), .A3(n8832), .A4(n8831), .ZN(n8836)
         );
  OAI211_X1 U10290 ( .C1(n8837), .C2(n8836), .A(n9329), .B(n8835), .ZN(n8838)
         );
  NAND2_X1 U10291 ( .A1(n8839), .A2(n8838), .ZN(n8842) );
  INV_X1 U10292 ( .A(n9289), .ZN(n8841) );
  AOI211_X1 U10293 ( .C1(n8843), .C2(n8842), .A(n8841), .B(n8840), .ZN(n8847)
         );
  OAI211_X1 U10294 ( .C1(n8847), .C2(n8846), .A(n8845), .B(n8844), .ZN(n8849)
         );
  AOI21_X1 U10295 ( .B1(n8850), .B2(n8849), .A(n8848), .ZN(n8854) );
  OAI211_X1 U10296 ( .C1(n8854), .C2(n8853), .A(n8852), .B(n8851), .ZN(n8856)
         );
  NAND2_X1 U10297 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  MUX2_X1 U10298 ( .A(n9671), .B(n8858), .S(n8857), .Z(n8859) );
  NOR2_X1 U10299 ( .A1(n8862), .A2(n8861), .ZN(n8865) );
  OAI21_X1 U10300 ( .B1(n8866), .B2(n8863), .A(P1_B_REG_SCAN_IN), .ZN(n8864)
         );
  OAI22_X1 U10301 ( .A1(n8867), .A2(n8866), .B1(n8865), .B2(n8864), .ZN(
        P1_U3242) );
  MUX2_X1 U10302 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9073), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10303 ( .A(n8868), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8869), .Z(
        P1_U3583) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9075), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9116), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9113), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9111), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9107), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9104), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9099), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9096), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9091), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9088), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9083), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10315 ( .A(n9082), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8869), .Z(
        P1_U3570) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9077), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8870), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8871), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10319 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8872), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8873), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10321 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8874), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n4646), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n4649), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10324 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8875), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8876), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8877), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8878), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8879), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8880), .S(P1_U3973), .Z(
        P1_U3556) );
  INV_X1 U10330 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8881) );
  OAI22_X1 U10331 ( .A1(n9650), .A2(n8881), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4397), .ZN(n8882) );
  AOI21_X1 U10332 ( .B1(n8883), .B2(n9630), .A(n8882), .ZN(n8892) );
  AND2_X1 U10333 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8885) );
  OAI211_X1 U10334 ( .C1(n8886), .C2(n8885), .A(n9634), .B(n8884), .ZN(n8891)
         );
  OAI211_X1 U10335 ( .C1(n8889), .C2(n8888), .A(n9642), .B(n8887), .ZN(n8890)
         );
  NAND3_X1 U10336 ( .A1(n8892), .A2(n8891), .A3(n8890), .ZN(P1_U3244) );
  INV_X1 U10337 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8893) );
  OAI22_X1 U10338 ( .A1(n9650), .A2(n8893), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9653), .ZN(n8894) );
  AOI21_X1 U10339 ( .B1(n8895), .B2(n9630), .A(n8894), .ZN(n8904) );
  OAI211_X1 U10340 ( .C1(n8898), .C2(n8897), .A(n9642), .B(n8896), .ZN(n8903)
         );
  OAI211_X1 U10341 ( .C1(n8901), .C2(n8900), .A(n9634), .B(n8899), .ZN(n8902)
         );
  NAND4_X1 U10342 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(
        P1_U3245) );
  AOI211_X1 U10343 ( .C1(n4321), .C2(n8907), .A(n8906), .B(n9619), .ZN(n8908)
         );
  INV_X1 U10344 ( .A(n8908), .ZN(n8918) );
  INV_X1 U10345 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U10346 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n8909) );
  OAI21_X1 U10347 ( .B1(n9650), .B2(n8910), .A(n8909), .ZN(n8911) );
  AOI21_X1 U10348 ( .B1(n8912), .B2(n9630), .A(n8911), .ZN(n8917) );
  OAI211_X1 U10349 ( .C1(n8915), .C2(n8914), .A(n9642), .B(n8913), .ZN(n8916)
         );
  NAND3_X1 U10350 ( .A1(n8918), .A2(n8917), .A3(n8916), .ZN(P1_U3246) );
  AOI211_X1 U10351 ( .C1(n8921), .C2(n8920), .A(n9619), .B(n8919), .ZN(n8922)
         );
  INV_X1 U10352 ( .A(n8922), .ZN(n8932) );
  INV_X1 U10353 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n8924) );
  OAI21_X1 U10354 ( .B1(n9650), .B2(n8924), .A(n8923), .ZN(n8925) );
  AOI21_X1 U10355 ( .B1(n8926), .B2(n9630), .A(n8925), .ZN(n8931) );
  OAI211_X1 U10356 ( .C1(n8929), .C2(n8928), .A(n9642), .B(n8927), .ZN(n8930)
         );
  NAND3_X1 U10357 ( .A1(n8932), .A2(n8931), .A3(n8930), .ZN(P1_U3248) );
  AOI211_X1 U10358 ( .C1(n8935), .C2(n8934), .A(n9619), .B(n8933), .ZN(n8936)
         );
  INV_X1 U10359 ( .A(n8936), .ZN(n8946) );
  INV_X1 U10360 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8938) );
  OAI21_X1 U10361 ( .B1(n9650), .B2(n8938), .A(n8937), .ZN(n8939) );
  AOI21_X1 U10362 ( .B1(n8940), .B2(n9630), .A(n8939), .ZN(n8945) );
  OAI211_X1 U10363 ( .C1(n8943), .C2(n8942), .A(n9642), .B(n8941), .ZN(n8944)
         );
  NAND3_X1 U10364 ( .A1(n8946), .A2(n8945), .A3(n8944), .ZN(P1_U3249) );
  AOI211_X1 U10365 ( .C1(n8949), .C2(n8948), .A(n9619), .B(n8947), .ZN(n8950)
         );
  INV_X1 U10366 ( .A(n8950), .ZN(n8960) );
  INV_X1 U10367 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8952) );
  OAI21_X1 U10368 ( .B1(n9650), .B2(n8952), .A(n8951), .ZN(n8953) );
  AOI21_X1 U10369 ( .B1(n8954), .B2(n9630), .A(n8953), .ZN(n8959) );
  OAI211_X1 U10370 ( .C1(n8957), .C2(n8956), .A(n9642), .B(n8955), .ZN(n8958)
         );
  NAND3_X1 U10371 ( .A1(n8960), .A2(n8959), .A3(n8958), .ZN(P1_U3250) );
  AOI211_X1 U10372 ( .C1(n8963), .C2(n8962), .A(n9619), .B(n8961), .ZN(n8964)
         );
  INV_X1 U10373 ( .A(n8964), .ZN(n8974) );
  INV_X1 U10374 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8966) );
  OAI21_X1 U10375 ( .B1(n9650), .B2(n8966), .A(n8965), .ZN(n8967) );
  AOI21_X1 U10376 ( .B1(n8968), .B2(n9630), .A(n8967), .ZN(n8973) );
  OAI211_X1 U10377 ( .C1(n8971), .C2(n8970), .A(n9642), .B(n8969), .ZN(n8972)
         );
  NAND3_X1 U10378 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(P1_U3251) );
  OAI21_X1 U10379 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n8978) );
  NAND2_X1 U10380 ( .A1(n8978), .A2(n9634), .ZN(n8988) );
  AOI21_X1 U10381 ( .B1(n9014), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8979), .ZN(
        n8987) );
  OAI21_X1 U10382 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8983) );
  NAND2_X1 U10383 ( .A1(n8983), .A2(n9642), .ZN(n8986) );
  NAND2_X1 U10384 ( .A1(n9630), .A2(n8984), .ZN(n8985) );
  NAND4_X1 U10385 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(
        P1_U3252) );
  AOI22_X1 U10386 ( .A1(n9013), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9999), .B2(
        n9004), .ZN(n8994) );
  XNOR2_X1 U10387 ( .A(n9593), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9591) );
  OR2_X1 U10388 ( .A1(n8999), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8990) );
  XNOR2_X1 U10389 ( .A(n9608), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U10390 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  NOR2_X1 U10391 ( .A1(n8991), .A2(n9002), .ZN(n8992) );
  NOR2_X1 U10392 ( .A1(n9621), .A2(n9622), .ZN(n9620) );
  OAI21_X1 U10393 ( .B1(n8994), .B2(n8993), .A(n9011), .ZN(n9009) );
  NAND2_X1 U10394 ( .A1(n9014), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8995) );
  OAI211_X1 U10395 ( .C1(n9646), .C2(n9004), .A(n8996), .B(n8995), .ZN(n9008)
         );
  AOI22_X1 U10396 ( .A1(n9593), .A2(n5317), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n8997), .ZN(n9595) );
  OAI21_X1 U10397 ( .B1(n8999), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8998), .ZN(
        n9596) );
  NOR2_X1 U10398 ( .A1(n9595), .A2(n9596), .ZN(n9594) );
  AOI21_X1 U10399 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9593), .A(n9594), .ZN(
        n9610) );
  AOI22_X1 U10400 ( .A1(n9608), .A2(n5348), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n9000), .ZN(n9611) );
  NOR2_X1 U10401 ( .A1(n9610), .A2(n9611), .ZN(n9609) );
  AOI21_X1 U10402 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9608), .A(n9609), .ZN(
        n9001) );
  NOR2_X1 U10403 ( .A1(n9001), .A2(n9002), .ZN(n9003) );
  XNOR2_X1 U10404 ( .A(n9002), .B(n9001), .ZN(n9626) );
  NOR2_X1 U10405 ( .A1(n9625), .A2(n9626), .ZN(n9624) );
  NOR2_X1 U10406 ( .A1(n9003), .A2(n9624), .ZN(n9006) );
  AOI22_X1 U10407 ( .A1(n9013), .A2(n9347), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9004), .ZN(n9005) );
  NOR2_X1 U10408 ( .A1(n9006), .A2(n9005), .ZN(n9012) );
  INV_X1 U10409 ( .A(n9642), .ZN(n9623) );
  AOI211_X1 U10410 ( .C1(n9006), .C2(n9005), .A(n9012), .B(n9623), .ZN(n9007)
         );
  AOI211_X1 U10411 ( .C1(n9634), .C2(n9009), .A(n9008), .B(n9007), .ZN(n9010)
         );
  INV_X1 U10412 ( .A(n9010), .ZN(P1_U3259) );
  INV_X1 U10413 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9430) );
  XNOR2_X1 U10414 ( .A(n9031), .B(n9430), .ZN(n9023) );
  XOR2_X1 U10415 ( .A(n9023), .B(n9024), .Z(n9021) );
  INV_X1 U10416 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9323) );
  XNOR2_X1 U10417 ( .A(n9031), .B(n9323), .ZN(n9030) );
  AOI21_X1 U10418 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9013), .A(n9012), .ZN(
        n9029) );
  XNOR2_X1 U10419 ( .A(n9030), .B(n9029), .ZN(n9019) );
  NAND2_X1 U10420 ( .A1(n9014), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9015) );
  OAI211_X1 U10421 ( .C1(n9646), .C2(n9017), .A(n9016), .B(n9015), .ZN(n9018)
         );
  AOI21_X1 U10422 ( .B1(n9642), .B2(n9019), .A(n9018), .ZN(n9020) );
  OAI21_X1 U10423 ( .B1(n9021), .B2(n9619), .A(n9020), .ZN(P1_U3260) );
  NOR2_X1 U10424 ( .A1(n9031), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9022) );
  AOI21_X1 U10425 ( .B1(n9024), .B2(n9023), .A(n9022), .ZN(n9637) );
  NAND2_X1 U10426 ( .A1(n9028), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9026) );
  OAI21_X1 U10427 ( .B1(n9028), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9026), .ZN(
        n9025) );
  INV_X1 U10428 ( .A(n9025), .ZN(n9636) );
  NAND2_X1 U10429 ( .A1(n9637), .A2(n9636), .ZN(n9635) );
  NAND2_X1 U10430 ( .A1(n9635), .A2(n9026), .ZN(n9027) );
  INV_X1 U10431 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9420) );
  XNOR2_X1 U10432 ( .A(n9027), .B(n9420), .ZN(n9037) );
  NAND2_X1 U10433 ( .A1(n9028), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9034) );
  OAI21_X1 U10434 ( .B1(n9028), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9034), .ZN(
        n9638) );
  NAND2_X1 U10435 ( .A1(n9030), .A2(n9029), .ZN(n9033) );
  OR2_X1 U10436 ( .A1(n9031), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U10437 ( .A1(n9033), .A2(n9032), .ZN(n9639) );
  NAND2_X1 U10438 ( .A1(n9641), .A2(n9034), .ZN(n9035) );
  XNOR2_X1 U10439 ( .A(n9035), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9039) );
  INV_X1 U10440 ( .A(n9039), .ZN(n9036) );
  AOI22_X1 U10441 ( .A1(n9037), .A2(n9634), .B1(n9642), .B2(n9036), .ZN(n9042)
         );
  NOR2_X1 U10442 ( .A1(n9037), .A2(n9619), .ZN(n9038) );
  AOI211_X1 U10443 ( .C1(n9642), .C2(n9039), .A(n9630), .B(n9038), .ZN(n9041)
         );
  MUX2_X1 U10444 ( .A(n9042), .B(n9041), .S(n9040), .Z(n9044) );
  NAND2_X1 U10445 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9043) );
  OAI211_X1 U10446 ( .C1(n9045), .C2(n9650), .A(n9044), .B(n9043), .ZN(
        P1_U3262) );
  NOR2_X1 U10447 ( .A1(n9048), .A2(n9342), .ZN(n9355) );
  NAND2_X1 U10448 ( .A1(n9355), .A2(n9350), .ZN(n9054) );
  INV_X1 U10449 ( .A(n9523), .ZN(n9049) );
  AND2_X1 U10450 ( .A1(n9049), .A2(P1_B_REG_SCAN_IN), .ZN(n9050) );
  NOR2_X1 U10451 ( .A1(n9051), .A2(n9050), .ZN(n9072) );
  AND2_X1 U10452 ( .A1(n9052), .A2(n9072), .ZN(n9354) );
  INV_X1 U10453 ( .A(n9354), .ZN(n9358) );
  NOR2_X1 U10454 ( .A1(n9304), .A2(n9358), .ZN(n9058) );
  AOI21_X1 U10455 ( .B1(n9304), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9058), .ZN(
        n9053) );
  OAI211_X1 U10456 ( .C1(n9451), .C2(n9345), .A(n9054), .B(n9053), .ZN(
        P1_U3263) );
  NAND2_X1 U10457 ( .A1(n9060), .A2(n9123), .ZN(n9055) );
  NAND2_X1 U10458 ( .A1(n9055), .A2(n9216), .ZN(n9056) );
  OR2_X1 U10459 ( .A1(n4348), .A2(n9056), .ZN(n9359) );
  NOR2_X1 U10460 ( .A1(n9678), .A2(n9057), .ZN(n9059) );
  AOI211_X1 U10461 ( .C1(n9060), .C2(n9657), .A(n9059), .B(n9058), .ZN(n9061)
         );
  OAI21_X1 U10462 ( .B1(n9359), .B2(n9660), .A(n9061), .ZN(P1_U3264) );
  INV_X1 U10463 ( .A(n9120), .ZN(n9071) );
  NAND2_X1 U10464 ( .A1(n9173), .A2(n9178), .ZN(n9172) );
  NAND3_X1 U10465 ( .A1(n9172), .A2(n9160), .A3(n9155), .ZN(n9067) );
  NAND2_X1 U10466 ( .A1(n9067), .A2(n9066), .ZN(n9145) );
  INV_X1 U10467 ( .A(n9144), .ZN(n9142) );
  NAND2_X1 U10468 ( .A1(n9145), .A2(n9142), .ZN(n9069) );
  NAND2_X1 U10469 ( .A1(n9069), .A2(n9068), .ZN(n9130) );
  INV_X1 U10470 ( .A(n9134), .ZN(n9131) );
  AOI22_X1 U10471 ( .A1(n9075), .A2(n9074), .B1(n9073), .B2(n9072), .ZN(n9076)
         );
  NAND2_X1 U10472 ( .A1(n9321), .A2(n9083), .ZN(n9084) );
  NAND2_X1 U10473 ( .A1(n9087), .A2(n9086), .ZN(n9287) );
  NAND2_X1 U10474 ( .A1(n9101), .A2(n9100), .ZN(n9102) );
  NAND2_X1 U10475 ( .A1(n9103), .A2(n4927), .ZN(n9223) );
  NOR2_X1 U10476 ( .A1(n9201), .A2(n9110), .ZN(n9112) );
  NOR2_X1 U10477 ( .A1(n9180), .A2(n9113), .ZN(n9115) );
  AND2_X1 U10478 ( .A1(n9164), .A2(n9116), .ZN(n9117) );
  NAND2_X1 U10479 ( .A1(n9365), .A2(n9339), .ZN(n9128) );
  OAI22_X1 U10480 ( .A1(n9678), .A2(n9122), .B1(n9121), .B2(n9673), .ZN(n9126)
         );
  INV_X1 U10481 ( .A(n9046), .ZN(n9124) );
  OAI211_X1 U10482 ( .C1(n9124), .C2(n4307), .A(n9216), .B(n9123), .ZN(n9362)
         );
  NOR2_X1 U10483 ( .A1(n9362), .A2(n9660), .ZN(n9125) );
  AOI211_X1 U10484 ( .C1(n9657), .C2(n9046), .A(n9126), .B(n9125), .ZN(n9127)
         );
  OAI211_X1 U10485 ( .C1(n9363), .C2(n9304), .A(n9128), .B(n9127), .ZN(
        P1_U3356) );
  OAI21_X1 U10486 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9133) );
  AOI21_X1 U10487 ( .B1(n9133), .B2(n9333), .A(n9132), .ZN(n9375) );
  OR2_X1 U10488 ( .A1(n9135), .A2(n9134), .ZN(n9371) );
  NAND3_X1 U10489 ( .A1(n9371), .A2(n9370), .A3(n9339), .ZN(n9141) );
  AOI211_X1 U10490 ( .C1(n9373), .C2(n9148), .A(n9342), .B(n4307), .ZN(n9372)
         );
  AOI22_X1 U10491 ( .A1(n9304), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9137), .B2(
        n9302), .ZN(n9138) );
  OAI21_X1 U10492 ( .B1(n9047), .B2(n9345), .A(n9138), .ZN(n9139) );
  AOI21_X1 U10493 ( .B1(n9372), .B2(n9350), .A(n9139), .ZN(n9140) );
  OAI211_X1 U10494 ( .C1(n9304), .C2(n9375), .A(n9141), .B(n9140), .ZN(
        P1_U3265) );
  XNOR2_X1 U10495 ( .A(n9143), .B(n9142), .ZN(n9381) );
  XNOR2_X1 U10496 ( .A(n9145), .B(n9144), .ZN(n9147) );
  OAI21_X1 U10497 ( .B1(n9147), .B2(n9240), .A(n9146), .ZN(n9378) );
  AOI211_X1 U10498 ( .C1(n9379), .C2(n9162), .A(n9342), .B(n9136), .ZN(n9377)
         );
  NAND2_X1 U10499 ( .A1(n9377), .A2(n9350), .ZN(n9151) );
  AOI22_X1 U10500 ( .A1(n9304), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9149), .B2(
        n9302), .ZN(n9150) );
  OAI211_X1 U10501 ( .C1(n9152), .C2(n9345), .A(n9151), .B(n9150), .ZN(n9153)
         );
  AOI21_X1 U10502 ( .B1(n9378), .B2(n9678), .A(n9153), .ZN(n9154) );
  OAI21_X1 U10503 ( .B1(n9381), .B2(n9309), .A(n9154), .ZN(P1_U3266) );
  NAND2_X1 U10504 ( .A1(n9172), .A2(n9155), .ZN(n9156) );
  XNOR2_X1 U10505 ( .A(n9156), .B(n9160), .ZN(n9157) );
  OR2_X1 U10506 ( .A1(n9157), .A2(n9240), .ZN(n9159) );
  NAND2_X1 U10507 ( .A1(n9159), .A2(n9158), .ZN(n9382) );
  INV_X1 U10508 ( .A(n9382), .ZN(n9171) );
  XNOR2_X1 U10509 ( .A(n9161), .B(n9160), .ZN(n9384) );
  NAND2_X1 U10510 ( .A1(n9384), .A2(n9339), .ZN(n9170) );
  INV_X1 U10511 ( .A(n9162), .ZN(n9163) );
  AOI211_X1 U10512 ( .C1(n9164), .C2(n4625), .A(n9342), .B(n9163), .ZN(n9383)
         );
  NOR2_X1 U10513 ( .A1(n9464), .A2(n9345), .ZN(n9168) );
  OAI22_X1 U10514 ( .A1(n9678), .A2(n9166), .B1(n9165), .B2(n9673), .ZN(n9167)
         );
  AOI211_X1 U10515 ( .C1(n9383), .C2(n9350), .A(n9168), .B(n9167), .ZN(n9169)
         );
  OAI211_X1 U10516 ( .C1(n9304), .C2(n9171), .A(n9170), .B(n9169), .ZN(
        P1_U3267) );
  OAI211_X1 U10517 ( .C1(n9178), .C2(n9173), .A(n9172), .B(n9333), .ZN(n9176)
         );
  INV_X1 U10518 ( .A(n9174), .ZN(n9175) );
  NAND2_X1 U10519 ( .A1(n9176), .A2(n9175), .ZN(n9387) );
  INV_X1 U10520 ( .A(n9387), .ZN(n9187) );
  XOR2_X1 U10521 ( .A(n9178), .B(n9177), .Z(n9389) );
  NAND2_X1 U10522 ( .A1(n9389), .A2(n9339), .ZN(n9186) );
  AOI211_X1 U10523 ( .C1(n9180), .C2(n9196), .A(n9342), .B(n9179), .ZN(n9388)
         );
  NOR2_X1 U10524 ( .A1(n4623), .A2(n9345), .ZN(n9184) );
  OAI22_X1 U10525 ( .A1(n9182), .A2(n9673), .B1(n9181), .B2(n9678), .ZN(n9183)
         );
  AOI211_X1 U10526 ( .C1(n9388), .C2(n9350), .A(n9184), .B(n9183), .ZN(n9185)
         );
  OAI211_X1 U10527 ( .C1(n9304), .C2(n9187), .A(n9186), .B(n9185), .ZN(
        P1_U3268) );
  XOR2_X1 U10528 ( .A(n9189), .B(n9188), .Z(n9396) );
  AOI21_X1 U10529 ( .B1(n9190), .B2(n9207), .A(n9189), .ZN(n9195) );
  NAND2_X1 U10530 ( .A1(n9191), .A2(n9333), .ZN(n9194) );
  INV_X1 U10531 ( .A(n9192), .ZN(n9193) );
  OAI21_X1 U10532 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9392) );
  INV_X1 U10533 ( .A(n9196), .ZN(n9197) );
  AOI211_X1 U10534 ( .C1(n9394), .C2(n9215), .A(n9342), .B(n9197), .ZN(n9393)
         );
  NAND2_X1 U10535 ( .A1(n9393), .A2(n9350), .ZN(n9200) );
  AOI22_X1 U10536 ( .A1(n9198), .A2(n9302), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9304), .ZN(n9199) );
  OAI211_X1 U10537 ( .C1(n9201), .C2(n9345), .A(n9200), .B(n9199), .ZN(n9202)
         );
  AOI21_X1 U10538 ( .B1(n9678), .B2(n9392), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10539 ( .B1(n9396), .B2(n9309), .A(n9203), .ZN(P1_U3269) );
  INV_X1 U10540 ( .A(n9212), .ZN(n9206) );
  NAND2_X1 U10541 ( .A1(n9227), .A2(n9204), .ZN(n9205) );
  NAND2_X1 U10542 ( .A1(n9206), .A2(n9205), .ZN(n9208) );
  NAND2_X1 U10543 ( .A1(n9208), .A2(n9207), .ZN(n9210) );
  AOI21_X1 U10544 ( .B1(n9210), .B2(n9333), .A(n9209), .ZN(n9398) );
  XOR2_X1 U10545 ( .A(n9212), .B(n9211), .Z(n9399) );
  OR2_X1 U10546 ( .A1(n9399), .A2(n9309), .ZN(n9221) );
  OAI22_X1 U10547 ( .A1(n9214), .A2(n9673), .B1(n9213), .B2(n9678), .ZN(n9218)
         );
  OAI211_X1 U10548 ( .C1(n9472), .C2(n9230), .A(n9216), .B(n9215), .ZN(n9397)
         );
  NOR2_X1 U10549 ( .A1(n9397), .A2(n9660), .ZN(n9217) );
  AOI211_X1 U10550 ( .C1(n9657), .C2(n9219), .A(n9218), .B(n9217), .ZN(n9220)
         );
  OAI211_X1 U10551 ( .C1(n9304), .C2(n9398), .A(n9221), .B(n9220), .ZN(
        P1_U3270) );
  XNOR2_X1 U10552 ( .A(n9223), .B(n9222), .ZN(n9405) );
  INV_X1 U10553 ( .A(n9405), .ZN(n9237) );
  NAND2_X1 U10554 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND3_X1 U10555 ( .A1(n9227), .A2(n9333), .A3(n9226), .ZN(n9229) );
  NAND2_X1 U10556 ( .A1(n9229), .A2(n9228), .ZN(n9403) );
  AOI211_X1 U10557 ( .C1(n9231), .C2(n9244), .A(n9342), .B(n9230), .ZN(n9404)
         );
  NAND2_X1 U10558 ( .A1(n9404), .A2(n9350), .ZN(n9234) );
  AOI22_X1 U10559 ( .A1(n9232), .A2(n9302), .B1(n9304), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9233) );
  OAI211_X1 U10560 ( .C1(n9476), .C2(n9345), .A(n9234), .B(n9233), .ZN(n9235)
         );
  AOI21_X1 U10561 ( .B1(n9678), .B2(n9403), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10562 ( .B1(n9237), .B2(n9309), .A(n9236), .ZN(P1_U3271) );
  XNOR2_X1 U10563 ( .A(n9238), .B(n9242), .ZN(n9241) );
  OAI21_X1 U10564 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9407) );
  INV_X1 U10565 ( .A(n9407), .ZN(n9253) );
  XNOR2_X1 U10566 ( .A(n9243), .B(n9242), .ZN(n9409) );
  NAND2_X1 U10567 ( .A1(n9409), .A2(n9339), .ZN(n9252) );
  INV_X1 U10568 ( .A(n9244), .ZN(n9245) );
  AOI211_X1 U10569 ( .C1(n9246), .C2(n9261), .A(n9342), .B(n9245), .ZN(n9408)
         );
  NOR2_X1 U10570 ( .A1(n9101), .A2(n9345), .ZN(n9250) );
  OAI22_X1 U10571 ( .A1(n9248), .A2(n9673), .B1(n9678), .B2(n9247), .ZN(n9249)
         );
  AOI211_X1 U10572 ( .C1(n9408), .C2(n9350), .A(n9250), .B(n9249), .ZN(n9251)
         );
  OAI211_X1 U10573 ( .C1(n9304), .C2(n9253), .A(n9252), .B(n9251), .ZN(
        P1_U3272) );
  XOR2_X1 U10574 ( .A(n9256), .B(n9254), .Z(n9414) );
  INV_X1 U10575 ( .A(n9414), .ZN(n9269) );
  OAI211_X1 U10576 ( .C1(n9258), .C2(n4430), .A(n9257), .B(n9333), .ZN(n9260)
         );
  NAND2_X1 U10577 ( .A1(n9260), .A2(n9259), .ZN(n9412) );
  INV_X1 U10578 ( .A(n9261), .ZN(n9262) );
  AOI211_X1 U10579 ( .C1(n9263), .C2(n9277), .A(n9342), .B(n9262), .ZN(n9413)
         );
  NAND2_X1 U10580 ( .A1(n9413), .A2(n9350), .ZN(n9266) );
  AOI22_X1 U10581 ( .A1(n9304), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9264), .B2(
        n9302), .ZN(n9265) );
  OAI211_X1 U10582 ( .C1(n9483), .C2(n9345), .A(n9266), .B(n9265), .ZN(n9267)
         );
  AOI21_X1 U10583 ( .B1(n9678), .B2(n9412), .A(n9267), .ZN(n9268) );
  OAI21_X1 U10584 ( .B1(n9269), .B2(n9309), .A(n9268), .ZN(P1_U3273) );
  XNOR2_X1 U10585 ( .A(n9271), .B(n9272), .ZN(n9419) );
  INV_X1 U10586 ( .A(n9419), .ZN(n9286) );
  XNOR2_X1 U10587 ( .A(n9273), .B(n9272), .ZN(n9274) );
  NAND2_X1 U10588 ( .A1(n9274), .A2(n9333), .ZN(n9276) );
  NAND2_X1 U10589 ( .A1(n9276), .A2(n9275), .ZN(n9417) );
  INV_X1 U10590 ( .A(n9277), .ZN(n9278) );
  AOI211_X1 U10591 ( .C1(n9279), .C2(n4633), .A(n9342), .B(n9278), .ZN(n9418)
         );
  NAND2_X1 U10592 ( .A1(n9418), .A2(n9350), .ZN(n9283) );
  INV_X1 U10593 ( .A(n9280), .ZN(n9281) );
  AOI22_X1 U10594 ( .A1(n9304), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9281), .B2(
        n9302), .ZN(n9282) );
  OAI211_X1 U10595 ( .C1(n9487), .C2(n9345), .A(n9283), .B(n9282), .ZN(n9284)
         );
  AOI21_X1 U10596 ( .B1(n9678), .B2(n9417), .A(n9284), .ZN(n9285) );
  OAI21_X1 U10597 ( .B1(n9286), .B2(n9309), .A(n9285), .ZN(P1_U3274) );
  XNOR2_X1 U10598 ( .A(n9288), .B(n9290), .ZN(n9424) );
  INV_X1 U10599 ( .A(n9424), .ZN(n9310) );
  NAND2_X1 U10600 ( .A1(n9311), .A2(n9289), .ZN(n9292) );
  INV_X1 U10601 ( .A(n9290), .ZN(n9291) );
  NAND2_X1 U10602 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  NAND2_X1 U10603 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U10604 ( .A1(n9295), .A2(n9333), .ZN(n9298) );
  INV_X1 U10605 ( .A(n9296), .ZN(n9297) );
  NAND2_X1 U10606 ( .A1(n9298), .A2(n9297), .ZN(n9422) );
  AOI211_X1 U10607 ( .C1(n9300), .C2(n9318), .A(n9342), .B(n9299), .ZN(n9423)
         );
  NAND2_X1 U10608 ( .A1(n9423), .A2(n9350), .ZN(n9306) );
  INV_X1 U10609 ( .A(n9301), .ZN(n9303) );
  AOI22_X1 U10610 ( .A1(n9304), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9303), .B2(
        n9302), .ZN(n9305) );
  OAI211_X1 U10611 ( .C1(n9491), .C2(n9345), .A(n9306), .B(n9305), .ZN(n9307)
         );
  AOI21_X1 U10612 ( .B1(n9678), .B2(n9422), .A(n9307), .ZN(n9308) );
  OAI21_X1 U10613 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(P1_U3275) );
  OAI211_X1 U10614 ( .C1(n9313), .C2(n9312), .A(n9311), .B(n9333), .ZN(n9315)
         );
  NAND2_X1 U10615 ( .A1(n9315), .A2(n9314), .ZN(n9427) );
  INV_X1 U10616 ( .A(n9427), .ZN(n9328) );
  XNOR2_X1 U10617 ( .A(n9317), .B(n9316), .ZN(n9429) );
  NAND2_X1 U10618 ( .A1(n9429), .A2(n9339), .ZN(n9327) );
  INV_X1 U10619 ( .A(n9341), .ZN(n9320) );
  INV_X1 U10620 ( .A(n9318), .ZN(n9319) );
  AOI211_X1 U10621 ( .C1(n9321), .C2(n9320), .A(n9342), .B(n9319), .ZN(n9428)
         );
  NOR2_X1 U10622 ( .A1(n9495), .A2(n9345), .ZN(n9325) );
  OAI22_X1 U10623 ( .A1(n9678), .A2(n9323), .B1(n9322), .B2(n9673), .ZN(n9324)
         );
  AOI211_X1 U10624 ( .C1(n9428), .C2(n9350), .A(n9325), .B(n9324), .ZN(n9326)
         );
  OAI211_X1 U10625 ( .C1(n9304), .C2(n9328), .A(n9327), .B(n9326), .ZN(
        P1_U3276) );
  NAND2_X1 U10626 ( .A1(n9330), .A2(n9329), .ZN(n9332) );
  INV_X1 U10627 ( .A(n9337), .ZN(n9331) );
  XNOR2_X1 U10628 ( .A(n9332), .B(n9331), .ZN(n9334) );
  NAND2_X1 U10629 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  NAND2_X1 U10630 ( .A1(n9336), .A2(n9335), .ZN(n9432) );
  INV_X1 U10631 ( .A(n9432), .ZN(n9353) );
  XOR2_X1 U10632 ( .A(n9338), .B(n9337), .Z(n9434) );
  NAND2_X1 U10633 ( .A1(n9434), .A2(n9339), .ZN(n9352) );
  INV_X1 U10634 ( .A(n9340), .ZN(n9343) );
  AOI211_X1 U10635 ( .C1(n9344), .C2(n9343), .A(n9342), .B(n9341), .ZN(n9433)
         );
  NOR2_X1 U10636 ( .A1(n9499), .A2(n9345), .ZN(n9349) );
  OAI22_X1 U10637 ( .A1(n9678), .A2(n9347), .B1(n9346), .B2(n9673), .ZN(n9348)
         );
  AOI211_X1 U10638 ( .C1(n9433), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9351)
         );
  OAI211_X1 U10639 ( .C1(n9304), .C2(n9353), .A(n9352), .B(n9351), .ZN(
        P1_U3277) );
  NOR2_X1 U10640 ( .A1(n9355), .A2(n9354), .ZN(n9448) );
  MUX2_X1 U10641 ( .A(n9356), .B(n9448), .S(n9712), .Z(n9357) );
  OAI21_X1 U10642 ( .B1(n9451), .B2(n9440), .A(n9357), .ZN(P1_U3553) );
  AND2_X1 U10643 ( .A1(n9359), .A2(n9358), .ZN(n9453) );
  MUX2_X1 U10644 ( .A(n9360), .B(n9453), .S(n9712), .Z(n9361) );
  OAI21_X1 U10645 ( .B1(n8720), .B2(n9440), .A(n9361), .ZN(P1_U3552) );
  NAND2_X1 U10646 ( .A1(n9046), .A2(n9367), .ZN(n9368) );
  NAND2_X1 U10647 ( .A1(n9369), .A2(n9368), .ZN(P1_U3551) );
  NAND3_X1 U10648 ( .A1(n9371), .A2(n9370), .A3(n9695), .ZN(n9376) );
  AOI21_X1 U10649 ( .B1(n9443), .B2(n9373), .A(n9372), .ZN(n9374) );
  NAND3_X1 U10650 ( .A1(n9376), .A2(n9375), .A3(n9374), .ZN(n9459) );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9459), .S(n9712), .Z(
        P1_U3550) );
  AOI211_X1 U10652 ( .C1(n9443), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9380)
         );
  OAI21_X1 U10653 ( .B1(n9381), .B2(n9446), .A(n9380), .ZN(n9460) );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9460), .S(n9712), .Z(
        P1_U3549) );
  AOI211_X1 U10655 ( .C1(n9384), .C2(n9695), .A(n9383), .B(n9382), .ZN(n9461)
         );
  MUX2_X1 U10656 ( .A(n9385), .B(n9461), .S(n9712), .Z(n9386) );
  OAI21_X1 U10657 ( .B1(n9464), .B2(n9440), .A(n9386), .ZN(P1_U3548) );
  AOI211_X1 U10658 ( .C1(n9389), .C2(n9695), .A(n9388), .B(n9387), .ZN(n9465)
         );
  MUX2_X1 U10659 ( .A(n9390), .B(n9465), .S(n9712), .Z(n9391) );
  OAI21_X1 U10660 ( .B1(n4623), .B2(n9440), .A(n9391), .ZN(P1_U3547) );
  AOI211_X1 U10661 ( .C1(n9443), .C2(n9394), .A(n9393), .B(n9392), .ZN(n9395)
         );
  OAI21_X1 U10662 ( .B1(n9396), .B2(n9446), .A(n9395), .ZN(n9468) );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9468), .S(n9712), .Z(
        P1_U3546) );
  OAI211_X1 U10664 ( .C1(n9399), .C2(n9446), .A(n9398), .B(n9397), .ZN(n9400)
         );
  INV_X1 U10665 ( .A(n9400), .ZN(n9469) );
  MUX2_X1 U10666 ( .A(n9401), .B(n9469), .S(n9712), .Z(n9402) );
  OAI21_X1 U10667 ( .B1(n9472), .B2(n9440), .A(n9402), .ZN(P1_U3545) );
  AOI211_X1 U10668 ( .C1(n9405), .C2(n9695), .A(n9404), .B(n9403), .ZN(n9473)
         );
  MUX2_X1 U10669 ( .A(n9945), .B(n9473), .S(n9712), .Z(n9406) );
  OAI21_X1 U10670 ( .B1(n9476), .B2(n9440), .A(n9406), .ZN(P1_U3544) );
  AOI211_X1 U10671 ( .C1(n9409), .C2(n9695), .A(n9408), .B(n9407), .ZN(n9477)
         );
  MUX2_X1 U10672 ( .A(n9410), .B(n9477), .S(n9712), .Z(n9411) );
  OAI21_X1 U10673 ( .B1(n9101), .B2(n9440), .A(n9411), .ZN(P1_U3543) );
  AOI211_X1 U10674 ( .C1(n9414), .C2(n9695), .A(n9413), .B(n9412), .ZN(n9480)
         );
  MUX2_X1 U10675 ( .A(n9415), .B(n9480), .S(n9712), .Z(n9416) );
  OAI21_X1 U10676 ( .B1(n9483), .B2(n9440), .A(n9416), .ZN(P1_U3542) );
  AOI211_X1 U10677 ( .C1(n9419), .C2(n9695), .A(n9418), .B(n9417), .ZN(n9484)
         );
  MUX2_X1 U10678 ( .A(n9420), .B(n9484), .S(n9712), .Z(n9421) );
  OAI21_X1 U10679 ( .B1(n9487), .B2(n9440), .A(n9421), .ZN(P1_U3541) );
  INV_X1 U10680 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9425) );
  AOI211_X1 U10681 ( .C1(n9424), .C2(n9695), .A(n9423), .B(n9422), .ZN(n9488)
         );
  MUX2_X1 U10682 ( .A(n9425), .B(n9488), .S(n9712), .Z(n9426) );
  OAI21_X1 U10683 ( .B1(n9491), .B2(n9440), .A(n9426), .ZN(P1_U3540) );
  AOI211_X1 U10684 ( .C1(n9429), .C2(n9695), .A(n9428), .B(n9427), .ZN(n9492)
         );
  MUX2_X1 U10685 ( .A(n9430), .B(n9492), .S(n9712), .Z(n9431) );
  OAI21_X1 U10686 ( .B1(n9495), .B2(n9440), .A(n9431), .ZN(P1_U3539) );
  AOI211_X1 U10687 ( .C1(n9434), .C2(n9695), .A(n9433), .B(n9432), .ZN(n9496)
         );
  MUX2_X1 U10688 ( .A(n9999), .B(n9496), .S(n9712), .Z(n9435) );
  OAI21_X1 U10689 ( .B1(n9499), .B2(n9440), .A(n9435), .ZN(P1_U3538) );
  AOI211_X1 U10690 ( .C1(n9438), .C2(n9695), .A(n9437), .B(n9436), .ZN(n9500)
         );
  MUX2_X1 U10691 ( .A(n9621), .B(n9500), .S(n9712), .Z(n9439) );
  OAI21_X1 U10692 ( .B1(n9504), .B2(n9440), .A(n9439), .ZN(P1_U3537) );
  AOI21_X1 U10693 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9444) );
  OAI211_X1 U10694 ( .C1(n9447), .C2(n9446), .A(n9445), .B(n9444), .ZN(n9505)
         );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9505), .S(n9712), .Z(
        P1_U3536) );
  MUX2_X1 U10696 ( .A(n9449), .B(n9448), .S(n9707), .Z(n9450) );
  OAI21_X1 U10697 ( .B1(n9451), .B2(n9503), .A(n9450), .ZN(P1_U3521) );
  MUX2_X1 U10698 ( .A(n9453), .B(n9452), .S(n9706), .Z(n9454) );
  OAI21_X1 U10699 ( .B1(n8720), .B2(n9503), .A(n9454), .ZN(P1_U3520) );
  NAND2_X1 U10700 ( .A1(n9046), .A2(n9456), .ZN(n9457) );
  NAND2_X1 U10701 ( .A1(n9458), .A2(n9457), .ZN(P1_U3519) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9459), .S(n9707), .Z(
        P1_U3518) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9460), .S(n9707), .Z(
        P1_U3517) );
  MUX2_X1 U10704 ( .A(n9462), .B(n9461), .S(n9707), .Z(n9463) );
  OAI21_X1 U10705 ( .B1(n9464), .B2(n9503), .A(n9463), .ZN(P1_U3516) );
  MUX2_X1 U10706 ( .A(n9466), .B(n9465), .S(n9707), .Z(n9467) );
  OAI21_X1 U10707 ( .B1(n4623), .B2(n9503), .A(n9467), .ZN(P1_U3515) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9468), .S(n9707), .Z(
        P1_U3514) );
  MUX2_X1 U10709 ( .A(n9470), .B(n9469), .S(n9707), .Z(n9471) );
  OAI21_X1 U10710 ( .B1(n9472), .B2(n9503), .A(n9471), .ZN(P1_U3513) );
  MUX2_X1 U10711 ( .A(n9474), .B(n9473), .S(n9707), .Z(n9475) );
  OAI21_X1 U10712 ( .B1(n9476), .B2(n9503), .A(n9475), .ZN(P1_U3512) );
  MUX2_X1 U10713 ( .A(n9478), .B(n9477), .S(n9707), .Z(n9479) );
  OAI21_X1 U10714 ( .B1(n9101), .B2(n9503), .A(n9479), .ZN(P1_U3511) );
  MUX2_X1 U10715 ( .A(n9481), .B(n9480), .S(n9707), .Z(n9482) );
  OAI21_X1 U10716 ( .B1(n9483), .B2(n9503), .A(n9482), .ZN(P1_U3510) );
  INV_X1 U10717 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9485) );
  MUX2_X1 U10718 ( .A(n9485), .B(n9484), .S(n9707), .Z(n9486) );
  OAI21_X1 U10719 ( .B1(n9487), .B2(n9503), .A(n9486), .ZN(P1_U3509) );
  MUX2_X1 U10720 ( .A(n9489), .B(n9488), .S(n9707), .Z(n9490) );
  OAI21_X1 U10721 ( .B1(n9491), .B2(n9503), .A(n9490), .ZN(P1_U3507) );
  INV_X1 U10722 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U10723 ( .A(n9493), .B(n9492), .S(n9707), .Z(n9494) );
  OAI21_X1 U10724 ( .B1(n9495), .B2(n9503), .A(n9494), .ZN(P1_U3504) );
  MUX2_X1 U10725 ( .A(n9497), .B(n9496), .S(n9707), .Z(n9498) );
  OAI21_X1 U10726 ( .B1(n9499), .B2(n9503), .A(n9498), .ZN(P1_U3501) );
  MUX2_X1 U10727 ( .A(n9501), .B(n9500), .S(n9707), .Z(n9502) );
  OAI21_X1 U10728 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(P1_U3498) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9505), .S(n9707), .Z(
        P1_U3495) );
  MUX2_X1 U10730 ( .A(n9506), .B(P1_D_REG_1__SCAN_IN), .S(n9681), .Z(P1_U3440)
         );
  NOR3_X1 U10731 ( .A1(n9507), .A2(n5386), .A3(P1_U3086), .ZN(n9508) );
  AOI21_X1 U10732 ( .B1(n9509), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9508), .ZN(
        n9510) );
  OAI21_X1 U10733 ( .B1(n9511), .B2(n9514), .A(n9510), .ZN(P1_U3324) );
  OAI222_X1 U10734 ( .A1(n9522), .A2(n9515), .B1(n9514), .B2(n9513), .C1(
        P1_U3086), .C2(n9512), .ZN(P1_U3325) );
  OAI222_X1 U10735 ( .A1(n9514), .A2(n9518), .B1(P1_U3086), .B2(n9516), .C1(
        n9956), .C2(n9522), .ZN(P1_U3326) );
  OAI222_X1 U10736 ( .A1(n9514), .A2(n9521), .B1(n9520), .B2(P1_U3086), .C1(
        n9519), .C2(n9522), .ZN(P1_U3327) );
  OAI222_X1 U10737 ( .A1(n9514), .A2(n9524), .B1(P1_U3086), .B2(n9523), .C1(
        n9933), .C2(n9522), .ZN(P1_U3328) );
  MUX2_X1 U10738 ( .A(n9525), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10739 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9536) );
  AOI211_X1 U10740 ( .C1(n9528), .C2(n9527), .A(n9526), .B(n9623), .ZN(n9533)
         );
  AOI211_X1 U10741 ( .C1(n9531), .C2(n9530), .A(n9529), .B(n9619), .ZN(n9532)
         );
  AOI211_X1 U10742 ( .C1(n9630), .C2(n9534), .A(n9533), .B(n9532), .ZN(n9535)
         );
  NAND2_X1 U10743 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9563) );
  OAI211_X1 U10744 ( .C1(n9650), .C2(n9536), .A(n9535), .B(n9563), .ZN(
        P1_U3253) );
  XNOR2_X1 U10745 ( .A(n9537), .B(n4589), .ZN(n9557) );
  INV_X1 U10746 ( .A(n9538), .ZN(n9539) );
  NOR2_X1 U10747 ( .A1(n9539), .A2(n9793), .ZN(n9556) );
  INV_X1 U10748 ( .A(n9556), .ZN(n9543) );
  OAI22_X1 U10749 ( .A1(n9543), .A2(n9542), .B1(n9541), .B2(n9540), .ZN(n9551)
         );
  XNOR2_X1 U10750 ( .A(n9544), .B(n4589), .ZN(n9545) );
  OAI222_X1 U10751 ( .A1(n9550), .A2(n9549), .B1(n9548), .B2(n9547), .C1(n9546), .C2(n9545), .ZN(n9555) );
  AOI211_X1 U10752 ( .C1(n9557), .C2(n9552), .A(n9551), .B(n9555), .ZN(n9553)
         );
  AOI22_X1 U10753 ( .A1(n9757), .A2(n9554), .B1(n9553), .B2(n8268), .ZN(
        P2_U3220) );
  AOI211_X1 U10754 ( .C1(n9557), .C2(n9811), .A(n9556), .B(n9555), .ZN(n9558)
         );
  AOI22_X1 U10755 ( .A1(n4275), .A2(n9558), .B1(n7388), .B2(n9833), .ZN(
        P2_U3472) );
  INV_X1 U10756 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10757 ( .A1(n9819), .A2(n9559), .B1(n9558), .B2(n9817), .ZN(
        P2_U3429) );
  OAI21_X1 U10758 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9572) );
  INV_X1 U10759 ( .A(n9563), .ZN(n9564) );
  AOI21_X1 U10760 ( .B1(n9566), .B2(n9565), .A(n9564), .ZN(n9567) );
  OAI21_X1 U10761 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9570) );
  AOI21_X1 U10762 ( .B1(n9572), .B2(n9571), .A(n9570), .ZN(n9573) );
  OAI21_X1 U10763 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(P1_U3217) );
  XNOR2_X1 U10764 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10765 ( .A(P2_RD_REG_SCAN_IN), .B(n4579), .Z(U126) );
  INV_X1 U10766 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9588) );
  OAI211_X1 U10767 ( .C1(n9578), .C2(n9577), .A(n9634), .B(n9576), .ZN(n9585)
         );
  NAND2_X1 U10768 ( .A1(n9630), .A2(n9579), .ZN(n9584) );
  OAI211_X1 U10769 ( .C1(n9582), .C2(n9581), .A(n9642), .B(n9580), .ZN(n9583)
         );
  AND3_X1 U10770 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(n9587) );
  NAND2_X1 U10771 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9586) );
  OAI211_X1 U10772 ( .C1(n9650), .C2(n9588), .A(n9587), .B(n9586), .ZN(
        P1_U3254) );
  INV_X1 U10773 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9603) );
  AOI21_X1 U10774 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(n9592) );
  NAND2_X1 U10775 ( .A1(n9634), .A2(n9592), .ZN(n9600) );
  NAND2_X1 U10776 ( .A1(n9630), .A2(n9593), .ZN(n9599) );
  AOI21_X1 U10777 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9597) );
  NAND2_X1 U10778 ( .A1(n9642), .A2(n9597), .ZN(n9598) );
  AND3_X1 U10779 ( .A1(n9600), .A2(n9599), .A3(n9598), .ZN(n9602) );
  NAND2_X1 U10780 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9601) );
  OAI211_X1 U10781 ( .C1(n9650), .C2(n9603), .A(n9602), .B(n9601), .ZN(
        P1_U3256) );
  INV_X1 U10782 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9618) );
  AOI21_X1 U10783 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  NAND2_X1 U10784 ( .A1(n9634), .A2(n9607), .ZN(n9615) );
  NAND2_X1 U10785 ( .A1(n9630), .A2(n9608), .ZN(n9614) );
  AOI21_X1 U10786 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9612) );
  NAND2_X1 U10787 ( .A1(n9642), .A2(n9612), .ZN(n9613) );
  AND3_X1 U10788 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n9617) );
  NAND2_X1 U10789 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9616) );
  OAI211_X1 U10790 ( .C1(n9650), .C2(n9618), .A(n9617), .B(n9616), .ZN(
        P1_U3257) );
  INV_X1 U10791 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9633) );
  AOI211_X1 U10792 ( .C1(n9622), .C2(n9621), .A(n9620), .B(n9619), .ZN(n9628)
         );
  AOI211_X1 U10793 ( .C1(n9626), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9627)
         );
  AOI211_X1 U10794 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9632)
         );
  NAND2_X1 U10795 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9631) );
  OAI211_X1 U10796 ( .C1(n9650), .C2(n9633), .A(n9632), .B(n9631), .ZN(
        P1_U3258) );
  OAI211_X1 U10797 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9644)
         );
  NAND2_X1 U10798 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  NAND3_X1 U10799 ( .A1(n9642), .A2(n9641), .A3(n9640), .ZN(n9643) );
  OAI211_X1 U10800 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9647)
         );
  INV_X1 U10801 ( .A(n9647), .ZN(n9649) );
  NAND2_X1 U10802 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9648) );
  OAI211_X1 U10803 ( .C1(n9650), .C2(n9841), .A(n9649), .B(n9648), .ZN(
        P1_U3261) );
  NAND2_X1 U10804 ( .A1(n9652), .A2(n9651), .ZN(n9664) );
  OAI22_X1 U10805 ( .A1(n9678), .A2(n9654), .B1(n9653), .B2(n9673), .ZN(n9655)
         );
  INV_X1 U10806 ( .A(n9655), .ZN(n9663) );
  NAND2_X1 U10807 ( .A1(n9657), .A2(n9656), .ZN(n9662) );
  INV_X1 U10808 ( .A(n9658), .ZN(n9659) );
  OR2_X1 U10809 ( .A1(n9660), .A2(n9659), .ZN(n9661) );
  AND4_X1 U10810 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9665)
         );
  OAI21_X1 U10811 ( .B1(n9304), .B2(n9666), .A(n9665), .ZN(P1_U3291) );
  INV_X1 U10812 ( .A(n9667), .ZN(n9677) );
  INV_X1 U10813 ( .A(n9668), .ZN(n9676) );
  INV_X1 U10814 ( .A(n9669), .ZN(n9670) );
  OAI22_X1 U10815 ( .A1(n9673), .A2(n9672), .B1(n9671), .B2(n9670), .ZN(n9674)
         );
  AOI211_X1 U10816 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9679)
         );
  AOI22_X1 U10817 ( .A1(n9304), .A2(n5039), .B1(n9679), .B2(n9678), .ZN(
        P1_U3293) );
  AND2_X1 U10818 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9681), .ZN(P1_U3294) );
  AND2_X1 U10819 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9681), .ZN(P1_U3295) );
  AND2_X1 U10820 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9681), .ZN(P1_U3296) );
  AND2_X1 U10821 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9681), .ZN(P1_U3297) );
  AND2_X1 U10822 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9681), .ZN(P1_U3298) );
  AND2_X1 U10823 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9681), .ZN(P1_U3299) );
  AND2_X1 U10824 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9681), .ZN(P1_U3300) );
  AND2_X1 U10825 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9681), .ZN(P1_U3301) );
  INV_X1 U10826 ( .A(n9681), .ZN(n9680) );
  INV_X1 U10827 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9983) );
  NOR2_X1 U10828 ( .A1(n9680), .A2(n9983), .ZN(P1_U3302) );
  AND2_X1 U10829 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9681), .ZN(P1_U3303) );
  AND2_X1 U10830 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9681), .ZN(P1_U3304) );
  AND2_X1 U10831 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9681), .ZN(P1_U3305) );
  AND2_X1 U10832 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9681), .ZN(P1_U3306) );
  AND2_X1 U10833 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9681), .ZN(P1_U3307) );
  AND2_X1 U10834 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9681), .ZN(P1_U3308) );
  AND2_X1 U10835 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9681), .ZN(P1_U3309) );
  AND2_X1 U10836 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9681), .ZN(P1_U3310) );
  AND2_X1 U10837 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9681), .ZN(P1_U3311) );
  AND2_X1 U10838 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9681), .ZN(P1_U3312) );
  INV_X1 U10839 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U10840 ( .A1(n9680), .A2(n9918), .ZN(P1_U3313) );
  AND2_X1 U10841 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9681), .ZN(P1_U3314) );
  AND2_X1 U10842 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9681), .ZN(P1_U3315) );
  AND2_X1 U10843 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9681), .ZN(P1_U3316) );
  AND2_X1 U10844 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9681), .ZN(P1_U3317) );
  AND2_X1 U10845 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9681), .ZN(P1_U3318) );
  AND2_X1 U10846 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9681), .ZN(P1_U3319) );
  AND2_X1 U10847 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9681), .ZN(P1_U3320) );
  AND2_X1 U10848 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9681), .ZN(P1_U3321) );
  AND2_X1 U10849 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9681), .ZN(P1_U3322) );
  AND2_X1 U10850 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9681), .ZN(P1_U3323) );
  AOI22_X1 U10851 ( .A1(n9707), .A2(n9682), .B1(n5038), .B2(n9706), .ZN(
        P1_U3453) );
  OAI21_X1 U10852 ( .B1(n9684), .B2(n9698), .A(n9683), .ZN(n9685) );
  AOI21_X1 U10853 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  AOI22_X1 U10854 ( .A1(n9707), .A2(n9708), .B1(n5158), .B2(n9706), .ZN(
        P1_U3474) );
  OAI211_X1 U10855 ( .C1(n4647), .C2(n9698), .A(n9692), .B(n9691), .ZN(n9693)
         );
  AOI21_X1 U10856 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9709) );
  AOI22_X1 U10857 ( .A1(n9707), .A2(n9709), .B1(n5213), .B2(n9706), .ZN(
        P1_U3480) );
  OAI211_X1 U10858 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9703)
         );
  INV_X1 U10859 ( .A(n9704), .ZN(n9701) );
  NOR2_X1 U10860 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  AOI211_X1 U10861 ( .C1(n9705), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9711)
         );
  AOI22_X1 U10862 ( .A1(n9707), .A2(n9711), .B1(n5271), .B2(n9706), .ZN(
        P1_U3486) );
  AOI22_X1 U10863 ( .A1(n9712), .A2(n9708), .B1(n6898), .B2(n9710), .ZN(
        P1_U3529) );
  AOI22_X1 U10864 ( .A1(n9712), .A2(n9709), .B1(n5208), .B2(n9710), .ZN(
        P1_U3531) );
  AOI22_X1 U10865 ( .A1(n9712), .A2(n9711), .B1(n5268), .B2(n9710), .ZN(
        P1_U3533) );
  AOI22_X1 U10866 ( .A1(n9882), .A2(n9714), .B1(n9713), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9727) );
  OAI21_X1 U10867 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9716), .A(n9715), .ZN(
        n9721) );
  XNOR2_X1 U10868 ( .A(n9718), .B(n9717), .ZN(n9719) );
  AOI22_X1 U10869 ( .A1(n9721), .A2(n9720), .B1(n9887), .B2(n9719), .ZN(n9726)
         );
  NAND2_X1 U10870 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n9725) );
  NOR2_X1 U10871 ( .A1(n4286), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9723) );
  OAI21_X1 U10872 ( .B1(n9723), .B2(n9722), .A(n9874), .ZN(n9724) );
  NAND4_X1 U10873 ( .A1(n9727), .A2(n9726), .A3(n9725), .A4(n9724), .ZN(
        P2_U3199) );
  XOR2_X1 U10874 ( .A(n9728), .B(n9732), .Z(n9731) );
  AOI222_X1 U10875 ( .A1(n9748), .A2(n9731), .B1(n9730), .B2(n9745), .C1(n9729), .C2(n9743), .ZN(n9788) );
  INV_X1 U10876 ( .A(n9732), .ZN(n9733) );
  NAND3_X1 U10877 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n9736) );
  NAND2_X1 U10878 ( .A1(n9737), .A2(n9736), .ZN(n9790) );
  INV_X1 U10879 ( .A(n9790), .ZN(n9739) );
  AOI222_X1 U10880 ( .A1(n9740), .A2(n9752), .B1(n9739), .B2(n9754), .C1(n9738), .C2(n9750), .ZN(n9741) );
  OAI221_X1 U10881 ( .B1(n9757), .B2(n9788), .C1(n8291), .C2(n6765), .A(n9741), 
        .ZN(P2_U3225) );
  XOR2_X1 U10882 ( .A(n9742), .B(n9749), .Z(n9747) );
  AOI222_X1 U10883 ( .A1(n9748), .A2(n9747), .B1(n9746), .B2(n9745), .C1(n9744), .C2(n9743), .ZN(n9762) );
  INV_X1 U10884 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9753) );
  AOI222_X1 U10885 ( .A1(n9764), .A2(n9754), .B1(n9753), .B2(n9752), .C1(n9751), .C2(n9750), .ZN(n9755) );
  OAI221_X1 U10886 ( .B1(n9757), .B2(n9762), .C1(n8268), .C2(n9756), .A(n9755), 
        .ZN(P2_U3230) );
  INV_X1 U10887 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9759) );
  AOI22_X1 U10888 ( .A1(n9819), .A2(n9759), .B1(n9758), .B2(n9817), .ZN(
        P2_U3393) );
  INV_X1 U10889 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U10890 ( .A1(n9819), .A2(n9761), .B1(n9760), .B2(n9817), .ZN(
        P2_U3396) );
  INV_X1 U10891 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9765) );
  OAI21_X1 U10892 ( .B1(n4522), .B2(n9793), .A(n9762), .ZN(n9763) );
  AOI21_X1 U10893 ( .B1(n9811), .B2(n9764), .A(n9763), .ZN(n9821) );
  AOI22_X1 U10894 ( .A1(n9819), .A2(n9765), .B1(n9821), .B2(n9817), .ZN(
        P2_U3399) );
  NOR2_X1 U10895 ( .A1(n9766), .A2(n9793), .ZN(n9768) );
  AOI211_X1 U10896 ( .C1(n9811), .C2(n9769), .A(n9768), .B(n9767), .ZN(n9823)
         );
  AOI22_X1 U10897 ( .A1(n9819), .A2(n5849), .B1(n9823), .B2(n9817), .ZN(
        P2_U3402) );
  INV_X1 U10898 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9962) );
  INV_X1 U10899 ( .A(n9770), .ZN(n9774) );
  OAI21_X1 U10900 ( .B1(n9772), .B2(n9793), .A(n9771), .ZN(n9773) );
  AOI21_X1 U10901 ( .B1(n9774), .B2(n9811), .A(n9773), .ZN(n9825) );
  AOI22_X1 U10902 ( .A1(n9819), .A2(n9962), .B1(n9825), .B2(n9817), .ZN(
        P2_U3405) );
  INV_X1 U10903 ( .A(n9775), .ZN(n9779) );
  OAI22_X1 U10904 ( .A1(n9777), .A2(n9804), .B1(n9776), .B2(n9793), .ZN(n9778)
         );
  NOR2_X1 U10905 ( .A1(n9779), .A2(n9778), .ZN(n9827) );
  AOI22_X1 U10906 ( .A1(n9819), .A2(n5872), .B1(n9827), .B2(n9817), .ZN(
        P2_U3408) );
  INV_X1 U10907 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9787) );
  INV_X1 U10908 ( .A(n9785), .ZN(n9781) );
  OAI22_X1 U10909 ( .A1(n9781), .A2(n9798), .B1(n9780), .B2(n9793), .ZN(n9784)
         );
  INV_X1 U10910 ( .A(n9782), .ZN(n9783) );
  AOI211_X1 U10911 ( .C1(n9786), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9828)
         );
  AOI22_X1 U10912 ( .A1(n9819), .A2(n9787), .B1(n9828), .B2(n9817), .ZN(
        P2_U3411) );
  INV_X1 U10913 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9976) );
  INV_X1 U10914 ( .A(n9788), .ZN(n9792) );
  OAI22_X1 U10915 ( .A1(n9790), .A2(n9804), .B1(n9789), .B2(n9793), .ZN(n9791)
         );
  NOR2_X1 U10916 ( .A1(n9792), .A2(n9791), .ZN(n9829) );
  AOI22_X1 U10917 ( .A1(n9819), .A2(n9976), .B1(n9829), .B2(n9817), .ZN(
        P2_U3414) );
  OAI22_X1 U10918 ( .A1(n9795), .A2(n9798), .B1(n9794), .B2(n9793), .ZN(n9796)
         );
  NOR2_X1 U10919 ( .A1(n9797), .A2(n9796), .ZN(n9830) );
  AOI22_X1 U10920 ( .A1(n9819), .A2(n5910), .B1(n9830), .B2(n9817), .ZN(
        P2_U3417) );
  INV_X1 U10921 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9803) );
  NOR2_X1 U10922 ( .A1(n9799), .A2(n9798), .ZN(n9801) );
  AOI211_X1 U10923 ( .C1(n9816), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9831)
         );
  AOI22_X1 U10924 ( .A1(n9819), .A2(n9803), .B1(n9831), .B2(n9817), .ZN(
        P2_U3420) );
  INV_X1 U10925 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U10926 ( .A1(n9805), .A2(n9804), .ZN(n9807) );
  AOI211_X1 U10927 ( .C1(n9816), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9832)
         );
  AOI22_X1 U10928 ( .A1(n9819), .A2(n9809), .B1(n9832), .B2(n9817), .ZN(
        P2_U3423) );
  INV_X1 U10929 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9818) );
  AND3_X1 U10930 ( .A1(n9812), .A2(n9811), .A3(n9810), .ZN(n9814) );
  AOI211_X1 U10931 ( .C1(n9816), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9834)
         );
  AOI22_X1 U10932 ( .A1(n9819), .A2(n9818), .B1(n9834), .B2(n9817), .ZN(
        P2_U3426) );
  INV_X1 U10933 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9820) );
  AOI22_X1 U10934 ( .A1(n4275), .A2(n9821), .B1(n9820), .B2(n9833), .ZN(
        P2_U3462) );
  AOI22_X1 U10935 ( .A1(n4275), .A2(n9823), .B1(n9822), .B2(n9833), .ZN(
        P2_U3463) );
  INV_X1 U10936 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U10937 ( .A1(n4275), .A2(n9825), .B1(n9824), .B2(n9833), .ZN(
        P2_U3464) );
  AOI22_X1 U10938 ( .A1(n4275), .A2(n9827), .B1(n9826), .B2(n9833), .ZN(
        P2_U3465) );
  AOI22_X1 U10939 ( .A1(n4275), .A2(n9828), .B1(n6748), .B2(n9833), .ZN(
        P2_U3466) );
  AOI22_X1 U10940 ( .A1(n4275), .A2(n9829), .B1(n6764), .B2(n9833), .ZN(
        P2_U3467) );
  AOI22_X1 U10941 ( .A1(n4275), .A2(n9830), .B1(n6834), .B2(n9833), .ZN(
        P2_U3468) );
  AOI22_X1 U10942 ( .A1(n4275), .A2(n9831), .B1(n7040), .B2(n9833), .ZN(
        P2_U3469) );
  AOI22_X1 U10943 ( .A1(n4275), .A2(n9832), .B1(n7069), .B2(n9833), .ZN(
        P2_U3470) );
  AOI22_X1 U10944 ( .A1(n4275), .A2(n9834), .B1(n7227), .B2(n9833), .ZN(
        P2_U3471) );
  OAI222_X1 U10945 ( .A1(n9839), .A2(n9838), .B1(n9839), .B2(n9837), .C1(n9836), .C2(n9835), .ZN(ADD_1068_U5) );
  XOR2_X1 U10946 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U10947 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9843) );
  XOR2_X1 U10948 ( .A(n9843), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55) );
  OAI21_X1 U10949 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(ADD_1068_U56) );
  OAI21_X1 U10950 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(ADD_1068_U57) );
  OAI21_X1 U10951 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(ADD_1068_U58) );
  OAI21_X1 U10952 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(ADD_1068_U59) );
  OAI21_X1 U10953 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(ADD_1068_U60) );
  OAI21_X1 U10954 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(ADD_1068_U61) );
  OAI21_X1 U10955 ( .B1(n9864), .B2(n9863), .A(n9862), .ZN(ADD_1068_U62) );
  OAI21_X1 U10956 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(ADD_1068_U63) );
  AOI21_X1 U10957 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9892) );
  INV_X1 U10958 ( .A(n9871), .ZN(n9883) );
  INV_X1 U10959 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9879) );
  AND3_X1 U10960 ( .A1(n9873), .A2(n9872), .A3(n4355), .ZN(n9875) );
  OAI21_X1 U10961 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9878) );
  OAI211_X1 U10962 ( .C1(n9880), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9881)
         );
  AOI21_X1 U10963 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9890) );
  OAI21_X1 U10964 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9888) );
  NAND2_X1 U10965 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  OAI211_X1 U10966 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9889), .ZN(n10041)
         );
  NOR4_X1 U10967 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(P2_REG1_REG_30__SCAN_IN), 
        .A3(P2_REG2_REG_26__SCAN_IN), .A4(P2_REG2_REG_15__SCAN_IN), .ZN(n9914)
         );
  NAND3_X1 U10968 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_DATAO_REG_29__SCAN_IN), 
        .A3(P1_DATAO_REG_24__SCAN_IN), .ZN(n9895) );
  NAND4_X1 U10969 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P1_DATAO_REG_29__SCAN_IN), .A3(P2_DATAO_REG_22__SCAN_IN), .A4(P2_DATAO_REG_13__SCAN_IN), .ZN(n9894) );
  NAND4_X1 U10970 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        SI_27_), .A4(P2_DATAO_REG_11__SCAN_IN), .ZN(n9893) );
  NOR4_X1 U10971 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9895), .A3(n9894), .A4(
        n9893), .ZN(n9913) );
  NAND4_X1 U10972 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .A3(P2_DATAO_REG_20__SCAN_IN), .A4(P2_REG0_REG_8__SCAN_IN), .ZN(n9899)
         );
  NAND4_X1 U10973 ( .A1(SI_21_), .A2(SI_19_), .A3(P1_IR_REG_29__SCAN_IN), .A4(
        P1_REG1_REG_22__SCAN_IN), .ZN(n9898) );
  NAND4_X1 U10974 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), 
        .A3(P1_REG3_REG_11__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n9897)
         );
  NAND4_X1 U10975 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P2_REG2_REG_22__SCAN_IN), .A3(P1_REG2_REG_23__SCAN_IN), .A4(P1_REG1_REG_16__SCAN_IN), .ZN(n9896) );
  NOR4_X1 U10976 ( .A1(n9899), .A2(n9898), .A3(n9897), .A4(n9896), .ZN(n9912)
         );
  NOR4_X1 U10977 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(P1_REG1_REG_29__SCAN_IN), .ZN(n9903)
         );
  NOR4_X1 U10978 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_REG3_REG_15__SCAN_IN), .A4(P1_REG0_REG_10__SCAN_IN), .ZN(n9902) );
  NOR4_X1 U10979 ( .A1(P1_RD_REG_SCAN_IN), .A2(P1_REG2_REG_3__SCAN_IN), .A3(
        P2_DATAO_REG_31__SCAN_IN), .A4(P1_ADDR_REG_12__SCAN_IN), .ZN(n9901) );
  NOR4_X1 U10980 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(P2_DATAO_REG_23__SCAN_IN), .A3(P1_DATAO_REG_23__SCAN_IN), .A4(P2_REG1_REG_17__SCAN_IN), .ZN(n9900) );
  NAND4_X1 U10981 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9910)
         );
  NOR4_X1 U10982 ( .A1(SI_15_), .A2(SI_1_), .A3(P1_DATAO_REG_0__SCAN_IN), .A4(
        P2_REG0_REG_5__SCAN_IN), .ZN(n9904) );
  NAND4_X1 U10983 ( .A1(n9905), .A2(P1_ADDR_REG_4__SCAN_IN), .A3(n9904), .A4(
        n9916), .ZN(n9909) );
  NAND4_X1 U10984 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n10007), .A3(n10024), 
        .A4(n9991), .ZN(n9906) );
  NOR3_X1 U10985 ( .A1(SI_20_), .A2(P2_REG0_REG_21__SCAN_IN), .A3(n9906), .ZN(
        n9907) );
  NAND3_X1 U10986 ( .A1(n9907), .A2(n9937), .A3(n9992), .ZN(n9908) );
  NOR3_X1 U10987 ( .A1(n9910), .A2(n9909), .A3(n9908), .ZN(n9911) );
  NAND4_X1 U10988 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n10039) );
  AOI22_X1 U10989 ( .A1(n8618), .A2(keyinput21), .B1(keyinput58), .B2(n9916), 
        .ZN(n9915) );
  OAI221_X1 U10990 ( .B1(n8618), .B2(keyinput21), .C1(n9916), .C2(keyinput58), 
        .A(n9915), .ZN(n9926) );
  AOI22_X1 U10991 ( .A1(n6764), .A2(keyinput45), .B1(keyinput61), .B2(n9918), 
        .ZN(n9917) );
  OAI221_X1 U10992 ( .B1(n6764), .B2(keyinput45), .C1(n9918), .C2(keyinput61), 
        .A(n9917), .ZN(n9925) );
  AOI22_X1 U10993 ( .A1(n6412), .A2(keyinput28), .B1(n9920), .B2(keyinput12), 
        .ZN(n9919) );
  OAI221_X1 U10994 ( .B1(n6412), .B2(keyinput28), .C1(n9920), .C2(keyinput12), 
        .A(n9919), .ZN(n9924) );
  XOR2_X1 U10995 ( .A(n7070), .B(keyinput33), .Z(n9922) );
  XNOR2_X1 U10996 ( .A(SI_1_), .B(keyinput14), .ZN(n9921) );
  NAND2_X1 U10997 ( .A1(n9922), .A2(n9921), .ZN(n9923) );
  NOR4_X1 U10998 ( .A1(n9926), .A2(n9925), .A3(n9924), .A4(n9923), .ZN(n9973)
         );
  AOI22_X1 U10999 ( .A1(n8107), .A2(keyinput25), .B1(n9928), .B2(keyinput23), 
        .ZN(n9927) );
  OAI221_X1 U11000 ( .B1(n8107), .B2(keyinput25), .C1(n9928), .C2(keyinput23), 
        .A(n9927), .ZN(n9941) );
  AOI22_X1 U11001 ( .A1(n9931), .A2(keyinput8), .B1(keyinput10), .B2(n9930), 
        .ZN(n9929) );
  OAI221_X1 U11002 ( .B1(n9931), .B2(keyinput8), .C1(n9930), .C2(keyinput10), 
        .A(n9929), .ZN(n9940) );
  AOI22_X1 U11003 ( .A1(n9934), .A2(keyinput24), .B1(n9933), .B2(keyinput2), 
        .ZN(n9932) );
  OAI221_X1 U11004 ( .B1(n9934), .B2(keyinput24), .C1(n9933), .C2(keyinput2), 
        .A(n9932), .ZN(n9939) );
  AOI22_X1 U11005 ( .A1(n9937), .A2(keyinput20), .B1(n9936), .B2(keyinput49), 
        .ZN(n9935) );
  OAI221_X1 U11006 ( .B1(n9937), .B2(keyinput20), .C1(n9936), .C2(keyinput49), 
        .A(n9935), .ZN(n9938) );
  NOR4_X1 U11007 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9972)
         );
  AOI22_X1 U11008 ( .A1(n9943), .A2(keyinput16), .B1(n6001), .B2(keyinput37), 
        .ZN(n9942) );
  OAI221_X1 U11009 ( .B1(n9943), .B2(keyinput16), .C1(n6001), .C2(keyinput37), 
        .A(n9942), .ZN(n9954) );
  AOI22_X1 U11010 ( .A1(n9946), .A2(keyinput1), .B1(keyinput41), .B2(n9945), 
        .ZN(n9944) );
  OAI221_X1 U11011 ( .B1(n9946), .B2(keyinput1), .C1(n9945), .C2(keyinput41), 
        .A(n9944), .ZN(n9953) );
  AOI22_X1 U11012 ( .A1(n8128), .A2(keyinput32), .B1(n9948), .B2(keyinput3), 
        .ZN(n9947) );
  OAI221_X1 U11013 ( .B1(n8128), .B2(keyinput32), .C1(n9948), .C2(keyinput3), 
        .A(n9947), .ZN(n9952) );
  XNOR2_X1 U11014 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput35), .ZN(n9950) );
  XNOR2_X1 U11015 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput27), .ZN(n9949) );
  NAND2_X1 U11016 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  NOR4_X1 U11017 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n9971)
         );
  AOI22_X1 U11018 ( .A1(n9957), .A2(keyinput26), .B1(keyinput36), .B2(n9956), 
        .ZN(n9955) );
  OAI221_X1 U11019 ( .B1(n9957), .B2(keyinput26), .C1(n9956), .C2(keyinput36), 
        .A(n9955), .ZN(n9969) );
  AOI22_X1 U11020 ( .A1(n9960), .A2(keyinput51), .B1(n9959), .B2(keyinput34), 
        .ZN(n9958) );
  OAI221_X1 U11021 ( .B1(n9960), .B2(keyinput51), .C1(n9959), .C2(keyinput34), 
        .A(n9958), .ZN(n9968) );
  AOI22_X1 U11022 ( .A1(n9963), .A2(keyinput53), .B1(keyinput19), .B2(n9962), 
        .ZN(n9961) );
  OAI221_X1 U11023 ( .B1(n9963), .B2(keyinput53), .C1(n9962), .C2(keyinput19), 
        .A(n9961), .ZN(n9967) );
  AOI22_X1 U11024 ( .A1(n9213), .A2(keyinput13), .B1(n9965), .B2(keyinput46), 
        .ZN(n9964) );
  OAI221_X1 U11025 ( .B1(n9213), .B2(keyinput13), .C1(n9965), .C2(keyinput46), 
        .A(n9964), .ZN(n9966) );
  NOR4_X1 U11026 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9970)
         );
  NAND4_X1 U11027 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n10037) );
  AOI22_X1 U11028 ( .A1(n9976), .A2(keyinput48), .B1(keyinput44), .B2(n9975), 
        .ZN(n9974) );
  OAI221_X1 U11029 ( .B1(n9976), .B2(keyinput48), .C1(n9975), .C2(keyinput44), 
        .A(n9974), .ZN(n9987) );
  AOI22_X1 U11030 ( .A1(n9979), .A2(keyinput11), .B1(n9978), .B2(keyinput30), 
        .ZN(n9977) );
  OAI221_X1 U11031 ( .B1(n9979), .B2(keyinput11), .C1(n9978), .C2(keyinput30), 
        .A(n9977), .ZN(n9986) );
  AOI22_X1 U11032 ( .A1(n7091), .A2(keyinput47), .B1(keyinput62), .B2(n5240), 
        .ZN(n9980) );
  OAI221_X1 U11033 ( .B1(n7091), .B2(keyinput47), .C1(n5240), .C2(keyinput62), 
        .A(n9980), .ZN(n9985) );
  AOI22_X1 U11034 ( .A1(n9983), .A2(keyinput57), .B1(n9982), .B2(keyinput42), 
        .ZN(n9981) );
  OAI221_X1 U11035 ( .B1(n9983), .B2(keyinput57), .C1(n9982), .C2(keyinput42), 
        .A(n9981), .ZN(n9984) );
  NOR4_X1 U11036 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n10035)
         );
  INV_X1 U11037 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U11038 ( .A1(n9990), .A2(keyinput17), .B1(n9989), .B2(keyinput0), 
        .ZN(n9988) );
  OAI221_X1 U11039 ( .B1(n9990), .B2(keyinput17), .C1(n9989), .C2(keyinput0), 
        .A(n9988), .ZN(n9995) );
  XNOR2_X1 U11040 ( .A(n9991), .B(keyinput52), .ZN(n9994) );
  XNOR2_X1 U11041 ( .A(n9992), .B(keyinput56), .ZN(n9993) );
  OR3_X1 U11042 ( .A1(n9995), .A2(n9994), .A3(n9993), .ZN(n10002) );
  AOI22_X1 U11043 ( .A1(n5072), .A2(keyinput22), .B1(keyinput29), .B2(n8054), 
        .ZN(n9996) );
  OAI221_X1 U11044 ( .B1(n5072), .B2(keyinput22), .C1(n8054), .C2(keyinput29), 
        .A(n9996), .ZN(n10001) );
  AOI22_X1 U11045 ( .A1(n9999), .A2(keyinput40), .B1(n9998), .B2(keyinput55), 
        .ZN(n9997) );
  OAI221_X1 U11046 ( .B1(n9999), .B2(keyinput40), .C1(n9998), .C2(keyinput55), 
        .A(n9997), .ZN(n10000) );
  NOR3_X1 U11047 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(n10034) );
  AOI22_X1 U11048 ( .A1(n10005), .A2(keyinput15), .B1(keyinput9), .B2(n10004), 
        .ZN(n10003) );
  OAI221_X1 U11049 ( .B1(n10005), .B2(keyinput15), .C1(n10004), .C2(keyinput9), 
        .A(n10003), .ZN(n10017) );
  AOI22_X1 U11050 ( .A1(n10008), .A2(keyinput59), .B1(n10007), .B2(keyinput18), 
        .ZN(n10006) );
  OAI221_X1 U11051 ( .B1(n10008), .B2(keyinput59), .C1(n10007), .C2(keyinput18), .A(n10006), .ZN(n10016) );
  INV_X1 U11052 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U11053 ( .A1(n10011), .A2(keyinput38), .B1(n10010), .B2(keyinput39), 
        .ZN(n10009) );
  OAI221_X1 U11054 ( .B1(n10011), .B2(keyinput38), .C1(n10010), .C2(keyinput39), .A(n10009), .ZN(n10015) );
  XOR2_X1 U11055 ( .A(n4579), .B(keyinput6), .Z(n10013) );
  XNOR2_X1 U11056 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput7), .ZN(n10012) );
  NAND2_X1 U11057 ( .A1(n10013), .A2(n10012), .ZN(n10014) );
  NOR4_X1 U11058 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n10033) );
  AOI22_X1 U11059 ( .A1(n10019), .A2(keyinput5), .B1(n5505), .B2(keyinput31), 
        .ZN(n10018) );
  OAI221_X1 U11060 ( .B1(n10019), .B2(keyinput5), .C1(n5505), .C2(keyinput31), 
        .A(n10018), .ZN(n10031) );
  INV_X1 U11061 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U11062 ( .A1(n10022), .A2(keyinput54), .B1(n10021), .B2(keyinput63), 
        .ZN(n10020) );
  OAI221_X1 U11063 ( .B1(n10022), .B2(keyinput54), .C1(n10021), .C2(keyinput63), .A(n10020), .ZN(n10030) );
  AOI22_X1 U11064 ( .A1(n10025), .A2(keyinput50), .B1(n10024), .B2(keyinput43), 
        .ZN(n10023) );
  OAI221_X1 U11065 ( .B1(n10025), .B2(keyinput50), .C1(n10024), .C2(keyinput43), .A(n10023), .ZN(n10029) );
  XNOR2_X1 U11066 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput60), .ZN(n10027)
         );
  XNOR2_X1 U11067 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput4), .ZN(n10026) );
  NAND2_X1 U11068 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NOR4_X1 U11069 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10032) );
  NAND4_X1 U11070 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10036) );
  NOR2_X1 U11071 ( .A1(n10037), .A2(n10036), .ZN(n10038) );
  XOR2_X1 U11072 ( .A(n10039), .B(n10038), .Z(n10040) );
  XNOR2_X1 U11073 ( .A(n10041), .B(n10040), .ZN(P2_U3188) );
  OAI21_X1 U11074 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(ADD_1068_U50) );
  OAI21_X1 U11075 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(ADD_1068_U51) );
  OAI21_X1 U11076 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(ADD_1068_U47) );
  OAI21_X1 U11077 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(ADD_1068_U49) );
  OAI21_X1 U11078 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(ADD_1068_U48) );
  AOI21_X1 U11079 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(ADD_1068_U54) );
  AOI21_X1 U11080 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(ADD_1068_U53) );
  OAI21_X1 U11081 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4935 ( .A(n6798), .Z(n4421) );
  CLKBUF_X1 U5118 ( .A(n8236), .Z(n4416) );
  CLKBUF_X2 U5220 ( .A(n5815), .Z(n4412) );
  CLKBUF_X1 U5336 ( .A(n5805), .Z(n6443) );
  AND4_X1 U5897 ( .A1(n4946), .A2(n4969), .A3(n4979), .A4(n5716), .ZN(n10068)
         );
endmodule

