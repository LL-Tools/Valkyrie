

module b14_C_AntiSAT_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727;

  OR2_X1 U2296 ( .A1(n2528), .A2(n3671), .ZN(n2537) );
  CLKBUF_X2 U2299 ( .A(n2275), .Z(n2609) );
  CLKBUF_X1 U2300 ( .A(n3757), .Z(n2054) );
  NOR2_X1 U2301 ( .A1(n2849), .A2(n4381), .ZN(n3757) );
  OR2_X1 U2302 ( .A1(n3529), .A2(n3528), .ZN(n3678) );
  INV_X1 U2303 ( .A(n2983), .ZN(n2286) );
  INV_X1 U2304 ( .A(n3597), .ZN(n3613) );
  NAND3_X1 U2305 ( .A1(n2742), .A2(n2734), .A3(n2739), .ZN(n2897) );
  INV_X1 U2306 ( .A(IR_REG_31__SCAN_IN), .ZN(n2754) );
  INV_X1 U2307 ( .A(n2634), .ZN(n3907) );
  NAND3_X1 U2309 ( .A1(n2226), .A2(n2281), .A3(n2280), .ZN(n2288) );
  NAND2_X1 U2310 ( .A1(n3280), .A2(n3259), .ZN(n3301) );
  XNOR2_X1 U2311 ( .A(n2259), .B(n2258), .ZN(n2723) );
  NAND2_X2 U2312 ( .A1(n4372), .A2(n2080), .ZN(n2200) );
  NAND2_X2 U2313 ( .A1(n3460), .A2(n2452), .ZN(n4372) );
  NAND2_X2 U2314 ( .A1(n4347), .A2(n2479), .ZN(n4304) );
  NAND2_X2 U2315 ( .A1(n2200), .A2(n2063), .ZN(n4347) );
  NAND2_X2 U2316 ( .A1(n3306), .A2(n3305), .ZN(n3342) );
  NAND2_X2 U2317 ( .A1(n2329), .A2(n2328), .ZN(n3074) );
  OAI21_X2 U2318 ( .B1(n3540), .B2(n2162), .A(n2159), .ZN(n3646) );
  NAND3_X2 U2319 ( .A1(n3535), .A2(n3534), .A3(n3533), .ZN(n3540) );
  XNOR2_X2 U2320 ( .A(n2566), .B(n2565), .ZN(n2634) );
  AND2_X1 U2321 ( .A1(n3678), .A2(n3677), .ZN(n3676) );
  CLKBUF_X1 U2322 ( .A(n2272), .Z(n2823) );
  NAND4_X1 U2323 ( .A1(n2308), .A2(n2307), .A3(n2306), .A4(n2305), .ZN(n3127)
         );
  NAND2_X2 U2324 ( .A1(n3911), .A2(n3907), .ZN(n3059) );
  CLKBUF_X3 U2325 ( .A(n2069), .Z(n3828) );
  AND2_X1 U2326 ( .A1(n2489), .A2(n2561), .ZN(n4362) );
  XNOR2_X1 U2327 ( .A(n2249), .B(IR_REG_29__SCAN_IN), .ZN(n2253) );
  NAND2_X1 U2328 ( .A1(n2115), .A2(n2614), .ZN(n2618) );
  AND2_X1 U2329 ( .A1(n2669), .A2(n2105), .ZN(n2674) );
  AND2_X1 U2330 ( .A1(n2195), .A2(n2076), .ZN(n4180) );
  NAND2_X1 U2331 ( .A1(n2366), .A2(n2365), .ZN(n3189) );
  AND2_X2 U2332 ( .A1(n2554), .A2(n2553), .ZN(n4404) );
  NAND2_X1 U2333 ( .A1(n4167), .A2(n2549), .ZN(n2554) );
  AND2_X1 U2334 ( .A1(n2548), .A2(n4157), .ZN(n4167) );
  BUF_X2 U2335 ( .A(n3344), .Z(n3544) );
  NAND2_X1 U2336 ( .A1(n3772), .A2(n3775), .ZN(n3864) );
  AND2_X2 U2337 ( .A1(n2897), .A2(n2696), .ZN(n2994) );
  NAND4_X2 U2338 ( .A1(n2295), .A2(n2294), .A3(n2293), .A4(n2292), .ZN(n3936)
         );
  INV_X1 U2339 ( .A(n4362), .ZN(n4146) );
  AND3_X1 U2340 ( .A1(n2124), .A2(n2126), .A3(n2064), .ZN(n2961) );
  MUX2_X1 U2341 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2056), .Z(n2867) );
  OR2_X1 U2342 ( .A1(n2810), .A2(n2127), .ZN(n2124) );
  NAND2_X1 U2343 ( .A1(n2251), .A2(n2250), .ZN(n2278) );
  NAND2_X1 U2344 ( .A1(n2561), .A2(IR_REG_31__SCAN_IN), .ZN(n2563) );
  AND2_X1 U2345 ( .A1(n2628), .A2(n2627), .ZN(n2734) );
  NAND2_X1 U2346 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  BUF_X1 U2347 ( .A(n2253), .Z(n2752) );
  OR2_X1 U2348 ( .A1(n2564), .A2(IR_REG_21__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U2349 ( .A1(n2627), .A2(n2262), .ZN(n2664) );
  NAND2_X1 U2350 ( .A1(n2228), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  OR2_X1 U2351 ( .A1(n2572), .A2(n2754), .ZN(n2249) );
  AND2_X1 U2352 ( .A1(n2621), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  AND2_X1 U2353 ( .A1(n2382), .A2(REG3_REG_10__SCAN_IN), .ZN(n2390) );
  AND2_X1 U2354 ( .A1(n2062), .A2(n2107), .ZN(n2106) );
  AND2_X1 U2355 ( .A1(n2207), .A2(n2247), .ZN(n2062) );
  AND2_X1 U2356 ( .A1(n2243), .A2(n2557), .ZN(n2620) );
  AND2_X1 U2357 ( .A1(n2622), .A2(n2244), .ZN(n2245) );
  OR2_X1 U2358 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2475)
         );
  OR2_X1 U2359 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2242)
         );
  NOR2_X1 U2360 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2231)
         );
  NOR2_X1 U2361 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2233)
         );
  NOR2_X1 U2362 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2234)
         );
  INV_X1 U2363 ( .A(IR_REG_3__SCAN_IN), .ZN(n2309) );
  INV_X1 U2364 ( .A(IR_REG_4__SCAN_IN), .ZN(n2312) );
  NOR2_X1 U2365 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2232)
         );
  INV_X1 U2366 ( .A(IR_REG_14__SCAN_IN), .ZN(n2240) );
  INV_X1 U2367 ( .A(IR_REG_2__SCAN_IN), .ZN(n2283) );
  AND4_X2 U2368 ( .A1(n2234), .A2(n2233), .A3(n2232), .A4(n2231), .ZN(n2420)
         );
  AOI21_X2 U2369 ( .B1(n3174), .B2(n2182), .A(n2179), .ZN(n3217) );
  NAND2_X2 U2370 ( .A1(n2577), .A2(n3764), .ZN(n2575) );
  OAI211_X2 U2371 ( .C1(n3629), .C2(n2609), .A(n2545), .B(n2544), .ZN(n4200)
         );
  MUX2_X1 U2372 ( .A(n2665), .B(n2664), .S(IR_REG_28__SCAN_IN), .Z(n2056) );
  OAI22_X1 U2373 ( .A1(n2655), .A2(n3851), .B1(n4404), .B2(n4170), .ZN(n2656)
         );
  NAND2_X2 U2374 ( .A1(n2265), .A2(n2264), .ZN(n2577) );
  AOI22_X2 U2375 ( .A1(n2823), .A2(n2057), .B1(n2994), .B2(n2264), .ZN(n2904)
         );
  INV_X2 U2376 ( .A(n3161), .ZN(n2264) );
  AND2_X1 U2377 ( .A1(n3610), .A2(n3085), .ZN(n2057) );
  AND2_X1 U2378 ( .A1(n3610), .A2(n3085), .ZN(n2058) );
  AND2_X1 U2379 ( .A1(n3610), .A2(n3085), .ZN(n3344) );
  NAND2_X1 U2380 ( .A1(n2251), .A2(n2250), .ZN(n2059) );
  AOI22_X2 U2381 ( .A1(n4234), .A2(n2527), .B1(n4255), .B2(n4241), .ZN(n4211)
         );
  AOI21_X2 U2382 ( .B1(n4247), .B2(n2520), .A(n2081), .ZN(n4234) );
  INV_X1 U2383 ( .A(IR_REG_23__SCAN_IN), .ZN(n2622) );
  NOR2_X1 U2384 ( .A1(n2776), .A2(n2074), .ZN(n2787) );
  OR2_X1 U2385 ( .A1(n3318), .A2(n3291), .ZN(n2204) );
  NAND2_X1 U2386 ( .A1(n2821), .A2(n2634), .ZN(n2833) );
  NOR2_X1 U2387 ( .A1(n3627), .A2(n2174), .ZN(n2173) );
  XNOR2_X1 U2388 ( .A(n2787), .B(n2211), .ZN(n2777) );
  OR2_X1 U2389 ( .A1(n2777), .A2(n2778), .ZN(n2210) );
  AOI21_X1 U2390 ( .B1(n2785), .B2(REG2_REG_3__SCAN_IN), .A(n2133), .ZN(n2811)
         );
  AND2_X1 U2391 ( .A1(n2134), .A2(n2790), .ZN(n2133) );
  NAND2_X1 U2392 ( .A1(n4582), .A2(n4583), .ZN(n4581) );
  XNOR2_X1 U2393 ( .A(n3498), .B(n2123), .ZN(n4594) );
  NAND2_X1 U2394 ( .A1(n3324), .A2(n2411), .ZN(n2413) );
  NAND2_X1 U2395 ( .A1(n2488), .A2(n2487), .ZN(n2561) );
  INV_X1 U2396 ( .A(IR_REG_19__SCAN_IN), .ZN(n2487) );
  OR2_X1 U2397 ( .A1(n2833), .A2(n3911), .ZN(n4331) );
  INV_X1 U2398 ( .A(IR_REG_24__SCAN_IN), .ZN(n2244) );
  OAI22_X1 U2399 ( .A1(n2667), .A2(n4336), .B1(n3836), .B2(n4152), .ZN(n4160)
         );
  INV_X1 U2400 ( .A(IR_REG_16__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2401 ( .A1(n3420), .A2(n2158), .ZN(n2156) );
  NOR2_X1 U2402 ( .A1(n2158), .A2(n3420), .ZN(n2157) );
  OR2_X1 U2403 ( .A1(n2821), .A2(n4362), .ZN(n2841) );
  OR2_X1 U2404 ( .A1(n4436), .A2(n4282), .ZN(n4251) );
  AND2_X1 U2405 ( .A1(n4300), .A2(n2597), .ZN(n3888) );
  NOR2_X1 U2406 ( .A1(n3807), .A2(n2102), .ZN(n2101) );
  OR2_X1 U2407 ( .A1(n3936), .A2(n3094), .ZN(n3771) );
  NOR2_X1 U2408 ( .A1(n4203), .A2(n2534), .ZN(n2112) );
  NOR2_X1 U2409 ( .A1(n2109), .A2(n4474), .ZN(n2108) );
  INV_X1 U2410 ( .A(n2110), .ZN(n2109) );
  AND2_X1 U2411 ( .A1(n3069), .A2(n3068), .ZN(n3022) );
  NAND2_X1 U2412 ( .A1(n2246), .A2(n2260), .ZN(n2208) );
  AOI21_X1 U2413 ( .B1(n2157), .B2(n2156), .A(n2154), .ZN(n2153) );
  INV_X1 U2414 ( .A(n3433), .ZN(n2154) );
  NAND2_X1 U2415 ( .A1(n3215), .A2(n3216), .ZN(n2182) );
  NAND2_X1 U2416 ( .A1(n2181), .A2(n2180), .ZN(n2179) );
  NAND2_X1 U2417 ( .A1(n3149), .A2(n2185), .ZN(n2180) );
  AND2_X1 U2418 ( .A1(n3576), .A2(n3575), .ZN(n3707) );
  INV_X1 U2419 ( .A(n2156), .ZN(n2155) );
  INV_X1 U2420 ( .A(n2157), .ZN(n2152) );
  NAND2_X1 U2421 ( .A1(n3302), .A2(n3304), .ZN(n3305) );
  INV_X1 U2422 ( .A(n3303), .ZN(n3304) );
  NOR2_X2 U2423 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2282)
         );
  NAND2_X1 U2424 ( .A1(n2812), .A2(n2813), .ZN(n2131) );
  NAND2_X1 U2425 ( .A1(n2128), .A2(REG2_REG_4__SCAN_IN), .ZN(n2127) );
  INV_X1 U2426 ( .A(n2814), .ZN(n2128) );
  OR2_X1 U2427 ( .A1(n2131), .A2(n2814), .ZN(n2126) );
  AND2_X1 U2428 ( .A1(n2210), .A2(n2209), .ZN(n2805) );
  NAND2_X1 U2429 ( .A1(n2789), .A2(n2790), .ZN(n2209) );
  OR2_X1 U2430 ( .A1(n2809), .A2(n2808), .ZN(n2217) );
  INV_X1 U2431 ( .A(n3006), .ZN(n2212) );
  NAND2_X1 U2432 ( .A1(n4562), .A2(n3494), .ZN(n3495) );
  NAND2_X1 U2433 ( .A1(n4572), .A2(n3479), .ZN(n4582) );
  NAND2_X1 U2434 ( .A1(n4598), .A2(n3482), .ZN(n3485) );
  NAND2_X1 U2435 ( .A1(n3485), .A2(n3484), .ZN(n4128) );
  NAND2_X1 U2436 ( .A1(n4584), .A2(n3497), .ZN(n3498) );
  NAND2_X1 U2437 ( .A1(n4594), .A2(REG2_REG_12__SCAN_IN), .ZN(n4593) );
  OAI22_X1 U2438 ( .A1(n4117), .A2(n4116), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4115), .ZN(n4118) );
  NOR2_X1 U2439 ( .A1(n4612), .A2(n2122), .ZN(n4121) );
  AND2_X1 U2440 ( .A1(n4126), .A2(REG2_REG_15__SCAN_IN), .ZN(n2122) );
  NAND2_X1 U2441 ( .A1(n4637), .A2(n2142), .ZN(n2141) );
  OR2_X1 U2442 ( .A1(n4138), .A2(REG2_REG_17__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2443 ( .A1(n2220), .A2(n2224), .ZN(n2221) );
  AND2_X1 U2444 ( .A1(n2194), .A2(n2536), .ZN(n2189) );
  NAND2_X1 U2445 ( .A1(n2187), .A2(n2071), .ZN(n2186) );
  NOR2_X1 U2446 ( .A1(n2535), .A2(n2192), .ZN(n2191) );
  INV_X1 U2447 ( .A(n3848), .ZN(n2192) );
  AND2_X1 U2448 ( .A1(n4181), .A2(n3820), .ZN(n2099) );
  NAND2_X1 U2449 ( .A1(n4194), .A2(n3815), .ZN(n2100) );
  NAND2_X1 U2450 ( .A1(n4268), .A2(n2513), .ZN(n4247) );
  INV_X1 U2451 ( .A(n4354), .ZN(n2478) );
  NAND2_X1 U2452 ( .A1(n2091), .A2(n2090), .ZN(n2593) );
  AOI21_X1 U2453 ( .B1(n2093), .B2(n2095), .A(n2083), .ZN(n2090) );
  AND2_X1 U2454 ( .A1(n3397), .A2(n2078), .ZN(n2198) );
  AOI21_X1 U2455 ( .B1(n2203), .B2(n2389), .A(n2072), .ZN(n2202) );
  NAND2_X1 U2456 ( .A1(n2390), .A2(REG3_REG_11__SCAN_IN), .ZN(n2401) );
  AND2_X1 U2457 ( .A1(n3865), .A2(n2204), .ZN(n2203) );
  OR2_X1 U2458 ( .A1(n3257), .A2(n2389), .ZN(n2205) );
  NAND2_X1 U2459 ( .A1(n2205), .A2(n2204), .ZN(n3272) );
  OAI21_X1 U2460 ( .B1(n3195), .B2(n3785), .A(n3781), .ZN(n3266) );
  NAND2_X1 U2461 ( .A1(n2580), .A2(n3788), .ZN(n3075) );
  OR2_X1 U2462 ( .A1(n3018), .A2(n3016), .ZN(n2580) );
  AND2_X1 U2463 ( .A1(n2607), .A2(n2606), .ZN(n4336) );
  OR2_X1 U2464 ( .A1(n2275), .A2(n2274), .ZN(n2277) );
  OR2_X1 U2465 ( .A1(n2834), .A2(n2835), .ZN(n3055) );
  INV_X1 U2466 ( .A(n4336), .ZN(n4370) );
  NAND2_X1 U2467 ( .A1(n2672), .A2(n4163), .ZN(n4394) );
  NOR2_X1 U2468 ( .A1(n2113), .A2(n3619), .ZN(n2672) );
  NOR2_X1 U2469 ( .A1(n4338), .A2(n4444), .ZN(n4309) );
  AND2_X1 U2470 ( .A1(n3470), .A2(n3469), .ZN(n4376) );
  INV_X1 U2471 ( .A(n2631), .ZN(n2623) );
  AOI21_X1 U2472 ( .B1(n2163), .B2(n2161), .A(n2160), .ZN(n2159) );
  INV_X1 U2473 ( .A(n2163), .ZN(n2162) );
  INV_X1 U2474 ( .A(n3728), .ZN(n2160) );
  NOR2_X1 U2475 ( .A1(n3738), .A2(n2177), .ZN(n2176) );
  INV_X1 U2476 ( .A(n3666), .ZN(n2177) );
  NAND2_X1 U2477 ( .A1(n3626), .A2(n2171), .ZN(n2170) );
  NAND2_X1 U2478 ( .A1(n2172), .A2(n2230), .ZN(n2171) );
  INV_X1 U2479 ( .A(n2173), .ZN(n2172) );
  INV_X1 U2480 ( .A(n4279), .ZN(n4421) );
  OAI211_X1 U2481 ( .C1(n3740), .C2(n2609), .A(n2541), .B(n2540), .ZN(n4401)
         );
  NAND4_X1 U2482 ( .A1(n2448), .A2(n2447), .A3(n2446), .A4(n2445), .ZN(n4378)
         );
  NAND4_X1 U2483 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .ZN(n3927)
         );
  XNOR2_X1 U2484 ( .A(n3495), .B(n2121), .ZN(n4575) );
  NAND2_X1 U2485 ( .A1(n4575), .A2(REG2_REG_10__SCAN_IN), .ZN(n4574) );
  XNOR2_X1 U2486 ( .A(n4121), .B(n4134), .ZN(n4624) );
  NAND2_X1 U2487 ( .A1(n4624), .A2(n4623), .ZN(n4622) );
  INV_X1 U2488 ( .A(n2221), .ZN(n4643) );
  INV_X1 U2489 ( .A(n2140), .ZN(n2139) );
  AOI21_X1 U2490 ( .B1(n2141), .B2(n4648), .A(n4646), .ZN(n2140) );
  AOI21_X1 U2491 ( .B1(n4650), .B2(ADDR_REG_18__SCAN_IN), .A(n4649), .ZN(n2138) );
  NOR2_X1 U2492 ( .A1(n2141), .A2(n4648), .ZN(n4647) );
  NOR2_X1 U2493 ( .A1(n4643), .A2(n4139), .ZN(n4653) );
  NAND2_X1 U2494 ( .A1(n2221), .A2(n2222), .ZN(n4651) );
  NAND2_X1 U2495 ( .A1(n4162), .A2(n2118), .ZN(n2117) );
  NAND2_X1 U2496 ( .A1(n3334), .A2(n2119), .ZN(n2118) );
  INV_X1 U2497 ( .A(n4163), .ZN(n2119) );
  NAND2_X1 U2498 ( .A1(n2848), .A2(n2847), .ZN(n4658) );
  AND2_X1 U2499 ( .A1(n4365), .A2(n3101), .ZN(n4374) );
  AOI21_X1 U2500 ( .B1(n4164), .B2(n4713), .A(n2668), .ZN(n2105) );
  OAI21_X1 U2501 ( .B1(n2672), .B2(n4163), .A(n4394), .ZN(n4158) );
  AND2_X1 U2502 ( .A1(n2649), .A2(n2648), .ZN(n2760) );
  INV_X1 U2503 ( .A(IR_REG_29__SCAN_IN), .ZN(n2107) );
  INV_X1 U2504 ( .A(n4125), .ZN(n4686) );
  NAND2_X1 U2505 ( .A1(n2183), .A2(n2184), .ZN(n2181) );
  OR2_X1 U2506 ( .A1(n3149), .A2(n2185), .ZN(n2183) );
  OR4_X1 U2507 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3903) );
  AND2_X1 U2508 ( .A1(n4229), .A2(n3847), .ZN(n3894) );
  OR2_X1 U2509 ( .A1(n2059), .A2(n2252), .ZN(n2257) );
  NAND2_X1 U2510 ( .A1(n2886), .A2(REG1_REG_5__SCAN_IN), .ZN(n2216) );
  AND2_X1 U2511 ( .A1(n2546), .A2(n2076), .ZN(n2194) );
  NAND2_X1 U2512 ( .A1(n2194), .A2(n2188), .ZN(n2187) );
  INV_X1 U2513 ( .A(n2191), .ZN(n2188) );
  INV_X1 U2514 ( .A(n2094), .ZN(n2093) );
  OAI21_X1 U2515 ( .B1(n3799), .B2(n2095), .A(n3872), .ZN(n2094) );
  NOR2_X1 U2516 ( .A1(n3347), .A2(n3413), .ZN(n2110) );
  AND2_X1 U2517 ( .A1(n3144), .A2(n3083), .ZN(n2114) );
  AND2_X1 U2518 ( .A1(n2462), .A2(n2241), .ZN(n2243) );
  AND2_X1 U2519 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2262)
         );
  INV_X1 U2520 ( .A(IR_REG_6__SCAN_IN), .ZN(n2347) );
  NOR2_X1 U2521 ( .A1(n3727), .A2(n2164), .ZN(n2163) );
  INV_X1 U2522 ( .A(n3549), .ZN(n2164) );
  INV_X1 U2523 ( .A(n2166), .ZN(n2161) );
  INV_X1 U2524 ( .A(n3130), .ZN(n3001) );
  OR2_X1 U2525 ( .A1(n3527), .A2(n3526), .ZN(n3535) );
  XNOR2_X1 U2526 ( .A(n2919), .B(n3597), .ZN(n2920) );
  INV_X1 U2527 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2528 ( .A1(n3540), .A2(n2166), .ZN(n2165) );
  OR2_X1 U2529 ( .A1(n2543), .A2(n2547), .ZN(n3629) );
  OR2_X1 U2530 ( .A1(n2609), .A2(n4274), .ZN(n2508) );
  OR2_X1 U2531 ( .A1(n2278), .A2(n2267), .ZN(n2268) );
  NOR3_X1 U2532 ( .A1(n2690), .A2(n2689), .A3(n4699), .ZN(n2711) );
  NAND2_X1 U2533 ( .A1(n2136), .A2(n2709), .ZN(n2774) );
  OR2_X1 U2534 ( .A1(n2711), .A2(n2710), .ZN(n2136) );
  NAND2_X1 U2535 ( .A1(n2774), .A2(n2135), .ZN(n2134) );
  NAND2_X1 U2536 ( .A1(n4552), .A2(REG2_REG_2__SCAN_IN), .ZN(n2135) );
  XNOR2_X1 U2537 ( .A(n2215), .B(n4551), .ZN(n2887) );
  OAI21_X1 U2538 ( .B1(n3476), .B2(n3475), .A(n2213), .ZN(n4561) );
  NAND2_X1 U2539 ( .A1(n4581), .A2(n3480), .ZN(n3481) );
  CLKBUF_X1 U2540 ( .A(n2322), .Z(n2323) );
  NAND2_X1 U2541 ( .A1(n4128), .A2(n4129), .ZN(n4131) );
  AND2_X1 U2542 ( .A1(n4654), .A2(n2223), .ZN(n2222) );
  INV_X1 U2543 ( .A(n4139), .ZN(n2223) );
  INV_X1 U2544 ( .A(n2222), .ZN(n2219) );
  AOI21_X1 U2545 ( .B1(n2099), .B2(n3897), .A(n2097), .ZN(n2096) );
  INV_X1 U2546 ( .A(n2099), .ZN(n2098) );
  INV_X1 U2547 ( .A(n3825), .ZN(n2097) );
  AND2_X1 U2548 ( .A1(n3826), .A2(n3819), .ZN(n3851) );
  AND2_X1 U2549 ( .A1(n4277), .A2(n2502), .ZN(n2206) );
  AND2_X1 U2550 ( .A1(n4250), .A2(n4249), .ZN(n4278) );
  NAND2_X1 U2551 ( .A1(n2103), .A2(n2066), .ZN(n4301) );
  AND2_X1 U2552 ( .A1(n2480), .A2(REG3_REG_19__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U2553 ( .A1(n2103), .A2(n2101), .ZN(n4325) );
  OR2_X1 U2554 ( .A1(n2456), .A2(n2455), .ZN(n2466) );
  NOR2_X1 U2555 ( .A1(n2466), .A2(n3732), .ZN(n2480) );
  NAND2_X1 U2556 ( .A1(n2436), .A2(REG3_REG_15__SCAN_IN), .ZN(n2456) );
  AOI21_X1 U2557 ( .B1(n2198), .B2(n2427), .A(n2061), .ZN(n2197) );
  NAND2_X1 U2558 ( .A1(n2092), .A2(n3802), .ZN(n3881) );
  NAND2_X1 U2559 ( .A1(n3325), .A2(n3799), .ZN(n2092) );
  OAI21_X1 U2560 ( .B1(n3325), .B2(n2095), .A(n2093), .ZN(n3444) );
  INV_X1 U2561 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3426) );
  OR2_X1 U2562 ( .A1(n2414), .A2(n3426), .ZN(n2429) );
  NAND2_X1 U2563 ( .A1(n2585), .A2(n3797), .ZN(n3325) );
  NAND2_X1 U2564 ( .A1(n3266), .A2(n3798), .ZN(n2585) );
  NAND2_X1 U2565 ( .A1(n2584), .A2(n3791), .ZN(n3195) );
  NAND2_X1 U2566 ( .A1(n2581), .A2(n3777), .ZN(n3114) );
  NAND2_X1 U2567 ( .A1(n3084), .A2(n3083), .ZN(n3112) );
  NOR2_X1 U2568 ( .A1(n2330), .A2(n2883), .ZN(n2339) );
  INV_X1 U2569 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2883) );
  OAI21_X1 U2570 ( .B1(n3061), .B2(n2579), .A(n3775), .ZN(n3018) );
  AND2_X1 U2571 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2317) );
  NAND2_X1 U2572 ( .A1(n2976), .A2(n3771), .ZN(n3061) );
  INV_X1 U2573 ( .A(n2575), .ZN(n2862) );
  NOR2_X1 U2574 ( .A1(n4394), .A2(n4396), .ZN(n4393) );
  AND2_X1 U2575 ( .A1(n2112), .A2(n4186), .ZN(n2111) );
  INV_X1 U2576 ( .A(n4197), .ZN(n4203) );
  NAND2_X1 U2577 ( .A1(n4236), .A2(n2112), .ZN(n4205) );
  NAND2_X1 U2578 ( .A1(n4236), .A2(n4221), .ZN(n4223) );
  AND2_X1 U2579 ( .A1(n4260), .A2(n4241), .ZN(n4236) );
  INV_X1 U2580 ( .A(n4254), .ZN(n4259) );
  NOR2_X1 U2581 ( .A1(n4273), .A2(n4259), .ZN(n4260) );
  OR2_X1 U2582 ( .A1(n4291), .A2(n2512), .ZN(n4273) );
  NAND2_X1 U2583 ( .A1(n4309), .A2(n4295), .ZN(n4291) );
  INV_X1 U2584 ( .A(n4316), .ZN(n4444) );
  NAND2_X1 U2585 ( .A1(n4376), .A2(n2086), .ZN(n4338) );
  NAND2_X1 U2586 ( .A1(n4376), .A2(n2068), .ZN(n4350) );
  NAND2_X1 U2587 ( .A1(n4376), .A2(n4386), .ZN(n4375) );
  AND2_X1 U2588 ( .A1(n3330), .A2(n2067), .ZN(n3470) );
  NAND2_X1 U2589 ( .A1(n3330), .A2(n2108), .ZN(n3449) );
  NAND2_X1 U2590 ( .A1(n3330), .A2(n2110), .ZN(n3401) );
  AND2_X1 U2591 ( .A1(n3330), .A2(n3379), .ZN(n3370) );
  INV_X1 U2592 ( .A(n4478), .ZN(n4400) );
  INV_X1 U2593 ( .A(n3319), .ZN(n3307) );
  NOR2_X1 U2594 ( .A1(n3280), .A2(n3307), .ZN(n3330) );
  OR2_X1 U2595 ( .A1(n3258), .A2(n3263), .ZN(n3280) );
  INV_X1 U2596 ( .A(n3231), .ZN(n3227) );
  NAND2_X1 U2597 ( .A1(n2077), .A2(n3084), .ZN(n3226) );
  AND2_X1 U2598 ( .A1(n3084), .A2(n2114), .ZN(n3228) );
  AND2_X1 U2599 ( .A1(n3022), .A2(n3001), .ZN(n3084) );
  NOR2_X1 U2600 ( .A1(n2982), .A2(n2651), .ZN(n3069) );
  MUX2_X1 U2601 ( .A(n2790), .B(DATAI_3_), .S(n3831), .Z(n2986) );
  NAND2_X1 U2602 ( .A1(n3100), .A2(n2568), .ZN(n4713) );
  INV_X1 U2603 ( .A(n4331), .ZN(n4473) );
  OR2_X1 U2604 ( .A1(n4554), .A2(n2835), .ZN(n4478) );
  AND3_X1 U2605 ( .A1(n2647), .A2(n2646), .A3(n2830), .ZN(n2670) );
  INV_X1 U2606 ( .A(n2208), .ZN(n2207) );
  INV_X1 U2607 ( .A(IR_REG_21__SCAN_IN), .ZN(n2565) );
  INV_X1 U2608 ( .A(IR_REG_20__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U2609 ( .A(n2408), .B(IR_REG_11__SCAN_IN), .ZN(n3490) );
  OR3_X1 U2610 ( .A1(n2374), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2377) );
  NOR2_X1 U2611 ( .A1(n2377), .A2(IR_REG_9__SCAN_IN), .ZN(n2397) );
  INV_X1 U2612 ( .A(IR_REG_7__SCAN_IN), .ZN(n2360) );
  AOI21_X1 U2613 ( .B1(n3421), .B2(n2153), .A(n2149), .ZN(n2148) );
  NAND2_X1 U2614 ( .A1(n2150), .A2(n3435), .ZN(n2149) );
  NAND2_X1 U2615 ( .A1(n2153), .A2(n2155), .ZN(n2150) );
  INV_X1 U2616 ( .A(n3263), .ZN(n3291) );
  AND2_X1 U2617 ( .A1(n3249), .A2(n3246), .ZN(n3247) );
  INV_X1 U2618 ( .A(n2986), .ZN(n3094) );
  AND4_X1 U2619 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n4255)
         );
  INV_X1 U2620 ( .A(n4460), .ZN(n4386) );
  INV_X1 U2621 ( .A(n2867), .ZN(n2953) );
  NAND2_X1 U2622 ( .A1(n3563), .A2(n3562), .ZN(n3654) );
  AOI21_X1 U2623 ( .B1(n3421), .B2(n2152), .A(n2155), .ZN(n2151) );
  AND2_X1 U2624 ( .A1(n3578), .A2(n2145), .ZN(n2144) );
  NAND2_X1 U2625 ( .A1(n2147), .A2(n3708), .ZN(n2143) );
  OR2_X1 U2626 ( .A1(n2146), .A2(n3562), .ZN(n2145) );
  INV_X1 U2627 ( .A(n3076), .ZN(n3083) );
  NAND2_X1 U2628 ( .A1(n2901), .A2(n2900), .ZN(n3745) );
  INV_X1 U2629 ( .A(n3747), .ZN(n3752) );
  INV_X1 U2630 ( .A(n3742), .ZN(n3759) );
  OR2_X1 U2631 ( .A1(n2519), .A2(n2518), .ZN(n4279) );
  NAND4_X1 U2632 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n4333)
         );
  NAND4_X1 U2633 ( .A1(n2485), .A2(n2484), .A3(n2483), .A4(n2482), .ZN(n4357)
         );
  NAND4_X1 U2634 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n4461)
         );
  NAND4_X1 U2635 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n4476)
         );
  NAND4_X1 U2636 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(n3928)
         );
  NAND4_X1 U2637 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n3929)
         );
  OR2_X1 U2638 ( .A1(n2342), .A2(n3358), .ZN(n2393) );
  NAND4_X1 U2639 ( .A1(n2387), .A2(n2386), .A3(n2385), .A4(n2384), .ZN(n3930)
         );
  OR2_X1 U2640 ( .A1(n2342), .A2(n2381), .ZN(n2385) );
  NAND4_X1 U2641 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n3931)
         );
  NAND4_X1 U2642 ( .A1(n2359), .A2(n2358), .A3(n2357), .A4(n2356), .ZN(n3932)
         );
  NAND4_X1 U2643 ( .A1(n2346), .A2(n2345), .A3(n2344), .A4(n2343), .ZN(n3933)
         );
  OR2_X1 U2644 ( .A1(n2609), .A2(n3070), .ZN(n2306) );
  OR2_X1 U2645 ( .A1(n2282), .A2(n2754), .ZN(n2284) );
  XNOR2_X1 U2646 ( .A(n2134), .B(n2211), .ZN(n2785) );
  INV_X1 U2647 ( .A(n2210), .ZN(n2788) );
  OR2_X1 U2648 ( .A1(n2810), .A2(n2132), .ZN(n2125) );
  NAND2_X1 U2649 ( .A1(n2124), .A2(n2126), .ZN(n2882) );
  NOR2_X1 U2650 ( .A1(n2806), .A2(n2073), .ZN(n2809) );
  INV_X1 U2651 ( .A(n2217), .ZN(n2885) );
  AOI22_X1 U2652 ( .A1(n2963), .A2(REG2_REG_6__SCAN_IN), .B1(n4551), .B2(n2962), .ZN(n2965) );
  XNOR2_X1 U2653 ( .A(n2214), .B(n3491), .ZN(n3476) );
  NAND2_X1 U2654 ( .A1(n4574), .A2(n3496), .ZN(n4585) );
  XNOR2_X1 U2655 ( .A(n3481), .B(n2123), .ZN(n4599) );
  NAND2_X1 U2656 ( .A1(n4593), .A2(n3499), .ZN(n4117) );
  XNOR2_X1 U2657 ( .A(n4131), .B(n4694), .ZN(n4609) );
  NAND2_X1 U2658 ( .A1(n4622), .A2(n4122), .ZN(n4636) );
  OAI21_X1 U2659 ( .B1(n2220), .B2(n2219), .A(n2218), .ZN(n4143) );
  AOI21_X1 U2660 ( .B1(n2222), .B2(n4641), .A(n2225), .ZN(n2218) );
  NAND2_X1 U2661 ( .A1(n2193), .A2(n2191), .ZN(n2195) );
  NAND2_X1 U2662 ( .A1(n2100), .A2(n2099), .ZN(n4179) );
  NAND2_X1 U2663 ( .A1(n2100), .A2(n3820), .ZN(n4177) );
  INV_X1 U2664 ( .A(n2535), .ZN(n2190) );
  NAND2_X1 U2665 ( .A1(n2200), .A2(n2464), .ZN(n4349) );
  NAND2_X1 U2666 ( .A1(n2103), .A2(n3885), .ZN(n4369) );
  NAND2_X1 U2667 ( .A1(n2199), .A2(n2198), .ZN(n3396) );
  AND2_X1 U2668 ( .A1(n2199), .A2(n2078), .ZN(n3398) );
  OR2_X1 U2669 ( .A1(n3369), .A2(n2427), .ZN(n2199) );
  NAND2_X1 U2670 ( .A1(n2205), .A2(n2203), .ZN(n3274) );
  CLKBUF_X1 U2671 ( .A(n3049), .Z(n3051) );
  INV_X1 U2672 ( .A(n4341), .ZN(n4664) );
  NAND2_X1 U2673 ( .A1(n2069), .A2(REG1_REG_2__SCAN_IN), .ZN(n2281) );
  INV_X1 U2674 ( .A(n4658), .ZN(n4381) );
  NAND2_X1 U2675 ( .A1(n2755), .A2(IR_REG_31__SCAN_IN), .ZN(n2248) );
  XNOR2_X1 U2676 ( .A(n2624), .B(IR_REG_24__SCAN_IN), .ZN(n2739) );
  INV_X1 U2677 ( .A(n3490), .ZN(n4696) );
  INV_X1 U2678 ( .A(IR_REG_1__SCAN_IN), .ZN(n2258) );
  INV_X1 U2679 ( .A(IR_REG_0__SCAN_IN), .ZN(n4699) );
  AND2_X1 U2680 ( .A1(n2230), .A2(n2176), .ZN(n2168) );
  INV_X1 U2681 ( .A(n2137), .ZN(n4656) );
  OAI21_X1 U2682 ( .B1(n4647), .B2(n2139), .A(n2138), .ZN(n2137) );
  AOI21_X1 U2683 ( .B1(n4164), .B2(n4374), .A(n2117), .ZN(n2116) );
  OR2_X1 U2684 ( .A1(n4496), .A2(n4486), .ZN(n2653) );
  OAI21_X1 U2685 ( .B1(n2674), .B2(n4718), .A(n2104), .ZN(U3515) );
  AND2_X1 U2686 ( .A1(n2673), .A2(n2087), .ZN(n2104) );
  OR2_X1 U2687 ( .A1(n4158), .A2(n4546), .ZN(n2673) );
  INV_X1 U2688 ( .A(n3216), .ZN(n2185) );
  AND2_X1 U2689 ( .A1(n2215), .A2(n4551), .ZN(n2060) );
  XNOR2_X1 U2690 ( .A(n2284), .B(n2283), .ZN(n2775) );
  NOR2_X1 U2691 ( .A1(n3452), .A2(n4474), .ZN(n2061) );
  INV_X1 U2692 ( .A(n3113), .ZN(n3873) );
  AND2_X1 U2693 ( .A1(n2478), .A2(n2464), .ZN(n2063) );
  OR2_X1 U2694 ( .A1(n2130), .A2(n2129), .ZN(n2064) );
  OR2_X1 U2695 ( .A1(n2060), .A2(n2212), .ZN(n2065) );
  INV_X1 U2696 ( .A(n3802), .ZN(n2095) );
  INV_X1 U2697 ( .A(n3347), .ZN(n3379) );
  AND2_X1 U2698 ( .A1(n2082), .A2(n2101), .ZN(n2066) );
  AND2_X1 U2699 ( .A1(n2108), .A2(n3756), .ZN(n2067) );
  INV_X1 U2700 ( .A(n4436), .ZN(n3661) );
  NAND4_X1 U2701 ( .A1(n2511), .A2(n2510), .A3(n2509), .A4(n2508), .ZN(n4436)
         );
  AND2_X1 U2702 ( .A1(n4352), .A2(n4386), .ZN(n2068) );
  INV_X1 U2703 ( .A(n4641), .ZN(n2224) );
  AND2_X1 U2705 ( .A1(n2251), .A2(n2752), .ZN(n2069) );
  OR2_X1 U2706 ( .A1(n2275), .A2(n2266), .ZN(n2070) );
  XNOR2_X1 U2707 ( .A(n2248), .B(IR_REG_30__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U2708 ( .A1(n2165), .A2(n3549), .ZN(n3726) );
  NAND2_X1 U2709 ( .A1(n2503), .A2(n2502), .ZN(n4269) );
  NAND2_X1 U2710 ( .A1(n4200), .A2(n4399), .ZN(n2071) );
  NOR2_X1 U2711 ( .A1(n3929), .A2(n3307), .ZN(n2072) );
  AND2_X1 U2712 ( .A1(n2807), .A2(n2813), .ZN(n2073) );
  AND2_X1 U2713 ( .A1(n4552), .A2(REG1_REG_2__SCAN_IN), .ZN(n2074) );
  NAND2_X1 U2714 ( .A1(n2217), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2715 ( .A1(n3717), .A2(n3718), .ZN(n3635) );
  AND2_X1 U2716 ( .A1(n2193), .A2(n2190), .ZN(n2075) );
  AND3_X1 U2717 ( .A1(n2240), .A2(n2239), .A3(n2238), .ZN(n2462) );
  INV_X1 U2718 ( .A(n4277), .ZN(n4270) );
  INV_X1 U2719 ( .A(IR_REG_26__SCAN_IN), .ZN(n2246) );
  OR2_X1 U2720 ( .A1(n4401), .A2(n4203), .ZN(n2076) );
  INV_X1 U2721 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2129) );
  INV_X1 U2722 ( .A(n2151), .ZN(n3434) );
  AND2_X1 U2723 ( .A1(n2114), .A2(n3227), .ZN(n2077) );
  INV_X1 U2724 ( .A(n3737), .ZN(n2174) );
  NAND2_X1 U2725 ( .A1(n3927), .A2(n3413), .ZN(n2078) );
  AND2_X1 U2726 ( .A1(n3517), .A2(n3752), .ZN(n2079) );
  INV_X1 U2727 ( .A(n3413), .ZN(n3428) );
  NAND2_X1 U2728 ( .A1(n4236), .A2(n2111), .ZN(n2113) );
  OR2_X1 U2729 ( .A1(n3682), .A2(n4460), .ZN(n2080) );
  INV_X1 U2730 ( .A(n3708), .ZN(n2146) );
  INV_X1 U2731 ( .A(n3577), .ZN(n2147) );
  AND2_X1 U2732 ( .A1(n4279), .A2(n4259), .ZN(n2081) );
  AND2_X1 U2733 ( .A1(n4327), .A2(n2594), .ZN(n2082) );
  OR2_X1 U2734 ( .A1(n3861), .A2(n2592), .ZN(n2083) );
  INV_X1 U2735 ( .A(n3144), .ZN(n3171) );
  INV_X1 U2736 ( .A(n4198), .ZN(n4418) );
  AND4_X1 U2737 ( .A1(n2533), .A2(n2532), .A3(n2531), .A4(n2530), .ZN(n4198)
         );
  AND2_X1 U2738 ( .A1(n2173), .A2(n2079), .ZN(n2084) );
  INV_X1 U2739 ( .A(n3885), .ZN(n2102) );
  NOR2_X1 U2740 ( .A1(n3174), .A2(n3149), .ZN(n2085) );
  NOR2_X1 U2741 ( .A1(n2618), .A2(n2208), .ZN(n2569) );
  INV_X1 U2742 ( .A(IR_REG_15__SCAN_IN), .ZN(n2239) );
  AND2_X1 U2743 ( .A1(n2068), .A2(n4339), .ZN(n2086) );
  INV_X1 U2744 ( .A(n4130), .ZN(n4694) );
  OR2_X1 U2745 ( .A1(n4719), .A2(n2671), .ZN(n2087) );
  INV_X1 U2746 ( .A(n4186), .ZN(n4399) );
  AND2_X1 U2747 ( .A1(n2125), .A2(n2131), .ZN(n2088) );
  INV_X1 U2748 ( .A(n2790), .ZN(n2211) );
  INV_X1 U2749 ( .A(n4592), .ZN(n2123) );
  INV_X1 U2750 ( .A(n4571), .ZN(n2121) );
  AND2_X1 U2751 ( .A1(n2326), .A2(n2325), .ZN(n2886) );
  OR2_X1 U2752 ( .A1(n3009), .A2(REG1_REG_7__SCAN_IN), .ZN(n2089) );
  NAND3_X1 U2753 ( .A1(n2251), .A2(n2752), .A3(REG1_REG_1__SCAN_IN), .ZN(n2256) );
  NAND2_X1 U2754 ( .A1(n2069), .A2(REG1_REG_0__SCAN_IN), .ZN(n2270) );
  NAND2_X1 U2755 ( .A1(n3325), .A2(n2093), .ZN(n2091) );
  OAI21_X1 U2756 ( .B1(n4194), .B2(n2098), .A(n2096), .ZN(n2658) );
  NAND2_X1 U2757 ( .A1(n3463), .A2(n3874), .ZN(n2103) );
  AND3_X1 U2758 ( .A1(n2115), .A2(n2062), .A3(n2614), .ZN(n2572) );
  NAND3_X1 U2759 ( .A1(n2115), .A2(n2614), .A3(n2106), .ZN(n2755) );
  INV_X1 U2760 ( .A(n2113), .ZN(n4182) );
  NAND3_X1 U2761 ( .A1(n2077), .A2(n3084), .A3(n3221), .ZN(n3258) );
  OR2_X2 U2762 ( .A1(n2618), .A2(IR_REG_26__SCAN_IN), .ZN(n2627) );
  AND2_X2 U2763 ( .A1(n2424), .A2(n4077), .ZN(n2115) );
  AND2_X2 U2764 ( .A1(n2620), .A2(n2245), .ZN(n2614) );
  NAND2_X1 U2765 ( .A1(n2120), .A2(n2116), .ZN(U3354) );
  OAI21_X1 U2766 ( .B1(n4160), .B2(n4159), .A(n4365), .ZN(n2120) );
  NAND2_X1 U2767 ( .A1(n4230), .A2(n3894), .ZN(n4213) );
  MUX2_X2 U2768 ( .A(n2055), .B(n2263), .S(n2271), .Z(n3161) );
  INV_X1 U2769 ( .A(n4160), .ZN(n2669) );
  MUX2_X2 U2770 ( .A(n2665), .B(n2664), .S(IR_REG_28__SCAN_IN), .Z(n2271) );
  INV_X1 U2771 ( .A(n2886), .ZN(n2130) );
  INV_X1 U2772 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2132) );
  OAI22_X2 U2773 ( .A1(n3563), .A2(n2143), .B1(n2144), .B2(n3577), .ZN(n3717)
         );
  INV_X1 U2774 ( .A(n2148), .ZN(n3520) );
  INV_X1 U2775 ( .A(n3423), .ZN(n2158) );
  NAND2_X1 U2776 ( .A1(n3540), .A2(n3539), .ZN(n3692) );
  NOR2_X1 U2777 ( .A1(n3547), .A2(n2167), .ZN(n2166) );
  INV_X1 U2778 ( .A(n3539), .ZN(n2167) );
  NAND2_X1 U2779 ( .A1(n3602), .A2(n2176), .ZN(n2175) );
  NAND2_X1 U2780 ( .A1(n2175), .A2(n2084), .ZN(n2178) );
  AOI21_X1 U2781 ( .B1(n3602), .B2(n2168), .A(n2170), .ZN(n2169) );
  NAND2_X1 U2782 ( .A1(n2175), .A2(n3737), .ZN(n3628) );
  NAND2_X1 U2783 ( .A1(n3602), .A2(n3666), .ZN(n3736) );
  NAND2_X1 U2784 ( .A1(n2178), .A2(n2169), .ZN(U3217) );
  INV_X1 U2785 ( .A(n3215), .ZN(n2184) );
  NAND2_X1 U2786 ( .A1(n4211), .A2(n2536), .ZN(n2193) );
  AOI21_X2 U2787 ( .B1(n4211), .B2(n2189), .A(n2186), .ZN(n2655) );
  NAND2_X1 U2788 ( .A1(n3369), .A2(n2198), .ZN(n2196) );
  NAND2_X1 U2789 ( .A1(n2196), .A2(n2197), .ZN(n3448) );
  NAND2_X1 U2790 ( .A1(n3257), .A2(n2203), .ZN(n2201) );
  NAND2_X1 U2791 ( .A1(n2201), .A2(n2202), .ZN(n3324) );
  NAND2_X1 U2792 ( .A1(n2503), .A2(n2206), .ZN(n4268) );
  OAI21_X1 U2793 ( .B1(n2966), .B2(n2065), .A(n2089), .ZN(n2214) );
  NOR2_X1 U2794 ( .A1(n2966), .A2(n2060), .ZN(n3007) );
  OR2_X1 U2795 ( .A1(n2214), .A2(n3491), .ZN(n2213) );
  INV_X1 U2796 ( .A(n4642), .ZN(n2220) );
  NOR2_X1 U2797 ( .A1(n4686), .A2(n4140), .ZN(n2225) );
  NAND2_X1 U2798 ( .A1(n2578), .A2(n3769), .ZN(n3863) );
  NAND2_X1 U2799 ( .A1(n4548), .A2(n2253), .ZN(n2275) );
  XNOR2_X1 U2800 ( .A(n2055), .B(n2682), .ZN(n2686) );
  AND2_X1 U2801 ( .A1(n2277), .A2(n2276), .ZN(n2226) );
  NAND2_X1 U2802 ( .A1(n2287), .A2(n2286), .ZN(n2578) );
  AND2_X1 U2803 ( .A1(n2309), .A2(n2312), .ZN(n2227) );
  NAND2_X1 U2804 ( .A1(n2556), .A2(n2476), .ZN(n2228) );
  AND2_X1 U2805 ( .A1(n4306), .A2(n3856), .ZN(n2229) );
  AND3_X1 U2806 ( .A1(n3622), .A2(n3623), .A3(n3752), .ZN(n2230) );
  INV_X2 U2807 ( .A(n2994), .ZN(n3615) );
  INV_X1 U2808 ( .A(IR_REG_13__SCAN_IN), .ZN(n2235) );
  INV_X1 U2809 ( .A(IR_REG_25__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U2810 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
  AOI21_X1 U2811 ( .B1(n3520), .B2(n3519), .A(n3518), .ZN(n3529) );
  NAND2_X1 U2812 ( .A1(n3690), .A2(n3548), .ZN(n3549) );
  NOR2_X1 U2813 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  INV_X1 U2814 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2353) );
  INV_X1 U2815 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U2816 ( .A1(n2490), .A2(REG3_REG_20__SCAN_IN), .ZN(n2506) );
  NOR2_X1 U2817 ( .A1(n4198), .A2(n4221), .ZN(n2535) );
  NAND2_X1 U2818 ( .A1(n4436), .A2(n2512), .ZN(n2513) );
  OR2_X1 U2819 ( .A1(n3452), .A2(n3406), .ZN(n3804) );
  NAND2_X1 U2820 ( .A1(n2339), .A2(REG3_REG_7__SCAN_IN), .ZN(n2354) );
  INV_X1 U2821 ( .A(n4352), .ZN(n4356) );
  INV_X1 U2822 ( .A(IR_REG_28__SCAN_IN), .ZN(n2247) );
  OR2_X1 U2823 ( .A1(n2506), .A2(n2505), .ZN(n2515) );
  AOI21_X2 U2824 ( .B1(n3342), .B2(n3341), .A(n3340), .ZN(n3421) );
  AND2_X1 U2825 ( .A1(n2928), .A2(n2931), .ZN(n2929) );
  OR2_X1 U2826 ( .A1(n2354), .A2(n2353), .ZN(n2368) );
  OR2_X1 U2827 ( .A1(n2401), .A2(n2400), .ZN(n2414) );
  NOR2_X1 U2828 ( .A1(n2429), .A2(n2428), .ZN(n2436) );
  AND2_X1 U2829 ( .A1(n3609), .A2(n2843), .ZN(n3917) );
  OR2_X1 U2830 ( .A1(n2537), .A2(n3741), .ZN(n2542) );
  INV_X1 U2831 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U2832 ( .A1(n4351), .A2(n4146), .ZN(n3085) );
  INV_X1 U2833 ( .A(n3851), .ZN(n2555) );
  INV_X1 U2834 ( .A(n3406), .ZN(n4474) );
  AND2_X1 U2835 ( .A1(n2629), .A2(n2734), .ZN(n2758) );
  NOR2_X1 U2836 ( .A1(n2323), .A2(IR_REG_5__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U2837 ( .A1(n3248), .A2(n3247), .ZN(n3306) );
  NAND2_X1 U2838 ( .A1(n2317), .A2(REG3_REG_5__SCAN_IN), .ZN(n2330) );
  NOR2_X1 U2839 ( .A1(n2368), .A2(n2367), .ZN(n2382) );
  AND3_X1 U2840 ( .A1(n3056), .A2(n2832), .A3(n2831), .ZN(n2852) );
  OR2_X1 U2841 ( .A1(n2609), .A2(n3659), .ZN(n2498) );
  NAND4_X1 U2842 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(n3452)
         );
  AOI21_X1 U2843 ( .B1(n2715), .B2(REG1_REG_1__SCAN_IN), .A(n2714), .ZN(n2717)
         );
  INV_X1 U2844 ( .A(n4627), .ZN(n4652) );
  AND2_X1 U2845 ( .A1(n4326), .A2(n4327), .ZN(n4354) );
  AOI21_X1 U2846 ( .B1(n3448), .B2(n2444), .A(n2443), .ZN(n3462) );
  AOI21_X1 U2847 ( .B1(n2758), .B2(n3964), .A(n2760), .ZN(n2832) );
  AND2_X1 U2848 ( .A1(n3916), .A2(n2821), .ZN(n4711) );
  INV_X1 U2849 ( .A(n3053), .ZN(n2848) );
  INV_X1 U2850 ( .A(n2821), .ZN(n3920) );
  INV_X1 U2851 ( .A(n3489), .ZN(n4115) );
  AND2_X1 U2852 ( .A1(n2685), .A2(n2683), .ZN(n4650) );
  NAND2_X1 U2853 ( .A1(n2852), .A2(n2837), .ZN(n3747) );
  INV_X1 U2854 ( .A(n3745), .ZN(n3763) );
  INV_X1 U2855 ( .A(n4404), .ZN(n4161) );
  NAND4_X1 U2856 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n4445)
         );
  OR2_X1 U2857 ( .A1(n2772), .A2(n2850), .ZN(n4657) );
  INV_X1 U2858 ( .A(n4374), .ZN(n4368) );
  OR2_X1 U2859 ( .A1(n4158), .A2(n4486), .ZN(n2676) );
  NAND2_X1 U2860 ( .A1(n4727), .A2(n4351), .ZN(n4486) );
  INV_X1 U2861 ( .A(n4727), .ZN(n4724) );
  NAND2_X1 U2862 ( .A1(n4719), .A2(n4351), .ZN(n4546) );
  INV_X1 U2863 ( .A(n4719), .ZN(n4718) );
  INV_X1 U2864 ( .A(n4682), .ZN(n4681) );
  NAND2_X1 U2865 ( .A1(n2759), .A2(n2848), .ZN(n4682) );
  AND2_X1 U2866 ( .A1(n2896), .A2(STATE_REG_SCAN_IN), .ZN(n4683) );
  INV_X1 U2867 ( .A(n4134), .ZN(n4690) );
  NOR2_X1 U2868 ( .A1(n2378), .A2(n2397), .ZN(n4558) );
  INV_X1 U2869 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U2870 ( .A1(n2420), .A2(n2235), .ZN(n2237) );
  NAND2_X1 U2871 ( .A1(n2282), .A2(n2283), .ZN(n2296) );
  INV_X1 U2872 ( .A(n2296), .ZN(n2236) );
  NAND2_X1 U2873 ( .A1(n2236), .A2(n2227), .ZN(n2322) );
  NOR2_X2 U2874 ( .A1(n2237), .A2(n2322), .ZN(n2424) );
  NOR2_X1 U2875 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2241)
         );
  NOR2_X2 U2876 ( .A1(n2475), .A2(n2242), .ZN(n2557) );
  INV_X1 U2877 ( .A(n4548), .ZN(n2251) );
  INV_X1 U2878 ( .A(n2253), .ZN(n2250) );
  INV_X1 U2879 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2252) );
  AND2_X2 U2880 ( .A1(n4548), .A2(n2250), .ZN(n2290) );
  NAND2_X1 U2881 ( .A1(n2290), .A2(REG2_REG_1__SCAN_IN), .ZN(n2255) );
  INV_X1 U2882 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3160) );
  OR2_X1 U2883 ( .A1(n2275), .A2(n3160), .ZN(n2254) );
  NAND4_X1 U2884 ( .A1(n2257), .A2(n2256), .A3(n2255), .A4(n2254), .ZN(n2272)
         );
  INV_X1 U2885 ( .A(n2272), .ZN(n2265) );
  NAND2_X1 U2886 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2259)
         );
  INV_X1 U2887 ( .A(DATAI_1_), .ZN(n2263) );
  NAND2_X1 U2888 ( .A1(n2627), .A2(IR_REG_31__SCAN_IN), .ZN(n2261) );
  INV_X1 U2889 ( .A(IR_REG_27__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2890 ( .A1(n2261), .A2(n2260), .ZN(n2665) );
  NAND2_X1 U2891 ( .A1(n2272), .A2(n3161), .ZN(n3764) );
  INV_X1 U2892 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2893 ( .A1(n2290), .A2(REG2_REG_0__SCAN_IN), .ZN(n2269) );
  INV_X1 U2894 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2267) );
  NAND4_X2 U2895 ( .A1(n2270), .A2(n2070), .A3(n2269), .A4(n2268), .ZN(n2576)
         );
  AND2_X1 U2896 ( .A1(n2576), .A2(n2867), .ZN(n2859) );
  NAND2_X1 U2897 ( .A1(n2575), .A2(n2859), .ZN(n2858) );
  NAND2_X1 U2898 ( .A1(n2823), .A2(n2264), .ZN(n2273) );
  AND2_X2 U2899 ( .A1(n2858), .A2(n2273), .ZN(n2872) );
  INV_X1 U2900 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2274) );
  NAND2_X1 U2901 ( .A1(n2290), .A2(REG2_REG_2__SCAN_IN), .ZN(n2276) );
  INV_X1 U2902 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2279) );
  OR2_X1 U2903 ( .A1(n2278), .A2(n2279), .ZN(n2280) );
  INV_X1 U2904 ( .A(n2288), .ZN(n2287) );
  INV_X1 U2905 ( .A(DATAI_2_), .ZN(n2285) );
  MUX2_X1 U2906 ( .A(n2775), .B(n2285), .S(n2056), .Z(n2983) );
  NAND2_X1 U2907 ( .A1(n2288), .A2(n2983), .ZN(n3769) );
  NAND2_X1 U2908 ( .A1(n2872), .A2(n3863), .ZN(n2871) );
  OR2_X1 U2909 ( .A1(n2288), .A2(n2286), .ZN(n2289) );
  NAND2_X1 U2910 ( .A1(n2871), .A2(n2289), .ZN(n2975) );
  NAND2_X1 U2911 ( .A1(n3828), .A2(REG1_REG_3__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2912 ( .A1(n3827), .A2(REG2_REG_3__SCAN_IN), .ZN(n2294) );
  OR2_X1 U2913 ( .A1(n2609), .A2(REG3_REG_3__SCAN_IN), .ZN(n2293) );
  INV_X1 U2914 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2291) );
  OR2_X1 U2915 ( .A1(n2278), .A2(n2291), .ZN(n2292) );
  NAND2_X1 U2916 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .ZN(n2310) );
  XNOR2_X1 U2917 ( .A(n2310), .B(IR_REG_3__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U2918 ( .A1(n3936), .A2(n2986), .ZN(n2297) );
  NAND2_X1 U2919 ( .A1(n2975), .A2(n2297), .ZN(n2299) );
  OR2_X1 U2920 ( .A1(n3936), .A2(n2986), .ZN(n2298) );
  NAND2_X1 U2921 ( .A1(n2299), .A2(n2298), .ZN(n3049) );
  INV_X1 U2922 ( .A(n3049), .ZN(n2314) );
  NAND2_X1 U2923 ( .A1(n3827), .A2(REG2_REG_4__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2924 ( .A1(n2069), .A2(REG1_REG_4__SCAN_IN), .ZN(n2307) );
  INV_X1 U2925 ( .A(n2317), .ZN(n2303) );
  INV_X1 U2926 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2301) );
  INV_X1 U2927 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2300) );
  NAND2_X1 U2928 ( .A1(n2301), .A2(n2300), .ZN(n2302) );
  NAND2_X1 U2929 ( .A1(n2303), .A2(n2302), .ZN(n3070) );
  INV_X1 U2930 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2304) );
  OR2_X1 U2931 ( .A1(n2278), .A2(n2304), .ZN(n2305) );
  NAND2_X1 U2932 ( .A1(n2310), .A2(n2309), .ZN(n2311) );
  NAND2_X1 U2933 ( .A1(n2311), .A2(IR_REG_31__SCAN_IN), .ZN(n2313) );
  XNOR2_X1 U2934 ( .A(n2313), .B(n2312), .ZN(n2791) );
  INV_X1 U2935 ( .A(DATAI_4_), .ZN(n2725) );
  MUX2_X1 U2936 ( .A(n2791), .B(n2725), .S(n3831), .Z(n3068) );
  OR2_X1 U2937 ( .A1(n3127), .A2(n3068), .ZN(n3772) );
  NAND2_X1 U2938 ( .A1(n3127), .A2(n3068), .ZN(n3775) );
  NAND2_X1 U2939 ( .A1(n2314), .A2(n3864), .ZN(n3048) );
  INV_X1 U2940 ( .A(n3068), .ZN(n2923) );
  NAND2_X1 U2941 ( .A1(n3127), .A2(n2923), .ZN(n2315) );
  NAND2_X1 U2942 ( .A1(n3048), .A2(n2315), .ZN(n3017) );
  NAND2_X1 U2943 ( .A1(n3828), .A2(REG1_REG_5__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2944 ( .A1(n3827), .A2(REG2_REG_5__SCAN_IN), .ZN(n2320) );
  INV_X1 U2945 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2316) );
  OR2_X1 U2946 ( .A1(n2278), .A2(n2316), .ZN(n2319) );
  OAI21_X1 U2947 ( .B1(n2317), .B2(REG3_REG_5__SCAN_IN), .A(n2330), .ZN(n3128)
         );
  OR2_X1 U2948 ( .A1(n2609), .A2(n3128), .ZN(n2318) );
  NAND4_X1 U2949 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n3935)
         );
  NAND2_X1 U2950 ( .A1(n2323), .A2(IR_REG_31__SCAN_IN), .ZN(n2324) );
  MUX2_X1 U2951 ( .A(IR_REG_31__SCAN_IN), .B(n2324), .S(IR_REG_5__SCAN_IN), 
        .Z(n2326) );
  INV_X1 U2952 ( .A(n2348), .ZN(n2325) );
  MUX2_X1 U2953 ( .A(n2886), .B(DATAI_5_), .S(n3831), .Z(n3130) );
  OR2_X1 U2954 ( .A1(n3935), .A2(n3130), .ZN(n2327) );
  NAND2_X1 U2955 ( .A1(n3017), .A2(n2327), .ZN(n2329) );
  NAND2_X1 U2956 ( .A1(n3935), .A2(n3130), .ZN(n2328) );
  NAND2_X1 U2957 ( .A1(n3827), .A2(REG2_REG_6__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U2958 ( .A1(n3828), .A2(REG1_REG_6__SCAN_IN), .ZN(n2335) );
  AND2_X1 U2959 ( .A1(n2330), .A2(n2883), .ZN(n2331) );
  OR2_X1 U2960 ( .A1(n2331), .A2(n2339), .ZN(n3087) );
  OR2_X1 U2961 ( .A1(n2609), .A2(n3087), .ZN(n2334) );
  INV_X1 U2962 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2332) );
  OR2_X1 U2963 ( .A1(n2278), .A2(n2332), .ZN(n2333) );
  NAND4_X1 U2964 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n3934)
         );
  OR2_X1 U2965 ( .A1(n2348), .A2(n2754), .ZN(n2337) );
  XNOR2_X1 U2966 ( .A(n2337), .B(IR_REG_6__SCAN_IN), .ZN(n4551) );
  MUX2_X1 U2967 ( .A(n4551), .B(DATAI_6_), .S(n3831), .Z(n3076) );
  AND2_X1 U2968 ( .A1(n3934), .A2(n3076), .ZN(n2338) );
  OAI22_X1 U2969 ( .A1(n3074), .A2(n2338), .B1(n3076), .B2(n3934), .ZN(n3122)
         );
  INV_X1 U2970 ( .A(n3122), .ZN(n2350) );
  NAND2_X1 U2971 ( .A1(n3827), .A2(REG2_REG_7__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2972 ( .A1(n3828), .A2(REG1_REG_7__SCAN_IN), .ZN(n2345) );
  OR2_X1 U2973 ( .A1(n2339), .A2(REG3_REG_7__SCAN_IN), .ZN(n2340) );
  NAND2_X1 U2974 ( .A1(n2354), .A2(n2340), .ZN(n3170) );
  OR2_X1 U2975 ( .A1(n2609), .A2(n3170), .ZN(n2344) );
  INV_X1 U2976 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2341) );
  OR2_X1 U2977 ( .A1(n2342), .A2(n2341), .ZN(n2343) );
  NAND2_X1 U2978 ( .A1(n2348), .A2(n2347), .ZN(n2374) );
  NAND2_X1 U2979 ( .A1(n2374), .A2(IR_REG_31__SCAN_IN), .ZN(n2361) );
  XNOR2_X1 U2980 ( .A(n2361), .B(n2360), .ZN(n2971) );
  INV_X1 U2981 ( .A(DATAI_7_), .ZN(n2349) );
  MUX2_X1 U2982 ( .A(n2971), .B(n2349), .S(n3831), .Z(n3144) );
  OR2_X1 U2983 ( .A1(n3933), .A2(n3144), .ZN(n2582) );
  NAND2_X1 U2984 ( .A1(n3933), .A2(n3144), .ZN(n3787) );
  NAND2_X1 U2985 ( .A1(n2582), .A2(n3787), .ZN(n3113) );
  NAND2_X1 U2986 ( .A1(n2350), .A2(n3113), .ZN(n3121) );
  NAND2_X1 U2987 ( .A1(n3933), .A2(n3171), .ZN(n2351) );
  NAND2_X1 U2988 ( .A1(n3121), .A2(n2351), .ZN(n3229) );
  NAND2_X1 U2989 ( .A1(n3828), .A2(REG1_REG_8__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U2990 ( .A1(n3827), .A2(REG2_REG_8__SCAN_IN), .ZN(n2358) );
  INV_X1 U2991 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2352) );
  OR2_X1 U2992 ( .A1(n2342), .A2(n2352), .ZN(n2357) );
  NAND2_X1 U2993 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  NAND2_X1 U2994 ( .A1(n2368), .A2(n2355), .ZN(n4659) );
  OR2_X1 U2995 ( .A1(n2609), .A2(n4659), .ZN(n2356) );
  NAND2_X1 U2996 ( .A1(n2361), .A2(n2360), .ZN(n2362) );
  NAND2_X1 U2997 ( .A1(n2362), .A2(IR_REG_31__SCAN_IN), .ZN(n2363) );
  XNOR2_X1 U2998 ( .A(n2363), .B(IR_REG_8__SCAN_IN), .ZN(n4550) );
  MUX2_X1 U2999 ( .A(n4550), .B(DATAI_8_), .S(n3831), .Z(n3231) );
  OR2_X1 U3000 ( .A1(n3932), .A2(n3231), .ZN(n2364) );
  NAND2_X1 U3001 ( .A1(n3229), .A2(n2364), .ZN(n2366) );
  NAND2_X1 U3002 ( .A1(n3932), .A2(n3231), .ZN(n2365) );
  NAND2_X1 U3003 ( .A1(n3828), .A2(REG1_REG_9__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3004 ( .A1(n3827), .A2(REG2_REG_9__SCAN_IN), .ZN(n2372) );
  AND2_X1 U3005 ( .A1(n2368), .A2(n2367), .ZN(n2369) );
  OR2_X1 U3006 ( .A1(n2369), .A2(n2382), .ZN(n3225) );
  OR2_X1 U3007 ( .A1(n2609), .A2(n3225), .ZN(n2371) );
  INV_X1 U3008 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3210) );
  OR2_X1 U3009 ( .A1(n2342), .A2(n3210), .ZN(n2370) );
  NAND2_X1 U3010 ( .A1(n2377), .A2(IR_REG_31__SCAN_IN), .ZN(n2375) );
  MUX2_X1 U3011 ( .A(IR_REG_31__SCAN_IN), .B(n2375), .S(IR_REG_9__SCAN_IN), 
        .Z(n2376) );
  INV_X1 U3012 ( .A(n2376), .ZN(n2378) );
  MUX2_X1 U3013 ( .A(n4558), .B(DATAI_9_), .S(n3831), .Z(n3214) );
  AND2_X1 U3014 ( .A1(n3931), .A2(n3214), .ZN(n2380) );
  OR2_X1 U3015 ( .A1(n3931), .A2(n3214), .ZN(n2379) );
  OAI21_X2 U3016 ( .B1(n3189), .B2(n2380), .A(n2379), .ZN(n3257) );
  NAND2_X1 U3017 ( .A1(n3828), .A2(REG1_REG_10__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U3018 ( .A1(n3827), .A2(REG2_REG_10__SCAN_IN), .ZN(n2386) );
  INV_X1 U3019 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2381) );
  NOR2_X1 U3020 ( .A1(n2382), .A2(REG3_REG_10__SCAN_IN), .ZN(n2383) );
  OR2_X1 U3021 ( .A1(n2390), .A2(n2383), .ZN(n3260) );
  OR2_X1 U3022 ( .A1(n2609), .A2(n3260), .ZN(n2384) );
  OR2_X1 U3023 ( .A1(n2397), .A2(n2754), .ZN(n2388) );
  XNOR2_X1 U3024 ( .A(n2388), .B(IR_REG_10__SCAN_IN), .ZN(n4571) );
  MUX2_X1 U3025 ( .A(n4571), .B(DATAI_10_), .S(n3831), .Z(n3263) );
  NOR2_X1 U3026 ( .A1(n3930), .A2(n3263), .ZN(n2389) );
  INV_X1 U3027 ( .A(n3930), .ZN(n3318) );
  NAND2_X1 U3028 ( .A1(n3828), .A2(REG1_REG_11__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3029 ( .A1(n3827), .A2(REG2_REG_11__SCAN_IN), .ZN(n2394) );
  INV_X1 U3030 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3358) );
  OR2_X1 U3031 ( .A1(n2390), .A2(REG3_REG_11__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3032 ( .A1(n2401), .A2(n2391), .ZN(n3323) );
  OR2_X1 U3033 ( .A1(n2609), .A2(n3323), .ZN(n2392) );
  INV_X1 U3034 ( .A(IR_REG_10__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3035 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  NAND2_X1 U3036 ( .A1(n2398), .A2(IR_REG_31__SCAN_IN), .ZN(n2408) );
  INV_X1 U3037 ( .A(DATAI_11_), .ZN(n2399) );
  MUX2_X1 U3038 ( .A(n4696), .B(n2399), .S(n3831), .Z(n3319) );
  OR2_X1 U3039 ( .A1(n3929), .A2(n3319), .ZN(n3327) );
  NAND2_X1 U3040 ( .A1(n3929), .A2(n3319), .ZN(n2587) );
  NAND2_X1 U3041 ( .A1(n3327), .A2(n2587), .ZN(n3865) );
  INV_X1 U3042 ( .A(n3865), .ZN(n3271) );
  NAND2_X1 U3043 ( .A1(n3827), .A2(REG2_REG_12__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3044 ( .A1(n3828), .A2(REG1_REG_12__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3045 ( .A1(n2401), .A2(n2400), .ZN(n2402) );
  NAND2_X1 U3046 ( .A1(n2414), .A2(n2402), .ZN(n3346) );
  OR2_X1 U3047 ( .A1(n2609), .A2(n3346), .ZN(n2404) );
  INV_X1 U3048 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3383) );
  OR2_X1 U3049 ( .A1(n2342), .A2(n3383), .ZN(n2403) );
  INV_X1 U3050 ( .A(IR_REG_11__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3051 ( .A1(n2408), .A2(n2407), .ZN(n2409) );
  NAND2_X1 U3052 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U3053 ( .A(n2410), .B(IR_REG_12__SCAN_IN), .ZN(n4592) );
  MUX2_X1 U3054 ( .A(n4592), .B(DATAI_12_), .S(n3831), .Z(n3347) );
  NAND2_X1 U3055 ( .A1(n3928), .A2(n3347), .ZN(n2411) );
  OR2_X1 U3056 ( .A1(n3928), .A2(n3347), .ZN(n2412) );
  NAND2_X1 U3057 ( .A1(n2413), .A2(n2412), .ZN(n3369) );
  NAND2_X1 U3058 ( .A1(n3828), .A2(REG1_REG_13__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3059 ( .A1(n3827), .A2(REG2_REG_13__SCAN_IN), .ZN(n2418) );
  INV_X1 U3060 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3391) );
  OR2_X1 U3061 ( .A1(n2342), .A2(n3391), .ZN(n2417) );
  NAND2_X1 U3062 ( .A1(n2414), .A2(n3426), .ZN(n2415) );
  NAND2_X1 U3063 ( .A1(n2429), .A2(n2415), .ZN(n3432) );
  OR2_X1 U3064 ( .A1(n2609), .A2(n3432), .ZN(n2416) );
  INV_X1 U3065 ( .A(n2420), .ZN(n2421) );
  NOR2_X1 U3066 ( .A1(n2323), .A2(n2421), .ZN(n2422) );
  NOR2_X1 U3067 ( .A1(n2422), .A2(n2754), .ZN(n2423) );
  MUX2_X1 U3068 ( .A(n2754), .B(n2423), .S(IR_REG_13__SCAN_IN), .Z(n2426) );
  BUF_X1 U3069 ( .A(n2424), .Z(n2425) );
  OR2_X1 U3070 ( .A1(n2426), .A2(n2425), .ZN(n3489) );
  MUX2_X1 U3071 ( .A(n4115), .B(DATAI_13_), .S(n3831), .Z(n3413) );
  NOR2_X1 U3072 ( .A1(n3927), .A2(n3413), .ZN(n2427) );
  NAND2_X1 U3073 ( .A1(n3828), .A2(REG1_REG_14__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3074 ( .A1(n3827), .A2(REG2_REG_14__SCAN_IN), .ZN(n2433) );
  INV_X1 U3075 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4544) );
  OR2_X1 U3076 ( .A1(n2342), .A2(n4544), .ZN(n2432) );
  INV_X1 U3077 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2428) );
  AND2_X1 U3078 ( .A1(n2429), .A2(n2428), .ZN(n2430) );
  OR2_X1 U3079 ( .A1(n2430), .A2(n2436), .ZN(n3403) );
  OR2_X1 U3080 ( .A1(n2609), .A2(n3403), .ZN(n2431) );
  OR2_X1 U3081 ( .A1(n2425), .A2(n2754), .ZN(n2435) );
  XNOR2_X1 U3082 ( .A(n2435), .B(IR_REG_14__SCAN_IN), .ZN(n4130) );
  INV_X1 U3083 ( .A(DATAI_14_), .ZN(n4693) );
  MUX2_X1 U3084 ( .A(n4694), .B(n4693), .S(n3831), .Z(n3406) );
  NAND2_X1 U3085 ( .A1(n3452), .A2(n3406), .ZN(n3783) );
  NAND2_X1 U3086 ( .A1(n3804), .A2(n3783), .ZN(n3397) );
  NAND2_X1 U3087 ( .A1(n3827), .A2(REG2_REG_15__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3088 ( .A1(n3828), .A2(REG1_REG_15__SCAN_IN), .ZN(n2440) );
  OR2_X1 U3089 ( .A1(n2436), .A2(REG3_REG_15__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3090 ( .A1(n2456), .A2(n2437), .ZN(n3762) );
  OR2_X1 U3091 ( .A1(n2609), .A2(n3762), .ZN(n2439) );
  INV_X1 U3092 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3508) );
  OR2_X1 U3093 ( .A1(n2342), .A2(n3508), .ZN(n2438) );
  NAND2_X1 U3094 ( .A1(n2425), .A2(n2240), .ZN(n2442) );
  NAND2_X1 U3095 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  XNOR2_X1 U3096 ( .A(n2449), .B(IR_REG_15__SCAN_IN), .ZN(n4126) );
  MUX2_X1 U3097 ( .A(n4126), .B(DATAI_15_), .S(n3831), .Z(n3523) );
  NAND2_X1 U3098 ( .A1(n4476), .A2(n3523), .ZN(n2444) );
  NOR2_X1 U3099 ( .A1(n4476), .A2(n3523), .ZN(n2443) );
  NAND2_X1 U3100 ( .A1(n3827), .A2(REG2_REG_16__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3101 ( .A1(n3828), .A2(REG1_REG_16__SCAN_IN), .ZN(n2447) );
  INV_X1 U3102 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2454) );
  XNOR2_X1 U3103 ( .A(n2456), .B(n2454), .ZN(n3681) );
  OR2_X1 U3104 ( .A1(n2609), .A2(n3681), .ZN(n2446) );
  INV_X1 U3105 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4540) );
  OR2_X1 U3106 ( .A1(n2342), .A2(n4540), .ZN(n2445) );
  NAND2_X1 U3107 ( .A1(n2449), .A2(n2239), .ZN(n2450) );
  NAND2_X1 U3108 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2451) );
  XNOR2_X1 U3109 ( .A(n2451), .B(IR_REG_16__SCAN_IN), .ZN(n4134) );
  INV_X1 U3110 ( .A(DATAI_16_), .ZN(n4689) );
  MUX2_X1 U3111 ( .A(n4690), .B(n4689), .S(n3831), .Z(n3469) );
  OR2_X1 U3112 ( .A1(n4378), .A2(n3469), .ZN(n3882) );
  NAND2_X1 U3113 ( .A1(n4378), .A2(n3469), .ZN(n3885) );
  NAND2_X1 U3114 ( .A1(n3882), .A2(n3885), .ZN(n3461) );
  NAND2_X1 U3115 ( .A1(n3462), .A2(n3461), .ZN(n3460) );
  INV_X1 U3116 ( .A(n3469), .ZN(n3683) );
  NAND2_X1 U3117 ( .A1(n4378), .A2(n3683), .ZN(n2452) );
  NAND2_X1 U3118 ( .A1(n3828), .A2(REG1_REG_17__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3119 ( .A1(n3827), .A2(REG2_REG_17__SCAN_IN), .ZN(n2460) );
  INV_X1 U3120 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4536) );
  OR2_X1 U3121 ( .A1(n2342), .A2(n4536), .ZN(n2459) );
  INV_X1 U3122 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2453) );
  OAI21_X1 U3123 ( .B1(n2456), .B2(n2454), .A(n2453), .ZN(n2457) );
  NAND2_X1 U3124 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2455) );
  NAND2_X1 U3125 ( .A1(n2457), .A2(n2466), .ZN(n4380) );
  OR2_X1 U3126 ( .A1(n2609), .A2(n4380), .ZN(n2458) );
  NAND4_X1 U3127 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3682)
         );
  AND2_X2 U3128 ( .A1(n2425), .A2(n2462), .ZN(n2556) );
  INV_X1 U3129 ( .A(n2556), .ZN(n2472) );
  NAND2_X1 U3130 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2463) );
  XNOR2_X1 U3131 ( .A(n2463), .B(IR_REG_17__SCAN_IN), .ZN(n4138) );
  MUX2_X1 U3132 ( .A(n4138), .B(DATAI_17_), .S(n3831), .Z(n4460) );
  NAND2_X1 U3133 ( .A1(n3682), .A2(n4460), .ZN(n2464) );
  NAND2_X1 U3134 ( .A1(n3828), .A2(REG1_REG_18__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3135 ( .A1(n3827), .A2(REG2_REG_18__SCAN_IN), .ZN(n2470) );
  INV_X1 U3136 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2465) );
  OR2_X1 U3137 ( .A1(n2342), .A2(n2465), .ZN(n2469) );
  INV_X1 U3138 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3732) );
  AND2_X1 U3139 ( .A1(n2466), .A2(n3732), .ZN(n2467) );
  OR2_X1 U3140 ( .A1(n2467), .A2(n2480), .ZN(n4363) );
  OR2_X1 U3141 ( .A1(n2609), .A2(n4363), .ZN(n2468) );
  OR2_X1 U3142 ( .A1(n2472), .A2(IR_REG_17__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3143 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  MUX2_X1 U3144 ( .A(IR_REG_31__SCAN_IN), .B(n2474), .S(IR_REG_18__SCAN_IN), 
        .Z(n2477) );
  INV_X1 U3145 ( .A(n2475), .ZN(n2476) );
  AND2_X1 U3146 ( .A1(n2477), .A2(n2228), .ZN(n4125) );
  INV_X1 U3147 ( .A(DATAI_18_), .ZN(n4685) );
  MUX2_X1 U31480 ( .A(n4686), .B(n4685), .S(n3831), .Z(n4352) );
  OR2_X1 U31490 ( .A1(n4461), .A2(n4352), .ZN(n4326) );
  NAND2_X1 U3150 ( .A1(n4461), .A2(n4352), .ZN(n4327) );
  OR2_X1 U3151 ( .A1(n4461), .A2(n4356), .ZN(n2479) );
  NAND2_X1 U3152 ( .A1(n3828), .A2(REG1_REG_19__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3153 ( .A1(n3827), .A2(REG2_REG_19__SCAN_IN), .ZN(n2484) );
  INV_X1 U3154 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4531) );
  OR2_X1 U3155 ( .A1(n2342), .A2(n4531), .ZN(n2483) );
  NOR2_X1 U3156 ( .A1(n2480), .A2(REG3_REG_19__SCAN_IN), .ZN(n2481) );
  OR2_X1 U3157 ( .A1(n2490), .A2(n2481), .ZN(n4342) );
  OR2_X1 U3158 ( .A1(n2609), .A2(n4342), .ZN(n2482) );
  INV_X1 U3159 ( .A(n2488), .ZN(n2486) );
  NAND2_X1 U3160 ( .A1(n2486), .A2(IR_REG_19__SCAN_IN), .ZN(n2489) );
  MUX2_X1 U3161 ( .A(n4362), .B(DATAI_19_), .S(n3831), .Z(n3648) );
  NOR2_X1 U3162 ( .A1(n4357), .A2(n3648), .ZN(n4305) );
  NAND2_X1 U3163 ( .A1(n4357), .A2(n3648), .ZN(n4306) );
  NAND2_X1 U3164 ( .A1(n3828), .A2(REG1_REG_20__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3165 ( .A1(n3827), .A2(REG2_REG_20__SCAN_IN), .ZN(n2494) );
  OR2_X1 U3166 ( .A1(n2490), .A2(REG3_REG_20__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3167 ( .A1(n2506), .A2(n2491), .ZN(n3711) );
  OR2_X1 U3168 ( .A1(n2609), .A2(n3711), .ZN(n2493) );
  INV_X1 U3169 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4527) );
  OR2_X1 U3170 ( .A1(n2342), .A2(n4527), .ZN(n2492) );
  NAND2_X1 U3171 ( .A1(n3831), .A2(DATAI_20_), .ZN(n4316) );
  NAND2_X1 U3172 ( .A1(n4333), .A2(n4444), .ZN(n3856) );
  OAI21_X1 U3173 ( .B1(n4304), .B2(n4305), .A(n2229), .ZN(n2496) );
  OR2_X1 U3174 ( .A1(n4333), .A2(n4444), .ZN(n3857) );
  NAND2_X1 U3175 ( .A1(n2496), .A2(n3857), .ZN(n4290) );
  NAND2_X1 U3176 ( .A1(n3827), .A2(REG2_REG_21__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3177 ( .A1(n3828), .A2(REG1_REG_21__SCAN_IN), .ZN(n2499) );
  INV_X1 U3178 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3660) );
  XNOR2_X1 U3179 ( .A(n2506), .B(n3660), .ZN(n3659) );
  INV_X1 U3180 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4523) );
  OR2_X1 U3181 ( .A1(n2342), .A2(n4523), .ZN(n2497) );
  NAND2_X1 U3182 ( .A1(n3831), .A2(DATAI_21_), .ZN(n4295) );
  INV_X1 U3183 ( .A(n4295), .ZN(n4435) );
  NAND2_X1 U3184 ( .A1(n4445), .A2(n4435), .ZN(n2501) );
  NAND2_X1 U3185 ( .A1(n4290), .A2(n2501), .ZN(n2503) );
  OR2_X1 U3186 ( .A1(n4445), .A2(n4435), .ZN(n2502) );
  NAND2_X1 U3187 ( .A1(n3828), .A2(REG1_REG_22__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U3188 ( .A1(n3827), .A2(REG2_REG_22__SCAN_IN), .ZN(n2510) );
  INV_X1 U3189 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4093) );
  OR2_X1 U3190 ( .A1(n2342), .A2(n4093), .ZN(n2509) );
  INV_X1 U3191 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2504) );
  OAI21_X1 U3192 ( .B1(n2506), .B2(n3660), .A(n2504), .ZN(n2507) );
  NAND2_X1 U3193 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2505) );
  NAND2_X1 U3194 ( .A1(n2507), .A2(n2515), .ZN(n4274) );
  NAND2_X1 U3195 ( .A1(n3831), .A2(DATAI_22_), .ZN(n4282) );
  NAND2_X1 U3196 ( .A1(n4436), .A2(n4282), .ZN(n2600) );
  NAND2_X1 U3197 ( .A1(n4251), .A2(n2600), .ZN(n4277) );
  INV_X1 U3198 ( .A(n4282), .ZN(n2512) );
  INV_X1 U3199 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U3200 ( .A1(n3828), .A2(REG1_REG_23__SCAN_IN), .ZN(n2514) );
  OAI21_X1 U3201 ( .B1(n2342), .B2(n4514), .A(n2514), .ZN(n2519) );
  INV_X1 U3202 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3641) );
  AND2_X1 U3203 ( .A1(n2515), .A2(n3641), .ZN(n2516) );
  NOR2_X2 U3204 ( .A1(n2515), .A2(n3641), .ZN(n2521) );
  OR2_X1 U3205 ( .A1(n2516), .A2(n2521), .ZN(n4262) );
  NAND2_X1 U3206 ( .A1(n3827), .A2(REG2_REG_23__SCAN_IN), .ZN(n2517) );
  OAI21_X1 U3207 ( .B1(n4262), .B2(n2609), .A(n2517), .ZN(n2518) );
  NAND2_X1 U3208 ( .A1(n3831), .A2(DATAI_23_), .ZN(n4254) );
  NAND2_X1 U3209 ( .A1(n4421), .A2(n4254), .ZN(n2520) );
  NAND2_X1 U32100 ( .A1(n3827), .A2(REG2_REG_24__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32110 ( .A1(n3828), .A2(REG1_REG_24__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32120 ( .A1(n2521), .A2(REG3_REG_24__SCAN_IN), .ZN(n2528) );
  OR2_X1 U32130 ( .A1(n2521), .A2(REG3_REG_24__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32140 ( .A1(n2528), .A2(n2522), .ZN(n3701) );
  OR2_X1 U32150 ( .A1(n3701), .A2(n2609), .ZN(n2524) );
  INV_X1 U32160 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4510) );
  OR2_X1 U32170 ( .A1(n2342), .A2(n4510), .ZN(n2523) );
  INV_X1 U32180 ( .A(n4255), .ZN(n4218) );
  NAND2_X1 U32190 ( .A1(n3831), .A2(DATAI_24_), .ZN(n4241) );
  INV_X1 U32200 ( .A(n4241), .ZN(n4417) );
  NAND2_X1 U32210 ( .A1(n4218), .A2(n4417), .ZN(n2527) );
  INV_X1 U32220 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U32230 ( .A1(n2528), .A2(n3671), .ZN(n2529) );
  NAND2_X1 U32240 ( .A1(n2537), .A2(n2529), .ZN(n3670) );
  OR2_X1 U32250 ( .A1(n3670), .A2(n2609), .ZN(n2533) );
  NAND2_X1 U32260 ( .A1(n3828), .A2(REG1_REG_25__SCAN_IN), .ZN(n2532) );
  INV_X1 U32270 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4506) );
  OR2_X1 U32280 ( .A1(n2342), .A2(n4506), .ZN(n2531) );
  NAND2_X1 U32290 ( .A1(n3827), .A2(REG2_REG_25__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32300 ( .A1(n3831), .A2(DATAI_25_), .ZN(n4221) );
  NAND2_X1 U32310 ( .A1(n4198), .A2(n4221), .ZN(n2536) );
  INV_X1 U32320 ( .A(n4221), .ZN(n2534) );
  INV_X1 U32330 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U32340 ( .A1(n2537), .A2(n3741), .ZN(n2538) );
  NAND2_X1 U32350 ( .A1(n2542), .A2(n2538), .ZN(n3740) );
  INV_X1 U32360 ( .A(n2278), .ZN(n2539) );
  AOI22_X1 U32370 ( .A1(n2539), .A2(REG0_REG_26__SCAN_IN), .B1(n3828), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32380 ( .A1(n3827), .A2(REG2_REG_26__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32390 ( .A1(n3831), .A2(DATAI_26_), .ZN(n4197) );
  NAND2_X1 U32400 ( .A1(n4401), .A2(n4203), .ZN(n3848) );
  INV_X1 U32410 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3630) );
  AND2_X1 U32420 ( .A1(n2542), .A2(n3630), .ZN(n2543) );
  NOR2_X2 U32430 ( .A1(n2542), .A2(n3630), .ZN(n2547) );
  AOI22_X1 U32440 ( .A1(n2539), .A2(REG0_REG_27__SCAN_IN), .B1(n3828), .B2(
        REG1_REG_27__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32450 ( .A1(n3827), .A2(REG2_REG_27__SCAN_IN), .ZN(n2544) );
  INV_X1 U32460 ( .A(n4200), .ZN(n3824) );
  NAND2_X1 U32470 ( .A1(n3831), .A2(DATAI_27_), .ZN(n4186) );
  NAND2_X1 U32480 ( .A1(n3824), .A2(n4186), .ZN(n2546) );
  OR2_X1 U32490 ( .A1(n2547), .A2(REG3_REG_28__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32500 ( .A1(n2547), .A2(REG3_REG_28__SCAN_IN), .ZN(n4157) );
  INV_X1 U32510 ( .A(n2609), .ZN(n2549) );
  INV_X1 U32520 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4494) );
  NAND2_X1 U32530 ( .A1(n3828), .A2(REG1_REG_28__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32540 ( .A1(n3827), .A2(REG2_REG_28__SCAN_IN), .ZN(n2550) );
  OAI211_X1 U32550 ( .C1(n2342), .C2(n4494), .A(n2551), .B(n2550), .ZN(n2552)
         );
  INV_X1 U32560 ( .A(n2552), .ZN(n2553) );
  NAND2_X1 U32570 ( .A1(n3831), .A2(DATAI_28_), .ZN(n4170) );
  INV_X1 U32580 ( .A(n4170), .ZN(n3619) );
  NAND2_X1 U32590 ( .A1(n4404), .A2(n3619), .ZN(n3826) );
  NAND2_X1 U32600 ( .A1(n4161), .A2(n4170), .ZN(n3819) );
  XNOR2_X1 U32610 ( .A(n2655), .B(n2555), .ZN(n4165) );
  NAND2_X1 U32620 ( .A1(n2557), .A2(n2556), .ZN(n2564) );
  INV_X1 U32630 ( .A(IR_REG_22__SCAN_IN), .ZN(n2559) );
  XNOR2_X2 U32640 ( .A(n2560), .B(n2559), .ZN(n2821) );
  XNOR2_X2 U32650 ( .A(n2563), .B(n2562), .ZN(n3911) );
  NAND2_X1 U32660 ( .A1(n2564), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  XNOR2_X1 U32670 ( .A(n3920), .B(n3059), .ZN(n2567) );
  NAND2_X1 U32680 ( .A1(n2567), .A2(n4146), .ZN(n3100) );
  AND2_X1 U32690 ( .A1(n3911), .A2(n4362), .ZN(n3916) );
  INV_X1 U32700 ( .A(n4711), .ZN(n2568) );
  NOR2_X1 U32710 ( .A1(n2569), .A2(n2754), .ZN(n2570) );
  MUX2_X1 U32720 ( .A(n2754), .B(n2570), .S(IR_REG_28__SCAN_IN), .Z(n2571) );
  INV_X1 U32730 ( .A(n2571), .ZN(n2574) );
  INV_X1 U32740 ( .A(n2572), .ZN(n2573) );
  NAND2_X1 U32750 ( .A1(n2574), .A2(n2573), .ZN(n4554) );
  NAND2_X1 U32760 ( .A1(n3920), .A2(n3907), .ZN(n2835) );
  OR2_X1 U32770 ( .A1(n2576), .A2(n2953), .ZN(n2798) );
  INV_X1 U32780 ( .A(n2798), .ZN(n3766) );
  NAND2_X1 U32790 ( .A1(n2862), .A2(n3766), .ZN(n2861) );
  NAND2_X1 U32800 ( .A1(n2861), .A2(n2577), .ZN(n2875) );
  INV_X1 U32810 ( .A(n3863), .ZN(n2876) );
  NAND2_X1 U32820 ( .A1(n2875), .A2(n2876), .ZN(n2874) );
  NAND2_X1 U32830 ( .A1(n2874), .A2(n2578), .ZN(n2977) );
  NAND2_X1 U32840 ( .A1(n3936), .A2(n3094), .ZN(n3768) );
  NAND2_X1 U32850 ( .A1(n3771), .A2(n3768), .ZN(n3868) );
  INV_X1 U32860 ( .A(n3868), .ZN(n2978) );
  NAND2_X1 U32870 ( .A1(n2977), .A2(n2978), .ZN(n2976) );
  INV_X1 U32880 ( .A(n3772), .ZN(n2579) );
  AND2_X1 U32890 ( .A1(n3935), .A2(n3001), .ZN(n3016) );
  OR2_X1 U32900 ( .A1(n3935), .A2(n3001), .ZN(n3788) );
  NAND2_X1 U32910 ( .A1(n3934), .A2(n3083), .ZN(n3790) );
  NAND2_X1 U32920 ( .A1(n3075), .A2(n3790), .ZN(n2581) );
  OR2_X1 U32930 ( .A1(n3934), .A2(n3083), .ZN(n3777) );
  INV_X1 U32940 ( .A(n2582), .ZN(n2583) );
  OAI21_X1 U32950 ( .B1(n3114), .B2(n2583), .A(n3787), .ZN(n3230) );
  OR2_X1 U32960 ( .A1(n3932), .A2(n3227), .ZN(n3780) );
  NAND2_X1 U32970 ( .A1(n3230), .A2(n3780), .ZN(n2584) );
  NAND2_X1 U32980 ( .A1(n3932), .A2(n3227), .ZN(n3791) );
  INV_X1 U32990 ( .A(n3214), .ZN(n3221) );
  AND2_X1 U33000 ( .A1(n3931), .A2(n3221), .ZN(n3785) );
  OR2_X1 U33010 ( .A1(n3931), .A2(n3221), .ZN(n3781) );
  NAND2_X1 U33020 ( .A1(n3930), .A2(n3291), .ZN(n3798) );
  OR2_X1 U33030 ( .A1(n3930), .A2(n3291), .ZN(n3797) );
  NAND2_X1 U33040 ( .A1(n3928), .A2(n3379), .ZN(n3362) );
  NAND2_X1 U33050 ( .A1(n3927), .A2(n3428), .ZN(n2586) );
  NAND2_X1 U33060 ( .A1(n3362), .A2(n2586), .ZN(n2588) );
  INV_X1 U33070 ( .A(n2587), .ZN(n3326) );
  NOR2_X1 U33080 ( .A1(n2588), .A2(n3326), .ZN(n3799) );
  INV_X1 U33090 ( .A(n2588), .ZN(n2591) );
  OR2_X1 U33100 ( .A1(n3928), .A2(n3379), .ZN(n3361) );
  NAND2_X1 U33110 ( .A1(n3327), .A2(n3361), .ZN(n2590) );
  NOR2_X1 U33120 ( .A1(n3927), .A2(n3428), .ZN(n2589) );
  AOI21_X1 U33130 ( .B1(n2591), .B2(n2590), .A(n2589), .ZN(n3802) );
  INV_X1 U33140 ( .A(n3397), .ZN(n3872) );
  INV_X1 U33150 ( .A(n3523), .ZN(n3756) );
  OR2_X1 U33160 ( .A1(n4476), .A2(n3756), .ZN(n3803) );
  NAND2_X1 U33170 ( .A1(n4476), .A2(n3756), .ZN(n3784) );
  NAND2_X1 U33180 ( .A1(n3803), .A2(n3784), .ZN(n3861) );
  INV_X1 U33190 ( .A(n3804), .ZN(n2592) );
  NAND2_X1 U33200 ( .A1(n2593), .A2(n3784), .ZN(n3463) );
  INV_X1 U33210 ( .A(n3461), .ZN(n3874) );
  AND2_X1 U33220 ( .A1(n3682), .A2(n4386), .ZN(n3807) );
  INV_X1 U33230 ( .A(n3648), .ZN(n4339) );
  NAND2_X1 U33240 ( .A1(n4357), .A2(n4339), .ZN(n2594) );
  OR2_X1 U33250 ( .A1(n3682), .A2(n4386), .ZN(n4324) );
  NAND2_X1 U33260 ( .A1(n4326), .A2(n4324), .ZN(n2596) );
  NOR2_X1 U33270 ( .A1(n4357), .A2(n4339), .ZN(n2595) );
  AOI21_X1 U33280 ( .B1(n2082), .B2(n2596), .A(n2595), .ZN(n4300) );
  OR2_X1 U33290 ( .A1(n4333), .A2(n4316), .ZN(n2597) );
  NAND2_X1 U33300 ( .A1(n4301), .A2(n3888), .ZN(n2598) );
  NAND2_X1 U33310 ( .A1(n4333), .A2(n4316), .ZN(n3810) );
  NAND2_X1 U33320 ( .A1(n2598), .A2(n3810), .ZN(n4287) );
  OR2_X1 U33330 ( .A1(n4445), .A2(n4295), .ZN(n4249) );
  NAND2_X1 U33340 ( .A1(n4251), .A2(n4249), .ZN(n3891) );
  INV_X1 U33350 ( .A(n3891), .ZN(n2599) );
  NAND2_X1 U33360 ( .A1(n4287), .A2(n2599), .ZN(n2604) );
  NAND2_X1 U33370 ( .A1(n4279), .A2(n4254), .ZN(n2601) );
  NAND2_X1 U33380 ( .A1(n2601), .A2(n2600), .ZN(n3813) );
  INV_X1 U33390 ( .A(n3813), .ZN(n2603) );
  AND2_X1 U33400 ( .A1(n4445), .A2(n4295), .ZN(n4248) );
  NAND2_X1 U33410 ( .A1(n4248), .A2(n4251), .ZN(n2602) );
  AND2_X1 U33420 ( .A1(n2603), .A2(n2602), .ZN(n3890) );
  NAND2_X1 U33430 ( .A1(n2604), .A2(n3890), .ZN(n4230) );
  NAND2_X1 U33440 ( .A1(n4421), .A2(n4259), .ZN(n4229) );
  NAND2_X1 U33450 ( .A1(n4255), .A2(n4417), .ZN(n3847) );
  OR2_X1 U33460 ( .A1(n4255), .A2(n4417), .ZN(n4212) );
  NAND2_X1 U33470 ( .A1(n4418), .A2(n4221), .ZN(n3846) );
  NAND2_X1 U33480 ( .A1(n4212), .A2(n3846), .ZN(n3893) );
  INV_X1 U33490 ( .A(n3893), .ZN(n3816) );
  NAND2_X1 U33500 ( .A1(n4213), .A2(n3816), .ZN(n4194) );
  OR2_X1 U33510 ( .A1(n4401), .A2(n4197), .ZN(n2605) );
  OR2_X1 U33520 ( .A1(n4418), .A2(n4221), .ZN(n4193) );
  AND2_X1 U3353 ( .A1(n2605), .A2(n4193), .ZN(n3815) );
  NAND2_X1 U33540 ( .A1(n4401), .A2(n4197), .ZN(n3820) );
  XNOR2_X1 U3355 ( .A(n4200), .B(n4399), .ZN(n4181) );
  INV_X1 U3356 ( .A(n4181), .ZN(n4176) );
  OR2_X1 U3357 ( .A1(n4200), .A2(n4186), .ZN(n3825) );
  XNOR2_X1 U3358 ( .A(n2658), .B(n3851), .ZN(n2608) );
  NAND2_X1 U3359 ( .A1(n3920), .A2(n4362), .ZN(n2607) );
  INV_X1 U3360 ( .A(n3911), .ZN(n2747) );
  NAND2_X1 U3361 ( .A1(n2747), .A2(n3907), .ZN(n2606) );
  NAND2_X1 U3362 ( .A1(n2608), .A2(n4370), .ZN(n4175) );
  INV_X1 U3363 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2671) );
  OR2_X1 U3364 ( .A1(n4157), .A2(n2609), .ZN(n2611) );
  AOI22_X1 U3365 ( .A1(REG1_REG_29__SCAN_IN), .A2(n3828), .B1(n3827), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n2610) );
  OAI211_X1 U3366 ( .C1(n2342), .C2(n2671), .A(n2611), .B(n2610), .ZN(n4166)
         );
  INV_X1 U3367 ( .A(n2835), .ZN(n2680) );
  AND2_X2 U3368 ( .A1(n4554), .A2(n2680), .ZN(n4475) );
  AOI22_X1 U3369 ( .A1(n4166), .A2(n4475), .B1(n4473), .B2(n3619), .ZN(n2612)
         );
  OAI211_X1 U3370 ( .C1(n3824), .C2(n4478), .A(n4175), .B(n2612), .ZN(n2613)
         );
  AOI21_X1 U3371 ( .B1(n4165), .B2(n4713), .A(n2613), .ZN(n4493) );
  AND2_X1 U3372 ( .A1(n2425), .A2(n2614), .ZN(n2615) );
  NOR2_X1 U3373 ( .A1(n2615), .A2(n2754), .ZN(n2616) );
  MUX2_X1 U3374 ( .A(n2754), .B(n2616), .S(IR_REG_25__SCAN_IN), .Z(n2617) );
  INV_X1 U3375 ( .A(n2617), .ZN(n2619) );
  NAND2_X1 U3376 ( .A1(n2619), .A2(n2618), .ZN(n2630) );
  NAND2_X1 U3377 ( .A1(n2630), .A2(B_REG_SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3378 ( .A1(n2425), .A2(n2620), .ZN(n2621) );
  NAND2_X1 U3379 ( .A1(n2623), .A2(n2622), .ZN(n2632) );
  NAND2_X1 U3380 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2624) );
  MUX2_X1 U3381 ( .A(n2625), .B(B_REG_SCAN_IN), .S(n2739), .Z(n2629) );
  NAND2_X1 U3382 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2626) );
  MUX2_X1 U3383 ( .A(IR_REG_31__SCAN_IN), .B(n2626), .S(IR_REG_26__SCAN_IN), 
        .Z(n2628) );
  INV_X1 U3384 ( .A(D_REG_1__SCAN_IN), .ZN(n4078) );
  NAND2_X1 U3385 ( .A1(n2758), .A2(n4078), .ZN(n2831) );
  INV_X1 U3386 ( .A(n2734), .ZN(n2649) );
  NAND2_X1 U3387 ( .A1(n2630), .A2(n2649), .ZN(n2829) );
  NAND2_X1 U3388 ( .A1(n2831), .A2(n2829), .ZN(n2647) );
  INV_X1 U3389 ( .A(n2630), .ZN(n2742) );
  NAND2_X1 U3390 ( .A1(n2631), .A2(IR_REG_23__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3391 ( .A1(n2633), .A2(n2632), .ZN(n2896) );
  NAND2_X1 U3392 ( .A1(n2897), .A2(n4683), .ZN(n3053) );
  NAND2_X1 U3393 ( .A1(n4711), .A2(n2634), .ZN(n2846) );
  AND2_X1 U3394 ( .A1(n3911), .A2(n4146), .ZN(n2834) );
  NAND2_X1 U3395 ( .A1(n2846), .A2(n3055), .ZN(n2635) );
  NOR2_X1 U3396 ( .A1(n3053), .A2(n2635), .ZN(n2646) );
  NOR4_X1 U3397 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2639) );
  NOR4_X1 U3398 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2638) );
  NOR4_X1 U3399 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2637) );
  NOR4_X1 U3400 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2636) );
  NAND4_X1 U3401 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n2645)
         );
  NOR2_X1 U3402 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_25__SCAN_IN), .ZN(n2643)
         );
  NOR4_X1 U3403 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2642) );
  NOR4_X1 U3404 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2641) );
  NOR4_X1 U3405 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2640) );
  NAND4_X1 U3406 ( .A1(n2643), .A2(n2642), .A3(n2641), .A4(n2640), .ZN(n2644)
         );
  OAI21_X1 U3407 ( .B1(n2645), .B2(n2644), .A(n2758), .ZN(n2830) );
  INV_X1 U3408 ( .A(D_REG_0__SCAN_IN), .ZN(n3964) );
  INV_X1 U3409 ( .A(n2739), .ZN(n2648) );
  AND2_X2 U3410 ( .A1(n2670), .A2(n2832), .ZN(n4727) );
  MUX2_X1 U3411 ( .A(n2650), .B(n4493), .S(n4727), .Z(n2654) );
  NAND2_X1 U3412 ( .A1(n3161), .A2(n2953), .ZN(n2982) );
  NAND2_X1 U3413 ( .A1(n2983), .A2(n3094), .ZN(n2651) );
  INV_X1 U3414 ( .A(n2672), .ZN(n2652) );
  OAI21_X1 U3415 ( .B1(n4182), .B2(n4170), .A(n2652), .ZN(n4496) );
  INV_X1 U3416 ( .A(n2833), .ZN(n2799) );
  AND2_X2 U3417 ( .A1(n2799), .A2(n3911), .ZN(n4351) );
  NAND2_X1 U3418 ( .A1(n2654), .A2(n2653), .ZN(U3546) );
  NAND2_X1 U3419 ( .A1(n3831), .A2(DATAI_29_), .ZN(n4163) );
  XOR2_X1 U3420 ( .A(n4163), .B(n4166), .Z(n3852) );
  XNOR2_X1 U3421 ( .A(n2656), .B(n3852), .ZN(n4164) );
  INV_X1 U3422 ( .A(n3826), .ZN(n2657) );
  AOI21_X1 U3423 ( .B1(n2658), .B2(n3819), .A(n2657), .ZN(n2659) );
  XNOR2_X1 U3424 ( .A(n2659), .B(n3852), .ZN(n2667) );
  NAND2_X1 U3425 ( .A1(n3828), .A2(REG1_REG_30__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3426 ( .A1(n3827), .A2(REG2_REG_30__SCAN_IN), .ZN(n2662) );
  INV_X1 U3427 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2660) );
  OR2_X1 U3428 ( .A1(n2342), .A2(n2660), .ZN(n2661) );
  AND3_X1 U3429 ( .A1(n2663), .A2(n2662), .A3(n2661), .ZN(n3836) );
  INV_X1 U3430 ( .A(B_REG_SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3431 ( .A1(n2665), .A2(n2664), .ZN(n2703) );
  OAI21_X1 U3432 ( .B1(n2666), .B2(n2703), .A(n4475), .ZN(n4152) );
  OAI22_X1 U3433 ( .A1(n4404), .A2(n4478), .B1(n4163), .B2(n4331), .ZN(n2668)
         );
  INV_X1 U3434 ( .A(n2832), .ZN(n3057) );
  AND2_X2 U3435 ( .A1(n2670), .A2(n3057), .ZN(n4719) );
  INV_X1 U3436 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2675) );
  MUX2_X1 U3437 ( .A(n2675), .B(n2674), .S(n4727), .Z(n2677) );
  NAND2_X1 U3438 ( .A1(n2677), .A2(n2676), .ZN(U3547) );
  INV_X1 U3439 ( .A(n4683), .ZN(n2678) );
  OR2_X1 U3440 ( .A1(n2897), .A2(n2678), .ZN(n3925) );
  INV_X2 U3441 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3442 ( .A(n2896), .ZN(n2679) );
  NAND2_X1 U3443 ( .A1(n2679), .A2(STATE_REG_SCAN_IN), .ZN(n3923) );
  NAND2_X1 U3444 ( .A1(n3053), .A2(n3923), .ZN(n2685) );
  NAND2_X1 U3445 ( .A1(n2680), .A2(n2896), .ZN(n2681) );
  NAND2_X1 U3446 ( .A1(n3831), .A2(n2681), .ZN(n2683) );
  INV_X1 U3447 ( .A(n4650), .ZN(n4635) );
  INV_X1 U3448 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n3942) );
  NOR2_X1 U3449 ( .A1(n4635), .A2(n3942), .ZN(n2694) );
  NAND2_X1 U3450 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2687) );
  INV_X1 U3451 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2769) );
  NOR3_X1 U3452 ( .A1(n2686), .A2(n4699), .A3(n2769), .ZN(n2714) );
  INV_X1 U3453 ( .A(n2683), .ZN(n2684) );
  NAND2_X1 U3454 ( .A1(n2685), .A2(n2684), .ZN(n2772) );
  INV_X1 U3455 ( .A(n2703), .ZN(n4549) );
  OR2_X1 U3456 ( .A1(n2772), .A2(n4549), .ZN(n4627) );
  AOI211_X1 U3457 ( .C1(n2687), .C2(n2686), .A(n2714), .B(n4627), .ZN(n2693)
         );
  NAND2_X1 U34580 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n2704) );
  INV_X1 U34590 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2688) );
  MUX2_X1 U3460 ( .A(REG2_REG_1__SCAN_IN), .B(n2688), .S(n2723), .Z(n2690) );
  INV_X1 U3461 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2689) );
  OR2_X1 U3462 ( .A1(n4554), .A2(n2703), .ZN(n3918) );
  NOR2_X1 U3463 ( .A1(n3918), .A2(n2772), .ZN(n4631) );
  INV_X1 U3464 ( .A(n4631), .ZN(n4646) );
  AOI211_X1 U3465 ( .C1(n2704), .C2(n2690), .A(n2711), .B(n4646), .ZN(n2692)
         );
  INV_X1 U3466 ( .A(n4554), .ZN(n2850) );
  OAI22_X1 U34670 ( .A1(n4657), .A2(n2055), .B1(STATE_REG_SCAN_IN), .B2(n3160), 
        .ZN(n2691) );
  OR4_X1 U3468 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(U3241) );
  NOR2_X1 U34690 ( .A1(n2703), .A2(REG2_REG_0__SCAN_IN), .ZN(n2695) );
  NOR2_X1 U3470 ( .A1(n4554), .A2(n2695), .ZN(n2767) );
  INV_X1 U34710 ( .A(n3059), .ZN(n2696) );
  NAND2_X1 U3472 ( .A1(n2576), .A2(n2994), .ZN(n2698) );
  AND2_X4 U34730 ( .A1(n2897), .A2(n3059), .ZN(n3610) );
  NAND2_X1 U3474 ( .A1(n2867), .A2(n3610), .ZN(n2697) );
  NAND2_X1 U34750 ( .A1(n2698), .A2(n2697), .ZN(n2825) );
  NOR2_X1 U3476 ( .A1(n2897), .A2(n2769), .ZN(n2699) );
  OR2_X1 U34770 ( .A1(n2825), .A2(n2699), .ZN(n2828) );
  NAND2_X1 U3478 ( .A1(n2576), .A2(n2058), .ZN(n2702) );
  INV_X1 U34790 ( .A(n2897), .ZN(n2700) );
  AOI22_X1 U3480 ( .A1(n2867), .A2(n2994), .B1(IR_REG_0__SCAN_IN), .B2(n2700), 
        .ZN(n2701) );
  NAND2_X1 U34810 ( .A1(n2702), .A2(n2701), .ZN(n2827) );
  XNOR2_X1 U3482 ( .A(n2828), .B(n2827), .ZN(n2957) );
  NAND3_X1 U34830 ( .A1(n2957), .A2(n2850), .A3(n2703), .ZN(n2707) );
  OAI21_X1 U3484 ( .B1(n3918), .B2(n2704), .A(U4043), .ZN(n2705) );
  INV_X1 U34850 ( .A(n2705), .ZN(n2706) );
  OAI211_X1 U3486 ( .C1(IR_REG_0__SCAN_IN), .C2(n2767), .A(n2707), .B(n2706), 
        .ZN(n2795) );
  INV_X1 U34870 ( .A(n2795), .ZN(n2722) );
  NOR2_X1 U3488 ( .A1(n2055), .A2(n2688), .ZN(n2710) );
  INV_X1 U34890 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2708) );
  MUX2_X1 U3490 ( .A(n2708), .B(REG2_REG_2__SCAN_IN), .S(n2775), .Z(n2709) );
  INV_X1 U34910 ( .A(n2774), .ZN(n2713) );
  NOR3_X1 U3492 ( .A1(n2711), .A2(n2710), .A3(n2709), .ZN(n2712) );
  NOR3_X1 U34930 ( .A1(n4646), .A2(n2713), .A3(n2712), .ZN(n2721) );
  INV_X1 U3494 ( .A(n2055), .ZN(n2715) );
  XOR2_X1 U34950 ( .A(REG1_REG_2__SCAN_IN), .B(n2775), .Z(n2716) );
  NOR2_X1 U3496 ( .A1(n2717), .A2(n2716), .ZN(n2776) );
  AOI211_X1 U34970 ( .C1(n2717), .C2(n2716), .A(n2776), .B(n4627), .ZN(n2720)
         );
  AOI22_X1 U3498 ( .A1(n4650), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2718) );
  OAI21_X1 U34990 ( .B1(n4657), .B2(n2775), .A(n2718), .ZN(n2719) );
  OR4_X1 U3500 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .ZN(U3242) );
  MUX2_X1 U35010 ( .A(n2055), .B(n2263), .S(U3149), .Z(n2724) );
  INV_X1 U3502 ( .A(n2724), .ZN(U3351) );
  MUX2_X1 U35030 ( .A(n2725), .B(n2791), .S(STATE_REG_SCAN_IN), .Z(n2726) );
  INV_X1 U3504 ( .A(n2726), .ZN(U3348) );
  INV_X1 U35050 ( .A(DATAI_3_), .ZN(n2727) );
  MUX2_X1 U35060 ( .A(n2727), .B(n2211), .S(STATE_REG_SCAN_IN), .Z(n2728) );
  INV_X1 U35070 ( .A(n2728), .ZN(U3349) );
  INV_X1 U35080 ( .A(DATAI_5_), .ZN(n2729) );
  MUX2_X1 U35090 ( .A(n2130), .B(n2729), .S(U3149), .Z(n2730) );
  INV_X1 U35100 ( .A(n2730), .ZN(U3347) );
  MUX2_X1 U35110 ( .A(n2349), .B(n2971), .S(STATE_REG_SCAN_IN), .Z(n2731) );
  INV_X1 U35120 ( .A(n2731), .ZN(U3345) );
  INV_X1 U35130 ( .A(DATAI_13_), .ZN(n2733) );
  NAND2_X1 U35140 ( .A1(n4115), .A2(STATE_REG_SCAN_IN), .ZN(n2732) );
  OAI21_X1 U35150 ( .B1(STATE_REG_SCAN_IN), .B2(n2733), .A(n2732), .ZN(U3339)
         );
  INV_X1 U35160 ( .A(DATAI_26_), .ZN(n2736) );
  NAND2_X1 U35170 ( .A1(n2734), .A2(STATE_REG_SCAN_IN), .ZN(n2735) );
  OAI21_X1 U35180 ( .B1(STATE_REG_SCAN_IN), .B2(n2736), .A(n2735), .ZN(U3326)
         );
  INV_X1 U35190 ( .A(DATAI_21_), .ZN(n2738) );
  NAND2_X1 U35200 ( .A1(n3907), .A2(STATE_REG_SCAN_IN), .ZN(n2737) );
  OAI21_X1 U35210 ( .B1(STATE_REG_SCAN_IN), .B2(n2738), .A(n2737), .ZN(U3331)
         );
  INV_X1 U35220 ( .A(DATAI_24_), .ZN(n2741) );
  NAND2_X1 U35230 ( .A1(n2739), .A2(STATE_REG_SCAN_IN), .ZN(n2740) );
  OAI21_X1 U35240 ( .B1(STATE_REG_SCAN_IN), .B2(n2741), .A(n2740), .ZN(U3328)
         );
  INV_X1 U35250 ( .A(DATAI_25_), .ZN(n2744) );
  NAND2_X1 U35260 ( .A1(n2742), .A2(STATE_REG_SCAN_IN), .ZN(n2743) );
  OAI21_X1 U35270 ( .B1(STATE_REG_SCAN_IN), .B2(n2744), .A(n2743), .ZN(U3327)
         );
  INV_X1 U35280 ( .A(DATAI_22_), .ZN(n2746) );
  NAND2_X1 U35290 ( .A1(n3920), .A2(STATE_REG_SCAN_IN), .ZN(n2745) );
  OAI21_X1 U35300 ( .B1(STATE_REG_SCAN_IN), .B2(n2746), .A(n2745), .ZN(U3330)
         );
  INV_X1 U35310 ( .A(DATAI_20_), .ZN(n2749) );
  NAND2_X1 U35320 ( .A1(n2747), .A2(STATE_REG_SCAN_IN), .ZN(n2748) );
  OAI21_X1 U35330 ( .B1(STATE_REG_SCAN_IN), .B2(n2749), .A(n2748), .ZN(U3332)
         );
  INV_X1 U35340 ( .A(DATAI_19_), .ZN(n2750) );
  MUX2_X1 U35350 ( .A(n4146), .B(n2750), .S(U3149), .Z(n2751) );
  INV_X1 U35360 ( .A(n2751), .ZN(U3333) );
  INV_X1 U35370 ( .A(DATAI_29_), .ZN(n4059) );
  NAND2_X1 U35380 ( .A1(n2752), .A2(STATE_REG_SCAN_IN), .ZN(n2753) );
  OAI21_X1 U35390 ( .B1(STATE_REG_SCAN_IN), .B2(n4059), .A(n2753), .ZN(U3323)
         );
  INV_X1 U35400 ( .A(DATAI_31_), .ZN(n2757) );
  OR4_X1 U35410 ( .A1(n2755), .A2(IR_REG_30__SCAN_IN), .A3(n2754), .A4(U3149), 
        .ZN(n2756) );
  OAI21_X1 U35420 ( .B1(STATE_REG_SCAN_IN), .B2(n2757), .A(n2756), .ZN(U3321)
         );
  INV_X1 U35430 ( .A(n2758), .ZN(n2759) );
  AOI22_X1 U35440 ( .A1(n4682), .A2(n3964), .B1(n2760), .B2(n4683), .ZN(U3458)
         );
  INV_X1 U35450 ( .A(n2829), .ZN(n2761) );
  AOI22_X1 U35460 ( .A1(n4682), .A2(n4078), .B1(n2761), .B2(n4683), .ZN(U3459)
         );
  NOR2_X1 U35470 ( .A1(n4650), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U35480 ( .A1(n3925), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2762) );
  OAI21_X1 U35490 ( .B1(n3836), .B2(n3925), .A(n2762), .ZN(U3580) );
  INV_X2 U35500 ( .A(n3925), .ZN(U4043) );
  INV_X1 U35510 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U35520 ( .A1(n3127), .A2(U4043), .ZN(n2763) );
  OAI21_X1 U35530 ( .B1(U4043), .B2(n2764), .A(n2763), .ZN(U3554) );
  INV_X1 U35540 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4057) );
  NAND2_X1 U35550 ( .A1(n3682), .A2(U4043), .ZN(n2765) );
  OAI21_X1 U35560 ( .B1(U4043), .B2(n4057), .A(n2765), .ZN(U3567) );
  INV_X1 U35570 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3953) );
  NAND2_X1 U35580 ( .A1(n3452), .A2(U4043), .ZN(n2766) );
  OAI21_X1 U35590 ( .B1(U4043), .B2(n3953), .A(n2766), .ZN(U3564) );
  OAI21_X1 U35600 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4549), .A(n2767), .ZN(n2768) );
  MUX2_X1 U35610 ( .A(n2768), .B(n2767), .S(IR_REG_0__SCAN_IN), .Z(n2773) );
  AOI22_X1 U35620 ( .A1(n4650), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2771) );
  NAND3_X1 U35630 ( .A1(n4652), .A2(IR_REG_0__SCAN_IN), .A3(n2769), .ZN(n2770)
         );
  OAI211_X1 U35640 ( .C1(n2773), .C2(n2772), .A(n2771), .B(n2770), .ZN(U3240)
         );
  INV_X1 U35650 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3093) );
  XNOR2_X1 U35660 ( .A(n2785), .B(n3093), .ZN(n2780) );
  INV_X1 U35670 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2778) );
  INV_X1 U35680 ( .A(n2775), .ZN(n4552) );
  AOI211_X1 U35690 ( .C1(n2778), .C2(n2777), .A(n2788), .B(n4627), .ZN(n2779)
         );
  AOI21_X1 U35700 ( .B1(n4631), .B2(n2780), .A(n2779), .ZN(n2782) );
  AOI22_X1 U35710 ( .A1(n4650), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2781) );
  OAI211_X1 U35720 ( .C1(n2211), .C2(n4657), .A(n2782), .B(n2781), .ZN(U3243)
         );
  INV_X1 U35730 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U35740 ( .A1(n4333), .A2(U4043), .ZN(n2783) );
  OAI21_X1 U35750 ( .B1(U4043), .B2(n2784), .A(n2783), .ZN(U3570) );
  XNOR2_X1 U35760 ( .A(n2811), .B(n2791), .ZN(n2810) );
  XOR2_X1 U35770 ( .A(REG2_REG_4__SCAN_IN), .B(n2810), .Z(n2797) );
  INV_X1 U35780 ( .A(n4657), .ZN(n2890) );
  INV_X1 U35790 ( .A(n2791), .ZN(n2813) );
  AND2_X1 U35800 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2935) );
  INV_X1 U35810 ( .A(n2935), .ZN(n2786) );
  OAI21_X1 U3582 ( .B1(n4635), .B2(n3941), .A(n2786), .ZN(n2794) );
  INV_X1 U3583 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4720) );
  INV_X1 U3584 ( .A(n2787), .ZN(n2789) );
  XNOR2_X1 U3585 ( .A(n2805), .B(n2791), .ZN(n2792) );
  NOR2_X1 U3586 ( .A1(n2792), .A2(n4720), .ZN(n2806) );
  AOI211_X1 U3587 ( .C1(n4720), .C2(n2792), .A(n4627), .B(n2806), .ZN(n2793)
         );
  AOI211_X1 U3588 ( .C1(n2890), .C2(n2813), .A(n2794), .B(n2793), .ZN(n2796)
         );
  OAI211_X1 U3589 ( .C1(n2797), .C2(n4646), .A(n2796), .B(n2795), .ZN(U3244)
         );
  NAND2_X1 U3590 ( .A1(n2576), .A2(n2953), .ZN(n3765) );
  NAND2_X1 U3591 ( .A1(n2798), .A2(n3765), .ZN(n3860) );
  NAND2_X1 U3592 ( .A1(n2867), .A2(n2799), .ZN(n3106) );
  INV_X1 U3593 ( .A(n3106), .ZN(n2801) );
  INV_X1 U3594 ( .A(n4475), .ZN(n4403) );
  INV_X1 U3595 ( .A(n3100), .ZN(n3400) );
  OAI21_X1 U3596 ( .B1(n3400), .B2(n4370), .A(n3860), .ZN(n2800) );
  OAI21_X1 U3597 ( .B1(n2265), .B2(n4403), .A(n2800), .ZN(n3108) );
  AOI211_X1 U3598 ( .C1(n4711), .C2(n3860), .A(n2801), .B(n3108), .ZN(n4700)
         );
  NAND2_X1 U3599 ( .A1(n4724), .A2(REG1_REG_0__SCAN_IN), .ZN(n2802) );
  OAI21_X1 U3600 ( .B1(n4700), .B2(n4724), .A(n2802), .ZN(U3518) );
  INV_X1 U3601 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3602 ( .A1(n4279), .A2(U4043), .ZN(n2803) );
  OAI21_X1 U3603 ( .B1(U4043), .B2(n2804), .A(n2803), .ZN(U3573) );
  INV_X1 U3604 ( .A(n2805), .ZN(n2807) );
  XNOR2_X1 U3605 ( .A(n2886), .B(REG1_REG_5__SCAN_IN), .ZN(n2808) );
  AOI211_X1 U3606 ( .C1(n2809), .C2(n2808), .A(n4627), .B(n2885), .ZN(n2818)
         );
  INV_X1 U3607 ( .A(n2811), .ZN(n2812) );
  MUX2_X1 U3608 ( .A(n2129), .B(REG2_REG_5__SCAN_IN), .S(n2886), .Z(n2814) );
  AOI211_X1 U3609 ( .C1(n2088), .C2(n2814), .A(n2882), .B(n4646), .ZN(n2817)
         );
  AND2_X1 U3610 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3003) );
  AOI21_X1 U3611 ( .B1(n4650), .B2(ADDR_REG_5__SCAN_IN), .A(n3003), .ZN(n2815)
         );
  OAI21_X1 U3612 ( .B1(n4657), .B2(n2130), .A(n2815), .ZN(n2816) );
  OR3_X1 U3613 ( .A1(n2818), .A2(n2817), .A3(n2816), .ZN(U3245) );
  NAND2_X1 U3614 ( .A1(n2823), .A2(n2994), .ZN(n2820) );
  NAND2_X1 U3615 ( .A1(n2264), .A2(n3610), .ZN(n2819) );
  NAND2_X1 U3616 ( .A1(n2820), .A2(n2819), .ZN(n2822) );
  NAND2_X4 U3617 ( .A1(n2841), .A2(n3059), .ZN(n3597) );
  XNOR2_X1 U3618 ( .A(n2822), .B(n3597), .ZN(n2902) );
  INV_X1 U3619 ( .A(n2904), .ZN(n2824) );
  XNOR2_X1 U3620 ( .A(n2902), .B(n2824), .ZN(n2905) );
  INV_X1 U3621 ( .A(n2825), .ZN(n2826) );
  AOI22_X1 U3622 ( .A1(n2828), .A2(n2827), .B1(n2826), .B2(n3613), .ZN(n2906)
         );
  XNOR2_X1 U3623 ( .A(n2905), .B(n2906), .ZN(n2856) );
  AND2_X1 U3624 ( .A1(n2830), .A2(n2829), .ZN(n3056) );
  OR2_X1 U3625 ( .A1(n2834), .A2(n2833), .ZN(n2836) );
  NAND2_X1 U3626 ( .A1(n2836), .A2(n2835), .ZN(n2838) );
  NOR2_X1 U3627 ( .A1(n3053), .A2(n2838), .ZN(n2837) );
  INV_X1 U3628 ( .A(n2852), .ZN(n2845) );
  NAND2_X1 U3629 ( .A1(n2838), .A2(n4331), .ZN(n2839) );
  NAND2_X1 U3630 ( .A1(n2845), .A2(n2839), .ZN(n2840) );
  NAND2_X1 U3631 ( .A1(n2840), .A2(n3055), .ZN(n2899) );
  INV_X1 U3632 ( .A(n2899), .ZN(n2844) );
  INV_X4 U3633 ( .A(n3615), .ZN(n3609) );
  INV_X1 U3634 ( .A(n2841), .ZN(n2842) );
  AND2_X1 U3635 ( .A1(n4683), .A2(n2842), .ZN(n2843) );
  NAND2_X1 U3636 ( .A1(n2845), .A2(n3917), .ZN(n2900) );
  NAND3_X1 U3637 ( .A1(n2844), .A2(n2848), .A3(n2900), .ZN(n2955) );
  NOR3_X1 U3638 ( .A1(n2845), .A2(n4331), .A3(n3053), .ZN(n2849) );
  INV_X1 U3639 ( .A(n2846), .ZN(n2847) );
  NAND3_X1 U3640 ( .A1(n2852), .A2(n2850), .A3(n3917), .ZN(n3754) );
  INV_X1 U3641 ( .A(n3754), .ZN(n3719) );
  AND2_X1 U3642 ( .A1(n3917), .A2(n4554), .ZN(n2851) );
  NAND2_X1 U3643 ( .A1(n2852), .A2(n2851), .ZN(n3742) );
  AOI22_X1 U3644 ( .A1(n3719), .A2(n2576), .B1(n3759), .B2(n2288), .ZN(n2853)
         );
  OAI21_X1 U3645 ( .B1(n2054), .B2(n3161), .A(n2853), .ZN(n2854) );
  AOI21_X1 U3646 ( .B1(REG3_REG_1__SCAN_IN), .B2(n2955), .A(n2854), .ZN(n2855)
         );
  OAI21_X1 U3647 ( .B1(n2856), .B2(n3747), .A(n2855), .ZN(U3219) );
  INV_X1 U3648 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U3649 ( .A1(n4418), .A2(U4043), .ZN(n2857) );
  OAI21_X1 U3650 ( .B1(U4043), .B2(n3938), .A(n2857), .ZN(U3575) );
  OAI21_X1 U3651 ( .B1(n2575), .B2(n2859), .A(n2858), .ZN(n3169) );
  INV_X1 U3652 ( .A(n3169), .ZN(n2866) );
  INV_X1 U3653 ( .A(n2576), .ZN(n3163) );
  AOI22_X1 U3654 ( .A1(n2288), .A2(n4475), .B1(n4473), .B2(n2264), .ZN(n2860)
         );
  OAI21_X1 U3655 ( .B1(n3163), .B2(n4478), .A(n2860), .ZN(n2865) );
  OAI21_X1 U3656 ( .B1(n2862), .B2(n3766), .A(n2861), .ZN(n2863) );
  NAND2_X1 U3657 ( .A1(n2863), .A2(n4370), .ZN(n2864) );
  OAI21_X1 U3658 ( .B1(n3169), .B2(n3100), .A(n2864), .ZN(n3158) );
  AOI211_X1 U3659 ( .C1(n4711), .C2(n2866), .A(n2865), .B(n3158), .ZN(n2960)
         );
  INV_X1 U3660 ( .A(n4486), .ZN(n3023) );
  NAND2_X1 U3661 ( .A1(n2264), .A2(n2867), .ZN(n2868) );
  NAND2_X1 U3662 ( .A1(n2868), .A2(n2982), .ZN(n3162) );
  INV_X1 U3663 ( .A(n3162), .ZN(n2869) );
  AOI22_X1 U3664 ( .A1(n3023), .A2(n2869), .B1(REG1_REG_1__SCAN_IN), .B2(n4724), .ZN(n2870) );
  OAI21_X1 U3665 ( .B1(n2960), .B2(n4724), .A(n2870), .ZN(U3519) );
  OAI21_X1 U3666 ( .B1(n2872), .B2(n3863), .A(n2871), .ZN(n3187) );
  AOI22_X1 U3667 ( .A1(n3936), .A2(n4475), .B1(n2286), .B2(n4473), .ZN(n2873)
         );
  OAI21_X1 U3668 ( .B1(n2265), .B2(n4478), .A(n2873), .ZN(n2880) );
  OAI21_X1 U3669 ( .B1(n2876), .B2(n2875), .A(n2874), .ZN(n2877) );
  NAND2_X1 U3670 ( .A1(n2877), .A2(n4370), .ZN(n2879) );
  NAND2_X1 U3671 ( .A1(n3187), .A2(n3400), .ZN(n2878) );
  NAND2_X1 U3672 ( .A1(n2879), .A2(n2878), .ZN(n3184) );
  AOI211_X1 U3673 ( .C1(n4711), .C2(n3187), .A(n2880), .B(n3184), .ZN(n2895)
         );
  XNOR2_X1 U3674 ( .A(n2982), .B(n2286), .ZN(n3183) );
  INV_X1 U3675 ( .A(n3183), .ZN(n2893) );
  AOI22_X1 U3676 ( .A1(n3023), .A2(n2893), .B1(REG1_REG_2__SCAN_IN), .B2(n4724), .ZN(n2881) );
  OAI21_X1 U3677 ( .B1(n2895), .B2(n4724), .A(n2881), .ZN(U3520) );
  XNOR2_X1 U3678 ( .A(n2961), .B(n4551), .ZN(n2963) );
  XNOR2_X1 U3679 ( .A(n2963), .B(REG2_REG_6__SCAN_IN), .ZN(n2892) );
  NOR2_X1 U3680 ( .A1(STATE_REG_SCAN_IN), .A2(n2883), .ZN(n3045) );
  AOI21_X1 U3681 ( .B1(n4650), .B2(ADDR_REG_6__SCAN_IN), .A(n3045), .ZN(n2884)
         );
  INV_X1 U3682 ( .A(n2884), .ZN(n2889) );
  INV_X1 U3683 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4722) );
  NOR2_X1 U3684 ( .A1(n2887), .A2(n4722), .ZN(n2966) );
  AOI211_X1 U3685 ( .C1(n4722), .C2(n2887), .A(n4627), .B(n2966), .ZN(n2888)
         );
  AOI211_X1 U3686 ( .C1(n2890), .C2(n4551), .A(n2889), .B(n2888), .ZN(n2891)
         );
  OAI21_X1 U3687 ( .B1(n2892), .B2(n4646), .A(n2891), .ZN(U3246) );
  INV_X1 U3688 ( .A(n4546), .ZN(n3025) );
  AOI22_X1 U3689 ( .A1(n3025), .A2(n2893), .B1(REG0_REG_2__SCAN_IN), .B2(n4718), .ZN(n2894) );
  OAI21_X1 U3690 ( .B1(n2895), .B2(n4718), .A(n2894), .ZN(U3471) );
  NAND2_X1 U3691 ( .A1(n2897), .A2(n2896), .ZN(n2898) );
  OAI21_X1 U3692 ( .B1(n2899), .B2(n2898), .A(STATE_REG_SCAN_IN), .ZN(n2901)
         );
  INV_X1 U3693 ( .A(n2902), .ZN(n2903) );
  OAI22_X1 U3694 ( .A1(n2906), .A2(n2905), .B1(n2904), .B2(n2903), .ZN(n2945)
         );
  INV_X1 U3695 ( .A(n2945), .ZN(n2915) );
  NAND2_X1 U3696 ( .A1(n2288), .A2(n2994), .ZN(n2908) );
  NAND2_X1 U3697 ( .A1(n2286), .A2(n3610), .ZN(n2907) );
  NAND2_X1 U3698 ( .A1(n2908), .A2(n2907), .ZN(n2909) );
  XNOR2_X1 U3699 ( .A(n2909), .B(n3613), .ZN(n2913) );
  INV_X1 U3700 ( .A(n2994), .ZN(n2910) );
  NOR2_X1 U3701 ( .A1(n2983), .A2(n2910), .ZN(n2911) );
  AOI21_X1 U3702 ( .B1(n2288), .B2(n3344), .A(n2911), .ZN(n2912) );
  NAND2_X1 U3703 ( .A1(n2913), .A2(n2912), .ZN(n2916) );
  OAI21_X1 U3704 ( .B1(n2913), .B2(n2912), .A(n2916), .ZN(n2948) );
  INV_X1 U3705 ( .A(n2948), .ZN(n2914) );
  NAND2_X1 U3706 ( .A1(n2915), .A2(n2914), .ZN(n2946) );
  NAND2_X1 U3707 ( .A1(n2946), .A2(n2916), .ZN(n2938) );
  NAND2_X1 U3708 ( .A1(n3936), .A2(n2994), .ZN(n2918) );
  NAND2_X1 U3709 ( .A1(n2986), .A2(n3610), .ZN(n2917) );
  AOI22_X1 U3710 ( .A1(n3936), .A2(n3344), .B1(n3609), .B2(n2986), .ZN(n2921)
         );
  XNOR2_X1 U3711 ( .A(n2920), .B(n2921), .ZN(n2939) );
  NAND2_X1 U3712 ( .A1(n2938), .A2(n2939), .ZN(n2930) );
  INV_X1 U3713 ( .A(n2920), .ZN(n2922) );
  NAND2_X1 U3714 ( .A1(n2922), .A2(n2921), .ZN(n2928) );
  AND2_X1 U3715 ( .A1(n2930), .A2(n2928), .ZN(n2932) );
  NAND2_X1 U3716 ( .A1(n3127), .A2(n2994), .ZN(n2925) );
  NAND2_X1 U3717 ( .A1(n2923), .A2(n3610), .ZN(n2924) );
  NAND2_X1 U3718 ( .A1(n2925), .A2(n2924), .ZN(n2926) );
  XNOR2_X1 U3719 ( .A(n2926), .B(n3597), .ZN(n2996) );
  NOR2_X1 U3720 ( .A1(n3068), .A2(n2910), .ZN(n2927) );
  AOI21_X1 U3721 ( .B1(n3127), .B2(n3544), .A(n2927), .ZN(n2999) );
  XNOR2_X1 U3722 ( .A(n2996), .B(n2999), .ZN(n2931) );
  NAND2_X1 U3723 ( .A1(n2930), .A2(n2929), .ZN(n2997) );
  OAI211_X1 U3724 ( .C1(n2932), .C2(n2931), .A(n3752), .B(n2997), .ZN(n2937)
         );
  INV_X1 U3725 ( .A(n3936), .ZN(n2933) );
  OAI22_X1 U3726 ( .A1(n2054), .A2(n3068), .B1(n2933), .B2(n3754), .ZN(n2934)
         );
  AOI211_X1 U3727 ( .C1(n3759), .C2(n3935), .A(n2935), .B(n2934), .ZN(n2936)
         );
  OAI211_X1 U3728 ( .C1(n3763), .C2(n3070), .A(n2937), .B(n2936), .ZN(U3227)
         );
  OAI21_X1 U3729 ( .B1(n2939), .B2(n2938), .A(n2930), .ZN(n2943) );
  MUX2_X1 U3730 ( .A(n3763), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n2941) );
  AOI22_X1 U3731 ( .A1(n3719), .A2(n2288), .B1(n3759), .B2(n3127), .ZN(n2940)
         );
  OAI211_X1 U3732 ( .C1(n2054), .C2(n3094), .A(n2941), .B(n2940), .ZN(n2942)
         );
  AOI21_X1 U3733 ( .B1(n2943), .B2(n3752), .A(n2942), .ZN(n2944) );
  INV_X1 U3734 ( .A(n2944), .ZN(U3215) );
  INV_X1 U3735 ( .A(n2946), .ZN(n2947) );
  AOI21_X1 U3736 ( .B1(n2945), .B2(n2948), .A(n2947), .ZN(n2952) );
  AOI22_X1 U3737 ( .A1(n3719), .A2(n2823), .B1(n3759), .B2(n3936), .ZN(n2949)
         );
  OAI21_X1 U3738 ( .B1(n2054), .B2(n2983), .A(n2949), .ZN(n2950) );
  AOI21_X1 U3739 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2955), .A(n2950), .ZN(n2951)
         );
  OAI21_X1 U3740 ( .B1(n2952), .B2(n3747), .A(n2951), .ZN(U3234) );
  OAI22_X1 U3741 ( .A1(n2054), .A2(n2953), .B1(n2265), .B2(n3742), .ZN(n2954)
         );
  AOI21_X1 U3742 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2955), .A(n2954), .ZN(n2956)
         );
  OAI21_X1 U3743 ( .B1(n3747), .B2(n2957), .A(n2956), .ZN(U3229) );
  CLKBUF_X1 U3744 ( .A(n4546), .Z(n4520) );
  OAI22_X1 U3745 ( .A1(n4520), .A2(n3162), .B1(n4719), .B2(n2252), .ZN(n2958)
         );
  INV_X1 U3746 ( .A(n2958), .ZN(n2959) );
  OAI21_X1 U3747 ( .B1(n2960), .B2(n4718), .A(n2959), .ZN(U3469) );
  INV_X1 U3748 ( .A(n2961), .ZN(n2962) );
  INV_X1 U3749 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3119) );
  MUX2_X1 U3750 ( .A(REG2_REG_7__SCAN_IN), .B(n3119), .S(n2971), .Z(n2964) );
  NOR2_X1 U3751 ( .A1(n2965), .A2(n2964), .ZN(n3008) );
  AOI211_X1 U3752 ( .C1(n2965), .C2(n2964), .A(n4646), .B(n3008), .ZN(n2974)
         );
  INV_X1 U3753 ( .A(n2971), .ZN(n3009) );
  NAND2_X1 U3754 ( .A1(n3009), .A2(REG1_REG_7__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U3755 ( .A1(n2089), .A2(n3006), .ZN(n2968) );
  OAI21_X1 U3756 ( .B1(n3007), .B2(n2968), .A(n4652), .ZN(n2967) );
  AOI21_X1 U3757 ( .B1(n3007), .B2(n2968), .A(n2967), .ZN(n2973) );
  NAND2_X1 U3758 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3172) );
  INV_X1 U3759 ( .A(n3172), .ZN(n2969) );
  AOI21_X1 U3760 ( .B1(n4650), .B2(ADDR_REG_7__SCAN_IN), .A(n2969), .ZN(n2970)
         );
  OAI21_X1 U3761 ( .B1(n4657), .B2(n2971), .A(n2970), .ZN(n2972) );
  OR3_X1 U3762 ( .A1(n2974), .A2(n2973), .A3(n2972), .ZN(U3247) );
  XNOR2_X1 U3763 ( .A(n2975), .B(n3868), .ZN(n3102) );
  INV_X1 U3764 ( .A(n3127), .ZN(n3095) );
  OAI22_X1 U3765 ( .A1(n3095), .A2(n4403), .B1(n4331), .B2(n3094), .ZN(n2981)
         );
  OAI21_X1 U3766 ( .B1(n2978), .B2(n2977), .A(n2976), .ZN(n2979) );
  AOI22_X1 U3767 ( .A1(n2979), .A2(n4370), .B1(n4400), .B2(n2288), .ZN(n3105)
         );
  INV_X1 U3768 ( .A(n3105), .ZN(n2980) );
  AOI211_X1 U3769 ( .C1(n4713), .C2(n3102), .A(n2981), .B(n2980), .ZN(n2989)
         );
  INV_X1 U3770 ( .A(n2982), .ZN(n2984) );
  NAND2_X1 U3771 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  AOI21_X1 U3772 ( .B1(n2986), .B2(n2985), .A(n3069), .ZN(n3098) );
  AOI22_X1 U3773 ( .A1(n3098), .A2(n3025), .B1(REG0_REG_3__SCAN_IN), .B2(n4718), .ZN(n2987) );
  OAI21_X1 U3774 ( .B1(n2989), .B2(n4718), .A(n2987), .ZN(U3473) );
  AOI22_X1 U3775 ( .A1(n3098), .A2(n3023), .B1(REG1_REG_3__SCAN_IN), .B2(n4724), .ZN(n2988) );
  OAI21_X1 U3776 ( .B1(n2989), .B2(n4724), .A(n2988), .ZN(U3521) );
  INV_X1 U3777 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U3778 ( .A1(n4200), .A2(U4043), .ZN(n2990) );
  OAI21_X1 U3779 ( .B1(U4043), .B2(n4091), .A(n2990), .ZN(U3577) );
  NAND2_X1 U3780 ( .A1(n3935), .A2(n3609), .ZN(n2992) );
  NAND2_X1 U3781 ( .A1(n3130), .A2(n3610), .ZN(n2991) );
  NAND2_X1 U3782 ( .A1(n2992), .A2(n2991), .ZN(n2993) );
  XNOR2_X1 U3783 ( .A(n2993), .B(n3597), .ZN(n3030) );
  NOR2_X1 U3784 ( .A1(n3001), .A2(n2910), .ZN(n2995) );
  AOI21_X1 U3785 ( .B1(n3935), .B2(n3544), .A(n2995), .ZN(n3032) );
  XNOR2_X1 U3786 ( .A(n3030), .B(n3032), .ZN(n3028) );
  INV_X1 U3787 ( .A(n2996), .ZN(n2998) );
  OAI21_X1 U3788 ( .B1(n2999), .B2(n2998), .A(n2997), .ZN(n3029) );
  XOR2_X1 U3789 ( .A(n3028), .B(n3029), .Z(n3000) );
  NAND2_X1 U3790 ( .A1(n3000), .A2(n3752), .ZN(n3005) );
  OAI22_X1 U3791 ( .A1(n2054), .A2(n3001), .B1(n3095), .B2(n3754), .ZN(n3002)
         );
  AOI211_X1 U3792 ( .C1(n3759), .C2(n3934), .A(n3003), .B(n3002), .ZN(n3004)
         );
  OAI211_X1 U3793 ( .C1(n3763), .C2(n3128), .A(n3005), .B(n3004), .ZN(U3224)
         );
  XOR2_X1 U3794 ( .A(REG1_REG_8__SCAN_IN), .B(n3476), .Z(n3015) );
  AOI21_X1 U3795 ( .B1(REG2_REG_7__SCAN_IN), .B2(n3009), .A(n3008), .ZN(n3492)
         );
  INV_X1 U3796 ( .A(n4550), .ZN(n3491) );
  XNOR2_X1 U3797 ( .A(n3492), .B(n3491), .ZN(n3493) );
  XNOR2_X1 U3798 ( .A(REG2_REG_8__SCAN_IN), .B(n3493), .ZN(n3010) );
  NAND2_X1 U3799 ( .A1(n4631), .A2(n3010), .ZN(n3011) );
  NAND2_X1 U3800 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3152) );
  NAND2_X1 U3801 ( .A1(n3011), .A2(n3152), .ZN(n3013) );
  NOR2_X1 U3802 ( .A1(n4657), .A2(n3491), .ZN(n3012) );
  AOI211_X1 U3803 ( .C1(n4650), .C2(ADDR_REG_8__SCAN_IN), .A(n3013), .B(n3012), 
        .ZN(n3014) );
  OAI21_X1 U3804 ( .B1(n3015), .B2(n4627), .A(n3014), .ZN(U3248) );
  INV_X1 U3805 ( .A(n3016), .ZN(n3774) );
  AND2_X1 U3806 ( .A1(n3774), .A2(n3788), .ZN(n3859) );
  XNOR2_X1 U3807 ( .A(n3017), .B(n3859), .ZN(n3135) );
  XOR2_X1 U3808 ( .A(n3859), .B(n3018), .Z(n3019) );
  NAND2_X1 U3809 ( .A1(n3019), .A2(n4370), .ZN(n3137) );
  AOI22_X1 U3810 ( .A1(n3934), .A2(n4475), .B1(n4473), .B2(n3130), .ZN(n3020)
         );
  OAI211_X1 U3811 ( .C1(n3095), .C2(n4478), .A(n3137), .B(n3020), .ZN(n3021)
         );
  AOI21_X1 U3812 ( .B1(n3135), .B2(n4713), .A(n3021), .ZN(n3027) );
  INV_X1 U3813 ( .A(n3022), .ZN(n3067) );
  AOI21_X1 U3814 ( .B1(n3130), .B2(n3067), .A(n3084), .ZN(n3126) );
  AOI22_X1 U3815 ( .A1(n3126), .A2(n3023), .B1(REG1_REG_5__SCAN_IN), .B2(n4724), .ZN(n3024) );
  OAI21_X1 U3816 ( .B1(n3027), .B2(n4724), .A(n3024), .ZN(U3523) );
  AOI22_X1 U3817 ( .A1(n3126), .A2(n3025), .B1(REG0_REG_5__SCAN_IN), .B2(n4718), .ZN(n3026) );
  OAI21_X1 U3818 ( .B1(n3027), .B2(n4718), .A(n3026), .ZN(U3477) );
  NAND2_X1 U3819 ( .A1(n3029), .A2(n3028), .ZN(n3034) );
  INV_X1 U3820 ( .A(n3030), .ZN(n3031) );
  OR2_X1 U3821 ( .A1(n3032), .A2(n3031), .ZN(n3033) );
  NAND2_X1 U3822 ( .A1(n3034), .A2(n3033), .ZN(n3140) );
  NAND2_X1 U3823 ( .A1(n3934), .A2(n3609), .ZN(n3036) );
  NAND2_X1 U3824 ( .A1(n3076), .A2(n3610), .ZN(n3035) );
  NAND2_X1 U3825 ( .A1(n3036), .A2(n3035), .ZN(n3037) );
  XNOR2_X1 U3826 ( .A(n3037), .B(n3613), .ZN(n3040) );
  NOR2_X1 U3827 ( .A1(n3083), .A2(n2910), .ZN(n3038) );
  AOI21_X1 U3828 ( .B1(n3934), .B2(n3544), .A(n3038), .ZN(n3039) );
  NOR2_X1 U3829 ( .A1(n3040), .A2(n3039), .ZN(n3139) );
  INV_X1 U3830 ( .A(n3139), .ZN(n3041) );
  NAND2_X1 U3831 ( .A1(n3040), .A2(n3039), .ZN(n3138) );
  NAND2_X1 U3832 ( .A1(n3041), .A2(n3138), .ZN(n3042) );
  XNOR2_X1 U3833 ( .A(n3140), .B(n3042), .ZN(n3043) );
  NAND2_X1 U3834 ( .A1(n3043), .A2(n3752), .ZN(n3047) );
  INV_X1 U3835 ( .A(n3935), .ZN(n3078) );
  OAI22_X1 U3836 ( .A1(n2054), .A2(n3083), .B1(n3078), .B2(n3754), .ZN(n3044)
         );
  AOI211_X1 U3837 ( .C1(n3759), .C2(n3933), .A(n3045), .B(n3044), .ZN(n3046)
         );
  OAI211_X1 U3838 ( .C1(n3763), .C2(n3087), .A(n3047), .B(n3046), .ZN(U3236)
         );
  INV_X1 U3839 ( .A(n3864), .ZN(n3050) );
  NAND2_X1 U3840 ( .A1(n3051), .A2(n3050), .ZN(n3052) );
  NAND2_X1 U3841 ( .A1(n3048), .A2(n3052), .ZN(n4701) );
  OAI21_X1 U3842 ( .B1(n4078), .B2(n3053), .A(n4682), .ZN(n3054) );
  NAND4_X1 U3843 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3058)
         );
  NAND2_X2 U3844 ( .A1(n3058), .A2(n4658), .ZN(n4365) );
  OR2_X1 U3845 ( .A1(n3059), .A2(n4146), .ZN(n3099) );
  INV_X1 U3846 ( .A(n3099), .ZN(n3060) );
  NAND2_X1 U3847 ( .A1(n4365), .A2(n3060), .ZN(n3168) );
  XNOR2_X1 U3848 ( .A(n3061), .B(n3864), .ZN(n3066) );
  NAND2_X1 U3849 ( .A1(n3936), .A2(n4400), .ZN(n3062) );
  OAI21_X1 U3850 ( .B1(n4331), .B2(n3068), .A(n3062), .ZN(n3064) );
  NOR2_X1 U3851 ( .A1(n4701), .A2(n3100), .ZN(n3063) );
  AOI211_X1 U3852 ( .C1(n4475), .C2(n3935), .A(n3064), .B(n3063), .ZN(n3065)
         );
  OAI21_X1 U3853 ( .B1(n4336), .B2(n3066), .A(n3065), .ZN(n4703) );
  OAI211_X1 U3854 ( .C1(n3069), .C2(n3068), .A(n3067), .B(n4351), .ZN(n4702)
         );
  OAI22_X1 U3855 ( .A1(n4702), .A2(n4362), .B1(n4658), .B2(n3070), .ZN(n3071)
         );
  OAI21_X1 U3856 ( .B1(n4703), .B2(n3071), .A(n4365), .ZN(n3073) );
  INV_X2 U3857 ( .A(n4365), .ZN(n4670) );
  NAND2_X1 U3858 ( .A1(n4670), .A2(REG2_REG_4__SCAN_IN), .ZN(n3072) );
  OAI211_X1 U3859 ( .C1(n4701), .C2(n3168), .A(n3073), .B(n3072), .ZN(U3286)
         );
  NAND2_X1 U3860 ( .A1(n3777), .A2(n3790), .ZN(n3867) );
  XNOR2_X1 U3861 ( .A(n3074), .B(n3867), .ZN(n3082) );
  XOR2_X1 U3862 ( .A(n3867), .B(n3075), .Z(n3080) );
  AOI22_X1 U3863 ( .A1(n3933), .A2(n4475), .B1(n4473), .B2(n3076), .ZN(n3077)
         );
  OAI21_X1 U3864 ( .B1(n3078), .B2(n4478), .A(n3077), .ZN(n3079) );
  AOI21_X1 U3865 ( .B1(n3080), .B2(n4370), .A(n3079), .ZN(n3081) );
  OAI21_X1 U3866 ( .B1(n3100), .B2(n3082), .A(n3081), .ZN(n4709) );
  INV_X1 U3867 ( .A(n4709), .ZN(n3092) );
  INV_X1 U3868 ( .A(n3082), .ZN(n4712) );
  INV_X1 U3869 ( .A(n3168), .ZN(n4665) );
  NOR2_X1 U3870 ( .A1(n3084), .A2(n3083), .ZN(n4708) );
  INV_X1 U3871 ( .A(n3112), .ZN(n4707) );
  INV_X1 U3872 ( .A(n3085), .ZN(n3086) );
  NAND2_X1 U3873 ( .A1(n4365), .A2(n3086), .ZN(n4341) );
  NOR3_X1 U3874 ( .A1(n4708), .A2(n4707), .A3(n4341), .ZN(n3090) );
  INV_X1 U3875 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3088) );
  OAI22_X1 U3876 ( .A1(n4365), .A2(n3088), .B1(n3087), .B2(n4658), .ZN(n3089)
         );
  AOI211_X1 U3877 ( .C1(n4712), .C2(n4665), .A(n3090), .B(n3089), .ZN(n3091)
         );
  OAI21_X1 U3878 ( .B1(n3092), .B2(n4670), .A(n3091), .ZN(U3284) );
  OAI22_X1 U3879 ( .A1(n4365), .A2(n3093), .B1(REG3_REG_3__SCAN_IN), .B2(n4658), .ZN(n3097) );
  AND2_X1 U3880 ( .A1(n4365), .A2(n4475), .ZN(n4377) );
  INV_X1 U3881 ( .A(n4377), .ZN(n4315) );
  NAND2_X1 U3882 ( .A1(n4365), .A2(n4473), .ZN(n4385) );
  OAI22_X1 U3883 ( .A1(n4315), .A2(n3095), .B1(n4385), .B2(n3094), .ZN(n3096)
         );
  AOI211_X1 U3884 ( .C1(n4664), .C2(n3098), .A(n3097), .B(n3096), .ZN(n3104)
         );
  NAND2_X1 U3885 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
  NAND2_X1 U3886 ( .A1(n3102), .A2(n4374), .ZN(n3103) );
  OAI211_X1 U3887 ( .C1(n3105), .C2(n4670), .A(n3104), .B(n3103), .ZN(U3287)
         );
  INV_X1 U3888 ( .A(n3860), .ZN(n3111) );
  NOR2_X1 U3889 ( .A1(n3106), .A2(n3916), .ZN(n3107) );
  OAI21_X1 U3890 ( .B1(n3108), .B2(n3107), .A(n4365), .ZN(n3110) );
  AOI22_X1 U3891 ( .A1(n4670), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4381), .ZN(n3109) );
  OAI211_X1 U3892 ( .C1(n3111), .C2(n3168), .A(n3110), .B(n3109), .ZN(U3290)
         );
  INV_X1 U3893 ( .A(n4351), .ZN(n4706) );
  AOI211_X1 U3894 ( .C1(n3171), .C2(n3112), .A(n4706), .B(n3228), .ZN(n4716)
         );
  XNOR2_X1 U3895 ( .A(n3114), .B(n3113), .ZN(n3118) );
  NOR2_X1 U3896 ( .A1(n3144), .A2(n4331), .ZN(n3115) );
  AOI21_X1 U3897 ( .B1(n3932), .B2(n4475), .A(n3115), .ZN(n3117) );
  NAND2_X1 U3898 ( .A1(n3934), .A2(n4400), .ZN(n3116) );
  OAI211_X1 U3899 ( .C1(n3118), .C2(n4336), .A(n3117), .B(n3116), .ZN(n4717)
         );
  AOI21_X1 U3900 ( .B1(n4716), .B2(n4146), .A(n4717), .ZN(n3125) );
  OAI22_X1 U3901 ( .A1(n4365), .A2(n3119), .B1(n3170), .B2(n4658), .ZN(n3120)
         );
  INV_X1 U3902 ( .A(n3120), .ZN(n3124) );
  NAND2_X1 U3903 ( .A1(n3122), .A2(n3873), .ZN(n4714) );
  NAND3_X1 U3904 ( .A1(n3121), .A2(n4714), .A3(n4374), .ZN(n3123) );
  OAI211_X1 U3905 ( .C1(n3125), .C2(n4670), .A(n3124), .B(n3123), .ZN(U3283)
         );
  INV_X1 U3906 ( .A(n3126), .ZN(n3133) );
  AND2_X1 U3907 ( .A1(n4365), .A2(n4400), .ZN(n4379) );
  AOI22_X1 U3908 ( .A1(n4379), .A2(n3127), .B1(n4377), .B2(n3934), .ZN(n3132)
         );
  INV_X1 U3909 ( .A(n4385), .ZN(n3334) );
  OAI22_X1 U3910 ( .A1(n4365), .A2(n2129), .B1(n3128), .B2(n4658), .ZN(n3129)
         );
  AOI21_X1 U3911 ( .B1(n3130), .B2(n3334), .A(n3129), .ZN(n3131) );
  OAI211_X1 U3912 ( .C1(n3133), .C2(n4341), .A(n3132), .B(n3131), .ZN(n3134)
         );
  AOI21_X1 U3913 ( .B1(n3135), .B2(n4374), .A(n3134), .ZN(n3136) );
  OAI21_X1 U3914 ( .B1(n3137), .B2(n4670), .A(n3136), .ZN(U3285) );
  OAI21_X2 U3915 ( .B1(n3140), .B2(n3139), .A(n3138), .ZN(n3175) );
  NAND2_X1 U3916 ( .A1(n3933), .A2(n3609), .ZN(n3142) );
  NAND2_X1 U3917 ( .A1(n3171), .A2(n3610), .ZN(n3141) );
  NAND2_X1 U3918 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  XNOR2_X1 U3919 ( .A(n3143), .B(n3597), .ZN(n3148) );
  NOR2_X1 U3920 ( .A1(n3144), .A2(n3615), .ZN(n3145) );
  AOI21_X1 U3921 ( .B1(n3933), .B2(n3544), .A(n3145), .ZN(n3146) );
  XOR2_X1 U3922 ( .A(n3148), .B(n3146), .Z(n3176) );
  NOR2_X1 U3923 ( .A1(n3175), .A2(n3176), .ZN(n3174) );
  INV_X1 U3924 ( .A(n3146), .ZN(n3147) );
  AND2_X1 U3925 ( .A1(n3148), .A2(n3147), .ZN(n3149) );
  AOI22_X1 U3926 ( .A1(n3932), .A2(n3609), .B1(n3610), .B2(n3231), .ZN(n3150)
         );
  XNOR2_X1 U3927 ( .A(n3150), .B(n3597), .ZN(n3215) );
  AOI22_X1 U3928 ( .A1(n3932), .A2(n3544), .B1(n3609), .B2(n3231), .ZN(n3216)
         );
  XNOR2_X1 U3929 ( .A(n3215), .B(n3216), .ZN(n3151) );
  XNOR2_X1 U3930 ( .A(n2085), .B(n3151), .ZN(n3157) );
  INV_X1 U3931 ( .A(n4659), .ZN(n3155) );
  INV_X1 U3932 ( .A(n3931), .ZN(n3252) );
  INV_X1 U3933 ( .A(n2054), .ZN(n3720) );
  AOI22_X1 U3934 ( .A1(n3720), .A2(n3231), .B1(n3719), .B2(n3933), .ZN(n3153)
         );
  OAI211_X1 U3935 ( .C1(n3252), .C2(n3742), .A(n3153), .B(n3152), .ZN(n3154)
         );
  AOI21_X1 U3936 ( .B1(n3155), .B2(n3745), .A(n3154), .ZN(n3156) );
  OAI21_X1 U3937 ( .B1(n3157), .B2(n3747), .A(n3156), .ZN(U3218) );
  MUX2_X1 U3938 ( .A(n3158), .B(REG2_REG_1__SCAN_IN), .S(n4670), .Z(n3159) );
  INV_X1 U3939 ( .A(n3159), .ZN(n3167) );
  OAI22_X1 U3940 ( .A1(n4385), .A2(n3161), .B1(n3160), .B2(n4658), .ZN(n3165)
         );
  INV_X1 U3941 ( .A(n4379), .ZN(n4317) );
  OAI22_X1 U3942 ( .A1(n4317), .A2(n3163), .B1(n3162), .B2(n4341), .ZN(n3164)
         );
  AOI211_X1 U3943 ( .C1(n4377), .C2(n2288), .A(n3165), .B(n3164), .ZN(n3166)
         );
  OAI211_X1 U3944 ( .C1(n3169), .C2(n3168), .A(n3167), .B(n3166), .ZN(U3289)
         );
  INV_X1 U3945 ( .A(n3170), .ZN(n3179) );
  INV_X1 U3946 ( .A(n3932), .ZN(n3220) );
  AOI22_X1 U3947 ( .A1(n3720), .A2(n3171), .B1(n3719), .B2(n3934), .ZN(n3173)
         );
  OAI211_X1 U3948 ( .C1(n3220), .C2(n3742), .A(n3173), .B(n3172), .ZN(n3178)
         );
  AOI211_X1 U3949 ( .C1(n3176), .C2(n3175), .A(n3747), .B(n3174), .ZN(n3177)
         );
  AOI211_X1 U3950 ( .C1(n3179), .C2(n3745), .A(n3178), .B(n3177), .ZN(n3180)
         );
  INV_X1 U3951 ( .A(n3180), .ZN(U3210) );
  AOI22_X1 U3952 ( .A1(n4377), .A2(n3936), .B1(n4379), .B2(n2823), .ZN(n3182)
         );
  AOI22_X1 U3953 ( .A1(n3334), .A2(n2286), .B1(REG3_REG_2__SCAN_IN), .B2(n4381), .ZN(n3181) );
  OAI211_X1 U3954 ( .C1(n3183), .C2(n4341), .A(n3182), .B(n3181), .ZN(n3186)
         );
  MUX2_X1 U3955 ( .A(n3184), .B(REG2_REG_2__SCAN_IN), .S(n4670), .Z(n3185) );
  AOI211_X1 U3956 ( .C1(n4665), .C2(n3187), .A(n3186), .B(n3185), .ZN(n3188)
         );
  INV_X1 U3957 ( .A(n3188), .ZN(U3288) );
  INV_X1 U3958 ( .A(n3785), .ZN(n3792) );
  AND2_X1 U3959 ( .A1(n3792), .A2(n3781), .ZN(n3843) );
  XNOR2_X1 U3960 ( .A(n3189), .B(n3843), .ZN(n3200) );
  NAND2_X1 U3961 ( .A1(n3226), .A2(n3214), .ZN(n3190) );
  NAND2_X1 U3962 ( .A1(n3258), .A2(n3190), .ZN(n3212) );
  INV_X1 U3963 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3951) );
  OAI22_X1 U3964 ( .A1(n3225), .A2(n4658), .B1(n3951), .B2(n4365), .ZN(n3191)
         );
  AOI21_X1 U3965 ( .B1(n3334), .B2(n3214), .A(n3191), .ZN(n3193) );
  AOI22_X1 U3966 ( .A1(n4379), .A2(n3932), .B1(n4377), .B2(n3930), .ZN(n3192)
         );
  OAI211_X1 U3967 ( .C1(n3212), .C2(n4341), .A(n3193), .B(n3192), .ZN(n3198)
         );
  INV_X1 U3968 ( .A(n3843), .ZN(n3194) );
  XNOR2_X1 U3969 ( .A(n3195), .B(n3194), .ZN(n3196) );
  NAND2_X1 U3970 ( .A1(n3196), .A2(n4370), .ZN(n3205) );
  NOR2_X1 U3971 ( .A1(n3205), .A2(n4670), .ZN(n3197) );
  AOI211_X1 U3972 ( .C1(n3200), .C2(n4374), .A(n3198), .B(n3197), .ZN(n3199)
         );
  INV_X1 U3973 ( .A(n3199), .ZN(U3281) );
  INV_X1 U3974 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U3975 ( .A1(n3200), .A2(n4713), .ZN(n3206) );
  NAND2_X1 U3976 ( .A1(n3932), .A2(n4400), .ZN(n3202) );
  NAND2_X1 U3977 ( .A1(n3930), .A2(n4475), .ZN(n3201) );
  OAI211_X1 U3978 ( .C1(n4331), .C2(n3221), .A(n3202), .B(n3201), .ZN(n3203)
         );
  INV_X1 U3979 ( .A(n3203), .ZN(n3204) );
  AND3_X1 U3980 ( .A1(n3206), .A2(n3205), .A3(n3204), .ZN(n3209) );
  MUX2_X1 U3981 ( .A(n3207), .B(n3209), .S(n4727), .Z(n3208) );
  OAI21_X1 U3982 ( .B1(n4486), .B2(n3212), .A(n3208), .ZN(U3527) );
  MUX2_X1 U3983 ( .A(n3210), .B(n3209), .S(n4719), .Z(n3211) );
  OAI21_X1 U3984 ( .B1(n3212), .B2(n4546), .A(n3211), .ZN(U3485) );
  AOI22_X1 U3985 ( .A1(n3931), .A2(n3609), .B1(n3610), .B2(n3214), .ZN(n3213)
         );
  XNOR2_X1 U3986 ( .A(n3213), .B(n3597), .ZN(n3241) );
  AOI22_X1 U3987 ( .A1(n3931), .A2(n3544), .B1(n3609), .B2(n3214), .ZN(n3240)
         );
  XOR2_X1 U3988 ( .A(n3241), .B(n3240), .Z(n3218) );
  NAND2_X1 U3989 ( .A1(n3217), .A2(n3218), .ZN(n3248) );
  OAI21_X1 U3990 ( .B1(n3218), .B2(n3217), .A(n3248), .ZN(n3219) );
  NAND2_X1 U3991 ( .A1(n3219), .A2(n3752), .ZN(n3224) );
  AND2_X1 U3992 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4569) );
  OAI22_X1 U3993 ( .A1(n2054), .A2(n3221), .B1(n3220), .B2(n3754), .ZN(n3222)
         );
  AOI211_X1 U3994 ( .C1(n3759), .C2(n3930), .A(n4569), .B(n3222), .ZN(n3223)
         );
  OAI211_X1 U3995 ( .C1(n3763), .C2(n3225), .A(n3224), .B(n3223), .ZN(U3228)
         );
  OAI21_X1 U3996 ( .B1(n3228), .B2(n3227), .A(n3226), .ZN(n4662) );
  AND2_X1 U3997 ( .A1(n3780), .A2(n3791), .ZN(n3842) );
  XNOR2_X1 U3998 ( .A(n3229), .B(n3842), .ZN(n4666) );
  XNOR2_X1 U3999 ( .A(n3230), .B(n3842), .ZN(n3234) );
  AOI22_X1 U4000 ( .A1(n3933), .A2(n4400), .B1(n4473), .B2(n3231), .ZN(n3233)
         );
  NAND2_X1 U4001 ( .A1(n3931), .A2(n4475), .ZN(n3232) );
  OAI211_X1 U4002 ( .C1(n3234), .C2(n4336), .A(n3233), .B(n3232), .ZN(n3235)
         );
  AOI21_X1 U4003 ( .B1(n3400), .B2(n4666), .A(n3235), .ZN(n4669) );
  INV_X1 U4004 ( .A(n4669), .ZN(n3236) );
  AOI21_X1 U4005 ( .B1(n4711), .B2(n4666), .A(n3236), .ZN(n3238) );
  MUX2_X1 U4006 ( .A(n3475), .B(n3238), .S(n4727), .Z(n3237) );
  OAI21_X1 U4007 ( .B1(n4662), .B2(n4486), .A(n3237), .ZN(U3526) );
  MUX2_X1 U4008 ( .A(n2352), .B(n3238), .S(n4719), .Z(n3239) );
  OAI21_X1 U4009 ( .B1(n4662), .B2(n4520), .A(n3239), .ZN(U3483) );
  NAND2_X1 U4010 ( .A1(n3241), .A2(n3240), .ZN(n3246) );
  AND2_X1 U4011 ( .A1(n3248), .A2(n3246), .ZN(n3250) );
  NAND2_X1 U4012 ( .A1(n3930), .A2(n3609), .ZN(n3243) );
  NAND2_X1 U4013 ( .A1(n3263), .A2(n3610), .ZN(n3242) );
  NAND2_X1 U4014 ( .A1(n3243), .A2(n3242), .ZN(n3244) );
  XNOR2_X1 U4015 ( .A(n3244), .B(n3597), .ZN(n3302) );
  NOR2_X1 U4016 ( .A1(n3291), .A2(n2910), .ZN(n3245) );
  AOI21_X1 U4017 ( .B1(n3930), .B2(n3544), .A(n3245), .ZN(n3303) );
  XNOR2_X1 U4018 ( .A(n3302), .B(n3303), .ZN(n3249) );
  OAI211_X1 U4019 ( .C1(n3250), .C2(n3249), .A(n3752), .B(n3306), .ZN(n3255)
         );
  INV_X1 U4020 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3251) );
  NOR2_X1 U4021 ( .A1(STATE_REG_SCAN_IN), .A2(n3251), .ZN(n4579) );
  OAI22_X1 U4022 ( .A1(n2054), .A2(n3291), .B1(n3252), .B2(n3754), .ZN(n3253)
         );
  AOI211_X1 U4023 ( .C1(n3759), .C2(n3929), .A(n4579), .B(n3253), .ZN(n3254)
         );
  OAI211_X1 U4024 ( .C1(n3763), .C2(n3260), .A(n3255), .B(n3254), .ZN(U3214)
         );
  AND2_X1 U4025 ( .A1(n3797), .A2(n3798), .ZN(n3844) );
  INV_X1 U4026 ( .A(n3844), .ZN(n3256) );
  XNOR2_X1 U4027 ( .A(n3257), .B(n3256), .ZN(n3288) );
  NAND2_X1 U4028 ( .A1(n3258), .A2(n3263), .ZN(n3259) );
  INV_X1 U4029 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3261) );
  OAI22_X1 U4030 ( .A1(n4365), .A2(n3261), .B1(n3260), .B2(n4658), .ZN(n3262)
         );
  AOI21_X1 U4031 ( .B1(n4377), .B2(n3929), .A(n3262), .ZN(n3265) );
  AOI22_X1 U4032 ( .A1(n3334), .A2(n3263), .B1(n4379), .B2(n3931), .ZN(n3264)
         );
  OAI211_X1 U4033 ( .C1(n3301), .C2(n4341), .A(n3265), .B(n3264), .ZN(n3269)
         );
  XNOR2_X1 U4034 ( .A(n3266), .B(n3844), .ZN(n3267) );
  NAND2_X1 U4035 ( .A1(n3267), .A2(n4370), .ZN(n3294) );
  NOR2_X1 U4036 ( .A1(n3294), .A2(n4670), .ZN(n3268) );
  AOI211_X1 U4037 ( .C1(n4374), .C2(n3288), .A(n3269), .B(n3268), .ZN(n3270)
         );
  INV_X1 U4038 ( .A(n3270), .ZN(U3280) );
  XNOR2_X1 U4039 ( .A(n3325), .B(n3865), .ZN(n3279) );
  NAND2_X1 U4040 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  NAND2_X1 U4041 ( .A1(n3274), .A2(n3273), .ZN(n3354) );
  NAND2_X1 U4042 ( .A1(n3928), .A2(n4475), .ZN(n3276) );
  NAND2_X1 U40430 ( .A1(n3930), .A2(n4400), .ZN(n3275) );
  OAI211_X1 U4044 ( .C1(n4331), .C2(n3319), .A(n3276), .B(n3275), .ZN(n3277)
         );
  AOI21_X1 U4045 ( .B1(n3354), .B2(n3400), .A(n3277), .ZN(n3278) );
  OAI21_X1 U4046 ( .B1(n4336), .B2(n3279), .A(n3278), .ZN(n3353) );
  INV_X1 U4047 ( .A(n3353), .ZN(n3287) );
  INV_X1 U4048 ( .A(n3330), .ZN(n3282) );
  NAND2_X1 U4049 ( .A1(n3280), .A2(n3307), .ZN(n3281) );
  NAND2_X1 U4050 ( .A1(n3282), .A2(n3281), .ZN(n3360) );
  NOR2_X1 U4051 ( .A1(n3360), .A2(n4341), .ZN(n3285) );
  INV_X1 U4052 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3283) );
  OAI22_X1 U4053 ( .A1(n4365), .A2(n3283), .B1(n3323), .B2(n4658), .ZN(n3284)
         );
  AOI211_X1 U4054 ( .C1(n3354), .C2(n4665), .A(n3285), .B(n3284), .ZN(n3286)
         );
  OAI21_X1 U4055 ( .B1(n3287), .B2(n4670), .A(n3286), .ZN(U3279) );
  NAND2_X1 U4056 ( .A1(n3288), .A2(n4713), .ZN(n3295) );
  NAND2_X1 U4057 ( .A1(n3931), .A2(n4400), .ZN(n3290) );
  NAND2_X1 U4058 ( .A1(n3929), .A2(n4475), .ZN(n3289) );
  OAI211_X1 U4059 ( .C1(n4331), .C2(n3291), .A(n3290), .B(n3289), .ZN(n3292)
         );
  INV_X1 U4060 ( .A(n3292), .ZN(n3293) );
  NAND3_X1 U4061 ( .A1(n3295), .A2(n3294), .A3(n3293), .ZN(n3298) );
  MUX2_X1 U4062 ( .A(REG0_REG_10__SCAN_IN), .B(n3298), .S(n4719), .Z(n3296) );
  INV_X1 U4063 ( .A(n3296), .ZN(n3297) );
  OAI21_X1 U4064 ( .B1(n3301), .B2(n4546), .A(n3297), .ZN(U3487) );
  MUX2_X1 U4065 ( .A(REG1_REG_10__SCAN_IN), .B(n3298), .S(n4727), .Z(n3299) );
  INV_X1 U4066 ( .A(n3299), .ZN(n3300) );
  OAI21_X1 U4067 ( .B1(n4486), .B2(n3301), .A(n3300), .ZN(U3528) );
  NAND2_X1 U4068 ( .A1(n3929), .A2(n3609), .ZN(n3309) );
  NAND2_X1 U4069 ( .A1(n3307), .A2(n3610), .ZN(n3308) );
  NAND2_X1 U4070 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  XNOR2_X1 U4071 ( .A(n3310), .B(n3613), .ZN(n3313) );
  NOR2_X1 U4072 ( .A1(n3319), .A2(n3615), .ZN(n3311) );
  AOI21_X1 U4073 ( .B1(n3929), .B2(n3544), .A(n3311), .ZN(n3312) );
  NOR2_X1 U4074 ( .A1(n3313), .A2(n3312), .ZN(n3340) );
  INV_X1 U4075 ( .A(n3340), .ZN(n3314) );
  NAND2_X1 U4076 ( .A1(n3313), .A2(n3312), .ZN(n3341) );
  NAND2_X1 U4077 ( .A1(n3314), .A2(n3341), .ZN(n3315) );
  XNOR2_X1 U4078 ( .A(n3342), .B(n3315), .ZN(n3316) );
  NAND2_X1 U4079 ( .A1(n3316), .A2(n3752), .ZN(n3322) );
  INV_X1 U4080 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3317) );
  NOR2_X1 U4081 ( .A1(STATE_REG_SCAN_IN), .A2(n3317), .ZN(n4590) );
  OAI22_X1 U4082 ( .A1(n2054), .A2(n3319), .B1(n3318), .B2(n3754), .ZN(n3320)
         );
  AOI211_X1 U4083 ( .C1(n3759), .C2(n3928), .A(n4590), .B(n3320), .ZN(n3321)
         );
  OAI211_X1 U4084 ( .C1(n3763), .C2(n3323), .A(n3322), .B(n3321), .ZN(U3233)
         );
  AND2_X1 U4085 ( .A1(n3361), .A2(n3362), .ZN(n3845) );
  XOR2_X1 U4086 ( .A(n3845), .B(n3324), .Z(n3382) );
  INV_X1 U4087 ( .A(n3382), .ZN(n3339) );
  INV_X1 U4088 ( .A(n3325), .ZN(n3328) );
  AOI21_X1 U4089 ( .B1(n3328), .B2(n3327), .A(n3326), .ZN(n3364) );
  XOR2_X1 U4090 ( .A(n3845), .B(n3364), .Z(n3329) );
  NOR2_X1 U4091 ( .A1(n3329), .A2(n4336), .ZN(n3380) );
  NOR2_X1 U4092 ( .A1(n3330), .A2(n3379), .ZN(n3331) );
  OR2_X1 U4093 ( .A1(n3370), .A2(n3331), .ZN(n3388) );
  INV_X1 U4094 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3332) );
  OAI22_X1 U4095 ( .A1(n4365), .A2(n3332), .B1(n3346), .B2(n4658), .ZN(n3333)
         );
  AOI21_X1 U4096 ( .B1(n3347), .B2(n3334), .A(n3333), .ZN(n3336) );
  AOI22_X1 U4097 ( .A1(n4379), .A2(n3929), .B1(n4377), .B2(n3927), .ZN(n3335)
         );
  OAI211_X1 U4098 ( .C1(n3388), .C2(n4341), .A(n3336), .B(n3335), .ZN(n3337)
         );
  AOI21_X1 U4099 ( .B1(n3380), .B2(n4365), .A(n3337), .ZN(n3338) );
  OAI21_X1 U4100 ( .B1(n3339), .B2(n4368), .A(n3338), .ZN(U3278) );
  AOI22_X1 U4101 ( .A1(n3928), .A2(n3609), .B1(n3610), .B2(n3347), .ZN(n3343)
         );
  XNOR2_X1 U4102 ( .A(n3343), .B(n3597), .ZN(n3420) );
  INV_X1 U4103 ( .A(n3420), .ZN(n3422) );
  INV_X1 U4104 ( .A(n3928), .ZN(n3427) );
  INV_X1 U4105 ( .A(n3344), .ZN(n3599) );
  OAI22_X1 U4106 ( .A1(n3427), .A2(n3599), .B1(n2910), .B2(n3379), .ZN(n3423)
         );
  XNOR2_X1 U4107 ( .A(n3422), .B(n3423), .ZN(n3345) );
  XNOR2_X1 U4108 ( .A(n3421), .B(n3345), .ZN(n3352) );
  INV_X1 U4109 ( .A(n3346), .ZN(n3350) );
  INV_X1 U4110 ( .A(n3927), .ZN(n4479) );
  AOI22_X1 U4111 ( .A1(n3720), .A2(n3347), .B1(n3719), .B2(n3929), .ZN(n3348)
         );
  NAND2_X1 U4112 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4595) );
  OAI211_X1 U4113 ( .C1(n4479), .C2(n3742), .A(n3348), .B(n4595), .ZN(n3349)
         );
  AOI21_X1 U4114 ( .B1(n3350), .B2(n3745), .A(n3349), .ZN(n3351) );
  OAI21_X1 U4115 ( .B1(n3352), .B2(n3747), .A(n3351), .ZN(U3221) );
  INV_X1 U4116 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3355) );
  AOI21_X1 U4117 ( .B1(n4711), .B2(n3354), .A(n3353), .ZN(n3357) );
  MUX2_X1 U4118 ( .A(n3355), .B(n3357), .S(n4727), .Z(n3356) );
  OAI21_X1 U4119 ( .B1(n4486), .B2(n3360), .A(n3356), .ZN(U3529) );
  MUX2_X1 U4120 ( .A(n3358), .B(n3357), .S(n4719), .Z(n3359) );
  OAI21_X1 U4121 ( .B1(n3360), .B2(n4546), .A(n3359), .ZN(U3489) );
  INV_X1 U4122 ( .A(n3361), .ZN(n3363) );
  OAI21_X1 U4123 ( .B1(n3364), .B2(n3363), .A(n3362), .ZN(n3365) );
  XNOR2_X1 U4124 ( .A(n3927), .B(n3413), .ZN(n3875) );
  XNOR2_X1 U4125 ( .A(n3365), .B(n3875), .ZN(n3368) );
  INV_X1 U4126 ( .A(n3452), .ZN(n3755) );
  OAI22_X1 U4127 ( .A1(n3755), .A2(n4403), .B1(n4331), .B2(n3428), .ZN(n3366)
         );
  AOI21_X1 U4128 ( .B1(n4400), .B2(n3928), .A(n3366), .ZN(n3367) );
  OAI21_X1 U4129 ( .B1(n3368), .B2(n4336), .A(n3367), .ZN(n3389) );
  INV_X1 U4130 ( .A(n3389), .ZN(n3376) );
  XOR2_X1 U4131 ( .A(n3875), .B(n3369), .Z(n3390) );
  OR2_X1 U4132 ( .A1(n3370), .A2(n3428), .ZN(n3371) );
  NAND2_X1 U4133 ( .A1(n3401), .A2(n3371), .ZN(n3395) );
  NOR2_X1 U4134 ( .A1(n3395), .A2(n4341), .ZN(n3374) );
  INV_X1 U4135 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3372) );
  OAI22_X1 U4136 ( .A1(n4365), .A2(n3372), .B1(n3432), .B2(n4658), .ZN(n3373)
         );
  AOI211_X1 U4137 ( .C1(n3390), .C2(n4374), .A(n3374), .B(n3373), .ZN(n3375)
         );
  OAI21_X1 U4138 ( .B1(n3376), .B2(n4670), .A(n3375), .ZN(U3277) );
  NAND2_X1 U4139 ( .A1(n3929), .A2(n4400), .ZN(n3378) );
  NAND2_X1 U4140 ( .A1(n3927), .A2(n4475), .ZN(n3377) );
  OAI211_X1 U4141 ( .C1(n4331), .C2(n3379), .A(n3378), .B(n3377), .ZN(n3381)
         );
  AOI211_X1 U4142 ( .C1(n4713), .C2(n3382), .A(n3381), .B(n3380), .ZN(n3385)
         );
  MUX2_X1 U4143 ( .A(n3383), .B(n3385), .S(n4719), .Z(n3384) );
  OAI21_X1 U4144 ( .B1(n3388), .B2(n4546), .A(n3384), .ZN(U3491) );
  INV_X1 U4145 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3386) );
  MUX2_X1 U4146 ( .A(n3386), .B(n3385), .S(n4727), .Z(n3387) );
  OAI21_X1 U4147 ( .B1(n4486), .B2(n3388), .A(n3387), .ZN(U3530) );
  AOI21_X1 U4148 ( .B1(n4713), .B2(n3390), .A(n3389), .ZN(n3393) );
  MUX2_X1 U4149 ( .A(n3391), .B(n3393), .S(n4719), .Z(n3392) );
  OAI21_X1 U4150 ( .B1(n3395), .B2(n4520), .A(n3392), .ZN(U3493) );
  INV_X1 U4151 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3483) );
  MUX2_X1 U4152 ( .A(n3483), .B(n3393), .S(n4727), .Z(n3394) );
  OAI21_X1 U4153 ( .B1(n4486), .B2(n3395), .A(n3394), .ZN(U3531) );
  OAI21_X1 U4154 ( .B1(n3398), .B2(n3397), .A(n3396), .ZN(n4483) );
  OAI21_X1 U4155 ( .B1(n3872), .B2(n3881), .A(n3444), .ZN(n3399) );
  AOI22_X1 U4156 ( .A1(n4483), .A2(n3400), .B1(n4370), .B2(n3399), .ZN(n4480)
         );
  INV_X1 U4157 ( .A(n3401), .ZN(n3402) );
  OAI21_X1 U4158 ( .B1(n3402), .B2(n3406), .A(n3449), .ZN(n4547) );
  NOR2_X1 U4159 ( .A1(n4547), .A2(n4341), .ZN(n3408) );
  AOI22_X1 U4160 ( .A1(n4377), .A2(n4476), .B1(n4379), .B2(n3927), .ZN(n3405)
         );
  INV_X1 U4161 ( .A(n3403), .ZN(n3441) );
  AOI22_X1 U4162 ( .A1(n4670), .A2(REG2_REG_14__SCAN_IN), .B1(n3441), .B2(
        n4381), .ZN(n3404) );
  OAI211_X1 U4163 ( .C1(n3406), .C2(n4385), .A(n3405), .B(n3404), .ZN(n3407)
         );
  AOI211_X1 U4164 ( .C1(n4483), .C2(n4665), .A(n3408), .B(n3407), .ZN(n3409)
         );
  OAI21_X1 U4165 ( .B1(n4480), .B2(n4670), .A(n3409), .ZN(U3276) );
  NAND2_X1 U4166 ( .A1(n3927), .A2(n3609), .ZN(n3411) );
  NAND2_X1 U4167 ( .A1(n3413), .A2(n3610), .ZN(n3410) );
  NAND2_X1 U4168 ( .A1(n3411), .A2(n3410), .ZN(n3412) );
  XNOR2_X1 U4169 ( .A(n3412), .B(n3597), .ZN(n3416) );
  NAND2_X1 U4170 ( .A1(n3927), .A2(n3544), .ZN(n3415) );
  NAND2_X1 U4171 ( .A1(n3413), .A2(n3609), .ZN(n3414) );
  NAND2_X1 U4172 ( .A1(n3415), .A2(n3414), .ZN(n3417) );
  NAND2_X1 U4173 ( .A1(n3416), .A2(n3417), .ZN(n3433) );
  INV_X1 U4174 ( .A(n3416), .ZN(n3419) );
  INV_X1 U4175 ( .A(n3417), .ZN(n3418) );
  NAND2_X1 U4176 ( .A1(n3419), .A2(n3418), .ZN(n3435) );
  NAND2_X1 U4177 ( .A1(n3433), .A2(n3435), .ZN(n3424) );
  XOR2_X1 U4178 ( .A(n3424), .B(n3434), .Z(n3425) );
  NAND2_X1 U4179 ( .A1(n3425), .A2(n3752), .ZN(n3431) );
  NOR2_X1 U4180 ( .A1(STATE_REG_SCAN_IN), .A2(n3426), .ZN(n3486) );
  OAI22_X1 U4181 ( .A1(n2054), .A2(n3428), .B1(n3427), .B2(n3754), .ZN(n3429)
         );
  AOI211_X1 U4182 ( .C1(n3759), .C2(n3452), .A(n3486), .B(n3429), .ZN(n3430)
         );
  OAI211_X1 U4183 ( .C1(n3763), .C2(n3432), .A(n3431), .B(n3430), .ZN(U3231)
         );
  AOI22_X1 U4184 ( .A1(n3452), .A2(n3609), .B1(n3610), .B2(n4474), .ZN(n3436)
         );
  XNOR2_X1 U4185 ( .A(n3436), .B(n3597), .ZN(n3519) );
  AOI22_X1 U4186 ( .A1(n3452), .A2(n3544), .B1(n3609), .B2(n4474), .ZN(n3518)
         );
  XNOR2_X1 U4187 ( .A(n3519), .B(n3518), .ZN(n3437) );
  XNOR2_X1 U4188 ( .A(n3520), .B(n3437), .ZN(n3443) );
  INV_X1 U4189 ( .A(n4476), .ZN(n3439) );
  AOI22_X1 U4190 ( .A1(n3720), .A2(n4474), .B1(n3719), .B2(n3927), .ZN(n3438)
         );
  NAND2_X1 U4191 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4602) );
  OAI211_X1 U4192 ( .C1(n3439), .C2(n3742), .A(n3438), .B(n4602), .ZN(n3440)
         );
  AOI21_X1 U4193 ( .B1(n3441), .B2(n3745), .A(n3440), .ZN(n3442) );
  OAI21_X1 U4194 ( .B1(n3443), .B2(n3747), .A(n3442), .ZN(U3212) );
  NAND2_X1 U4195 ( .A1(n3444), .A2(n3804), .ZN(n3446) );
  INV_X1 U4196 ( .A(n3861), .ZN(n3445) );
  XNOR2_X1 U4197 ( .A(n3446), .B(n3445), .ZN(n3447) );
  NAND2_X1 U4198 ( .A1(n3447), .A2(n4370), .ZN(n3505) );
  XNOR2_X1 U4199 ( .A(n3448), .B(n3861), .ZN(n3507) );
  NAND2_X1 U4200 ( .A1(n3507), .A2(n4374), .ZN(n3459) );
  INV_X1 U4201 ( .A(n3449), .ZN(n3451) );
  INV_X1 U4202 ( .A(n3470), .ZN(n3450) );
  OAI21_X1 U4203 ( .B1(n3451), .B2(n3756), .A(n3450), .ZN(n3513) );
  INV_X1 U4204 ( .A(n3513), .ZN(n3457) );
  AOI22_X1 U4205 ( .A1(n4379), .A2(n3452), .B1(n4377), .B2(n4378), .ZN(n3455)
         );
  INV_X1 U4206 ( .A(n3762), .ZN(n3453) );
  AOI22_X1 U4207 ( .A1(n4670), .A2(REG2_REG_15__SCAN_IN), .B1(n3453), .B2(
        n4381), .ZN(n3454) );
  OAI211_X1 U4208 ( .C1(n3756), .C2(n4385), .A(n3455), .B(n3454), .ZN(n3456)
         );
  AOI21_X1 U4209 ( .B1(n3457), .B2(n4664), .A(n3456), .ZN(n3458) );
  OAI211_X1 U4210 ( .C1(n4670), .C2(n3505), .A(n3459), .B(n3458), .ZN(U3275)
         );
  OAI21_X1 U4211 ( .B1(n3462), .B2(n3461), .A(n3460), .ZN(n4468) );
  XNOR2_X1 U4212 ( .A(n3463), .B(n3874), .ZN(n3467) );
  NOR2_X1 U4213 ( .A1(n3469), .A2(n4331), .ZN(n3464) );
  AOI21_X1 U4214 ( .B1(n3682), .B2(n4475), .A(n3464), .ZN(n3466) );
  NAND2_X1 U4215 ( .A1(n4476), .A2(n4400), .ZN(n3465) );
  OAI211_X1 U4216 ( .C1(n3467), .C2(n4336), .A(n3466), .B(n3465), .ZN(n4469)
         );
  INV_X1 U4217 ( .A(n4376), .ZN(n3468) );
  OAI21_X1 U4218 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n4542) );
  NOR2_X1 U4219 ( .A1(n4542), .A2(n4341), .ZN(n3472) );
  OAI22_X1 U4220 ( .A1(n4365), .A2(n4623), .B1(n3681), .B2(n4658), .ZN(n3471)
         );
  AOI211_X1 U4221 ( .C1(n4469), .C2(n4365), .A(n3472), .B(n3471), .ZN(n3473)
         );
  OAI21_X1 U4222 ( .B1(n4468), .B2(n4368), .A(n3473), .ZN(U3274) );
  NAND2_X1 U4223 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3490), .ZN(n3480) );
  AOI22_X1 U4224 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3490), .B1(n4696), .B2(
        n3355), .ZN(n4583) );
  NAND2_X1 U4225 ( .A1(n4558), .A2(REG1_REG_9__SCAN_IN), .ZN(n3477) );
  MUX2_X1 U4226 ( .A(n3207), .B(REG1_REG_9__SCAN_IN), .S(n4558), .Z(n3474) );
  INV_X1 U4227 ( .A(n3474), .ZN(n4560) );
  INV_X1 U4228 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U4229 ( .A1(n4560), .A2(n4561), .ZN(n4559) );
  NAND2_X1 U4230 ( .A1(n3477), .A2(n4559), .ZN(n3478) );
  NAND2_X1 U4231 ( .A1(n4571), .A2(n3478), .ZN(n3479) );
  XOR2_X1 U4232 ( .A(n3478), .B(n4571), .Z(n4573) );
  NAND2_X1 U4233 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U4234 ( .A1(n4592), .A2(n3481), .ZN(n3482) );
  NAND2_X1 U4235 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4599), .ZN(n4598) );
  NOR2_X1 U4236 ( .A1(n3489), .A2(n3483), .ZN(n4127) );
  AOI21_X1 U4237 ( .B1(n3483), .B2(n3489), .A(n4127), .ZN(n3484) );
  OAI211_X1 U4238 ( .C1(n3485), .C2(n3484), .A(n4652), .B(n4128), .ZN(n3488)
         );
  AOI21_X1 U4239 ( .B1(n4650), .B2(ADDR_REG_13__SCAN_IN), .A(n3486), .ZN(n3487) );
  OAI211_X1 U4240 ( .C1(n4657), .C2(n3489), .A(n3488), .B(n3487), .ZN(n3503)
         );
  NOR2_X1 U4241 ( .A1(n3489), .A2(n3372), .ZN(n4116) );
  AOI21_X1 U4242 ( .B1(n3372), .B2(n3489), .A(n4116), .ZN(n3501) );
  NAND2_X1 U4243 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3490), .ZN(n3497) );
  AOI22_X1 U4244 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3490), .B1(n4696), .B2(
        n3283), .ZN(n4586) );
  NAND2_X1 U4245 ( .A1(n4558), .A2(REG2_REG_9__SCAN_IN), .ZN(n3494) );
  MUX2_X1 U4246 ( .A(REG2_REG_9__SCAN_IN), .B(n3951), .S(n4558), .Z(n4563) );
  INV_X1 U4247 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4660) );
  OAI22_X1 U4248 ( .A1(n3493), .A2(n4660), .B1(n3492), .B2(n3491), .ZN(n4564)
         );
  NAND2_X1 U4249 ( .A1(n4563), .A2(n4564), .ZN(n4562) );
  NAND2_X1 U4250 ( .A1(n4571), .A2(n3495), .ZN(n3496) );
  NAND2_X1 U4251 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U4252 ( .A1(n4592), .A2(n3498), .ZN(n3499) );
  OAI21_X1 U4253 ( .B1(n3501), .B2(n4117), .A(n4631), .ZN(n3500) );
  AOI21_X1 U4254 ( .B1(n3501), .B2(n4117), .A(n3500), .ZN(n3502) );
  OR2_X1 U4255 ( .A1(n3503), .A2(n3502), .ZN(U3253) );
  AOI22_X1 U4256 ( .A1(n4378), .A2(n4475), .B1(n4473), .B2(n3523), .ZN(n3504)
         );
  OAI211_X1 U4257 ( .C1(n3755), .C2(n4478), .A(n3505), .B(n3504), .ZN(n3506)
         );
  AOI21_X1 U4258 ( .B1(n3507), .B2(n4713), .A(n3506), .ZN(n3511) );
  MUX2_X1 U4259 ( .A(n3511), .B(n3508), .S(n4718), .Z(n3509) );
  OAI21_X1 U4260 ( .B1(n3513), .B2(n4520), .A(n3509), .ZN(U3497) );
  INV_X1 U4261 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3510) );
  MUX2_X1 U4262 ( .A(n3511), .B(n3510), .S(n4724), .Z(n3512) );
  OAI21_X1 U4263 ( .B1(n4486), .B2(n3513), .A(n3512), .ZN(U3533) );
  OAI22_X1 U4264 ( .A1(n4404), .A2(n3599), .B1(n4170), .B2(n2910), .ZN(n3514)
         );
  XNOR2_X1 U4265 ( .A(n3514), .B(n3613), .ZN(n3516) );
  INV_X1 U4266 ( .A(n3610), .ZN(n3596) );
  OAI22_X1 U4267 ( .A1(n4404), .A2(n2910), .B1(n4170), .B2(n3596), .ZN(n3515)
         );
  XNOR2_X1 U4268 ( .A(n3516), .B(n3515), .ZN(n3623) );
  INV_X1 U4269 ( .A(n3623), .ZN(n3517) );
  NOR2_X1 U4270 ( .A1(n3520), .A2(n3519), .ZN(n3528) );
  AOI22_X1 U4271 ( .A1(n4476), .A2(n3609), .B1(n3523), .B2(n3610), .ZN(n3521)
         );
  XOR2_X1 U4272 ( .A(n3521), .B(n3597), .Z(n3677) );
  OR2_X1 U4273 ( .A1(n3528), .A2(n3677), .ZN(n3522) );
  NOR2_X1 U4274 ( .A1(n3529), .A2(n3522), .ZN(n3527) );
  NAND2_X1 U4275 ( .A1(n4476), .A2(n3344), .ZN(n3525) );
  NAND2_X1 U4276 ( .A1(n3523), .A2(n3609), .ZN(n3524) );
  NAND2_X1 U4277 ( .A1(n3525), .A2(n3524), .ZN(n3750) );
  INV_X1 U4278 ( .A(n3750), .ZN(n3526) );
  INV_X1 U4279 ( .A(n3676), .ZN(n3534) );
  NAND2_X1 U4280 ( .A1(n4378), .A2(n3609), .ZN(n3531) );
  NAND2_X1 U4281 ( .A1(n3683), .A2(n3610), .ZN(n3530) );
  NAND2_X1 U4282 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XNOR2_X1 U4283 ( .A(n3532), .B(n3597), .ZN(n3536) );
  AOI22_X1 U4284 ( .A1(n4378), .A2(n3544), .B1(n3683), .B2(n3609), .ZN(n3537)
         );
  XOR2_X1 U4285 ( .A(n3536), .B(n3537), .Z(n3679) );
  INV_X1 U4286 ( .A(n3679), .ZN(n3533) );
  INV_X1 U4287 ( .A(n3536), .ZN(n3538) );
  NAND2_X1 U4288 ( .A1(n3538), .A2(n3537), .ZN(n3539) );
  NAND2_X1 U4289 ( .A1(n3682), .A2(n3609), .ZN(n3542) );
  NAND2_X1 U4290 ( .A1(n4460), .A2(n3610), .ZN(n3541) );
  NAND2_X1 U4291 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  XNOR2_X1 U4292 ( .A(n3543), .B(n3597), .ZN(n3690) );
  NAND2_X1 U4293 ( .A1(n3682), .A2(n3544), .ZN(n3546) );
  NAND2_X1 U4294 ( .A1(n4460), .A2(n3609), .ZN(n3545) );
  NAND2_X1 U4295 ( .A1(n3546), .A2(n3545), .ZN(n3548) );
  NOR2_X1 U4296 ( .A1(n3690), .A2(n3548), .ZN(n3547) );
  INV_X1 U4297 ( .A(n3548), .ZN(n3689) );
  NAND2_X1 U4298 ( .A1(n4461), .A2(n3609), .ZN(n3551) );
  NAND2_X1 U4299 ( .A1(n4356), .A2(n3610), .ZN(n3550) );
  NAND2_X1 U4300 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  XNOR2_X1 U4301 ( .A(n3552), .B(n3613), .ZN(n3555) );
  NOR2_X1 U4302 ( .A1(n4352), .A2(n2910), .ZN(n3553) );
  AOI21_X1 U4303 ( .B1(n4461), .B2(n3544), .A(n3553), .ZN(n3554) );
  NOR2_X1 U4304 ( .A1(n3555), .A2(n3554), .ZN(n3727) );
  NAND2_X1 U4305 ( .A1(n3555), .A2(n3554), .ZN(n3728) );
  NAND2_X1 U4306 ( .A1(n4357), .A2(n3609), .ZN(n3557) );
  NAND2_X1 U4307 ( .A1(n3648), .A2(n3610), .ZN(n3556) );
  NAND2_X1 U4308 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  XNOR2_X1 U4309 ( .A(n3558), .B(n3597), .ZN(n3559) );
  AOI22_X1 U4310 ( .A1(n4357), .A2(n3344), .B1(n3648), .B2(n3609), .ZN(n3560)
         );
  XNOR2_X1 U4311 ( .A(n3559), .B(n3560), .ZN(n3647) );
  NAND2_X1 U4312 ( .A1(n3646), .A2(n3647), .ZN(n3563) );
  INV_X1 U4313 ( .A(n3559), .ZN(n3561) );
  NAND2_X1 U4314 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  NAND2_X1 U4315 ( .A1(n4333), .A2(n3609), .ZN(n3565) );
  NAND2_X1 U4316 ( .A1(n4444), .A2(n3610), .ZN(n3564) );
  NAND2_X1 U4317 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  XNOR2_X1 U4318 ( .A(n3566), .B(n3597), .ZN(n3573) );
  NAND2_X1 U4319 ( .A1(n4333), .A2(n3344), .ZN(n3568) );
  NAND2_X1 U4320 ( .A1(n4444), .A2(n3609), .ZN(n3567) );
  NAND2_X1 U4321 ( .A1(n3568), .A2(n3567), .ZN(n3574) );
  NAND2_X1 U4322 ( .A1(n3573), .A2(n3574), .ZN(n3708) );
  NOR2_X1 U4323 ( .A1(n3615), .A2(n4295), .ZN(n3569) );
  AOI21_X1 U4324 ( .B1(n4445), .B2(n3344), .A(n3569), .ZN(n3656) );
  NAND2_X1 U4325 ( .A1(n4445), .A2(n3609), .ZN(n3571) );
  NAND2_X1 U4326 ( .A1(n4435), .A2(n3610), .ZN(n3570) );
  NAND2_X1 U4327 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  XNOR2_X1 U4328 ( .A(n3572), .B(n3613), .ZN(n3655) );
  INV_X1 U4329 ( .A(n3573), .ZN(n3576) );
  INV_X1 U4330 ( .A(n3574), .ZN(n3575) );
  AOI21_X1 U4331 ( .B1(n3656), .B2(n3655), .A(n3707), .ZN(n3578) );
  NOR2_X1 U4332 ( .A1(n3655), .A2(n3656), .ZN(n3577) );
  OAI22_X1 U4333 ( .A1(n3661), .A2(n3599), .B1(n4282), .B2(n3615), .ZN(n3580)
         );
  OAI22_X1 U4334 ( .A1(n3661), .A2(n2910), .B1(n4282), .B2(n3596), .ZN(n3579)
         );
  XNOR2_X1 U4335 ( .A(n3579), .B(n3597), .ZN(n3581) );
  XOR2_X1 U4336 ( .A(n3580), .B(n3581), .Z(n3718) );
  NOR2_X1 U4337 ( .A1(n3581), .A2(n3580), .ZN(n3637) );
  NAND2_X1 U4338 ( .A1(n4279), .A2(n3609), .ZN(n3583) );
  NAND2_X1 U4339 ( .A1(n4259), .A2(n3610), .ZN(n3582) );
  NAND2_X1 U4340 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  XNOR2_X1 U4341 ( .A(n3584), .B(n3613), .ZN(n3588) );
  NOR2_X1 U4342 ( .A1(n3615), .A2(n4254), .ZN(n3585) );
  AOI21_X1 U4343 ( .B1(n4279), .B2(n3344), .A(n3585), .ZN(n3587) );
  XNOR2_X1 U4344 ( .A(n3588), .B(n3587), .ZN(n3636) );
  NOR2_X1 U4345 ( .A1(n3637), .A2(n3636), .ZN(n3586) );
  NAND2_X1 U4346 ( .A1(n3635), .A2(n3586), .ZN(n3640) );
  NOR2_X1 U4347 ( .A1(n3588), .A2(n3587), .ZN(n3592) );
  INV_X1 U4348 ( .A(n3592), .ZN(n3589) );
  NAND2_X1 U4349 ( .A1(n3640), .A2(n3589), .ZN(n3590) );
  OAI22_X1 U4350 ( .A1(n4255), .A2(n3599), .B1(n3615), .B2(n4241), .ZN(n3591)
         );
  NAND2_X1 U4351 ( .A1(n3590), .A2(n3591), .ZN(n3698) );
  NAND2_X1 U4352 ( .A1(n3640), .A2(n3593), .ZN(n3697) );
  OAI22_X1 U4353 ( .A1(n4255), .A2(n3615), .B1(n3596), .B2(n4241), .ZN(n3594)
         );
  XNOR2_X1 U4354 ( .A(n3594), .B(n3597), .ZN(n3700) );
  NAND2_X1 U4355 ( .A1(n3697), .A2(n3700), .ZN(n3595) );
  NAND2_X1 U4356 ( .A1(n3698), .A2(n3595), .ZN(n3668) );
  OAI22_X1 U4357 ( .A1(n4198), .A2(n3615), .B1(n3596), .B2(n4221), .ZN(n3598)
         );
  XNOR2_X1 U4358 ( .A(n3598), .B(n3597), .ZN(n3601) );
  OAI22_X1 U4359 ( .A1(n4198), .A2(n3599), .B1(n3615), .B2(n4221), .ZN(n3600)
         );
  OR2_X1 U4360 ( .A1(n3601), .A2(n3600), .ZN(n3667) );
  NAND2_X1 U4361 ( .A1(n3668), .A2(n3667), .ZN(n3602) );
  NAND2_X1 U4362 ( .A1(n3601), .A2(n3600), .ZN(n3666) );
  NAND2_X1 U4363 ( .A1(n4401), .A2(n3609), .ZN(n3604) );
  NAND2_X1 U4364 ( .A1(n4203), .A2(n3610), .ZN(n3603) );
  NAND2_X1 U4365 ( .A1(n3604), .A2(n3603), .ZN(n3605) );
  XNOR2_X1 U4366 ( .A(n3605), .B(n3613), .ZN(n3608) );
  NOR2_X1 U4367 ( .A1(n2910), .A2(n4197), .ZN(n3606) );
  AOI21_X1 U4368 ( .B1(n4401), .B2(n3344), .A(n3606), .ZN(n3607) );
  NOR2_X1 U4369 ( .A1(n3608), .A2(n3607), .ZN(n3738) );
  NAND2_X1 U4370 ( .A1(n3608), .A2(n3607), .ZN(n3737) );
  NAND2_X1 U4371 ( .A1(n4200), .A2(n3609), .ZN(n3612) );
  NAND2_X1 U4372 ( .A1(n4399), .A2(n3610), .ZN(n3611) );
  NAND2_X1 U4373 ( .A1(n3612), .A2(n3611), .ZN(n3614) );
  XNOR2_X1 U4374 ( .A(n3614), .B(n3613), .ZN(n3618) );
  NOR2_X1 U4375 ( .A1(n3615), .A2(n4186), .ZN(n3616) );
  AOI21_X1 U4376 ( .B1(n4200), .B2(n3344), .A(n3616), .ZN(n3617) );
  XNOR2_X1 U4377 ( .A(n3618), .B(n3617), .ZN(n3627) );
  OR2_X1 U4378 ( .A1(n3618), .A2(n3617), .ZN(n3622) );
  AOI22_X1 U4379 ( .A1(n4166), .A2(n3759), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3621) );
  NAND2_X1 U4380 ( .A1(n3720), .A2(n3619), .ZN(n3620) );
  OAI211_X1 U4381 ( .C1(n3824), .C2(n3754), .A(n3621), .B(n3620), .ZN(n3625)
         );
  NOR3_X1 U4382 ( .A1(n3623), .A2(n3747), .A3(n3622), .ZN(n3624) );
  AOI211_X1 U4383 ( .C1(n4167), .C2(n3745), .A(n3625), .B(n3624), .ZN(n3626)
         );
  XNOR2_X1 U4384 ( .A(n3628), .B(n3627), .ZN(n3634) );
  INV_X1 U4385 ( .A(n3629), .ZN(n4184) );
  INV_X1 U4386 ( .A(n4401), .ZN(n4216) );
  OAI22_X1 U4387 ( .A1(n2054), .A2(n4186), .B1(n4216), .B2(n3754), .ZN(n3632)
         );
  OAI22_X1 U4388 ( .A1(n4404), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3630), 
        .ZN(n3631) );
  AOI211_X1 U4389 ( .C1(n4184), .C2(n3745), .A(n3632), .B(n3631), .ZN(n3633)
         );
  OAI21_X1 U4390 ( .B1(n3634), .B2(n3747), .A(n3633), .ZN(U3211) );
  INV_X1 U4391 ( .A(n3635), .ZN(n3638) );
  OAI21_X1 U4392 ( .B1(n3638), .B2(n3637), .A(n3636), .ZN(n3639) );
  NAND3_X1 U4393 ( .A1(n3640), .A2(n3639), .A3(n3752), .ZN(n3645) );
  OAI22_X1 U4394 ( .A1(n2054), .A2(n4254), .B1(n3661), .B2(n3754), .ZN(n3643)
         );
  OAI22_X1 U4395 ( .A1(n4255), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3641), 
        .ZN(n3642) );
  NOR2_X1 U4396 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  OAI211_X1 U4397 ( .C1(n3763), .C2(n4262), .A(n3645), .B(n3644), .ZN(U3213)
         );
  XOR2_X1 U4398 ( .A(n3647), .B(n3646), .Z(n3653) );
  INV_X1 U4399 ( .A(n4342), .ZN(n3651) );
  INV_X1 U4400 ( .A(n4333), .ZN(n4439) );
  AOI22_X1 U4401 ( .A1(n3720), .A2(n3648), .B1(n3719), .B2(n4461), .ZN(n3649)
         );
  NAND2_X1 U4402 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4145) );
  OAI211_X1 U4403 ( .C1(n4439), .C2(n3742), .A(n3649), .B(n4145), .ZN(n3650)
         );
  AOI21_X1 U4404 ( .B1(n3651), .B2(n3745), .A(n3650), .ZN(n3652) );
  OAI21_X1 U4405 ( .B1(n3653), .B2(n3747), .A(n3652), .ZN(U3216) );
  OAI21_X1 U4406 ( .B1(n3654), .B2(n3707), .A(n3708), .ZN(n3658) );
  XOR2_X1 U4407 ( .A(n3656), .B(n3655), .Z(n3657) );
  XNOR2_X1 U4408 ( .A(n3658), .B(n3657), .ZN(n3665) );
  INV_X1 U4409 ( .A(n3659), .ZN(n4292) );
  OAI22_X1 U4410 ( .A1(n3661), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3660), 
        .ZN(n3663) );
  OAI22_X1 U4411 ( .A1(n2054), .A2(n4295), .B1(n4439), .B2(n3754), .ZN(n3662)
         );
  AOI211_X1 U4412 ( .C1(n4292), .C2(n3745), .A(n3663), .B(n3662), .ZN(n3664)
         );
  OAI21_X1 U4413 ( .B1(n3665), .B2(n3747), .A(n3664), .ZN(U3220) );
  NAND2_X1 U4414 ( .A1(n3667), .A2(n3666), .ZN(n3669) );
  XOR2_X1 U4415 ( .A(n3669), .B(n3668), .Z(n3675) );
  INV_X1 U4416 ( .A(n3670), .ZN(n4224) );
  OAI22_X1 U4417 ( .A1(n4216), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3671), 
        .ZN(n3673) );
  OAI22_X1 U4418 ( .A1(n2054), .A2(n4221), .B1(n4255), .B2(n3754), .ZN(n3672)
         );
  AOI211_X1 U4419 ( .C1(n4224), .C2(n3745), .A(n3673), .B(n3672), .ZN(n3674)
         );
  OAI21_X1 U4420 ( .B1(n3675), .B2(n3747), .A(n3674), .ZN(U3222) );
  OR2_X1 U4421 ( .A1(n3678), .A2(n3677), .ZN(n3749) );
  OAI21_X1 U4422 ( .B1(n3676), .B2(n3750), .A(n3749), .ZN(n3680) );
  XNOR2_X1 U4423 ( .A(n3680), .B(n3679), .ZN(n3688) );
  INV_X1 U4424 ( .A(n3681), .ZN(n3686) );
  INV_X1 U4425 ( .A(n3682), .ZN(n4359) );
  AOI22_X1 U4426 ( .A1(n3720), .A2(n3683), .B1(n3719), .B2(n4476), .ZN(n3684)
         );
  NAND2_X1 U4427 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4632) );
  OAI211_X1 U4428 ( .C1(n4359), .C2(n3742), .A(n3684), .B(n4632), .ZN(n3685)
         );
  AOI21_X1 U4429 ( .B1(n3686), .B2(n3745), .A(n3685), .ZN(n3687) );
  OAI21_X1 U4430 ( .B1(n3688), .B2(n3747), .A(n3687), .ZN(U3223) );
  XNOR2_X1 U4431 ( .A(n3690), .B(n3689), .ZN(n3691) );
  XNOR2_X1 U4432 ( .A(n3692), .B(n3691), .ZN(n3693) );
  NAND2_X1 U4433 ( .A1(n3693), .A2(n3752), .ZN(n3696) );
  NOR2_X1 U4434 ( .A1(STATE_REG_SCAN_IN), .A2(n2453), .ZN(n4640) );
  INV_X1 U4435 ( .A(n4378), .ZN(n4464) );
  OAI22_X1 U4436 ( .A1(n2054), .A2(n4386), .B1(n4464), .B2(n3754), .ZN(n3694)
         );
  AOI211_X1 U4437 ( .C1(n3759), .C2(n4461), .A(n4640), .B(n3694), .ZN(n3695)
         );
  OAI211_X1 U4438 ( .C1(n3763), .C2(n4380), .A(n3696), .B(n3695), .ZN(U3225)
         );
  NAND2_X1 U4439 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  XOR2_X1 U4440 ( .A(n3700), .B(n3699), .Z(n3706) );
  INV_X1 U4441 ( .A(n3701), .ZN(n4238) );
  INV_X1 U4442 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3702) );
  OAI22_X1 U4443 ( .A1(n4198), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3702), 
        .ZN(n3704) );
  OAI22_X1 U4444 ( .A1(n2054), .A2(n4241), .B1(n4421), .B2(n3754), .ZN(n3703)
         );
  AOI211_X1 U4445 ( .C1(n4238), .C2(n3745), .A(n3704), .B(n3703), .ZN(n3705)
         );
  OAI21_X1 U4446 ( .B1(n3706), .B2(n3747), .A(n3705), .ZN(U3226) );
  INV_X1 U4447 ( .A(n3707), .ZN(n3709) );
  NAND2_X1 U4448 ( .A1(n3709), .A2(n3708), .ZN(n3710) );
  XNOR2_X1 U4449 ( .A(n3654), .B(n3710), .ZN(n3716) );
  INV_X1 U4450 ( .A(n3711), .ZN(n4312) );
  INV_X1 U4451 ( .A(n4445), .ZN(n4314) );
  INV_X1 U4452 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3712) );
  OAI22_X1 U4453 ( .A1(n4314), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3712), 
        .ZN(n3714) );
  INV_X1 U4454 ( .A(n4357), .ZN(n4448) );
  OAI22_X1 U4455 ( .A1(n2054), .A2(n4316), .B1(n4448), .B2(n3754), .ZN(n3713)
         );
  AOI211_X1 U4456 ( .C1(n4312), .C2(n3745), .A(n3714), .B(n3713), .ZN(n3715)
         );
  OAI21_X1 U4457 ( .B1(n3716), .B2(n3747), .A(n3715), .ZN(U3230) );
  OAI21_X1 U4458 ( .B1(n3718), .B2(n3717), .A(n3635), .ZN(n3724) );
  AOI22_X1 U4459 ( .A1(n3720), .A2(n2512), .B1(n3719), .B2(n4445), .ZN(n3722)
         );
  AOI22_X1 U4460 ( .A1(n3759), .A2(n4279), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3721) );
  OAI211_X1 U4461 ( .C1(n3763), .C2(n4274), .A(n3722), .B(n3721), .ZN(n3723)
         );
  AOI21_X1 U4462 ( .B1(n3724), .B2(n3752), .A(n3723), .ZN(n3725) );
  INV_X1 U4463 ( .A(n3725), .ZN(U3232) );
  INV_X1 U4464 ( .A(n3727), .ZN(n3729) );
  NAND2_X1 U4465 ( .A1(n3729), .A2(n3728), .ZN(n3730) );
  XNOR2_X1 U4466 ( .A(n3726), .B(n3730), .ZN(n3731) );
  NAND2_X1 U4467 ( .A1(n3731), .A2(n3752), .ZN(n3735) );
  NOR2_X1 U4468 ( .A1(STATE_REG_SCAN_IN), .A2(n3732), .ZN(n4649) );
  OAI22_X1 U4469 ( .A1(n2054), .A2(n4352), .B1(n4359), .B2(n3754), .ZN(n3733)
         );
  AOI211_X1 U4470 ( .C1(n3759), .C2(n4357), .A(n4649), .B(n3733), .ZN(n3734)
         );
  OAI211_X1 U4471 ( .C1(n3763), .C2(n4363), .A(n3735), .B(n3734), .ZN(U3235)
         );
  NOR2_X1 U4472 ( .A1(n3738), .A2(n2174), .ZN(n3739) );
  XNOR2_X1 U4473 ( .A(n3736), .B(n3739), .ZN(n3748) );
  INV_X1 U4474 ( .A(n3740), .ZN(n4206) );
  OAI22_X1 U4475 ( .A1(n2054), .A2(n4197), .B1(n4198), .B2(n3754), .ZN(n3744)
         );
  OAI22_X1 U4476 ( .A1(n3824), .A2(n3742), .B1(STATE_REG_SCAN_IN), .B2(n3741), 
        .ZN(n3743) );
  AOI211_X1 U4477 ( .C1(n4206), .C2(n3745), .A(n3744), .B(n3743), .ZN(n3746)
         );
  OAI21_X1 U4478 ( .B1(n3748), .B2(n3747), .A(n3746), .ZN(U3237) );
  NAND2_X1 U4479 ( .A1(n3534), .A2(n3749), .ZN(n3751) );
  XNOR2_X1 U4480 ( .A(n3751), .B(n3750), .ZN(n3753) );
  NAND2_X1 U4481 ( .A1(n3753), .A2(n3752), .ZN(n3761) );
  AND2_X1 U4482 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4616) );
  OAI22_X1 U4483 ( .A1(n2054), .A2(n3756), .B1(n3755), .B2(n3754), .ZN(n3758)
         );
  AOI211_X1 U4484 ( .C1(n3759), .C2(n4378), .A(n4616), .B(n3758), .ZN(n3760)
         );
  OAI211_X1 U4485 ( .C1(n3763), .C2(n3762), .A(n3761), .B(n3760), .ZN(U3238)
         );
  OAI211_X1 U4486 ( .C1(n3766), .C2(n3907), .A(n3765), .B(n3764), .ZN(n3767)
         );
  NAND3_X1 U4487 ( .A1(n3767), .A2(n2578), .A3(n2577), .ZN(n3770) );
  NAND3_X1 U4488 ( .A1(n3770), .A2(n3769), .A3(n3768), .ZN(n3773) );
  NAND3_X1 U4489 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3776) );
  NAND4_X1 U4490 ( .A1(n3776), .A2(n3775), .A3(n3790), .A4(n3774), .ZN(n3778)
         );
  NAND3_X1 U4491 ( .A1(n3778), .A2(n3873), .A3(n3777), .ZN(n3779) );
  NAND3_X1 U4492 ( .A1(n3779), .A2(n3787), .A3(n3791), .ZN(n3782) );
  AND3_X1 U4493 ( .A1(n3782), .A2(n3781), .A3(n3780), .ZN(n3786) );
  NAND2_X1 U4494 ( .A1(n3784), .A2(n3783), .ZN(n3794) );
  NOR3_X1 U4495 ( .A1(n3786), .A2(n3785), .A3(n3794), .ZN(n3801) );
  INV_X1 U4496 ( .A(n3787), .ZN(n3789) );
  NOR2_X1 U4497 ( .A1(n3789), .A2(n3788), .ZN(n3793) );
  NAND4_X1 U4498 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3796)
         );
  NAND2_X1 U4499 ( .A1(n3794), .A2(n3803), .ZN(n3879) );
  INV_X1 U4500 ( .A(n3879), .ZN(n3795) );
  AOI21_X1 U4501 ( .B1(n3797), .B2(n3796), .A(n3795), .ZN(n3800) );
  OAI211_X1 U4502 ( .C1(n3801), .C2(n3800), .A(n3799), .B(n3798), .ZN(n3806)
         );
  NAND2_X1 U4503 ( .A1(n3804), .A2(n3803), .ZN(n3880) );
  OAI21_X1 U4504 ( .B1(n2095), .B2(n3880), .A(n3879), .ZN(n3805) );
  AOI21_X1 U4505 ( .B1(n3806), .B2(n3805), .A(n2102), .ZN(n3809) );
  INV_X1 U4506 ( .A(n3882), .ZN(n3808) );
  INV_X1 U4507 ( .A(n3807), .ZN(n3884) );
  OAI211_X1 U4508 ( .C1(n3809), .C2(n3808), .A(n2082), .B(n3884), .ZN(n3811)
         );
  INV_X1 U4509 ( .A(n3810), .ZN(n3887) );
  AOI211_X1 U4510 ( .C1(n3811), .C2(n3888), .A(n3887), .B(n4248), .ZN(n3812)
         );
  NOR2_X1 U4511 ( .A1(n3812), .A2(n3891), .ZN(n3814) );
  OAI21_X1 U4512 ( .B1(n3814), .B2(n3813), .A(n3894), .ZN(n3817) );
  INV_X1 U4513 ( .A(n3815), .ZN(n3897) );
  AOI21_X1 U4514 ( .B1(n3817), .B2(n3816), .A(n3897), .ZN(n3835) );
  NAND2_X1 U4515 ( .A1(n4166), .A2(n4163), .ZN(n3818) );
  AND2_X1 U4516 ( .A1(n3819), .A2(n3818), .ZN(n3833) );
  INV_X1 U4517 ( .A(n3833), .ZN(n3822) );
  INV_X1 U4518 ( .A(n3820), .ZN(n3821) );
  OR2_X1 U4519 ( .A1(n3822), .A2(n3821), .ZN(n3901) );
  INV_X1 U4520 ( .A(n3901), .ZN(n3823) );
  OAI21_X1 U4521 ( .B1(n3824), .B2(n4399), .A(n3823), .ZN(n3834) );
  NAND2_X1 U4522 ( .A1(n3826), .A2(n3825), .ZN(n3898) );
  AND2_X1 U4523 ( .A1(n3831), .A2(DATAI_30_), .ZN(n4396) );
  NAND2_X1 U4524 ( .A1(n3836), .A2(n4396), .ZN(n3832) );
  INV_X1 U4525 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U4526 ( .A1(n3827), .A2(REG2_REG_31__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4527 ( .A1(n3828), .A2(REG1_REG_31__SCAN_IN), .ZN(n3829) );
  OAI211_X1 U4528 ( .C1(n2342), .C2(n4488), .A(n3830), .B(n3829), .ZN(n3926)
         );
  NAND2_X1 U4529 ( .A1(n3831), .A2(DATAI_31_), .ZN(n4151) );
  NAND2_X1 U4530 ( .A1(n3926), .A2(n4151), .ZN(n3838) );
  AND2_X1 U4531 ( .A1(n3832), .A2(n3838), .ZN(n3849) );
  OAI21_X1 U4532 ( .B1(n4166), .B2(n4163), .A(n3849), .ZN(n3896) );
  AOI21_X1 U4533 ( .B1(n3833), .B2(n3898), .A(n3896), .ZN(n3900) );
  OAI21_X1 U4534 ( .B1(n3835), .B2(n3834), .A(n3900), .ZN(n3841) );
  OR2_X1 U4535 ( .A1(n3836), .A2(n4396), .ZN(n3904) );
  OR2_X1 U4536 ( .A1(n3926), .A2(n4151), .ZN(n3837) );
  AND2_X1 U4537 ( .A1(n3904), .A2(n3837), .ZN(n3850) );
  INV_X1 U4538 ( .A(n3850), .ZN(n3839) );
  NAND2_X1 U4539 ( .A1(n3839), .A2(n3838), .ZN(n3840) );
  NAND2_X1 U4540 ( .A1(n3841), .A2(n3840), .ZN(n3915) );
  NAND4_X1 U4541 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3855)
         );
  AND2_X1 U4542 ( .A1(n4193), .A2(n3846), .ZN(n4214) );
  NAND2_X1 U4543 ( .A1(n4212), .A2(n3847), .ZN(n4235) );
  INV_X1 U4544 ( .A(n4235), .ZN(n4231) );
  NAND2_X1 U4545 ( .A1(n2076), .A2(n3848), .ZN(n4196) );
  NAND4_X1 U4546 ( .A1(n4214), .A2(n4231), .A3(n3849), .A4(n4196), .ZN(n3854)
         );
  NAND4_X1 U4547 ( .A1(n3852), .A2(n3851), .A3(n4181), .A4(n3850), .ZN(n3853)
         );
  NOR3_X1 U4548 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3858) );
  NAND2_X1 U4549 ( .A1(n3857), .A2(n3856), .ZN(n4307) );
  NAND4_X1 U4550 ( .A1(n3859), .A2(n4354), .A3(n3858), .A4(n4307), .ZN(n3862)
         );
  NOR3_X1 U4551 ( .A1(n3862), .A2(n3861), .A3(n3860), .ZN(n3871) );
  NOR4_X1 U4552 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n2575), .ZN(n3870)
         );
  INV_X1 U4553 ( .A(n4248), .ZN(n3866) );
  NAND2_X1 U4554 ( .A1(n3866), .A2(n4249), .ZN(n4289) );
  NAND2_X1 U4555 ( .A1(n3884), .A2(n4324), .ZN(n4373) );
  NOR4_X1 U4556 ( .A1(n4289), .A2(n4373), .A3(n3868), .A4(n3867), .ZN(n3869)
         );
  NAND3_X1 U4557 ( .A1(n3871), .A2(n3870), .A3(n3869), .ZN(n3878) );
  XNOR2_X1 U4558 ( .A(n4279), .B(n4259), .ZN(n4246) );
  INV_X1 U4559 ( .A(n4246), .ZN(n4252) );
  NAND4_X1 U4560 ( .A1(n4270), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3877)
         );
  XNOR2_X1 U4561 ( .A(n4357), .B(n4339), .ZN(n4323) );
  INV_X1 U4562 ( .A(n4323), .ZN(n4329) );
  NAND2_X1 U4563 ( .A1(n4329), .A2(n3875), .ZN(n3876) );
  NOR4_X1 U4564 ( .A1(n3878), .A2(n4252), .A3(n3877), .A4(n3876), .ZN(n3909)
         );
  OAI21_X1 U4565 ( .B1(n3881), .B2(n3880), .A(n3879), .ZN(n3883) );
  NAND2_X1 U4566 ( .A1(n3883), .A2(n3882), .ZN(n3886) );
  NAND4_X1 U4567 ( .A1(n3886), .A2(n2082), .A3(n3885), .A4(n3884), .ZN(n3889)
         );
  AOI21_X1 U4568 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n3892) );
  OAI21_X1 U4569 ( .B1(n3892), .B2(n3891), .A(n3890), .ZN(n3895) );
  AOI21_X1 U4570 ( .B1(n3895), .B2(n3894), .A(n3893), .ZN(n3899) );
  OAI21_X1 U4571 ( .B1(n3901), .B2(n4176), .A(n3900), .ZN(n3902) );
  INV_X1 U4572 ( .A(n3926), .ZN(n4153) );
  AOI22_X1 U4573 ( .A1(n3903), .A2(n3902), .B1(n4153), .B2(n4396), .ZN(n3906)
         );
  AOI21_X1 U4574 ( .B1(n3904), .B2(n3926), .A(n4151), .ZN(n3905) );
  NOR2_X1 U4575 ( .A1(n3906), .A2(n3905), .ZN(n3908) );
  MUX2_X1 U4576 ( .A(n3909), .B(n3908), .S(n3907), .Z(n3910) );
  NOR2_X1 U4577 ( .A1(n3910), .A2(n3911), .ZN(n3913) );
  AOI21_X1 U4578 ( .B1(n3911), .B2(n3915), .A(n3913), .ZN(n3912) );
  MUX2_X1 U4579 ( .A(n3913), .B(n3912), .S(n4146), .Z(n3914) );
  AOI21_X1 U4580 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3924) );
  INV_X1 U4581 ( .A(n3917), .ZN(n3919) );
  NOR2_X1 U4582 ( .A1(n3919), .A2(n3918), .ZN(n3922) );
  OAI21_X1 U4583 ( .B1(n3923), .B2(n3920), .A(B_REG_SCAN_IN), .ZN(n3921) );
  OAI22_X1 U4584 ( .A1(n3924), .A2(n3923), .B1(n3922), .B2(n3921), .ZN(U3239)
         );
  MUX2_X1 U4585 ( .A(n3926), .B(DATAO_REG_31__SCAN_IN), .S(n3925), .Z(U3581)
         );
  MUX2_X1 U4586 ( .A(DATAO_REG_29__SCAN_IN), .B(n4166), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4587 ( .A(DATAO_REG_28__SCAN_IN), .B(n4161), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4588 ( .A(DATAO_REG_26__SCAN_IN), .B(n4401), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4589 ( .A(DATAO_REG_24__SCAN_IN), .B(n4218), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4590 ( .A(DATAO_REG_22__SCAN_IN), .B(n4436), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4591 ( .A(DATAO_REG_21__SCAN_IN), .B(n4445), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4592 ( .A(DATAO_REG_19__SCAN_IN), .B(n4357), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4593 ( .A(DATAO_REG_18__SCAN_IN), .B(n4461), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4594 ( .A(DATAO_REG_16__SCAN_IN), .B(n4378), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4595 ( .A(DATAO_REG_15__SCAN_IN), .B(n4476), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4596 ( .A(DATAO_REG_13__SCAN_IN), .B(n3927), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4597 ( .A(DATAO_REG_12__SCAN_IN), .B(n3928), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4598 ( .A(DATAO_REG_11__SCAN_IN), .B(n3929), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4599 ( .A(DATAO_REG_10__SCAN_IN), .B(n3930), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4600 ( .A(DATAO_REG_9__SCAN_IN), .B(n3931), .S(U4043), .Z(U3559) );
  MUX2_X1 U4601 ( .A(DATAO_REG_8__SCAN_IN), .B(n3932), .S(U4043), .Z(U3558) );
  MUX2_X1 U4602 ( .A(DATAO_REG_7__SCAN_IN), .B(n3933), .S(U4043), .Z(U3557) );
  MUX2_X1 U4603 ( .A(DATAO_REG_6__SCAN_IN), .B(n3934), .S(U4043), .Z(U3556) );
  MUX2_X1 U4604 ( .A(DATAO_REG_5__SCAN_IN), .B(n3935), .S(U4043), .Z(U3555) );
  MUX2_X1 U4605 ( .A(DATAO_REG_3__SCAN_IN), .B(n3936), .S(U4043), .Z(n4110) );
  INV_X1 U4606 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4607 ( .A1(n3938), .A2(keyinput76), .B1(n4069), .B2(keyinput116), 
        .ZN(n3937) );
  OAI221_X1 U4608 ( .B1(n3938), .B2(keyinput76), .C1(n4069), .C2(keyinput116), 
        .A(n3937), .ZN(n3948) );
  INV_X1 U4609 ( .A(D_REG_8__SCAN_IN), .ZN(n4677) );
  INV_X1 U4610 ( .A(D_REG_9__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U4611 ( .A1(n4677), .A2(keyinput123), .B1(n4676), .B2(keyinput110), 
        .ZN(n3939) );
  OAI221_X1 U4612 ( .B1(n4677), .B2(keyinput123), .C1(n4676), .C2(keyinput110), 
        .A(n3939), .ZN(n3947) );
  INV_X1 U4613 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4614 ( .A1(n3942), .A2(keyinput80), .B1(n3941), .B2(keyinput105), 
        .ZN(n3940) );
  OAI221_X1 U4615 ( .B1(n3942), .B2(keyinput80), .C1(n3941), .C2(keyinput105), 
        .A(n3940), .ZN(n3946) );
  INV_X1 U4616 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n3944) );
  INV_X1 U4617 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U4618 ( .A1(n3944), .A2(keyinput119), .B1(n4634), .B2(keyinput70), 
        .ZN(n3943) );
  OAI221_X1 U4619 ( .B1(n3944), .B2(keyinput119), .C1(n4634), .C2(keyinput70), 
        .A(n3943), .ZN(n3945) );
  NOR4_X1 U4620 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3982)
         );
  INV_X1 U4621 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4137) );
  INV_X1 U4622 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U4623 ( .A1(n4137), .A2(keyinput127), .B1(keyinput104), .B2(n4424), 
        .ZN(n3949) );
  OAI221_X1 U4624 ( .B1(n4137), .B2(keyinput127), .C1(n4424), .C2(keyinput104), 
        .A(n3949), .ZN(n3959) );
  INV_X1 U4625 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4626 ( .A1(n3951), .A2(keyinput121), .B1(n4089), .B2(keyinput87), 
        .ZN(n3950) );
  OAI221_X1 U4627 ( .B1(n3951), .B2(keyinput121), .C1(n4089), .C2(keyinput87), 
        .A(n3950), .ZN(n3958) );
  AOI22_X1 U4628 ( .A1(n3953), .A2(keyinput98), .B1(keyinput126), .B2(n4057), 
        .ZN(n3952) );
  OAI221_X1 U4629 ( .B1(n3953), .B2(keyinput98), .C1(n4057), .C2(keyinput126), 
        .A(n3952), .ZN(n3957) );
  INV_X1 U4630 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4141) );
  INV_X1 U4631 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4632 ( .A1(n4141), .A2(keyinput108), .B1(n3955), .B2(keyinput106), 
        .ZN(n3954) );
  OAI221_X1 U4633 ( .B1(n4141), .B2(keyinput108), .C1(n3955), .C2(keyinput106), 
        .A(n3954), .ZN(n3956) );
  NOR4_X1 U4634 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3981)
         );
  INV_X1 U4635 ( .A(D_REG_5__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U4636 ( .A1(n3210), .A2(keyinput115), .B1(n4679), .B2(keyinput124), 
        .ZN(n3960) );
  OAI221_X1 U4637 ( .B1(n3210), .B2(keyinput115), .C1(n4679), .C2(keyinput124), 
        .A(n3960), .ZN(n3968) );
  INV_X1 U4638 ( .A(D_REG_29__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U4639 ( .A1(n4672), .A2(keyinput67), .B1(keyinput86), .B2(n2267), 
        .ZN(n3961) );
  OAI221_X1 U4640 ( .B1(n4672), .B2(keyinput67), .C1(n2267), .C2(keyinput86), 
        .A(n3961), .ZN(n3967) );
  INV_X1 U4641 ( .A(D_REG_17__SCAN_IN), .ZN(n4674) );
  INV_X1 U4642 ( .A(D_REG_14__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U4643 ( .A1(n4674), .A2(keyinput91), .B1(n4675), .B2(keyinput101), 
        .ZN(n3962) );
  OAI221_X1 U4644 ( .B1(n4674), .B2(keyinput91), .C1(n4675), .C2(keyinput101), 
        .A(n3962), .ZN(n3966) );
  AOI22_X1 U4645 ( .A1(n3964), .A2(keyinput88), .B1(n4078), .B2(keyinput69), 
        .ZN(n3963) );
  OAI221_X1 U4646 ( .B1(n3964), .B2(keyinput88), .C1(n4078), .C2(keyinput69), 
        .A(n3963), .ZN(n3965) );
  NOR4_X1 U4647 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3980)
         );
  INV_X1 U4648 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4649 ( .A1(n4076), .A2(keyinput81), .B1(n2453), .B2(keyinput99), 
        .ZN(n3969) );
  OAI221_X1 U4650 ( .B1(n4076), .B2(keyinput81), .C1(n2453), .C2(keyinput99), 
        .A(n3969), .ZN(n3978) );
  INV_X1 U4651 ( .A(DATAI_9_), .ZN(n3971) );
  AOI22_X1 U4652 ( .A1(n3971), .A2(keyinput65), .B1(n4693), .B2(keyinput84), 
        .ZN(n3970) );
  OAI221_X1 U4653 ( .B1(n3971), .B2(keyinput65), .C1(n4693), .C2(keyinput84), 
        .A(n3970), .ZN(n3977) );
  INV_X1 U4654 ( .A(DATAI_23_), .ZN(n4684) );
  XOR2_X1 U4655 ( .A(n4684), .B(keyinput82), .Z(n3975) );
  XNOR2_X1 U4656 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput112), .ZN(n3974) );
  XNOR2_X1 U4657 ( .A(IR_REG_25__SCAN_IN), .B(keyinput77), .ZN(n3973) );
  XNOR2_X1 U4658 ( .A(IR_REG_20__SCAN_IN), .B(keyinput90), .ZN(n3972) );
  NAND4_X1 U4659 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  NOR3_X1 U4660 ( .A1(n3978), .A2(n3977), .A3(n3976), .ZN(n3979) );
  AND4_X1 U4661 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n4108)
         );
  OAI22_X1 U4662 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput109), .B1(
        DATAO_REG_23__SCAN_IN), .B2(keyinput93), .ZN(n3983) );
  AOI221_X1 U4663 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput109), .C1(
        keyinput93), .C2(DATAO_REG_23__SCAN_IN), .A(n3983), .ZN(n3990) );
  OAI22_X1 U4664 ( .A1(REG1_REG_25__SCAN_IN), .A2(keyinput111), .B1(
        keyinput118), .B2(REG0_REG_30__SCAN_IN), .ZN(n3984) );
  AOI221_X1 U4665 ( .B1(REG1_REG_25__SCAN_IN), .B2(keyinput111), .C1(
        REG0_REG_30__SCAN_IN), .C2(keyinput118), .A(n3984), .ZN(n3989) );
  OAI22_X1 U4666 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput120), .B1(keyinput73), 
        .B2(DATAO_REG_4__SCAN_IN), .ZN(n3985) );
  AOI221_X1 U4667 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput120), .C1(
        DATAO_REG_4__SCAN_IN), .C2(keyinput73), .A(n3985), .ZN(n3988) );
  OAI22_X1 U4668 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput117), .B1(keyinput83), .B2(DATAO_REG_27__SCAN_IN), .ZN(n3986) );
  AOI221_X1 U4669 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput117), .C1(
        DATAO_REG_27__SCAN_IN), .C2(keyinput83), .A(n3986), .ZN(n3987) );
  NAND4_X1 U4670 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n4018)
         );
  OAI22_X1 U4671 ( .A1(REG2_REG_25__SCAN_IN), .A2(keyinput72), .B1(keyinput114), .B2(REG2_REG_7__SCAN_IN), .ZN(n3991) );
  AOI221_X1 U4672 ( .B1(REG2_REG_25__SCAN_IN), .B2(keyinput72), .C1(
        REG2_REG_7__SCAN_IN), .C2(keyinput114), .A(n3991), .ZN(n3998) );
  OAI22_X1 U4673 ( .A1(REG1_REG_29__SCAN_IN), .A2(keyinput122), .B1(keyinput92), .B2(REG2_REG_15__SCAN_IN), .ZN(n3992) );
  AOI221_X1 U4674 ( .B1(REG1_REG_29__SCAN_IN), .B2(keyinput122), .C1(
        REG2_REG_15__SCAN_IN), .C2(keyinput92), .A(n3992), .ZN(n3997) );
  OAI22_X1 U4675 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput64), .B1(
        REG0_REG_24__SCAN_IN), .B2(keyinput113), .ZN(n3993) );
  AOI221_X1 U4676 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput64), .C1(keyinput113), .C2(REG0_REG_24__SCAN_IN), .A(n3993), .ZN(n3996) );
  OAI22_X1 U4677 ( .A1(REG2_REG_20__SCAN_IN), .A2(keyinput78), .B1(
        REG2_REG_16__SCAN_IN), .B2(keyinput68), .ZN(n3994) );
  AOI221_X1 U4678 ( .B1(REG2_REG_20__SCAN_IN), .B2(keyinput78), .C1(keyinput68), .C2(REG2_REG_16__SCAN_IN), .A(n3994), .ZN(n3995) );
  NAND4_X1 U4679 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n4017)
         );
  OAI22_X1 U4680 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput107), .B1(
        REG0_REG_16__SCAN_IN), .B2(keyinput79), .ZN(n3999) );
  AOI221_X1 U4681 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput107), .C1(keyinput79), 
        .C2(REG0_REG_16__SCAN_IN), .A(n3999), .ZN(n4006) );
  OAI22_X1 U4682 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput100), .B1(keyinput125), 
        .B2(D_REG_30__SCAN_IN), .ZN(n4000) );
  AOI221_X1 U4683 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput100), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput125), .A(n4000), .ZN(n4005) );
  OAI22_X1 U4684 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput66), .B1(keyinput97), 
        .B2(D_REG_18__SCAN_IN), .ZN(n4001) );
  AOI221_X1 U4685 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput66), .C1(
        D_REG_18__SCAN_IN), .C2(keyinput97), .A(n4001), .ZN(n4004) );
  OAI22_X1 U4686 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput85), .B1(keyinput75), 
        .B2(REG0_REG_22__SCAN_IN), .ZN(n4002) );
  AOI221_X1 U4687 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput85), .C1(
        REG0_REG_22__SCAN_IN), .C2(keyinput75), .A(n4002), .ZN(n4003) );
  NAND4_X1 U4688 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4016)
         );
  OAI22_X1 U4689 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput94), .B1(DATAI_17_), 
        .B2(keyinput102), .ZN(n4007) );
  AOI221_X1 U4690 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput94), .C1(keyinput102), 
        .C2(DATAI_17_), .A(n4007), .ZN(n4014) );
  OAI22_X1 U4691 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput71), .B1(keyinput89), 
        .B2(REG3_REG_14__SCAN_IN), .ZN(n4008) );
  AOI221_X1 U4692 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput71), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput89), .A(n4008), .ZN(n4013) );
  OAI22_X1 U4693 ( .A1(DATAI_13_), .A2(keyinput74), .B1(keyinput96), .B2(
        DATAI_3_), .ZN(n4009) );
  AOI221_X1 U4694 ( .B1(DATAI_13_), .B2(keyinput74), .C1(DATAI_3_), .C2(
        keyinput96), .A(n4009), .ZN(n4012) );
  OAI22_X1 U4695 ( .A1(DATAI_29_), .A2(keyinput103), .B1(keyinput95), .B2(
        DATAI_30_), .ZN(n4010) );
  AOI221_X1 U4696 ( .B1(DATAI_29_), .B2(keyinput103), .C1(DATAI_30_), .C2(
        keyinput95), .A(n4010), .ZN(n4011) );
  NAND4_X1 U4697 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  NOR4_X1 U4698 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4107)
         );
  AOI22_X1 U4699 ( .A1(ADDR_REG_4__SCAN_IN), .A2(keyinput41), .B1(
        REG2_REG_9__SCAN_IN), .B2(keyinput57), .ZN(n4019) );
  OAI221_X1 U4700 ( .B1(ADDR_REG_4__SCAN_IN), .B2(keyinput41), .C1(
        REG2_REG_9__SCAN_IN), .C2(keyinput57), .A(n4019), .ZN(n4026) );
  AOI22_X1 U4701 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput9), .B1(
        REG0_REG_24__SCAN_IN), .B2(keyinput49), .ZN(n4020) );
  OAI221_X1 U4702 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput9), .C1(
        REG0_REG_24__SCAN_IN), .C2(keyinput49), .A(n4020), .ZN(n4025) );
  AOI22_X1 U4703 ( .A1(DATAI_9_), .A2(keyinput1), .B1(D_REG_14__SCAN_IN), .B2(
        keyinput37), .ZN(n4021) );
  OAI221_X1 U4704 ( .B1(DATAI_9_), .B2(keyinput1), .C1(D_REG_14__SCAN_IN), 
        .C2(keyinput37), .A(n4021), .ZN(n4024) );
  AOI22_X1 U4705 ( .A1(DATAO_REG_23__SCAN_IN), .A2(keyinput29), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput45), .ZN(n4022) );
  OAI221_X1 U4706 ( .B1(DATAO_REG_23__SCAN_IN), .B2(keyinput29), .C1(
        DATAO_REG_20__SCAN_IN), .C2(keyinput45), .A(n4022), .ZN(n4023) );
  NOR4_X1 U4707 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4054)
         );
  AOI22_X1 U4708 ( .A1(REG2_REG_16__SCAN_IN), .A2(keyinput4), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput8), .ZN(n4027) );
  OAI221_X1 U4709 ( .B1(REG2_REG_16__SCAN_IN), .B2(keyinput4), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput8), .A(n4027), .ZN(n4034) );
  AOI22_X1 U4710 ( .A1(ADDR_REG_1__SCAN_IN), .A2(keyinput16), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput25), .ZN(n4028) );
  OAI221_X1 U4711 ( .B1(ADDR_REG_1__SCAN_IN), .B2(keyinput16), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput25), .A(n4028), .ZN(n4033) );
  AOI22_X1 U4712 ( .A1(REG2_REG_15__SCAN_IN), .A2(keyinput28), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput36), .ZN(n4029) );
  OAI221_X1 U4713 ( .B1(REG2_REG_15__SCAN_IN), .B2(keyinput28), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput36), .A(n4029), .ZN(n4032) );
  AOI22_X1 U4714 ( .A1(DATAO_REG_25__SCAN_IN), .A2(keyinput12), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput24), .ZN(n4030) );
  OAI221_X1 U4715 ( .B1(DATAO_REG_25__SCAN_IN), .B2(keyinput12), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput24), .A(n4030), .ZN(n4031) );
  NOR4_X1 U4716 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4053)
         );
  AOI22_X1 U4717 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput50), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput58), .ZN(n4035) );
  OAI221_X1 U4718 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput50), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput58), .A(n4035), .ZN(n4042) );
  AOI22_X1 U4719 ( .A1(REG1_REG_22__SCAN_IN), .A2(keyinput42), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput46), .ZN(n4036) );
  OAI221_X1 U4720 ( .B1(REG1_REG_22__SCAN_IN), .B2(keyinput42), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput46), .A(n4036), .ZN(n4041) );
  AOI22_X1 U4721 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput34), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput26), .ZN(n4037) );
  OAI221_X1 U4722 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput34), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput26), .A(n4037), .ZN(n4040) );
  AOI22_X1 U4723 ( .A1(ADDR_REG_16__SCAN_IN), .A2(keyinput6), .B1(DATAI_13_), 
        .B2(keyinput10), .ZN(n4038) );
  OAI221_X1 U4724 ( .B1(ADDR_REG_16__SCAN_IN), .B2(keyinput6), .C1(DATAI_13_), 
        .C2(keyinput10), .A(n4038), .ZN(n4039) );
  NOR4_X1 U4725 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4052)
         );
  AOI22_X1 U4726 ( .A1(DATAI_3_), .A2(keyinput32), .B1(REG0_REG_16__SCAN_IN), 
        .B2(keyinput15), .ZN(n4043) );
  OAI221_X1 U4727 ( .B1(DATAI_3_), .B2(keyinput32), .C1(REG0_REG_16__SCAN_IN), 
        .C2(keyinput15), .A(n4043), .ZN(n4050) );
  AOI22_X1 U4728 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput56), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput43), .ZN(n4044) );
  OAI221_X1 U4729 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput56), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput43), .A(n4044), .ZN(n4049) );
  AOI22_X1 U4730 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput59), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput27), .ZN(n4045) );
  OAI221_X1 U4731 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput59), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput27), .A(n4045), .ZN(n4048) );
  AOI22_X1 U4732 ( .A1(ADDR_REG_14__SCAN_IN), .A2(keyinput55), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput35), .ZN(n4046) );
  OAI221_X1 U4733 ( .B1(ADDR_REG_14__SCAN_IN), .B2(keyinput55), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput35), .A(n4046), .ZN(n4047) );
  NOR4_X1 U4734 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4051)
         );
  NAND4_X1 U4735 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4106)
         );
  AOI22_X1 U4736 ( .A1(n4137), .A2(keyinput63), .B1(keyinput54), .B2(n2660), 
        .ZN(n4055) );
  OAI221_X1 U4737 ( .B1(n4137), .B2(keyinput63), .C1(n2660), .C2(keyinput54), 
        .A(n4055), .ZN(n4065) );
  AOI22_X1 U4738 ( .A1(n4722), .A2(keyinput0), .B1(keyinput62), .B2(n4057), 
        .ZN(n4056) );
  OAI221_X1 U4739 ( .B1(n4722), .B2(keyinput0), .C1(n4057), .C2(keyinput62), 
        .A(n4056), .ZN(n4064) );
  INV_X1 U4740 ( .A(DATAI_17_), .ZN(n4687) );
  AOI22_X1 U4741 ( .A1(n4059), .A2(keyinput39), .B1(keyinput38), .B2(n4687), 
        .ZN(n4058) );
  OAI221_X1 U4742 ( .B1(n4059), .B2(keyinput39), .C1(n4687), .C2(keyinput38), 
        .A(n4058), .ZN(n4063) );
  INV_X1 U4743 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4744 ( .A1(n3210), .A2(keyinput51), .B1(n4061), .B2(keyinput47), 
        .ZN(n4060) );
  OAI221_X1 U4745 ( .B1(n3210), .B2(keyinput51), .C1(n4061), .C2(keyinput47), 
        .A(n4060), .ZN(n4062) );
  NOR4_X1 U4746 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4104)
         );
  INV_X1 U4747 ( .A(D_REG_30__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U4748 ( .A1(n4671), .A2(keyinput61), .B1(keyinput20), .B2(n4693), 
        .ZN(n4066) );
  OAI221_X1 U4749 ( .B1(n4671), .B2(keyinput61), .C1(n4693), .C2(keyinput20), 
        .A(n4066), .ZN(n4074) );
  AOI22_X1 U4750 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput48), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput7), .ZN(n4067) );
  OAI221_X1 U4751 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput48), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput7), .A(n4067), .ZN(n4073) );
  AOI22_X1 U4752 ( .A1(n4069), .A2(keyinput52), .B1(n4679), .B2(keyinput60), 
        .ZN(n4068) );
  OAI221_X1 U4753 ( .B1(n4069), .B2(keyinput52), .C1(n4679), .C2(keyinput60), 
        .A(n4068), .ZN(n4072) );
  AOI22_X1 U4754 ( .A1(n4141), .A2(keyinput44), .B1(keyinput40), .B2(n4424), 
        .ZN(n4070) );
  OAI221_X1 U4755 ( .B1(n4141), .B2(keyinput44), .C1(n4424), .C2(keyinput40), 
        .A(n4070), .ZN(n4071) );
  NOR4_X1 U4756 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4103)
         );
  INV_X1 U4757 ( .A(D_REG_3__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U4758 ( .A1(n4076), .A2(keyinput17), .B1(n4680), .B2(keyinput21), 
        .ZN(n4075) );
  OAI221_X1 U4759 ( .B1(n4076), .B2(keyinput17), .C1(n4680), .C2(keyinput21), 
        .A(n4075), .ZN(n4081) );
  XNOR2_X1 U4760 ( .A(n4077), .B(keyinput13), .ZN(n4080) );
  XNOR2_X1 U4761 ( .A(n4078), .B(keyinput5), .ZN(n4079) );
  OR3_X1 U4762 ( .A1(n4081), .A2(n4080), .A3(n4079), .ZN(n4087) );
  INV_X1 U4763 ( .A(D_REG_18__SCAN_IN), .ZN(n4673) );
  INV_X1 U4764 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4765 ( .A1(n4673), .A2(keyinput33), .B1(keyinput53), .B2(n4083), 
        .ZN(n4082) );
  OAI221_X1 U4766 ( .B1(n4673), .B2(keyinput33), .C1(n4083), .C2(keyinput53), 
        .A(n4082), .ZN(n4086) );
  INV_X1 U4767 ( .A(D_REG_7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U4768 ( .A1(n4672), .A2(keyinput3), .B1(keyinput2), .B2(n4678), 
        .ZN(n4084) );
  OAI221_X1 U4769 ( .B1(n4672), .B2(keyinput3), .C1(n4678), .C2(keyinput2), 
        .A(n4084), .ZN(n4085) );
  NOR3_X1 U4770 ( .A1(n4087), .A2(n4086), .A3(n4085), .ZN(n4102) );
  AOI22_X1 U4771 ( .A1(n4089), .A2(keyinput23), .B1(keyinput22), .B2(n2267), 
        .ZN(n4088) );
  OAI221_X1 U4772 ( .B1(n4089), .B2(keyinput23), .C1(n2267), .C2(keyinput22), 
        .A(n4088), .ZN(n4100) );
  AOI22_X1 U4773 ( .A1(n4091), .A2(keyinput19), .B1(n4684), .B2(keyinput18), 
        .ZN(n4090) );
  OAI221_X1 U4774 ( .B1(n4091), .B2(keyinput19), .C1(n4684), .C2(keyinput18), 
        .A(n4090), .ZN(n4099) );
  INV_X1 U4775 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4776 ( .A1(n4094), .A2(keyinput14), .B1(n4093), .B2(keyinput11), 
        .ZN(n4092) );
  OAI221_X1 U4777 ( .B1(n4094), .B2(keyinput14), .C1(n4093), .C2(keyinput11), 
        .A(n4092), .ZN(n4098) );
  XNOR2_X1 U4778 ( .A(IR_REG_17__SCAN_IN), .B(keyinput30), .ZN(n4096) );
  XNOR2_X1 U4779 ( .A(DATAI_30_), .B(keyinput31), .ZN(n4095) );
  NAND2_X1 U4780 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  NOR4_X1 U4781 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4101)
         );
  NAND4_X1 U4782 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  AOI211_X1 U4783 ( .C1(n4108), .C2(n4107), .A(n4106), .B(n4105), .ZN(n4109)
         );
  XOR2_X1 U4784 ( .A(n4110), .B(n4109), .Z(U3553) );
  MUX2_X1 U4785 ( .A(DATAO_REG_2__SCAN_IN), .B(n2288), .S(U4043), .Z(U3552) );
  MUX2_X1 U4786 ( .A(DATAO_REG_1__SCAN_IN), .B(n2823), .S(U4043), .Z(U3551) );
  MUX2_X1 U4787 ( .A(DATAO_REG_0__SCAN_IN), .B(n2576), .S(U4043), .Z(U3550) );
  INV_X1 U4788 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4112) );
  MUX2_X1 U4789 ( .A(REG2_REG_19__SCAN_IN), .B(n4112), .S(n4362), .Z(n4124) );
  INV_X1 U4790 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4791 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4686), .B1(n4125), .B2(
        n4113), .ZN(n4648) );
  NOR2_X1 U4792 ( .A1(n4138), .A2(REG2_REG_17__SCAN_IN), .ZN(n4114) );
  AOI21_X1 U4793 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4138), .A(n4114), .ZN(n4638) );
  NOR2_X1 U4794 ( .A1(n4694), .A2(n4118), .ZN(n4119) );
  INV_X1 U4795 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4605) );
  XNOR2_X1 U4796 ( .A(n4694), .B(n4118), .ZN(n4604) );
  NOR2_X1 U4797 ( .A1(n4605), .A2(n4604), .ZN(n4603) );
  NOR2_X1 U4798 ( .A1(n4119), .A2(n4603), .ZN(n4614) );
  NAND2_X1 U4799 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4126), .ZN(n4120) );
  OAI21_X1 U4800 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4126), .A(n4120), .ZN(n4613) );
  NOR2_X1 U4801 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U4802 ( .A1(n4121), .A2(n4690), .ZN(n4122) );
  INV_X1 U4803 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U4804 ( .A1(n4638), .A2(n4636), .ZN(n4637) );
  AOI21_X1 U4805 ( .B1(n4125), .B2(REG2_REG_18__SCAN_IN), .A(n4647), .ZN(n4123) );
  XOR2_X1 U4806 ( .A(n4124), .B(n4123), .Z(n4150) );
  INV_X1 U4807 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4808 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4125), .B1(n4686), .B2(
        n4140), .ZN(n4654) );
  NOR2_X1 U4809 ( .A1(n4138), .A2(REG1_REG_17__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U4810 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4126), .ZN(n4133) );
  INV_X1 U4811 ( .A(n4126), .ZN(n4692) );
  AOI22_X1 U4812 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4126), .B1(n4692), .B2(
        n3510), .ZN(n4619) );
  INV_X1 U4813 ( .A(n4127), .ZN(n4129) );
  NAND2_X1 U4814 ( .A1(n4130), .A2(n4131), .ZN(n4132) );
  NAND2_X1 U4815 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4609), .ZN(n4608) );
  NAND2_X1 U4816 ( .A1(n4132), .A2(n4608), .ZN(n4618) );
  NAND2_X1 U4817 ( .A1(n4619), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U4818 ( .A1(n4133), .A2(n4617), .ZN(n4135) );
  NOR2_X1 U4819 ( .A1(n4134), .A2(n4135), .ZN(n4136) );
  XNOR2_X1 U4820 ( .A(n4135), .B(n4134), .ZN(n4626) );
  NOR2_X1 U4821 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4626), .ZN(n4625) );
  NOR2_X1 U4822 ( .A1(n4136), .A2(n4625), .ZN(n4642) );
  INV_X1 U4823 ( .A(n4138), .ZN(n4688) );
  AOI22_X1 U4824 ( .A1(n4138), .A2(n4137), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4688), .ZN(n4641) );
  MUX2_X1 U4825 ( .A(n4141), .B(REG1_REG_19__SCAN_IN), .S(n4362), .Z(n4142) );
  XNOR2_X1 U4826 ( .A(n4143), .B(n4142), .ZN(n4148) );
  NAND2_X1 U4827 ( .A1(n4650), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4144) );
  OAI211_X1 U4828 ( .C1(n4657), .C2(n4146), .A(n4145), .B(n4144), .ZN(n4147)
         );
  AOI21_X1 U4829 ( .B1(n4148), .B2(n4652), .A(n4147), .ZN(n4149) );
  OAI21_X1 U4830 ( .B1(n4150), .B2(n4646), .A(n4149), .ZN(U3259) );
  XNOR2_X1 U4831 ( .A(n4393), .B(n4151), .ZN(n4490) );
  INV_X1 U4832 ( .A(n4151), .ZN(n4154) );
  NOR2_X1 U4833 ( .A1(n4153), .A2(n4152), .ZN(n4395) );
  AOI21_X1 U4834 ( .B1(n4154), .B2(n4473), .A(n4395), .ZN(n4487) );
  NOR2_X1 U4835 ( .A1(n4487), .A2(n4670), .ZN(n4155) );
  AOI21_X1 U4836 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4670), .A(n4155), .ZN(n4156) );
  OAI21_X1 U4837 ( .B1(n4490), .B2(n4341), .A(n4156), .ZN(U3260) );
  OAI22_X1 U4838 ( .A1(n4158), .A2(n4341), .B1(n4157), .B2(n4658), .ZN(n4159)
         );
  AOI22_X1 U4839 ( .A1(n4161), .A2(n4379), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4670), .ZN(n4162) );
  NAND2_X1 U4840 ( .A1(n4165), .A2(n4374), .ZN(n4174) );
  INV_X1 U4841 ( .A(n4496), .ZN(n4172) );
  AOI22_X1 U4842 ( .A1(n4200), .A2(n4379), .B1(n4166), .B2(n4377), .ZN(n4169)
         );
  AOI22_X1 U4843 ( .A1(n4167), .A2(n4381), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4670), .ZN(n4168) );
  OAI211_X1 U4844 ( .C1(n4170), .C2(n4385), .A(n4169), .B(n4168), .ZN(n4171)
         );
  AOI21_X1 U4845 ( .B1(n4172), .B2(n4664), .A(n4171), .ZN(n4173) );
  OAI211_X1 U4846 ( .C1(n4670), .C2(n4175), .A(n4174), .B(n4173), .ZN(U3262)
         );
  NAND2_X1 U4847 ( .A1(n4177), .A2(n4176), .ZN(n4178) );
  AOI21_X1 U4848 ( .B1(n4179), .B2(n4178), .A(n4336), .ZN(n4406) );
  INV_X1 U4849 ( .A(n4406), .ZN(n4192) );
  XNOR2_X1 U4850 ( .A(n4180), .B(n4181), .ZN(n4407) );
  NAND2_X1 U4851 ( .A1(n4407), .A2(n4374), .ZN(n4191) );
  INV_X1 U4852 ( .A(n4205), .ZN(n4183) );
  OAI21_X1 U4853 ( .B1(n4183), .B2(n4186), .A(n2113), .ZN(n4500) );
  INV_X1 U4854 ( .A(n4500), .ZN(n4189) );
  AOI22_X1 U4855 ( .A1(n4184), .A2(n4381), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4670), .ZN(n4185) );
  OAI21_X1 U4856 ( .B1(n4186), .B2(n4385), .A(n4185), .ZN(n4188) );
  OAI22_X1 U4857 ( .A1(n4404), .A2(n4315), .B1(n4216), .B2(n4317), .ZN(n4187)
         );
  AOI211_X1 U4858 ( .C1(n4189), .C2(n4664), .A(n4188), .B(n4187), .ZN(n4190)
         );
  OAI211_X1 U4859 ( .C1(n4670), .C2(n4192), .A(n4191), .B(n4190), .ZN(U3263)
         );
  XOR2_X1 U4860 ( .A(n4196), .B(n2075), .Z(n4411) );
  INV_X1 U4861 ( .A(n4411), .ZN(n4210) );
  NAND2_X1 U4862 ( .A1(n4194), .A2(n4193), .ZN(n4195) );
  XOR2_X1 U4863 ( .A(n4196), .B(n4195), .Z(n4202) );
  OAI22_X1 U4864 ( .A1(n4198), .A2(n4478), .B1(n4197), .B2(n4331), .ZN(n4199)
         );
  AOI21_X1 U4865 ( .B1(n4200), .B2(n4475), .A(n4199), .ZN(n4201) );
  OAI21_X1 U4866 ( .B1(n4202), .B2(n4336), .A(n4201), .ZN(n4410) );
  NAND2_X1 U4867 ( .A1(n4223), .A2(n4203), .ZN(n4204) );
  NAND2_X1 U4868 ( .A1(n4205), .A2(n4204), .ZN(n4504) );
  AOI22_X1 U4869 ( .A1(n4670), .A2(REG2_REG_26__SCAN_IN), .B1(n4206), .B2(
        n4381), .ZN(n4207) );
  OAI21_X1 U4870 ( .B1(n4504), .B2(n4341), .A(n4207), .ZN(n4208) );
  AOI21_X1 U4871 ( .B1(n4410), .B2(n4365), .A(n4208), .ZN(n4209) );
  OAI21_X1 U4872 ( .B1(n4210), .B2(n4368), .A(n4209), .ZN(U3264) );
  XNOR2_X1 U4873 ( .A(n4211), .B(n4214), .ZN(n4415) );
  INV_X1 U4874 ( .A(n4415), .ZN(n4228) );
  NAND2_X1 U4875 ( .A1(n4213), .A2(n4212), .ZN(n4215) );
  XNOR2_X1 U4876 ( .A(n4215), .B(n4214), .ZN(n4220) );
  OAI22_X1 U4877 ( .A1(n4216), .A2(n4403), .B1(n4331), .B2(n4221), .ZN(n4217)
         );
  AOI21_X1 U4878 ( .B1(n4400), .B2(n4218), .A(n4217), .ZN(n4219) );
  OAI21_X1 U4879 ( .B1(n4220), .B2(n4336), .A(n4219), .ZN(n4414) );
  OR2_X1 U4880 ( .A1(n4236), .A2(n4221), .ZN(n4222) );
  NAND2_X1 U4881 ( .A1(n4223), .A2(n4222), .ZN(n4508) );
  AOI22_X1 U4882 ( .A1(n4670), .A2(REG2_REG_25__SCAN_IN), .B1(n4224), .B2(
        n4381), .ZN(n4225) );
  OAI21_X1 U4883 ( .B1(n4508), .B2(n4341), .A(n4225), .ZN(n4226) );
  AOI21_X1 U4884 ( .B1(n4414), .B2(n4365), .A(n4226), .ZN(n4227) );
  OAI21_X1 U4885 ( .B1(n4228), .B2(n4368), .A(n4227), .ZN(U3265) );
  NAND2_X1 U4886 ( .A1(n4230), .A2(n4229), .ZN(n4232) );
  XNOR2_X1 U4887 ( .A(n4232), .B(n4231), .ZN(n4233) );
  NAND2_X1 U4888 ( .A1(n4233), .A2(n4370), .ZN(n4420) );
  XNOR2_X1 U4889 ( .A(n4234), .B(n4235), .ZN(n4423) );
  NAND2_X1 U4890 ( .A1(n4423), .A2(n4374), .ZN(n4245) );
  INV_X1 U4891 ( .A(n4236), .ZN(n4237) );
  OAI21_X1 U4892 ( .B1(n4260), .B2(n4241), .A(n4237), .ZN(n4512) );
  INV_X1 U4893 ( .A(n4512), .ZN(n4243) );
  AOI22_X1 U4894 ( .A1(n4418), .A2(n4377), .B1(n4379), .B2(n4279), .ZN(n4240)
         );
  AOI22_X1 U4895 ( .A1(n4670), .A2(REG2_REG_24__SCAN_IN), .B1(n4238), .B2(
        n4381), .ZN(n4239) );
  OAI211_X1 U4896 ( .C1(n4241), .C2(n4385), .A(n4240), .B(n4239), .ZN(n4242)
         );
  AOI21_X1 U4897 ( .B1(n4243), .B2(n4664), .A(n4242), .ZN(n4244) );
  OAI211_X1 U4898 ( .C1(n4670), .C2(n4420), .A(n4245), .B(n4244), .ZN(U3266)
         );
  XNOR2_X1 U4899 ( .A(n4247), .B(n4246), .ZN(n4427) );
  INV_X1 U4900 ( .A(n4427), .ZN(n4267) );
  OR2_X1 U4901 ( .A1(n4287), .A2(n4248), .ZN(n4250) );
  OAI21_X1 U4902 ( .B1(n4278), .B2(n4277), .A(n4251), .ZN(n4253) );
  XNOR2_X1 U4903 ( .A(n4253), .B(n4252), .ZN(n4258) );
  OAI22_X1 U4904 ( .A1(n4255), .A2(n4403), .B1(n4331), .B2(n4254), .ZN(n4256)
         );
  AOI21_X1 U4905 ( .B1(n4400), .B2(n4436), .A(n4256), .ZN(n4257) );
  OAI21_X1 U4906 ( .B1(n4258), .B2(n4336), .A(n4257), .ZN(n4426) );
  AND2_X1 U4907 ( .A1(n4273), .A2(n4259), .ZN(n4261) );
  OR2_X1 U4908 ( .A1(n4261), .A2(n4260), .ZN(n4516) );
  INV_X1 U4909 ( .A(n4262), .ZN(n4263) );
  AOI22_X1 U4910 ( .A1(n4670), .A2(REG2_REG_23__SCAN_IN), .B1(n4263), .B2(
        n4381), .ZN(n4264) );
  OAI21_X1 U4911 ( .B1(n4516), .B2(n4341), .A(n4264), .ZN(n4265) );
  AOI21_X1 U4912 ( .B1(n4426), .B2(n4365), .A(n4265), .ZN(n4266) );
  OAI21_X1 U4913 ( .B1(n4267), .B2(n4368), .A(n4266), .ZN(U3267) );
  NAND2_X1 U4914 ( .A1(n4269), .A2(n4270), .ZN(n4271) );
  NAND2_X1 U4915 ( .A1(n4268), .A2(n4271), .ZN(n4430) );
  NAND2_X1 U4916 ( .A1(n4291), .A2(n2512), .ZN(n4272) );
  NAND2_X1 U4917 ( .A1(n4273), .A2(n4272), .ZN(n4521) );
  INV_X1 U4918 ( .A(n4521), .ZN(n4276) );
  OAI22_X1 U4919 ( .A1(n4365), .A2(n4089), .B1(n4274), .B2(n4658), .ZN(n4275)
         );
  AOI21_X1 U4920 ( .B1(n4276), .B2(n4664), .A(n4275), .ZN(n4286) );
  XNOR2_X1 U4921 ( .A(n4278), .B(n4277), .ZN(n4284) );
  NAND2_X1 U4922 ( .A1(n4279), .A2(n4475), .ZN(n4281) );
  NAND2_X1 U4923 ( .A1(n4445), .A2(n4400), .ZN(n4280) );
  OAI211_X1 U4924 ( .C1(n4331), .C2(n4282), .A(n4281), .B(n4280), .ZN(n4283)
         );
  AOI21_X1 U4925 ( .B1(n4284), .B2(n4370), .A(n4283), .ZN(n4431) );
  OR2_X1 U4926 ( .A1(n4431), .A2(n4670), .ZN(n4285) );
  OAI211_X1 U4927 ( .C1(n4430), .C2(n4368), .A(n4286), .B(n4285), .ZN(U3268)
         );
  XNOR2_X1 U4928 ( .A(n4287), .B(n4289), .ZN(n4288) );
  NAND2_X1 U4929 ( .A1(n4288), .A2(n4370), .ZN(n4438) );
  XNOR2_X1 U4930 ( .A(n4290), .B(n4289), .ZN(n4441) );
  NAND2_X1 U4931 ( .A1(n4441), .A2(n4374), .ZN(n4299) );
  OAI21_X1 U4932 ( .B1(n4309), .B2(n4295), .A(n4291), .ZN(n4525) );
  INV_X1 U4933 ( .A(n4525), .ZN(n4297) );
  AOI22_X1 U4934 ( .A1(n4379), .A2(n4333), .B1(n4377), .B2(n4436), .ZN(n4294)
         );
  AOI22_X1 U4935 ( .A1(n4670), .A2(REG2_REG_21__SCAN_IN), .B1(n4292), .B2(
        n4381), .ZN(n4293) );
  OAI211_X1 U4936 ( .C1(n4295), .C2(n4385), .A(n4294), .B(n4293), .ZN(n4296)
         );
  AOI21_X1 U4937 ( .B1(n4297), .B2(n4664), .A(n4296), .ZN(n4298) );
  OAI211_X1 U4938 ( .C1(n4670), .C2(n4438), .A(n4299), .B(n4298), .ZN(U3269)
         );
  NAND2_X1 U4939 ( .A1(n4301), .A2(n4300), .ZN(n4302) );
  XNOR2_X1 U4940 ( .A(n4302), .B(n4307), .ZN(n4303) );
  NAND2_X1 U4941 ( .A1(n4303), .A2(n4370), .ZN(n4447) );
  AOI21_X1 U4942 ( .B1(n4304), .B2(n4306), .A(n4305), .ZN(n4308) );
  XNOR2_X1 U4943 ( .A(n4308), .B(n4307), .ZN(n4450) );
  NAND2_X1 U4944 ( .A1(n4450), .A2(n4374), .ZN(n4322) );
  INV_X1 U4945 ( .A(n4338), .ZN(n4311) );
  INV_X1 U4946 ( .A(n4309), .ZN(n4310) );
  OAI21_X1 U4947 ( .B1(n4311), .B2(n4316), .A(n4310), .ZN(n4529) );
  INV_X1 U4948 ( .A(n4529), .ZN(n4320) );
  AOI22_X1 U4949 ( .A1(n4670), .A2(REG2_REG_20__SCAN_IN), .B1(n4312), .B2(
        n4381), .ZN(n4313) );
  OAI21_X1 U4950 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4319) );
  OAI22_X1 U4951 ( .A1(n4317), .A2(n4448), .B1(n4316), .B2(n4385), .ZN(n4318)
         );
  AOI211_X1 U4952 ( .C1(n4320), .C2(n4664), .A(n4319), .B(n4318), .ZN(n4321)
         );
  OAI211_X1 U4953 ( .C1(n4670), .C2(n4447), .A(n4322), .B(n4321), .ZN(U3270)
         );
  XNOR2_X1 U4954 ( .A(n4304), .B(n4323), .ZN(n4454) );
  INV_X1 U4955 ( .A(n4454), .ZN(n4346) );
  NAND2_X1 U4956 ( .A1(n4325), .A2(n4324), .ZN(n4355) );
  INV_X1 U4957 ( .A(n4326), .ZN(n4328) );
  OAI21_X1 U4958 ( .B1(n4355), .B2(n4328), .A(n4327), .ZN(n4330) );
  XNOR2_X1 U4959 ( .A(n4330), .B(n4329), .ZN(n4337) );
  NOR2_X1 U4960 ( .A1(n4339), .A2(n4331), .ZN(n4332) );
  AOI21_X1 U4961 ( .B1(n4333), .B2(n4475), .A(n4332), .ZN(n4335) );
  NAND2_X1 U4962 ( .A1(n4461), .A2(n4400), .ZN(n4334) );
  OAI211_X1 U4963 ( .C1(n4337), .C2(n4336), .A(n4335), .B(n4334), .ZN(n4453)
         );
  INV_X1 U4964 ( .A(n4350), .ZN(n4340) );
  OAI21_X1 U4965 ( .B1(n4340), .B2(n4339), .A(n4338), .ZN(n4533) );
  NOR2_X1 U4966 ( .A1(n4533), .A2(n4341), .ZN(n4344) );
  OAI22_X1 U4967 ( .A1(n4365), .A2(n4112), .B1(n4342), .B2(n4658), .ZN(n4343)
         );
  AOI211_X1 U4968 ( .C1(n4453), .C2(n4365), .A(n4344), .B(n4343), .ZN(n4345)
         );
  OAI21_X1 U4969 ( .B1(n4346), .B2(n4368), .A(n4345), .ZN(U3271) );
  INV_X1 U4970 ( .A(n4347), .ZN(n4348) );
  AOI21_X1 U4971 ( .B1(n4354), .B2(n4349), .A(n4348), .ZN(n4459) );
  INV_X1 U4972 ( .A(n4375), .ZN(n4353) );
  OAI211_X1 U4973 ( .C1(n4353), .C2(n4352), .A(n4351), .B(n4350), .ZN(n4456)
         );
  XNOR2_X1 U4974 ( .A(n4355), .B(n4354), .ZN(n4361) );
  AOI22_X1 U4975 ( .A1(n4357), .A2(n4475), .B1(n4473), .B2(n4356), .ZN(n4358)
         );
  OAI21_X1 U4976 ( .B1(n4359), .B2(n4478), .A(n4358), .ZN(n4360) );
  AOI21_X1 U4977 ( .B1(n4361), .B2(n4370), .A(n4360), .ZN(n4457) );
  OAI21_X1 U4978 ( .B1(n4362), .B2(n4456), .A(n4457), .ZN(n4366) );
  OAI22_X1 U4979 ( .A1(n4365), .A2(n4113), .B1(n4363), .B2(n4658), .ZN(n4364)
         );
  AOI21_X1 U4980 ( .B1(n4366), .B2(n4365), .A(n4364), .ZN(n4367) );
  OAI21_X1 U4981 ( .B1(n4459), .B2(n4368), .A(n4367), .ZN(U3272) );
  XNOR2_X1 U4982 ( .A(n4369), .B(n4373), .ZN(n4371) );
  NAND2_X1 U4983 ( .A1(n4371), .A2(n4370), .ZN(n4463) );
  XOR2_X1 U4984 ( .A(n4373), .B(n4372), .Z(n4466) );
  NAND2_X1 U4985 ( .A1(n4466), .A2(n4374), .ZN(n4390) );
  OAI21_X1 U4986 ( .B1(n4376), .B2(n4386), .A(n4375), .ZN(n4538) );
  INV_X1 U4987 ( .A(n4538), .ZN(n4388) );
  AOI22_X1 U4988 ( .A1(n4379), .A2(n4378), .B1(n4377), .B2(n4461), .ZN(n4384)
         );
  INV_X1 U4989 ( .A(n4380), .ZN(n4382) );
  AOI22_X1 U4990 ( .A1(n4670), .A2(REG2_REG_17__SCAN_IN), .B1(n4382), .B2(
        n4381), .ZN(n4383) );
  OAI211_X1 U4991 ( .C1(n4386), .C2(n4385), .A(n4384), .B(n4383), .ZN(n4387)
         );
  AOI21_X1 U4992 ( .B1(n4388), .B2(n4664), .A(n4387), .ZN(n4389) );
  OAI211_X1 U4993 ( .C1(n4670), .C2(n4463), .A(n4390), .B(n4389), .ZN(U3273)
         );
  NOR2_X1 U4994 ( .A1(n4487), .A2(n4724), .ZN(n4391) );
  AOI21_X1 U4995 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4724), .A(n4391), .ZN(n4392) );
  OAI21_X1 U4996 ( .B1(n4490), .B2(n4486), .A(n4392), .ZN(U3549) );
  AOI21_X1 U4997 ( .B1(n4396), .B2(n4394), .A(n4393), .ZN(n4555) );
  INV_X1 U4998 ( .A(n4555), .ZN(n4492) );
  INV_X1 U4999 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4397) );
  AOI21_X1 U5000 ( .B1(n4396), .B2(n4473), .A(n4395), .ZN(n4557) );
  MUX2_X1 U5001 ( .A(n4397), .B(n4557), .S(n4727), .Z(n4398) );
  OAI21_X1 U5002 ( .B1(n4492), .B2(n4486), .A(n4398), .ZN(U3548) );
  INV_X1 U5003 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U5004 ( .A1(n4401), .A2(n4400), .B1(n4399), .B2(n4473), .ZN(n4402)
         );
  OAI21_X1 U5005 ( .B1(n4404), .B2(n4403), .A(n4402), .ZN(n4405) );
  AOI211_X1 U5006 ( .C1(n4407), .C2(n4713), .A(n4406), .B(n4405), .ZN(n4497)
         );
  MUX2_X1 U5007 ( .A(n4408), .B(n4497), .S(n4727), .Z(n4409) );
  OAI21_X1 U5008 ( .B1(n4486), .B2(n4500), .A(n4409), .ZN(U3545) );
  INV_X1 U5009 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4412) );
  AOI21_X1 U5010 ( .B1(n4411), .B2(n4713), .A(n4410), .ZN(n4501) );
  MUX2_X1 U5011 ( .A(n4412), .B(n4501), .S(n4727), .Z(n4413) );
  OAI21_X1 U5012 ( .B1(n4486), .B2(n4504), .A(n4413), .ZN(U3544) );
  AOI21_X1 U5013 ( .B1(n4415), .B2(n4713), .A(n4414), .ZN(n4505) );
  MUX2_X1 U5014 ( .A(n4061), .B(n4505), .S(n4727), .Z(n4416) );
  OAI21_X1 U5015 ( .B1(n4486), .B2(n4508), .A(n4416), .ZN(U3543) );
  AOI22_X1 U5016 ( .A1(n4418), .A2(n4475), .B1(n4473), .B2(n4417), .ZN(n4419)
         );
  OAI211_X1 U5017 ( .C1(n4421), .C2(n4478), .A(n4420), .B(n4419), .ZN(n4422)
         );
  AOI21_X1 U5018 ( .B1(n4423), .B2(n4713), .A(n4422), .ZN(n4509) );
  MUX2_X1 U5019 ( .A(n4424), .B(n4509), .S(n4727), .Z(n4425) );
  OAI21_X1 U5020 ( .B1(n4486), .B2(n4512), .A(n4425), .ZN(U3542) );
  INV_X1 U5021 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4428) );
  AOI21_X1 U5022 ( .B1(n4427), .B2(n4713), .A(n4426), .ZN(n4513) );
  MUX2_X1 U5023 ( .A(n4428), .B(n4513), .S(n4727), .Z(n4429) );
  OAI21_X1 U5024 ( .B1(n4486), .B2(n4516), .A(n4429), .ZN(U3541) );
  INV_X1 U5025 ( .A(n4713), .ZN(n4458) );
  OR2_X1 U5026 ( .A1(n4430), .A2(n4458), .ZN(n4432) );
  NAND2_X1 U5027 ( .A1(n4432), .A2(n4431), .ZN(n4517) );
  MUX2_X1 U5028 ( .A(REG1_REG_22__SCAN_IN), .B(n4517), .S(n4727), .Z(n4433) );
  INV_X1 U5029 ( .A(n4433), .ZN(n4434) );
  OAI21_X1 U5030 ( .B1(n4486), .B2(n4521), .A(n4434), .ZN(U3540) );
  INV_X1 U5031 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U5032 ( .A1(n4436), .A2(n4475), .B1(n4473), .B2(n4435), .ZN(n4437)
         );
  OAI211_X1 U5033 ( .C1(n4439), .C2(n4478), .A(n4438), .B(n4437), .ZN(n4440)
         );
  AOI21_X1 U5034 ( .B1(n4441), .B2(n4713), .A(n4440), .ZN(n4522) );
  MUX2_X1 U5035 ( .A(n4442), .B(n4522), .S(n4727), .Z(n4443) );
  OAI21_X1 U5036 ( .B1(n4486), .B2(n4525), .A(n4443), .ZN(U3539) );
  INV_X1 U5037 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U5038 ( .A1(n4445), .A2(n4475), .B1(n4444), .B2(n4473), .ZN(n4446)
         );
  OAI211_X1 U5039 ( .C1(n4448), .C2(n4478), .A(n4447), .B(n4446), .ZN(n4449)
         );
  AOI21_X1 U5040 ( .B1(n4450), .B2(n4713), .A(n4449), .ZN(n4526) );
  MUX2_X1 U5041 ( .A(n4451), .B(n4526), .S(n4727), .Z(n4452) );
  OAI21_X1 U5042 ( .B1(n4486), .B2(n4529), .A(n4452), .ZN(U3538) );
  AOI21_X1 U5043 ( .B1(n4454), .B2(n4713), .A(n4453), .ZN(n4530) );
  MUX2_X1 U5044 ( .A(n4141), .B(n4530), .S(n4727), .Z(n4455) );
  OAI21_X1 U5045 ( .B1(n4486), .B2(n4533), .A(n4455), .ZN(U3537) );
  OAI211_X1 U5046 ( .C1(n4459), .C2(n4458), .A(n4457), .B(n4456), .ZN(n4534)
         );
  MUX2_X1 U5047 ( .A(REG1_REG_18__SCAN_IN), .B(n4534), .S(n4727), .Z(U3536) );
  AOI22_X1 U5048 ( .A1(n4461), .A2(n4475), .B1(n4473), .B2(n4460), .ZN(n4462)
         );
  OAI211_X1 U5049 ( .C1(n4464), .C2(n4478), .A(n4463), .B(n4462), .ZN(n4465)
         );
  AOI21_X1 U5050 ( .B1(n4466), .B2(n4713), .A(n4465), .ZN(n4535) );
  MUX2_X1 U5051 ( .A(n4137), .B(n4535), .S(n4727), .Z(n4467) );
  OAI21_X1 U5052 ( .B1(n4486), .B2(n4538), .A(n4467), .ZN(U3535) );
  INV_X1 U5053 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4471) );
  INV_X1 U5054 ( .A(n4468), .ZN(n4470) );
  AOI21_X1 U5055 ( .B1(n4470), .B2(n4713), .A(n4469), .ZN(n4539) );
  MUX2_X1 U5056 ( .A(n4471), .B(n4539), .S(n4727), .Z(n4472) );
  OAI21_X1 U5057 ( .B1(n4486), .B2(n4542), .A(n4472), .ZN(U3534) );
  INV_X1 U5058 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5059 ( .A1(n4476), .A2(n4475), .B1(n4474), .B2(n4473), .ZN(n4477)
         );
  OAI21_X1 U5060 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(n4482) );
  INV_X1 U5061 ( .A(n4480), .ZN(n4481) );
  AOI211_X1 U5062 ( .C1(n4711), .C2(n4483), .A(n4482), .B(n4481), .ZN(n4543)
         );
  MUX2_X1 U5063 ( .A(n4484), .B(n4543), .S(n4727), .Z(n4485) );
  OAI21_X1 U5064 ( .B1(n4486), .B2(n4547), .A(n4485), .ZN(U3532) );
  MUX2_X1 U5065 ( .A(n4488), .B(n4487), .S(n4719), .Z(n4489) );
  OAI21_X1 U5066 ( .B1(n4490), .B2(n4546), .A(n4489), .ZN(U3517) );
  MUX2_X1 U5067 ( .A(n2660), .B(n4557), .S(n4719), .Z(n4491) );
  OAI21_X1 U5068 ( .B1(n4492), .B2(n4546), .A(n4491), .ZN(U3516) );
  MUX2_X1 U5069 ( .A(n4494), .B(n4493), .S(n4719), .Z(n4495) );
  OAI21_X1 U5070 ( .B1(n4496), .B2(n4546), .A(n4495), .ZN(U3514) );
  INV_X1 U5071 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4498) );
  MUX2_X1 U5072 ( .A(n4498), .B(n4497), .S(n4719), .Z(n4499) );
  OAI21_X1 U5073 ( .B1(n4500), .B2(n4546), .A(n4499), .ZN(U3513) );
  INV_X1 U5074 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4502) );
  MUX2_X1 U5075 ( .A(n4502), .B(n4501), .S(n4719), .Z(n4503) );
  OAI21_X1 U5076 ( .B1(n4504), .B2(n4546), .A(n4503), .ZN(U3512) );
  MUX2_X1 U5077 ( .A(n4506), .B(n4505), .S(n4719), .Z(n4507) );
  OAI21_X1 U5078 ( .B1(n4508), .B2(n4520), .A(n4507), .ZN(U3511) );
  MUX2_X1 U5079 ( .A(n4510), .B(n4509), .S(n4719), .Z(n4511) );
  OAI21_X1 U5080 ( .B1(n4512), .B2(n4546), .A(n4511), .ZN(U3510) );
  MUX2_X1 U5081 ( .A(n4514), .B(n4513), .S(n4719), .Z(n4515) );
  OAI21_X1 U5082 ( .B1(n4516), .B2(n4546), .A(n4515), .ZN(U3509) );
  MUX2_X1 U5083 ( .A(REG0_REG_22__SCAN_IN), .B(n4517), .S(n4719), .Z(n4518) );
  INV_X1 U5084 ( .A(n4518), .ZN(n4519) );
  OAI21_X1 U5085 ( .B1(n4521), .B2(n4520), .A(n4519), .ZN(U3508) );
  MUX2_X1 U5086 ( .A(n4523), .B(n4522), .S(n4719), .Z(n4524) );
  OAI21_X1 U5087 ( .B1(n4525), .B2(n4546), .A(n4524), .ZN(U3507) );
  MUX2_X1 U5088 ( .A(n4527), .B(n4526), .S(n4719), .Z(n4528) );
  OAI21_X1 U5089 ( .B1(n4529), .B2(n4546), .A(n4528), .ZN(U3506) );
  MUX2_X1 U5090 ( .A(n4531), .B(n4530), .S(n4719), .Z(n4532) );
  OAI21_X1 U5091 ( .B1(n4533), .B2(n4546), .A(n4532), .ZN(U3505) );
  MUX2_X1 U5092 ( .A(REG0_REG_18__SCAN_IN), .B(n4534), .S(n4719), .Z(U3503) );
  MUX2_X1 U5093 ( .A(n4536), .B(n4535), .S(n4719), .Z(n4537) );
  OAI21_X1 U5094 ( .B1(n4538), .B2(n4546), .A(n4537), .ZN(U3501) );
  MUX2_X1 U5095 ( .A(n4540), .B(n4539), .S(n4719), .Z(n4541) );
  OAI21_X1 U5096 ( .B1(n4542), .B2(n4546), .A(n4541), .ZN(U3499) );
  MUX2_X1 U5097 ( .A(n4544), .B(n4543), .S(n4719), .Z(n4545) );
  OAI21_X1 U5098 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(U3495) );
  MUX2_X1 U5099 ( .A(n4548), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5100 ( .A(DATAI_27_), .B(n4549), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5101 ( .A(n4558), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5102 ( .A(DATAI_8_), .B(n4550), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5103 ( .A(n4551), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5104 ( .A(n4552), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5105 ( .A(DATAI_28_), .ZN(n4553) );
  AOI22_X1 U5106 ( .A1(STATE_REG_SCAN_IN), .A2(n4554), .B1(n4553), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5107 ( .A1(n4555), .A2(n4664), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4670), .ZN(n4556) );
  OAI21_X1 U5108 ( .B1(n4670), .B2(n4557), .A(n4556), .ZN(U3261) );
  INV_X1 U5109 ( .A(n4558), .ZN(n4567) );
  OAI211_X1 U5110 ( .C1(n4561), .C2(n4560), .A(n4652), .B(n4559), .ZN(n4566)
         );
  OAI211_X1 U5111 ( .C1(n4564), .C2(n4563), .A(n4631), .B(n4562), .ZN(n4565)
         );
  OAI211_X1 U5112 ( .C1(n4657), .C2(n4567), .A(n4566), .B(n4565), .ZN(n4568)
         );
  AOI211_X1 U5113 ( .C1(n4650), .C2(ADDR_REG_9__SCAN_IN), .A(n4569), .B(n4568), 
        .ZN(n4570) );
  INV_X1 U5114 ( .A(n4570), .ZN(U3249) );
  OAI211_X1 U5115 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4573), .A(n4652), .B(n4572), .ZN(n4577) );
  OAI211_X1 U5116 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4575), .A(n4631), .B(n4574), .ZN(n4576) );
  OAI211_X1 U5117 ( .C1(n4657), .C2(n2121), .A(n4577), .B(n4576), .ZN(n4578)
         );
  AOI211_X1 U5118 ( .C1(n4650), .C2(ADDR_REG_10__SCAN_IN), .A(n4579), .B(n4578), .ZN(n4580) );
  INV_X1 U5119 ( .A(n4580), .ZN(U3250) );
  OAI211_X1 U5120 ( .C1(n4583), .C2(n4582), .A(n4652), .B(n4581), .ZN(n4588)
         );
  OAI211_X1 U5121 ( .C1(n4586), .C2(n4585), .A(n4631), .B(n4584), .ZN(n4587)
         );
  OAI211_X1 U5122 ( .C1(n4657), .C2(n4696), .A(n4588), .B(n4587), .ZN(n4589)
         );
  AOI211_X1 U5123 ( .C1(n4650), .C2(ADDR_REG_11__SCAN_IN), .A(n4590), .B(n4589), .ZN(n4591) );
  INV_X1 U5124 ( .A(n4591), .ZN(U3251) );
  OAI211_X1 U5125 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4594), .A(n4631), .B(n4593), .ZN(n4596) );
  NAND2_X1 U5126 ( .A1(n4596), .A2(n4595), .ZN(n4597) );
  AOI21_X1 U5127 ( .B1(n4650), .B2(ADDR_REG_12__SCAN_IN), .A(n4597), .ZN(n4601) );
  OAI211_X1 U5128 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4599), .A(n4652), .B(n4598), .ZN(n4600) );
  OAI211_X1 U5129 ( .C1(n4657), .C2(n2123), .A(n4601), .B(n4600), .ZN(U3252)
         );
  INV_X1 U5130 ( .A(n4602), .ZN(n4607) );
  AOI211_X1 U5131 ( .C1(n4605), .C2(n4604), .A(n4603), .B(n4646), .ZN(n4606)
         );
  AOI211_X1 U5132 ( .C1(n4650), .C2(ADDR_REG_14__SCAN_IN), .A(n4607), .B(n4606), .ZN(n4611) );
  OAI211_X1 U5133 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4609), .A(n4652), .B(n4608), .ZN(n4610) );
  OAI211_X1 U5134 ( .C1(n4657), .C2(n4694), .A(n4611), .B(n4610), .ZN(U3254)
         );
  AOI211_X1 U5135 ( .C1(n4614), .C2(n4613), .A(n4612), .B(n4646), .ZN(n4615)
         );
  AOI211_X1 U5136 ( .C1(n4650), .C2(ADDR_REG_15__SCAN_IN), .A(n4616), .B(n4615), .ZN(n4621) );
  OAI211_X1 U5137 ( .C1(n4619), .C2(n4618), .A(n4652), .B(n4617), .ZN(n4620)
         );
  OAI211_X1 U5138 ( .C1(n4657), .C2(n4692), .A(n4621), .B(n4620), .ZN(U3255)
         );
  OAI21_X1 U5139 ( .B1(n4624), .B2(n4623), .A(n4622), .ZN(n4630) );
  AOI21_X1 U5140 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4626), .A(n4625), .ZN(n4628) );
  OAI22_X1 U5141 ( .A1(n4628), .A2(n4627), .B1(n4690), .B2(n4657), .ZN(n4629)
         );
  AOI21_X1 U5142 ( .B1(n4631), .B2(n4630), .A(n4629), .ZN(n4633) );
  OAI211_X1 U5143 ( .C1(n4635), .C2(n4634), .A(n4633), .B(n4632), .ZN(U3256)
         );
  AOI221_X1 U5144 ( .B1(n4638), .B2(n4637), .C1(n4636), .C2(n4637), .A(n4646), 
        .ZN(n4639) );
  AOI211_X1 U5145 ( .C1(n4650), .C2(ADDR_REG_17__SCAN_IN), .A(n4640), .B(n4639), .ZN(n4645) );
  OAI221_X1 U5146 ( .B1(n4643), .B2(n4642), .C1(n4643), .C2(n4641), .A(n4652), 
        .ZN(n4644) );
  OAI211_X1 U5147 ( .C1(n4657), .C2(n4688), .A(n4645), .B(n4644), .ZN(U3257)
         );
  OAI211_X1 U5148 ( .C1(n4654), .C2(n4653), .A(n4652), .B(n4651), .ZN(n4655)
         );
  OAI211_X1 U5149 ( .C1(n4657), .C2(n4686), .A(n4656), .B(n4655), .ZN(U3258)
         );
  OAI22_X1 U5150 ( .A1(n4365), .A2(n4660), .B1(n4659), .B2(n4658), .ZN(n4661)
         );
  INV_X1 U5151 ( .A(n4661), .ZN(n4668) );
  INV_X1 U5152 ( .A(n4662), .ZN(n4663) );
  AOI22_X1 U5153 ( .A1(n4666), .A2(n4665), .B1(n4664), .B2(n4663), .ZN(n4667)
         );
  OAI211_X1 U5154 ( .C1(n4670), .C2(n4669), .A(n4668), .B(n4667), .ZN(U3282)
         );
  AND2_X1 U5155 ( .A1(D_REG_31__SCAN_IN), .A2(n4682), .ZN(U3291) );
  NOR2_X1 U5156 ( .A1(n4681), .A2(n4671), .ZN(U3292) );
  NOR2_X1 U5157 ( .A1(n4681), .A2(n4672), .ZN(U3293) );
  AND2_X1 U5158 ( .A1(D_REG_28__SCAN_IN), .A2(n4682), .ZN(U3294) );
  AND2_X1 U5159 ( .A1(D_REG_27__SCAN_IN), .A2(n4682), .ZN(U3295) );
  AND2_X1 U5160 ( .A1(D_REG_26__SCAN_IN), .A2(n4682), .ZN(U3296) );
  AND2_X1 U5161 ( .A1(n4682), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  AND2_X1 U5162 ( .A1(D_REG_24__SCAN_IN), .A2(n4682), .ZN(U3298) );
  AND2_X1 U5163 ( .A1(n4682), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  AND2_X1 U5164 ( .A1(D_REG_22__SCAN_IN), .A2(n4682), .ZN(U3300) );
  AND2_X1 U5165 ( .A1(D_REG_21__SCAN_IN), .A2(n4682), .ZN(U3301) );
  AND2_X1 U5166 ( .A1(D_REG_20__SCAN_IN), .A2(n4682), .ZN(U3302) );
  AND2_X1 U5167 ( .A1(D_REG_19__SCAN_IN), .A2(n4682), .ZN(U3303) );
  NOR2_X1 U5168 ( .A1(n4681), .A2(n4673), .ZN(U3304) );
  NOR2_X1 U5169 ( .A1(n4681), .A2(n4674), .ZN(U3305) );
  AND2_X1 U5170 ( .A1(D_REG_16__SCAN_IN), .A2(n4682), .ZN(U3306) );
  AND2_X1 U5171 ( .A1(D_REG_15__SCAN_IN), .A2(n4682), .ZN(U3307) );
  NOR2_X1 U5172 ( .A1(n4681), .A2(n4675), .ZN(U3308) );
  AND2_X1 U5173 ( .A1(D_REG_13__SCAN_IN), .A2(n4682), .ZN(U3309) );
  AND2_X1 U5174 ( .A1(D_REG_12__SCAN_IN), .A2(n4682), .ZN(U3310) );
  AND2_X1 U5175 ( .A1(D_REG_11__SCAN_IN), .A2(n4682), .ZN(U3311) );
  AND2_X1 U5176 ( .A1(D_REG_10__SCAN_IN), .A2(n4682), .ZN(U3312) );
  NOR2_X1 U5177 ( .A1(n4681), .A2(n4676), .ZN(U3313) );
  NOR2_X1 U5178 ( .A1(n4681), .A2(n4677), .ZN(U3314) );
  NOR2_X1 U5179 ( .A1(n4681), .A2(n4678), .ZN(U3315) );
  AND2_X1 U5180 ( .A1(D_REG_6__SCAN_IN), .A2(n4682), .ZN(U3316) );
  NOR2_X1 U5181 ( .A1(n4681), .A2(n4679), .ZN(U3317) );
  AND2_X1 U5182 ( .A1(D_REG_4__SCAN_IN), .A2(n4682), .ZN(U3318) );
  NOR2_X1 U5183 ( .A1(n4681), .A2(n4680), .ZN(U3319) );
  AND2_X1 U5184 ( .A1(D_REG_2__SCAN_IN), .A2(n4682), .ZN(U3320) );
  AOI21_X1 U5185 ( .B1(U3149), .B2(n4684), .A(n4683), .ZN(U3329) );
  AOI22_X1 U5186 ( .A1(STATE_REG_SCAN_IN), .A2(n4686), .B1(n4685), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5187 ( .A1(STATE_REG_SCAN_IN), .A2(n4688), .B1(n4687), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5188 ( .A1(STATE_REG_SCAN_IN), .A2(n4690), .B1(n4689), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5189 ( .A(DATAI_15_), .ZN(n4691) );
  AOI22_X1 U5190 ( .A1(STATE_REG_SCAN_IN), .A2(n4692), .B1(n4691), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5191 ( .A1(STATE_REG_SCAN_IN), .A2(n4694), .B1(n4693), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5192 ( .A(DATAI_12_), .ZN(n4695) );
  AOI22_X1 U5193 ( .A1(STATE_REG_SCAN_IN), .A2(n2123), .B1(n4695), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5194 ( .A1(STATE_REG_SCAN_IN), .A2(n4696), .B1(n2399), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5195 ( .A(DATAI_10_), .ZN(n4697) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n2121), .B1(n4697), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5197 ( .A(DATAI_0_), .ZN(n4698) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4699), .B1(n4698), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5199 ( .A1(n4719), .A2(n4700), .B1(n2267), .B2(n4718), .ZN(U3467)
         );
  INV_X1 U5200 ( .A(n4701), .ZN(n4705) );
  INV_X1 U5201 ( .A(n4702), .ZN(n4704) );
  AOI211_X1 U5202 ( .C1(n4705), .C2(n4711), .A(n4704), .B(n4703), .ZN(n4721)
         );
  AOI22_X1 U5203 ( .A1(n4719), .A2(n4721), .B1(n2304), .B2(n4718), .ZN(U3475)
         );
  NOR3_X1 U5204 ( .A1(n4708), .A2(n4707), .A3(n4706), .ZN(n4710) );
  AOI211_X1 U5205 ( .C1(n4712), .C2(n4711), .A(n4710), .B(n4709), .ZN(n4723)
         );
  AOI22_X1 U5206 ( .A1(n4719), .A2(n4723), .B1(n2332), .B2(n4718), .ZN(U3479)
         );
  AND3_X1 U5207 ( .A1(n3121), .A2(n4714), .A3(n4713), .ZN(n4715) );
  NOR3_X1 U5208 ( .A1(n4717), .A2(n4716), .A3(n4715), .ZN(n4726) );
  AOI22_X1 U5209 ( .A1(n4719), .A2(n4726), .B1(n2341), .B2(n4718), .ZN(U3481)
         );
  AOI22_X1 U5210 ( .A1(n4727), .A2(n4721), .B1(n4720), .B2(n4724), .ZN(U3522)
         );
  AOI22_X1 U5211 ( .A1(n4727), .A2(n4723), .B1(n4722), .B2(n4724), .ZN(U3524)
         );
  INV_X1 U5212 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5213 ( .A1(n4727), .A2(n4726), .B1(n4725), .B2(n4724), .ZN(U3525)
         );
  CLKBUF_X3 U2297 ( .A(n2290), .Z(n3827) );
  CLKBUF_X3 U2298 ( .A(n2271), .Z(n3831) );
  CLKBUF_X1 U2308 ( .A(n2278), .Z(n2342) );
  CLKBUF_X1 U2704 ( .A(n2723), .Z(n2055) );
endmodule

