
module b21_C_2inp_gates_syn ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN,
    ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966;
  wire n13995, n11811, n12487, n17409, n16014, n17227, n9355, n10698, n12524,
    n13606, n14977, n16310, n13384, n17505, n12581, n16320, n15080, n15024,
    n16274, n11216, n12439, n15869, n15930, n15972, n13546, n15286, n11249,
    n13164, n11063, n8992, n12788, n13972, n15016, n13974, n9827, n15198,
    n17041, n17095, n17399, n16516, n16078, n8987, n10828, n11802, n11200,
    n11196, n12395, n11973, n13105, n12706, n13980, n14012, n14345, n13558,
    n14266, n9171, n14567, n9609, n14529, n9272, n15047, n13984, n15035,
    n14006, n11032, n13644, n14017, n15069, n14049, n13690, n11785, n14789,
    n13757, n13020, n13825, n12299, n14933, n9556, n14936, n14060, n15145,
    n14071, n9643, n9595, n12660, n15841, n15155, n14363, n14091, n14114,
    n11467, n15365, n16955, n15209, n9483, n9491, n15396, n16487, n17067,
    n17419, n15954, n15411, n12098, n16625, n17387, n12430, n11864, n16046,
    n8995, n16283, n12624, n11923, n11391, n8990, n16463, n9959, n12248,
    n12102, n9957, n9484, n8988, n10101, n16251, n10089, n13191, n10234,
    n11181, n11285, n10012, n12791, n11243, n12422, n10815, n11204, n10207,
    n10361, n11229, n14227, n10812, n11198, n10467, n11543, n9844, n9845,
    n11211, n9978, n11162, n11175, n11176, n11169, n11208, n10018, n9977,
    n9602, n11164, n11165, n11163, n10016, n11166, n11144, n9970, n10814,
    n14500, n17185, n13329, n13541, n12268, n11289, n14663, n10481, n8989,
    n8991, n12429, n14573, n14552, n14621, n11295, n8993, n8994, n11299,
    n8996, n11068, n12725, n9307, n9800, n9801, n9743, n9522, n13064,
    n13075, n11069, n9933, n9618, n9619, n9426, n9893, n9834, n9836, n9284,
    n9285, n9809, n9557, n13833, n9289, n9985, n9984, n10339, n9788,
    n13098, n9903, n9885, n9886, n14559, n13169, n12647, n9336, n10271,
    n10242, n9941, n9942, n16943, n17033, n13748, n9215, n9275, n9320,
    n10562, n10514, n9439, n9440, n11816, n9437, n9449, n9450, n9222,
    n9730, n11307, n9872, n9392, n12241, n12242, n9855, n9589, n9865,
    n9591, n14881, n9607, n9342, n9343, n9344, n10380, n10345, n9776,
    n9777, n9778, n9779, n14323, n11851, n16074, n12294, n12835, n9402,
    n9403, n9396, n9397, n9503, n9703, n9724, n9231, n9369, n11106, n9471,
    n9408, n13044, n13047, n9328, n9704, n9467, n9539, n12806, n9528,
    n9529, n9532, n9533, n9534, n9535, n9742, n9525, n9526, n9523, n9416,
    n9465, n9209, n9210, n9211, n9917, n9939, n9555, n9948, n9310, n9580,
    n9548, n9305, n9876, n9878, n13134, n10711, n9261, n9750, n9751,
    n10319, n9306, n9278, n13538, n11094, n9817, n11088, n9958, n9752,
    n9286, n9288, n9579, n9219, n9549, n9926, n9217, n9569, n13204, n9441,
    n11303, n11367, n13126, n12815, n9540, n9541, n9542, n9612, n9899,
    n12238, n9615, n9424, n9425, n9617, n12680, n14609, n9390, n9860,
    n9862, n13041, n13021, n9476, n14856, n12959, n12222, n13143, n12736,
    n9361, n9672, n9915, n9916, n10408, n10232, n9474, n9640, n9823, n9821,
    n9242, n12445, n10822, n10041, n9746, n12522, n9379, n9380, n9830,
    n12512, n12460, n13317, n9710, n9337, n9208, n9708, n9709, n9196,
    n9246, n9253, n9259, n9260, n9257, n13260, n13665, n9759, n9796,
    n11000, n10999, n9763, n10498, n9755, n9756, n10254, n13280, n9919,
    n9311, n9312, n11050, n9216, n9293, n9570, n9574, n9294, n9295, n9273,
    n9274, n9568, n9987, n10214, n10441, n10094, n9434, n11461, n11389,
    n9667, n9668, n13180, n9502, n9496, n15780, n9695, n9696, n9420, n9421,
    n13010, n12997, n12895, n15891, n9384, n9482, n16042, n14587, n12824,
    n16023, n14616, n14633, n12674, n9585, n9869, n9882, n15961, n9520,
    n9519, n9737, n9738, n9356, n9358, n9357, n9359, n10648, n10651,
    n11182, n10647, n9908, n9907, n16124, n9234, n9459, n9914, n10382,
    n9662, n10295, n9202, n9458, n9381, n12610, n12511, n9493, n10306,
    n9494, n14102, n14113, n12597, n16626, n9313, n12586, n9268, n9249,
    n9266, n9265, n9221, n9567, n17150, n17191, n13945, n9339, n9340,
    n13539, n13258, n13259, n9812, n17487, n11130, n17225, n9323, n9319,
    n10780, n10816, n9207, n17272, n9597, n9770, n14252, n9455, n9456,
    n11824, n9784, n14327, n15091, n11551, n9781, n9782, n11943, n9401,
    n15604, n15719, n12085, n13082, n15025, n11454, n15023, n16357, n16309,
    n12295, n12289, n12290, n16245, n11870, n11231, n10803, n10763, n10716,
    n9194, n12346, n10629, n11194, n11195, n16922, n16794, n15421, n16426,
    n15686, n16241, n17638, n17630, n9497, n9410, n9411, n10865, n9728,
    n10888, n12974, n9332, n9472, n9735, n9736, n9509, n9726, n9469, n9723,
    n9365, n9362, n9363, n12726, n13049, n9229, n9230, n9707, n13161,
    n9366, n9368, n9530, n9521, n9511, n9937, n13068, n9406, n9741, n11073,
    n11072, n9324, n9718, n9330, n9326, n9936, n9981, n9982, n9983, n9536,
    n9537, n9538, n12811, n9531, n9524, n9897, n9898, n9896, n9417, n10719,
    n11167, n9665, n11158, n11159, n10015, n9241, n9489, n9633, n9634,
    n9832, n9338, n9946, n9944, n9945, n9513, n11114, n9200, n9201, n9551,
    n11090, n9309, n13678, n9929, n9931, n9575, n13895, n9299, n10518,
    n9447, n9443, n9446, n9451, n9452, n9623, n9732, n9423, n9393, n9874,
    n15918, n9383, n9729, n9856, n9852, n9853, n14605, n13175, n9682,
    n9588, n9887, n9867, n9690, n12661, n9605, n9606, n9394, n9594, n9881,
    n9883, n9889, n9891, n15893, n15896, n10717, n10694, n11203, n10434,
    n9912, n10328, n10241, n9842, n12515, n10702, n9247, n13505, n13569,
    n10664, n10635, n9762, n10622, n10595, n10569, n9757, n9758, n10447,
    n17008, n9271, n9805, n17074, n9276, n9279, n13207, n13287, n9814,
    n13253, n13588, n9283, n9218, n9811, n13631, n9947, n13244, n9220,
    n9213, n9212, n9753, n9754, n9819, n17096, n16489, n17373, n10817,
    n10543, n9674, n9675, n9321, n10522, n10386, n9775, n9772, n9767,
    n9768, n9445, n9444, n9442, n15392, n14411, n11270, n9785, n14289,
    n9790, n11631, n9544, n9545, n12820, n15792, n11855, n9176, n9610,
    n14713, n9678, n11733, n14792, n11666, n15969, n16025, n9599, n9600,
    n12650, n9614, n9386, n9863, n9864, n14660, n14681, n9900, n9683,
    n14790, n14735, n9680, n9679, n14749, n14871, n9685, n9686, n9688,
    n9608, n14992, n9492, n12245, n12406, n12652, n15956, n16296, n16020,
    n16055, n11212, n11205, n10657, n10610, n10582, n11199, n10460, n11592,
    n10270, n11472, n9560, n11382, n10147, n9480, n16628, n9637, n9645,
    n16501, n16583, n9174, n16608, n17432, n9656, n13494, n13495, n9345,
    n9205, n9348, n13806, n12005, n13898, n10921, n12026, n9954, n16655,
    n9251, n10334, n9256, n13531, n9581, n9583, n13713, n9233, n13926,
    n10312, n17362, n17081, n17134, n9748, n9298, n12571, n13953, n13986,
    n13701, n9799, n9807, n14107, n9290, n16929, n16983, n10191, n17224,
    n9699, n11143, n10824, n10818, n10819, n10811, n17334, n14586, n14237,
    n14269, n15348, n14320, n9429, n14375, n14378, n15412, n9487, n15188,
    n14470, n15134, n15429, n12792, n9400, n14751, n13011, n14828, n14804,
    n14364, n14937, n14965, n14993, n14964, n15847, n9373, n9374, n12908,
    n15848, n15437, n15326, n9404, n11247, n9179, n9177, n9182, n15748,
    n9187, n9188, n9693, n9694, n15034, n9880, n14296, n9372, n11504,
    n9385, n12237, n15926, n9473, n16108, n12400, n14594, n15065, n14689,
    n9592, n16261, n9677, n9517, n11172, n9354, n10760, n9170, n9464,
    n15319, n9206, n11190, n11188, n17245, n9913, n17265, n17284, n10210,
    n10203, n17305, n15489, n16226, n16569, n13344, n9378, n9824, n9826,
    n13392, n13393, n13419, n16617, n9479, n16575, n17585, n17561, n13395,
    n13838, n13871, n13935, n16506, n16592, n16505, n16559, n16477, n16558,
    n16627, n17342, n16913, n16811, n16868, n9264, n17209, n12582, n17130,
    n17553, n17555, n14175, n17501, n13291, n17514, n17358, n17352, n11132,
    n17351, n9991, n12569, n11145, n10782, n9793, n9795, n9454, n14329,
    n14843, n14466, n15457, n13198, n13120, n9486, n16419, n16416, n16413,
    n14703, n14774, n14859, n14533, n14908, n14907, n15903, n15929, n15585,
    n9190, n16011, n16003, n16109, n16119, n16393, n16395, n12419, n12700,
    n16349, n16363, n16239, n16234, n16233, n15276, n15275, n15309, n12334,
    n16128, n16225, n15502, n17646, n17634, n17626, n9563, n9508, n8997,
    n8998, n11077, n11093, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n11008, n9010, n9173, n9011, n13837,
    n13897, n9012, n9577, n12902, n9765, n9013, n17087, n9014, n9015,
    n9016, n12800, n9017, n9018, n9019, n9020, n13813, n9021, n15958,
    n9022, n9364, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n17582, n9036, n10428, n9572, n9037,
    n9038, n10523, n9039, n9040, n14905, n14701, n13559, n13774, n9041,
    n9042, n9043, n9044, n13583, n9045, n9046, n13933, n9047, n13964,
    n9749, n9048, n9049, n9050, n9051, n9052, n13680, n9053, n9054, n9055,
    n9056, n9057, n13107, n9058, n13679, n9059, n9510, n14799, n9060,
    n9061, n9062, n12737, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n13622, n9076, n9077, n13572,
    n9078, n13892, n9079, n9080, n9081, n9082, n9083, n11230, n9084, n9085,
    n9697, n13920, n9086, n9760, n9761, n9087, n9088, n9407, n9089, n9901,
    n9902, n11228, n9350, n9090, n13714, n15277, n9091, n12759, n9092,
    n9093, n9094, n9095, n17588, n9918, n9797, n9798, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n14464, n9103, n9104, n9105, n9414, n16244,
    n16087, n9106, n13608, n9107, n9108, n9109, n10091, n9262, n14922,
    n9687, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9192, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9462, n9235, n9133, n10004, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9843, n9145, n9146, n9147, n9148, n9149, n9500, n11082, n9689, n17028,
    n9684, n9150, n13932, n17009, n13432, n13835, n9512, n9151, n9764,
    n9698, n9152, n13142, n9153, n9322, n9154, n9155, n9156, n9157, n9158,
    n9159, n15925, n16076, n10825, n9160, n13192, n9161, n16088, n9162,
    n17098, n13537, n16924, n9657, n9291, n10159, n10267, n9292, n9573,
    n13629, n13237, n9460, n9237, n12967, n9163, n12984, n9164, n9658,
    n9490, n10663, n9552, n11155, n9165, n12345, n9527, n9341, n9226,
    n12703, n14213, n9616, n10013, n13168, n9166, n13132, n9282, n13179,
    n9167, n13190, n9168, n9169, n13630, n14208, n13106, n13121, n12532,
    n11123, n13266, n9172, n9238, n9377, n13073, n10034, n12438, n9175,
    n9601, n15374, n11281, n14503, n17039, n13615, n11634, n14654, n9676,
    n9613, n9183, n15541, n15543, n9178, n9180, n15531, n9181, n15794,
    n9184, n9185, n9186, n15582, n15607, n15749, n9189, n9191, n9193,
    n11251, n9195, n9197, n9198, n9199, n9203, n9204, n10587, n10618,
    n10652, n12322, n11119, n13832, n13230, n13231, n13827, n9214, n9506,
    n13103, n9223, n9224, n9225, n9227, n9228, n12609, n9840, n13405,
    n9232, n9240, n9236, n9239, n9375, n9243, n9244, n9254, n9250, n9245,
    n9252, n12127, n9248, n16693, n16695, n16746, n9255, n16744, n9258,
    n10047, n16812, n9263, n12117, n9267, n12185, n16869, n9269, n16848,
    n9270, n17026, n13725, n9578, n13224, n9280, n17114, n17105, n9277,
    n13254, n9281, n9810, n9287, n9296, n13891, n13293, n13961, n9297,
    n17161, n10061, n17363, n17189, n16574, n9304, n10105, n9302, n9300,
    n9301, n17147, n17091, n9303, n16964, n9501, n13800, n13803, n9308,
    n10745, n11085, n9713, n9314, n9315, n9316, n9468, n9317, n9318,
    n10781, n9727, n9325, n9327, n9329, n11031, n9331, n9335, n9333, n9334,
    n10955, n9516, n9376, n10661, n9920, n10747, n9346, n9347, n9349,
    n9351, n9352, n9353, n9360, n11286, n12761, n12769, n9367, n12789,
    n9370, n9371, n13446, n17238, n9828, n9382, n16299, n15927, n15867,
    n12678, n9387, n9388, n14711, n9389, n9391, n9593, n9395, n12929,
    n12916, n9398, n9399, n9624, n9405, n9409, n9412, n12894, n9413,
    n11232, n9625, n9415, n16021, n9418, n14724, n9419, n9422, n12646,
    n14772, n9427, n14584, n9428, n12645, n12644, n11569, n14447, n12307,
    n15352, n9430, n15375, n15427, n9431, n9432, n14531, n9433, n11276,
    n9435, n9436, n9438, n9789, n9783, n9448, n14306, n9453, n9769, n9457,
    n14239, n11929, n15333, n12073, n11201, n10202, n9649, n9586, n9596,
    n15177, n9647, n16526, n12648, n11304, n10536, n9952, n12427, n10429,
    n12474, n9461, n13379, n9669, n13634, n9611, n9546, n9922, n14361,
    n9463, n16070, n9604, n10036, n9488, n10081, n10511, n10075, n9648,
    n9847, n9846, n11628, n11466, n9466, n12847, n12830, n14254, n9794,
    n11944, n11134, n9706, n9498, n12826, n9990, n9992, n14139, n9470,
    n9620, n9858, n15031, n15894, n11101, n11110, n13104, n9543, n16006,
    n10237, n9475, n12829, n9477, n9622, n12856, n9478, n12994, n9631,
    n11271, n9651, n9820, n10354, n12538, n9773, n14757, n12684, n9485,
    n9481, n12694, n12236, n16041, n14642, n12664, n14834, n14731, n12882,
    n9505, n12831, n11259, n9739, n15394, n9504, n11122, n14141, n9905,
    n9553, n10083, n17298, n11430, n9660, n15875, n14975, n9871, n11401,
    n9495, n10546, n12839, n9774, n9787, n9791, n9661, n10726, n13110,
    n13605, n9499, n13599, n12110, n13845, n13593, n11272, n10010, n17048,
    n9923, n9895, n10920, n10836, n9515, n9507, n9771, n9636, n9747,
    n10321, n11115, n9514, n11768, n10539, n9518, n9547, n9550, n9554,
    n13610, n13607, n10508, n10175, n9559, n9558, n9562, n10233, n9561,
    n9564, n9565, n9566, n13234, n9571, n9576, n16961, n9582, n9584,
    n14868, n9587, n14917, n9590, n9879, n9598, n14568, n11191, n11636,
    n9603, n14560, n9621, n9626, n9627, n9628, n9629, n9630, n16430,
    n16474, n9632, n9635, n9822, n9638, n12494, n9639, n9641, n9642,
    n16503, n9644, n12534, n13460, n9646, n9650, n9652, n13359, n9653,
    n9654, n9655, n9910, n17333, n10056, n9911, n9659, n10324, n9663,
    n9664, n12771, n12776, n9666, n9670, n9671, n9673, n15101, n12401,
    n9681, n14733, n14920, n9691, n9692, n12695, n14596, n9988, n9921,
    n9956, n9700, n9701, n9702, n9705, n9711, n10905, n9712, n9714, n11049,
    n9715, n9716, n9719, n9717, n10837, n9720, n9721, n9722, n9725, n16071,
    n9733, n9731, n9734, n13002, n13015, n9740, n11214, n11227, n9744,
    n13202, n10080, n12961, n11581, n13951, n14135, n9745, n10100, n10125,
    n10732, n17142, n13908, n11921, n11241, n9766, n12205, n14519, n9780,
    n9786, n11522, n9792, n9802, n17057, n9803, n9804, n13773, n9806,
    n13799, n9808, n9815, n9813, n13554, n9816, n9818, n10005, n12643,
    n9825, n12629, n16584, n9829, n9831, n16445, n9833, n9835, n13294,
    n9837, n9838, n9839, n9841, n10465, n9848, n16620, n9849, n9850, n9851,
    n9854, n9857, n14661, n9859, n9861, n9866, n14884, n9868, n9870, n9873,
    n14963, n9875, n9877, n14959, n14989, n9884, n9888, n9890, n15845,
    n9892, n9894, n14604, n9904, n17291, n9906, n10563, n9909, n10140,
    n10143, n10402, n10678, n11142, n17082, n9924, n9925, n9927, n9930,
    n13702, n9928, n13726, n9932, n9938, n9934, n9935, n9940, n17116,
    n9943, n9949, n13654, n9950, n9951, n9953, n13017, n13787, n10017,
    n14737, n11924, n12247, n13102, n14220, n17197, n11988, n10062, n10245,
    n9996, n13330, n9993, n10060, n10049, n10258, n11263, n14187, n9955,
    n9989, n12584, n11126, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n10177, n10357, n10163, n9979, n13174, n12774, n11168,
    n10581, n13226, n10521, n11913, n10720, n10650, n11336, n10000, n13279,
    n13219, n11138, n10517, n14562, n11903, n11233, n11747, n16077, n11213,
    n10675, n10433, n11125, n13255, n16490, n16605, n13274, n10683, n10552,
    n13805, n17504, n17493, n10542, n11711, n11713, n11825, n12287, n16084,
    n14935, n15175, n16045, n12288, n11215, n10605, n11129, n16624, n13557,
    n17173, n13801, n13510, n13639, n17212, n13290, n17239, n15438, n15378,
    n14608, n13109, n11658, n16116, n12693, n11185, n10660, n10355, n12588,
    n16554, n13491, n16472, n12152, n17068, n13948, n13949, n12329, n15419,
    n15441, n15447, n15442, n15653, n15996, n14918, n12291, n16122, n11187,
    n16622, n16631, n17595, n17564, n16872, n17206, n17186, n17218, n14184,
    n17340, n17347, n15402, n15414, n16404, n14509, n15881, n15816, n16040,
    n16105, n16104, n15317, n17647, n17643, n17594, n17350, n16425, n17650,
    n17642, n9969, n9972, n9971, n9976, n9974, n9973, n9975, n10090,
    n11133, n10212, n10438, n9980, n9986, n10440, n9994, n14196, n9995,
    n10777, n10003, n9997, n10068, n9999, n10065, n9998, n10001, n10002,
    n10826, n11147, n10006, n10009, n10007, n10008, n10011, n14214, n10021,
    n10014, n10054, n10019, n11966, n10020, n16568, n10026, n10023, n10022,
    n10024, n10025, n10027, n10042, n10085, n10028, n10031, n10029, n10030,
    n10032, n10033, n10035, n10079, n10038, n10037, n10039, n10073, n10050,
    n17341, n10040, n10063, n10046, n10044, n10043, n10045, n11976, n12194,
    n10048, n10053, n10051, n10052, n10058, n10055, n10076, n10057, n11972,
    n10059, n11095, n10064, n10396, n10067, n10066, n10072, n10070, n16456,
    n10069, n10071, n16541, n10074, n10078, n10077, n10084, n10082, n10087,
    n10086, n10123, n10088, n10122, n10098, n10092, n10093, n10096, n10095,
    n10097, n10099, n10104, n10102, n10103, n17141, n10106, n10108, n10107,
    n10114, n10112, n16534, n10109, n10153, n17125, n10110, n10111, n10113,
    n16517, n10866, n10115, n10118, n10116, n17327, n10117, n10126, n10120,
    n10119, n10141, n10121, n10139, n10124, n17326, n17133, n10127, n17102,
    n10129, n10128, n10133, n10131, n10130, n10132, n13214, n10768, n10134,
    n10138, n10135, n10168, n10136, n17320, n10137, n10148, n10142, n10145,
    n10144, n10160, n10146, n10158, n17319, n11097, n10149, n11096, n10151,
    n10150, n10157, n10684, n10152, n10192, n16618, n17069, n10155, n10154,
    n10156, n10162, n10161, n10165, n12394, n10164, n10176, n10166, n10174,
    n17312, n10167, n10171, n10169, n17313, n10170, n10172, n10173, n10230,
    n10179, n11975, n10178, n10181, n10180, n10235, n10182, n10229, n10200,
    n10183, n10189, n10185, n10184, n10186, n10187, n17306, n10188, n10190,
    n17443, n10194, n10221, n17054, n10193, n10198, n10196, n10195, n10197,
    n10889, n10199, n10890, n17032, n10201, n10205, n10204, n10206, n10236,
    n10208, n10209, n10219, n10211, n10217, n10213, n10248, n10215, n17299,
    n10216, n10218, n10220, n17023, n10223, n10222, n10227, n10225, n10224,
    n10226, n13220, n10228, n16989, n16435, n16990, n10231, n10238, n10240,
    n10239, n10266, n10243, n10244, n10264, n10253, n10246, n10251, n10247,
    n10249, n17292, n10250, n10252, n17465, n10281, n10255, n17005, n10257,
    n10256, n10262, n10260, n10259, n10261, n10288, n16991, n10263, n10291,
    n10265, n10269, n10268, n10296, n10272, n10273, n10293, n10280, n10274,
    n10275, n10300, n17285, n10278, n10276, n10277, n10279, n17476, n16443,
    n16980, n10283, n10282, n10287, n10285, n10284, n10286, n16591, n10289,
    n10913, n10290, n10292, n10294, n10298, n10297, n10322, n10320, n17278,
    n10299, n10301, n10331, n16779, n10304, n10302, n10303, n10305, n10308,
    n10307, n10318, n10316, n10310, n10309, n10313, n10311, n10393, n16950,
    n10314, n10315, n10317, n11105, n10323, n10326, n10325, n10327, n10356,
    n10329, n10330, n17271, n10332, n10333, n10335, n10337, n10338, n10336,
    n10340, n10385, n10343, n10341, n10342, n10344, n10347, n16940, n10346,
    n10351, n10349, n10348, n10350, n10353, n10931, n16931, n10352, n10932,
    n10359, n10358, n10360, n10381, n10362, n10363, n10378, n10364, n16817,
    n10367, n10365, n10366, n10368, n10369, n10370, n13923, n10372, n10371,
    n10376, n10374, n10373, n10375, n10377, n10379, n10384, n10383, n10403,
    n10401, n17258, n10391, n10412, n17259, n10389, n10387, n10388, n10390,
    n10392, n13910, n10395, n10394, n10400, n10398, n10397, n10399, n13893,
    n10404, n10406, n10405, n10407, n10430, n10409, n10410, n17252, n10419,
    n10411, n10413, n10414, n17253, n10417, n10415, n10416, n10418, n10421,
    n10420, n10427, n10422, n10423, n13881, n10425, n10424, n10426, n10947,
    n10432, n10431, n10461, n10435, n10436, n10458, n10437, n10444, n10439,
    n10442, n17246, n10443, n10445, n10446, n13856, n10449, n10448, n10453,
    n10451, n10450, n10452, n10456, n13830, n10454, n10455, n10457, n10459,
    n10463, n10462, n10488, n10464, n10474, n10466, n10472, n10468, n10470,
    n10469, n10471, n10473, n10475, n10476, n10478, n10477, n13818, n10480,
    n10479, n10485, n10483, n10482, n10484, n10487, n13778, n10486, n10490,
    n10489, n10512, n10509, n16131, n10496, n10491, n10494, n10492, n16916,
    n10493, n10495, n10497, n10532, n10499, n13789, n10501, n10500, n10505,
    n10503, n10502, n10504, n10506, n10507, n13749, n10510, n10513, n10516,
    n10515, n10538, n10519, n10520, n10537, n10526, n10524, n10525, n10527,
    n10529, n10528, n10531, n10530, n10535, n13766, n10533, n10534, n17558,
    n13777, n11112, n11111, n10541, n10540, n10544, n10545, n10547, n10549,
    n10548, n10551, n12197, n10550, n10553, n13738, n10555, n10554, n10559,
    n10557, n10556, n10558, n13752, n10560, n10561, n10565, n10564, n10585,
    n10604, n10568, n10566, n10567, n14038, n10570, n13715, n10572, n10571,
    n10576, n10574, n10573, n10575, n10577, n13729, n10578, n10580, n10579,
    n10603, n10583, n10584, n10588, n10586, n10592, n10590, n10589, n10591,
    n11769, n10594, n12358, n10593, n13691, n10601, n10597, n10596, n10599,
    n10598, n10600, n17567, n13656, n10602, n10606, n10615, n10613, n10608,
    n10607, n10609, n10644, n10611, n10612, n10614, n10619, n10617, n10616,
    n10649, n10621, n12336, n10620, n13667, n10628, n10624, n10623, n10626,
    n10625, n10627, n17570, n13408, n11014, n11015, n10632, n10631, n10630,
    n10653, n10643, n14226, n10634, n14228, n10633, n10636, n13645, n10642,
    n10638, n10637, n10640, n10639, n10641, n17573, n11022, n13655, n11023,
    n13246, n10645, n10646, n10655, n10654, n10656, n10671, n10658, n10659,
    n12340, n10662, n13623, n10670, n10666, n10665, n10668, n10667, n10669,
    n17576, n13249, n11033, n10673, n10672, n10674, n10724, n10676, n10677,
    n10679, n10680, n10714, n10682, n14221, n10681, n13478, n13476, n10690,
    n10686, n10685, n10688, n10687, n10689, n17579, n13251, n11089, n10697,
    n10692, n10691, n10693, n10722, n10695, n10696, n10707, n14215, n10699,
    n10701, n10700, n10706, n10737, n13573, n10704, n10703, n10705, n11051,
    n13560, n10728, n10709, n10708, n10710, n10746, n10712, n10713, n10715,
    n10718, n10721, n10723, n10727, n10725, n10731, n10729, n10730, n10735,
    n10733, n10734, n10736, n10754, n10738, n13547, n10740, n10739, n10744,
    n10742, n10741, n10743, n11087, n10749, n10748, n10761, n10750, n14202,
    n14203, n10751, n10753, n10752, n10759, n10757, n13532, n10755, n10756,
    n10758, n10762, n10765, n10764, n10799, n10766, n10767, n14195, n10770,
    n14197, n10769, n13506, n10772, n10771, n10774, n10773, n17591, n13273,
    n10776, n10775, n10779, n10778, n13514, n12424, n12423, n10806, n10784,
    n10783, n10786, n10785, n10788, n10787, n10791, n10789, n10790, n10798,
    n10801, n10792, n10796, n10794, n10793, n10795, n10797, n10800, n10802,
    n10804, n10805, n11078, n10808, n10807, n10809, n11074, n10810, n10829,
    n10813, n10820, n11124, n12431, n10821, n10823, n17365, n16570, n17163,
    n10827, n10830, n10832, n10831, n10835, n10833, n10834, n10842, n10839,
    n10838, n10840, n17170, n10841, n10846, n10844, n10843, n10845, n10850,
    n10848, n10847, n10849, n10852, n10851, n10861, n10859, n10854, n10853,
    n10868, n13212, n10860, n16603, n10856, n10855, n10857, n10858, n10863,
    n10862, n10864, n10867, n10872, n10870, n10869, n10871, n10874, n10873,
    n10880, n12459, n10875, n10879, n10877, n10876, n10878, n10881, n13217,
    n10882, n10883, n10884, n10886, n10885, n10897, n10887, n10896, n10894,
    n10892, n10891, n10893, n10895, n10898, n10900, n10899, n10910, n13223,
    n10904, n10902, n10901, n10903, n10914, n16442, n10906, n10907, n10909,
    n10908, n10918, n10911, n10912, n10916, n10915, n10917, n10919, n10927,
    n10923, n10922, n10925, n10924, n10926, n10929, n10928, n10930, n10934,
    n10933, n10935, n14125, n10937, n10936, n10939, n10938, n10940, n10942,
    n10941, n10951, n10944, n10943, n10950, n10945, n10946, n10949, n10948,
    n10953, n10952, n10954, n10959, n10957, n10956, n10958, n10965, n10961,
    n10960, n10967, n10963, n10962, n10966, n10964, n10969, n10968, n10970,
    n10972, n10971, n10975, n10973, n10974, n10976, n13235, n10977, n10979,
    n10978, n10983, n10981, n10980, n10982, n10985, n10984, n10987, n10986,
    n10989, n10988, n10994, n11091, n10993, n10991, n10990, n10992, n13240,
    n10995, n10997, n10996, n11003, n13241, n10998, n11002, n11001, n11006,
    n11004, n13242, n11005, n11007, n11010, n11009, n11012, n11011, n11013,
    n11017, n11016, n11019, n11018, n11020, n13245, n11021, n11025, n11024,
    n11026, n11028, n11027, n11030, n11029, n11035, n11034, n11036, n11038,
    n11037, n11040, n11039, n11041, n11043, n11042, n11044, n11046, n11045,
    n11048, n11047, n11053, n11052, n11054, n11056, n11055, n11058, n11057,
    n11059, n11061, n11060, n11062, n11065, n11064, n11067, n11066, n11071,
    n11070, n11076, n11075, n11080, n11079, n11081, n13269, n11083, n11084,
    n12580, n11086, n13267, n11117, n13555, n13587, n13250, n13727, n11092,
    n13232, n11098, n17106, n11099, n13211, n17117, n17198, n17148, n11100,
    n11102, n11103, n17058, n11104, n17015, n16963, n16934, n11107, n11108,
    n11109, n11113, n13750, n13775, n13703, n11116, n11118, n12595, n11120,
    n11121, n12335, n11127, n11128, n11153, n11131, n11135, n11136, n11137,
    n11140, n11139, n11141, n11146, n12101, n12598, n11148, n11149, n11151,
    n11150, n11152, n11154, n13271, n11157, n11156, n11161, n11160, n11337,
    n11210, n11170, n11171, n11173, n11186, n11174, n11183, n11178, n11177,
    n11179, n11180, n15310, n11184, n11189, n11192, n11193, n11197, n16125,
    n11202, n11206, n11207, n11209, n15494, n11218, n12402, n15312, n11217,
    n14622, n11359, n11219, n11374, n11409, n11220, n11221, n11222, n11223,
    n11608, n11224, n11225, n11710, n11772, n11800, n11788, n14399, n11828,
    n11226, n14623, n11239, n11235, n11234, n11237, n11236, n11238, n16410,
    n11240, n11242, n11845, n11245, n12246, n11244, n11846, n14520, n11246,
    n11248, n11250, n11702, n11257, n11252, n11255, n11253, n11254, n11256,
    n11258, n11260, n11280, n11262, n11261, n11267, n11264, n11265, n11969,
    n11266, n11268, n11269, n11275, n11273, n11274, n11277, n11279, n11278,
    n15376, n11284, n11283, n11282, n11288, n11287, n11290, n11297, n11983,
    n11292, n11291, n11294, n11293, n15420, n11296, n11298, n11302, n11301,
    n11300, n15424, n11306, n11305, n15425, n11309, n11308, n11314, n11312,
    n11310, n11311, n11313, n11322, n11315, n11318, n11316, n16219, n11317,
    n11320, n11319, n11321, n11323, n11327, n11325, n11324, n11326, n15349,
    n15347, n11328, n15982, n11330, n11329, n11334, n11332, n11331, n11333,
    n11344, n11335, n11340, n11353, n11338, n16213, n11339, n11342, n11341,
    n12861, n11343, n11345, n11348, n11347, n11346, n11349, n15395, n11351,
    n11350, n11358, n11352, n11356, n11354, n16207, n11355, n11357, n15959,
    n11361, n11360, n11365, n11363, n11362, n11364, n11366, n11368, n12204,
    n11370, n11369, n12208, n11371, n11852, n11373, n11372, n11380, n11378,
    n11375, n15943, n11376, n11377, n11379, n11387, n11381, n11385, n11425,
    n11383, n15588, n11384, n11386, n15946, n11388, n11390, n11397, n11393,
    n11392, n11398, n15450, n12202, n11394, n11395, n11396, n11400, n11399,
    n15451, n11402, n11407, n11403, n11404, n11405, n16196, n11406, n11408,
    n11417, n11411, n15914, n11410, n11415, n11413, n11412, n11414, n11416,
    n11418, n11422, n11420, n11419, n11421, n15331, n11423, n11428, n11424,
    n11445, n11426, n16190, n11427, n11429, n16334, n11439, n11432, n11431,
    n11437, n11435, n11453, n15878, n11433, n11434, n11436, n11438, n11440,
    n14410, n11442, n11441, n11443, n11450, n11444, n11448, n11446, n15657,
    n11447, n11449, n16353, n11462, n11452, n11451, n11460, n11458, n11455,
    n11456, n15836, n14419, n11457, n11459, n11463, n11468, n11465, n11464,
    n11469, n14417, n11470, n11471, n11480, n11496, n11473, n11474, n11475,
    n16173, n11478, n11476, n11477, n11479, n11492, n11482, n11481, n11490,
    n11486, n11484, n11483, n11485, n15005, n11488, n11487, n11489, n11491,
    n11493, n11516, n11495, n11494, n11517, n14482, n11497, n15672, n11500,
    n11498, n11499, n11501, n11509, n11502, n11503, n14292, n11506, n11505,
    n11507, n11508, n11510, n14287, n11512, n11511, n14483, n11513, n11514,
    n11515, n11520, n11519, n11518, n14481, n11521, n11528, n11523, n11526,
    n11524, n16167, n11525, n11527, n11537, n11530, n11529, n11535, n11531,
    n14980, n11533, n11532, n11534, n11536, n11538, n11564, n11540, n11539,
    n11565, n14445, n11548, n11541, n11546, n11542, n11576, n11544, n16161,
    n11545, n11547, n11560, n11550, n11549, n11558, n11553, n11552, n11554,
    n14948, n11556, n11555, n11557, n11559, n11561, n11570, n11563, n11562,
    n11571, n14448, n11567, n11566, n12306, n11568, n11574, n11573, n11572,
    n14449, n11575, n11579, n11577, n16155, n11578, n11580, n11589, n11583,
    n11582, n11587, n14924, n11585, n11584, n11586, n11588, n11590, n11604,
    n11591, n11602, n11594, n11593, n11595, n11596, n11599, n11597, n11598,
    n11600, n16150, n11601, n11603, n15166, n11617, n11606, n11605, n11615,
    n11607, n11610, n11609, n11611, n14895, n11613, n11612, n11614, n11616,
    n11618, n11629, n11624, n11620, n11619, n11622, n11621, n14251, n11623,
    n11626, n11625, n14530, n11627, n11633, n11630, n11632, n11641, n11635,
    n11639, n11637, n16144, n11638, n11640, n11649, n11643, n11642, n11647,
    n14872, n11645, n11644, n11646, n11648, n11650, n11653, n11652, n11651,
    n11654, n14358, n11656, n11655, n14359, n11662, n11657, n11660, n11699,
    n16138, n11659, n11661, n11675, n11664, n11663, n11673, n11665, n11668,
    n11667, n11669, n14844, n11671, n11670, n11672, n11674, n11676, n11680,
    n11678, n11677, n11679, n14374, n11685, n11681, n11683, n11682, n11684,
    n15123, n11694, n11686, n14780, n11688, n11687, n11692, n11690, n11689,
    n11691, n11693, n11695, n11726, n11697, n11696, n11727, n14318, n11707,
    n11698, n11700, n11701, n16132, n11705, n11703, n11704, n11706, n11719,
    n11709, n11708, n11717, n11712, n14817, n11715, n11714, n11716, n11718,
    n11720, n14303, n11722, n11721, n14504, n11723, n11724, n11725, n11730,
    n11729, n11728, n11732, n12301, n11731, n15112, n11742, n11734, n14763,
    n11801, n11736, n11735, n11740, n11738, n11737, n11739, n11741, n11743,
    n11759, n11745, n11744, n11760, n12324, n11746, n11755, n14738, n11753,
    n11749, n11748, n11751, n11750, n11752, n11754, n11756, n11764, n11758,
    n11757, n11765, n14326, n11762, n11761, n14322, n11763, n11767, n11766,
    n11771, n12353, n11770, n11780, n14715, n14469, n11778, n11774, n11773,
    n11776, n11775, n11777, n16398, n11779, n11781, n11783, n11782, n14463,
    n15321, n11784, n11794, n11787, n11786, n11792, n14669, n11790, n11789,
    n11791, n11793, n11795, n11818, n11797, n11796, n11819, n14394, n11799,
    n12330, n11798, n11810, n14692, n11808, n11804, n11803, n11806, n11805,
    n11807, n16401, n11809, n11812, n14265, n11814, n11813, n11815, n11817,
    n11822, n11821, n11820, n14393, n11823, n11827, n12348, n11826, n15059,
    n11837, n14645, n11829, n11835, n11831, n11830, n11833, n11832, n11834,
    n16407, n11836, n11838, n11841, n11840, n11839, n11842, n14344, n11844,
    n11843, n14343, n11848, n11847, n11849, n15305, n11850, n11862, n11854,
    n11853, n11860, n11856, n14597, n11858, n11857, n11859, n11861, n11863,
    n11868, n11866, n11865, n11867, n14235, n11869, n11871, n11872, n11873,
    n11874, n11880, n11878, n11876, n11875, n11877, n11879, n11896, n11882,
    n11881, n11886, n11884, n11883, n11885, n11894, n11888, n11887, n11892,
    n11890, n11889, n11891, n11893, n11895, n11901, n11898, n11897, n11899,
    n11900, n11902, n11904, n11906, n11905, n12258, n11907, n11908, n13114,
    n11909, n11911, n11910, n11912, n11952, n14574, n11915, n11914, n11919,
    n11917, n11916, n11918, n11920, n11922, n11928, n11926, n11925, n11927,
    n11930, n11932, n11931, n11964, n16059, n16238, n11935, n11934, n16337,
    n11933, n11962, n12709, n16113, n13112, n11936, n15379, n11937, n15380,
    n11938, n11940, n11939, n11941, n11942, n11960, n11948, n11945, n12251,
    n11947, n11946, n11958, n11950, n11949, n11956, n11954, n11951, n12711,
    n11953, n11955, n11957, n11959, n11961, n11963, n11965, n11968, n11967,
    n11971, n11970, n11981, n11980, n11974, n11978, n14229, n11977, n11979,
    n11987, n11982, n11985, n11984, n11986, n11990, n11989, n11992, n11991,
    n11994, n11993, n11996, n11995, n11998, n11997, n12000, n11999, n12002,
    n12001, n12004, n12003, n12007, n12006, n12009, n12008, n12011, n12010,
    n12013, n12012, n12015, n12014, n12017, n12016, n12019, n12018, n12021,
    n12020, n12023, n12022, n12025, n12024, n12028, n12027, n12030, n12029,
    n12032, n12031, n12034, n12033, n12036, n12035, n12038, n12037, n12040,
    n12039, n12042, n12041, n14453, n12044, n12043, n12046, n12045, n12048,
    n12047, n12050, n12049, n12052, n12051, n14535, n12054, n12053, n12056,
    n12055, n14490, n12058, n12057, n12060, n12059, n12062, n12061, n12064,
    n12063, n12066, n12065, n12654, n12068, n12067, n12070, n12069, n14775,
    n12072, n12071, n12074, n12075, n12086, n15341, n12097, n15830, n12076,
    n15484, n15480, n15479, n12077, n12079, n12078, n15485, n12081, n12080,
    n15515, n12082, n15514, n12083, n12084, n12096, n15818, n12094, n15465,
    n15496, n12087, n15508, n15472, n15473, n12089, n12088, n15507, n15506,
    n12090, n12091, n15530, n12092, n12093, n12095, n12100, n12099, n16556,
    n12103, n12105, n12104, n12106, n12151, n12109, n14210, n12107, n12108,
    n12111, n12143, n12145, n16921, n12170, n16650, n16638, n12171, n12113,
    n12112, n12184, n12114, n12115, n16656, n12116, n16671, n12118, n16672,
    n12120, n12119, n12156, n12121, n12157, n12123, n12122, n16694, n12124,
    n12125, n16704, n12126, n16720, n16719, n12128, n12129, n16743, n12130,
    n12149, n12173, n17219, n12174, n12132, n12131, n12187, n12188, n12134,
    n12133, n16661, n16660, n16662, n12135, n16677, n16676, n16678, n12136,
    n12159, n12137, n12160, n12139, n12138, n16688, n16687, n12140, n16709,
    n16708, n16710, n12141, n16725, n16724, n16726, n12142, n16737, n16735,
    n12147, n12144, n12146, n16911, n12148, n12150, n12154, n12153, n16520,
    n12155, n12165, n12158, n12163, n12161, n12162, n12164, n12167, n12166,
    n12169, n12168, n12179, n12172, n12177, n12175, n12176, n12178, n12181,
    n12180, n12183, n12182, n12193, n12186, n12191, n12189, n12190, n12192,
    n12196, n12195, n12201, n12199, n12198, n12200, n12220, n12218, n15539,
    n12216, n12203, n15452, n12206, n12207, n15454, n12209, n12210, n12214,
    n12212, n16026, n12211, n12213, n12215, n12217, n12219, n13133, n13140,
    n12228, n16053, n13149, n13148, n15920, n13154, n12868, n12221, n15861,
    n12896, n12733, n12731, n12804, n12805, n12732, n12223, n12226, n12225,
    n12224, n12257, n16083, n12227, n16051, n12834, n15986, n12229, n12742,
    n15989, n12231, n12230, n12232, n15987, n12233, n12852, n12234, n12235,
    n12859, n15890, n12888, n15865, n15864, n12240, n12239, n12243, n12244,
    n12267, n12250, n12249, n12255, n12253, n12252, n12254, n12256, n12285,
    n12259, n12262, n12260, n12261, n12263, n12266, n12264, n12265, n12278,
    n12279, n16095, n12276, n16037, n16039, n15938, n15874, n12269, n12270,
    n16350, n12281, n14979, n12274, n12272, n12271, n12273, n12275, n12277,
    n12283, n16352, n12280, n12282, n12284, n12296, n12286, n12293, n12292,
    n12298, n12297, n12300, n12305, n12303, n12302, n12304, n14444, n12317,
    n12308, n12315, n12313, n12311, n12309, n15689, n12310, n12312, n12314,
    n12316, n12321, n12319, n12318, n12320, n12323, n12328, n12326, n12325,
    n12327, n12333, n13113, n13197, n12331, n12332, n12339, n12337, n12338,
    n12344, n12342, n12341, n12343, n12352, n12347, n12350, n12349, n12351,
    n12357, n12355, n12354, n12356, n12362, n12360, n12359, n12361, n12391,
    n17620, n17619, n17624, n17623, n17628, n17627, n17632, n17631, n17636,
    n17635, n17640, n17639, n17644, n17648, n12381, n12379, n12377, n12375,
    n12373, n12371, n12369, n17614, n12367, n12364, n12363, n17599, n17598,
    n12365, n17616, n17615, n12366, n17613, n12368, n17612, n17611, n12370,
    n17610, n17609, n12372, n17608, n17607, n12374, n17606, n17605, n12376,
    n17604, n17603, n12378, n17602, n17601, n12380, n12382, n12383, n12384,
    n12385, n12386, n12387, n12388, n17622, n12389, n17618, n17617, n12390,
    n12393, n12392, n12397, n12396, n12398, n14545, n13090, n15287, n12399,
    n12404, n15293, n12403, n12405, n15003, n14919, n14815, n14762, n14666,
    n12407, n14544, n12416, n12414, n12408, n12690, n12413, n12410, n12409,
    n12412, n12411, n14546, n12415, n12418, n12417, n12421, n12420, n12426,
    n12425, n12428, n12432, n12433, n12437, n12434, n12436, n12435, n16486,
    n16598, n12440, n12441, n16600, n12444, n12443, n12442, n16599, n16460,
    n12446, n12447, n16458, n12450, n12449, n12448, n16459, n16536, n12451,
    n12452, n16538, n12455, n12454, n12453, n16537, n12458, n12457, n16522,
    n16523, n12461, n12465, n12463, n12462, n12464, n16621, n12468, n12466,
    n16431, n12467, n12469, n12470, n12471, n16475, n12472, n12473, n16550,
    n12475, n12476, n16552, n12478, n12477, n16551, n12479, n12480, n16446,
    n12481, n12482, n12483, n12484, n12486, n12485, n16582, n12488, n12489,
    n16500, n12491, n12490, n12493, n12492, n13433, n13309, n12495, n12496,
    n13310, n13307, n13372, n12497, n12498, n13374, n13371, n12499, n12500,
    n12509, n12501, n12502, n12510, n12504, n12503, n12505, n13377, n12506,
    n12507, n12508, n12513, n12514, n12516, n13459, n12517, n12519, n12518,
    n13345, n12521, n13420, n12520, n12523, n12525, n12526, n13358, n12527,
    n12528, n13445, n12529, n12530, n12531, n13331, n12533, n13406, n12535,
    n12537, n12536, n12611, n12613, n12579, n12539, n12573, n12545, n12543,
    n12541, n12540, n12542, n12544, n12561, n12547, n12546, n12551, n12549,
    n12548, n12550, n12559, n12553, n12552, n12557, n12555, n12554, n12556,
    n12558, n12560, n12566, n12563, n12562, n12564, n12565, n12567, n12568,
    n12570, n17357, n12576, n12572, n12574, n12575, n12577, n12578, n12606,
    n12583, n12604, n12585, n13286, n12587, n12589, n12590, n13321, n12591,
    n12592, n13475, n12594, n12593, n12602, n12596, n13314, n12600, n12599,
    n13612, n12601, n12603, n12605, n12607, n12608, n12612, n12614, n12615,
    n12617, n12616, n13472, n12620, n12618, n13295, n12622, n12619, n12621,
    n12623, n12630, n12625, n12627, n12626, n12628, n12633, n12631, n12632,
    n12634, n12635, n12637, n12636, n13543, n12641, n12639, n12638, n12640,
    n12642, n12810, n12925, n14958, n12753, n12933, n12955, n14916, n12756,
    n12940, n12662, n14854, n12766, n14885, n12975, n12989, n14800, n12990,
    n14803, n12777, n12727, n14331, n14714, n12796, n14468, n12795, n13167,
    n12677, n13171, n13177, n12793, n12722, n13074, n12649, n12721, n13127,
    n12651, n12905, n12653, n12655, n14962, n12656, n12657, n12659, n12658,
    n12799, n12798, n14867, n14833, n12981, n12663, n12814, n14809, n12666,
    n12665, n12667, n14786, n12668, n12669, n12670, n14730, n12671, n12672,
    n12673, n12675, n12676, n13043, n13048, n14641, n12679, n12681, n12682,
    n12683, n12720, n12685, n12692, n12687, n12686, n12689, n12688, n16422,
    n13125, n12691, n12699, n12710, n12697, n12696, n12698, n12702, n12701,
    n12705, n12704, n12708, n12707, n12719, n12717, n15940, n12715, n12713,
    n12712, n12714, n12716, n12718, n13085, n13094, n13183, n12723, n13131,
    n12724, n13129, n12797, n12728, n12729, n12767, n12730, n12751, n15839,
    n12808, n12734, n12735, n13160, n12738, n15917, n12739, n12740, n12741,
    n12749, n12743, n12744, n12745, n12746, n12747, n13153, n12748, n12750,
    n12768, n12765, n12752, n12754, n12755, n12757, n12763, n12758, n12760,
    n12762, n12764, n12770, n12772, n12785, n12773, n12775, n12783, n12780,
    n12778, n12779, n12781, n12782, n12784, n12787, n12786, n12790, n13123,
    n13189, n13122, n12827, n14614, n12794, n14690, n14680, n14710, n14756,
    n12816, n12958, n14883, n13135, n16115, n12801, n12803, n12802, n15840,
    n12807, n12809, n14991, n12812, n12813, n14835, n12817, n12818, n12819,
    n12821, n12822, n12823, n12825, n12828, n12832, n12833, n12837, n12836,
    n12838, n12842, n12840, n12841, n15388, n12846, n12844, n12843, n12845,
    n12849, n12848, n12854, n12851, n12850, n12860, n12853, n12855, n12867,
    n12858, n12857, n12871, n12865, n12863, n12862, n12864, n12866, n12877,
    n12870, n12869, n12875, n12873, n12872, n12874, n12876, n12879, n12878,
    n12881, n12880, n12884, n12883, n12885, n12887, n12886, n12889, n12890,
    n12892, n12891, n12893, n12898, n12897, n12899, n13003, n12901, n12900,
    n12907, n12904, n12903, n12913, n12906, n12910, n12909, n12911, n12912,
    n12922, n12915, n12914, n12921, n12920, n12918, n12917, n12919, n12931,
    n12923, n12924, n12927, n12926, n12928, n12930, n12932, n12935, n12934,
    n12937, n12936, n12971, n12939, n12938, n12970, n12944, n12942, n12941,
    n12943, n12969, n12946, n12945, n12963, n12948, n12947, n12962, n12952,
    n12950, n12949, n12951, n12953, n12954, n12957, n12956, n12960, n12965,
    n12964, n12966, n12968, n12973, n12972, n12977, n12976, n12978, n12980,
    n12979, n12982, n12983, n12988, n12986, n12985, n12987, n12992, n12991,
    n12993, n12996, n12995, n13001, n12999, n12998, n13000, n13007, n13005,
    n13004, n13006, n13008, n13009, n13013, n13012, n13014, n13019, n13016,
    n13018, n13025, n13023, n13022, n13024, n13027, n13026, n13028, n13030,
    n13029, n13031, n13033, n13032, n13038, n13035, n13034, n13037, n13036,
    n13040, n13039, n13042, n13046, n13045, n13051, n13050, n13052, n13054,
    n13053, n13055, n13057, n13056, n13058, n13060, n13059, n13061, n13067,
    n13063, n13066, n13065, n13062, n13070, n13069, n13071, n13072, n13079,
    n13077, n13076, n13078, n13081, n13080, n13084, n13083, n13086, n13087,
    n13089, n13088, n13093, n13091, n13092, n13097, n13095, n13096, n13101,
    n13099, n13100, n13108, n13111, n13118, n13116, n13115, n13117, n13200,
    n13119, n13124, n13188, n13128, n13187, n13130, n13182, n13138, n13136,
    n13137, n13139, n13141, n13145, n13144, n13147, n13146, n13152, n15921,
    n13150, n13151, n13158, n13156, n13155, n13157, n13159, n13162, n13163,
    n13165, n13166, n13170, n13172, n13173, n13176, n13178, n13181, n13185,
    n13184, n13186, n13194, n13193, n13196, n13195, n13199, n13201, n13203,
    n17169, n13205, n13206, n13209, n13208, n17143, n13210, n13213, n13216,
    n13215, n17077, n13218, n13221, n13222, n16960, n13225, n13227, n13228,
    n13826, n13229, n13233, n13236, n13238, n13239, n13243, n13247, n13248,
    n13584, n13474, n13252, n13256, n13257, n13264, n13262, n13261, n13263,
    n13265, n17446, n13285, n13270, n13268, n13278, n13272, n13515, n13276,
    n13275, n13277, n13529, n17059, n17001, n16984, n16953, n13909, n13847,
    n13788, n13666, n13643, n13530, n17502, n13282, n13281, n13283, n13284,
    n13288, n13508, n13289, n13292, n13296, n13306, n13304, n13298, n13297,
    n13562, n13302, n13300, n13299, n13301, n13303, n13305, n13308, n13312,
    n13311, n13313, n13328, n16604, n13462, n13316, n13448, n13315, n13326,
    n13324, n13318, n13319, n13320, n13322, n16816, n13323, n13325, n13327,
    n13332, n13333, n13343, n13341, n13337, n13335, n13334, n13336, n13339,
    n13338, n13340, n13342, n13346, n13347, n13357, n13351, n13348, n13349,
    n16915, n13350, n13353, n13352, n13355, n13354, n13356, n13360, n13370,
    n13368, n13364, n13362, n13361, n13363, n13366, n13365, n13367, n13369,
    n13373, n13490, n13376, n13375, n13489, n13378, n13380, n13381, n13391,
    n13383, n13382, n13389, n13387, n13385, n16852, n13386, n13388, n13390,
    n13394, n13404, n13398, n13396, n16865, n13397, n13402, n13400, n13399,
    n13401, n13403, n13407, n13418, n13416, n13412, n13410, n13409, n13411,
    n13414, n13413, n13415, n13417, n13421, n13431, n13425, n13423, n13422,
    n13424, n13427, n13426, n13429, n13428, n13430, n13434, n13435, n13444,
    n13437, n13436, n13442, n13440, n13438, n16798, n13439, n13441, n13443,
    n13447, n13458, n13456, n13452, n13450, n13449, n13451, n13454, n13453,
    n13455, n13457, n13461, n13471, n13465, n13463, n16891, n13464, n13467,
    n13466, n13469, n13468, n13470, n13473, n13488, n13486, n13477, n13596,
    n13480, n13479, n13484, n13482, n13481, n13590, n13483, n13485, n13487,
    n13492, n13493, n13504, n13497, n13496, n13502, n13500, n13498, n16830,
    n13499, n13501, n13503, n13522, n13507, n13944, n13513, n13509, n13511,
    n13512, n13521, n13519, n13946, n13954, n13523, n13516, n13517, n13518,
    n13520, n13952, n13528, n13526, n13524, n13525, n13527, n13536, n13534,
    n13533, n13535, n13568, n17213, n13677, n13540, n13542, n13544, n13968,
    n13545, n13553, n13963, n13552, n13550, n13548, n13549, n13551, n13962,
    n13556, n13565, n13561, n13563, n13564, n13567, n13566, n13582, n17176,
    n13580, n13571, n13570, n13973, n13578, n13576, n13574, n13575, n13577,
    n13579, n13581, n13585, n13586, n13983, n13602, n13589, n13592, n13591,
    n13988, n13594, n13595, n13597, n13598, n13600, n13601, n13603, n13604,
    n13993, n13619, n13609, n13611, n13614, n13613, n13999, n13994, n13616,
    n13617, n13618, n13621, n13620, n13628, n13626, n13624, n13625, n13627,
    n14004, n13640, n13632, n13633, n13638, n13636, n13635, n13637, n13642,
    n13641, n13653, n13651, n14005, n13649, n13647, n17190, n13646, n13648,
    n13650, n13652, n14015, n13662, n13660, n13658, n13657, n13659, n13661,
    n14023, n13664, n13663, n13676, n13674, n14016, n13672, n13670, n13668,
    n13669, n13671, n13673, n13675, n14026, n13700, n13683, n13681, n13682,
    n13687, n13685, n13684, n13686, n14031, n13689, n13688, n13698, n14027,
    n13696, n13694, n13692, n13693, n13695, n13697, n13699, n14036, n13710,
    n13704, n13708, n13706, n13705, n13707, n13709, n14044, n13712, n13711,
    n13724, n13722, n14037, n13720, n13718, n13716, n13717, n13719, n13721,
    n13723, n14047, n13735, n13728, n13733, n13731, n13730, n13732, n13734,
    n14055, n13737, n13736, n13747, n13745, n14048, n13743, n13741, n13739,
    n13740, n13742, n13744, n13746, n14058, n13762, n13751, n13756, n13754,
    n13753, n13755, n14064, n13758, n14059, n13759, n13760, n13761, n13765,
    n13763, n13764, n13772, n17144, n13770, n13768, n13767, n13769, n13771,
    n14069, n13784, n13776, n13782, n13780, n13779, n13781, n13783, n14077,
    n13786, n16896, n13785, n13798, n13796, n14070, n13794, n13792, n13790,
    n13791, n13793, n13795, n13797, n14080, n13812, n13802, n13804, n13810,
    n13808, n13807, n13809, n13811, n14087, n14081, n13814, n13815, n13817,
    n16877, n13816, n13824, n13822, n13820, n13819, n13821, n13823, n13863,
    n13828, n13829, n13855, n13844, n13831, n13867, n13866, n13865, n13834,
    n13836, n13842, n13840, n13839, n13841, n13843, n14096, n13851, n13846,
    n13848, n14093, n13849, n13850, n13854, n13852, n13853, n13862, n14090,
    n13860, n13858, n13857, n13859, n13861, n14100, n13864, n13877, n13870,
    n13868, n13869, n13875, n13873, n13872, n13874, n13876, n13880, n13878,
    n13879, n13890, n13888, n14101, n13886, n13884, n13882, n13883, n13885,
    n13887, n13889, n14111, n13904, n13894, n13896, n13902, n13900, n13899,
    n13901, n13903, n14120, n13907, n13905, n13906, n13919, n13917, n14112,
    n13915, n13913, n13911, n13912, n13914, n13916, n13918, n13922, n13921,
    n13925, n13924, n13931, n14123, n13929, n14124, n13927, n13928, n13930,
    n13943, n13941, n13934, n13939, n13937, n13936, n13938, n13940, n14131,
    n13942, n13947, n13950, n13957, n13955, n13956, n14136, n13959, n13958,
    n13960, n13966, n13965, n13967, n13969, n13971, n13970, n13978, n13976,
    n13975, n13977, n13979, n14142, n13982, n13981, n13990, n13985, n13987,
    n13989, n14145, n13992, n13991, n14001, n13997, n13996, n13998, n14000,
    n14148, n14003, n14002, n14010, n14008, n14007, n14009, n14011, n14151,
    n14014, n14013, n14021, n14019, n14018, n14020, n14022, n14154, n14025,
    n14024, n14033, n14029, n14028, n14030, n14032, n14157, n14035, n14034,
    n14042, n14040, n14039, n14041, n14043, n14160, n14046, n14045, n14053,
    n14051, n14050, n14052, n14054, n14163, n14057, n14056, n14066, n14062,
    n14061, n14063, n14065, n14166, n14068, n14067, n14075, n14073, n14072,
    n14074, n14076, n14169, n14079, n14078, n14085, n14083, n14082, n14084,
    n14086, n14172, n14089, n14088, n14095, n14092, n14094, n14097, n14099,
    n14098, n14106, n14104, n14103, n14105, n14108, n14178, n14110, n14109,
    n14118, n14116, n14115, n14117, n14119, n14181, n14122, n14121, n17481,
    n14129, n14127, n14126, n14128, n14130, n14133, n14132, n14134, n14138,
    n14137, n14140, n14144, n14143, n14147, n14146, n14150, n14149, n14153,
    n14152, n14156, n14155, n14159, n14158, n14162, n14161, n14165, n14164,
    n14168, n14167, n14171, n14170, n14174, n14173, n14177, n14176, n14180,
    n14179, n14183, n14182, n14186, n14185, n14194, n14188, n14189, n14192,
    n14190, n14191, n14193, n15285, n14201, n14199, n14198, n14200, n15292,
    n14207, n14205, n14204, n14206, n15298, n14212, n14209, n14211, n15304,
    n14219, n14217, n14216, n14218, n14225, n14223, n14222, n14224, n15318,
    n14234, n14232, n14230, n14231, n14233, n14236, n14238, n14240, n14250,
    n14248, n14246, n14244, n14242, n14241, n14243, n14245, n14247, n14249,
    n14253, n14255, n14264, n14262, n14260, n14256, n15722, n14258, n14257,
    n14259, n14261, n14263, n14268, n14392, n14267, n14391, n14273, n14271,
    n14270, n14272, n14274, n14285, n14691, n14283, n14275, n14281, n14279,
    n14277, n14276, n14278, n14280, n14282, n14284, n14286, n14486, n14288,
    n14484, n14290, n14291, n14302, n14300, n14293, n15646, n14295, n14294,
    n14298, n14297, n14299, n14301, n14305, n14304, n14502, n14319, n14307,
    n14308, n14317, n14315, n14313, n14309, n15808, n14311, n14310, n14312,
    n14314, n14316, n14321, n14430, n14429, n14325, n14324, n14328, n14330,
    n14342, n14340, n14335, n14333, n14332, n14334, n14338, n14336, n14337,
    n14339, n14341, n14346, n14347, n14357, n14644, n14355, n14351, n14349,
    n14348, n14350, n14353, n14352, n14354, n14356, n14360, n14362, n14373,
    n14371, n14369, n14367, n14365, n15755, n14366, n14368, n14370, n14372,
    n14380, n14376, n14377, n14379, n14381, n14390, n14388, n14386, n14382,
    n15774, n14384, n14383, n14385, n14387, n14389, n14396, n14395, n14397,
    n14409, n14407, n14405, n14398, n14401, n14400, n14403, n14402, n14404,
    n14406, n14408, n14413, n14412, n15364, n14415, n14414, n14416, n14418,
    n14428, n14426, n14420, n15635, n14422, n14421, n14424, n14423, n14425,
    n14427, n14431, n14443, n14441, n14432, n14439, n14435, n14433, n14434,
    n14437, n14436, n14438, n14440, n14442, n14446, n14451, n14450, n14452,
    n14462, n14460, n14458, n14454, n15702, n14456, n14455, n14457, n14459,
    n14461, n14465, n14467, n14480, n14478, n14476, n14474, n14472, n14471,
    n14473, n14475, n14477, n14479, n14488, n14485, n14487, n14489, n14499,
    n14497, n14495, n14491, n15677, n14493, n14492, n14494, n14496, n14498,
    n14501, n14507, n14505, n14506, n14508, n14518, n14816, n14516, n14514,
    n14510, n15791, n14512, n14511, n14513, n14515, n14517, n14528, n14526,
    n14524, n14522, n14521, n14523, n14525, n14527, n14532, n14543, n14541,
    n14539, n14534, n15736, n14537, n14536, n14538, n14540, n14542, n14551,
    n14549, n15017, n14554, n14547, n14548, n14550, n15015, n14558, n14556,
    n14553, n14555, n14557, n14561, n14566, n14564, n14563, n14565, n14570,
    n14569, n14572, n14571, n14583, n14581, n14579, n14577, n14575, n14576,
    n14578, n14580, n14582, n14585, n14591, n14589, n14588, n14590, n15039,
    n14593, n14592, n14603, n15040, n14595, n14643, n14601, n14599, n14598,
    n14600, n14602, n14606, n14607, n14613, n14611, n14610, n14612, n14618,
    n14615, n15045, n14617, n15053, n14620, n14619, n14632, n14630, n15046,
    n14628, n14626, n14624, n14625, n14627, n14629, n14631, n14634, n14638,
    n14636, n14635, n14637, n14640, n14639, n14653, n15057, n14651, n15058,
    n14649, n14647, n14646, n14648, n14650, n14652, n14655, n14659, n14657,
    n14656, n14658, n15075, n15068, n14662, n14732, n14675, n14664, n14665,
    n14668, n14667, n15071, n14673, n16092, n14671, n14670, n14672, n14674,
    n14676, n14677, n14679, n14678, n14682, n14686, n14684, n14683, n14685,
    n15086, n14688, n14687, n14700, n15078, n14698, n15079, n14696, n14694,
    n14693, n14695, n14697, n14699, n14702, n14707, n14705, n14704, n14706,
    n15097, n14709, n14708, n14723, n15089, n14721, n14712, n15090, n14719,
    n14717, n14716, n14718, n14720, n14722, n14725, n14729, n14727, n14726,
    n14728, n15107, n15100, n14744, n14734, n14736, n15103, n14742, n14740,
    n14739, n14741, n14743, n14745, n14746, n14748, n14747, n14750, n14755,
    n14753, n14752, n14754, n14759, n15110, n14758, n15118, n14761, n14760,
    n14771, n14769, n15111, n14767, n14765, n14764, n14766, n14768, n14770,
    n14773, n14779, n14777, n14776, n14778, n15129, n14781, n14782, n14783,
    n14785, n15827, n14784, n14798, n14787, n14788, n15121, n14796, n14791,
    n15122, n14794, n14793, n14795, n14797, n14801, n14802, n14808, n14806,
    n14805, n14807, n14811, n15132, n14810, n15140, n14814, n14812, n14813,
    n14826, n14824, n15133, n14822, n14820, n14818, n14819, n14821, n14823,
    n14825, n14827, n14832, n14830, n14829, n14831, n14839, n14837, n14836,
    n15143, n14838, n15151, n14842, n14840, n14841, n14853, n14851, n15144,
    n14849, n14847, n14845, n14846, n14848, n14850, n14852, n14855, n14857,
    n14858, n14863, n14861, n14860, n14862, n15161, n14866, n14864, n14865,
    n14880, n15154, n14878, n14869, n14870, n15157, n14876, n14874, n14873,
    n14875, n14877, n14879, n14882, n14891, n14894, n14889, n14887, n14886,
    n14888, n14890, n15172, n14893, n15741, n14892, n14904, n15164, n14902,
    n15165, n14900, n14898, n14896, n14897, n14899, n14901, n14903, n14906,
    n14912, n14910, n14909, n14911, n15183, n14915, n14913, n14914, n14932,
    n15176, n14930, n14921, n14923, n15179, n14928, n14926, n14925, n14927,
    n14929, n14931, n14934, n14943, n14947, n14941, n14939, n14938, n14940,
    n14942, n15194, n14946, n14944, n14945, n14957, n15186, n14955, n15187,
    n14953, n14951, n14949, n14950, n14952, n14954, n14956, n14960, n14961,
    n14971, n15197, n14969, n14967, n14966, n14968, n14970, n15204, n14974,
    n14972, n14973, n14988, n14986, n14976, n14978, n15200, n14984, n14982,
    n14981, n14983, n14985, n14987, n14990, n14999, n15002, n14997, n14995,
    n14994, n14996, n14998, n15215, n15001, n15675, n15000, n15014, n15207,
    n15012, n15208, n15010, n15004, n15008, n15006, n15007, n15009, n15011,
    n15013, n15020, n15018, n15019, n15218, n15022, n15021, n15029, n15027,
    n15026, n15028, n15030, n15221, n15033, n15032, n15037, n15036, n15038,
    n15042, n15056, n15041, n15224, n15044, n15043, n15051, n15049, n15048,
    n15050, n15052, n15227, n15055, n15054, n15063, n15061, n15060, n15062,
    n15064, n15230, n15067, n15066, n15073, n15070, n15072, n15074, n15233,
    n15077, n15076, n15084, n15082, n15081, n15083, n15085, n15236, n15088,
    n15087, n15095, n15093, n15092, n15094, n15096, n15239, n15099, n15098,
    n15105, n15102, n15104, n15106, n15242, n15109, n15108, n15116, n15114,
    n15113, n15115, n15117, n15245, n15120, n15119, n15127, n15125, n15124,
    n15126, n15128, n15248, n15131, n15130, n15138, n15136, n15135, n15137,
    n15139, n15251, n15142, n15141, n15149, n15147, n15146, n15148, n15150,
    n15254, n15153, n15152, n15159, n15156, n15158, n15160, n15257, n15163,
    n15162, n15170, n15168, n15167, n15169, n15171, n15260, n15174, n15173,
    n15181, n15178, n15180, n15182, n15263, n15185, n15184, n15192, n15190,
    n15189, n15191, n15193, n15266, n15196, n15195, n15202, n15199, n15201,
    n15203, n15269, n15206, n15205, n15213, n15211, n15210, n15212, n15214,
    n15272, n15217, n15216, n15220, n15219, n15223, n15222, n15226, n15225,
    n15229, n15228, n15232, n15231, n15235, n15234, n15238, n15237, n15241,
    n15240, n15244, n15243, n15247, n15246, n15250, n15249, n15253, n15252,
    n15256, n15255, n15259, n15258, n15262, n15261, n15265, n15264, n15268,
    n15267, n15271, n15270, n15274, n15273, n15284, n15278, n15279, n15282,
    n15280, n15281, n15283, n15291, n15289, n15288, n15290, n15297, n15295,
    n15294, n15296, n15303, n15301, n15299, n15300, n15302, n15308, n15306,
    n15307, n15316, n15311, n15314, n15313, n15315, n15325, n15320, n15323,
    n15322, n15324, n15329, n15327, n15328, n15340, n15330, n15595, n15338,
    n15332, n15334, n15336, n15335, n15337, n15339, n15342, n15346, n15344,
    n15343, n15345, n15358, n15350, n15353, n15351, n15354, n15356, n15355,
    n15357, n15359, n15611, n15363, n15361, n15360, n15362, n15370, n15366,
    n15368, n15367, n15369, n15371, n15373, n15372, n15387, n15377, n15385,
    n15381, n15434, n15383, n15382, n15384, n15386, n15390, n15389, n15408,
    n15391, n15523, n15406, n15393, n15400, n15398, n15397, n15399, n15401,
    n15404, n15403, n15405, n15407, n15410, n15409, n15416, n15413, n15495,
    n15415, n15418, n15417, n15423, n15422, n15433, n15426, n15428, n15431,
    n15430, n15432, n15436, n15435, n15440, n15439, n15556, n15446, n15981,
    n15444, n15443, n15445, n15449, n15448, n15460, n15456, n15453, n15455,
    n15458, n15459, n15461, n15499, n15462, n15463, n15464, n15467, n15466,
    n15469, n15468, n15471, n15470, n15478, n15474, n15476, n15475, n15477,
    n15483, n15481, n15482, n15486, n15488, n15487, n15493, n15491, n15490,
    n15492, n15513, n15498, n15497, n15500, n15503, n15501, n15505, n15504,
    n15535, n15510, n15509, n15511, n15512, n15517, n15516, n15520, n15550,
    n15518, n15519, n15551, n15521, n15522, n15524, n15528, n15526, n15525,
    n15527, n15537, n15542, n15529, n15540, n15532, n15533, n15534, n15536,
    n15538, n15549, n15559, n15544, n15558, n15545, n15547, n15546, n15548,
    n15555, n15570, n15552, n15569, n15553, n15554, n15647, n16202, n15557,
    n15580, n15561, n15560, n15564, n15581, n15562, n15563, n15565, n15566,
    n15568, n15567, n15578, n15572, n15571, n15574, n15573, n15576, n15590,
    n15575, n15577, n15579, n15603, n15583, n15584, n15586, n15587, n15602,
    n15589, n15592, n15911, n15591, n15593, n15613, n15594, n15596, n15600,
    n15598, n15597, n15599, n15601, n15625, n15605, n15606, n15608, n15626,
    n15609, n15624, n15610, n15622, n15612, n15616, n15636, n15614, n15615,
    n15637, n15617, n15618, n15620, n15619, n15621, n15623, n15630, n16185,
    n15627, n15650, n15628, n15629, n15652, n15632, n15631, n15633, n15644,
    n15634, n15642, n15655, n15656, n15638, n15640, n15639, n15641, n15643,
    n15645, n15649, n16179, n15648, n15667, n15668, n15651, n15669, n15654,
    n15665, n15660, n15659, n15658, n15661, n15663, n15673, n15662, n15664,
    n15666, n15685, n15670, n15671, n15684, n15674, n15690, n15691, n15676,
    n15678, n15682, n15680, n15679, n15681, n15683, n15703, n15687, n15700,
    n15688, n15698, n15693, n15692, n15712, n15711, n15694, n15696, n15695,
    n15697, n15699, n15701, n15710, n15718, n15705, n15704, n15706, n15708,
    n15707, n15709, n15717, n15724, n15714, n15713, n15723, n15715, n15716,
    n15747, n15720, n15734, n15721, n15732, n15726, n15725, n15737, n15740,
    n15738, n15727, n15728, n15730, n15729, n15731, n15733, n15735, n15746,
    n15739, n15756, n15757, n15742, n15744, n15761, n15743, n15745, n15753,
    n15750, n15762, n15763, n15751, n15752, n15754, n15770, n15776, n15759,
    n15758, n15775, n15760, n15768, n15781, n15765, n15764, n15766, n15767,
    n15769, n15772, n15771, n15773, n15787, n15802, n15778, n15777, n15801,
    n15779, n15785, n15793, n15782, n15783, n15784, n15786, n15789, n15788,
    n15790, n15800, n15795, n15811, n15810, n15796, n15798, n15797, n15799,
    n15807, n15824, n15804, n15803, n15823, n15805, n15806, n15809, n15822,
    n15813, n15812, n15815, n15814, n15817, n15820, n15819, n15821, n15833,
    n15826, n15825, n15829, n15828, n15831, n15832, n15835, n15834, n15838,
    n15837, n15858, n16351, n15843, n15844, n16356, n16017, n15842, n15856,
    n15846, n15854, n15852, n15850, n15849, n15851, n15853, n16362, n15855,
    n15857, n15860, n15859, n15887, n15862, n15863, n15873, n15866, n15868,
    n16341, n15871, n15870, n15872, n16346, n15884, n15877, n15876, n16338,
    n15880, n15879, n15882, n16335, n15883, n15885, n15886, n15889, n15888,
    n15892, n16323, n15909, n15895, n15897, n15899, n15898, n15901, n15900,
    n16331, n15902, n16327, n15906, n15904, n16321, n15905, n15907, n15908,
    n15910, n15913, n15912, n15916, n15915, n15919, n15970, n15922, n15923,
    n15924, n15936, n15928, n16313, n15934, n15932, n15931, n15933, n15935,
    n16315, n15937, n15939, n16308, n15941, n15942, n15950, n15945, n15944,
    n15948, n15947, n15949, n15953, n15951, n15952, n15955, n15957, n16303,
    n15965, n16298, n15960, n15963, n15962, n15964, n15968, n15966, n15967,
    n15977, n15971, n15976, n15974, n15973, n15975, n16305, n15978, n15980,
    n15979, n16285, n15983, n15984, n15994, n15985, n15993, n16016, n15988,
    n16002, n15991, n15990, n15992, n16293, n15995, n16001, n15999, n15997,
    n15998, n16000, n16005, n16289, n16004, n16008, n16286, n16007, n16010,
    n16009, n16013, n16012, n16036, n16273, n16019, n16015, n16271, n16018,
    n16034, n16022, n16032, n16030, n16024, n16028, n16027, n16029, n16031,
    n16280, n16033, n16035, n16038, n16260, n16067, n16044, n16043, n16264,
    n16050, n16048, n16047, n16049, n16058, n16052, n16054, n16056, n16057,
    n16266, n16060, n16062, n16061, n16064, n16063, n16065, n16066, n16069,
    n16068, n16073, n16072, n16075, n16082, n16080, n16079, n16081, n16086,
    n16250, n16085, n16255, n16089, n16256, n16091, n16100, n16094, n16093,
    n16098, n16096, n16097, n16099, n16101, n16103, n16102, n16107, n16106,
    n16112, n16110, n16111, n16121, n16114, n16118, n16117, n16247, n16120,
    n16123, n17226, n16127, n16126, n16130, n16230, n16129, n17232, n16135,
    n16133, n16134, n16137, n16136, n16141, n16139, n16140, n16143, n16142,
    n16147, n16145, n16146, n16149, n16148, n16152, n16151, n16154, n16153,
    n16158, n16156, n16157, n16160, n16159, n16164, n16162, n16163, n16166,
    n16165, n16170, n16168, n16169, n16172, n16171, n16176, n16174, n16175,
    n16178, n16177, n16181, n16180, n16183, n16182, n16187, n16186, n16189,
    n16188, n16193, n16191, n16192, n16195, n16194, n16199, n16197, n16198,
    n16201, n16200, n16204, n16203, n16206, n16205, n16210, n16208, n16209,
    n16212, n16211, n16216, n16214, n16215, n16218, n16217, n16222, n16220,
    n16221, n16224, n16223, n16229, n16227, n16228, n16232, n16231, n16237,
    n16235, n16236, n16243, n16240, n16242, n16249, n16246, n16366, n16248,
    n16259, n16324, n16253, n16252, n16254, n16257, n16369, n16258, n16270,
    n16263, n16262, n16268, n16265, n16267, n16372, n16269, n16282, n16272,
    n16278, n16276, n16275, n16277, n16279, n16375, n16281, n16295, n16284,
    n16288, n16287, n16291, n16290, n16292, n16378, n16294, n16307, n16297,
    n16301, n16300, n16302, n16304, n16381, n16306, n16319, n16312, n16311,
    n16317, n16314, n16316, n16384, n16318, n16333, n16322, n16329, n16325,
    n16326, n16328, n16330, n16387, n16332, n16348, n16336, n16340, n16339,
    n16344, n16342, n16343, n16345, n16390, n16347, n16365, n16355, n16354,
    n16360, n16358, n16359, n16361, n16394, n16364, n16368, n16367, n16371,
    n16370, n16374, n16373, n16377, n16376, n16380, n16379, n16383, n16382,
    n16386, n16385, n16389, n16388, n16392, n16391, n16397, n16396, n16400,
    n16399, n16403, n16402, n16406, n16405, n16409, n16408, n16412, n16411,
    n16415, n16414, n16418, n16417, n16421, n16420, n16424, n16423, n16428,
    n16427, n17052, n16429, n16703, n16441, n16432, n16434, n16433, n16439,
    n16437, n16436, n17050, n16438, n16440, n16444, n16734, n16455, n16447,
    n16453, n16451, n16449, n16448, n16995, n16450, n16452, n16454, n16457,
    n16654, n16471, n16461, n16462, n16467, n16465, n16464, n17154, n16466,
    n16469, n16588, n16468, n16470, n17454, n16473, n16718, n16485, n16476,
    n16483, n16481, n16479, n16478, n17035, n16480, n16482, n16484, n16488,
    n16494, n16492, n16491, n17378, n16493, n16499, n16612, n16495, n16497,
    n16496, n16498, n16502, n16504, n16515, n16778, n16508, n16507, n16936,
    n16509, n16513, n16511, n16510, n16512, n16514, n17421, n16518, n17093,
    n16519, n16533, n16521, n16531, n16524, n16525, n16527, n16529, n16528,
    n16530, n16532, n16535, n16670, n16549, n16539, n16540, n16545, n16543,
    n16542, n17119, n16544, n16547, n16546, n16548, n16553, n16555, n16567,
    n16557, n16565, n16563, n16561, n16560, n17017, n16562, n16564, n16566,
    n16577, n16572, n16571, n16573, n16576, n16579, n17208, n16578, n16581,
    n17367, n16580, n16586, n16585, n16587, n16590, n16589, n16597, n17488,
    n16595, n16760, n16970, n16956, n17489, n16593, n16594, n16596, n16601,
    n16602, n16610, n16607, n16606, n17167, n16609, n16616, n16611, n16614,
    n16613, n16615, n16619, n16686, n16637, n16623, n16635, n16633, n16630,
    n16629, n17084, n16632, n16634, n16636, n16639, n16641, n16640, n16642,
    n16646, n16644, n16643, n16645, n16652, n16648, n16647, n16649, n16651,
    n16653, n16668, n16659, n16657, n16658, n16666, n16664, n16663, n16665,
    n16667, n16669, n16684, n16675, n16673, n16674, n16682, n16680, n16679,
    n16681, n16683, n16685, n16701, n16689, n16690, n16692, n16691, n16699,
    n16697, n16696, n16698, n16700, n16702, n16716, n16707, n16705, n16706,
    n16714, n16712, n16711, n16713, n16715, n16717, n16732, n16723, n16721,
    n16722, n16730, n16728, n16727, n16729, n16731, n16733, n16753, n16755,
    n16736, n16739, n16738, n16754, n16740, n16742, n16741, n16751, n16745,
    n16747, n16761, n16749, n16748, n16750, n16752, n16757, n16756, n16781,
    n17279, n16780, n16758, n16769, n16759, n16767, n16771, n16762, n16770,
    n16763, n16765, n16764, n16766, n16768, n16773, n16772, n16795, n16775,
    n16774, n16793, n16776, n16792, n16777, n16790, n16788, n16783, n16782,
    n16800, n16802, n16785, n16784, n16799, n16786, n16787, n16789, n16791,
    n16810, n16796, n16809, n16797, n16807, n16805, n16801, n16819, n17266,
    n16818, n16803, n16804, n16806, n16808, n16831, n16813, n16832, n16814,
    n16828, n16815, n16826, n16824, n16821, n16820, n16841, n16840, n16822,
    n16823, n16825, n16827, n16829, n16839, n16834, n16833, n16847, n16835,
    n16837, n16836, n16838, n16846, n16843, n16842, n16853, n16854, n16844,
    n16845, n16867, n16849, n16850, n16863, n16851, n16861, n16879, n16856,
    n16855, n16878, n16857, n16859, n16858, n16860, n16862, n16864, n16876,
    n16866, n16885, n16870, n16886, n16871, n16874, n16873, n16875, n16884,
    n16893, n16881, n16880, n16892, n16882, n16883, n16888, n16887, n16917,
    n16918, n16889, n16904, n16890, n16902, n16895, n16894, n16905, n16907,
    n17233, n16906, n16897, n16898, n16900, n16899, n16901, n16903, n16908,
    n16909, n16910, n16912, n16928, n16914, n16926, n16920, n16919, n16923,
    n16925, n16927, n17509, n16930, n16938, n16967, n16932, n16933, n16935,
    n16937, n17513, n16939, n16949, n16942, n16941, n16947, n17503, n16945,
    n16944, n16946, n16948, n16952, n16951, n16977, n16954, n17497, n16959,
    n16957, n16958, n16972, n16962, n17494, n16969, n16965, n16966, n16968,
    n17492, n16971, n16973, n16975, n16974, n16976, n16979, n16978, n16982,
    n16981, n16988, n17482, n16986, n17475, n16985, n16987, n17000, n17014,
    n16992, n16993, n16994, n16996, n16998, n16997, n17480, n16999, n17004,
    n17002, n17003, n17007, n17006, n17013, n17464, n17011, n17470, n17010,
    n17012, n17022, n17016, n17018, n17020, n17019, n17469, n17021, n17025,
    n17024, n17030, n17027, n17031, n17457, n17029, n17047, n17038, n17034,
    n17036, n17037, n17459, n17040, n17456, n17043, n17042, n17044, n17045,
    n17046, n17049, n17051, n17449, n17100, n17053, n17056, n17055, n17063,
    n17447, n17061, n17442, n17060, n17062, n17064, n17066, n17065, n17073,
    n17071, n17070, n17072, n17076, n17431, n17075, n17079, n17435, n17078,
    n17090, n17080, n17086, n17083, n17085, n17439, n17088, n17089, n17092,
    n17094, n17424, n17097, n17427, n17099, n17110, n17101, n17104, n17103,
    n17108, n17422, n17199, n17107, n17109, n17111, n17113, n17112, n17412,
    n17115, n17121, n17118, n17120, n17416, n17122, n17129, n17124, n17123,
    n17127, n17126, n17128, n17132, n17131, n17136, n17408, n17135, n17138,
    n17137, n17140, n17139, n17158, n17398, n17146, n17396, n17145, n17156,
    n17149, n17152, n17151, n17153, n17405, n17155, n17157, n17160, n17159,
    n17184, n17162, n17164, n17165, n17166, n17168, n17175, n17171, n17172,
    n17177, n17385, n17174, n17393, n17181, n17179, n17178, n17180, n17182,
    n17183, n17188, n17386, n17187, n17381, n17195, n17372, n17193, n17192,
    n17194, n17196, n17201, n17376, n17200, n17202, n17203, n17205, n17204,
    n17207, n17211, n17210, n17223, n17215, n17214, n17216, n17217, n17221,
    n17220, n17222, n17359, n17353, n17229, n17228, n17231, n17230, n17235,
    n17234, n17237, n17236, n17242, n17240, n17241, n17244, n17243, n17249,
    n17247, n17248, n17251, n17250, n17255, n17254, n17257, n17256, n17262,
    n17260, n17261, n17264, n17263, n17268, n17267, n17270, n17269, n17275,
    n17273, n17274, n17277, n17276, n17281, n17280, n17283, n17282, n17288,
    n17286, n17287, n17290, n17289, n17295, n17293, n17294, n17297, n17296,
    n17302, n17300, n17301, n17304, n17303, n17309, n17307, n17308, n17311,
    n17310, n17316, n17314, n17315, n17318, n17317, n17323, n17321, n17322,
    n17325, n17324, n17330, n17328, n17329, n17332, n17331, n17337, n17335,
    n17336, n17339, n17338, n17346, n17344, n17345, n17349, n17348, n17356,
    n17354, n17355, n17361, n17360, n17371, n17508, n17364, n17369, n17366,
    n17368, n17517, n17370, n17384, n17375, n17374, n17380, n17377, n17379,
    n17382, n17520, n17383, n17395, n17391, n17389, n17388, n17390, n17392,
    n17523, n17394, n17407, n17397, n17403, n17401, n17400, n17402, n17404,
    n17526, n17406, n17418, n17411, n17410, n17414, n17413, n17415, n17529,
    n17417, n17430, n17420, n17426, n17423, n17425, n17428, n17532, n17429,
    n17441, n17434, n17433, n17437, n17436, n17438, n17535, n17440, n17453,
    n17445, n17444, n17451, n17448, n17450, n17538, n17452, n17463, n17455,
    n17461, n17458, n17460, n17541, n17462, n17474, n17467, n17466, n17468,
    n17472, n17471, n17544, n17473, n17486, n17478, n17477, n17479, n17484,
    n17483, n17547, n17485, n17500, n17490, n17491, n17496, n17495, n17498,
    n17550, n17499, n17516, n17507, n17506, n17511, n17510, n17512, n17554,
    n17515, n17519, n17518, n17522, n17521, n17525, n17524, n17528, n17527,
    n17531, n17530, n17534, n17533, n17537, n17536, n17540, n17539, n17543,
    n17542, n17546, n17545, n17549, n17548, n17552, n17551, n17557, n17556,
    n17560, n17559, n17563, n17562, n17566, n17565, n17569, n17568, n17572,
    n17571, n17575, n17574, n17578, n17577, n17581, n17580, n17584, n17583,
    n17587, n17586, n17590, n17589, n17593, n17592, n17597, n17596, n17600,
    n17621, n17625, n17629, n17633, n17637, n17641, n17645, n17649, n16090;
  assign n13995 = ~n10663 | ~n10662;
  assign n11811 = ~n11923;
  assign n12487 = n12431;
  assign n17409 = ~n17133;
  assign n16014 = n11320 & n11319;
  assign n17227 = ~n10812 ^ n10811;
  assign n9355 = n9360 & n9356;
  assign n10698 = n10245;
  assign n12524 = ~n12624;
  assign n13606 = ~n11032 | ~n11033;
  assign n14977 = n14975 | n15198;
  assign n16310 = ~n15946;
  assign n13384 = ~n14091;
  assign n17505 = ~n10345 | ~n10344;
  assign n12581 = ~n13537 | ~n11082;
  assign n16320 = ~n9597 | ~n11408;
  assign n15080 = ~n11799 | ~n11798;
  assign n15024 = n15025 ^ n14573;
  assign n16274 = ~n16014;
  assign n11216 = ~n11214 | ~P1_IR_REG_31__SCAN_IN;
  assign n12439 = ~n17387;
  assign n15869 = ~n12895 | ~n12896;
  assign n15930 = n11365 | n11364;
  assign n15972 = n11334 | n11333;
  assign n13546 = ~n13968 & ~n17218;
  assign n15286 = ~n9355 | ~n9353;
  assign n11249 = ~n9957 | ~n9959;
  assign n13164 = ~n12776 & ~n12728;
  assign n11063 = ~n10828;
  assign n8992 = n11285;
  assign n12788 = n15035 | n14609;
  assign n13972 = ~n13558 ^ n13557;
  assign n15016 = n12400 & n12399;
  assign n13974 = ~n9202 | ~n10699;
  assign n9827 = ~n12520 | ~n13345;
  assign n15198 = ~n11528 | ~n11527;
  assign n17041 = ~n10219 | ~n10218;
  assign n17095 = ~n10148 | ~n10147;
  assign n17399 = ~n17141;
  assign n16516 = n10157 & n10156;
  assign n16078 = ~n9502 | ~n9095;
  assign n8987 = ~n12902;
  assign n10828 = n10825 & n13538;
  assign n11802 = ~n11307;
  assign n11200 = ~n11192 | ~P1_IR_REG_31__SCAN_IN;
  assign n11196 = ~n11543 | ~n11191;
  assign n12395 = n10357;
  assign n11973 = ~n10177;
  assign n13105 = n13103 & n9498;
  assign n12706 = n9485 & n9858;
  assign n13980 = ~n13565 & ~n13564;
  assign n14012 = ~n13640 & ~n13639;
  assign n14345 = ~n11824 | ~n11823;
  assign n13558 = n13254 | n13253;
  assign n14266 = n9444 & n9445;
  assign n9171 = n9240 & n9238;
  assign n14567 = ~n14559;
  assign n9609 = n14724 | n9611;
  assign n14529 = ~n11632 | ~n11633;
  assign n9272 = ~n13748 | ~n13238;
  assign n15047 = ~n11218 | ~n11217;
  assign n13984 = ~n10682 | ~n10681;
  assign n15035 = ~n11851 | ~n11850;
  assign n14006 = ~n13644;
  assign n11032 = n13995 | n13249;
  assign n13644 = n10634 & n10633;
  assign n14017 = ~n10621 | ~n10620;
  assign n15069 = ~n11785 | ~n11784;
  assign n14049 = ~n10551 | ~n10550;
  assign n13690 = n10594 & n10593;
  assign n11785 = n14226 | n12401;
  assign n14789 = n12777 & n12727;
  assign n13757 = ~n13787 | ~n13788;
  assign n13020 = ~n15101 & ~n14751;
  assign n13825 = n9028 | n9291;
  assign n12299 = ~n10549 | ~n10563;
  assign n14933 = ~n9428 | ~n9099;
  assign n9556 = n10506 & n10487;
  assign n14936 = ~n9392 | ~n9872;
  assign n14060 = ~n9233 | ~n10527;
  assign n15145 = ~n11662 | ~n11661;
  assign n14071 = ~n10496 | ~n10495;
  assign n9643 = n9636 & n16500;
  assign n9595 = ~n15841 | ~n12243;
  assign n12660 = n15177 | n14535;
  assign n15841 = ~n12241 | ~n12242;
  assign n15155 = ~n14363;
  assign n14363 = n11641 & n11640;
  assign n14091 = ~n9221 | ~n10445;
  assign n14114 = ~n10391 | ~n10390;
  assign n11467 = n11466 & n14417;
  assign n15365 = n11442 & n11441;
  assign n16955 = ~n10306 | ~n10305;
  assign n15209 = ~n11480 | ~n11479;
  assign n9483 = n9477 & n12234;
  assign n9491 = ~n15938 & ~n16320;
  assign n15396 = n11351 | n11350;
  assign n16487 = ~n12437 | ~n12434;
  assign n17067 = ~n17432;
  assign n17419 = ~n17095;
  assign n15954 = ~n16006 & ~n12861;
  assign n15411 = n11272 & n11271;
  assign n12098 = ~n12097 & ~n12251;
  assign n16625 = n10133 | n10132;
  assign n17387 = ~n10060 | ~n10059;
  assign n12430 = ~n10026 | ~n10025;
  assign n11864 = ~n11391;
  assign n16046 = n11314 | n11313;
  assign n8995 = n11299;
  assign n16283 = n11342 & n11341;
  assign n12624 = n12445;
  assign n11923 = ~n12248 | ~n12268;
  assign n11391 = n9766 | n12246;
  assign n8990 = ~n8989;
  assign n16463 = ~n10045 | ~n10046;
  assign n9959 = n11248 & n11247;
  assign n12248 = n13107 | n16090;
  assign n12102 = n10089;
  assign n9957 = n9463 & n11246;
  assign n9484 = ~n11290 & ~n9063;
  assign n8988 = n11289;
  assign n10101 = ~n12110 | ~n12394;
  assign n16251 = ~n9517 | ~n9677;
  assign n10089 = ~n12110;
  assign n13191 = n13192 & n16125;
  assign n10234 = ~n10209 | ~n10236;
  assign n11181 = ~n11180 | ~P1_IR_REG_31__SCAN_IN;
  assign n11285 = ~n15286 & ~n11232;
  assign n10012 = ~n10009 | ~n10008;
  assign n12791 = ~n11200 ^ n11199;
  assign n11243 = ~n11204 ^ n11203;
  assign n12422 = ~n10815 ^ n10814;
  assign n10815 = ~n10813 | ~P2_IR_REG_31__SCAN_IN;
  assign n11204 = ~n11202 | ~P1_IR_REG_31__SCAN_IN;
  assign n10207 = n10205 & n10204;
  assign n10361 = n10359 & n10358;
  assign n11229 = n11231 | n11228;
  assign n14227 = ~n11973 & ~P2_STATE_REG_SCAN_IN;
  assign n10812 = n10781 | n10523;
  assign n11198 = ~n11196 | ~P1_IR_REG_31__SCAN_IN;
  assign n10467 = ~n9844 | ~n9845;
  assign n11543 = n11210 & n11208;
  assign n9844 = n10441 & n10466;
  assign n9845 = n10440 & n10439;
  assign n11211 = ~n11176 & ~n11175;
  assign n9978 = ~n9976 & ~n9975;
  assign n11162 = ~n11161 & ~n11160;
  assign n11175 = ~n11169 | ~n11168;
  assign n11176 = ~n9602 | ~n11174;
  assign n11169 = n11166 & n11167;
  assign n11208 = n11163 & n11336;
  assign n10018 = ~n10014 | ~n10013;
  assign n9977 = n10094 & n10090;
  assign n9602 = n11164 & n11165;
  assign n11164 = ~P1_IR_REG_13__SCAN_IN & ~P1_IR_REG_12__SCAN_IN;
  assign n11165 = ~P1_IR_REG_14__SCAN_IN & ~P1_IR_REG_15__SCAN_IN;
  assign P2_U3152 = ~P2_STATE_REG_SCAN_IN;
  assign n11163 = ~P1_IR_REG_5__SCAN_IN & ~P1_IR_REG_4__SCAN_IN;
  assign n10016 = ~P1_ADDR_REG_19__SCAN_IN & ~P1_RD_REG_SCAN_IN;
  assign n11166 = ~P1_IR_REG_20__SCAN_IN & ~P1_IR_REG_19__SCAN_IN;
  assign n11144 = ~P2_IR_REG_25__SCAN_IN;
  assign n9970 = ~P2_IR_REG_23__SCAN_IN & ~P2_IR_REG_22__SCAN_IN;
  assign n10814 = ~P2_IR_REG_20__SCAN_IN;
  assign n14500 = ~n14503 | ~n14304;
  assign n17185 = ~n17373 & ~n16568;
  assign n13329 = ~n12532 & ~n12531;
  assign n13541 = n9311 & n11050;
  assign n12268 = ~n9504 | ~n11243;
  assign n11289 = n9414 & n11232;
  assign n14663 = ~n14713 & ~n15080;
  assign n10481 = ~n10396;
  assign n8989 = ~n10258;
  assign n8991 = ~n11923;
  assign n12429 = ~n10822;
  assign n14573 = n14621 & n9694;
  assign n14552 = n14621 & n9140;
  assign n14621 = ~n14666 & ~n15059;
  assign n11295 = ~n9766;
  assign n8993 = ~n11391;
  assign n8994 = n11299;
  assign n11299 = ~n11924;
  assign n8996 = ~n12581;
  assign n11068 = n13280 & n9918;
  assign n12725 = n15091 & n14331;
  assign n9307 = ~n9950 | ~n9064;
  assign n9800 = n9801 & n13218;
  assign n9801 = ~n9047 | ~n9802;
  assign n9743 = ~n9744 | ~n13052;
  assign n9522 = ~n9743 | ~n13055;
  assign n13064 = ~n13063 | ~n13062;
  assign n13075 = n15025 & n16416;
  assign n11069 = ~n13280 & ~n9918;
  assign n9933 = ~n9937 & ~n9934;
  assign n9618 = ~n9619 & ~n13075;
  assign n9619 = ~n12788;
  assign n9426 = ~n12648 | ~n9010;
  assign n9893 = n9894 & n12731;
  assign n9834 = n16446 & n9835;
  assign n9836 = ~n16552;
  assign n9284 = ~n9285 | ~n13248;
  assign n9285 = ~n9286;
  assign n9809 = n13246 & n13245;
  assign n9557 = n13801 & n10457;
  assign n13833 = n14102 | n13897;
  assign n9289 = ~n9292 | ~n9293;
  assign n9985 = n9984 & n9983;
  assign n9984 = ~P2_IR_REG_13__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n10339 = n10334 & n10333;
  assign n9788 = ~n9791 | ~n11471;
  assign n13098 = ~n15016 & ~n13094;
  assign n9903 = ~n13021;
  assign n9885 = n9886 & n12774;
  assign n9886 = ~n9002 | ~n12766;
  assign n14559 = ~n12720 | ~n12649;
  assign n13169 = ~n13041 | ~n16404;
  assign n12647 = n14724 | n13020;
  assign n9336 = ~n10460 | ~n10459;
  assign n10271 = n10269 & n10268;
  assign n10242 = n10240 & n10239;
  assign n9941 = ~n9942 | ~n11077;
  assign n9942 = ~n9020 | ~n9946;
  assign n16943 = n16953 | n16955;
  assign n17033 = ~n13220 | ~n10228;
  assign n13748 = ~n13237 | ~n13236;
  assign n9215 = ~n9216 | ~n13235;
  assign n9275 = ~n17028 | ~n9108;
  assign n9320 = ~n9321;
  assign n10562 = ~n10543 | ~n10542;
  assign n10514 = ~n10511 | ~n10510;
  assign n9439 = n9440 & n11467;
  assign n9440 = ~n15331 | ~n9441;
  assign n11816 = ~n14394 & ~n11815;
  assign n9437 = ~n16078 | ~n8994;
  assign n9449 = n9450 & n9022;
  assign n9450 = ~n9003 | ~n9453;
  assign n9222 = ~n9733 | ~n9016;
  assign n9730 = ~n9031 | ~n9015;
  assign n11307 = ~n15286 | ~n11232;
  assign n9872 = n9873 & n12656;
  assign n9392 = ~n9394 | ~n9393;
  assign n12241 = n12240 & n12239;
  assign n12242 = ~n9384 | ~n9030;
  assign n9855 = ~n9856 | ~n12682;
  assign n9589 = n9865 & n9590;
  assign n9865 = n9866 & n12798;
  assign n9591 = ~n12658;
  assign n14881 = ~n9604 | ~n9124;
  assign n9607 = ~n14916 & ~n9364;
  assign n9342 = ~n9344 & ~n9343;
  assign n9343 = ~n10746;
  assign n9344 = ~n9960;
  assign n10380 = ~n9911 | ~n10356;
  assign n10345 = n17271 | n10698;
  assign n9776 = ~n9778 | ~n9777;
  assign n9777 = ~n11849;
  assign n9778 = ~n9780;
  assign n9779 = ~n14344;
  assign n14323 = n11759 | n11760;
  assign n11851 = n14213 | n12401;
  assign n16074 = n12225 & n12224;
  assign n12294 = n11874 & n16234;
  assign n12835 = ~n12833 | ~n9402;
  assign n9402 = ~n9403 | ~n9484;
  assign n9403 = n12902 & n9404;
  assign n9396 = ~n9628 | ~n9626;
  assign n9397 = ~n9398 | ~n12931;
  assign n9503 = n9703 & n10935;
  assign n9703 = ~n10940 | ~n9098;
  assign n9724 = ~n9032 | ~n9725;
  assign n9231 = ~n11784;
  assign n9369 = n12764 | n12765;
  assign n11106 = ~n9471 | ~n9046;
  assign n9471 = n9509 & n9572;
  assign n9408 = ~n13028 | ~n9409;
  assign n13044 = ~n13043 | ~n13047;
  assign n13047 = ~n13049;
  assign n9328 = n9704 & n11021;
  assign n9704 = n9705 & n11013;
  assign n9467 = n11007 & n9104;
  assign n9539 = ~n14867;
  assign n12806 = ~n9529 & ~n9528;
  assign n9528 = n15925 | n15891;
  assign n9529 = ~n9530 | ~n9079;
  assign n9532 = ~n14962 & ~n9533;
  assign n9533 = ~n12809 | ~n9534;
  assign n9534 = ~n15869;
  assign n9535 = ~n14991;
  assign n9742 = ~n9743;
  assign n9525 = n9526 & n13061;
  assign n9526 = ~n9522 | ~n9521;
  assign n9523 = ~n13064 | ~n9084;
  assign n9416 = n9417 & n12229;
  assign n9465 = ~n13703;
  assign n9209 = ~n9210 | ~n10602;
  assign n9210 = n11113 & n9211;
  assign n9211 = ~n9947 & ~n9038;
  assign n9917 = ~n9001 | ~n9056;
  assign n9939 = n11090 & n11032;
  assign n9555 = ~n11022;
  assign n9948 = ~n10999;
  assign n9310 = n9548 & n11015;
  assign n9580 = ~n9581;
  assign n9548 = n10602 & n10578;
  assign n9305 = ~n10866 | ~n17409;
  assign n9876 = n14962 & n9877;
  assign n9878 = ~n12653;
  assign n13134 = ~n16088 | ~n11249;
  assign n10711 = n10709 & n10708;
  assign n9261 = ~n12129;
  assign n9750 = ~n13974 & ~n9751;
  assign n9751 = ~n9752;
  assign n10319 = n9306 & n10292;
  assign n9306 = ~n10291 | ~n10290;
  assign n9278 = ~n13210;
  assign n13538 = ~n12424 & ~n17227;
  assign n11094 = ~n9055 | ~n10045;
  assign n9817 = n9818 & n13555;
  assign n11088 = n13964 | n13274;
  assign n9958 = n13250 | n13584;
  assign n9752 = ~n13984 & ~n13995;
  assign n9286 = n9287 & n13247;
  assign n9288 = ~n9811;
  assign n9579 = ~n9580 | ~n9798;
  assign n9219 = ~n9272 | ~n9580;
  assign n9549 = ~n9925 | ~n9926;
  assign n9926 = n10577 & n9927;
  assign n9217 = n9569 & n9120;
  assign n9569 = ~n13825 | ~n9118;
  assign n13204 = ~n11095 | ~n11094;
  assign n9441 = ~n9021;
  assign n11303 = ~n11300 | ~n11301;
  assign n11367 = ~n16296 | ~n11295;
  assign n13126 = ~n15016;
  assign n12815 = ~n12812 & ~n9536;
  assign n9540 = ~n9541 | ~n14680;
  assign n9541 = ~n9542 & ~n14710;
  assign n9542 = n14641 | n14730;
  assign n9612 = n9899 & n9613;
  assign n9899 = n12796 & n9904;
  assign n12238 = n15869 & n15864;
  assign n9615 = ~n9618 | ~n9616;
  assign n9424 = ~n9617 & ~n9425;
  assign n9425 = ~n9897;
  assign n9617 = ~n9618;
  assign n12680 = ~n14642 | ~n14641;
  assign n14609 = ~n16413;
  assign n9390 = n14730 | n9391;
  assign n9860 = n9861 & n13043;
  assign n9862 = ~n9863;
  assign n13041 = ~n15069;
  assign n13021 = ~n15101 | ~n14751;
  assign n9476 = ~n14815 & ~n15134;
  assign n14856 = ~n14881 & ~n12940;
  assign n12959 = n15188 | n14965;
  assign n12222 = n9625 & n9091;
  assign n13143 = ~n16046 & ~n16014;
  assign n12736 = n16046 & n16014;
  assign n9361 = ~P1_IR_REG_30__SCAN_IN | ~P1_IR_REG_31__SCAN_IN;
  assign n9672 = n9673 & n9117;
  assign n9915 = n10401 | n9916;
  assign n9916 = ~n10381;
  assign n10408 = n10406 & n10405;
  assign n10232 = ~n10234 & ~n10231;
  assign n9474 = ~n10235;
  assign n9640 = ~n9643 | ~n9641;
  assign n9823 = ~n9968;
  assign n9821 = ~n16501;
  assign n9242 = ~n13445;
  assign n12445 = ~n12428 | ~n12427;
  assign n10822 = ~n10041 | ~n10040;
  assign n10041 = n10034 & n10033;
  assign n9746 = ~n17319;
  assign n12522 = ~n14049 ^ n12624;
  assign n9379 = n9380 | n9041;
  assign n9380 = ~n9965;
  assign n9830 = n9831 & n12482;
  assign n12512 = ~n13813 ^ n12524;
  assign n12460 = ~n17067 ^ n12624;
  assign n13317 = ~n13287 & ~n12577;
  assign n9710 = ~n9036 | ~n11081;
  assign n9337 = ~n9338 | ~n11077;
  assign n9208 = n11117 & n9093;
  assign n9708 = n9710 & n13537;
  assign n9709 = ~n9196 | ~n9199;
  assign n9196 = n9197 & n9122;
  assign n9246 = ~n16694 | ~n9253;
  assign n9253 = ~n12122;
  assign n9259 = ~n9260 & ~n16743;
  assign n9260 = ~n12128 & ~n9261;
  assign n9257 = ~n9259 | ~n9261;
  assign n13260 = n10825 | n12424;
  assign n13665 = ~n13757 & ~n9759;
  assign n9759 = ~n9760 | ~n13690;
  assign n9796 = ~n9797 | ~n13727;
  assign n11000 = ~n11008 | ~n13656;
  assign n10999 = ~n13690 | ~n17567;
  assign n9763 = ~n9765 | ~n9764;
  assign n10498 = n10447 | n10446;
  assign n9755 = ~n9756 | ~n13909;
  assign n9756 = ~n9757;
  assign n10254 = n10221 | n10220;
  assign n13280 = ~n9919 | ~n10751;
  assign n9919 = n14202 | n10698;
  assign n9311 = ~n9312 | ~n9550;
  assign n9312 = n9551 & n13557;
  assign n11050 = ~n9202 | ~n9086;
  assign n9216 = n9808 | n13801;
  assign n9293 = ~n9570 | ~n13228;
  assign n9570 = ~n9574 | ~n9571;
  assign n9574 = ~n9577 & ~n9575;
  assign n9294 = ~n9573 & ~n9295;
  assign n9295 = ~n13228;
  assign n9273 = ~n9510 & ~n9274;
  assign n9274 = ~n13222;
  assign n9568 = n9271 & n13219;
  assign n9987 = ~n10438 & ~n9980;
  assign n10214 = n10168 | P2_IR_REG_5__SCAN_IN;
  assign n10441 = n10091 & n9977;
  assign n10094 = ~P2_IR_REG_3__SCAN_IN;
  assign n9434 = ~n9436 & ~n9435;
  assign n11461 = n12908 | n11924;
  assign n11389 = n15326 | n11924;
  assign n9667 = ~n13098 & ~n9668;
  assign n9668 = ~n13127;
  assign n13180 = n12788 & n12722;
  assign n9502 = n9496 & n11261;
  assign n9496 = n11262 & n9432;
  assign n15780 = ~n15764 | ~n15765;
  assign n9695 = ~n9698 & ~n9696;
  assign n9696 = ~n9697 | ~n14622;
  assign n9420 = n9421 & n12997;
  assign n9421 = ~n9053 | ~n9423;
  assign n13010 = ~n15112 | ~n13011;
  assign n12997 = n15112 | n13011;
  assign n12895 = n16334 | n15848;
  assign n15891 = ~n12882 | ~n15861;
  assign n9384 = ~n12236 | ~n12859;
  assign n9482 = ~n15969;
  assign n16042 = n9382 & n12227;
  assign n14587 = ~n16416;
  assign n12824 = ~n12721 | ~n13127;
  assign n16023 = n13102 | n11945;
  assign n14616 = ~n12680 | ~n12679;
  assign n14633 = n12648 & n13171;
  assign n12674 = ~n14711 | ~n12672;
  assign n9585 = n9586 & n14867;
  assign n9869 = n9870 & n12799;
  assign n9882 = ~n12753 | ~n9883;
  assign n15961 = ~n16296;
  assign n9520 = n12401 | n17341;
  assign n9519 = ~n11702 | ~n16226;
  assign n9737 = n9739 & n9738;
  assign n9738 = ~n11175 & ~P1_IR_REG_27__SCAN_IN;
  assign n9356 = n9358 & n9357;
  assign n9358 = ~n9359 | ~P1_IR_REG_29__SCAN_IN;
  assign n9357 = ~n15277 | ~n11228;
  assign n9359 = ~n9361;
  assign n10648 = n10647 | n10646;
  assign n10651 = n10650 & n10649;
  assign n11182 = ~n11179 | ~P1_IR_REG_31__SCAN_IN;
  assign n10647 = n10604 | n10606;
  assign n9908 = ~n10514 | ~n9119;
  assign n9907 = ~n10538;
  assign n16124 = ~n9234 ^ n10537;
  assign n9234 = ~n10514 | ~n10513;
  assign n9459 = ~n9376 ^ n9089;
  assign n9914 = ~n9915;
  assign n10382 = ~n10380 | ~n10379;
  assign n9662 = ~n10296;
  assign n10295 = ~n10267 | ~n10266;
  assign n9202 = n14213 | n10698;
  assign n9458 = n9647 & n9650;
  assign n9381 = ~n13379 | ~n9647;
  assign n12610 = n12624 ^ n13644;
  assign n12511 = ~n12512 ^ n9004;
  assign n9493 = n9828;
  assign n10306 = ~n9747 | ~n10732;
  assign n9494 = n13379;
  assign n14102 = ~n10419 | ~n10418;
  assign n14113 = ~n17487;
  assign n12597 = n13317 & n17225;
  assign n16626 = ~n16605;
  assign n9313 = ~n9709 | ~n9710;
  assign n12586 = ~n17352 | ~n11146;
  assign n9268 = ~P2_REG1_REG_2__SCAN_IN;
  assign n9249 = n9250 & n16704;
  assign n9266 = ~n16919 & ~n16920;
  assign n9265 = ~n17098 ^ P2_REG1_REG_19__SCAN_IN;
  assign n9221 = n17245 | n10698;
  assign n9567 = n17265 | n10698;
  assign n17150 = ~n17173;
  assign n17191 = n11082 & n12580;
  assign n13945 = ~n9339 | ~n12110;
  assign n9339 = ~n9340 | ~n10805;
  assign n9340 = ~n15275 | ~n12395;
  assign n13539 = ~n13259 ^ n13258;
  assign n13258 = ~n13267;
  assign n13259 = ~n9815 | ~n9812;
  assign n9812 = n9813 & n13257;
  assign n17487 = ~n17504;
  assign n11130 = ~n11125 | ~P2_IR_REG_31__SCAN_IN;
  assign n17225 = n12586 & n17358;
  assign n9323 = ~n9319 | ~n9087;
  assign n9319 = ~n10467;
  assign n10780 = ~P2_IR_REG_20__SCAN_IN & ~P2_IR_REG_19__SCAN_IN;
  assign n10816 = ~P2_IR_REG_21__SCAN_IN;
  assign n9207 = ~n9908 | ~n9092;
  assign n17272 = n10340 & n10385;
  assign n9597 = n17305 | n12401;
  assign n9770 = n11396 & n9771;
  assign n14252 = ~n11590 ^ n11923;
  assign n9455 = n9776 & n9456;
  assign n9456 = ~n14237;
  assign n11824 = ~n14266 | ~n11816;
  assign n9784 = n9785 & n14323;
  assign n14327 = n11767 | n11766;
  assign n15091 = ~n11771 | ~n11770;
  assign n11551 = n11504 & n11222;
  assign n9781 = ~n14343;
  assign n9782 = ~n14345 | ~n14344;
  assign n11943 = n12294 & n12258;
  assign n9401 = ~n9507;
  assign n15604 = ~n9186 | ~n9112;
  assign n15719 = ~n15704 & ~n15705;
  assign n12085 = ~n11186 & ~n12073;
  assign n13082 = ~n12404 | ~n12403;
  assign n15025 = ~n11912 | ~n11264;
  assign n11454 = n11409 | n11220;
  assign n15023 = ~n14568 ^ n14567;
  assign n16357 = ~n13003 | ~n13192;
  assign n16309 = n16245 | n13191;
  assign n12295 = ~n12290 & ~n12289;
  assign n12289 = ~n12288 | ~n16239;
  assign n12290 = n12286 | n15378;
  assign n16245 = n13114 | n9504;
  assign n11870 = n15319 | P1_B_REG_SCAN_IN;
  assign n11231 = ~n11227 & ~P1_IR_REG_28__SCAN_IN;
  assign n10803 = ~n10763 | ~n10762;
  assign n10763 = ~n9341 | ~n9156;
  assign n10716 = ~n9194 | ~n10671;
  assign n9194 = ~n9920 | ~n10660;
  assign n12346 = ~n11182 ^ P1_IR_REG_25__SCAN_IN;
  assign n10629 = n10649 | n10618;
  assign n11194 = ~P1_IR_REG_22__SCAN_IN;
  assign n11195 = ~n11193 | ~P1_IR_REG_31__SCAN_IN;
  assign n16922 = n16872;
  assign n16794 = ~n16772 | ~n16773;
  assign n15421 = ~n15442;
  assign n16426 = n12412 | n12411;
  assign n15686 = ~n9191 & ~n15670;
  assign n16241 = n11907 & n12073;
  assign n17638 = ~n17640 & ~n12384;
  assign n17630 = ~n17632 & ~n12386;
  assign n9497 = ~n12834 | ~n12835;
  assign n9410 = n12876 & n12885;
  assign n9411 = n12890 & n9413;
  assign n10865 = ~n10850 | ~n10849;
  assign n9728 = ~n12907;
  assign n10888 = n17041 | n11063;
  assign n12974 = ~n12973 & ~n12972;
  assign n9332 = n9503 & n9333;
  assign n9472 = n11100 & n17117;
  assign n9735 = ~n9736 & ~n13001;
  assign n9736 = ~n12993;
  assign n9509 = n16934 & n9510;
  assign n9726 = ~n10974;
  assign n9469 = ~n9723 | ~n9039;
  assign n9723 = n9724 & n10977;
  assign n9365 = ~n12808 | ~n12805;
  assign n9362 = ~n9364 & ~n9363;
  assign n9363 = ~n12933 | ~n12810;
  assign n12726 = n13021 & n13010;
  assign n13049 = ~n9229 | ~n13042;
  assign n9229 = ~n11785 | ~n9230;
  assign n9230 = ~n13003 & ~n9231;
  assign n9707 = ~n9018 | ~n10998;
  assign n13161 = ~n9367 | ~n9366;
  assign n9366 = ~n12767;
  assign n9368 = ~n12766;
  assign n9530 = ~n15840 & ~n12803;
  assign n9521 = n9527 & n13058;
  assign n9511 = ~n13801 | ~n9512;
  assign n9937 = ~n10932;
  assign n13068 = n15035 | n8987;
  assign n9406 = ~n13031 | ~n9407;
  assign n9741 = n13044 & n13036;
  assign n11073 = ~n11072;
  assign n11072 = n13506 | n13273;
  assign n9324 = ~n11054;
  assign n9718 = ~n11036;
  assign n9330 = n11026 & n9331;
  assign n9326 = n9327 & n11059;
  assign n9936 = ~n10352 & ~n9937;
  assign n9981 = ~P2_IR_REG_15__SCAN_IN & ~P2_IR_REG_9__SCAN_IN;
  assign n9982 = ~P2_IR_REG_14__SCAN_IN & ~P2_IR_REG_12__SCAN_IN;
  assign n9983 = ~P2_IR_REG_11__SCAN_IN & ~P2_IR_REG_8__SCAN_IN;
  assign n9536 = ~n9537 | ~n12813;
  assign n9537 = ~n9538 & ~n14883;
  assign n9538 = ~n9539 | ~n14835;
  assign n12811 = ~n9531 & ~n12807;
  assign n9531 = ~n9535 | ~n9532;
  assign n9524 = ~n13064 | ~n9742;
  assign n9897 = ~n9898 | ~n12793;
  assign n9898 = ~n13174;
  assign n9896 = ~n12229 | ~n12736;
  assign n9417 = ~n13143 & ~n9418;
  assign n10719 = n10746 & n10713;
  assign n11167 = ~P1_IR_REG_22__SCAN_IN & ~P1_IR_REG_21__SCAN_IN;
  assign n9665 = ~n9089;
  assign n11158 = ~P1_IR_REG_7__SCAN_IN;
  assign n11159 = ~P1_IR_REG_8__SCAN_IN;
  assign n10015 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n9241 = ~n9052 | ~n13445;
  assign n9489 = n9846 & n12469;
  assign n9633 = n16475 & n9634;
  assign n9634 = n9635 | n16431;
  assign n9832 = ~n16551;
  assign n9338 = ~n11073 & ~n10828;
  assign n9946 = ~n9014 | ~n11068;
  assign n9944 = ~n10810 & ~n9945;
  assign n9945 = ~n9014;
  assign n9513 = n13250 & n13631;
  assign n11114 = ~n9209 & ~n9085;
  assign n9200 = n9201 & n9026;
  assign n9201 = ~n9917 | ~n9106;
  assign n9551 = n9552 & n11089;
  assign n11090 = n13984 | n13251;
  assign n9309 = ~n9310 | ~n9549;
  assign n13678 = ~n9549 | ~n9548;
  assign n9929 = n9930 & n10561;
  assign n9931 = ~n11111;
  assign n9575 = ~n13227;
  assign n13895 = ~n9953 | ~n9952;
  assign n9299 = ~n9300 | ~n10127;
  assign n10518 = n10516 & n10515;
  assign n9447 = ~n14463;
  assign n9443 = ~n14327;
  assign n9446 = n14464 & n9447;
  assign n9451 = ~n9767 | ~n9452;
  assign n9452 = ~n14358;
  assign n9623 = ~n9016;
  assign n9732 = n13078 & n9015;
  assign n9423 = ~n14789;
  assign n9393 = n9876 & n12905;
  assign n9874 = ~n12655;
  assign n15918 = ~n15972 & ~n16283;
  assign n9383 = ~n16083;
  assign n9729 = n9502 & n16087;
  assign n9856 = ~n12681;
  assign n9852 = ~n9857 & ~n9853;
  assign n9853 = ~n12679;
  assign n14605 = n15059 | n14608;
  assign n13175 = ~n15059 | ~n14608;
  assign n9682 = ~n9683;
  assign n9588 = ~n9869;
  assign n9887 = n14856 | n12766;
  assign n9867 = ~n12661;
  assign n9690 = ~n9691;
  assign n12661 = ~n15177 | ~n14535;
  assign n9605 = ~n12756 & ~n9606;
  assign n9606 = ~n12959;
  assign n9394 = ~n9595 | ~n9594;
  assign n9594 = n9881 & n12244;
  assign n9881 = ~n12652;
  assign n9883 = ~n12223 | ~n12810;
  assign n9889 = n9890 & n12804;
  assign n9891 = ~n12895;
  assign n15893 = ~n15891;
  assign n15896 = ~n15894 | ~n15893;
  assign n10717 = n10728 & n10719;
  assign n10694 = n10692 & n10691;
  assign n11203 = ~P1_IR_REG_20__SCAN_IN;
  assign n10434 = n10432 & n10431;
  assign n9912 = n10355 & n10323;
  assign n10328 = n10326 & n10325;
  assign n10241 = ~SI_9_;
  assign n9842 = ~n13472;
  assign n12515 = ~n14071 ^ n12524;
  assign n10702 = n10683 & P2_REG3_REG_25__SCAN_IN;
  assign n9247 = ~n9248 | ~n12123;
  assign n13505 = n13615 & n9136;
  assign n13569 = ~n13615 | ~n9750;
  assign n10664 = n10635 & P2_REG3_REG_23__SCAN_IN;
  assign n10635 = n10622 & P2_REG3_REG_22__SCAN_IN;
  assign n9762 = ~n9763;
  assign n10622 = n10595 & P2_REG3_REG_21__SCAN_IN;
  assign n10595 = n10569 & P2_REG3_REG_20__SCAN_IN;
  assign n10569 = n10552 & P2_REG3_REG_19__SCAN_IN;
  assign n9757 = ~n14125 | ~n9758;
  assign n9758 = ~n17505;
  assign n10447 = n10393 | n10392;
  assign n17008 = ~n17039 & ~n17041;
  assign n9271 = ~n17077 | ~n9047;
  assign n9805 = ~n17067 ^ n16516;
  assign n17074 = n17096 & n17419;
  assign n9276 = n9277 & n13212;
  assign n9279 = ~n17143 | ~n9051;
  assign n13207 = n13204 & n13203;
  assign n13287 = ~n17224 & ~n12568;
  assign n9814 = ~n13256;
  assign n13253 = ~n9958 | ~n13252;
  assign n13588 = ~n13610 | ~n11032;
  assign n9283 = ~n9090 | ~n9219;
  assign n9218 = n9809 & n13680;
  assign n9811 = n9947 & n13243;
  assign n13631 = ~n13246;
  assign n9947 = ~n11014 | ~n11015;
  assign n13244 = ~n9220 | ~n9219;
  assign n9220 = n9579 & n13680;
  assign n9213 = n13827 & n13833;
  assign n9212 = n11093 & n13835;
  assign n9753 = ~n9755 & ~n14102;
  assign n9754 = ~n16943;
  assign n9819 = n13226 & n13225;
  assign n17096 = ~n17134 & ~n17409;
  assign n16489 = ~n16463;
  assign n17373 = n10822;
  assign n10817 = ~n9323;
  assign n10543 = n10541 & n10540;
  assign n9674 = n9675 & n10513;
  assign n9675 = ~n10537;
  assign n9321 = ~n10521 | ~n9322;
  assign n10522 = ~n10467 & ~P2_IR_REG_17__SCAN_IN;
  assign n10386 = n10385 | P2_IR_REG_13__SCAN_IN;
  assign n9775 = ~n11371;
  assign n9772 = ~n15396;
  assign n9767 = ~n14374 & ~n9768;
  assign n9768 = ~n14359;
  assign n9445 = n14464 | n9447;
  assign n9444 = ~n11768 | ~n9442;
  assign n9442 = ~n9446 & ~n9443;
  assign n15392 = ~n15394 | ~n15395;
  assign n14411 = ~n8997 | ~n15331;
  assign n11270 = n11924 | n16244;
  assign n9785 = ~n9022 | ~n11724;
  assign n14289 = ~n9789 | ~n9790;
  assign n9790 = ~n9788;
  assign n11631 = ~n11620 | ~n11619;
  assign n9544 = ~n13122 & ~n9545;
  assign n9545 = ~n9037 | ~n14567;
  assign n12820 = ~n12819 & ~n9540;
  assign n15792 = ~n9184 | ~n15782;
  assign n11855 = n11828 & P1_REG3_REG_25__SCAN_IN;
  assign n9176 = n9610 & n13167;
  assign n9610 = ~n9612 | ~n9902;
  assign n14713 = ~n9476 | ~n9678;
  assign n9678 = ~n9681 & ~n15091;
  assign n11733 = n11713 & P1_REG3_REG_19__SCAN_IN;
  assign n14792 = ~n14790 & ~n15123;
  assign n11666 = n11608 | n11224;
  assign n15969 = n13148 & n12235;
  assign n16025 = n13102 | n12251;
  assign n9599 = ~n14567 & ~n9600;
  assign n9600 = ~n12683;
  assign n12650 = ~n9427 | ~n9614;
  assign n9614 = n9615 & n12649;
  assign n9386 = n9388 & n9860;
  assign n9863 = ~n12675 & ~n9864;
  assign n9864 = ~n12673;
  assign n14660 = n13169 & n13171;
  assign n14681 = ~n9900 | ~n12796;
  assign n9900 = ~n12647 | ~n9901;
  assign n9683 = ~n14762 | ~n9684;
  assign n14790 = ~n9476;
  assign n14735 = ~n9680 | ~n9679;
  assign n9680 = ~n9681;
  assign n9679 = ~n14790;
  assign n14749 = n12646 & n12727;
  assign n14871 = ~n14977 & ~n9685;
  assign n9685 = ~n9690 | ~n9686;
  assign n9686 = ~n15166 & ~n15155;
  assign n9688 = ~n9690 | ~n9689;
  assign n9608 = ~n14933 | ~n12959;
  assign n14992 = n9394 & n12905;
  assign n9492 = ~n15003 & ~n15209;
  assign n12245 = ~n9595 | ~n12244;
  assign n12406 = n15874 & n12269;
  assign n12652 = n12805 & n12223;
  assign n15956 = n15954 & n15961;
  assign n16296 = ~n11358 | ~n11357;
  assign n16020 = ~n12231 | ~n12230;
  assign n16055 = ~n16074;
  assign n11212 = ~P1_IR_REG_28__SCAN_IN;
  assign n11205 = ~P1_IR_REG_25__SCAN_IN;
  assign n10657 = n10655 & n10654;
  assign n10610 = n10608 & n10607;
  assign n10582 = n10580 & n10579;
  assign n11199 = ~P1_IR_REG_21__SCAN_IN;
  assign n10460 = ~n9670 | ~n9115;
  assign n11592 = n11576 | P1_IR_REG_13__SCAN_IN;
  assign n10270 = ~SI_10_;
  assign n11472 = n11445 | P1_IR_REG_8__SCAN_IN;
  assign n9560 = n10238 & n9558;
  assign n11382 = n11353 | P1_IR_REG_4__SCAN_IN;
  assign n10147 = ~n9746 | ~n10732;
  assign n9480 = ~n12610;
  assign n16628 = n13314;
  assign n9637 = ~n16583;
  assign n9645 = ~n16585;
  assign n16501 = n12491 | n12490;
  assign n16583 = n12483 | n12484;
  assign n9174 = ~n16486;
  assign n16608 = ~n16631;
  assign n17432 = ~n9656 | ~n10172;
  assign n9656 = n17312 | n10698;
  assign n13494 = ~n16608 & ~n16604;
  assign n13495 = ~n13448;
  assign n9345 = ~n11123 & ~n9955;
  assign n9205 = ~n9709 | ~n9708;
  assign n9348 = ~n9313 & ~n11084;
  assign n13806 = n10453 & n10452;
  assign n12005 = n10400 & n10399;
  assign n13898 = n10376 & n10375;
  assign n10921 = n10318 & n10317;
  assign n12026 = n10198 & n10197;
  assign n9954 = n10777 & P2_REG1_REG_2__SCAN_IN;
  assign n16655 = ~n9267 | ~n12114;
  assign n9251 = ~n12123 & ~n9254;
  assign n10334 = n10248 & n10247;
  assign n9256 = n9257 & n16745;
  assign n13531 = ~n13280;
  assign n9581 = ~n9088 | ~n9582;
  assign n9583 = ~n13239;
  assign n13713 = ~n13757 & ~n9763;
  assign n9233 = ~n16124 | ~n10732;
  assign n13926 = ~n16943 & ~n17505;
  assign n10312 = n10281 & P2_REG3_REG_9__SCAN_IN;
  assign n17362 = ~n17212;
  assign n17081 = ~n9805;
  assign n17134 = ~n9748 | ~n17141;
  assign n9748 = ~n17142;
  assign n9298 = ~n16490 | ~n16568;
  assign n12571 = ~P2_D_REG_1__SCAN_IN & ~n17224;
  assign n13953 = ~n13506;
  assign n13986 = n9023 | n13595;
  assign n13701 = n9799 & n13240;
  assign n9799 = n13725 | n13727;
  assign n9807 = ~n9216;
  assign n14107 = n13877 & n13876;
  assign n9290 = ~n9296 | ~n9294;
  assign n16929 = ~n16961 | ~n13225;
  assign n16983 = ~n9275 | ~n13222;
  assign n10191 = n17305 | n10698;
  assign n17224 = ~n17351 | ~n12573;
  assign n9699 = ~n11133 & ~P2_IR_REG_28__SCAN_IN;
  assign n11143 = n11133 | n11134;
  assign n10824 = ~n10819 ^ n10818;
  assign n10818 = ~P2_IR_REG_22__SCAN_IN;
  assign n10819 = ~n11124 | ~P2_IR_REG_31__SCAN_IN;
  assign n10811 = ~P2_IR_REG_19__SCAN_IN;
  assign n17334 = n10098 & n10097;
  assign n14586 = ~n16410;
  assign n14237 = ~n11868 & ~n11867;
  assign n14269 = n11814 & n11813;
  assign n15348 = ~n9430 | ~n9515;
  assign n14320 = n11729 | n11728;
  assign n9429 = ~n11522 | ~n11521;
  assign n14375 = n11680 | n11679;
  assign n14378 = ~n9769 | ~n14359;
  assign n15412 = ~n9437 | ~n9017;
  assign n9487 = n16087;
  assign n15188 = ~n11548 | ~n11547;
  assign n14470 = ~P1_REG3_REG_22__SCAN_IN;
  assign n15134 = ~n11707 | ~n11706;
  assign n15429 = n11948 & n12251;
  assign n12792 = n9349 & n13124;
  assign n9400 = ~n9507 & ~n13102;
  assign n14751 = n11753 & n11752;
  assign n13011 = n11740 & n11739;
  assign n14828 = n11717 & n11716;
  assign n14804 = n11673 & n11672;
  assign n14364 = n11615 & n11614;
  assign n14937 = n11587 & n11586;
  assign n14965 = n11558 & n11557;
  assign n14993 = n11535 & n11534;
  assign n14964 = n11490 & n11489;
  assign n15847 = n9373 & n11507;
  assign n9373 = n9374 & n11502;
  assign n9374 = ~n11286 | ~P1_REG1_REG_10__SCAN_IN;
  assign n12908 = n11460 & n11459;
  assign n15848 = n11437 & n11436;
  assign n15437 = n11415 & n11414;
  assign n15326 = n11380 & n11379;
  assign n9404 = ~n8988 | ~P1_REG2_REG_2__SCAN_IN;
  assign n11247 = ~n11289 | ~P1_REG2_REG_1__SCAN_IN;
  assign n9179 = ~n9177 | ~n15530;
  assign n9177 = ~n15506;
  assign n9182 = ~n12090;
  assign n15748 = n9187 & n9161;
  assign n9187 = ~n9189 | ~n9188;
  assign n9188 = ~n15718;
  assign n9693 = ~n13082;
  assign n9694 = ~n9696;
  assign n15034 = ~n14596 ^ n9697;
  assign n9880 = ~n8998 & ~n9044;
  assign n14296 = ~n9372 | ~n11501;
  assign n9372 = n17284 | n12401;
  assign n11504 = ~n11454 & ~n11221;
  assign n9385 = ~n15864;
  assign n12237 = ~n15890 | ~n15891;
  assign n15926 = ~n9384;
  assign n9473 = ~n16039 & ~n16274;
  assign n16108 = ~n15996;
  assign n12400 = n14195 | n12401;
  assign n14594 = ~n9854 | ~n12682;
  assign n15065 = ~n14638 & ~n14637;
  assign n14689 = ~n12674 | ~n12673;
  assign n9592 = ~n12659;
  assign n16261 = n11294 & n11293;
  assign n9677 = n12402 | n11250;
  assign n9517 = n9520 & n9519;
  assign n11172 = ~P1_IR_REG_23__SCAN_IN;
  assign n9354 = n11230 & n15277;
  assign n10760 = ~n9341 | ~n9342;
  assign n9170 = n10731 & n10730;
  assign n9464 = n10651 | n9154;
  assign n15319 = ~n11184 ^ P1_IR_REG_24__SCAN_IN;
  assign n9206 = ~n10604;
  assign n11190 = n11189 & n11188;
  assign n11188 = ~P1_IR_REG_18__SCAN_IN;
  assign n17245 = ~n10460 ^ n10458;
  assign n9913 = ~n10382 | ~n9914;
  assign n17265 = ~n10380 ^ n10378;
  assign n17284 = ~n10295 ^ n10293;
  assign n10210 = ~n10203 | ~n10235;
  assign n10203 = n10202 | n10201;
  assign n17305 = ~n10202 ^ n10200;
  assign n15489 = ~n9193 ^ n9192;
  assign n16226 = n11257 & n11256;
  assign n16569 = ~n16617;
  assign n13344 = ~n9378 | ~n9381;
  assign n9378 = ~n9458 & ~n9041;
  assign n9824 = n9825 & n9049;
  assign n9826 = ~n9827;
  assign n13392 = ~n12511;
  assign n13393 = ~n9494 | ~n12510;
  assign n13419 = ~n9493 | ~n13345;
  assign n16617 = n12583 & n17209;
  assign n9479 = ~n12608;
  assign n16575 = n12597 & n12578;
  assign n17585 = n10744 | n10743;
  assign n17561 = n10559 | n10558;
  assign n13395 = n10505 | n10504;
  assign n13838 = n10485 | n10484;
  assign n13871 = ~n13806;
  assign n13935 = ~n12005;
  assign n16506 = ~n13898;
  assign n16592 = n10351 | n10350;
  assign n16505 = ~n10921;
  assign n16559 = n10287 | n10286;
  assign n16477 = n10262 | n10261;
  assign n16558 = n10227 | n10226;
  assign n16627 = ~n12026;
  assign n17342 = n9262 & n10032;
  assign n16913 = ~n12105 | ~n12104;
  assign n16811 = ~n9263 & ~n16795;
  assign n16868 = ~n9269 | ~n16849;
  assign n9264 = ~n9266 ^ n9265;
  assign n17209 = ~n17225 | ~n12582;
  assign n12582 = ~n13290;
  assign n17130 = ~n17087 | ~n17176;
  assign n17553 = ~n13949 | ~n13948;
  assign n17555 = ~n17553;
  assign n14175 = n14097 | n14096;
  assign n17501 = ~n13291 | ~n13949;
  assign n13291 = ~n13948;
  assign n17514 = ~n17501;
  assign n17358 = ~n11187;
  assign n17352 = ~n11132 ^ P2_IR_REG_24__SCAN_IN;
  assign n11132 = ~n11131 | ~P2_IR_REG_31__SCAN_IN;
  assign n17351 = ~n14220;
  assign n9991 = ~P2_IR_REG_30__SCAN_IN;
  assign n12569 = ~n11145 ^ n11144;
  assign n11145 = ~n11143 | ~P2_IR_REG_31__SCAN_IN;
  assign n10782 = ~n9323 | ~P2_IR_REG_31__SCAN_IN;
  assign n9793 = ~n9072 | ~n11930;
  assign n9795 = n9457 & n9454;
  assign n9454 = n9455 & n9094;
  assign n14329 = ~n14325 & ~n14324;
  assign n14843 = ~n15145;
  assign n14466 = ~n11768 | ~n14327;
  assign n15457 = n11943 & n11909;
  assign n13198 = n13196 | n13195;
  assign n13120 = ~n13110 | ~n9486;
  assign n9486 = ~n13119 & ~n13192;
  assign n16419 = n11956 | n11955;
  assign n16416 = n11919 | n11918;
  assign n16413 = n11860 | n11859;
  assign n14703 = ~n14751;
  assign n14774 = ~n13011;
  assign n14859 = ~n14804;
  assign n14533 = n11647 | n11646;
  assign n14908 = ~n14364;
  assign n14907 = ~n14965;
  assign n15903 = ~n15848;
  assign n15929 = ~n15437;
  assign n15585 = ~n15582 | ~n15581;
  assign n9190 = n15686 | n15685;
  assign n16011 = n16337 | n11933;
  assign n16003 = n16104 | n16095;
  assign n16109 = ~n16040;
  assign n16119 = ~n16104;
  assign n16393 = ~n12295 | ~n12294;
  assign n16395 = ~n16393;
  assign n12419 = n12416 | n12415;
  assign n12700 = ~n12699 & ~n12698;
  assign n16349 = ~n12295 | ~n12291;
  assign n16363 = ~n16349;
  assign n16239 = ~n11906 | ~n11905;
  assign n16234 = n15310 | n15319;
  assign n16233 = ~n16123 | ~n16241;
  assign n15276 = ~n11231 | ~n11230;
  assign n15275 = ~n9019 | ~n10798;
  assign n15309 = ~n10680 | ~n10726;
  assign n12334 = ~n10619 | ~n10629;
  assign n16128 = ~n12395 | ~P1_U3084;
  assign n16225 = ~n15317;
  assign n15502 = P1_IR_REG_0__SCAN_IN;
  assign n17646 = ~n17648 & ~n12382;
  assign n17634 = ~n17636 & ~n12385;
  assign n17626 = ~n17628 & ~n12387;
  assign n9563 = n13540 & n9102;
  assign n9508 = ~n9081 | ~n9000;
  assign n8997 = n15333 | n9441;
  assign n8998 = ~n12667 & ~n14786;
  assign n11077 = n13945 | n17595;
  assign n11093 = ~n14102 | ~n13897;
  assign n8999 = n9110 & n9390;
  assign n9000 = ~n9782 | ~n9780;
  assign n9001 = n11069 | n11063;
  assign n9002 = n9035 & n12975;
  assign n9003 = n9451 & n14375;
  assign n9004 = n12487 & n13838;
  assign n9005 = n11119 & n17227;
  assign n9006 = n11093 & n9952;
  assign n9007 = n9889 & n9101;
  assign n9008 = n13944 | n12581;
  assign n9009 = n10872 | n10871;
  assign n11008 = ~n13690;
  assign n9010 = n9096 & n12793;
  assign n9173 = ~n10101;
  assign n9011 = n9190 & n9151;
  assign n13837 = ~n13897;
  assign n13897 = n10427 & n10426;
  assign n9012 = n9841 & n9842;
  assign n9577 = ~n13933;
  assign n12902 = n13107 & n16090;
  assign n9765 = ~n14049;
  assign n9013 = ~n9155 & ~n12736;
  assign n17087 = ~n13511 | ~n17209;
  assign n9014 = n10784 & n10783;
  assign n9015 = n13084 | n13083;
  assign n9016 = n13089 & n13088;
  assign n12800 = n13134 & n12829;
  assign n9017 = n11274 & n11275;
  assign n9018 = n10995 | n10994;
  assign n9019 = n10804 & n10797;
  assign n9020 = n10809 & n11074;
  assign n13813 = n9460 & n10475;
  assign n9021 = ~n11422 | ~n11421;
  assign n15958 = ~n15326;
  assign n9022 = n11730 & n14320;
  assign n9364 = ~n12955;
  assign n9023 = n13615 & n9752;
  assign n9024 = n12511 & n12510;
  assign n9025 = ~n17313 & ~P2_REG2_REG_6__SCAN_IN;
  assign n9026 = n11071 | n11070;
  assign n9027 = n9654 & n13358;
  assign n9028 = n16960 & n9293;
  assign n9029 = n12627 | n12626;
  assign n9030 = n15865 & n15869;
  assign n9031 = n13081 & n13080;
  assign n9032 = n10974 & n10964;
  assign n9033 = n13010 & n12727;
  assign n9034 = n11076 | n11075;
  assign n9035 = ~n15155 | ~n14885;
  assign n17582 = n10706 | n10705;
  assign n9036 = n9034 & n9337;
  assign n10428 = n10430 & n10410;
  assign n9572 = ~n16963;
  assign n9037 = n13126 ^ n13125;
  assign n9038 = n13750 | n13775;
  assign n10523 = ~P2_IR_REG_31__SCAN_IN;
  assign n9039 = n10983 | n10982;
  assign n9040 = n9840 & n9843;
  assign n14905 = ~n9608 | ~n12955;
  assign n14701 = ~n12647 | ~n13021;
  assign n13559 = n9550 & n9551;
  assign n13774 = n13803 & n10487;
  assign n9041 = ~n12517 & ~n12516;
  assign n9042 = n9576 & n13227;
  assign n9043 = n11232 & P1_REG2_REG_0__SCAN_IN;
  assign n9044 = n15123 & n14509;
  assign n13583 = ~n9283 | ~n9286;
  assign n9045 = n12664 & n12814;
  assign n9046 = n11104 & n17015;
  assign n13933 = ~n13920 ^ n13898;
  assign n9047 = n9804 & n17058;
  assign n13964 = ~n10735 | ~n10734;
  assign n9749 = ~n13964;
  assign n9048 = n10985 | n10984;
  assign n9049 = n12628 | n16575;
  assign n9050 = n12692 | n12691;
  assign n9051 = n13211 & n17148;
  assign n9052 = n13690 ^ n12624;
  assign n13680 = ~n10999 | ~n11000;
  assign n9053 = n9033 & n9422;
  assign n9054 = n15040 & n14643;
  assign n9055 = n10046 & n17387;
  assign n9056 = n11068 | n10828;
  assign n9057 = n9236 & n9244;
  assign n13107 = ~n11195 ^ n11194;
  assign n9058 = ~n13189 & ~n13108;
  assign n13679 = ~n9549 | ~n10578;
  assign n9059 = n17476 ^ n16559;
  assign n9510 = ~n9059;
  assign n14799 = ~n9887 | ~n9002;
  assign n9060 = ~n14603 & ~n9054;
  assign n9061 = ~n11849 & ~n9779;
  assign n9062 = n11123 & n10821;
  assign n12737 = n15972 & n16283;
  assign n9063 = n11802 & P1_REG0_REG_2__SCAN_IN;
  assign n9064 = n10456 & n10455;
  assign n9065 = n11030 & n11029;
  assign n9066 = n13123 | n13085;
  assign n9067 = n9223 & n9224;
  assign n9068 = n9195 & n11062;
  assign n9069 = n9715 & n11044;
  assign n9070 = n9734 & n13000;
  assign n9071 = n11119 | n11118;
  assign n9072 = n14235 & n15457;
  assign n9073 = n11116 & n13557;
  assign n9074 = n9769 & n9767;
  assign n9075 = n11121 & n9071;
  assign n13622 = ~n13995;
  assign n9076 = n10859 | n10858;
  assign n9077 = n14361 | n9453;
  assign n13572 = ~n13974;
  assign n9078 = n12974 & n9399;
  assign n13892 = ~n9546 | ~n10377;
  assign n9079 = n12802 & n15969;
  assign n9080 = n12881 & n12880;
  assign n9081 = n9514 & n15457;
  assign n9082 = n9947 | n9948;
  assign n9083 = n9701 & n9700;
  assign n11230 = ~P1_IR_REG_29__SCAN_IN;
  assign n9084 = n13058 | n9527;
  assign n9085 = n13606 | n9465;
  assign n9697 = ~n15035;
  assign n13920 = ~n9567 | ~n10368;
  assign n9086 = n17582 & n10699;
  assign n9760 = ~n9761;
  assign n9761 = ~n13714 | ~n9762;
  assign n9087 = n9320 & n10780;
  assign n9088 = n9796 & n13242;
  assign n9407 = ~n13028;
  assign n9089 = n10488 ^ SI_17_;
  assign n9901 = ~n9902;
  assign n9902 = n12725 | n9903;
  assign n11228 = ~P1_IR_REG_31__SCAN_IN;
  assign n9350 = ~n13189;
  assign n9090 = n9579 & n9218;
  assign n13714 = ~n14038;
  assign n15277 = ~P1_IR_REG_30__SCAN_IN;
  assign n9091 = n13149 & n13148;
  assign n12759 = ~n15847 & ~n14296;
  assign n9092 = n9906 & n10562;
  assign n9093 = n11072 & n11074;
  assign n9094 = n11932 & n15457;
  assign n9095 = ~n11286 | ~P1_REG1_REG_0__SCAN_IN;
  assign n17588 = n10759 | n10758;
  assign n9918 = ~n17588;
  assign n9797 = ~n9798;
  assign n9798 = ~n13241 | ~n13240;
  assign n9096 = n13171 & n13175;
  assign n9097 = n11249 | n16251;
  assign n9098 = n10937 & n10936;
  assign n9099 = n9882 & n12933;
  assign n9100 = n13757 | n14060;
  assign n9101 = n12753 & n12805;
  assign n9102 = n13536 & n13535;
  assign n14464 = ~n11781 ^ n11811;
  assign n9103 = n10965 & n9722;
  assign n9104 = n10993 & n10992;
  assign n9105 = n10864 & n10865;
  assign n9414 = ~n15286;
  assign n16244 = n11267 & n11266;
  assign n16087 = ~n16244;
  assign n9106 = n11067 & n11066;
  assign n13608 = ~n13606;
  assign n9107 = n12788 & n13174;
  assign n9108 = n13221 & n13220;
  assign n9109 = n12465 & n16523;
  assign n10091 = ~P2_IR_REG_1__SCAN_IN & ~P2_IR_REG_0__SCAN_IN;
  assign n9262 = ~n10091;
  assign n14922 = ~n9687;
  assign n9687 = ~n14977 & ~n9691;
  assign n9110 = n12676 & n12672;
  assign n9111 = n10879 & n10878;
  assign n9112 = n15584 & n9185;
  assign n9113 = ~n10987 | ~n10986;
  assign n9114 = ~n16516 & ~n17432;
  assign n9115 = n9671 & n10430;
  assign n9116 = n9581 | n9578;
  assign n9117 = n10428 & n10404;
  assign n9118 = n13235 & n13229;
  assign n9119 = n9674 & n10548;
  assign n9120 = ~n14071 | ~n13395;
  assign n9121 = n13101 & n13100;
  assign n9122 = n11081 & n9093;
  assign n9192 = ~P1_IR_REG_2__SCAN_IN;
  assign n9123 = n13552 & n13551;
  assign n9124 = n9607 | n12756;
  assign n9125 = n13248 & n9809;
  assign n9126 = n13947 & n13946;
  assign n9127 = n12935 & n12934;
  assign n9128 = n11048 & n11047;
  assign n9129 = n9839 & n9964;
  assign n9130 = n13040 & n13039;
  assign n9131 = n9092 & n9206;
  assign n9132 = n11017 & n11016;
  assign n9462 = ~n9235;
  assign n9235 = ~n9651 | ~n12528;
  assign n9133 = ~n9665 & ~n9664;
  assign n10004 = ~P2_IR_REG_28__SCAN_IN;
  assign n9134 = n9616 & n9855;
  assign n9135 = n13244 & n13243;
  assign n9136 = n9750 & n9749;
  assign n9137 = n12899 & n9728;
  assign n9138 = n12621 & n9029;
  assign n9139 = n9887 & n9035;
  assign n9140 = n9695 & n9693;
  assign n9141 = n9702 & n10945;
  assign n9142 = n9659 & n9912;
  assign n9143 = ~n13757 & ~n9761;
  assign n9144 = n9896 & n12742;
  assign n9843 = ~n12615;
  assign n9145 = n11050 & n11088;
  assign n9146 = n9408 & n13024;
  assign n9147 = n14977 | n9688;
  assign n9148 = ~n9522 | ~n13058;
  assign n9149 = ~n9031 | ~n13078;
  assign n9500 = n12791;
  assign n11082 = n10824 & n12424;
  assign n9689 = ~n15166;
  assign n17028 = ~n9568 | ~n9800;
  assign n9684 = ~n15123;
  assign n9150 = n10761 | SI_29_;
  assign n13932 = ~n9935 | ~n10932;
  assign n17009 = ~n17028 | ~n13220;
  assign n13432 = ~n9822 | ~n16501;
  assign n13835 = n13232 & n11092;
  assign n9512 = ~n13835;
  assign n9151 = n16173 | P1_REG1_REG_11__SCAN_IN;
  assign n9764 = ~n14060;
  assign n9698 = ~n15025;
  assign n9152 = n17087 | P2_REG2_REG_29__SCAN_IN;
  assign n13142 = n16261 | n16076;
  assign n9153 = ~n10488 | ~SI_17_;
  assign n9322 = ~P2_IR_REG_17__SCAN_IN;
  assign n9154 = n10653 & SI_24_;
  assign n9155 = n16053 & n9417;
  assign n9156 = n9342 & n9150;
  assign n9157 = n14528 & n14527;
  assign n9158 = n9889 & n12805;
  assign n9159 = n16943 | n9755;
  assign n15925 = ~n12868 | ~n13149;
  assign n16076 = ~n9484 | ~n9404;
  assign n10825 = n10824;
  assign n9160 = ~n15494 & ~P1_U3084;
  assign n13192 = n11243;
  assign n9161 = n16161 | P1_REG1_REG_13__SCAN_IN;
  assign n16088 = ~n16251;
  assign n9162 = n9252 | n9251;
  assign n17098 = ~n17227;
  assign n13537 = n12422;
  assign n16924 = ~n9264 | ~n16921;
  assign n9657 = ~n10083 | ~n10084;
  assign n9291 = ~n9289 | ~n13893;
  assign n10159 = ~n10143 | ~n10142;
  assign n10267 = ~n9905 | ~n10265;
  assign n9292 = ~n9294;
  assign n9573 = ~n9819;
  assign n13629 = n9810 & n13245;
  assign n13237 = ~n9217 | ~n9215;
  assign n9460 = ~n9459 | ~n10732;
  assign n9237 = ~n9243 | ~n9242;
  assign n12967 = ~n9163 | ~n12958;
  assign n9163 = ~n12957 | ~n12956;
  assign n12984 = ~n9164 | ~n12978;
  assign n9164 = ~n9078 | ~n9397;
  assign n9658 = ~n10054;
  assign P2_U3268 = n13553 | n9169;
  assign n9490 = ~n10295;
  assign n10663 = ~n12345 | ~n10732;
  assign n9552 = ~n9553 | ~n13606;
  assign n11155 = ~n9165 | ~n11126;
  assign n9165 = ~n9346 | ~n9172;
  assign n12345 = ~n9194 | ~n10661;
  assign n9527 = ~n13055;
  assign n9341 = ~n10716 | ~n10715;
  assign n9226 = ~n9228 | ~n9227;
  assign n12703 = ~n12706 | ~n12700;
  assign n14213 = ~n10697 ^ n10707;
  assign n9616 = ~n13180;
  assign n10013 = ~P2_RD_REG_SCAN_IN;
  assign n13168 = ~n9166 | ~n13166;
  assign n9166 = ~n13132;
  assign n13132 = ~n12782 | ~n12783;
  assign n9282 = ~n13244;
  assign n13179 = ~n9167 | ~n13178;
  assign n9167 = ~n13173 | ~n13174;
  assign n13190 = ~n9168 | ~n13188;
  assign n9168 = ~n13186 | ~n13187;
  assign n9169 = ~n13556 | ~n9123;
  assign n13630 = ~n9309 | ~n9308;
  assign n14208 = ~n9170 | ~n10747;
  assign n13106 = ~n12828 & ~n16090;
  assign n13121 = ~n13106 & ~n13105;
  assign n12532 = ~n9171 | ~n9237;
  assign n11123 = ~n9943 | ~n9941;
  assign n13266 = ~n10745 | ~n11087;
  assign n9172 = n9203 & n9204;
  assign n9238 = ~n9239 | ~n9244;
  assign n9377 = ~n9458 & ~n9379;
  assign n13073 = ~n9225 | ~n9067;
  assign n10034 = ~n9173 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n12438 = ~n9175 | ~n9174;
  assign n9175 = ~n16487;
  assign n9601 = ~n9598 | ~n12685;
  assign n15374 = ~n11281 | ~n11280;
  assign n11281 = ~n11277 | ~n11276;
  assign n14503 = n14306 | n14305;
  assign n17039 = n17059 | n17443;
  assign n13615 = ~n13643 & ~n14006;
  assign n11634 = ~n9433 | ~n14530;
  assign n14654 = ~n9176 | ~n9609;
  assign n9676 = n12322 | n12401;
  assign n9613 = ~n9901 | ~n13020;
  assign n9183 = ~n9179;
  assign n15541 = n9183 | n9180;
  assign n15543 = ~n9179 | ~n9178;
  assign n9178 = ~n9180 & ~n15540;
  assign n9180 = ~n9181 | ~n15532;
  assign n15531 = ~n15506 | ~n12090;
  assign n9181 = ~n15530 | ~n9182;
  assign n15794 = ~n15792 | ~n15793;
  assign n9184 = ~n15780 | ~n15781;
  assign n9185 = ~n15563 | ~n15581;
  assign n9186 = ~n15564 | ~n15581;
  assign n15582 = n15564 | n15563;
  assign n15607 = ~n15604 | ~n15603;
  assign n15749 = ~n15748 & ~n15747;
  assign n9189 = ~n15719;
  assign n9191 = ~n15669 & ~n15668;
  assign n9193 = ~n11251 & ~n11228;
  assign n11251 = ~P1_IR_REG_1__SCAN_IN & ~P1_IR_REG_0__SCAN_IN;
  assign n9195 = ~n9326 | ~n9324;
  assign n9197 = ~n9200 | ~n9198;
  assign n9198 = ~n9917;
  assign n9199 = ~n9727 | ~n9200;
  assign n9203 = ~n9345 & ~n9062;
  assign n9204 = ~n9075 | ~n9205;
  assign n10587 = ~n9908 | ~n9131;
  assign n10618 = ~n9207 & ~n10647;
  assign n10652 = ~n9207 & ~n10648;
  assign n12322 = ~n9207 ^ n10604;
  assign n11119 = ~n9073 | ~n9208;
  assign n13832 = ~n13833 | ~n11093;
  assign n13230 = n13827 & n13835;
  assign n13231 = ~n9213 | ~n9212;
  assign n13827 = ~n9214 | ~n13897;
  assign n9214 = ~n14102;
  assign n9506 = ~n9401 | ~n9222;
  assign n13103 = ~n9400 | ~n9222;
  assign n9223 = ~n9525 | ~n9148;
  assign n9224 = ~n9523 | ~n9524;
  assign n9225 = ~n9226 | ~n9466;
  assign n9227 = ~n9525;
  assign n9228 = ~n9523;
  assign n12609 = ~n9232;
  assign n9840 = ~n9232 | ~n9479;
  assign n13405 = ~n9232 ^ n9480;
  assign n9232 = n12533 | n13330;
  assign n9240 = ~n9235 | ~n9241;
  assign n9236 = ~n9462 | ~n9652;
  assign n9239 = ~n9652;
  assign n9375 = ~n9243 & ~n9235;
  assign n9243 = ~n9652 | ~n9052;
  assign n9244 = ~n9052;
  assign n9254 = ~n16694;
  assign n9250 = n16694 | n9245;
  assign n9245 = ~n12124;
  assign n9252 = ~n9246 | ~n12124;
  assign n12127 = ~n9249 | ~n9247;
  assign n9248 = ~n9252;
  assign n16693 = ~n16695 | ~n16694;
  assign n16695 = ~n12123 | ~n12122;
  assign n16746 = ~n9255 | ~n9256;
  assign n9255 = ~n16720 | ~n9259;
  assign n16744 = ~n9258 | ~n12129;
  assign n9258 = ~n16720 | ~n12128;
  assign n10047 = ~n9262 | ~P2_IR_REG_31__SCAN_IN;
  assign n16812 = ~n16811 & ~n16810;
  assign n9263 = ~n16793 & ~n16794;
  assign n12117 = ~n16655 | ~n16656;
  assign n9267 = ~n12184 | ~n12185;
  assign n12185 = ~n12194 ^ n9268;
  assign n16869 = ~n16868 & ~n16867;
  assign n9269 = ~n16848 | ~P2_REG1_REG_15__SCAN_IN;
  assign n16848 = ~n16847 ^ n9270;
  assign n9270 = ~n17253;
  assign n17026 = ~n9800 | ~n9271;
  assign n13725 = ~n9272 | ~n13239;
  assign n9578 = ~n9272 & ~n9798;
  assign n13224 = ~n9275 | ~n9273;
  assign n9280 = ~n17143 | ~n17148;
  assign n17114 = ~n9280 | ~n13210;
  assign n17105 = ~n9279 | ~n9276;
  assign n9277 = ~n13211 | ~n9278;
  assign n13254 = ~n9281 | ~n9284;
  assign n9281 = ~n9282 | ~n9125;
  assign n9810 = ~n13244 | ~n9811;
  assign n9287 = ~n9809 | ~n9288;
  assign n9296 = ~n16960;
  assign n13891 = ~n9290 | ~n9293;
  assign n13293 = ~n9297 | ~n17514;
  assign n13961 = ~n9297 | ~n17555;
  assign n9297 = ~n13284 | ~n13285;
  assign n17161 = ~n9298;
  assign n10061 = ~n12430 | ~n9298;
  assign n17363 = ~n16570 | ~n9298;
  assign n17189 = ~n17198 ^ n9298;
  assign n16574 = ~n16573 | ~n9298;
  assign n9304 = n9966 & n9305;
  assign n10105 = n10064 & n11094;
  assign n9302 = ~n9301 | ~n9299;
  assign n9300 = ~n9305;
  assign n9301 = ~n10106 | ~n10127;
  assign n17147 = ~n10105;
  assign n17091 = ~n9303 | ~n9302;
  assign n9303 = ~n10105 | ~n9304;
  assign n16964 = ~n10319;
  assign n9501 = ~n10319 | ~n9933;
  assign n13800 = n9307 & n10457;
  assign n13803 = ~n9307 | ~n9557;
  assign n9308 = ~n9082 | ~n11015;
  assign n10745 = ~n9311 | ~n9145;
  assign n11085 = ~n9313 | ~n13269;
  assign n9713 = ~n9711 | ~n9314;
  assign n9314 = ~n9315 | ~n9111;
  assign n9315 = ~n9076 | ~n9316;
  assign n9316 = ~n9105 & ~n9009;
  assign n9468 = ~n9317 | ~n9113;
  assign n9317 = ~n9318 | ~n9048;
  assign n9318 = n9103 | n9469;
  assign n10781 = ~n10467 & ~n9321;
  assign n9727 = ~n9325 | ~n9068;
  assign n9325 = ~n11049 | ~n9326;
  assign n9327 = ~n11054 | ~n9128;
  assign n9329 = ~n9706 | ~n9328;
  assign n11031 = ~n9329 | ~n9330;
  assign n9331 = ~n9132 | ~n11021;
  assign n9335 = ~n9334 | ~n9332;
  assign n9333 = ~n10930 | ~n10926;
  assign n9334 = ~n10927 | ~n10930;
  assign n10955 = ~n9335 | ~n9141;
  assign n9516 = ~n9336 | ~n9133;
  assign n9376 = ~n9336 | ~n10461;
  assign n10661 = n9920 | n10660;
  assign n9920 = ~n10652 & ~n9464;
  assign n10747 = n9341 & n9960;
  assign n9346 = ~n9347 | ~n11085;
  assign n9347 = ~n9348 & ~n12580;
  assign n9349 = ~n9351 | ~n9350;
  assign n9351 = ~n9352 | ~n9066;
  assign n9352 = ~n9669 | ~n9667;
  assign n9353 = ~n11231 | ~n9354;
  assign n9360 = n11231 | n9361;
  assign n11286 = n11233 & n15286;
  assign n12761 = ~n9365 | ~n9362;
  assign n12769 = ~n12768 | ~n13161;
  assign n9367 = ~n9369 | ~n9368;
  assign n12789 = ~n9370 | ~n13129;
  assign n9370 = ~n9371 | ~n9107;
  assign n9371 = ~n12787 | ~n12786;
  assign n13446 = ~n9057 & ~n9375;
  assign n17238 = ~n9459;
  assign n9828 = ~n9377 | ~n9381;
  assign n9382 = ~n9097 | ~n9383;
  assign n16299 = ~n9483 ^ n15969;
  assign n15927 = n15926 & n15925;
  assign n15867 = n15926 & n9385;
  assign n12678 = ~n9387 | ~n9386;
  assign n9387 = ~n14731 | ~n8999;
  assign n9388 = ~n8999 | ~n9391;
  assign n14711 = ~n9389 | ~n12671;
  assign n9389 = ~n14731 | ~n14730;
  assign n9391 = ~n12671;
  assign n9593 = ~n12664 | ~n9395;
  assign n9395 = n12665 & n12814;
  assign n12929 = ~n9396 | ~n12924;
  assign n12916 = ~n9396 | ~n12922;
  assign n9398 = n12930 & n12954;
  assign n9399 = ~n12954 | ~n9127;
  assign n9624 = ~n9405 | ~n9406;
  assign n9405 = ~n13025 | ~n9146;
  assign n9409 = ~n13031;
  assign n9412 = ~n12877 | ~n9410;
  assign n12894 = ~n9412 | ~n9411;
  assign n9413 = ~n9080 | ~n12885;
  assign n11232 = ~n11229 ^ n11230;
  assign n9625 = ~n9415 | ~n9144;
  assign n9415 = ~n9416 | ~n16053;
  assign n16021 = ~n16053 | ~n13142;
  assign n9418 = ~n13142;
  assign n14724 = ~n9419 | ~n9420;
  assign n9419 = ~n9603 | ~n9053;
  assign n9422 = ~n14789 | ~n12773;
  assign n12646 = ~n14772 | ~n14789;
  assign n14772 = ~n9603 | ~n12990;
  assign n9427 = ~n9424 | ~n9426;
  assign n14584 = ~n9426 | ~n9897;
  assign n9428 = ~n9888 | ~n9007;
  assign n12645 = n9158 & n9888;
  assign n12644 = ~n9888 | ~n9889;
  assign n11569 = ~n9429 | ~n14445;
  assign n14447 = ~n9429 & ~n14444;
  assign n12307 = ~n9429 ^ n14444;
  assign n15352 = ~n15351 & ~n9430;
  assign n9430 = n11306 & n15425;
  assign n15375 = ~n9431 | ~n15374;
  assign n15427 = ~n11284 | ~n9431;
  assign n9431 = ~n11282 | ~n11283;
  assign n9432 = ~n9414 | ~n9043;
  assign n14531 = ~n14529 | ~n9433;
  assign n9433 = ~n11623 | ~n11624;
  assign n11276 = ~n9437 | ~n9434;
  assign n9435 = ~n11274;
  assign n9436 = ~n11275 | ~n11923;
  assign n9438 = ~n15333 | ~n15331;
  assign n9789 = ~n9439 | ~n9438;
  assign n9783 = ~n9448 | ~n9449;
  assign n9448 = ~n14361 | ~n9003;
  assign n14306 = ~n9077 | ~n9003;
  assign n9453 = ~n9767;
  assign n9769 = ~n14361 | ~n14358;
  assign n9457 = ~n14345 | ~n9061;
  assign n14239 = ~n9457 | ~n9776;
  assign n11929 = n9457 & n9455;
  assign n15333 = ~n11401 | ~n15451;
  assign n12073 = ~n15310 | ~n11185;
  assign n11201 = ~n11196 & ~P1_IR_REG_19__SCAN_IN;
  assign n10202 = ~n10233 | ~n10230;
  assign n9649 = ~n9024 & ~n9650;
  assign n9586 = ~n9589 | ~n9588;
  assign n9596 = ~n15437 & ~n16320;
  assign n15177 = ~n11581 | ~n11580;
  assign n9647 = ~n9649 & ~n9648;
  assign n16526 = ~n12455 | ~n16537;
  assign n12648 = ~n14654 | ~n13169;
  assign n11304 = ~n11303;
  assign n10536 = ~n13749 | ~n11112;
  assign n9952 = ~n13893;
  assign n12427 = ~n11082;
  assign n10429 = ~n9913 | ~n10404;
  assign n12474 = ~n9461 | ~n9633;
  assign n9461 = ~n9848 | ~n9489;
  assign n13379 = ~n12509 | ~n12508;
  assign n9669 = n12790 | n13183;
  assign n13634 = ~n13630 | ~n13631;
  assign n9611 = ~n9612;
  assign n9546 = ~n9501 | ~n9547;
  assign n9922 = ~n10149 | ~n9923;
  assign n14361 = ~n11634 | ~n14529;
  assign n9463 = ~n11802 | ~P1_REG0_REG_1__SCAN_IN;
  assign n16070 = ~n12800 | ~n16071;
  assign n9604 = ~n14933 | ~n9605;
  assign n10036 = ~n9658 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n9488 = ~n10081 | ~n10080;
  assign n10081 = ~n10077 | ~n10076;
  assign n10511 = ~n9516 | ~n9153;
  assign n10075 = ~n10056 | ~n10055;
  assign n9648 = ~n13459;
  assign n9847 = ~n16621 | ~n9850;
  assign n9846 = ~n9847 | ~n12465;
  assign n11628 = ~n14254 | ~n14252;
  assign n11466 = n14410 | n15365;
  assign n9466 = n9624 & n9741;
  assign n12847 = ~n12839 | ~n12838;
  assign n12830 = ~n9729 | ~n9095;
  assign n14254 = n11574 & n14449;
  assign n9794 = ~n9795 & ~n11965;
  assign n11944 = ~n11213 ^ n11212;
  assign n11134 = ~n9845;
  assign n9706 = ~n9468 | ~n9467;
  assign n9498 = ~n13104 & ~n16125;
  assign n12826 = ~n12823 & ~n9543;
  assign n9990 = ~n9992;
  assign n9992 = ~n9699 | ~n9921;
  assign n14139 = ~n9470 | ~n13969;
  assign n9470 = ~n13962 | ~n17446;
  assign n9620 = ~n14584 | ~n13180;
  assign n9858 = ~n12693 & ~n9050;
  assign n15031 = ~n14570 & ~n14569;
  assign n15894 = ~n12222 & ~n12221;
  assign n11101 = ~n11099 | ~n9472;
  assign n11110 = ~n11109 & ~n9511;
  assign n13104 = ~n12826 & ~n9504;
  assign n9543 = ~n12825 | ~n9544;
  assign n16006 = ~n9473;
  assign n10237 = ~n9475 | ~n9474;
  assign n9475 = ~n10234;
  assign P1_U3264 = ~n14602 | ~n9060;
  assign n12829 = ~n9518 | ~n16251;
  assign n9477 = ~n12232 | ~n15986;
  assign n9622 = ~n9623 & ~n9149;
  assign n12856 = ~n9478 | ~n12846;
  assign n9478 = ~n12845 | ~n16046;
  assign n12994 = ~n12988 | ~n12987;
  assign n9631 = ~n12894 | ~n12893;
  assign n11271 = n11270 & n11269;
  assign n9651 = ~n9027 | ~n9655;
  assign n9820 = ~n9823 & ~n9821;
  assign n10354 = ~n10324 | ~n10323;
  assign n12538 = ~n12535 & ~n12534;
  assign n9773 = ~n9775 & ~n9774;
  assign n14757 = ~n9593 | ~n9880;
  assign n12684 = ~n9851 | ~n9134;
  assign n9485 = ~n9481 | ~n16084;
  assign n9481 = ~n12694;
  assign n12694 = ~n9601 ^ n12824;
  assign n12236 = ~n9483 | ~n9482;
  assign n16041 = ~n16042 | ~n16051;
  assign n14642 = ~n12678 | ~n13048;
  assign n12664 = ~n14834 | ~n12663;
  assign n14834 = ~n9584 | ~n9585;
  assign n14731 = ~n9879 | ~n12669;
  assign n12882 = ~n9596;
  assign n9505 = ~n12832 ^ n12902;
  assign n12831 = ~n12829 | ~n12830;
  assign n11259 = ~n8994 | ~n11249;
  assign n9739 = ~n11176;
  assign n15394 = ~n15348 | ~n15347;
  assign n9504 = ~n12791;
  assign n11122 = ~n13538;
  assign n14141 = ~n14139 | ~n17514;
  assign n9905 = ~n9562 | ~n9560;
  assign n9553 = n9554 & n9939;
  assign n10083 = n9488 & n10082;
  assign n17298 = ~n10210 ^ n10234;
  assign n11430 = n17298 | n12401;
  assign n9660 = ~n9490 | ~n9661;
  assign n15875 = ~n9491;
  assign n14975 = ~n9492;
  assign n9871 = ~n12660;
  assign n11401 = ~n9495 | ~n9770;
  assign n9495 = ~n15394 | ~n9773;
  assign n10546 = ~n9909;
  assign n12839 = ~n9505 | ~n9497;
  assign n9774 = ~n15395;
  assign n9787 = ~n9788 & ~n11514;
  assign n9791 = ~n11467 | ~n11443;
  assign n9661 = ~n10320 & ~n9662;
  assign n10726 = ~n10716 | ~n10714;
  assign n13110 = ~n9506 | ~n9058;
  assign n13605 = ~n9499 | ~n13603;
  assign n9499 = ~n13601 | ~n13602;
  assign n13599 = n13986 | n17098;
  assign n12110 = ~n11147 | ~n14214;
  assign n13845 = ~n9754 | ~n9753;
  assign n13593 = ~n13615 | ~n13622;
  assign n11272 = ~n16078 | ~n8993;
  assign n10010 = n9921 & n9988;
  assign n17048 = ~n9922 | ~n10173;
  assign n9923 = ~n9114 & ~n9924;
  assign n9895 = ~n12733;
  assign n10920 = ~n10905 & ~n10914;
  assign n10836 = ~n10835 & ~n10834;
  assign n9515 = ~n15349;
  assign n9507 = ~n9621 | ~n9121;
  assign P1_U3238 = ~n9508 | ~n9157;
  assign n9771 = ~n9772 | ~n11371;
  assign n9636 = ~n9637 | ~n16582;
  assign n9747 = ~n17278;
  assign n10321 = ~n9663 | ~n10296;
  assign n11115 = ~n11114 | ~n9513;
  assign n9514 = ~n14519 | ~n14520;
  assign n11768 = ~n9786 | ~n11763;
  assign n10539 = ~n10514 | ~n9674;
  assign n9518 = ~n11249;
  assign n9547 = ~n9936 & ~n13933;
  assign n9550 = ~n13634 | ~n9553;
  assign n9554 = ~n13608 | ~n9555;
  assign n13610 = ~n13607 | ~n13608;
  assign n13607 = ~n13634 | ~n11022;
  assign n10508 = ~n13803 | ~n9556;
  assign n10175 = ~n10162 | ~n10161;
  assign n9559 = n10232 & n10161;
  assign n9558 = ~n10232 | ~n9561;
  assign n9562 = ~n10162 | ~n9559;
  assign n10233 = ~n10175 | ~n10174;
  assign n9561 = ~n10174;
  assign P2_U3267 = ~n9564 | ~n9563;
  assign n9564 = ~n9565 | ~n9152;
  assign n9565 = ~n9566 | ~n17087;
  assign n9566 = ~n13529;
  assign n13234 = ~n13825 | ~n13229;
  assign n9571 = ~n9572 | ~n9819;
  assign n9576 = ~n16961 | ~n9819;
  assign n16961 = ~n16960 | ~n16963;
  assign n9582 = ~n9797 | ~n9583;
  assign n9584 = ~n12659 | ~n9589;
  assign n14868 = ~n9587 | ~n9589;
  assign n9587 = ~n9592 | ~n9869;
  assign n14917 = ~n12659 | ~n12658;
  assign n9590 = ~n9869 | ~n9591;
  assign n9879 = ~n14757 | ~n12668;
  assign n9598 = ~n12684 | ~n9599;
  assign n14568 = ~n12684 | ~n12683;
  assign n11191 = n11190 & n9602;
  assign n11636 = ~n11543 | ~n9602;
  assign n9603 = ~n9884 | ~n9885;
  assign n14560 = ~n9620 | ~n12788;
  assign n9621 = ~n13079 | ~n9622;
  assign n9626 = n9627 & n12906;
  assign n9627 = ~n9631 | ~n9137;
  assign n9628 = ~n9629 | ~n12911;
  assign n9629 = ~n9630 | ~n12907;
  assign n9630 = ~n9631 | ~n12899;
  assign n16430 = ~n9846 | ~n9848;
  assign n16474 = ~n9632 | ~n12469;
  assign n9632 = ~n16430 | ~n16431;
  assign n9635 = ~n12469;
  assign n9822 = ~n9638 | ~n9643;
  assign n9638 = ~n9645 | ~n16582;
  assign n12494 = ~n9642 | ~n9639;
  assign n9639 = n9640 & n9820;
  assign n9641 = ~n16582;
  assign n9642 = ~n16584 | ~n9643;
  assign n16503 = ~n9644 | ~n16582;
  assign n9644 = ~n16585 | ~n16583;
  assign n12534 = ~n12609 & ~n12610;
  assign n13460 = ~n9646 | ~n12514;
  assign n9646 = ~n9494 | ~n9024;
  assign n9650 = ~n12514;
  assign n9652 = ~n9828 | ~n9027;
  assign n13359 = ~n9653 | ~n12523;
  assign n9653 = ~n9493 | ~n9826;
  assign n9654 = ~n9827 | ~n12523;
  assign n9655 = ~n12523;
  assign n9910 = ~n9657 | ~n10122;
  assign n17333 = ~n9657 ^ n10122;
  assign n10056 = ~n9658 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n9911 = ~n9660 | ~n9142;
  assign n9659 = ~n9661 | ~n10293;
  assign n10324 = ~n9663 | ~n9661;
  assign n9663 = ~n10295 | ~n10294;
  assign n9664 = ~n10461;
  assign n12771 = ~n13164 | ~n12770;
  assign n12776 = ~n9666 | ~n12797;
  assign n9666 = n12726 | n13020;
  assign n9670 = ~n10380 | ~n9672;
  assign n9671 = ~n9672 | ~n9915;
  assign n9673 = ~n9914 | ~n10378;
  assign n15101 = ~n9676 | ~n11746;
  assign n12401 = ~n11263 | ~n11973;
  assign n9681 = ~n9682 | ~n14737;
  assign n14733 = ~n14790 & ~n9683;
  assign n14920 = ~n14977 & ~n15188;
  assign n9691 = ~n14919 | ~n9692;
  assign n9692 = ~n15188;
  assign n12695 = ~n14621 | ~n9695;
  assign n14596 = ~n14621 | ~n14622;
  assign n9988 = ~n11133;
  assign n9921 = n9956 & n10007;
  assign n9956 = n9987 & n10440;
  assign n9700 = ~n10940;
  assign n9701 = ~n9098;
  assign n9702 = ~n9083 | ~n9703;
  assign n9705 = ~n11007 | ~n9707;
  assign n9711 = ~n10898 & ~n10884;
  assign n10905 = ~n9713 | ~n9712;
  assign n9712 = ~n10895 | ~n9714;
  assign n9714 = ~n10898;
  assign n11049 = ~n9716 | ~n9069;
  assign n9715 = ~n9719 | ~n9718;
  assign n9716 = ~n11031 | ~n9719;
  assign n9719 = n9717 & n11041;
  assign n9717 = ~n11036 | ~n9065;
  assign n10837 = ~n10827 | ~n9720;
  assign n9720 = n9721 | n10823;
  assign n9721 = ~n16570 | ~n10828;
  assign n9722 = ~n10970 & ~n9726;
  assign n9725 = ~n10970;
  assign n16071 = ~n12830;
  assign n9733 = ~n9731 | ~n9730;
  assign n9731 = ~n13079 | ~n9732;
  assign n9734 = ~n12994 | ~n9735;
  assign n13002 = ~n12994 | ~n12993;
  assign n13015 = ~n13008 | ~n9070;
  assign n9740 = n11210 & n11209;
  assign n11214 = ~n9740 | ~n11211;
  assign n11227 = ~n9740 | ~n9737;
  assign n9744 = ~n13044 | ~n9130;
  assign n13202 = ~n13121 & ~n13120;
  assign n10080 = n10079 & SI_1_;
  assign n12961 = n12963 | n14535;
  assign n11581 = n17258 | n12401;
  assign n13951 = ~n9745 | ~n17555;
  assign n14135 = ~n9745 | ~n17514;
  assign n9745 = ~n9008 | ~n9126;
  assign n10100 = n10245 | n17333;
  assign n10125 = n17326 | n10245;
  assign n10732 = ~n10245;
  assign n17142 = ~n17185 | ~n12439;
  assign n13908 = ~n16943 & ~n9757;
  assign n11921 = ~n15025 & ~n9766;
  assign n11241 = ~n14622 & ~n9766;
  assign n9766 = ~n12268 | ~n12073;
  assign n12205 = ~n15392 | ~n15396;
  assign n14519 = ~n9782 | ~n14343;
  assign n9780 = ~n14520 & ~n9781;
  assign n9786 = ~n9783 | ~n9784;
  assign n11522 = ~n9789 | ~n9787;
  assign P1_U3218 = ~n9794 | ~n9792;
  assign n9792 = n11929 | n9793;
  assign n9802 = ~n13217;
  assign n17057 = ~n9803 | ~n13217;
  assign n9803 = ~n17077 | ~n17081;
  assign n9804 = ~n9805 | ~n13217;
  assign n13773 = ~n9806 | ~n13235;
  assign n9806 = ~n13234 | ~n9807;
  assign n13799 = ~n13234 | ~n13233;
  assign n9808 = ~n13233;
  assign n9815 = ~n13558 | ~n9817;
  assign n9813 = ~n9817 | ~n9814;
  assign n13554 = ~n9816 | ~n13256;
  assign n9816 = ~n13558 | ~n13560;
  assign n9818 = ~n13557 | ~n13256;
  assign n10005 = n10010 | n10523;
  assign n12643 = ~n9824 | ~n12635;
  assign n9825 = ~n12622 | ~n9138;
  assign n12629 = ~n12622 | ~n12621;
  assign n16584 = ~n9829 | ~n9830;
  assign n9829 = ~n16550 | ~n9834;
  assign n9831 = ~n9834 | ~n9832;
  assign n16445 = ~n9833 | ~n16551;
  assign n9833 = ~n16554 | ~n16552;
  assign n9835 = ~n9836 | ~n16551;
  assign n13294 = ~n9837 | ~n9129;
  assign n9837 = ~n9838 | ~n9012;
  assign n9838 = ~n12609;
  assign n9839 = ~n9012 | ~n12615;
  assign n9841 = ~n12608 | ~n9843;
  assign n10465 = ~n9845 | ~n10441;
  assign n9848 = ~n16526 | ~n9109;
  assign n16620 = ~n9849 | ~n16523;
  assign n9849 = n16526 | n16522;
  assign n9850 = ~n16522 | ~n16523;
  assign n9851 = ~n12680 | ~n9852;
  assign n9854 = ~n14616 | ~n12681;
  assign n9857 = ~n12682;
  assign n14661 = ~n9859 | ~n12676;
  assign n9859 = ~n12674 | ~n9863;
  assign n9861 = ~n9862 | ~n12676;
  assign n9866 = ~n9869 | ~n9867;
  assign n14884 = ~n9868 | ~n12661;
  assign n9868 = ~n14917 | ~n12660;
  assign n9870 = ~n9871 | ~n12661;
  assign n9873 = ~n9876 | ~n9874;
  assign n14963 = ~n9875 | ~n12655;
  assign n9875 = ~n14992 | ~n12653;
  assign n9877 = ~n9878 | ~n12655;
  assign n14959 = n12645 | n9883;
  assign n14989 = ~n12645 & ~n12732;
  assign n9884 = ~n14856 | ~n9002;
  assign n9888 = ~n15896 | ~n9893;
  assign n9890 = ~n9893 | ~n9891;
  assign n15845 = ~n9892 | ~n12895;
  assign n9892 = ~n15896 | ~n12733;
  assign n9894 = ~n9895 | ~n12895;
  assign n14604 = ~n12648 | ~n9096;
  assign n9904 = ~n12795;
  assign n17291 = ~n9905 ^ n10264;
  assign n9906 = ~n10548 | ~n9907;
  assign n10563 = ~n9909 | ~n10548;
  assign n9909 = ~n10539 | ~n10538;
  assign n10140 = ~n9910 | ~n10124;
  assign n10143 = ~n10140 | ~n10139;
  assign n10402 = ~n10382 | ~n10381;
  assign n10678 = ~n10716;
  assign n11142 = ~n9988 | ~n9956;
  assign n17082 = ~n10149 | ~n11096;
  assign n9924 = ~n11096;
  assign n9925 = ~n10536 | ~n9929;
  assign n9927 = ~n9929 | ~n9932;
  assign n9930 = ~n10560 | ~n9931;
  assign n13702 = ~n9928 | ~n9929;
  assign n9928 = n10536 | n9932;
  assign n13726 = ~n10536 | ~n11111;
  assign n9932 = ~n10560;
  assign n9938 = ~n10319 | ~n11105;
  assign n9934 = ~n11105;
  assign n9935 = ~n9938 | ~n10352;
  assign n9940 = ~n10105 | ~n9966;
  assign n17116 = ~n9940 | ~n10106;
  assign n9943 = ~n13266 | ~n9944;
  assign n9949 = ~n13678 | ~n10999;
  assign n13654 = ~n9949 ^ n9947;
  assign n9950 = ~n9951 | ~n9006;
  assign n9951 = ~n13892;
  assign n9953 = ~n13892;
  assign n13017 = n13020 | n13003;
  assign n13787 = ~n13847 & ~n13279;
  assign n10017 = ~n10016 | ~n10015;
  assign n14737 = ~n15101;
  assign n11924 = ~n12247 | ~n12073;
  assign n12247 = ~n12268;
  assign n13102 = n13107 | n9500;
  assign n14220 = ~n11142 | ~n11141;
  assign n17197 = n10826 & n16568;
  assign n11988 = n10826;
  assign n10062 = n11095 & n10061;
  assign n10245 = ~n12110 | ~n10357;
  assign n9996 = ~n9993 ^ n9989;
  assign n13330 = ~n12529 & ~n12530;
  assign n9993 = ~n9992 | ~P2_IR_REG_31__SCAN_IN;
  assign n10060 = n10049 & n10048;
  assign n10049 = n10101 | n11976;
  assign n10258 = n14196 & n9996;
  assign n11263 = ~n11944 | ~n15494;
  assign n14187 = ~n9990 | ~n9989;
  assign n9955 = n11122 | n13537;
  assign n9989 = ~P2_IR_REG_29__SCAN_IN;
  assign n12584 = ~n13260;
  assign n11126 = ~n12335;
  assign n9960 = n10721 & n10720;
  assign n9961 = n10065 & P2_REG2_REG_1__SCAN_IN;
  assign n9962 = n10065 & P2_REG2_REG_2__SCAN_IN;
  assign n9963 = n11154 | n13271;
  assign n9964 = n12617 | n12616;
  assign n9965 = ~n12519 | ~n12518;
  assign n9966 = n16541 | n17141;
  assign n9967 = n12611 & n12613;
  assign n9968 = ~n12493 | ~n12492;
  assign n10177 = n9658;
  assign n10357 = ~n10085;
  assign n10163 = ~n10085;
  assign n9979 = ~P2_IR_REG_5__SCAN_IN & ~P2_IR_REG_4__SCAN_IN;
  assign n13174 = n13177 & n14605;
  assign n12774 = n12989 & n14800;
  assign n11168 = ~P1_IR_REG_17__SCAN_IN & ~P1_IR_REG_18__SCAN_IN;
  assign n10581 = ~SI_22_;
  assign n13226 = ~n16934;
  assign n10521 = ~P2_IR_REG_18__SCAN_IN;
  assign n11913 = n11855 & P1_REG3_REG_26__SCAN_IN;
  assign n10720 = n10723 | n10722;
  assign n10650 = n10645 & n10644;
  assign n11336 = ~P1_IR_REG_3__SCAN_IN;
  assign n10000 = n10258 & P2_REG0_REG_0__SCAN_IN;
  assign n13279 = ~n13813;
  assign n13219 = ~n17033;
  assign n11138 = ~P2_IR_REG_26__SCAN_IN;
  assign n10517 = ~SI_19_;
  assign n14562 = ~n16419;
  assign n11903 = P1_D_REG_29__SCAN_IN | n11902;
  assign n11233 = ~n11232;
  assign n11747 = n11733 & P1_REG3_REG_20__SCAN_IN;
  assign n16077 = ~n16023;
  assign n11213 = ~n11227 | ~P1_IR_REG_31__SCAN_IN;
  assign n10675 = n10673 & n10672;
  assign n10433 = ~SI_16_;
  assign n11125 = n11124 | P2_IR_REG_22__SCAN_IN;
  assign n13255 = ~n17582;
  assign n16490 = ~n10826;
  assign n16605 = ~n12584 | ~n12598;
  assign n13274 = ~n17585;
  assign n10683 = n10664 & P2_REG3_REG_24__SCAN_IN;
  assign n10552 = n10532 & P2_REG3_REG_18__SCAN_IN;
  assign n13805 = ~n13395;
  assign n17504 = n11082 & n12595;
  assign n17493 = ~n13265 | ~n10825;
  assign n10542 = ~SI_20_;
  assign n11711 = n11666 | n11225;
  assign n11713 = ~n11711 & ~n11710;
  assign n11825 = ~n12401;
  assign n12287 = n16122 & n11903;
  assign n16084 = ~n16045;
  assign n14935 = n12959 & n12955;
  assign n15175 = ~n15056;
  assign n16045 = n12250 & n12249;
  assign n12288 = ~n12287;
  assign n11215 = ~P1_IR_REG_27__SCAN_IN;
  assign n10605 = n10588 & n10586;
  assign n11129 = ~P2_IR_REG_23__SCAN_IN;
  assign n16624 = ~n13321 | ~n13320;
  assign n13557 = ~n13560;
  assign n17173 = ~n13264 | ~n13263;
  assign n13801 = n10487 & n10486;
  assign n13510 = ~n17357 & ~n12571;
  assign n13639 = n13638 | n13637;
  assign n17212 = ~n13269 | ~n13268;
  assign n13290 = n12581 | n17227;
  assign n17239 = n10472 & n10471;
  assign n15438 = ~n11948 | ~n11945;
  assign n15378 = ~n12260 | ~n16241;
  assign n14608 = ~n16407;
  assign n13109 = ~n13192;
  assign n11658 = ~n11636 & ~P1_IR_REG_16__SCAN_IN;
  assign n16116 = ~n16025;
  assign n12693 = ~n12651 & ~n16074;
  assign n11185 = n12346 & n15319;
  assign n10660 = n10671 & n10659;
  assign n10355 = n10356 & n10330;
  assign n12588 = ~n11130 ^ n11129;
  assign n16554 = n16550;
  assign n13491 = n13837 & n12487;
  assign n16472 = ~P2_REG3_REG_8__SCAN_IN;
  assign n12152 = ~n12144 & ~P2_U3966;
  assign n17068 = ~n17087 | ~n17191;
  assign n13948 = ~n12576 | ~n12575;
  assign n13949 = n13290 & n13289;
  assign n12329 = ~n11173 ^ n11172;
  assign n15419 = ~n15438;
  assign n15441 = ~n15429;
  assign n15447 = ~n15402;
  assign n15442 = n11934 & n16011;
  assign n15653 = n15465 | n15496;
  assign n15996 = n16104 | n16059;
  assign n14918 = ~n14643;
  assign n12291 = ~n12294;
  assign n16122 = n11872 & n15310;
  assign n11187 = ~n12588 | ~P2_STATE_REG_SCAN_IN;
  assign n16622 = ~n16575;
  assign n16631 = n12597 & n12596;
  assign n17595 = n10779 | n10778;
  assign n17564 = n10576 | n10575;
  assign n16872 = ~n12152 & ~n12598;
  assign n17206 = ~n17068;
  assign n17186 = n17087 & n13512;
  assign n17218 = ~n17087;
  assign n14184 = n14131 | n14130;
  assign n17340 = ~n14227;
  assign n17347 = ~n14229;
  assign n15402 = n15379 | n11942;
  assign n15414 = ~n15457;
  assign n16404 = n11792 | n11791;
  assign n14509 = n11692 | n11691;
  assign n15881 = ~n12908;
  assign n15816 = ~n15653;
  assign n16040 = n16104 | n15940;
  assign n16105 = ~n16011;
  assign n16104 = n12263 & n16011;
  assign n15317 = n11973 & P1_U3084;
  assign n17647 = P1_ADDR_REG_10__SCAN_IN & P2_ADDR_REG_10__SCAN_IN;
  assign n17643 = P1_ADDR_REG_11__SCAN_IN & P2_ADDR_REG_11__SCAN_IN;
  assign n17594 = n12586 | n11187;
  assign n17350 = ~n17225 | ~n17224;
  assign n16425 = ~n12085 | ~P1_STATE_REG_SCAN_IN;
  assign n17650 = ~n12381 & ~n12380;
  assign n17642 = ~n17644 & ~n12383;
  assign P2_U3966 = ~n17594;
  assign P1_U4006 = ~n16425;
  assign n9969 = ~P2_IR_REG_24__SCAN_IN;
  assign n9972 = n9970 & n9969;
  assign n9971 = ~P2_IR_REG_17__SCAN_IN & ~P2_IR_REG_16__SCAN_IN;
  assign n9976 = ~n9972 | ~n9971;
  assign n9974 = ~P2_IR_REG_21__SCAN_IN & ~P2_IR_REG_20__SCAN_IN;
  assign n9973 = ~P2_IR_REG_19__SCAN_IN & ~P2_IR_REG_18__SCAN_IN;
  assign n9975 = ~n9974 | ~n9973;
  assign n10090 = ~P2_IR_REG_2__SCAN_IN;
  assign n11133 = ~n9978 | ~n10441;
  assign n10212 = ~P2_IR_REG_6__SCAN_IN & ~P2_IR_REG_7__SCAN_IN;
  assign n10438 = ~n9979 | ~n10212;
  assign n9980 = ~n11144 | ~n11138;
  assign n9986 = n9982 & n9981;
  assign n10440 = n9986 & n9985;
  assign n9994 = ~n14187 | ~P2_IR_REG_31__SCAN_IN;
  assign n14196 = ~n9994 ^ n9991;
  assign n9995 = ~n9996;
  assign n10777 = n14196 & n9995;
  assign n10003 = ~n10777 | ~P2_REG1_REG_0__SCAN_IN;
  assign n9997 = ~n9994 ^ P2_IR_REG_30__SCAN_IN;
  assign n10068 = n9997 & n9995;
  assign n9999 = ~n10068 | ~P2_REG3_REG_0__SCAN_IN;
  assign n10065 = n9997 & n9996;
  assign n9998 = ~n10065 | ~P2_REG2_REG_0__SCAN_IN;
  assign n10001 = ~n9999 | ~n9998;
  assign n10002 = ~n10001 & ~n10000;
  assign n10826 = ~n10003 | ~n10002;
  assign n11147 = ~n10005 ^ n10004;
  assign n10006 = ~n11142 | ~P2_IR_REG_31__SCAN_IN;
  assign n10009 = ~n10006 | ~P2_IR_REG_27__SCAN_IN;
  assign n10007 = ~P2_IR_REG_27__SCAN_IN;
  assign n10008 = ~n10007 | ~P2_IR_REG_31__SCAN_IN;
  assign n10011 = ~n10010;
  assign n14214 = ~n10012 | ~n10011;
  assign n10021 = ~n10089 | ~P2_IR_REG_0__SCAN_IN;
  assign n10014 = P2_ADDR_REG_19__SCAN_IN & P1_ADDR_REG_19__SCAN_IN;
  assign n10054 = ~n10018 | ~n10017;
  assign n10019 = ~n10177 | ~SI_0_;
  assign n11966 = ~n10019 ^ P1_DATAO_REG_0__SCAN_IN;
  assign n10020 = ~n12110 | ~n11966;
  assign n16568 = ~n10021 | ~n10020;
  assign n10026 = ~n10777 | ~P2_REG1_REG_1__SCAN_IN;
  assign n10023 = ~n10258 | ~P2_REG0_REG_1__SCAN_IN;
  assign n10022 = ~n10068 | ~P2_REG3_REG_1__SCAN_IN;
  assign n10024 = ~n10023 | ~n10022;
  assign n10025 = ~n10024 & ~n9961;
  assign n10027 = ~n12430;
  assign n10042 = ~n17161 | ~n10027;
  assign n10085 = n10054;
  assign n10028 = ~P2_IR_REG_1__SCAN_IN;
  assign n10031 = ~n10028 | ~P2_IR_REG_31__SCAN_IN;
  assign n10029 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign n10030 = ~n10029 | ~P2_IR_REG_1__SCAN_IN;
  assign n10032 = ~n10031 | ~n10030;
  assign n10033 = ~n10089 | ~n17342;
  assign n10035 = ~n10054 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n10079 = ~n10036 | ~n10035;
  assign n10038 = ~n9658 | ~P1_DATAO_REG_0__SCAN_IN;
  assign n10037 = ~n10054 | ~P2_DATAO_REG_0__SCAN_IN;
  assign n10039 = ~n10038 | ~n10037;
  assign n10073 = ~n10039 | ~SI_0_;
  assign n10050 = ~n10073 ^ SI_1_;
  assign n17341 = ~n10079 ^ n10050;
  assign n10040 = n10245 | n17341;
  assign n10063 = ~n10042 | ~n12429;
  assign n10046 = ~n9954 & ~n9962;
  assign n10044 = ~n10258 | ~P2_REG0_REG_2__SCAN_IN;
  assign n10043 = ~n10068 | ~P2_REG3_REG_2__SCAN_IN;
  assign n10045 = n10044 & n10043;
  assign n11976 = ~P1_DATAO_REG_2__SCAN_IN;
  assign n12194 = ~n10047 ^ P2_IR_REG_2__SCAN_IN;
  assign n10048 = ~n10089 | ~n12194;
  assign n10053 = ~n10050 | ~n10079;
  assign n10051 = ~n10073;
  assign n10052 = ~n10051 | ~SI_1_;
  assign n10058 = ~n10053 | ~n10052;
  assign n10055 = ~n10054 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n10076 = ~SI_2_;
  assign n10057 = ~n10075 ^ n10076;
  assign n11972 = ~n10058 ^ n10057;
  assign n10059 = n10245 | n11972;
  assign n11095 = ~n16463 | ~n12439;
  assign n10064 = ~n10063 | ~n10062;
  assign n10396 = ~n10065;
  assign n10067 = ~n10481 | ~P2_REG2_REG_3__SCAN_IN;
  assign n10066 = ~n10777 | ~P2_REG1_REG_3__SCAN_IN;
  assign n10072 = ~n10067 | ~n10066;
  assign n10070 = ~n10258 | ~P2_REG0_REG_3__SCAN_IN;
  assign n16456 = ~P2_REG3_REG_3__SCAN_IN;
  assign n10069 = ~n10068 | ~n16456;
  assign n10071 = ~n10070 | ~n10069;
  assign n16541 = n10072 | n10071;
  assign n10074 = ~n10079 & ~SI_1_;
  assign n10078 = ~n10074 & ~n10073;
  assign n10077 = ~n10075;
  assign n10084 = ~n10078 | ~n10081;
  assign n10082 = ~n10075 | ~SI_2_;
  assign n10087 = ~n10163 | ~P1_DATAO_REG_3__SCAN_IN;
  assign n10086 = ~n10085 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n10123 = ~n10087 | ~n10086;
  assign n10088 = ~SI_3_;
  assign n10122 = ~n10123 ^ n10088;
  assign n10098 = ~n10441;
  assign n10092 = n10091 & n10090;
  assign n10093 = n10092 | n10523;
  assign n10096 = ~n10093 | ~P2_IR_REG_3__SCAN_IN;
  assign n10095 = ~n10094 | ~P2_IR_REG_31__SCAN_IN;
  assign n10097 = ~n10096 | ~n10095;
  assign n10099 = ~n12102 | ~n17334;
  assign n10104 = n10100 & n10099;
  assign n10102 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n10103 = n10768 | n10102;
  assign n17141 = n10104 & n10103;
  assign n10106 = ~n16541 | ~n17141;
  assign n10108 = ~n10481 | ~P2_REG2_REG_4__SCAN_IN;
  assign n10107 = ~n10777 | ~P2_REG1_REG_4__SCAN_IN;
  assign n10114 = ~n10108 | ~n10107;
  assign n10112 = ~n10258 | ~P2_REG0_REG_4__SCAN_IN;
  assign n16534 = ~P2_REG3_REG_4__SCAN_IN;
  assign n10109 = ~n16456 | ~n16534;
  assign n10153 = ~P2_REG3_REG_4__SCAN_IN | ~P2_REG3_REG_3__SCAN_IN;
  assign n17125 = ~n10109 | ~n10153;
  assign n10110 = ~n17125;
  assign n10111 = ~n10068 | ~n10110;
  assign n10113 = ~n10112 | ~n10111;
  assign n16517 = n10114 | n10113;
  assign n10866 = ~n16517;
  assign n10115 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n10118 = n10101 | n10115;
  assign n10116 = n10441 | n10523;
  assign n17327 = ~n10116 ^ P2_IR_REG_4__SCAN_IN;
  assign n10117 = ~n12102 | ~n17327;
  assign n10126 = n10118 & n10117;
  assign n10120 = ~n10177 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n10119 = ~n11975 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n10141 = ~n10120 | ~n10119;
  assign n10121 = ~SI_4_;
  assign n10139 = ~n10141 ^ n10121;
  assign n10124 = ~n10123 | ~SI_3_;
  assign n17326 = ~n10140 ^ n10139;
  assign n17133 = n10126 & n10125;
  assign n10127 = ~n16517 | ~n17133;
  assign n17102 = ~n10153 ^ P2_REG3_REG_5__SCAN_IN;
  assign n10129 = ~n10684 | ~n17102;
  assign n10128 = ~n10777 | ~P2_REG1_REG_5__SCAN_IN;
  assign n10133 = ~n10129 | ~n10128;
  assign n10131 = ~n10258 | ~P2_REG0_REG_5__SCAN_IN;
  assign n10130 = ~n10481 | ~P2_REG2_REG_5__SCAN_IN;
  assign n10132 = ~n10131 | ~n10130;
  assign n13214 = ~n16625;
  assign n10768 = ~n9173;
  assign n10134 = ~P1_DATAO_REG_5__SCAN_IN;
  assign n10138 = n10768 | n10134;
  assign n10135 = ~P2_IR_REG_4__SCAN_IN;
  assign n10168 = ~n10441 | ~n10135;
  assign n10136 = ~n10168 | ~P2_IR_REG_31__SCAN_IN;
  assign n17320 = ~n10136 ^ P2_IR_REG_5__SCAN_IN;
  assign n10137 = ~n12102 | ~n17320;
  assign n10148 = n10138 & n10137;
  assign n10142 = ~n10141 | ~SI_4_;
  assign n10145 = ~n10357 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n10144 = ~n11973 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n10160 = ~n10145 | ~n10144;
  assign n10146 = ~SI_5_;
  assign n10158 = ~n10160 ^ n10146;
  assign n17319 = ~n10159 ^ n10158;
  assign n11097 = ~n13214 | ~n17095;
  assign n10149 = ~n17091 | ~n11097;
  assign n11096 = ~n16625 | ~n17419;
  assign n10151 = ~n10258 | ~P2_REG0_REG_6__SCAN_IN;
  assign n10150 = ~n10481 | ~P2_REG2_REG_6__SCAN_IN;
  assign n10157 = n10151 & n10150;
  assign n10684 = n10068;
  assign n10152 = ~P2_REG3_REG_5__SCAN_IN;
  assign n10192 = ~n10153 & ~n10152;
  assign n16618 = ~P2_REG3_REG_6__SCAN_IN;
  assign n17069 = ~n10192 ^ n16618;
  assign n10155 = ~n10684 | ~n17069;
  assign n10154 = ~n10777 | ~P2_REG1_REG_6__SCAN_IN;
  assign n10156 = n10155 & n10154;
  assign n10162 = ~n10159 | ~n10158;
  assign n10161 = ~n10160 | ~SI_5_;
  assign n10165 = ~n10357 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n12394 = ~n10163;
  assign n10164 = ~n12394 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n10176 = ~n10165 | ~n10164;
  assign n10166 = ~SI_6_;
  assign n10174 = ~n10176 ^ n10166;
  assign n17312 = ~n10175 ^ n10174;
  assign n10167 = ~P1_DATAO_REG_6__SCAN_IN;
  assign n10171 = n10768 | n10167;
  assign n10169 = ~n10214 | ~P2_IR_REG_31__SCAN_IN;
  assign n17313 = ~n10169 ^ P2_IR_REG_6__SCAN_IN;
  assign n10170 = ~n12102 | ~n17313;
  assign n10172 = n10171 & n10170;
  assign n10173 = ~n16516 | ~n17432;
  assign n10230 = ~n10176 | ~SI_6_;
  assign n10179 = ~n10357 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n11975 = ~n10163;
  assign n10178 = ~n11975 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n10181 = n10179 & n10178;
  assign n10180 = ~SI_7_;
  assign n10235 = ~n10181 | ~n10180;
  assign n10182 = ~n10181;
  assign n10229 = ~n10182 | ~SI_7_;
  assign n10200 = n10235 & n10229;
  assign n10183 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n10189 = n10768 | n10183;
  assign n10185 = ~n10214;
  assign n10184 = ~P2_IR_REG_6__SCAN_IN;
  assign n10186 = ~n10185 | ~n10184;
  assign n10187 = ~n10186 | ~P2_IR_REG_31__SCAN_IN;
  assign n17306 = ~n10187 ^ P2_IR_REG_7__SCAN_IN;
  assign n10188 = ~n12102 | ~n17306;
  assign n10190 = n10189 & n10188;
  assign n17443 = ~n10191 | ~n10190;
  assign n10194 = ~n10258 | ~P2_REG0_REG_7__SCAN_IN;
  assign n10221 = ~n10192 | ~P2_REG3_REG_6__SCAN_IN;
  assign n17054 = ~n10221 ^ P2_REG3_REG_7__SCAN_IN;
  assign n10193 = ~n10684 | ~n17054;
  assign n10198 = n10194 & n10193;
  assign n10196 = ~n10481 | ~P2_REG2_REG_7__SCAN_IN;
  assign n10195 = ~n10777 | ~P2_REG1_REG_7__SCAN_IN;
  assign n10197 = n10196 & n10195;
  assign n10889 = n17443 | n12026;
  assign n10199 = ~n17048 | ~n10889;
  assign n10890 = ~n17443 | ~n12026;
  assign n17032 = ~n10199 | ~n10890;
  assign n10201 = ~n10200;
  assign n10205 = ~n10357 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n10204 = ~n11975 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n10206 = ~SI_8_;
  assign n10236 = ~n10207 | ~n10206;
  assign n10208 = ~n10207;
  assign n10209 = ~n10208 | ~SI_8_;
  assign n10219 = n17298 | n10698;
  assign n10211 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n10217 = n10768 | n10211;
  assign n10213 = ~n10212;
  assign n10248 = ~n10214 & ~n10213;
  assign n10215 = n10248 | n10523;
  assign n17299 = ~n10215 ^ P2_IR_REG_8__SCAN_IN;
  assign n10216 = ~n12102 | ~n17299;
  assign n10218 = n10217 & n10216;
  assign n10220 = ~P2_REG3_REG_7__SCAN_IN;
  assign n17023 = ~n10254 ^ P2_REG3_REG_8__SCAN_IN;
  assign n10223 = ~n10068 | ~n17023;
  assign n10222 = ~n10777 | ~P2_REG1_REG_8__SCAN_IN;
  assign n10227 = ~n10223 | ~n10222;
  assign n10225 = ~n8990 | ~P2_REG0_REG_8__SCAN_IN;
  assign n10224 = ~n10481 | ~P2_REG2_REG_8__SCAN_IN;
  assign n10226 = ~n10225 | ~n10224;
  assign n13220 = ~n17041 | ~n16558;
  assign n10228 = n17041 | n16558;
  assign n16989 = ~n17032 | ~n17033;
  assign n16435 = ~n16558;
  assign n16990 = ~n17041 | ~n16435;
  assign n10231 = ~n10230 | ~n10229;
  assign n10238 = n10237 & n10236;
  assign n10240 = ~n10177 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n10239 = ~n11973 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n10266 = ~n10242 | ~n10241;
  assign n10243 = ~n10242;
  assign n10244 = ~n10243 | ~SI_9_;
  assign n10264 = ~n10266 | ~n10244;
  assign n10253 = n17291 | n10698;
  assign n10246 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n10251 = n10768 | n10246;
  assign n10247 = ~P2_IR_REG_8__SCAN_IN;
  assign n10249 = n10334 | n10523;
  assign n17292 = ~n10249 ^ P2_IR_REG_9__SCAN_IN;
  assign n10250 = ~n17292 | ~n12102;
  assign n10252 = n10251 & n10250;
  assign n17465 = ~n10253 | ~n10252;
  assign n10281 = ~n10254 & ~n16472;
  assign n10255 = ~P2_REG3_REG_9__SCAN_IN;
  assign n17005 = ~n10281 ^ n10255;
  assign n10257 = ~n10684 | ~n17005;
  assign n10256 = ~n10481 | ~P2_REG2_REG_9__SCAN_IN;
  assign n10262 = ~n10257 | ~n10256;
  assign n10260 = ~n8990 | ~P2_REG0_REG_9__SCAN_IN;
  assign n10259 = ~n10777 | ~P2_REG1_REG_9__SCAN_IN;
  assign n10261 = ~n10260 | ~n10259;
  assign n10288 = ~n16477;
  assign n16991 = ~n17465 | ~n10288;
  assign n10263 = n16990 & n16991;
  assign n10291 = ~n16989 | ~n10263;
  assign n10265 = ~n10264;
  assign n10269 = ~n10177 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n10268 = ~n12394 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n10296 = ~n10271 | ~n10270;
  assign n10272 = ~n10271;
  assign n10273 = ~n10272 | ~SI_10_;
  assign n10293 = ~n10296 | ~n10273;
  assign n10280 = n17284 | n10698;
  assign n10274 = ~P2_IR_REG_9__SCAN_IN;
  assign n10275 = ~n10334 | ~n10274;
  assign n10300 = ~n10275 | ~P2_IR_REG_31__SCAN_IN;
  assign n17285 = ~n10300 ^ P2_IR_REG_10__SCAN_IN;
  assign n10278 = ~n17285 | ~n12102;
  assign n10276 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n10277 = n10768 | n10276;
  assign n10279 = n10278 & n10277;
  assign n17476 = ~n10280 | ~n10279;
  assign n16443 = ~P2_REG3_REG_10__SCAN_IN;
  assign n16980 = ~n10312 ^ n16443;
  assign n10283 = ~n10684 | ~n16980;
  assign n10282 = ~n10777 | ~P2_REG1_REG_10__SCAN_IN;
  assign n10287 = ~n10283 | ~n10282;
  assign n10285 = ~n10258 | ~P2_REG0_REG_10__SCAN_IN;
  assign n10284 = ~n10065 | ~P2_REG2_REG_10__SCAN_IN;
  assign n10286 = ~n10285 | ~n10284;
  assign n16591 = ~n16559;
  assign n10289 = n17476 | n16591;
  assign n10913 = n17465 | n10288;
  assign n10290 = n10289 & n10913;
  assign n10292 = ~n17476 | ~n16591;
  assign n10294 = ~n10293;
  assign n10298 = ~n12395 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n10297 = ~n11973 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n10322 = ~n10298 | ~n10297;
  assign n10320 = ~n10322 ^ SI_11_;
  assign n17278 = ~n10321 ^ n10320;
  assign n10299 = ~P2_IR_REG_10__SCAN_IN | ~P2_IR_REG_31__SCAN_IN;
  assign n10301 = ~n10300 | ~n10299;
  assign n10331 = ~P2_IR_REG_11__SCAN_IN;
  assign n16779 = ~n10301 ^ n10331;
  assign n10304 = ~n16779 | ~n12102;
  assign n10302 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n10303 = n10768 | n10302;
  assign n10305 = n10304 & n10303;
  assign n10308 = ~n10481 | ~P2_REG2_REG_11__SCAN_IN;
  assign n10307 = ~n10777 | ~P2_REG1_REG_11__SCAN_IN;
  assign n10318 = n10308 & n10307;
  assign n10316 = ~n8990 | ~P2_REG0_REG_11__SCAN_IN;
  assign n10310 = ~n10312 | ~P2_REG3_REG_10__SCAN_IN;
  assign n10309 = ~P2_REG3_REG_11__SCAN_IN;
  assign n10313 = ~n10310 | ~n10309;
  assign n10311 = P2_REG3_REG_10__SCAN_IN & P2_REG3_REG_11__SCAN_IN;
  assign n10393 = ~n10312 | ~n10311;
  assign n16950 = ~n10313 | ~n10393;
  assign n10314 = ~n16950;
  assign n10315 = ~n10684 | ~n10314;
  assign n10317 = n10316 & n10315;
  assign n11105 = ~n16955 | ~n10921;
  assign n10323 = ~n10322 | ~SI_11_;
  assign n10326 = ~n12395 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n10325 = ~n11973 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n10327 = ~SI_12_;
  assign n10356 = ~n10328 | ~n10327;
  assign n10329 = ~n10328;
  assign n10330 = ~n10329 | ~SI_12_;
  assign n17271 = ~n10354 ^ n10355;
  assign n10332 = ~P2_IR_REG_9__SCAN_IN & ~P2_IR_REG_10__SCAN_IN;
  assign n10333 = n10332 & n10331;
  assign n10335 = n10339 | n10523;
  assign n10337 = ~n10335 | ~P2_IR_REG_12__SCAN_IN;
  assign n10338 = ~P2_IR_REG_12__SCAN_IN;
  assign n10336 = ~n10338 | ~P2_IR_REG_31__SCAN_IN;
  assign n10340 = ~n10337 | ~n10336;
  assign n10385 = ~n10339 | ~n10338;
  assign n10343 = ~n17272 | ~n12102;
  assign n10341 = ~P1_DATAO_REG_12__SCAN_IN;
  assign n10342 = n10768 | n10341;
  assign n10344 = n10343 & n10342;
  assign n10347 = ~n8990 | ~P2_REG0_REG_12__SCAN_IN;
  assign n16940 = ~n10393 ^ P2_REG3_REG_12__SCAN_IN;
  assign n10346 = ~n10684 | ~n16940;
  assign n10351 = ~n10347 | ~n10346;
  assign n10349 = ~n10481 | ~P2_REG2_REG_12__SCAN_IN;
  assign n10348 = ~n10777 | ~P2_REG1_REG_12__SCAN_IN;
  assign n10350 = ~n10349 | ~n10348;
  assign n10353 = ~n16592;
  assign n10931 = n17505 | n10353;
  assign n16931 = n16955 | n10921;
  assign n10352 = n10931 & n16931;
  assign n10932 = ~n17505 | ~n10353;
  assign n10359 = ~n12395 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n10358 = ~n11975 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n10360 = ~SI_13_;
  assign n10381 = ~n10361 | ~n10360;
  assign n10362 = ~n10361;
  assign n10363 = ~n10362 | ~SI_13_;
  assign n10378 = ~n10381 | ~n10363;
  assign n10364 = ~n10385 | ~P2_IR_REG_31__SCAN_IN;
  assign n16817 = ~n10364 ^ P2_IR_REG_13__SCAN_IN;
  assign n10367 = ~n16817 | ~n12102;
  assign n10365 = ~P1_DATAO_REG_13__SCAN_IN;
  assign n10366 = n10768 | n10365;
  assign n10368 = n10367 & n10366;
  assign n10369 = ~P2_REG3_REG_12__SCAN_IN;
  assign n10370 = n10393 | n10369;
  assign n13923 = ~n10370 ^ P2_REG3_REG_13__SCAN_IN;
  assign n10372 = ~n10684 | ~n13923;
  assign n10371 = ~n10065 | ~P2_REG2_REG_13__SCAN_IN;
  assign n10376 = n10372 & n10371;
  assign n10374 = ~n8990 | ~P2_REG0_REG_13__SCAN_IN;
  assign n10373 = ~n10777 | ~P2_REG1_REG_13__SCAN_IN;
  assign n10375 = n10374 & n10373;
  assign n10377 = ~n13920 | ~n13898;
  assign n10379 = ~n10378;
  assign n10384 = ~n12395 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n10383 = ~n12394 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n10403 = ~n10384 | ~n10383;
  assign n10401 = ~n10403 ^ SI_14_;
  assign n17258 = ~n10402 ^ n10401;
  assign n10391 = n17258 | n10698;
  assign n10412 = ~n10386 | ~P2_IR_REG_31__SCAN_IN;
  assign n17259 = ~n10412 ^ P2_IR_REG_14__SCAN_IN;
  assign n10389 = ~n17259 | ~n12102;
  assign n10387 = ~P1_DATAO_REG_14__SCAN_IN;
  assign n10388 = n10768 | n10387;
  assign n10390 = n10389 & n10388;
  assign n10392 = ~P2_REG3_REG_12__SCAN_IN | ~P2_REG3_REG_13__SCAN_IN;
  assign n13910 = ~n10447 ^ P2_REG3_REG_14__SCAN_IN;
  assign n10395 = ~n10684 | ~n13910;
  assign n10394 = ~n10258 | ~P2_REG0_REG_14__SCAN_IN;
  assign n10400 = n10395 & n10394;
  assign n10398 = ~n10481 | ~P2_REG2_REG_14__SCAN_IN;
  assign n10397 = ~n10777 | ~P2_REG1_REG_14__SCAN_IN;
  assign n10399 = n10398 & n10397;
  assign n13893 = ~n14114 ^ n12005;
  assign n10404 = ~n10403 | ~SI_14_;
  assign n10406 = ~n12395 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n10405 = ~n11973 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n10407 = ~SI_15_;
  assign n10430 = ~n10408 | ~n10407;
  assign n10409 = ~n10408;
  assign n10410 = ~n10409 | ~SI_15_;
  assign n17252 = ~n10429 ^ n10428;
  assign n10419 = n17252 | n10698;
  assign n10411 = ~P2_IR_REG_14__SCAN_IN;
  assign n10413 = ~n10412 | ~n10411;
  assign n10414 = ~n10413 | ~P2_IR_REG_31__SCAN_IN;
  assign n17253 = ~n10414 ^ P2_IR_REG_15__SCAN_IN;
  assign n10417 = ~n17253 | ~n12102;
  assign n10415 = ~P1_DATAO_REG_15__SCAN_IN;
  assign n10416 = n10768 | n10415;
  assign n10418 = n10417 & n10416;
  assign n10421 = ~n8990 | ~P2_REG0_REG_15__SCAN_IN;
  assign n10420 = ~n10777 | ~P2_REG1_REG_15__SCAN_IN;
  assign n10427 = n10421 & n10420;
  assign n10422 = ~P2_REG3_REG_14__SCAN_IN;
  assign n10423 = n10447 | n10422;
  assign n13881 = ~n10423 ^ P2_REG3_REG_15__SCAN_IN;
  assign n10425 = ~n10684 | ~n13881;
  assign n10424 = ~n10065 | ~P2_REG2_REG_15__SCAN_IN;
  assign n10426 = n10425 & n10424;
  assign n10947 = ~n11093;
  assign n10432 = ~n12395 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n10431 = ~n12394 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n10461 = ~n10434 | ~n10433;
  assign n10435 = ~n10434;
  assign n10436 = ~n10435 | ~SI_16_;
  assign n10458 = ~n10461 | ~n10436;
  assign n10437 = ~P1_DATAO_REG_16__SCAN_IN;
  assign n10444 = n10768 | n10437;
  assign n10439 = ~n10438;
  assign n10442 = ~n10465 | ~P2_IR_REG_31__SCAN_IN;
  assign n17246 = ~n10442 ^ P2_IR_REG_16__SCAN_IN;
  assign n10443 = ~n12102 | ~n17246;
  assign n10445 = n10444 & n10443;
  assign n10446 = ~P2_REG3_REG_14__SCAN_IN | ~P2_REG3_REG_15__SCAN_IN;
  assign n13856 = ~n10498 ^ P2_REG3_REG_16__SCAN_IN;
  assign n10449 = ~n10684 | ~n13856;
  assign n10448 = ~n8990 | ~P2_REG0_REG_16__SCAN_IN;
  assign n10453 = n10449 & n10448;
  assign n10451 = ~n10065 | ~P2_REG2_REG_16__SCAN_IN;
  assign n10450 = ~n10777 | ~P2_REG1_REG_16__SCAN_IN;
  assign n10452 = n10451 & n10450;
  assign n10456 = ~n13384 | ~n13871;
  assign n13830 = ~n14114 & ~n12005;
  assign n10454 = ~n11093 | ~n13830;
  assign n10455 = n10454 & n13833;
  assign n10457 = ~n14091 | ~n13806;
  assign n10459 = ~n10458;
  assign n10463 = ~n12395 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n10462 = ~n11975 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n10488 = ~n10463 | ~n10462;
  assign n10464 = ~P1_DATAO_REG_17__SCAN_IN;
  assign n10474 = n10768 | n10464;
  assign n10466 = ~P2_IR_REG_16__SCAN_IN;
  assign n10472 = ~n10522;
  assign n10468 = ~n10467 | ~P2_IR_REG_31__SCAN_IN;
  assign n10470 = ~n10468 | ~P2_IR_REG_17__SCAN_IN;
  assign n10469 = ~n9322 | ~P2_IR_REG_31__SCAN_IN;
  assign n10471 = ~n10470 | ~n10469;
  assign n10473 = ~n12102 | ~n17239;
  assign n10475 = n10474 & n10473;
  assign n10476 = ~P2_REG3_REG_16__SCAN_IN;
  assign n10478 = ~n10498 & ~n10476;
  assign n10477 = ~P2_REG3_REG_17__SCAN_IN;
  assign n13818 = ~n10478 ^ n10477;
  assign n10480 = ~n10684 | ~n13818;
  assign n10479 = ~n8990 | ~P2_REG0_REG_17__SCAN_IN;
  assign n10485 = ~n10480 | ~n10479;
  assign n10483 = ~n10481 | ~P2_REG2_REG_17__SCAN_IN;
  assign n10482 = ~n10777 | ~P2_REG1_REG_17__SCAN_IN;
  assign n10484 = ~n10483 | ~n10482;
  assign n10487 = ~n13813 | ~n13838;
  assign n13778 = ~n13838;
  assign n10486 = ~n13279 | ~n13778;
  assign n10490 = ~n12395 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n10489 = ~n11973 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n10512 = ~n10490 | ~n10489;
  assign n10509 = ~n10512 ^ SI_18_;
  assign n16131 = ~n10511 ^ n10509;
  assign n10496 = ~n16131 | ~n10732;
  assign n10491 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n10494 = n10768 | n10491;
  assign n10492 = n10522 | n10523;
  assign n16916 = ~n10492 ^ P2_IR_REG_18__SCAN_IN;
  assign n10493 = ~n16916 | ~n12102;
  assign n10495 = n10494 & n10493;
  assign n10497 = ~P2_REG3_REG_16__SCAN_IN | ~P2_REG3_REG_17__SCAN_IN;
  assign n10532 = ~n10498 & ~n10497;
  assign n10499 = ~n10532;
  assign n13789 = ~n10499 ^ P2_REG3_REG_18__SCAN_IN;
  assign n10501 = ~n13789 | ~n10684;
  assign n10500 = ~n10481 | ~P2_REG2_REG_18__SCAN_IN;
  assign n10505 = ~n10501 | ~n10500;
  assign n10503 = ~n8990 | ~P2_REG0_REG_18__SCAN_IN;
  assign n10502 = ~n10777 | ~P2_REG1_REG_18__SCAN_IN;
  assign n10504 = ~n10503 | ~n10502;
  assign n10506 = n14071 | n13805;
  assign n10507 = ~n14071 | ~n13805;
  assign n13749 = ~n10508 | ~n10507;
  assign n10510 = ~n10509;
  assign n10513 = ~n10512 | ~SI_18_;
  assign n10516 = ~n12395 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n10515 = ~n12394 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n10538 = ~n10518 | ~n10517;
  assign n10519 = ~n10518;
  assign n10520 = ~n10519 | ~SI_19_;
  assign n10537 = ~n10538 | ~n10520;
  assign n10526 = n17227 | n12110;
  assign n10524 = ~P1_DATAO_REG_19__SCAN_IN;
  assign n10525 = n10768 | n10524;
  assign n10527 = n10526 & n10525;
  assign n10529 = ~n10481 | ~P2_REG2_REG_19__SCAN_IN;
  assign n10528 = ~n10777 | ~P2_REG1_REG_19__SCAN_IN;
  assign n10531 = ~n10529 | ~n10528;
  assign n10530 = n8990 & P2_REG0_REG_19__SCAN_IN;
  assign n10535 = ~n10531 & ~n10530;
  assign n13766 = ~n10552 ^ P2_REG3_REG_19__SCAN_IN;
  assign n10533 = ~n10684;
  assign n10534 = n13766 | n10533;
  assign n17558 = ~n10535 | ~n10534;
  assign n13777 = ~n17558;
  assign n11112 = n14060 | n13777;
  assign n11111 = ~n14060 | ~n13777;
  assign n10541 = ~n12395 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n10540 = ~n12394 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n10544 = ~n10543;
  assign n10545 = ~n10544 | ~SI_20_;
  assign n10547 = ~n10562 | ~n10545;
  assign n10549 = ~n10546 | ~n10547;
  assign n10548 = ~n10547;
  assign n10551 = ~n12299 | ~n10732;
  assign n12197 = ~P1_DATAO_REG_20__SCAN_IN;
  assign n10550 = n10768 | n12197;
  assign n10553 = ~n10569;
  assign n13738 = ~P2_REG3_REG_20__SCAN_IN ^ n10553;
  assign n10555 = ~n10684 | ~n13738;
  assign n10554 = ~n10777 | ~P2_REG1_REG_20__SCAN_IN;
  assign n10559 = ~n10555 | ~n10554;
  assign n10557 = ~n8990 | ~P2_REG0_REG_20__SCAN_IN;
  assign n10556 = ~n10481 | ~P2_REG2_REG_20__SCAN_IN;
  assign n10558 = ~n10557 | ~n10556;
  assign n13752 = ~n17561;
  assign n10560 = n14049 | n13752;
  assign n10561 = ~n14049 | ~n13752;
  assign n10565 = ~n12395 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n10564 = ~n11973 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n10585 = ~n10565 | ~n10564;
  assign n10604 = ~n10585 ^ SI_21_;
  assign n10568 = n12322 | n10698;
  assign n10566 = ~P1_DATAO_REG_21__SCAN_IN;
  assign n10567 = n10768 | n10566;
  assign n14038 = ~n10568 | ~n10567;
  assign n10570 = ~n10595;
  assign n13715 = ~P2_REG3_REG_21__SCAN_IN ^ n10570;
  assign n10572 = ~n10684 | ~n13715;
  assign n10571 = ~n10777 | ~P2_REG1_REG_21__SCAN_IN;
  assign n10576 = ~n10572 | ~n10571;
  assign n10574 = ~n8990 | ~P2_REG0_REG_21__SCAN_IN;
  assign n10573 = ~n10065 | ~P2_REG2_REG_21__SCAN_IN;
  assign n10575 = ~n10574 | ~n10573;
  assign n10577 = ~n13714 | ~n17564;
  assign n13729 = ~n17564;
  assign n10578 = ~n14038 | ~n13729;
  assign n10580 = ~n12395 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n10579 = ~n11973 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n10603 = ~n10582 | ~n10581;
  assign n10583 = ~n10582;
  assign n10584 = ~n10583 | ~SI_22_;
  assign n10588 = n10603 & n10584;
  assign n10586 = ~n10585 | ~SI_21_;
  assign n10592 = ~n10587 | ~n10605;
  assign n10590 = ~n10587 | ~n10586;
  assign n10589 = ~n10588;
  assign n10591 = ~n10590 | ~n10589;
  assign n11769 = ~n10592 | ~n10591;
  assign n10594 = ~n11769 | ~n10732;
  assign n12358 = ~P1_DATAO_REG_22__SCAN_IN;
  assign n10593 = n10768 | n12358;
  assign n13691 = P2_REG3_REG_22__SCAN_IN ^ n10622;
  assign n10601 = ~n13691 | ~n10684;
  assign n10597 = ~n10065 | ~P2_REG2_REG_22__SCAN_IN;
  assign n10596 = ~n10777 | ~P2_REG1_REG_22__SCAN_IN;
  assign n10599 = ~n10597 | ~n10596;
  assign n10598 = n8990 & P2_REG0_REG_22__SCAN_IN;
  assign n10600 = ~n10599 & ~n10598;
  assign n17567 = ~n10601 | ~n10600;
  assign n13656 = ~n17567;
  assign n10602 = ~n13680;
  assign n10606 = ~n10603;
  assign n10615 = ~n10606 & ~n10605;
  assign n10613 = n10618 | n10615;
  assign n10608 = ~n12395 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n10607 = ~n11973 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n10609 = ~SI_23_;
  assign n10644 = ~n10610 | ~n10609;
  assign n10611 = ~n10610;
  assign n10612 = ~n10611 | ~SI_23_;
  assign n10614 = ~n10644 | ~n10612;
  assign n10619 = ~n10613 | ~n10614;
  assign n10617 = ~n10614;
  assign n10616 = ~n10615;
  assign n10649 = ~n10617 | ~n10616;
  assign n10621 = ~n12334 | ~n10732;
  assign n12336 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n10620 = n10768 | n12336;
  assign n13667 = P2_REG3_REG_23__SCAN_IN ^ n10635;
  assign n10628 = ~n13667 | ~n10684;
  assign n10624 = ~n8990 | ~P2_REG0_REG_23__SCAN_IN;
  assign n10623 = ~n10481 | ~P2_REG2_REG_23__SCAN_IN;
  assign n10626 = ~n10624 | ~n10623;
  assign n10625 = n10777 & P2_REG1_REG_23__SCAN_IN;
  assign n10627 = ~n10626 & ~n10625;
  assign n17570 = ~n10628 | ~n10627;
  assign n13408 = ~n17570;
  assign n11014 = n14017 | n13408;
  assign n11015 = ~n14017 | ~n13408;
  assign n10632 = ~n10629 | ~n10644;
  assign n10631 = ~n12395 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n10630 = ~n12394 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n10653 = ~n10631 | ~n10630;
  assign n10643 = ~n10653 ^ SI_24_;
  assign n14226 = ~n10632 ^ n10643;
  assign n10634 = n14226 | n10698;
  assign n14228 = ~P1_DATAO_REG_24__SCAN_IN;
  assign n10633 = n10768 | n14228;
  assign n10636 = ~P2_REG3_REG_24__SCAN_IN;
  assign n13645 = ~n10664 ^ n10636;
  assign n10642 = ~n13645 | ~n10684;
  assign n10638 = ~n10481 | ~P2_REG2_REG_24__SCAN_IN;
  assign n10637 = ~n10777 | ~P2_REG1_REG_24__SCAN_IN;
  assign n10640 = ~n10638 | ~n10637;
  assign n10639 = n8990 & P2_REG0_REG_24__SCAN_IN;
  assign n10641 = ~n10640 & ~n10639;
  assign n17573 = ~n10642 | ~n10641;
  assign n11022 = ~n13644 | ~n17573;
  assign n13655 = ~n17573;
  assign n11023 = ~n14006 | ~n13655;
  assign n13246 = ~n11022 | ~n11023;
  assign n10645 = ~n10643;
  assign n10646 = ~n10650;
  assign n10655 = ~n12395 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n10654 = ~n11975 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n10656 = ~SI_25_;
  assign n10671 = ~n10657 | ~n10656;
  assign n10658 = ~n10657;
  assign n10659 = ~n10658 | ~SI_25_;
  assign n12340 = ~P1_DATAO_REG_25__SCAN_IN;
  assign n10662 = n10768 | n12340;
  assign n13623 = P2_REG3_REG_25__SCAN_IN ^ n10683;
  assign n10670 = ~n13623 | ~n10684;
  assign n10666 = ~n10777 | ~P2_REG1_REG_25__SCAN_IN;
  assign n10665 = ~n8990 | ~P2_REG0_REG_25__SCAN_IN;
  assign n10668 = ~n10666 | ~n10665;
  assign n10667 = n10481 & P2_REG2_REG_25__SCAN_IN;
  assign n10669 = ~n10668 & ~n10667;
  assign n17576 = ~n10670 | ~n10669;
  assign n13249 = ~n17576;
  assign n11033 = ~n13995 | ~n13249;
  assign n10673 = ~n12395 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n10672 = ~n11973 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n10674 = ~SI_26_;
  assign n10724 = ~n10675 | ~n10674;
  assign n10676 = ~n10675;
  assign n10677 = ~n10676 | ~SI_26_;
  assign n10679 = ~n10724 | ~n10677;
  assign n10680 = ~n10678 | ~n10679;
  assign n10714 = ~n10679;
  assign n10682 = ~n15309 | ~n10732;
  assign n14221 = ~P1_DATAO_REG_26__SCAN_IN;
  assign n10681 = n10768 | n14221;
  assign n13478 = ~P2_REG3_REG_26__SCAN_IN;
  assign n13476 = ~n10702 ^ n13478;
  assign n10690 = ~n13476 | ~n10684;
  assign n10686 = ~n10481 | ~P2_REG2_REG_26__SCAN_IN;
  assign n10685 = ~n8990 | ~P2_REG0_REG_26__SCAN_IN;
  assign n10688 = ~n10686 | ~n10685;
  assign n10687 = n10777 & P2_REG1_REG_26__SCAN_IN;
  assign n10689 = ~n10688 & ~n10687;
  assign n17579 = ~n10690 | ~n10689;
  assign n13251 = ~n17579;
  assign n11089 = ~n13984 | ~n13251;
  assign n10697 = ~n10726 | ~n10724;
  assign n10692 = ~n12395 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n10691 = ~n11973 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n10693 = ~SI_27_;
  assign n10722 = ~n10694 | ~n10693;
  assign n10695 = ~n10694;
  assign n10696 = ~n10695 | ~SI_27_;
  assign n10707 = ~n10722 | ~n10696;
  assign n14215 = ~P1_DATAO_REG_27__SCAN_IN;
  assign n10699 = n10768 | n14215;
  assign n10701 = ~n8990 | ~P2_REG0_REG_27__SCAN_IN;
  assign n10700 = ~n10777 | ~P2_REG1_REG_27__SCAN_IN;
  assign n10706 = ~n10701 | ~n10700;
  assign n10737 = ~n10702 | ~P2_REG3_REG_26__SCAN_IN;
  assign n13573 = ~P2_REG3_REG_27__SCAN_IN ^ n10737;
  assign n10704 = ~n10684 | ~n13573;
  assign n10703 = ~n10481 | ~P2_REG2_REG_27__SCAN_IN;
  assign n10705 = ~n10704 | ~n10703;
  assign n11051 = ~n13974 | ~n13255;
  assign n13560 = ~n11050 | ~n11051;
  assign n10728 = ~n10707;
  assign n10709 = ~n12395 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n10708 = ~n12394 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n10710 = ~SI_28_;
  assign n10746 = ~n10711 | ~n10710;
  assign n10712 = ~n10711;
  assign n10713 = ~n10712 | ~SI_28_;
  assign n10715 = n10714 & n10717;
  assign n10718 = ~n10717;
  assign n10721 = n10718 | n10724;
  assign n10723 = ~n10719;
  assign n10727 = n10723 & n10722;
  assign n10725 = n10724 & n10727;
  assign n10731 = ~n10726 | ~n10725;
  assign n10729 = ~n10727;
  assign n10730 = n10729 | n10728;
  assign n10735 = ~n14208 | ~n10732;
  assign n10733 = ~P1_DATAO_REG_28__SCAN_IN;
  assign n10734 = n10768 | n10733;
  assign n10736 = ~P2_REG3_REG_27__SCAN_IN;
  assign n10754 = ~n10737 & ~n10736;
  assign n10738 = ~n10754;
  assign n13547 = ~P2_REG3_REG_28__SCAN_IN ^ n10738;
  assign n10740 = ~n10684 | ~n13547;
  assign n10739 = ~n8990 | ~P2_REG0_REG_28__SCAN_IN;
  assign n10744 = ~n10740 | ~n10739;
  assign n10742 = ~n10481 | ~P2_REG2_REG_28__SCAN_IN;
  assign n10741 = ~n10777 | ~P2_REG1_REG_28__SCAN_IN;
  assign n10743 = ~n10742 | ~n10741;
  assign n11087 = ~n13964 | ~n13274;
  assign n10749 = ~n12395 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n10748 = ~n12394 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n10761 = ~n10749 | ~n10748;
  assign n10750 = ~n10761 ^ SI_29_;
  assign n14202 = ~n10760 ^ n10750;
  assign n14203 = ~P1_DATAO_REG_29__SCAN_IN;
  assign n10751 = n10768 | n14203;
  assign n10753 = ~n10065 | ~P2_REG2_REG_29__SCAN_IN;
  assign n10752 = ~n10777 | ~P2_REG1_REG_29__SCAN_IN;
  assign n10759 = ~n10753 | ~n10752;
  assign n10757 = ~n8990 | ~P2_REG0_REG_29__SCAN_IN;
  assign n13532 = ~n10754 | ~P2_REG3_REG_28__SCAN_IN;
  assign n10755 = ~n13532;
  assign n10756 = ~n10684 | ~n10755;
  assign n10758 = ~n10757 | ~n10756;
  assign n10762 = ~n10761 | ~SI_29_;
  assign n10765 = ~n12395 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n10764 = ~n12394 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n10799 = ~n10765 | ~n10764;
  assign n10766 = ~SI_30_;
  assign n10767 = ~n10799 ^ n10766;
  assign n14195 = ~n10803 ^ n10767;
  assign n10770 = n14195 | n10698;
  assign n14197 = ~P1_DATAO_REG_30__SCAN_IN;
  assign n10769 = n10768 | n14197;
  assign n13506 = ~n10770 | ~n10769;
  assign n10772 = ~n10777 | ~P2_REG1_REG_30__SCAN_IN;
  assign n10771 = ~n8990 | ~P2_REG0_REG_30__SCAN_IN;
  assign n10774 = ~n10772 | ~n10771;
  assign n10773 = n10481 & P2_REG2_REG_30__SCAN_IN;
  assign n17591 = n10774 | n10773;
  assign n13273 = ~n17591;
  assign n10776 = ~n10481 | ~P2_REG2_REG_31__SCAN_IN;
  assign n10775 = ~n8990 | ~P2_REG0_REG_31__SCAN_IN;
  assign n10779 = ~n10776 | ~n10775;
  assign n10778 = n10777 & P2_REG1_REG_31__SCAN_IN;
  assign n13514 = ~n17595;
  assign n12424 = ~n10782 ^ n10816;
  assign n12423 = ~n12424;
  assign n10806 = ~n13514 | ~n12423;
  assign n10784 = ~n11073 | ~n10806;
  assign n10783 = ~n11069;
  assign n10786 = ~n12395 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n10785 = ~n11973 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n10788 = ~n10786 | ~n10785;
  assign n10787 = ~SI_31_;
  assign n10791 = ~n10788 ^ n10787;
  assign n10789 = ~n10799 | ~SI_30_;
  assign n10790 = ~n10791 | ~n10789;
  assign n10798 = n10803 | n10790;
  assign n10801 = ~n10791;
  assign n10792 = ~n10801 | ~SI_30_;
  assign n10796 = ~n10792 | ~n10799;
  assign n10794 = n10801 | SI_30_;
  assign n10793 = ~n10799;
  assign n10795 = ~n10794 | ~n10793;
  assign n10797 = ~n10796 | ~n10795;
  assign n10800 = n10799 | SI_30_;
  assign n10802 = n10801 & n10800;
  assign n10804 = ~n10803 | ~n10802;
  assign n10805 = ~n11973 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n11078 = ~n13945 | ~n17595;
  assign n10808 = ~n11078;
  assign n10807 = ~n13953 & ~n10806;
  assign n10809 = ~n10808 & ~n10807;
  assign n11074 = ~n13506 | ~n13273;
  assign n10810 = ~n11077;
  assign n10829 = n12424 | n17098;
  assign n10813 = ~n10812 | ~n10811;
  assign n10820 = n10829 | n13537;
  assign n11124 = ~n10817 | ~n10816;
  assign n12431 = ~n8996 | ~n17227;
  assign n10821 = ~n10820 | ~n12487;
  assign n10823 = ~n10027 & ~n17373;
  assign n17365 = ~n16568;
  assign n16570 = ~n11988 | ~n17365;
  assign n17163 = ~n10027 | ~n17373;
  assign n10827 = ~n17163 | ~n11063;
  assign n10830 = ~n10828 & ~n17365;
  assign n10832 = ~n13260 | ~n10829;
  assign n10831 = ~n10830 & ~n10832;
  assign n10835 = ~n10831 & ~n11988;
  assign n10833 = ~n10832;
  assign n10834 = ~n10833 & ~n17365;
  assign n10842 = ~n10837 | ~n10836;
  assign n10839 = ~n10828 | ~n10027;
  assign n10838 = ~n11063 | ~n12429;
  assign n10840 = ~n10839 | ~n10838;
  assign n17170 = ~n10027 | ~n12429;
  assign n10841 = ~n10840 | ~n17170;
  assign n10846 = ~n10842 | ~n10841;
  assign n10844 = ~n11094 | ~n11063;
  assign n10843 = ~n10828 | ~n11095;
  assign n10845 = ~n10844 | ~n10843;
  assign n10850 = ~n10846 | ~n10845;
  assign n10848 = ~n11094 | ~n10828;
  assign n10847 = ~n11095 | ~n11063;
  assign n10849 = ~n10848 | ~n10847;
  assign n10852 = ~n10828 & ~n16541;
  assign n10851 = ~n11063 & ~n17399;
  assign n10861 = ~n10852 & ~n10851;
  assign n10859 = ~n10865 & ~n10861;
  assign n10854 = ~n10828 | ~n17133;
  assign n10853 = ~n10866 | ~n11063;
  assign n10868 = ~n10854 | ~n10853;
  assign n13212 = ~n10866 | ~n17133;
  assign n10860 = ~n10868 | ~n13212;
  assign n16603 = ~n16541;
  assign n10856 = ~n10828 | ~n16603;
  assign n10855 = ~n11063 | ~n17141;
  assign n10857 = ~n10856 | ~n10855;
  assign n10858 = ~n10860 | ~n10857;
  assign n10863 = ~n10860;
  assign n10862 = ~n10861;
  assign n10864 = ~n10863 & ~n10862;
  assign n10867 = ~n10866 & ~n17133;
  assign n10872 = ~n10868 & ~n10867;
  assign n10870 = ~n11097 | ~n10828;
  assign n10869 = ~n11096 | ~n11063;
  assign n10871 = n10870 & n10869;
  assign n10874 = ~n17067 | ~n11063;
  assign n10873 = ~n10828 | ~n16516;
  assign n10880 = n10874 & n10873;
  assign n12459 = ~n16516;
  assign n10875 = ~n12459 | ~n17432;
  assign n10879 = ~n10880 | ~n10875;
  assign n10877 = ~n11097 | ~n11063;
  assign n10876 = ~n10828 | ~n11096;
  assign n10878 = ~n10877 | ~n10876;
  assign n10881 = ~n10880;
  assign n13217 = ~n17067 | ~n16516;
  assign n10882 = ~n10881 | ~n13217;
  assign n10883 = n10882 & n10889;
  assign n10884 = ~n10883 | ~n10890;
  assign n10886 = n17041 | n10828;
  assign n10885 = ~n10828 | ~n16435;
  assign n10897 = n10886 & n10885;
  assign n10887 = ~n16435 | ~n11063;
  assign n10896 = ~n10888 | ~n10887;
  assign n10894 = ~n10897 | ~n10896;
  assign n10892 = ~n10889 | ~n10828;
  assign n10891 = ~n10890 | ~n11063;
  assign n10893 = ~n10892 | ~n10891;
  assign n10895 = ~n10894 | ~n10893;
  assign n10898 = ~n10897 & ~n10896;
  assign n10900 = ~n17476 & ~n10828;
  assign n10899 = ~n11063 & ~n16559;
  assign n10910 = ~n10900 & ~n10899;
  assign n13223 = ~n17476 | ~n16559;
  assign n10904 = ~n10910 | ~n13223;
  assign n10902 = ~n10913 | ~n10828;
  assign n10901 = ~n16991 | ~n11063;
  assign n10903 = ~n10902 | ~n10901;
  assign n10914 = ~n10904 | ~n10903;
  assign n16442 = ~n17476;
  assign n10906 = ~n10910 & ~n16442;
  assign n10907 = ~n10906 & ~n11063;
  assign n10909 = ~n10907 | ~n11105;
  assign n10908 = ~n10914 & ~n16991;
  assign n10918 = ~n10909 & ~n10908;
  assign n10911 = ~n10910 & ~n16591;
  assign n10912 = ~n10911 & ~n10828;
  assign n10916 = ~n10912 | ~n16931;
  assign n10915 = ~n10914 & ~n10913;
  assign n10917 = ~n10916 & ~n10915;
  assign n10919 = ~n10918 & ~n10917;
  assign n10927 = ~n10920 & ~n10919;
  assign n10923 = ~n16955 & ~n11063;
  assign n10922 = ~n16505 & ~n10828;
  assign n10925 = ~n10923 & ~n10922;
  assign n10924 = ~n16955 & ~n16505;
  assign n10926 = ~n10925 & ~n10924;
  assign n10929 = ~n10931 | ~n11063;
  assign n10928 = ~n10932 | ~n10828;
  assign n10930 = ~n10929 | ~n10928;
  assign n10934 = ~n10931 | ~n10828;
  assign n10933 = ~n10932 | ~n11063;
  assign n10935 = ~n10934 | ~n10933;
  assign n14125 = ~n13920;
  assign n10937 = ~n14125 | ~n11063;
  assign n10936 = ~n10828 | ~n13898;
  assign n10939 = ~n14125 | ~n10828;
  assign n10938 = ~n13898 | ~n11063;
  assign n10940 = ~n10939 | ~n10938;
  assign n10942 = n14114 | n11063;
  assign n10941 = ~n12005 | ~n11063;
  assign n10951 = n10942 & n10941;
  assign n10944 = n14114 | n10828;
  assign n10943 = ~n10828 | ~n12005;
  assign n10950 = ~n10944 | ~n10943;
  assign n10945 = ~n10951 | ~n10950;
  assign n10946 = ~n13833;
  assign n10949 = ~n10946 & ~n11063;
  assign n10948 = ~n10947 & ~n10828;
  assign n10953 = ~n10949 & ~n10948;
  assign n10952 = ~n10951 & ~n10950;
  assign n10954 = ~n10953 & ~n10952;
  assign n10959 = ~n10955 | ~n10954;
  assign n10957 = ~n13833 | ~n11063;
  assign n10956 = ~n11093 | ~n10828;
  assign n10958 = ~n10957 | ~n10956;
  assign n10965 = ~n10959 | ~n10958;
  assign n10961 = ~n14091 & ~n10828;
  assign n10960 = ~n13871 & ~n11063;
  assign n10967 = ~n10961 & ~n10960;
  assign n10963 = ~n13384 | ~n10828;
  assign n10962 = ~n13806 | ~n11063;
  assign n10966 = ~n10963 | ~n10962;
  assign n10964 = ~n10967 & ~n10966;
  assign n10969 = ~n10966;
  assign n10968 = ~n10967;
  assign n10970 = ~n10969 & ~n10968;
  assign n10972 = ~n13813 | ~n11063;
  assign n10971 = ~n10828 | ~n13778;
  assign n10975 = n10972 & n10971;
  assign n10973 = ~n13279 | ~n13838;
  assign n10974 = ~n10975 | ~n10973;
  assign n10976 = ~n10975;
  assign n13235 = ~n13813 | ~n13778;
  assign n10977 = ~n10976 | ~n13235;
  assign n10979 = n14071 | n10828;
  assign n10978 = ~n10828 | ~n13805;
  assign n10983 = n10979 & n10978;
  assign n10981 = n14071 | n11063;
  assign n10980 = ~n13805 | ~n11063;
  assign n10982 = ~n10981 | ~n10980;
  assign n10985 = ~n10982;
  assign n10984 = ~n10983;
  assign n10987 = ~n11112 | ~n11063;
  assign n10986 = ~n11111 | ~n10828;
  assign n10989 = n14049 | n11063;
  assign n10988 = ~n13752 | ~n11063;
  assign n10994 = ~n10989 | ~n10988;
  assign n11091 = n14049 | n17561;
  assign n10993 = ~n10994 | ~n11091;
  assign n10991 = ~n11112 | ~n10828;
  assign n10990 = ~n11111 | ~n11063;
  assign n10992 = ~n10991 | ~n10990;
  assign n13240 = ~n14049 | ~n17561;
  assign n10995 = ~n13240;
  assign n10997 = ~n14038 & ~n11063;
  assign n10996 = ~n10828 & ~n17564;
  assign n11003 = ~n10997 & ~n10996;
  assign n13241 = ~n14038 | ~n17564;
  assign n10998 = ~n11003 | ~n13241;
  assign n11002 = ~n10999 | ~n10828;
  assign n11001 = ~n11000 | ~n11063;
  assign n11006 = ~n11002 | ~n11001;
  assign n11004 = ~n11003;
  assign n13242 = ~n13714 | ~n13729;
  assign n11005 = ~n11004 | ~n13242;
  assign n11007 = n11006 & n11005;
  assign n11010 = ~n11008 | ~n10828;
  assign n11009 = ~n17567 | ~n11063;
  assign n11012 = ~n11010 | ~n11009;
  assign n11011 = ~n11008 | ~n17567;
  assign n11013 = ~n11012 | ~n11011;
  assign n11017 = ~n11014 | ~n10828;
  assign n11016 = ~n11015 | ~n11063;
  assign n11019 = ~n14017 | ~n10828;
  assign n11018 = ~n17570 | ~n11063;
  assign n11020 = ~n11019 | ~n11018;
  assign n13245 = ~n14017 | ~n17570;
  assign n11021 = ~n11020 | ~n13245;
  assign n11025 = ~n11022 | ~n10828;
  assign n11024 = ~n11023 | ~n11063;
  assign n11026 = ~n11025 | ~n11024;
  assign n11028 = ~n14006 | ~n10828;
  assign n11027 = ~n17573 | ~n11063;
  assign n11030 = ~n11028 | ~n11027;
  assign n11029 = ~n14006 | ~n17573;
  assign n11035 = ~n11032 | ~n10828;
  assign n11034 = ~n11033 | ~n11063;
  assign n11036 = ~n11035 | ~n11034;
  assign n11038 = ~n13995 | ~n10828;
  assign n11037 = ~n17576 | ~n11063;
  assign n11040 = ~n11038 | ~n11037;
  assign n11039 = ~n13995 | ~n17576;
  assign n11041 = ~n11040 | ~n11039;
  assign n11043 = ~n11090 | ~n10828;
  assign n11042 = ~n11089 | ~n11063;
  assign n11044 = ~n11043 | ~n11042;
  assign n11046 = ~n13984 | ~n10828;
  assign n11045 = ~n17579 | ~n11063;
  assign n11048 = ~n11046 | ~n11045;
  assign n11047 = ~n13984 | ~n17579;
  assign n11053 = ~n11050 | ~n10828;
  assign n11052 = ~n11051 | ~n11063;
  assign n11054 = ~n11053 | ~n11052;
  assign n11056 = ~n13974 | ~n10828;
  assign n11055 = ~n11063 | ~n17582;
  assign n11058 = ~n11056 | ~n11055;
  assign n11057 = ~n13974 | ~n17582;
  assign n11059 = ~n11058 | ~n11057;
  assign n11061 = ~n11088 | ~n10828;
  assign n11060 = ~n11087 | ~n11063;
  assign n11062 = ~n11061 | ~n11060;
  assign n11065 = ~n13964 | ~n10828;
  assign n11064 = ~n11063 | ~n17585;
  assign n11067 = ~n11065 | ~n11064;
  assign n11066 = ~n13964 | ~n17585;
  assign n11071 = ~n11068 & ~n11063;
  assign n11070 = ~n11069 & ~n10828;
  assign n11076 = ~n11078 | ~n10828;
  assign n11075 = ~n11074;
  assign n11080 = ~n11077 | ~n10828;
  assign n11079 = ~n11078 | ~n11063;
  assign n11081 = ~n11080 | ~n11079;
  assign n13269 = n10825 | n17227;
  assign n11083 = ~n13269;
  assign n11084 = ~n11083 & ~n11082;
  assign n12580 = ~n13537;
  assign n11086 = ~n13945 ^ n13514;
  assign n13267 = ~n13280 ^ n17588;
  assign n11117 = n11086 & n13267;
  assign n13555 = ~n11088 | ~n11087;
  assign n13587 = ~n11090 | ~n11089;
  assign n13250 = ~n13587;
  assign n13727 = ~n11091 | ~n13240;
  assign n11092 = ~n13384 | ~n13806;
  assign n13232 = ~n14091 | ~n13871;
  assign n11098 = n13204 | n17363;
  assign n17106 = ~n11097 | ~n11096;
  assign n11099 = ~n11098 & ~n17106;
  assign n13211 = ~n16517 ^ n17133;
  assign n17117 = ~n13211;
  assign n17198 = ~n12430 ^ n12429;
  assign n17148 = ~n16541 ^ n17141;
  assign n11100 = ~n17198 & ~n17148;
  assign n11102 = ~n11101 & ~n17081;
  assign n11103 = ~n11102 | ~n17033;
  assign n17058 = ~n17443 ^ n12026;
  assign n11104 = ~n11103 & ~n17058;
  assign n17015 = ~n17465 ^ n16477;
  assign n16963 = ~n16931 | ~n11105;
  assign n16934 = ~n17505 ^ n16592;
  assign n11107 = n11106 | n13933;
  assign n11108 = ~n13832 & ~n11107;
  assign n11109 = ~n11108 | ~n9952;
  assign n11113 = n13727 & n11110;
  assign n13750 = ~n11112 | ~n11111;
  assign n13775 = ~n14071 ^ n13805;
  assign n13703 = ~n14038 ^ n17564;
  assign n11116 = ~n13555 & ~n11115;
  assign n11118 = ~n12580 | ~n17098;
  assign n12595 = ~n13537 | ~n17227;
  assign n11120 = ~n12595 | ~n12424;
  assign n11121 = ~n9005 & ~n11120;
  assign n12335 = n12588 | P2_U3152;
  assign n11127 = ~n10825;
  assign n11128 = ~P2_U3152 & ~n11127;
  assign n11153 = ~n11128 & ~n12588;
  assign n11131 = ~n11130 | ~n11129;
  assign n11135 = ~n11143;
  assign n11136 = ~n11135 | ~n11144;
  assign n11137 = ~n11136 | ~P2_IR_REG_31__SCAN_IN;
  assign n11140 = ~n11137 | ~P2_IR_REG_26__SCAN_IN;
  assign n11139 = ~n11138 | ~P2_IR_REG_31__SCAN_IN;
  assign n11141 = ~n11140 | ~n11139;
  assign n11146 = ~n14220 & ~n12569;
  assign n12101 = ~n17225;
  assign n12598 = ~n11147;
  assign n11148 = ~n12595 & ~n14214;
  assign n11149 = ~n16626 | ~n11148;
  assign n11151 = ~n12101 & ~n11149;
  assign n11150 = ~n12588;
  assign n11152 = ~n11151 & ~n11150;
  assign n11154 = ~n11153 & ~n11152;
  assign n13271 = ~P2_B_REG_SCAN_IN;
  assign P2_U3244 = ~n11155 | ~n9963;
  assign n11157 = ~P1_IR_REG_6__SCAN_IN & ~P1_IR_REG_10__SCAN_IN;
  assign n11156 = ~P1_IR_REG_9__SCAN_IN & ~P1_IR_REG_11__SCAN_IN;
  assign n11161 = ~n11157 | ~n11156;
  assign n11160 = ~n11159 | ~n11158;
  assign n11337 = n11251 & n9192;
  assign n11210 = n11162 & n11337;
  assign n11170 = ~n11175;
  assign n11171 = ~n11658 | ~n11170;
  assign n11173 = ~n11171 | ~P1_IR_REG_31__SCAN_IN;
  assign n11186 = ~n12329;
  assign n11174 = ~P1_IR_REG_16__SCAN_IN & ~P1_IR_REG_23__SCAN_IN;
  assign n11183 = ~n11543 | ~n11211;
  assign n11178 = ~n11183;
  assign n11177 = ~P1_IR_REG_24__SCAN_IN;
  assign n11179 = ~n11178 | ~n11177;
  assign n11180 = ~n11182 | ~n11205;
  assign n15310 = ~n11181 ^ P1_IR_REG_26__SCAN_IN;
  assign n11184 = ~n11183 | ~P1_IR_REG_31__SCAN_IN;
  assign P1_U3084 = ~P1_STATE_REG_SCAN_IN;
  assign n11189 = ~P1_IR_REG_17__SCAN_IN & ~P1_IR_REG_16__SCAN_IN;
  assign n11192 = ~n11201 | ~n11203;
  assign n11193 = ~n11200 | ~n11199;
  assign n11197 = ~P1_IR_REG_19__SCAN_IN;
  assign n16125 = ~n11198 ^ n11197;
  assign n11202 = ~n11201;
  assign n11206 = ~P1_IR_REG_26__SCAN_IN & ~P1_IR_REG_24__SCAN_IN;
  assign n11207 = n11206 & n11205;
  assign n11209 = n11208 & n11207;
  assign n15494 = ~n11216 ^ n11215;
  assign n11218 = ~n15309 | ~n11825;
  assign n12402 = ~n11263 | ~n10357;
  assign n15312 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n11217 = n12402 | n15312;
  assign n14622 = ~n15047;
  assign n11359 = ~P1_REG3_REG_4__SCAN_IN | ~P1_REG3_REG_3__SCAN_IN;
  assign n11219 = ~P1_REG3_REG_5__SCAN_IN;
  assign n11374 = ~n11359 & ~n11219;
  assign n11409 = ~n11374 | ~P1_REG3_REG_6__SCAN_IN;
  assign n11220 = ~P1_REG3_REG_7__SCAN_IN;
  assign n11221 = ~P1_REG3_REG_8__SCAN_IN | ~P1_REG3_REG_9__SCAN_IN;
  assign n11222 = P1_REG3_REG_11__SCAN_IN & P1_REG3_REG_10__SCAN_IN;
  assign n11223 = P1_REG3_REG_13__SCAN_IN & P1_REG3_REG_12__SCAN_IN;
  assign n11608 = ~n11551 | ~n11223;
  assign n11224 = ~P1_REG3_REG_15__SCAN_IN | ~P1_REG3_REG_14__SCAN_IN;
  assign n11225 = ~P1_REG3_REG_17__SCAN_IN | ~P1_REG3_REG_16__SCAN_IN;
  assign n11710 = ~P1_REG3_REG_18__SCAN_IN;
  assign n11772 = ~n11747 | ~P1_REG3_REG_21__SCAN_IN;
  assign n11800 = ~n11772 & ~n14470;
  assign n11788 = ~n11800 | ~P1_REG3_REG_23__SCAN_IN;
  assign n14399 = ~P1_REG3_REG_24__SCAN_IN;
  assign n11828 = ~n11788 & ~n14399;
  assign n11226 = ~P1_REG3_REG_26__SCAN_IN;
  assign n14623 = ~n11855 ^ n11226;
  assign n11239 = ~n14623 | ~n8992;
  assign n11235 = ~n11852 | ~P1_REG0_REG_26__SCAN_IN;
  assign n11234 = ~n11286 | ~P1_REG1_REG_26__SCAN_IN;
  assign n11237 = ~n11235 | ~n11234;
  assign n11236 = n8988 & P1_REG2_REG_26__SCAN_IN;
  assign n11238 = ~n11237 & ~n11236;
  assign n16410 = ~n11239 | ~n11238;
  assign n11240 = ~n14586 & ~n11924;
  assign n11242 = ~n11241 & ~n11240;
  assign n11845 = n11923 ^ n11242;
  assign n11245 = ~n15047 | ~n8995;
  assign n12246 = n13107 & n13191;
  assign n11244 = ~n16410 | ~n11864;
  assign n11846 = ~n11245 | ~n11244;
  assign n14520 = ~n11845 ^ n11846;
  assign n11246 = ~n11285 | ~P1_REG3_REG_1__SCAN_IN;
  assign n11248 = ~n11286 | ~P1_REG1_REG_1__SCAN_IN;
  assign n11250 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n11702 = ~n11263;
  assign n11257 = ~n11251;
  assign n11252 = ~P1_IR_REG_1__SCAN_IN;
  assign n11255 = ~n11252 | ~P1_IR_REG_31__SCAN_IN;
  assign n11253 = ~P1_IR_REG_31__SCAN_IN | ~n15502;
  assign n11254 = ~n11253 | ~P1_IR_REG_1__SCAN_IN;
  assign n11256 = ~n11255 | ~n11254;
  assign n11258 = ~n16251 | ~n11295;
  assign n11260 = ~n11259 | ~n11258;
  assign n11280 = ~n11260 ^ n8991;
  assign n11262 = ~n11285 | ~P1_REG3_REG_0__SCAN_IN;
  assign n11261 = ~n11802 | ~P1_REG0_REG_0__SCAN_IN;
  assign n11267 = ~n11702 | ~n15502;
  assign n11264 = n11263;
  assign n11265 = ~n11973 | ~SI_0_;
  assign n11969 = ~n11265 ^ P2_DATAO_REG_0__SCAN_IN;
  assign n11266 = ~n11263 | ~n11969;
  assign n11268 = ~n15502;
  assign n11269 = n12073 | n11268;
  assign n11275 = ~n11295 | ~n16087;
  assign n11273 = ~P1_REG1_REG_0__SCAN_IN;
  assign n11274 = n12073 | n11273;
  assign n11277 = ~n15411 | ~n15412;
  assign n11279 = ~n11249 | ~n11864;
  assign n11278 = ~n16251 | ~n8995;
  assign n15376 = ~n11279 | ~n11278;
  assign n11284 = ~n15374 | ~n15376;
  assign n11283 = ~n11280;
  assign n11282 = ~n11281;
  assign n11288 = ~n11285 | ~P1_REG3_REG_2__SCAN_IN;
  assign n11287 = ~n11286 | ~P1_REG1_REG_2__SCAN_IN;
  assign n11290 = ~n11288 | ~n11287;
  assign n11297 = ~n16076 | ~n8994;
  assign n11983 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n11292 = n12402 | n11983;
  assign n11291 = ~n11702 | ~n15489;
  assign n11294 = n11292 & n11291;
  assign n11293 = n12401 | n11972;
  assign n15420 = ~n16261;
  assign n11296 = ~n15420 | ~n11295;
  assign n11298 = ~n11297 | ~n11296;
  assign n11302 = ~n11298 ^ n11923;
  assign n11301 = ~n16076 | ~n11864;
  assign n11300 = ~n15420 | ~n8995;
  assign n15424 = n11302 | n11303;
  assign n11306 = ~n15427 | ~n15424;
  assign n11305 = ~n11302;
  assign n15425 = n11305 | n11304;
  assign n11309 = ~n11802 | ~P1_REG0_REG_3__SCAN_IN;
  assign n11308 = ~n11286 | ~P1_REG1_REG_3__SCAN_IN;
  assign n11314 = ~n11309 | ~n11308;
  assign n11312 = ~n8988 | ~P1_REG2_REG_3__SCAN_IN;
  assign n11310 = ~P1_REG3_REG_3__SCAN_IN;
  assign n11311 = ~n8992 | ~n11310;
  assign n11313 = ~n11312 | ~n11311;
  assign n11322 = ~n16046 | ~n8995;
  assign n11315 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n11318 = n12402 | n11315;
  assign n11316 = n11337 | n11228;
  assign n16219 = ~n11316 ^ P1_IR_REG_3__SCAN_IN;
  assign n11317 = ~n11702 | ~n16219;
  assign n11320 = n11318 & n11317;
  assign n11319 = n12401 | n17333;
  assign n11321 = ~n16274 | ~n11295;
  assign n11323 = ~n11322 | ~n11321;
  assign n11327 = ~n11323 ^ n11923;
  assign n11325 = ~n16046 | ~n11864;
  assign n11324 = ~n16274 | ~n8995;
  assign n11326 = ~n11325 | ~n11324;
  assign n15349 = n11327 & n11326;
  assign n15347 = n11327 | n11326;
  assign n11328 = ~P1_REG3_REG_4__SCAN_IN;
  assign n15982 = ~n11328 ^ P1_REG3_REG_3__SCAN_IN;
  assign n11330 = ~n8992 | ~n15982;
  assign n11329 = ~n11286 | ~P1_REG1_REG_4__SCAN_IN;
  assign n11334 = ~n11330 | ~n11329;
  assign n11332 = ~n8988 | ~P1_REG2_REG_4__SCAN_IN;
  assign n11331 = ~n11802 | ~P1_REG0_REG_4__SCAN_IN;
  assign n11333 = ~n11332 | ~n11331;
  assign n11344 = ~n15972 | ~n8995;
  assign n11335 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n11340 = n12402 | n11335;
  assign n11353 = ~n11337 | ~n11336;
  assign n11338 = ~n11353 | ~P1_IR_REG_31__SCAN_IN;
  assign n16213 = ~n11338 ^ P1_IR_REG_4__SCAN_IN;
  assign n11339 = ~n11702 | ~n16213;
  assign n11342 = n11340 & n11339;
  assign n11341 = n17326 | n12401;
  assign n12861 = ~n16283;
  assign n11343 = ~n12861 | ~n11295;
  assign n11345 = ~n11344 | ~n11343;
  assign n11348 = ~n11345 ^ n11811;
  assign n11347 = ~n15972 | ~n11864;
  assign n11346 = ~n12861 | ~n8995;
  assign n11349 = n11347 & n11346;
  assign n15395 = n11348 | n11349;
  assign n11351 = ~n11348;
  assign n11350 = ~n11349;
  assign n11358 = n17319 | n12401;
  assign n11352 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n11356 = n12402 | n11352;
  assign n11354 = ~n11382 | ~P1_IR_REG_31__SCAN_IN;
  assign n16207 = ~n11354 ^ P1_IR_REG_5__SCAN_IN;
  assign n11355 = ~n11702 | ~n16207;
  assign n11357 = n11356 & n11355;
  assign n15959 = ~n11359 ^ P1_REG3_REG_5__SCAN_IN;
  assign n11361 = ~n8992 | ~n15959;
  assign n11360 = ~n11286 | ~P1_REG1_REG_5__SCAN_IN;
  assign n11365 = ~n11361 | ~n11360;
  assign n11363 = ~n8988 | ~P1_REG2_REG_5__SCAN_IN;
  assign n11362 = ~n11802 | ~P1_REG0_REG_5__SCAN_IN;
  assign n11364 = ~n11363 | ~n11362;
  assign n11366 = ~n15930 | ~n8995;
  assign n11368 = ~n11367 | ~n11366;
  assign n12204 = ~n11368 ^ n11811;
  assign n11370 = ~n16296 | ~n8995;
  assign n11369 = ~n15930 | ~n11864;
  assign n12208 = n11370 & n11369;
  assign n11371 = n12204 | n12208;
  assign n11852 = ~n11307;
  assign n11373 = ~n11852 | ~P1_REG0_REG_6__SCAN_IN;
  assign n11372 = ~n11286 | ~P1_REG1_REG_6__SCAN_IN;
  assign n11380 = n11373 & n11372;
  assign n11378 = ~n8988 | ~P1_REG2_REG_6__SCAN_IN;
  assign n11375 = n11374 | P1_REG3_REG_6__SCAN_IN;
  assign n15943 = ~n11409 | ~n11375;
  assign n11376 = ~n15943;
  assign n11377 = ~n11285 | ~n11376;
  assign n11379 = n11378 & n11377;
  assign n11387 = n17312 | n12401;
  assign n11381 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n11385 = n12402 | n11381;
  assign n11425 = ~n11382 & ~P1_IR_REG_5__SCAN_IN;
  assign n11383 = n11425 | n11228;
  assign n15588 = ~n11383 ^ P1_IR_REG_6__SCAN_IN;
  assign n11384 = ~n11702 | ~n15588;
  assign n11386 = n11385 & n11384;
  assign n15946 = ~n11387 | ~n11386;
  assign n11388 = ~n15946 | ~n11295;
  assign n11390 = ~n11389 | ~n11388;
  assign n11397 = ~n11390 ^ n11923;
  assign n11393 = n15326 | n11391;
  assign n11392 = ~n15946 | ~n8995;
  assign n11398 = ~n11393 | ~n11392;
  assign n15450 = n11397 | n11398;
  assign n12202 = ~n12204;
  assign n11394 = ~n12208;
  assign n11395 = n12202 | n11394;
  assign n11396 = n11395 & n15450;
  assign n11400 = ~n11397;
  assign n11399 = ~n11398;
  assign n15451 = n11400 | n11399;
  assign n11402 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n11407 = n12402 | n11402;
  assign n11403 = ~P1_IR_REG_6__SCAN_IN;
  assign n11404 = ~n11425 | ~n11403;
  assign n11405 = ~n11404 | ~P1_IR_REG_31__SCAN_IN;
  assign n16196 = ~n11405 ^ P1_IR_REG_7__SCAN_IN;
  assign n11406 = ~n11702 | ~n16196;
  assign n11408 = n11407 & n11406;
  assign n11417 = ~n16320 | ~n11295;
  assign n11411 = ~n8988 | ~P1_REG2_REG_7__SCAN_IN;
  assign n15914 = ~n11409 ^ P1_REG3_REG_7__SCAN_IN;
  assign n11410 = ~n8992 | ~n15914;
  assign n11415 = n11411 & n11410;
  assign n11413 = ~n11852 | ~P1_REG0_REG_7__SCAN_IN;
  assign n11412 = ~n11286 | ~P1_REG1_REG_7__SCAN_IN;
  assign n11414 = n11413 & n11412;
  assign n11416 = n15437 | n11924;
  assign n11418 = ~n11417 | ~n11416;
  assign n11422 = ~n11418 ^ n11923;
  assign n11420 = ~n16320 | ~n8995;
  assign n11419 = n15437 | n11391;
  assign n11421 = ~n11420 | ~n11419;
  assign n15331 = n11422 | n11421;
  assign n11423 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n11428 = n12402 | n11423;
  assign n11424 = ~P1_IR_REG_7__SCAN_IN & ~P1_IR_REG_6__SCAN_IN;
  assign n11445 = ~n11425 | ~n11424;
  assign n11426 = ~n11445 | ~P1_IR_REG_31__SCAN_IN;
  assign n16190 = ~n11426 ^ P1_IR_REG_8__SCAN_IN;
  assign n11427 = ~n11702 | ~n16190;
  assign n11429 = n11428 & n11427;
  assign n16334 = ~n11430 | ~n11429;
  assign n11439 = ~n16334 | ~n11295;
  assign n11432 = ~n11852 | ~P1_REG0_REG_8__SCAN_IN;
  assign n11431 = ~n11286 | ~P1_REG1_REG_8__SCAN_IN;
  assign n11437 = n11432 & n11431;
  assign n11435 = ~n8988 | ~P1_REG2_REG_8__SCAN_IN;
  assign n11453 = ~P1_REG3_REG_8__SCAN_IN;
  assign n15878 = ~n11454 ^ n11453;
  assign n11433 = ~n15878;
  assign n11434 = ~n8992 | ~n11433;
  assign n11436 = n11435 & n11434;
  assign n11438 = n15848 | n11924;
  assign n11440 = ~n11439 | ~n11438;
  assign n14410 = ~n11440 ^ n11811;
  assign n11442 = ~n16334 | ~n8995;
  assign n11441 = n15848 | n11391;
  assign n11443 = n14410 & n15365;
  assign n11450 = n17291 | n12401;
  assign n11444 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n11448 = n12402 | n11444;
  assign n11446 = ~n11472 | ~P1_IR_REG_31__SCAN_IN;
  assign n15657 = ~n11446 ^ P1_IR_REG_9__SCAN_IN;
  assign n11447 = ~n15657 | ~n11702;
  assign n11449 = n11448 & n11447;
  assign n16353 = ~n11450 | ~n11449;
  assign n11462 = ~n16353 | ~n11295;
  assign n11452 = ~n11852 | ~P1_REG0_REG_9__SCAN_IN;
  assign n11451 = ~n11286 | ~P1_REG1_REG_9__SCAN_IN;
  assign n11460 = n11452 & n11451;
  assign n11458 = ~n8988 | ~P1_REG2_REG_9__SCAN_IN;
  assign n11455 = ~n11454 & ~n11453;
  assign n11456 = ~n11455 & ~P1_REG3_REG_9__SCAN_IN;
  assign n15836 = n11456 | n11504;
  assign n14419 = ~n15836;
  assign n11457 = ~n8992 | ~n14419;
  assign n11459 = n11458 & n11457;
  assign n11463 = ~n11462 | ~n11461;
  assign n11468 = ~n11463 ^ n11811;
  assign n11465 = ~n16353 | ~n8995;
  assign n11464 = n12908 | n11391;
  assign n11469 = ~n11465 | ~n11464;
  assign n14417 = ~n11468 ^ n11469;
  assign n11470 = ~n11468;
  assign n11471 = n11470 | n11469;
  assign n11480 = n17278 | n12401;
  assign n11496 = ~n11472 & ~P1_IR_REG_9__SCAN_IN;
  assign n11473 = ~P1_IR_REG_10__SCAN_IN;
  assign n11474 = ~n11496 | ~n11473;
  assign n11475 = ~n11474 | ~P1_IR_REG_31__SCAN_IN;
  assign n16173 = ~n11475 ^ P1_IR_REG_11__SCAN_IN;
  assign n11478 = ~n16173 | ~n11702;
  assign n11476 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n11477 = n12402 | n11476;
  assign n11479 = n11478 & n11477;
  assign n11492 = ~n15209 | ~n11295;
  assign n11482 = ~n11802 | ~P1_REG0_REG_11__SCAN_IN;
  assign n11481 = ~n11286 | ~P1_REG1_REG_11__SCAN_IN;
  assign n11490 = n11482 & n11481;
  assign n11486 = ~n11551;
  assign n11484 = ~n11504 | ~P1_REG3_REG_10__SCAN_IN;
  assign n11483 = ~P1_REG3_REG_11__SCAN_IN;
  assign n11485 = ~n11484 | ~n11483;
  assign n15005 = n11486 & n11485;
  assign n11488 = ~n8992 | ~n15005;
  assign n11487 = ~n8988 | ~P1_REG2_REG_11__SCAN_IN;
  assign n11489 = n11488 & n11487;
  assign n11491 = n14964 | n11924;
  assign n11493 = ~n11492 | ~n11491;
  assign n11516 = ~n11493 ^ n11923;
  assign n11495 = ~n15209 | ~n8995;
  assign n11494 = n14964 | n11391;
  assign n11517 = ~n11495 | ~n11494;
  assign n14482 = n11516 | n11517;
  assign n11497 = n11496 | n11228;
  assign n15672 = ~n11497 ^ P1_IR_REG_10__SCAN_IN;
  assign n11500 = ~n15672 | ~n11702;
  assign n11498 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n11499 = n12402 | n11498;
  assign n11501 = n11500 & n11499;
  assign n11509 = ~n14296 | ~n11295;
  assign n11502 = ~n11802 | ~P1_REG0_REG_10__SCAN_IN;
  assign n11503 = ~P1_REG3_REG_10__SCAN_IN;
  assign n14292 = ~n11504 ^ n11503;
  assign n11506 = ~n8992 | ~n14292;
  assign n11505 = ~n8988 | ~P1_REG2_REG_10__SCAN_IN;
  assign n11507 = n11506 & n11505;
  assign n11508 = n15847 | n11924;
  assign n11510 = ~n11509 | ~n11508;
  assign n14287 = ~n11510 ^ n11923;
  assign n11512 = ~n14296 | ~n8995;
  assign n11511 = n15847 | n11391;
  assign n14483 = ~n11512 | ~n11511;
  assign n11513 = n14287 | n14483;
  assign n11514 = ~n14482 | ~n11513;
  assign n11515 = n14287 & n14483;
  assign n11520 = ~n14482 | ~n11515;
  assign n11519 = ~n11516;
  assign n11518 = ~n11517;
  assign n14481 = n11519 | n11518;
  assign n11521 = n11520 & n14481;
  assign n11528 = n17271 | n12401;
  assign n11523 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n11526 = n12402 | n11523;
  assign n11524 = n11543 | n11228;
  assign n16167 = ~n11524 ^ P1_IR_REG_12__SCAN_IN;
  assign n11525 = ~n11702 | ~n16167;
  assign n11527 = n11526 & n11525;
  assign n11537 = ~n15198 | ~n11295;
  assign n11530 = ~n11802 | ~P1_REG0_REG_12__SCAN_IN;
  assign n11529 = ~n11286 | ~P1_REG1_REG_12__SCAN_IN;
  assign n11535 = n11530 & n11529;
  assign n11531 = ~P1_REG3_REG_12__SCAN_IN;
  assign n14980 = ~n11551 ^ n11531;
  assign n11533 = ~n8992 | ~n14980;
  assign n11532 = ~n8988 | ~P1_REG2_REG_12__SCAN_IN;
  assign n11534 = n11533 & n11532;
  assign n11536 = n14993 | n11924;
  assign n11538 = ~n11537 | ~n11536;
  assign n11564 = ~n11538 ^ n11923;
  assign n11540 = ~n15198 | ~n8995;
  assign n11539 = n14993 | n11391;
  assign n11565 = ~n11540 | ~n11539;
  assign n14445 = n11564 | n11565;
  assign n11548 = n17265 | n12401;
  assign n11541 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n11546 = n12402 | n11541;
  assign n11542 = ~P1_IR_REG_12__SCAN_IN;
  assign n11576 = ~n11543 | ~n11542;
  assign n11544 = ~n11576 | ~P1_IR_REG_31__SCAN_IN;
  assign n16161 = ~n11544 ^ P1_IR_REG_13__SCAN_IN;
  assign n11545 = ~n11702 | ~n16161;
  assign n11547 = n11546 & n11545;
  assign n11560 = ~n15188 | ~n11295;
  assign n11550 = ~n11802 | ~P1_REG0_REG_13__SCAN_IN;
  assign n11549 = ~n11286 | ~P1_REG1_REG_13__SCAN_IN;
  assign n11558 = n11550 & n11549;
  assign n11553 = ~n11551 | ~P1_REG3_REG_12__SCAN_IN;
  assign n11552 = ~P1_REG3_REG_13__SCAN_IN;
  assign n11554 = ~n11553 | ~n11552;
  assign n14948 = n11554 & n11608;
  assign n11556 = ~n8992 | ~n14948;
  assign n11555 = ~n8988 | ~P1_REG2_REG_13__SCAN_IN;
  assign n11557 = n11556 & n11555;
  assign n11559 = n14965 | n11924;
  assign n11561 = ~n11560 | ~n11559;
  assign n11570 = ~n11561 ^ n11811;
  assign n11563 = ~n15188 | ~n8995;
  assign n11562 = n14965 | n11391;
  assign n11571 = n11563 & n11562;
  assign n14448 = n11570 | n11571;
  assign n11567 = ~n11564;
  assign n11566 = ~n11565;
  assign n12306 = n11567 | n11566;
  assign n11568 = n14448 & n12306;
  assign n11574 = ~n11569 | ~n11568;
  assign n11573 = ~n11570;
  assign n11572 = ~n11571;
  assign n14449 = n11573 | n11572;
  assign n11575 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n11579 = n12402 | n11575;
  assign n11577 = ~n11592 | ~P1_IR_REG_31__SCAN_IN;
  assign n16155 = ~n11577 ^ P1_IR_REG_14__SCAN_IN;
  assign n11578 = ~n11702 | ~n16155;
  assign n11580 = n11579 & n11578;
  assign n11589 = ~n15177 | ~n11295;
  assign n11583 = ~n11852 | ~P1_REG0_REG_14__SCAN_IN;
  assign n11582 = ~n11286 | ~P1_REG1_REG_14__SCAN_IN;
  assign n11587 = n11583 & n11582;
  assign n14924 = ~n11608 ^ P1_REG3_REG_14__SCAN_IN;
  assign n11585 = ~n8992 | ~n14924;
  assign n11584 = ~n8988 | ~P1_REG2_REG_14__SCAN_IN;
  assign n11586 = n11585 & n11584;
  assign n11588 = n14937 | n11924;
  assign n11590 = ~n11589 | ~n11588;
  assign n11604 = n17252 | n12401;
  assign n11591 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n11602 = n12402 | n11591;
  assign n11594 = ~n11592;
  assign n11593 = ~P1_IR_REG_14__SCAN_IN;
  assign n11595 = ~n11594 | ~n11593;
  assign n11596 = ~n11595 | ~P1_IR_REG_31__SCAN_IN;
  assign n11599 = ~n11596 | ~P1_IR_REG_15__SCAN_IN;
  assign n11597 = ~P1_IR_REG_15__SCAN_IN;
  assign n11598 = ~n11597 | ~P1_IR_REG_31__SCAN_IN;
  assign n11600 = ~n11599 | ~n11598;
  assign n16150 = ~n11600 | ~n11636;
  assign n11601 = n11264 | n16150;
  assign n11603 = n11602 & n11601;
  assign n15166 = ~n11604 | ~n11603;
  assign n11617 = ~n15166 | ~n11295;
  assign n11606 = ~n11852 | ~P1_REG0_REG_15__SCAN_IN;
  assign n11605 = ~n11286 | ~P1_REG1_REG_15__SCAN_IN;
  assign n11615 = n11606 & n11605;
  assign n11607 = ~P1_REG3_REG_14__SCAN_IN;
  assign n11610 = n11608 | n11607;
  assign n11609 = ~P1_REG3_REG_15__SCAN_IN;
  assign n11611 = ~n11610 | ~n11609;
  assign n14895 = n11611 & n11666;
  assign n11613 = ~n8992 | ~n14895;
  assign n11612 = ~n8988 | ~P1_REG2_REG_15__SCAN_IN;
  assign n11614 = n11613 & n11612;
  assign n11616 = n14364 | n11924;
  assign n11618 = ~n11617 | ~n11616;
  assign n11629 = ~n11618 ^ n11811;
  assign n11624 = n11628 & n11629;
  assign n11620 = ~n14254;
  assign n11619 = ~n14252;
  assign n11622 = ~n15177 | ~n8995;
  assign n11621 = n14937 | n11391;
  assign n14251 = ~n11622 | ~n11621;
  assign n11623 = ~n11631 | ~n14251;
  assign n11626 = ~n15166 | ~n8995;
  assign n11625 = n14364 | n11391;
  assign n14530 = ~n11626 | ~n11625;
  assign n11627 = ~n14251;
  assign n11633 = ~n11628 | ~n11627;
  assign n11630 = ~n11629;
  assign n11632 = n11631 & n11630;
  assign n11641 = n17245 | n12401;
  assign n11635 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n11639 = n12402 | n11635;
  assign n11637 = ~n11636 | ~P1_IR_REG_31__SCAN_IN;
  assign n16144 = ~n11637 ^ P1_IR_REG_16__SCAN_IN;
  assign n11638 = ~n11702 | ~n16144;
  assign n11640 = n11639 & n11638;
  assign n11649 = ~n15155 | ~n11295;
  assign n11643 = ~n11802 | ~P1_REG0_REG_16__SCAN_IN;
  assign n11642 = ~n11286 | ~P1_REG1_REG_16__SCAN_IN;
  assign n11647 = ~n11643 | ~n11642;
  assign n14872 = ~n11666 ^ P1_REG3_REG_16__SCAN_IN;
  assign n11645 = ~n8992 | ~n14872;
  assign n11644 = ~n8988 | ~P1_REG2_REG_16__SCAN_IN;
  assign n11646 = ~n11645 | ~n11644;
  assign n11648 = ~n14533 | ~n8995;
  assign n11650 = ~n11649 | ~n11648;
  assign n11653 = ~n11650 ^ n11923;
  assign n11652 = ~n15155 | ~n8995;
  assign n11651 = ~n14533 | ~n11864;
  assign n11654 = ~n11652 | ~n11651;
  assign n14358 = n11653 | n11654;
  assign n11656 = ~n11653;
  assign n11655 = ~n11654;
  assign n14359 = n11656 | n11655;
  assign n11662 = n17238 | n12401;
  assign n11657 = ~P2_DATAO_REG_17__SCAN_IN;
  assign n11660 = n12402 | n11657;
  assign n11699 = n11658 | n11228;
  assign n16138 = ~n11699 ^ P1_IR_REG_17__SCAN_IN;
  assign n11659 = ~n16138 | ~n11702;
  assign n11661 = n11660 & n11659;
  assign n11675 = ~n15145 | ~n11295;
  assign n11664 = ~n11802 | ~P1_REG0_REG_17__SCAN_IN;
  assign n11663 = ~n11286 | ~P1_REG1_REG_17__SCAN_IN;
  assign n11673 = n11664 & n11663;
  assign n11665 = ~P1_REG3_REG_16__SCAN_IN;
  assign n11668 = n11666 | n11665;
  assign n11667 = ~P1_REG3_REG_17__SCAN_IN;
  assign n11669 = ~n11668 | ~n11667;
  assign n14844 = n11669 & n11711;
  assign n11671 = ~n8992 | ~n14844;
  assign n11670 = ~n8988 | ~P1_REG2_REG_17__SCAN_IN;
  assign n11672 = n11671 & n11670;
  assign n11674 = n14804 | n11924;
  assign n11676 = ~n11675 | ~n11674;
  assign n11680 = ~n11676 ^ n11923;
  assign n11678 = ~n15145 | ~n8995;
  assign n11677 = n14804 | n11391;
  assign n11679 = ~n11678 | ~n11677;
  assign n14374 = n11680 & n11679;
  assign n11685 = ~n16124 | ~n11825;
  assign n11681 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n11683 = n12402 | n11681;
  assign n11682 = ~n11702 | ~n16090;
  assign n11684 = n11683 & n11682;
  assign n15123 = ~n11685 | ~n11684;
  assign n11694 = ~n15123 | ~n11295;
  assign n11686 = ~P1_REG3_REG_19__SCAN_IN;
  assign n14780 = ~n11713 ^ n11686;
  assign n11688 = ~n14780 | ~n8992;
  assign n11687 = ~n11852 | ~P1_REG0_REG_19__SCAN_IN;
  assign n11692 = ~n11688 | ~n11687;
  assign n11690 = ~n8988 | ~P1_REG2_REG_19__SCAN_IN;
  assign n11689 = ~n11286 | ~P1_REG1_REG_19__SCAN_IN;
  assign n11691 = ~n11690 | ~n11689;
  assign n11693 = ~n14509 | ~n8995;
  assign n11695 = ~n11694 | ~n11693;
  assign n11726 = ~n11695 ^ n11923;
  assign n11697 = ~n15123 | ~n8995;
  assign n11696 = ~n14509 | ~n11864;
  assign n11727 = ~n11697 | ~n11696;
  assign n14318 = n11726 | n11727;
  assign n11707 = ~n16131 | ~n11825;
  assign n11698 = ~P1_IR_REG_17__SCAN_IN;
  assign n11700 = ~n11699 | ~n11698;
  assign n11701 = ~n11700 | ~P1_IR_REG_31__SCAN_IN;
  assign n16132 = ~n11701 ^ P1_IR_REG_18__SCAN_IN;
  assign n11705 = ~n16132 | ~n11702;
  assign n11703 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n11704 = n12402 | n11703;
  assign n11706 = n11705 & n11704;
  assign n11719 = ~n15134 | ~n11295;
  assign n11709 = ~n11852 | ~P1_REG0_REG_18__SCAN_IN;
  assign n11708 = ~n11286 | ~P1_REG1_REG_18__SCAN_IN;
  assign n11717 = n11709 & n11708;
  assign n11712 = n11711 & n11710;
  assign n14817 = ~n11713 & ~n11712;
  assign n11715 = ~n8992 | ~n14817;
  assign n11714 = ~n8988 | ~P1_REG2_REG_18__SCAN_IN;
  assign n11716 = n11715 & n11714;
  assign n11718 = n14828 | n11924;
  assign n11720 = ~n11719 | ~n11718;
  assign n14303 = ~n11720 ^ n11923;
  assign n11722 = ~n15134 | ~n8995;
  assign n11721 = n14828 | n11391;
  assign n14504 = ~n11722 | ~n11721;
  assign n11723 = n14303 | n14504;
  assign n11724 = ~n14318 | ~n11723;
  assign n11725 = n14303 & n14504;
  assign n11730 = ~n14318 | ~n11725;
  assign n11729 = ~n11726;
  assign n11728 = ~n11727;
  assign n11732 = ~n12299 | ~n11825;
  assign n12301 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n11731 = n12402 | n12301;
  assign n15112 = ~n11732 | ~n11731;
  assign n11742 = ~n15112 | ~n11295;
  assign n11734 = ~n11733 & ~P1_REG3_REG_20__SCAN_IN;
  assign n14763 = n11747 | n11734;
  assign n11801 = ~n8992;
  assign n11736 = ~n14763 & ~n11801;
  assign n11735 = n8988 & P1_REG2_REG_20__SCAN_IN;
  assign n11740 = ~n11736 & ~n11735;
  assign n11738 = ~n11852 | ~P1_REG0_REG_20__SCAN_IN;
  assign n11737 = ~n11286 | ~P1_REG1_REG_20__SCAN_IN;
  assign n11739 = n11738 & n11737;
  assign n11741 = n13011 | n11924;
  assign n11743 = ~n11742 | ~n11741;
  assign n11759 = ~n11743 ^ n11923;
  assign n11745 = ~n15112 | ~n8995;
  assign n11744 = n13011 | n11391;
  assign n11760 = ~n11745 | ~n11744;
  assign n12324 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n11746 = n12402 | n12324;
  assign n11755 = ~n15101 | ~n11295;
  assign n14738 = ~n11747 ^ P1_REG3_REG_21__SCAN_IN;
  assign n11753 = n14738 | n11801;
  assign n11749 = ~n11802 | ~P1_REG0_REG_21__SCAN_IN;
  assign n11748 = ~n11286 | ~P1_REG1_REG_21__SCAN_IN;
  assign n11751 = ~n11749 | ~n11748;
  assign n11750 = n8988 & P1_REG2_REG_21__SCAN_IN;
  assign n11752 = ~n11751 & ~n11750;
  assign n11754 = ~n14703 | ~n8995;
  assign n11756 = ~n11755 | ~n11754;
  assign n11764 = ~n11756 ^ n11811;
  assign n11758 = ~n15101 | ~n8995;
  assign n11757 = ~n14703 | ~n11864;
  assign n11765 = n11758 & n11757;
  assign n14326 = n11764 | n11765;
  assign n11762 = ~n11759;
  assign n11761 = ~n11760;
  assign n14322 = n11762 | n11761;
  assign n11763 = n14326 & n14322;
  assign n11767 = ~n11764;
  assign n11766 = ~n11765;
  assign n11771 = ~n11769 | ~n11825;
  assign n12353 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n11770 = n12402 | n12353;
  assign n11780 = ~n15091 | ~n11295;
  assign n14715 = ~n14470 ^ n11772;
  assign n14469 = ~n14715;
  assign n11778 = ~n14469 | ~n8992;
  assign n11774 = ~n11852 | ~P1_REG0_REG_22__SCAN_IN;
  assign n11773 = ~n11286 | ~P1_REG1_REG_22__SCAN_IN;
  assign n11776 = ~n11774 | ~n11773;
  assign n11775 = n8988 & P1_REG2_REG_22__SCAN_IN;
  assign n11777 = ~n11776 & ~n11775;
  assign n16398 = ~n11778 | ~n11777;
  assign n11779 = ~n16398 | ~n8995;
  assign n11781 = ~n11780 | ~n11779;
  assign n11783 = ~n15091 | ~n8995;
  assign n11782 = ~n16398 | ~n11864;
  assign n14463 = ~n11783 | ~n11782;
  assign n15321 = ~P2_DATAO_REG_24__SCAN_IN;
  assign n11784 = n12402 | n15321;
  assign n11794 = ~n15069 | ~n11295;
  assign n11787 = ~n11852 | ~P1_REG0_REG_24__SCAN_IN;
  assign n11786 = ~n11286 | ~P1_REG1_REG_24__SCAN_IN;
  assign n11792 = ~n11787 | ~n11786;
  assign n14669 = ~P1_REG3_REG_24__SCAN_IN ^ n11788;
  assign n11790 = ~n8992 | ~n14669;
  assign n11789 = ~n8988 | ~P1_REG2_REG_24__SCAN_IN;
  assign n11791 = ~n11790 | ~n11789;
  assign n11793 = ~n16404 | ~n8995;
  assign n11795 = ~n11794 | ~n11793;
  assign n11818 = ~n11795 ^ n11811;
  assign n11797 = ~n15069 | ~n8995;
  assign n11796 = ~n16404 | ~n11864;
  assign n11819 = n11797 & n11796;
  assign n14394 = ~n11818 & ~n11819;
  assign n11799 = ~n12334 | ~n11825;
  assign n12330 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n11798 = n12402 | n12330;
  assign n11810 = ~n15080 | ~n11295;
  assign n14692 = ~n11800 ^ P1_REG3_REG_23__SCAN_IN;
  assign n11808 = n14692 | n11801;
  assign n11804 = ~n11852 | ~P1_REG0_REG_23__SCAN_IN;
  assign n11803 = ~n11286 | ~P1_REG1_REG_23__SCAN_IN;
  assign n11806 = ~n11804 | ~n11803;
  assign n11805 = n8988 & P1_REG2_REG_23__SCAN_IN;
  assign n11807 = ~n11806 & ~n11805;
  assign n16401 = ~n11808 | ~n11807;
  assign n11809 = ~n16401 | ~n8995;
  assign n11812 = ~n11810 | ~n11809;
  assign n14265 = ~n11812 ^ n11811;
  assign n11814 = ~n15080 | ~n8995;
  assign n11813 = ~n16401 | ~n11864;
  assign n11815 = ~n14265 & ~n14269;
  assign n11817 = ~n14265 | ~n14269;
  assign n11822 = ~n14394 & ~n11817;
  assign n11821 = ~n11818;
  assign n11820 = ~n11819;
  assign n14393 = ~n11821 & ~n11820;
  assign n11823 = ~n11822 & ~n14393;
  assign n11827 = ~n12345 | ~n11825;
  assign n12348 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n11826 = n12402 | n12348;
  assign n15059 = ~n11827 | ~n11826;
  assign n11837 = ~n15059 | ~n11295;
  assign n14645 = ~P1_REG3_REG_25__SCAN_IN ^ n11828;
  assign n11829 = ~n14645;
  assign n11835 = ~n11829 | ~n8992;
  assign n11831 = ~n11802 | ~P1_REG0_REG_25__SCAN_IN;
  assign n11830 = ~n11286 | ~P1_REG1_REG_25__SCAN_IN;
  assign n11833 = ~n11831 | ~n11830;
  assign n11832 = n8988 & P1_REG2_REG_25__SCAN_IN;
  assign n11834 = ~n11833 & ~n11832;
  assign n16407 = ~n11835 | ~n11834;
  assign n11836 = ~n16407 | ~n8995;
  assign n11838 = ~n11837 | ~n11836;
  assign n11841 = ~n11838 ^ n11923;
  assign n11840 = ~n15059 | ~n8995;
  assign n11839 = ~n16407 | ~n11864;
  assign n11842 = ~n11840 | ~n11839;
  assign n14344 = ~n11841 | ~n11842;
  assign n11844 = ~n11841;
  assign n11843 = ~n11842;
  assign n14343 = ~n11844 | ~n11843;
  assign n11848 = ~n11845;
  assign n11847 = ~n11846;
  assign n11849 = ~n11848 & ~n11847;
  assign n15305 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n11850 = n12402 | n15305;
  assign n11862 = ~n15035 | ~n11295;
  assign n11854 = ~n11852 | ~P1_REG0_REG_27__SCAN_IN;
  assign n11853 = ~n11286 | ~P1_REG1_REG_27__SCAN_IN;
  assign n11860 = ~n11854 | ~n11853;
  assign n11856 = ~n11913;
  assign n14597 = ~P1_REG3_REG_27__SCAN_IN ^ n11856;
  assign n11858 = ~n8992 | ~n14597;
  assign n11857 = ~n8988 | ~P1_REG2_REG_27__SCAN_IN;
  assign n11859 = ~n11858 | ~n11857;
  assign n11861 = ~n16413 | ~n8995;
  assign n11863 = ~n11862 | ~n11861;
  assign n11868 = ~n11863 ^ n11923;
  assign n11866 = ~n15035 | ~n8995;
  assign n11865 = ~n16413 | ~n11864;
  assign n11867 = ~n11866 | ~n11865;
  assign n14235 = ~n11868 | ~n11867;
  assign n11869 = n12346 | n15319;
  assign n11871 = ~n11869 | ~P1_B_REG_SCAN_IN;
  assign n11872 = ~n11871 | ~n11870;
  assign n11873 = ~P1_D_REG_0__SCAN_IN;
  assign n11874 = ~n16122 | ~n11873;
  assign n11880 = ~P1_D_REG_6__SCAN_IN & ~P1_D_REG_7__SCAN_IN;
  assign n11878 = P1_D_REG_8__SCAN_IN | P1_D_REG_9__SCAN_IN;
  assign n11876 = ~P1_D_REG_10__SCAN_IN & ~P1_D_REG_11__SCAN_IN;
  assign n11875 = ~P1_D_REG_12__SCAN_IN & ~P1_D_REG_13__SCAN_IN;
  assign n11877 = ~n11876 | ~n11875;
  assign n11879 = ~n11878 & ~n11877;
  assign n11896 = ~n11880 | ~n11879;
  assign n11882 = ~P1_D_REG_18__SCAN_IN & ~P1_D_REG_19__SCAN_IN;
  assign n11881 = ~P1_D_REG_20__SCAN_IN & ~P1_D_REG_21__SCAN_IN;
  assign n11886 = ~n11882 | ~n11881;
  assign n11884 = ~P1_D_REG_16__SCAN_IN & ~P1_D_REG_14__SCAN_IN;
  assign n11883 = ~P1_D_REG_15__SCAN_IN & ~P1_D_REG_17__SCAN_IN;
  assign n11885 = ~n11884 | ~n11883;
  assign n11894 = ~n11886 & ~n11885;
  assign n11888 = ~P1_D_REG_26__SCAN_IN & ~P1_D_REG_27__SCAN_IN;
  assign n11887 = ~P1_D_REG_28__SCAN_IN & ~P1_D_REG_31__SCAN_IN;
  assign n11892 = ~n11888 | ~n11887;
  assign n11890 = ~P1_D_REG_22__SCAN_IN & ~P1_D_REG_23__SCAN_IN;
  assign n11889 = ~P1_D_REG_24__SCAN_IN & ~P1_D_REG_25__SCAN_IN;
  assign n11891 = ~n11890 | ~n11889;
  assign n11893 = ~n11892 & ~n11891;
  assign n11895 = ~n11894 | ~n11893;
  assign n11901 = ~n11896 & ~n11895;
  assign n11898 = ~P1_D_REG_2__SCAN_IN & ~P1_D_REG_3__SCAN_IN;
  assign n11897 = ~P1_D_REG_4__SCAN_IN & ~P1_D_REG_5__SCAN_IN;
  assign n11899 = ~n11898 | ~n11897;
  assign n11900 = ~P1_D_REG_30__SCAN_IN & ~n11899;
  assign n11902 = ~n11901 | ~n11900;
  assign n11904 = ~P1_D_REG_1__SCAN_IN;
  assign n11906 = ~n16122 | ~n11904;
  assign n11905 = n15310 | n12346;
  assign n12258 = ~n12287 & ~n16239;
  assign n11907 = n12329 & P1_STATE_REG_SCAN_IN;
  assign n11908 = n16241 & n13102;
  assign n13114 = ~n13107;
  assign n11909 = n11908 & n16309;
  assign n11911 = ~n14208 | ~n12394;
  assign n11910 = ~n12395 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n11912 = ~n11911 | ~n11910;
  assign n11952 = ~n11913 | ~P1_REG3_REG_27__SCAN_IN;
  assign n14574 = ~P1_REG3_REG_28__SCAN_IN ^ n11952;
  assign n11915 = ~n8992 | ~n14574;
  assign n11914 = ~n11852 | ~P1_REG0_REG_28__SCAN_IN;
  assign n11919 = ~n11915 | ~n11914;
  assign n11917 = ~n8988 | ~P1_REG2_REG_28__SCAN_IN;
  assign n11916 = ~n11286 | ~P1_REG1_REG_28__SCAN_IN;
  assign n11918 = ~n11917 | ~n11916;
  assign n11920 = ~n14587 & ~n11924;
  assign n11922 = ~n11921 & ~n11920;
  assign n11928 = n11923 ^ n11922;
  assign n11926 = ~n15025 & ~n11924;
  assign n11925 = ~n14587 & ~n11391;
  assign n11927 = ~n11926 & ~n11925;
  assign n11930 = ~n11928 ^ n11927;
  assign n11932 = ~n11930;
  assign n11931 = ~n14235 & ~n15414;
  assign n11964 = ~n11932 | ~n11931;
  assign n16059 = n16245 | n13192;
  assign n16238 = ~n16241;
  assign n11935 = ~n16059 & ~n16238;
  assign n11934 = ~n11935 | ~n11943;
  assign n16337 = n16245 | n13109;
  assign n11933 = ~n16241 | ~n16090;
  assign n11962 = ~n15025 & ~n15442;
  assign n12709 = ~n13191;
  assign n16113 = n13102 | n12709;
  assign n13112 = ~n16113 & ~n16238;
  assign n11936 = ~n11935 & ~n13112;
  assign n15379 = ~n11943 & ~n11936;
  assign n11937 = ~n11943;
  assign n15380 = ~n11937 | ~n16309;
  assign n11938 = ~n15380 | ~n13102;
  assign n11940 = ~n11938 | ~n16113;
  assign n11939 = n12073 & n12329;
  assign n11941 = ~n11940 | ~n11939;
  assign n11942 = n11941 & P1_STATE_REG_SCAN_IN;
  assign n11960 = ~n15402 | ~n14574;
  assign n11948 = n13112 & n11943;
  assign n11945 = n11944;
  assign n12251 = ~n11945;
  assign n11947 = ~n15429 | ~n16413;
  assign n11946 = ~P1_U3084 | ~P1_REG3_REG_28__SCAN_IN;
  assign n11958 = ~n11947 | ~n11946;
  assign n11950 = ~n11802 | ~P1_REG0_REG_29__SCAN_IN;
  assign n11949 = ~n11286 | ~P1_REG1_REG_29__SCAN_IN;
  assign n11956 = ~n11950 | ~n11949;
  assign n11954 = ~n8988 | ~P1_REG2_REG_29__SCAN_IN;
  assign n11951 = ~P1_REG3_REG_28__SCAN_IN;
  assign n12711 = ~n11952 & ~n11951;
  assign n11953 = ~n8992 | ~n12711;
  assign n11955 = ~n11954 | ~n11953;
  assign n11957 = ~n15438 & ~n14562;
  assign n11959 = ~n11958 & ~n11957;
  assign n11961 = ~n11960 | ~n11959;
  assign n11963 = ~n11962 & ~n11961;
  assign n11965 = ~n11964 | ~n11963;
  assign n11968 = ~n11966 | ~P2_U3152;
  assign n11967 = ~P2_STATE_REG_SCAN_IN | ~P2_IR_REG_0__SCAN_IN;
  assign P2_U3358 = ~n11968 | ~n11967;
  assign n11971 = ~n11969 | ~P1_U3084;
  assign n11970 = ~n15502 | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3353 = ~n11971 | ~n11970;
  assign n11981 = ~n11972;
  assign n11980 = ~n11981 | ~n14227;
  assign n11974 = ~n12194;
  assign n11978 = ~n11974 & ~P2_U3152;
  assign n14229 = ~n11975 | ~P2_U3152;
  assign n11977 = ~n14229 & ~n11976;
  assign n11979 = ~n11978 & ~n11977;
  assign P2_U3356 = ~n11980 | ~n11979;
  assign n11987 = ~n11981 | ~n15317;
  assign n11982 = ~n15489;
  assign n11985 = ~n11982 & ~P1_U3084;
  assign n11984 = ~n16128 & ~n11983;
  assign n11986 = ~n11985 & ~n11984;
  assign P1_U3351 = ~n11987 | ~n11986;
  assign n11990 = ~P2_U3966 | ~n11988;
  assign n11989 = ~P2_DATAO_REG_0__SCAN_IN | ~n17594;
  assign P2_U3552 = ~n11990 | ~n11989;
  assign n11992 = ~P2_U3966 | ~n16463;
  assign n11991 = ~P2_DATAO_REG_2__SCAN_IN | ~n17594;
  assign P2_U3554 = ~n11992 | ~n11991;
  assign n11994 = ~P2_U3966 | ~n12430;
  assign n11993 = ~P2_DATAO_REG_1__SCAN_IN | ~n17594;
  assign P2_U3553 = ~n11994 | ~n11993;
  assign n11996 = ~P2_U3966 | ~n16558;
  assign n11995 = ~P2_DATAO_REG_8__SCAN_IN | ~n17594;
  assign P2_U3560 = ~n11996 | ~n11995;
  assign n11998 = ~P2_U3966 | ~n16592;
  assign n11997 = ~P2_DATAO_REG_12__SCAN_IN | ~n17594;
  assign P2_U3564 = ~n11998 | ~n11997;
  assign n12000 = ~P2_U3966 | ~n16505;
  assign n11999 = ~P2_DATAO_REG_11__SCAN_IN | ~n17594;
  assign P2_U3563 = ~n12000 | ~n11999;
  assign n12002 = ~P2_U3966 | ~n16477;
  assign n12001 = ~P2_DATAO_REG_9__SCAN_IN | ~n17594;
  assign P2_U3561 = ~n12002 | ~n12001;
  assign n12004 = ~P2_U3966 | ~n16506;
  assign n12003 = ~P2_DATAO_REG_13__SCAN_IN | ~n17594;
  assign P2_U3565 = ~n12004 | ~n12003;
  assign n12007 = ~P2_U3966 | ~n13935;
  assign n12006 = ~P2_DATAO_REG_14__SCAN_IN | ~n17594;
  assign P2_U3566 = ~n12007 | ~n12006;
  assign n12009 = ~P2_U3966 | ~n13837;
  assign n12008 = ~P2_DATAO_REG_15__SCAN_IN | ~n17594;
  assign P2_U3567 = ~n12009 | ~n12008;
  assign n12011 = ~P2_U3966 | ~n16559;
  assign n12010 = ~P2_DATAO_REG_10__SCAN_IN | ~n17594;
  assign P2_U3562 = ~n12011 | ~n12010;
  assign n12013 = ~P2_U3966 | ~n13871;
  assign n12012 = ~P2_DATAO_REG_16__SCAN_IN | ~n17594;
  assign P2_U3568 = ~n12013 | ~n12012;
  assign n12015 = ~P2_U3966 | ~n13838;
  assign n12014 = ~P2_DATAO_REG_17__SCAN_IN | ~n17594;
  assign P2_U3569 = ~n12015 | ~n12014;
  assign n12017 = ~P2_U3966 | ~n13395;
  assign n12016 = ~P2_DATAO_REG_18__SCAN_IN | ~n17594;
  assign P2_U3570 = ~n12017 | ~n12016;
  assign n12019 = ~P2_U3966 | ~n16541;
  assign n12018 = ~P2_DATAO_REG_3__SCAN_IN | ~n17594;
  assign P2_U3555 = ~n12019 | ~n12018;
  assign n12021 = ~P2_U3966 | ~n16517;
  assign n12020 = ~P2_DATAO_REG_4__SCAN_IN | ~n17594;
  assign P2_U3556 = ~n12021 | ~n12020;
  assign n12023 = ~P2_U3966 | ~n16625;
  assign n12022 = ~P2_DATAO_REG_5__SCAN_IN | ~n17594;
  assign P2_U3557 = ~n12023 | ~n12022;
  assign n12025 = ~P2_U3966 | ~n12459;
  assign n12024 = ~P2_DATAO_REG_6__SCAN_IN | ~n17594;
  assign P2_U3558 = ~n12025 | ~n12024;
  assign n12028 = ~P2_U3966 | ~n16627;
  assign n12027 = ~P2_DATAO_REG_7__SCAN_IN | ~n17594;
  assign P2_U3559 = ~n12028 | ~n12027;
  assign n12030 = ~P1_U4006 | ~n16046;
  assign n12029 = ~n16425 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P1_U3558 = ~n12030 | ~n12029;
  assign n12032 = ~P1_U4006 | ~n15930;
  assign n12031 = ~n16425 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P1_U3560 = ~n12032 | ~n12031;
  assign n12034 = ~P1_U4006 | ~n15972;
  assign n12033 = ~n16425 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P1_U3559 = ~n12034 | ~n12033;
  assign n12036 = ~P1_U4006 | ~n14533;
  assign n12035 = ~n16425 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P1_U3571 = ~n12036 | ~n12035;
  assign n12038 = ~P1_U4006 | ~n16078;
  assign n12037 = ~n16425 | ~P1_DATAO_REG_0__SCAN_IN;
  assign P1_U3555 = ~n12038 | ~n12037;
  assign n12040 = ~P1_U4006 | ~n11249;
  assign n12039 = ~n16425 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U3556 = ~n12040 | ~n12039;
  assign n12042 = ~P1_U4006 | ~n16076;
  assign n12041 = ~n16425 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P1_U3557 = ~n12042 | ~n12041;
  assign n14453 = ~n14993;
  assign n12044 = ~n14453 | ~P1_U4006;
  assign n12043 = ~n16425 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P1_U3567 = ~n12044 | ~n12043;
  assign n12046 = ~n15881 | ~P1_U4006;
  assign n12045 = ~n16425 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P1_U3564 = ~n12046 | ~n12045;
  assign n12048 = ~n14509 | ~P1_U4006;
  assign n12047 = ~n16425 | ~P1_DATAO_REG_19__SCAN_IN;
  assign P1_U3574 = ~n12048 | ~n12047;
  assign n12050 = ~n15929 | ~P1_U4006;
  assign n12049 = ~n16425 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P1_U3562 = ~n12050 | ~n12049;
  assign n12052 = ~n15958 | ~P1_U4006;
  assign n12051 = ~n16425 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P1_U3561 = ~n12052 | ~n12051;
  assign n14535 = ~n14937;
  assign n12054 = ~n14535 | ~P1_U4006;
  assign n12053 = ~n16425 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P1_U3569 = ~n12054 | ~n12053;
  assign n12056 = ~n14907 | ~P1_U4006;
  assign n12055 = ~n16425 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U3568 = ~n12056 | ~n12055;
  assign n14490 = ~n15847;
  assign n12058 = ~n14490 | ~P1_U4006;
  assign n12057 = ~n16425 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U3565 = ~n12058 | ~n12057;
  assign n12060 = ~n14859 | ~P1_U4006;
  assign n12059 = ~n16425 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P1_U3572 = ~n12060 | ~n12059;
  assign n12062 = ~n14703 | ~P1_U4006;
  assign n12061 = ~n16425 | ~P1_DATAO_REG_21__SCAN_IN;
  assign P1_U3576 = ~n12062 | ~n12061;
  assign n12064 = ~n15903 | ~P1_U4006;
  assign n12063 = ~n16425 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P1_U3563 = ~n12064 | ~n12063;
  assign n12066 = ~n14774 | ~P1_U4006;
  assign n12065 = ~n16425 | ~P1_DATAO_REG_20__SCAN_IN;
  assign P1_U3575 = ~n12066 | ~n12065;
  assign n12654 = ~n14964;
  assign n12068 = ~n12654 | ~P1_U4006;
  assign n12067 = ~n16425 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U3566 = ~n12068 | ~n12067;
  assign n12070 = ~n14908 | ~P1_U4006;
  assign n12069 = ~n16425 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P1_U3570 = ~n12070 | ~n12069;
  assign n14775 = ~n14828;
  assign n12072 = ~n14775 | ~P1_U4006;
  assign n12071 = ~n16425 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P1_U3573 = ~n12072 | ~n12071;
  assign n12074 = ~n13102 | ~n12073;
  assign n12075 = ~n12074 | ~n12329;
  assign n12086 = ~n12075 | ~n11264;
  assign P1_U3083 = ~n12086 | ~P1_STATE_REG_SCAN_IN;
  assign n15341 = ~P1_REG3_REG_3__SCAN_IN | ~P1_U3084;
  assign n12097 = ~n12075 | ~n9160;
  assign n15830 = ~n12097 & ~n11945;
  assign n12076 = ~P1_REG2_REG_2__SCAN_IN;
  assign n15484 = ~n15489 ^ n12076;
  assign n15480 = ~n16226 ^ P1_REG2_REG_1__SCAN_IN;
  assign n15479 = n15502 & P1_REG2_REG_0__SCAN_IN;
  assign n12077 = ~n15479;
  assign n12079 = n15480 | n12077;
  assign n12078 = ~n16226 | ~P1_REG2_REG_1__SCAN_IN;
  assign n15485 = ~n12079 | ~n12078;
  assign n12081 = ~n15484 | ~n15485;
  assign n12080 = ~n15489 | ~P1_REG2_REG_2__SCAN_IN;
  assign n15515 = ~n12081 | ~n12080;
  assign n12082 = ~P1_REG2_REG_3__SCAN_IN;
  assign n15514 = ~n16219 ^ n12082;
  assign n12083 = n15515 ^ n15514;
  assign n12084 = ~n15830 | ~n12083;
  assign n12096 = ~n15341 | ~n12084;
  assign n15818 = ~P1_U3083 & ~n12085;
  assign n12094 = ~P1_ADDR_REG_3__SCAN_IN | ~n15818;
  assign n15465 = n12086 | P1_U3084;
  assign n15496 = ~n15494;
  assign n12087 = ~P1_REG1_REG_2__SCAN_IN;
  assign n15508 = ~n15489 ^ n12087;
  assign n15472 = ~n16226 ^ P1_REG1_REG_1__SCAN_IN;
  assign n15473 = ~n15502 | ~P1_REG1_REG_0__SCAN_IN;
  assign n12089 = n15472 | n15473;
  assign n12088 = ~n16226 | ~P1_REG1_REG_1__SCAN_IN;
  assign n15507 = ~n12089 | ~n12088;
  assign n15506 = ~n15508 | ~n15507;
  assign n12090 = ~n15489 | ~P1_REG1_REG_2__SCAN_IN;
  assign n12091 = ~P1_REG1_REG_3__SCAN_IN;
  assign n15530 = ~n16219 ^ n12091;
  assign n12092 = n15531 ^ n15530;
  assign n12093 = ~n15816 | ~n12092;
  assign n12095 = ~n12094 | ~n12093;
  assign n12100 = ~n12096 & ~n12095;
  assign n12099 = ~n12098 | ~n16219;
  assign P1_U3244 = ~n12100 | ~n12099;
  assign n16556 = ~P2_REG3_REG_9__SCAN_IN | ~P2_U3152;
  assign n12103 = ~n12101 | ~n12335;
  assign n12105 = ~n12103 | ~n12102;
  assign n12104 = ~n17225 | ~n12584;
  assign n12106 = ~n16913 | ~P2_ADDR_REG_9__SCAN_IN;
  assign n12151 = ~n16556 | ~n12106;
  assign n12109 = ~n17225 | ~n13260;
  assign n14210 = n11147 | P2_U3152;
  assign n12107 = n12586 | n14210;
  assign n12108 = n12107 & n12335;
  assign n12111 = ~n12109 | ~n12108;
  assign n12143 = ~n12111 | ~n12110;
  assign n12145 = ~n14214;
  assign n16921 = ~n12143 & ~n12145;
  assign n12170 = P2_REG1_REG_1__SCAN_IN ^ n17342;
  assign n16650 = ~P2_IR_REG_0__SCAN_IN;
  assign n16638 = ~P2_REG1_REG_0__SCAN_IN;
  assign n12171 = ~n16650 & ~n16638;
  assign n12113 = ~n12170 | ~n12171;
  assign n12112 = ~n17342 | ~P2_REG1_REG_1__SCAN_IN;
  assign n12184 = ~n12113 | ~n12112;
  assign n12114 = ~n12194 | ~P2_REG1_REG_2__SCAN_IN;
  assign n12115 = ~P2_REG1_REG_3__SCAN_IN;
  assign n16656 = ~n17334 ^ n12115;
  assign n12116 = ~n17334 | ~P2_REG1_REG_3__SCAN_IN;
  assign n16671 = ~n12117 | ~n12116;
  assign n12118 = ~P2_REG1_REG_4__SCAN_IN;
  assign n16672 = ~n17327 ^ n12118;
  assign n12120 = ~n16671 | ~n16672;
  assign n12119 = ~n17327 | ~P2_REG1_REG_4__SCAN_IN;
  assign n12156 = ~n12120 | ~n12119;
  assign n12121 = ~P2_REG1_REG_5__SCAN_IN;
  assign n12157 = ~n17320 ^ n12121;
  assign n12123 = ~n12156 | ~n12157;
  assign n12122 = ~n17320 | ~P2_REG1_REG_5__SCAN_IN;
  assign n16694 = P2_REG1_REG_6__SCAN_IN ^ n17313;
  assign n12124 = ~n17313 | ~P2_REG1_REG_6__SCAN_IN;
  assign n12125 = ~P2_REG1_REG_7__SCAN_IN;
  assign n16704 = ~n17306 ^ n12125;
  assign n12126 = ~n17306 | ~P2_REG1_REG_7__SCAN_IN;
  assign n16720 = ~n12127 | ~n12126;
  assign n16719 = ~n17299 ^ P2_REG1_REG_8__SCAN_IN;
  assign n12128 = ~n16719;
  assign n12129 = ~n17299 | ~P2_REG1_REG_8__SCAN_IN;
  assign n16743 = ~n17292 ^ P2_REG1_REG_9__SCAN_IN;
  assign n12130 = ~n16744 ^ n16743;
  assign n12149 = ~n16921 | ~n12130;
  assign n12173 = P2_REG2_REG_1__SCAN_IN ^ n17342;
  assign n17219 = ~P2_REG2_REG_0__SCAN_IN;
  assign n12174 = ~n16650 & ~n17219;
  assign n12132 = ~n12173 | ~n12174;
  assign n12131 = ~n17342 | ~P2_REG2_REG_1__SCAN_IN;
  assign n12187 = ~n12132 | ~n12131;
  assign n12188 = P2_REG2_REG_2__SCAN_IN ^ n12194;
  assign n12134 = ~n12187 | ~n12188;
  assign n12133 = ~n12194 | ~P2_REG2_REG_2__SCAN_IN;
  assign n16661 = ~n12134 | ~n12133;
  assign n16660 = P2_REG2_REG_3__SCAN_IN ^ n17334;
  assign n16662 = ~n16661 | ~n16660;
  assign n12135 = ~n17334 | ~P2_REG2_REG_3__SCAN_IN;
  assign n16677 = ~n16662 | ~n12135;
  assign n16676 = P2_REG2_REG_4__SCAN_IN ^ n17327;
  assign n16678 = ~n16677 | ~n16676;
  assign n12136 = ~n17327 | ~P2_REG2_REG_4__SCAN_IN;
  assign n12159 = ~n16678 | ~n12136;
  assign n12137 = ~P2_REG2_REG_5__SCAN_IN;
  assign n12160 = ~n17320 ^ n12137;
  assign n12139 = ~n12159 | ~n12160;
  assign n12138 = ~n17320 | ~P2_REG2_REG_5__SCAN_IN;
  assign n16688 = ~n12139 | ~n12138;
  assign n16687 = n17313 & P2_REG2_REG_6__SCAN_IN;
  assign n12140 = ~n16688 & ~n16687;
  assign n16709 = ~n12140 & ~n9025;
  assign n16708 = P2_REG2_REG_7__SCAN_IN ^ n17306;
  assign n16710 = ~n16709 | ~n16708;
  assign n12141 = ~n17306 | ~P2_REG2_REG_7__SCAN_IN;
  assign n16725 = ~n16710 | ~n12141;
  assign n16724 = P2_REG2_REG_8__SCAN_IN ^ n17299;
  assign n16726 = ~n16725 | ~n16724;
  assign n12142 = ~n17299 | ~P2_REG2_REG_8__SCAN_IN;
  assign n16737 = ~n16726 | ~n12142;
  assign n16735 = ~n17292 ^ P2_REG2_REG_9__SCAN_IN;
  assign n12147 = ~n16737 ^ n16735;
  assign n12144 = ~n12143;
  assign n12146 = ~n12598 | ~n12145;
  assign n16911 = ~n12152 & ~n12146;
  assign n12148 = ~n12147 | ~n16911;
  assign n12150 = ~n12149 | ~n12148;
  assign n12154 = ~n12151 & ~n12150;
  assign n12153 = ~n16872 | ~n17292;
  assign P2_U3254 = ~n12154 | ~n12153;
  assign n16520 = ~P2_REG3_REG_5__SCAN_IN | ~P2_U3152;
  assign n12155 = ~n16913 | ~P2_ADDR_REG_5__SCAN_IN;
  assign n12165 = ~n16520 | ~n12155;
  assign n12158 = n12157 ^ n12156;
  assign n12163 = ~n16921 | ~n12158;
  assign n12161 = n12160 ^ n12159;
  assign n12162 = ~n12161 | ~n16911;
  assign n12164 = ~n12163 | ~n12162;
  assign n12167 = ~n12165 & ~n12164;
  assign n12166 = ~n16872 | ~n17320;
  assign P2_U3250 = ~n12167 | ~n12166;
  assign n12169 = ~P2_ADDR_REG_1__SCAN_IN | ~n16913;
  assign n12168 = ~P2_REG3_REG_1__SCAN_IN | ~P2_U3152;
  assign n12179 = ~n12169 | ~n12168;
  assign n12172 = n12171 ^ n12170;
  assign n12177 = ~n16921 | ~n12172;
  assign n12175 = n12174 ^ n12173;
  assign n12176 = ~n12175 | ~n16911;
  assign n12178 = ~n12177 | ~n12176;
  assign n12181 = ~n12179 & ~n12178;
  assign n12180 = ~n16922 | ~n17342;
  assign P2_U3246 = ~n12181 | ~n12180;
  assign n12183 = ~P2_ADDR_REG_2__SCAN_IN | ~n16913;
  assign n12182 = ~P2_REG3_REG_2__SCAN_IN | ~P2_U3152;
  assign n12193 = ~n12183 | ~n12182;
  assign n12186 = n12185 ^ n12184;
  assign n12191 = ~n16921 | ~n12186;
  assign n12189 = n12188 ^ n12187;
  assign n12190 = ~n12189 | ~n16911;
  assign n12192 = ~n12191 | ~n12190;
  assign n12196 = ~n12193 & ~n12192;
  assign n12195 = ~n16922 | ~n12194;
  assign P2_U3247 = ~n12196 | ~n12195;
  assign n12201 = ~n12299 | ~n14227;
  assign n12199 = ~n13537 & ~P2_U3152;
  assign n12198 = ~n14229 & ~n12197;
  assign n12200 = ~n12199 & ~n12198;
  assign P2_U3338 = ~n12201 | ~n12200;
  assign n12220 = ~n15402 | ~n15959;
  assign n12218 = ~n15419 | ~n15958;
  assign n15539 = ~P1_REG3_REG_5__SCAN_IN | ~P1_U3084;
  assign n12216 = ~n15539;
  assign n12203 = ~n12205;
  assign n15452 = ~n12203 & ~n12202;
  assign n12206 = ~n12205 & ~n12204;
  assign n12207 = ~n15452 & ~n12206;
  assign n15454 = ~n12207 | ~n12208;
  assign n12209 = n12208 | n12207;
  assign n12210 = ~n15454 | ~n12209;
  assign n12214 = ~n15457 | ~n12210;
  assign n12212 = ~n15961 & ~n15442;
  assign n16026 = ~n15972;
  assign n12211 = ~n16026 & ~n15441;
  assign n12213 = ~n12212 & ~n12211;
  assign n12215 = ~n12214 | ~n12213;
  assign n12217 = ~n12216 & ~n12215;
  assign n12219 = n12218 & n12217;
  assign P1_U3225 = ~n12220 | ~n12219;
  assign n13133 = ~n16070 | ~n12829;
  assign n13140 = ~n16076 | ~n16261;
  assign n12228 = n13142 & n13140;
  assign n16053 = ~n13133 | ~n12228;
  assign n13149 = ~n15326 | ~n15946;
  assign n13148 = n15961 | n15930;
  assign n15920 = n15930 & n15961;
  assign n13154 = ~n13149 | ~n15920;
  assign n12868 = ~n16310 | ~n15958;
  assign n12221 = ~n13154 | ~n12868;
  assign n15861 = ~n16320 | ~n15437;
  assign n12896 = ~n16334 | ~n15848;
  assign n12733 = n12896 & n15861;
  assign n12731 = ~n16353 | ~n12908;
  assign n12804 = n16353 | n12908;
  assign n12805 = ~n12759;
  assign n12732 = n14296 & n15847;
  assign n12223 = ~n12732;
  assign n12226 = ~n12644 ^ n12652;
  assign n12225 = n13107 | n16125;
  assign n12224 = n9500 | n13192;
  assign n12257 = ~n12226 & ~n16074;
  assign n16083 = ~n16078 | ~n16087;
  assign n12227 = ~n11249 | ~n16251;
  assign n16051 = ~n12228;
  assign n12834 = n16076 | n15420;
  assign n15986 = ~n16041 | ~n12834;
  assign n12229 = ~n15918;
  assign n12742 = ~n12737;
  assign n15989 = ~n12229 | ~n12742;
  assign n12231 = ~n13143;
  assign n12230 = ~n12736;
  assign n12232 = n15989 & n16020;
  assign n15987 = ~n16046 & ~n16274;
  assign n12233 = ~n15989 | ~n15987;
  assign n12852 = n15972 | n12861;
  assign n12234 = n12233 & n12852;
  assign n12235 = ~n15920;
  assign n12859 = ~n15930 | ~n16296;
  assign n15890 = ~n15946 & ~n15958;
  assign n12888 = n16320 | n15929;
  assign n15865 = n12237 & n12888;
  assign n15864 = ~n15891 | ~n15925;
  assign n12240 = ~n12238 | ~n15865;
  assign n12239 = ~n16334 | ~n15903;
  assign n12243 = n16353 | n15881;
  assign n12244 = ~n16353 | ~n15881;
  assign n12267 = ~n12245 ^ n12652;
  assign n12250 = ~n12246 | ~n9504;
  assign n12249 = n12248 | n12247;
  assign n12255 = ~n12267 | ~n16084;
  assign n12253 = ~n14964 & ~n16025;
  assign n12252 = ~n12908 & ~n16023;
  assign n12254 = ~n12253 & ~n12252;
  assign n12256 = ~n12255 | ~n12254;
  assign n12285 = ~n12257 & ~n12256;
  assign n12259 = ~n12258;
  assign n12262 = ~n12294 & ~n12259;
  assign n12260 = n13102 | n13191;
  assign n12261 = ~n15378;
  assign n12263 = ~n12262 | ~n12261;
  assign n12266 = ~n12285 | ~n16119;
  assign n12264 = ~P1_REG2_REG_10__SCAN_IN;
  assign n12265 = ~n16104 | ~n12264;
  assign n12278 = ~n12266 | ~n12265;
  assign n12279 = ~n12267;
  assign n16095 = n12268 | n16125;
  assign n12276 = ~n12279 & ~n16003;
  assign n16037 = ~n16251 & ~n9487;
  assign n16039 = ~n16037 | ~n16261;
  assign n15938 = ~n15956 | ~n16310;
  assign n15874 = ~n15875 & ~n16334;
  assign n12269 = ~n16353;
  assign n12270 = ~n12406 ^ n14296;
  assign n16350 = ~n16337;
  assign n12281 = ~n12270 | ~n16350;
  assign n14979 = n16104 | n16090;
  assign n12274 = ~n12281 & ~n14979;
  assign n12272 = ~n16108 | ~n14296;
  assign n12271 = ~n16105 | ~n14292;
  assign n12273 = ~n12272 | ~n12271;
  assign n12275 = n12274 | n12273;
  assign n12277 = ~n12276 & ~n12275;
  assign P1_U3281 = ~n12278 | ~n12277;
  assign n12283 = ~n12279 & ~n16357;
  assign n16352 = ~n16309;
  assign n12280 = ~n14296 | ~n16352;
  assign n12282 = ~n12281 | ~n12280;
  assign n12284 = ~n12283 & ~n12282;
  assign n12296 = ~n12285 | ~n12284;
  assign n12286 = ~n16337 & ~n16125;
  assign n12293 = ~n12296 | ~n16363;
  assign n12292 = ~n16349 | ~P1_REG0_REG_10__SCAN_IN;
  assign P1_U3484 = ~n12293 | ~n12292;
  assign n12298 = ~n12296 | ~n16395;
  assign n12297 = ~n16393 | ~P1_REG1_REG_10__SCAN_IN;
  assign P1_U3533 = ~n12298 | ~n12297;
  assign n12300 = ~n12299;
  assign n12305 = ~n12300 & ~n16225;
  assign n12303 = n13192 | P1_U3084;
  assign n12302 = n16128 | n12301;
  assign n12304 = ~n12303 | ~n12302;
  assign P1_U3333 = n12305 | n12304;
  assign n14444 = ~n14445 | ~n12306;
  assign n12317 = ~n12307 | ~n15457;
  assign n12308 = ~n15198;
  assign n12315 = ~n12308 & ~n15442;
  assign n12313 = ~n15402 | ~n14980;
  assign n12311 = ~n15441 & ~n14964;
  assign n12309 = ~n15419 | ~n14907;
  assign n15689 = ~P1_REG3_REG_12__SCAN_IN | ~P1_U3084;
  assign n12310 = ~n12309 | ~n15689;
  assign n12312 = ~n12311 & ~n12310;
  assign n12314 = ~n12313 | ~n12312;
  assign n12316 = ~n12315 & ~n12314;
  assign P1_U3222 = ~n12317 | ~n12316;
  assign n12321 = ~n12322 & ~n17340;
  assign n12319 = n12424 | P2_U3152;
  assign n12318 = ~n17347 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n12320 = ~n12319 | ~n12318;
  assign P2_U3337 = n12321 | n12320;
  assign n12323 = ~n12322;
  assign n12328 = ~n12323 | ~n15317;
  assign n12326 = ~n9500 & ~P1_U3084;
  assign n12325 = ~n16128 & ~n12324;
  assign n12327 = ~n12326 & ~n12325;
  assign P1_U3332 = ~n12328 | ~n12327;
  assign n12333 = ~n12334 | ~n15317;
  assign n13113 = n12329 | P1_U3084;
  assign n13197 = ~n13113;
  assign n12331 = ~n16128 & ~n12330;
  assign n12332 = ~n13197 & ~n12331;
  assign P1_U3330 = ~n12333 | ~n12332;
  assign n12339 = ~n12334 | ~n14227;
  assign n12337 = ~n14229 & ~n12336;
  assign n12338 = ~n11126 & ~n12337;
  assign P2_U3335 = ~n12339 | ~n12338;
  assign n12344 = ~n12345 | ~n14227;
  assign n12342 = ~n14229 & ~n12340;
  assign n12341 = ~P2_U3152 & ~n12569;
  assign n12343 = ~n12342 & ~n12341;
  assign P2_U3333 = ~n12344 | ~n12343;
  assign n12352 = ~n12345 | ~n15317;
  assign n12347 = ~n12346;
  assign n12350 = ~n12347 & ~P1_U3084;
  assign n12349 = ~n16128 & ~n12348;
  assign n12351 = ~n12350 & ~n12349;
  assign P1_U3328 = ~n12352 | ~n12351;
  assign n12357 = ~n11769 | ~n15317;
  assign n12355 = ~n13107 & ~P1_U3084;
  assign n12354 = ~n16128 & ~n12353;
  assign n12356 = ~n12355 & ~n12354;
  assign P1_U3331 = ~n12357 | ~n12356;
  assign n12362 = ~n11769 | ~n14227;
  assign n12360 = ~n10825 & ~P2_U3152;
  assign n12359 = ~n14229 & ~n12358;
  assign n12361 = ~n12360 & ~n12359;
  assign P2_U3336 = ~n12362 | ~n12361;
  assign n12391 = ~P1_ADDR_REG_18__SCAN_IN & ~P2_ADDR_REG_18__SCAN_IN;
  assign n17620 = ~P1_ADDR_REG_17__SCAN_IN & ~P2_ADDR_REG_17__SCAN_IN;
  assign n17619 = P1_ADDR_REG_17__SCAN_IN & P2_ADDR_REG_17__SCAN_IN;
  assign n17624 = ~P1_ADDR_REG_16__SCAN_IN & ~P2_ADDR_REG_16__SCAN_IN;
  assign n17623 = P1_ADDR_REG_16__SCAN_IN & P2_ADDR_REG_16__SCAN_IN;
  assign n17628 = ~P1_ADDR_REG_15__SCAN_IN & ~P2_ADDR_REG_15__SCAN_IN;
  assign n17627 = P1_ADDR_REG_15__SCAN_IN & P2_ADDR_REG_15__SCAN_IN;
  assign n17632 = ~P1_ADDR_REG_14__SCAN_IN & ~P2_ADDR_REG_14__SCAN_IN;
  assign n17631 = P1_ADDR_REG_14__SCAN_IN & P2_ADDR_REG_14__SCAN_IN;
  assign n17636 = ~P2_ADDR_REG_13__SCAN_IN & ~P1_ADDR_REG_13__SCAN_IN;
  assign n17635 = P2_ADDR_REG_13__SCAN_IN & P1_ADDR_REG_13__SCAN_IN;
  assign n17640 = ~P1_ADDR_REG_12__SCAN_IN & ~P2_ADDR_REG_12__SCAN_IN;
  assign n17639 = P1_ADDR_REG_12__SCAN_IN & P2_ADDR_REG_12__SCAN_IN;
  assign n17644 = ~P1_ADDR_REG_11__SCAN_IN & ~P2_ADDR_REG_11__SCAN_IN;
  assign n17648 = ~P1_ADDR_REG_10__SCAN_IN & ~P2_ADDR_REG_10__SCAN_IN;
  assign n12381 = ~P2_ADDR_REG_9__SCAN_IN & ~P1_ADDR_REG_9__SCAN_IN;
  assign n12379 = ~P2_ADDR_REG_8__SCAN_IN & ~P1_ADDR_REG_8__SCAN_IN;
  assign n12377 = ~P1_ADDR_REG_7__SCAN_IN & ~P2_ADDR_REG_7__SCAN_IN;
  assign n12375 = ~P2_ADDR_REG_6__SCAN_IN & ~P1_ADDR_REG_6__SCAN_IN;
  assign n12373 = ~P2_ADDR_REG_5__SCAN_IN & ~P1_ADDR_REG_5__SCAN_IN;
  assign n12371 = ~P2_ADDR_REG_4__SCAN_IN & ~P1_ADDR_REG_4__SCAN_IN;
  assign n12369 = ~P1_ADDR_REG_3__SCAN_IN | ~P2_ADDR_REG_3__SCAN_IN;
  assign n17614 = P1_ADDR_REG_3__SCAN_IN ^ P2_ADDR_REG_3__SCAN_IN;
  assign n12367 = ~P1_ADDR_REG_2__SCAN_IN | ~P2_ADDR_REG_2__SCAN_IN;
  assign n12364 = ~P1_ADDR_REG_1__SCAN_IN;
  assign n12363 = ~P1_ADDR_REG_0__SCAN_IN | ~P2_ADDR_REG_0__SCAN_IN;
  assign n17599 = n12364 & n12363;
  assign n17598 = ~n12364 & ~n12363;
  assign n12365 = ~P2_ADDR_REG_1__SCAN_IN & ~n17598;
  assign n17616 = ~n17599 & ~n12365;
  assign n17615 = P1_ADDR_REG_2__SCAN_IN ^ P2_ADDR_REG_2__SCAN_IN;
  assign n12366 = ~n17616 | ~n17615;
  assign n17613 = ~n12367 | ~n12366;
  assign n12368 = ~n17614 | ~n17613;
  assign n17612 = ~n12369 | ~n12368;
  assign n17611 = ~P2_ADDR_REG_4__SCAN_IN ^ P1_ADDR_REG_4__SCAN_IN;
  assign n12370 = ~n17612 & ~n17611;
  assign n17610 = ~n12371 & ~n12370;
  assign n17609 = ~P2_ADDR_REG_5__SCAN_IN ^ P1_ADDR_REG_5__SCAN_IN;
  assign n12372 = ~n17610 & ~n17609;
  assign n17608 = ~n12373 & ~n12372;
  assign n17607 = ~P2_ADDR_REG_6__SCAN_IN ^ P1_ADDR_REG_6__SCAN_IN;
  assign n12374 = ~n17608 & ~n17607;
  assign n17606 = ~n12375 & ~n12374;
  assign n17605 = ~P1_ADDR_REG_7__SCAN_IN ^ P2_ADDR_REG_7__SCAN_IN;
  assign n12376 = ~n17606 & ~n17605;
  assign n17604 = ~n12377 & ~n12376;
  assign n17603 = ~P2_ADDR_REG_8__SCAN_IN ^ P1_ADDR_REG_8__SCAN_IN;
  assign n12378 = ~n17604 & ~n17603;
  assign n17602 = ~n12379 & ~n12378;
  assign n17601 = ~P2_ADDR_REG_9__SCAN_IN ^ P1_ADDR_REG_9__SCAN_IN;
  assign n12380 = ~n17602 & ~n17601;
  assign n12382 = ~n17647 & ~n17650;
  assign n12383 = ~n17643 & ~n17646;
  assign n12384 = ~n17639 & ~n17642;
  assign n12385 = ~n17635 & ~n17638;
  assign n12386 = ~n17631 & ~n17634;
  assign n12387 = ~n17627 & ~n17630;
  assign n12388 = ~n17623 & ~n17626;
  assign n17622 = ~n17624 & ~n12388;
  assign n12389 = ~n17619 & ~n17622;
  assign n17618 = ~n17620 & ~n12389;
  assign n17617 = ~P1_ADDR_REG_18__SCAN_IN ^ P2_ADDR_REG_18__SCAN_IN;
  assign n12390 = ~n17618 & ~n17617;
  assign n12393 = ~n12391 & ~n12390;
  assign n12392 = ~P2_ADDR_REG_19__SCAN_IN ^ P1_ADDR_REG_19__SCAN_IN;
  assign ADD_1071_U4 = ~n12393 ^ n12392;
  assign n12397 = ~n15275 | ~n12394;
  assign n12396 = ~n12395 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n12398 = ~n12397 | ~n12396;
  assign n14545 = ~n12398 | ~n11264;
  assign n13090 = ~n14545;
  assign n15287 = ~P2_DATAO_REG_30__SCAN_IN;
  assign n12399 = n12402 | n15287;
  assign n12404 = n14202 | n12401;
  assign n15293 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n12403 = n12402 | n15293;
  assign n12405 = ~n14296;
  assign n15003 = ~n12406 | ~n12405;
  assign n14919 = ~n15177;
  assign n14815 = ~n14871 | ~n14843;
  assign n14762 = ~n15112;
  assign n14666 = ~n13041 | ~n14663;
  assign n12407 = ~n15016 | ~n14552;
  assign n14544 = ~n13090 ^ n12407;
  assign n12416 = ~n14544 & ~n16337;
  assign n12414 = n14545 | n16309;
  assign n12408 = n15496 & P1_B_REG_SCAN_IN;
  assign n12690 = n16025 | n12408;
  assign n12413 = ~n12690;
  assign n12410 = ~n11286 | ~P1_REG1_REG_31__SCAN_IN;
  assign n12409 = ~n8988 | ~P1_REG2_REG_31__SCAN_IN;
  assign n12412 = ~n12410 | ~n12409;
  assign n12411 = n11852 & P1_REG0_REG_31__SCAN_IN;
  assign n14546 = ~n12413 | ~n16426;
  assign n12415 = ~n12414 | ~n14546;
  assign n12418 = ~n12419 | ~n16395;
  assign n12417 = ~n16393 | ~P1_REG1_REG_31__SCAN_IN;
  assign P1_U3554 = ~n12418 | ~n12417;
  assign n12421 = ~n12419 | ~n16363;
  assign n12420 = ~n16349 | ~P1_REG0_REG_31__SCAN_IN;
  assign P1_U3522 = ~n12421 | ~n12420;
  assign n12426 = ~n12423 | ~n12422;
  assign n12425 = ~n12424 | ~n17227;
  assign n12428 = ~n12426 | ~n12425;
  assign n12432 = ~n12445 ^ n12429;
  assign n12433 = n12431 & n12430;
  assign n12437 = n12432 | n12433;
  assign n12434 = ~n12433 | ~n12432;
  assign n12436 = ~n17197 | ~n12487;
  assign n12435 = ~n12445 | ~n17365;
  assign n16486 = ~n12436 | ~n12435;
  assign n16598 = n12438 & n12437;
  assign n12440 = ~n12624 ^ n12439;
  assign n12441 = n16463 & n12487;
  assign n16600 = n12440 | n12441;
  assign n12444 = ~n16598 | ~n16600;
  assign n12443 = ~n12440;
  assign n12442 = ~n12441;
  assign n16599 = n12443 | n12442;
  assign n16460 = n12444 & n16599;
  assign n12446 = ~n12624 ^ n17399;
  assign n12447 = ~n12487 | ~n16541;
  assign n16458 = n12446 | n12447;
  assign n12450 = ~n16460 | ~n16458;
  assign n12449 = ~n12446;
  assign n12448 = ~n12447;
  assign n16459 = n12449 | n12448;
  assign n16536 = n12450 & n16459;
  assign n12451 = ~n12624 ^ n17133;
  assign n12452 = n12487 & n16517;
  assign n16538 = n12451 | n12452;
  assign n12455 = ~n16536 | ~n16538;
  assign n12454 = ~n12451;
  assign n12453 = ~n12452;
  assign n16537 = n12454 | n12453;
  assign n12458 = ~n12624 ^ n17419;
  assign n12457 = n12487 & n16625;
  assign n16522 = n12458 & n12457;
  assign n16523 = n12458 | n12457;
  assign n12461 = n12459 & n12487;
  assign n12465 = n12460 | n12461;
  assign n12463 = ~n12460;
  assign n12462 = ~n12461;
  assign n12464 = n12463 | n12462;
  assign n16621 = n12465 & n12464;
  assign n12468 = ~n17443 ^ n12624;
  assign n12466 = n16627 & n12487;
  assign n16431 = ~n12468 ^ n12466;
  assign n12467 = ~n12466;
  assign n12469 = n12468 | n12467;
  assign n12470 = ~n17041 ^ n12524;
  assign n12471 = ~n12487 | ~n16558;
  assign n16475 = ~n12470 ^ n12471;
  assign n12472 = ~n12470;
  assign n12473 = n12472 | n12471;
  assign n16550 = ~n12474 | ~n12473;
  assign n12475 = ~n17465 ^ n12524;
  assign n12476 = n12487 & n16477;
  assign n16552 = n12475 | n12476;
  assign n12478 = ~n12475;
  assign n12477 = ~n12476;
  assign n16551 = n12478 | n12477;
  assign n12479 = ~n17476 ^ n12524;
  assign n12480 = ~n12487 | ~n16559;
  assign n16446 = ~n12479 ^ n12480;
  assign n12481 = ~n12479;
  assign n12482 = n12481 | n12480;
  assign n12483 = ~n16955 ^ n12524;
  assign n12484 = n16505 & n12487;
  assign n12486 = ~n12483;
  assign n12485 = ~n12484;
  assign n16582 = n12486 | n12485;
  assign n12488 = ~n17505 ^ n12524;
  assign n12489 = n12487 & n16592;
  assign n16500 = n12488 | n12489;
  assign n12491 = ~n12488;
  assign n12490 = ~n12489;
  assign n12493 = ~n13920 ^ n12524;
  assign n12492 = n16506 & n12487;
  assign n13433 = n12493 | n12492;
  assign n13309 = ~n12494 | ~n13433;
  assign n12495 = ~n14114 ^ n12524;
  assign n12496 = ~n13935 | ~n12487;
  assign n13310 = ~n12495 ^ n12496;
  assign n13307 = ~n13309 | ~n13310;
  assign n13372 = ~n14102 ^ n12624;
  assign n12497 = ~n12495;
  assign n12498 = n12497 & n12496;
  assign n13374 = n13372 | n12498;
  assign n13371 = ~n12498;
  assign n12499 = ~n13371 | ~n13491;
  assign n12500 = ~n13374 | ~n12499;
  assign n12509 = ~n13307 | ~n12500;
  assign n12501 = ~n13384 ^ n12524;
  assign n12502 = ~n13871 | ~n12487;
  assign n12510 = ~n12501 | ~n12502;
  assign n12504 = ~n12501;
  assign n12503 = ~n12502;
  assign n12505 = ~n12504 | ~n12503;
  assign n13377 = ~n12510 | ~n12505;
  assign n12506 = ~n13372;
  assign n12507 = n12506 & n13491;
  assign n12508 = ~n13377 & ~n12507;
  assign n12513 = ~n12512;
  assign n12514 = ~n12513 | ~n9004;
  assign n12516 = ~n12487 | ~n13395;
  assign n13459 = ~n12515 ^ n12516;
  assign n12517 = ~n12515;
  assign n12519 = ~n14060 ^ n12524;
  assign n12518 = n17558 & n12487;
  assign n13345 = n12519 | n12518;
  assign n12521 = ~n12487 | ~n17561;
  assign n13420 = ~n12522 ^ n12521;
  assign n12520 = ~n13420;
  assign n12523 = n12522 | n12521;
  assign n12525 = ~n14038 ^ n12524;
  assign n12526 = ~n12487 | ~n17564;
  assign n13358 = ~n12525 ^ n12526;
  assign n12527 = ~n12525;
  assign n12528 = n12527 | n12526;
  assign n13445 = ~n17567 | ~n12487;
  assign n12529 = ~n12532;
  assign n12530 = ~n14017 ^ n12624;
  assign n12531 = ~n12530;
  assign n13331 = ~n17570 | ~n12487;
  assign n12533 = ~n13329 & ~n13331;
  assign n13406 = ~n17573 | ~n12487;
  assign n12535 = ~n13405 & ~n13406;
  assign n12537 = ~n13995 ^ n12624;
  assign n12536 = ~n17576 | ~n12487;
  assign n12611 = ~n12537 | ~n12536;
  assign n12613 = n12537 | n12536;
  assign n12579 = ~n12538 ^ n9967;
  assign n12539 = P2_B_REG_SCAN_IN ^ n17352;
  assign n12573 = ~n12569 | ~n12539;
  assign n12545 = ~P2_D_REG_6__SCAN_IN & ~P2_D_REG_7__SCAN_IN;
  assign n12543 = P2_D_REG_8__SCAN_IN | P2_D_REG_9__SCAN_IN;
  assign n12541 = ~P2_D_REG_10__SCAN_IN & ~P2_D_REG_11__SCAN_IN;
  assign n12540 = ~P2_D_REG_12__SCAN_IN & ~P2_D_REG_13__SCAN_IN;
  assign n12542 = ~n12541 | ~n12540;
  assign n12544 = ~n12543 & ~n12542;
  assign n12561 = ~n12545 | ~n12544;
  assign n12547 = ~P2_D_REG_18__SCAN_IN & ~P2_D_REG_19__SCAN_IN;
  assign n12546 = ~P2_D_REG_20__SCAN_IN & ~P2_D_REG_21__SCAN_IN;
  assign n12551 = ~n12547 | ~n12546;
  assign n12549 = ~P2_D_REG_16__SCAN_IN & ~P2_D_REG_14__SCAN_IN;
  assign n12548 = ~P2_D_REG_15__SCAN_IN & ~P2_D_REG_17__SCAN_IN;
  assign n12550 = ~n12549 | ~n12548;
  assign n12559 = ~n12551 & ~n12550;
  assign n12553 = ~P2_D_REG_26__SCAN_IN & ~P2_D_REG_27__SCAN_IN;
  assign n12552 = ~P2_D_REG_28__SCAN_IN & ~P2_D_REG_31__SCAN_IN;
  assign n12557 = ~n12553 | ~n12552;
  assign n12555 = ~P2_D_REG_22__SCAN_IN & ~P2_D_REG_23__SCAN_IN;
  assign n12554 = ~P2_D_REG_24__SCAN_IN & ~P2_D_REG_25__SCAN_IN;
  assign n12556 = ~n12555 | ~n12554;
  assign n12558 = ~n12557 & ~n12556;
  assign n12560 = ~n12559 | ~n12558;
  assign n12566 = ~n12561 & ~n12560;
  assign n12563 = ~P2_D_REG_2__SCAN_IN & ~P2_D_REG_3__SCAN_IN;
  assign n12562 = ~P2_D_REG_4__SCAN_IN & ~P2_D_REG_5__SCAN_IN;
  assign n12564 = ~n12563 | ~n12562;
  assign n12565 = ~P2_D_REG_30__SCAN_IN & ~n12564;
  assign n12567 = ~n12566 | ~n12565;
  assign n12568 = ~P2_D_REG_29__SCAN_IN & ~n12567;
  assign n12570 = ~n12569;
  assign n17357 = ~n17351 & ~n12570;
  assign n12576 = ~n17352 | ~n14220;
  assign n12572 = ~P2_D_REG_0__SCAN_IN;
  assign n12574 = ~n12573 | ~n12572;
  assign n12575 = ~n12574 | ~n17351;
  assign n12577 = ~n13510 | ~n13948;
  assign n12578 = ~n14113 & ~n12584;
  assign n12606 = ~n12579 | ~n16575;
  assign n12583 = ~n12597 | ~n17191;
  assign n12604 = ~n13622 & ~n16617;
  assign n12585 = ~n12584 | ~n12595;
  assign n13286 = ~n12586 | ~n12585;
  assign n12587 = ~n13317 & ~n14113;
  assign n12589 = ~n13286 & ~n12587;
  assign n12590 = ~n12589 | ~n12588;
  assign n13321 = ~P2_STATE_REG_SCAN_IN | ~n12590;
  assign n12591 = ~n13317 & ~P2_U3152;
  assign n12592 = ~n17191 | ~n12591;
  assign n13475 = ~n13321 | ~n12592;
  assign n12594 = ~n13475 | ~n13623;
  assign n12593 = ~P2_REG3_REG_25__SCAN_IN | ~P2_U3152;
  assign n12602 = n12594 & n12593;
  assign n12596 = ~n12595;
  assign n13314 = ~n13260 & ~n12598;
  assign n12600 = ~n17579 | ~n16628;
  assign n12599 = ~n17573 | ~n16626;
  assign n13612 = ~n12600 | ~n12599;
  assign n12601 = ~n16631 | ~n13612;
  assign n12603 = ~n12602 | ~n12601;
  assign n12605 = ~n12604 & ~n12603;
  assign P2_U3227 = ~n12606 | ~n12605;
  assign n12607 = ~n12610 | ~n13406;
  assign n12608 = ~n12611 | ~n12607;
  assign n12612 = ~n12610 & ~n13406;
  assign n12614 = ~n12612 | ~n12611;
  assign n12615 = ~n12614 | ~n12613;
  assign n12617 = ~n13984 ^ n12624;
  assign n12616 = ~n17579 | ~n12487;
  assign n13472 = ~n12617 ^ n12616;
  assign n12620 = n12624 ^ n13974;
  assign n12618 = ~n12487 | ~n17582;
  assign n13295 = ~n12620 ^ n12618;
  assign n12622 = ~n13294 | ~n13295;
  assign n12619 = ~n12618;
  assign n12621 = ~n12620 | ~n12619;
  assign n12623 = ~n12487 | ~n17585;
  assign n12630 = ~n12624 ^ n12623;
  assign n12625 = ~n16617 | ~n12630;
  assign n12627 = ~n9749 & ~n12625;
  assign n12626 = ~n13964 & ~n12630;
  assign n12628 = ~n9749 & ~n16617;
  assign n12633 = ~n9749 | ~n12630;
  assign n12631 = ~n16569 & ~n12630;
  assign n12632 = ~n13964 | ~n12631;
  assign n12634 = ~n12633 | ~n12632;
  assign n12635 = ~n12629 | ~n12634;
  assign n12637 = n16605 | n13255;
  assign n12636 = ~n16628 | ~n17588;
  assign n13543 = n12637 & n12636;
  assign n12641 = ~n16608 & ~n13543;
  assign n12639 = ~n13475 | ~n13547;
  assign n12638 = ~P2_U3152 | ~P2_REG3_REG_28__SCAN_IN;
  assign n12640 = ~n12639 | ~n12638;
  assign n12642 = ~n12641 & ~n12640;
  assign P2_U3222 = ~n12643 | ~n12642;
  assign n12810 = ~n15209 | ~n14964;
  assign n12925 = n15198 | n14993;
  assign n14958 = n15209 | n14964;
  assign n12753 = n12925 & n14958;
  assign n12933 = ~n15198 | ~n14993;
  assign n12955 = ~n15188 | ~n14965;
  assign n14916 = ~n15177 ^ n14937;
  assign n12756 = ~n15177 & ~n14937;
  assign n12940 = n15166 & n14364;
  assign n12662 = ~n14363 | ~n14533;
  assign n14854 = n15166 | n14364;
  assign n12766 = ~n12662 | ~n14854;
  assign n14885 = ~n14533;
  assign n12975 = ~n15145 | ~n14804;
  assign n12989 = n15134 | n14828;
  assign n14800 = ~n14843 | ~n14859;
  assign n12990 = ~n15134 | ~n14828;
  assign n14803 = ~n14509;
  assign n12777 = n15123 | n14803;
  assign n12727 = ~n15123 | ~n14803;
  assign n14331 = ~n16398;
  assign n14714 = ~n15091;
  assign n12796 = ~n14714 | ~n16398;
  assign n14468 = ~n16401;
  assign n12795 = ~n15080 & ~n14468;
  assign n13167 = ~n15080 | ~n14468;
  assign n12677 = ~n16404;
  assign n13171 = ~n15069 | ~n12677;
  assign n13177 = n15047 | n14586;
  assign n12793 = ~n15047 | ~n14586;
  assign n12722 = ~n15035 | ~n14609;
  assign n13074 = ~n15025 & ~n16416;
  assign n12649 = ~n13074;
  assign n12721 = n13082 | n14562;
  assign n13127 = ~n13082 | ~n14562;
  assign n12651 = ~n12650 ^ n12824;
  assign n12905 = n14296 | n14490;
  assign n12653 = n15209 | n12654;
  assign n12655 = ~n15209 | ~n12654;
  assign n14962 = ~n12925 | ~n12933;
  assign n12656 = ~n15198 | ~n14453;
  assign n12657 = n15188 | n14907;
  assign n12659 = ~n14936 | ~n12657;
  assign n12658 = ~n15188 | ~n14907;
  assign n12799 = n15166 | n14908;
  assign n12798 = ~n15166 | ~n14908;
  assign n14867 = ~n12662 | ~n9035;
  assign n14833 = ~n15155 | ~n14533;
  assign n12981 = ~n15145 | ~n14859;
  assign n12663 = n14833 & n12981;
  assign n12814 = ~n14843 | ~n14804;
  assign n14809 = ~n12989 | ~n12990;
  assign n12666 = n15123 | n14509;
  assign n12665 = n14809 & n12666;
  assign n12667 = ~n12666;
  assign n14786 = ~n15134 | ~n14775;
  assign n12668 = n15112 | n14774;
  assign n12669 = ~n15112 | ~n14774;
  assign n12670 = ~n13020;
  assign n14730 = ~n12670 | ~n13021;
  assign n12671 = ~n15101 | ~n14703;
  assign n12672 = ~n14714 | ~n14331;
  assign n12673 = ~n15091 | ~n16398;
  assign n12675 = n15080 & n16401;
  assign n12676 = n15080 | n16401;
  assign n13043 = ~n15069 | ~n16404;
  assign n13048 = ~n13041 | ~n12677;
  assign n14641 = ~n14605 | ~n13175;
  assign n12679 = n15059 | n16407;
  assign n12681 = ~n15047 | ~n16410;
  assign n12682 = n15047 | n16410;
  assign n12683 = n15035 | n16413;
  assign n12720 = ~n13075;
  assign n12685 = n15025 | n14587;
  assign n12692 = ~n14587 & ~n16023;
  assign n12687 = ~n8988 | ~P1_REG2_REG_30__SCAN_IN;
  assign n12686 = ~n11852 | ~P1_REG0_REG_30__SCAN_IN;
  assign n12689 = ~n12687 | ~n12686;
  assign n12688 = n11286 & P1_REG1_REG_30__SCAN_IN;
  assign n16422 = n12689 | n12688;
  assign n13125 = ~n16422;
  assign n12691 = ~n13125 & ~n12690;
  assign n12699 = ~n12694 & ~n16357;
  assign n12710 = n12695 ^ n13082;
  assign n12697 = ~n12710 | ~n16350;
  assign n12696 = ~n13082 | ~n16352;
  assign n12698 = ~n12697 | ~n12696;
  assign n12702 = ~n12703 | ~n16395;
  assign n12701 = ~n16393 | ~P1_REG1_REG_29__SCAN_IN;
  assign P1_U3552 = ~n12702 | ~n12701;
  assign n12705 = ~n12703 | ~n16363;
  assign n12704 = ~n16349 | ~P1_REG0_REG_29__SCAN_IN;
  assign P1_U3520 = ~n12705 | ~n12704;
  assign n12708 = ~n12706 | ~n16119;
  assign n12707 = n16119 | P1_REG2_REG_29__SCAN_IN;
  assign n12719 = ~n12708 | ~n12707;
  assign n12717 = ~n12694 & ~n16003;
  assign n15940 = n16245 | n12709;
  assign n12715 = ~n12710 | ~n16109;
  assign n12713 = ~n13082 | ~n16108;
  assign n12712 = ~n16105 | ~n12711;
  assign n12714 = n12713 & n12712;
  assign n12716 = ~n12715 | ~n12714;
  assign n12718 = ~n12717 & ~n12716;
  assign P1_U3355 = ~n12719 | ~n12718;
  assign n13085 = ~n16426;
  assign n13094 = ~n13125 & ~n13085;
  assign n13183 = ~n12721 | ~n12720;
  assign n12723 = ~n12722;
  assign n13131 = n13074 | n12723;
  assign n12724 = ~n12793;
  assign n13129 = ~n12788 | ~n12724;
  assign n12797 = ~n12725;
  assign n12728 = ~n12727;
  assign n12729 = n12975 & n9035;
  assign n12767 = ~n12990 | ~n12729;
  assign n12730 = n15177 & n14937;
  assign n12751 = ~n12940 & ~n12730;
  assign n15839 = ~n12731;
  assign n12808 = n12732 | n15839;
  assign n12734 = ~n12761 & ~n9895;
  assign n12735 = ~n12751 | ~n12734;
  assign n13160 = ~n12767 & ~n12735;
  assign n12738 = ~n12868;
  assign n15917 = n12737 | n12736;
  assign n12739 = ~n12738 & ~n15917;
  assign n12740 = ~n12739 | ~n13154;
  assign n12741 = ~n12740 & ~n9596;
  assign n12749 = ~n12741 | ~n16021;
  assign n12743 = n15918 | n13143;
  assign n12744 = ~n12743 | ~n12742;
  assign n12745 = n12744 | n15920;
  assign n12746 = n12745 & n13148;
  assign n12747 = ~n12746 | ~n13149;
  assign n13153 = n12882 & n12868;
  assign n12748 = ~n12747 | ~n13153;
  assign n12750 = n12749 & n12748;
  assign n12768 = ~n13160 | ~n12750;
  assign n12765 = ~n12751;
  assign n12752 = ~n12933;
  assign n12754 = ~n12753 & ~n12752;
  assign n12755 = ~n12754 | ~n12955;
  assign n12757 = ~n12755 | ~n12959;
  assign n12763 = n12757 | n12756;
  assign n12758 = ~n12895 | ~n12804;
  assign n12760 = ~n12759 & ~n12758;
  assign n12762 = ~n12761 & ~n12760;
  assign n12764 = ~n12763 & ~n12762;
  assign n12770 = n13167 & n12769;
  assign n12772 = n12771 & n9904;
  assign n12785 = n12772 & n13169;
  assign n12773 = ~n12990;
  assign n12775 = ~n12774 & ~n12773;
  assign n12783 = ~n13164 | ~n12775;
  assign n12780 = ~n12776;
  assign n12778 = ~n12997 | ~n12777;
  assign n12779 = n13020 | n12778;
  assign n12781 = ~n12780 | ~n12779;
  assign n12782 = n12781 & n12796;
  assign n12784 = ~n13132 | ~n13167;
  assign n12787 = ~n12785 | ~n12784;
  assign n12786 = n13175 & n13171;
  assign n12790 = ~n13131 & ~n12789;
  assign n13123 = n13126 | n13125;
  assign n13189 = n14545 & n16426;
  assign n13122 = ~n14545 & ~n16426;
  assign n12827 = ~n12792 & ~n9500;
  assign n14614 = ~n13177 | ~n12793;
  assign n12794 = ~n13167;
  assign n14690 = n12795 | n12794;
  assign n14680 = ~n14690;
  assign n14710 = ~n12797 | ~n12796;
  assign n14756 = ~n12997 | ~n13010;
  assign n12816 = ~n14809;
  assign n12958 = ~n12799 | ~n12798;
  assign n14883 = ~n12958;
  assign n13135 = n16078 & n16244;
  assign n16115 = ~n16071 & ~n13135;
  assign n12801 = ~n16115 | ~n12800;
  assign n12803 = n12801 | n16051;
  assign n12802 = ~n15989 & ~n16020;
  assign n15840 = ~n12804;
  assign n12807 = ~n12806 | ~n12805;
  assign n12809 = ~n12808;
  assign n14991 = ~n14958 | ~n12810;
  assign n12812 = ~n12811 | ~n14935;
  assign n12813 = ~n14916;
  assign n14835 = ~n12814 | ~n12981;
  assign n12817 = ~n12816 | ~n12815;
  assign n12818 = ~n14756 & ~n12817;
  assign n12819 = ~n12818 | ~n14789;
  assign n12821 = ~n12820 | ~n14660;
  assign n12822 = ~n14614 & ~n12821;
  assign n12823 = ~n13180 | ~n12822;
  assign n12825 = ~n13189 & ~n12824;
  assign n12828 = ~n12827 & ~n13104;
  assign n12832 = ~n12831 | ~n13134;
  assign n12833 = ~n16261 | ~n8987;
  assign n12837 = ~n12835;
  assign n12836 = ~n16076 | ~n15420;
  assign n12838 = ~n12837 | ~n12836;
  assign n12842 = n16014 & n12902;
  assign n12840 = ~n12847 | ~n12842;
  assign n12841 = ~n12840 | ~n13003;
  assign n15388 = ~n16046;
  assign n12846 = ~n12841 | ~n15388;
  assign n12844 = ~n12847 | ~n16274;
  assign n12843 = ~n12842;
  assign n12845 = ~n12844 | ~n12843;
  assign n12849 = ~n12847;
  assign n12848 = n16014 & n8987;
  assign n12854 = ~n12849 | ~n12848;
  assign n12851 = n15972 | n8987;
  assign n12850 = ~n16283 | ~n8987;
  assign n12860 = ~n12851 | ~n12850;
  assign n12853 = ~n12860 | ~n12852;
  assign n12855 = n12854 & n12853;
  assign n12867 = ~n12856 | ~n12855;
  assign n12858 = n15930 | n8987;
  assign n12857 = ~n15961 | ~n8987;
  assign n12871 = n12858 & n12857;
  assign n12865 = ~n12871 | ~n12859;
  assign n12863 = ~n12860;
  assign n12862 = ~n15972 | ~n12861;
  assign n12864 = ~n12863 | ~n12862;
  assign n12866 = n12865 & n12864;
  assign n12877 = ~n12867 | ~n12866;
  assign n12870 = ~n13149 | ~n13003;
  assign n12869 = ~n12868 | ~n8987;
  assign n12875 = ~n12870 | ~n12869;
  assign n12873 = ~n12871;
  assign n12872 = n16296 | n15930;
  assign n12874 = ~n12873 | ~n12872;
  assign n12876 = n12875 & n12874;
  assign n12879 = n15326 | n8987;
  assign n12878 = ~n15946 | ~n8987;
  assign n12881 = ~n12879 | ~n12878;
  assign n12880 = n16310 | n15326;
  assign n12884 = ~n12882 | ~n8987;
  assign n12883 = ~n15861 | ~n13003;
  assign n12885 = ~n12884 | ~n12883;
  assign n12887 = n16320 | n8987;
  assign n12886 = ~n15437 | ~n8987;
  assign n12889 = ~n12887 | ~n12886;
  assign n12890 = ~n12889 | ~n12888;
  assign n12892 = ~n12895 | ~n8987;
  assign n12891 = ~n12896 | ~n13003;
  assign n12893 = ~n12892 | ~n12891;
  assign n12898 = ~n12895 | ~n13003;
  assign n12897 = ~n12896 | ~n8987;
  assign n12899 = ~n12898 | ~n12897;
  assign n13003 = n12902;
  assign n12901 = n16353 | n13003;
  assign n12900 = ~n12908 | ~n13003;
  assign n12907 = n12901 & n12900;
  assign n12904 = n14296 | n13003;
  assign n12903 = ~n15847 | ~n13003;
  assign n12913 = ~n12904 | ~n12903;
  assign n12906 = ~n12913 | ~n12905;
  assign n12910 = ~n16353 | ~n13003;
  assign n12909 = n12908 | n13003;
  assign n12911 = ~n12910 | ~n12909;
  assign n12912 = n14296 & n14490;
  assign n12922 = n12913 | n12912;
  assign n12915 = n15209 | n13003;
  assign n12914 = ~n14964 | ~n13003;
  assign n12921 = n12915 & n12914;
  assign n12920 = ~n12916 | ~n12921;
  assign n12918 = ~n15209 | ~n13003;
  assign n12917 = n14964 | n13003;
  assign n12919 = ~n12918 | ~n12917;
  assign n12931 = ~n12920 | ~n12919;
  assign n12923 = ~n12921;
  assign n12924 = n12923 & n12922;
  assign n12927 = ~n12925 | ~n8987;
  assign n12926 = ~n12933 | ~n13003;
  assign n12928 = ~n12927 | ~n12926;
  assign n12930 = n12929 & n12928;
  assign n12932 = n15198 | n8987;
  assign n12935 = ~n12933 | ~n12932;
  assign n12934 = ~n14993 | ~n13003;
  assign n12937 = ~n14363 | ~n13003;
  assign n12936 = n14533 | n13003;
  assign n12971 = n12937 & n12936;
  assign n12939 = ~n14363 | ~n8987;
  assign n12938 = n14533 | n8987;
  assign n12970 = ~n12939 | ~n12938;
  assign n12944 = ~n12971 | ~n12970;
  assign n12942 = n12940 | n8987;
  assign n12941 = ~n14854 | ~n8987;
  assign n12943 = ~n12942 | ~n12941;
  assign n12969 = ~n12944 | ~n12943;
  assign n12946 = n15177 | n8987;
  assign n12945 = ~n14937 | ~n8987;
  assign n12963 = ~n12946 | ~n12945;
  assign n12948 = ~n15177 | ~n8987;
  assign n12947 = n14937 | n8987;
  assign n12962 = ~n12948 | ~n12947;
  assign n12952 = n12963 | n12962;
  assign n12950 = ~n12959 | ~n8987;
  assign n12949 = ~n12955 | ~n13003;
  assign n12951 = ~n12950 | ~n12949;
  assign n12953 = ~n12952 | ~n12951;
  assign n12954 = ~n12969 & ~n12953;
  assign n12957 = n12963 | n15177;
  assign n12956 = ~n12955 & ~n13003;
  assign n12960 = ~n12959 & ~n8987;
  assign n12965 = ~n12961 | ~n12960;
  assign n12964 = ~n12963 | ~n12962;
  assign n12966 = ~n12965 | ~n12964;
  assign n12968 = ~n12967 & ~n12966;
  assign n12973 = ~n12969 & ~n12968;
  assign n12972 = ~n12971 & ~n12970;
  assign n12977 = ~n14800 | ~n8987;
  assign n12976 = ~n12975 | ~n13003;
  assign n12978 = ~n12977 | ~n12976;
  assign n12980 = ~n15145 | ~n8987;
  assign n12979 = n14804 | n8987;
  assign n12982 = ~n12980 | ~n12979;
  assign n12983 = ~n12982 | ~n12981;
  assign n12988 = ~n12984 | ~n12983;
  assign n12986 = ~n12989 | ~n8987;
  assign n12985 = ~n12990 | ~n13003;
  assign n12987 = ~n12986 | ~n12985;
  assign n12992 = ~n12989 | ~n13003;
  assign n12991 = ~n12990 | ~n8987;
  assign n12993 = ~n12992 | ~n12991;
  assign n12996 = n15123 | n8987;
  assign n12995 = n14509 | n13003;
  assign n13001 = ~n12996 | ~n12995;
  assign n12999 = ~n12997 | ~n8987;
  assign n12998 = ~n13010 | ~n13003;
  assign n13000 = ~n12999 | ~n12998;
  assign n13007 = ~n13002 | ~n13001;
  assign n13005 = n15123 | n13003;
  assign n13004 = n14509 | n8987;
  assign n13006 = ~n13005 | ~n13004;
  assign n13008 = ~n13007 | ~n13006;
  assign n13009 = n15112 | n8987;
  assign n13013 = ~n13010 | ~n13009;
  assign n13012 = ~n13011 | ~n13003;
  assign n13014 = ~n13013 | ~n13012;
  assign n13019 = ~n13015 | ~n13014;
  assign n13016 = ~n13021 | ~n13003;
  assign n13018 = ~n13017 | ~n13016;
  assign n13025 = ~n13019 | ~n13018;
  assign n13023 = n13020 | n8987;
  assign n13022 = ~n13021 | ~n8987;
  assign n13024 = ~n13023 | ~n13022;
  assign n13027 = n15091 | n8987;
  assign n13026 = ~n14331 | ~n8987;
  assign n13028 = ~n13027 | ~n13026;
  assign n13030 = n15091 | n13003;
  assign n13029 = ~n14331 | ~n13003;
  assign n13031 = ~n13030 | ~n13029;
  assign n13033 = n15080 | n13003;
  assign n13032 = ~n14468 | ~n13003;
  assign n13038 = n13033 & n13032;
  assign n13035 = n15080 | n8987;
  assign n13034 = ~n14468 | ~n8987;
  assign n13037 = ~n13035 | ~n13034;
  assign n13036 = ~n13038 | ~n13037;
  assign n13040 = ~n13037;
  assign n13039 = ~n13038;
  assign n13042 = n16404 | n8987;
  assign n13046 = ~n14605 | ~n8987;
  assign n13045 = ~n13175 | ~n13003;
  assign n13051 = ~n13046 | ~n13045;
  assign n13050 = ~n13049 | ~n13048;
  assign n13052 = n13051 & n13050;
  assign n13054 = ~n14605 | ~n13003;
  assign n13053 = ~n13175 | ~n8987;
  assign n13055 = ~n13054 | ~n13053;
  assign n13057 = n15047 | n8987;
  assign n13056 = n16410 | n13003;
  assign n13058 = ~n13057 | ~n13056;
  assign n13060 = n15047 | n13003;
  assign n13059 = n16410 | n8987;
  assign n13061 = ~n13060 | ~n13059;
  assign n13067 = n16413 | n13003;
  assign n13063 = n13068 & n13067;
  assign n13066 = n15035 | n13003;
  assign n13065 = n16413 | n8987;
  assign n13062 = ~n13066 | ~n13065;
  assign n13070 = n13066 & n13065;
  assign n13069 = ~n13068 | ~n13067;
  assign n13071 = ~n13070 | ~n13069;
  assign n13072 = n14567 & n13071;
  assign n13079 = ~n13073 | ~n13072;
  assign n13077 = n13074 | n8987;
  assign n13076 = n13075 | n13003;
  assign n13078 = ~n13077 | ~n13076;
  assign n13081 = n13082 | n13003;
  assign n13080 = n16419 | n8987;
  assign n13084 = ~n13082 & ~n8987;
  assign n13083 = ~n16419 & ~n13003;
  assign n13086 = ~n13085 & ~n16422;
  assign n13087 = ~n14545 & ~n13086;
  assign n13089 = ~n13087 | ~n15016;
  assign n13088 = ~n13098;
  assign n13093 = ~n13090 & ~n16426;
  assign n13091 = ~n16426 & ~n8987;
  assign n13092 = ~n14545 & ~n13091;
  assign n13097 = ~n13093 & ~n13092;
  assign n13095 = ~n13094 | ~n13003;
  assign n13096 = ~n13126 & ~n13095;
  assign n13101 = ~n13097 & ~n13096;
  assign n13099 = ~n13122 & ~n13003;
  assign n13100 = ~n13099 | ~n13098;
  assign n13108 = ~n13107 | ~n9504;
  assign n13111 = ~n11945 & ~n15494;
  assign n13118 = ~n13112 | ~n13111;
  assign n13116 = ~n13114 & ~n13113;
  assign n13115 = ~P1_B_REG_SCAN_IN;
  assign n13117 = ~n13116 & ~n13115;
  assign n13200 = ~n13118 | ~n13117;
  assign n13119 = ~n13200;
  assign n13124 = ~n13122;
  assign n13188 = n13124 & n13123;
  assign n13128 = ~n13126 | ~n13125;
  assign n13187 = n13128 & n13127;
  assign n13130 = ~n13129;
  assign n13182 = ~n13131 & ~n13130;
  assign n13138 = ~n13134;
  assign n13136 = ~n13135;
  assign n13137 = ~n13136 | ~n9504;
  assign n13139 = ~n13138 & ~n13137;
  assign n13141 = n13133 | n13139;
  assign n13145 = ~n13141 | ~n13140;
  assign n13144 = ~n13143 & ~n9418;
  assign n13147 = ~n13145 | ~n13144;
  assign n13146 = ~n15917;
  assign n13152 = ~n13147 | ~n13146;
  assign n15921 = ~n13148;
  assign n13150 = ~n15918 & ~n15921;
  assign n13151 = n13150 & n13149;
  assign n13158 = ~n13152 | ~n13151;
  assign n13156 = ~n13153;
  assign n13155 = ~n13154;
  assign n13157 = ~n13156 & ~n13155;
  assign n13159 = ~n13158 | ~n13157;
  assign n13162 = ~n13160 | ~n13159;
  assign n13163 = ~n13162 | ~n13161;
  assign n13165 = ~n13164 | ~n13163;
  assign n13166 = n13165 & n9904;
  assign n13170 = ~n13168 | ~n13167;
  assign n13172 = ~n13170 | ~n13169;
  assign n13173 = ~n13172 | ~n13171;
  assign n13176 = ~n13175;
  assign n13178 = ~n13177 | ~n13176;
  assign n13181 = ~n13180 | ~n13179;
  assign n13185 = ~n13182 | ~n13181;
  assign n13184 = ~n13183;
  assign n13186 = ~n13185 | ~n13184;
  assign n13194 = ~n13190 | ~n9350;
  assign n13193 = ~n13194 | ~n13191;
  assign n13196 = ~n13193 | ~n13192;
  assign n13195 = ~n13194 & ~n16125;
  assign n13199 = ~n13198 | ~n13197;
  assign n13201 = n13200 & n13199;
  assign P1_U3240 = ~n13202 & ~n13201;
  assign n13203 = ~n17197 | ~n12430;
  assign n17169 = ~n17197;
  assign n13205 = ~n17169 | ~n10027;
  assign n13206 = ~n13205 | ~n17373;
  assign n13209 = ~n13207 | ~n13206;
  assign n13208 = ~n16489 | ~n12439;
  assign n17143 = ~n13209 | ~n13208;
  assign n13210 = ~n16603 | ~n17141;
  assign n13213 = ~n16625 | ~n17095;
  assign n13216 = ~n17105 | ~n13213;
  assign n13215 = ~n13214 | ~n17419;
  assign n17077 = ~n13216 | ~n13215;
  assign n13218 = n17443 | n16627;
  assign n13221 = ~n17015;
  assign n13222 = n17465 | n16477;
  assign n16960 = ~n13224 | ~n13223;
  assign n13225 = ~n16955 | ~n16505;
  assign n13227 = n17505 | n16592;
  assign n13228 = ~n13920 | ~n16506;
  assign n13826 = n14114 | n13935;
  assign n13229 = n13826 & n13230;
  assign n13233 = n13232 & n13231;
  assign n13236 = n14071 | n13395;
  assign n13238 = ~n14060 | ~n17558;
  assign n13239 = n14060 | n17558;
  assign n13243 = ~n13690 | ~n13656;
  assign n13247 = ~n13644 | ~n13655;
  assign n13248 = n13606 & n13587;
  assign n13584 = ~n13622 | ~n13249;
  assign n13474 = ~n13984;
  assign n13252 = ~n13474 | ~n13251;
  assign n13256 = ~n13572 | ~n13255;
  assign n13257 = ~n9749 | ~n13274;
  assign n13264 = ~n11082 & ~n17098;
  assign n13262 = ~n13260 | ~n13537;
  assign n13261 = n10825 | n13537;
  assign n13263 = ~n13262 | ~n13261;
  assign n13265 = n13537 & n17098;
  assign n17446 = ~n17173 | ~n17493;
  assign n13285 = ~n13539 | ~n17446;
  assign n13270 = ~n13266 ^ n13267;
  assign n13268 = n12424 | n13537;
  assign n13278 = ~n13270 | ~n17212;
  assign n13272 = n14214 | n13271;
  assign n13515 = ~n16628 | ~n13272;
  assign n13276 = ~n13515 & ~n13273;
  assign n13275 = ~n16605 & ~n13274;
  assign n13277 = ~n13276 & ~n13275;
  assign n13529 = ~n13278 | ~n13277;
  assign n17059 = ~n17074 | ~n17067;
  assign n17001 = ~n17465;
  assign n16984 = n17008 & n17001;
  assign n16953 = ~n16984 | ~n16442;
  assign n13909 = ~n14114;
  assign n13847 = n13845 | n14091;
  assign n13788 = ~n14071;
  assign n13666 = ~n14017;
  assign n13643 = ~n13665 | ~n13666;
  assign n13530 = ~n13280 ^ n13505;
  assign n17502 = ~n12581;
  assign n13282 = ~n13530 | ~n17502;
  assign n13281 = ~n13280 | ~n17504;
  assign n13283 = ~n13282 | ~n13281;
  assign n13284 = ~n13529 & ~n13283;
  assign n13288 = ~n13287 & ~n13286;
  assign n13508 = ~n17358 | ~n13288;
  assign n13289 = ~n13510 & ~n13508;
  assign n13292 = ~n17501 | ~P2_REG0_REG_29__SCAN_IN;
  assign P2_U3517 = ~n13293 | ~n13292;
  assign n13296 = n13295 ^ n13294;
  assign n13306 = ~n13296 | ~n16575;
  assign n13304 = ~n13974 | ~n16569;
  assign n13298 = ~n17579 | ~n16626;
  assign n13297 = ~n16628 | ~n17585;
  assign n13562 = n13298 & n13297;
  assign n13302 = ~n16608 & ~n13562;
  assign n13300 = ~n13475 | ~n13573;
  assign n13299 = ~P2_U3152 | ~P2_REG3_REG_27__SCAN_IN;
  assign n13301 = ~n13300 | ~n13299;
  assign n13303 = ~n13302 & ~n13301;
  assign n13305 = n13304 & n13303;
  assign P2_U3216 = ~n13306 | ~n13305;
  assign n13308 = n13307;
  assign n13312 = ~n13308;
  assign n13311 = ~n13309 & ~n13310;
  assign n13313 = ~n13312 & ~n13311;
  assign n13328 = ~n13313 & ~n16622;
  assign n16604 = ~n13314;
  assign n13462 = ~n13494;
  assign n13316 = ~n13462 & ~n13897;
  assign n13448 = ~n16631 | ~n16626;
  assign n13315 = ~n13448 & ~n13898;
  assign n13326 = ~n13316 & ~n13315;
  assign n13324 = ~n16617 & ~n13909;
  assign n13318 = ~n13317;
  assign n13319 = n17191 & n13318;
  assign n13320 = ~n17225 | ~n13319;
  assign n13322 = ~n16624 | ~n13910;
  assign n16816 = ~P2_REG3_REG_14__SCAN_IN | ~P2_U3152;
  assign n13323 = ~n13322 | ~n16816;
  assign n13325 = ~n13324 & ~n13323;
  assign n13327 = ~n13326 | ~n13325;
  assign P2_U3217 = n13328 | n13327;
  assign n13332 = ~n13330 & ~n13329;
  assign n13333 = ~n13332 ^ n13331;
  assign n13343 = ~n13333 | ~n16575;
  assign n13341 = ~n13666 & ~n16617;
  assign n13337 = ~n13448 & ~n13656;
  assign n13335 = ~n13475 | ~n13667;
  assign n13334 = ~P2_REG3_REG_23__SCAN_IN | ~P2_U3152;
  assign n13336 = ~n13335 | ~n13334;
  assign n13339 = ~n13337 & ~n13336;
  assign n13338 = ~n13494 | ~n17573;
  assign n13340 = ~n13339 | ~n13338;
  assign n13342 = ~n13341 & ~n13340;
  assign P2_U3218 = ~n13343 | ~n13342;
  assign n13346 = ~n9965 | ~n13345;
  assign n13347 = ~n13344 ^ n13346;
  assign n13357 = ~n13347 | ~n16575;
  assign n13351 = ~n13462 & ~n13752;
  assign n13348 = ~n13766;
  assign n13349 = ~n16624 | ~n13348;
  assign n16915 = ~P2_U3152 | ~P2_REG3_REG_19__SCAN_IN;
  assign n13350 = ~n13349 | ~n16915;
  assign n13353 = ~n13351 & ~n13350;
  assign n13352 = ~n13495 | ~n13395;
  assign n13355 = ~n13353 | ~n13352;
  assign n13354 = ~n9764 & ~n16617;
  assign n13356 = ~n13355 & ~n13354;
  assign P2_U3221 = ~n13357 | ~n13356;
  assign n13360 = n13359 ^ n13358;
  assign n13370 = ~n13360 | ~n16575;
  assign n13368 = ~n13714 & ~n16617;
  assign n13364 = ~n13462 & ~n13656;
  assign n13362 = ~n13475 | ~n13715;
  assign n13361 = ~P2_U3152 | ~P2_REG3_REG_21__SCAN_IN;
  assign n13363 = ~n13362 | ~n13361;
  assign n13366 = ~n13364 & ~n13363;
  assign n13365 = ~n13495 | ~n17561;
  assign n13367 = ~n13366 | ~n13365;
  assign n13369 = ~n13368 & ~n13367;
  assign P2_U3225 = ~n13370 | ~n13369;
  assign n13373 = ~n13308 | ~n13371;
  assign n13490 = ~n13373 | ~n13372;
  assign n13376 = ~n13490 | ~n13491;
  assign n13375 = ~n13374;
  assign n13489 = ~n13308 | ~n13375;
  assign n13378 = ~n13376 | ~n13489;
  assign n13380 = ~n13378 | ~n13377;
  assign n13381 = ~n13380 | ~n9494;
  assign n13391 = ~n13381 | ~n16575;
  assign n13383 = ~n13494 | ~n13838;
  assign n13382 = ~n13495 | ~n13837;
  assign n13389 = ~n13383 | ~n13382;
  assign n13387 = ~n16617 & ~n13384;
  assign n13385 = ~n16624 | ~n13856;
  assign n16852 = ~P2_REG3_REG_16__SCAN_IN | ~P2_U3152;
  assign n13386 = ~n13385 | ~n16852;
  assign n13388 = n13387 | n13386;
  assign n13390 = ~n13389 & ~n13388;
  assign P2_U3228 = ~n13391 | ~n13390;
  assign n13394 = n13392 ^ n13393;
  assign n13404 = ~n13394 | ~n16575;
  assign n13398 = ~n13494 | ~n13395;
  assign n13396 = ~n16624 | ~n13818;
  assign n16865 = ~P2_U3152 | ~P2_REG3_REG_17__SCAN_IN;
  assign n13397 = n13396 & n16865;
  assign n13402 = ~n13398 | ~n13397;
  assign n13400 = ~n13495 | ~n13871;
  assign n13399 = ~n16569 | ~n13279;
  assign n13401 = ~n13400 | ~n13399;
  assign n13403 = ~n13402 & ~n13401;
  assign P2_U3230 = ~n13404 | ~n13403;
  assign n13407 = n13406 ^ n13405;
  assign n13418 = ~n13407 | ~n16575;
  assign n13416 = ~n13644 & ~n16617;
  assign n13412 = ~n13448 & ~n13408;
  assign n13410 = ~n13475 | ~n13645;
  assign n13409 = ~P2_U3152 | ~P2_REG3_REG_24__SCAN_IN;
  assign n13411 = ~n13410 | ~n13409;
  assign n13414 = ~n13412 & ~n13411;
  assign n13413 = ~n13494 | ~n17576;
  assign n13415 = ~n13414 | ~n13413;
  assign n13417 = ~n13416 & ~n13415;
  assign P2_U3231 = ~n13418 | ~n13417;
  assign n13421 = n13420 ^ n13419;
  assign n13431 = ~n13421 | ~n16575;
  assign n13425 = ~n13462 & ~n13729;
  assign n13423 = ~n13475 | ~n13738;
  assign n13422 = ~P2_U3152 | ~P2_REG3_REG_20__SCAN_IN;
  assign n13424 = ~n13423 | ~n13422;
  assign n13427 = ~n13425 & ~n13424;
  assign n13426 = ~n13495 | ~n17558;
  assign n13429 = ~n13427 | ~n13426;
  assign n13428 = ~n9765 & ~n16617;
  assign n13430 = ~n13429 & ~n13428;
  assign P2_U3235 = ~n13431 | ~n13430;
  assign n13434 = ~n9968 | ~n13433;
  assign n13435 = ~n13432 ^ n13434;
  assign n13444 = ~n13435 | ~n16575;
  assign n13437 = ~n13494 | ~n13935;
  assign n13436 = ~n13495 | ~n16592;
  assign n13442 = ~n13437 | ~n13436;
  assign n13440 = ~n16617 & ~n14125;
  assign n13438 = ~n16624 | ~n13923;
  assign n16798 = ~P2_U3152 | ~P2_REG3_REG_13__SCAN_IN;
  assign n13439 = ~n13438 | ~n16798;
  assign n13441 = n13440 | n13439;
  assign n13443 = ~n13442 & ~n13441;
  assign P2_U3236 = ~n13444 | ~n13443;
  assign n13447 = ~n13446 ^ n13445;
  assign n13458 = ~n13447 | ~n16575;
  assign n13456 = ~n13690 & ~n16617;
  assign n13452 = ~n13448 & ~n13729;
  assign n13450 = ~n13475 | ~n13691;
  assign n13449 = ~P2_REG3_REG_22__SCAN_IN | ~P2_U3152;
  assign n13451 = ~n13450 | ~n13449;
  assign n13454 = ~n13452 & ~n13451;
  assign n13453 = ~n13494 | ~n17570;
  assign n13455 = ~n13454 | ~n13453;
  assign n13457 = ~n13456 & ~n13455;
  assign P2_U3237 = ~n13458 | ~n13457;
  assign n13461 = n13459 ^ n13460;
  assign n13471 = ~n13461 | ~n16575;
  assign n13465 = ~n13462 & ~n13777;
  assign n13463 = ~n16624 | ~n13789;
  assign n16891 = ~P2_U3152 | ~P2_REG3_REG_18__SCAN_IN;
  assign n13464 = ~n13463 | ~n16891;
  assign n13467 = ~n13465 & ~n13464;
  assign n13466 = ~n13495 | ~n13838;
  assign n13469 = ~n13467 | ~n13466;
  assign n13468 = ~n13788 & ~n16617;
  assign n13470 = ~n13469 & ~n13468;
  assign P2_U3240 = ~n13471 | ~n13470;
  assign n13473 = n13472 ^ n9040;
  assign n13488 = ~n13473 | ~n16575;
  assign n13486 = ~n13474 & ~n16617;
  assign n13477 = ~n13475;
  assign n13596 = ~n13476;
  assign n13480 = ~n13477 & ~n13596;
  assign n13479 = ~n13478 & ~P2_STATE_REG_SCAN_IN;
  assign n13484 = ~n13480 & ~n13479;
  assign n13482 = ~n17576 | ~n16626;
  assign n13481 = ~n16628 | ~n17582;
  assign n13590 = ~n13482 | ~n13481;
  assign n13483 = ~n16631 | ~n13590;
  assign n13485 = ~n13484 | ~n13483;
  assign n13487 = ~n13486 & ~n13485;
  assign P2_U3242 = ~n13488 | ~n13487;
  assign n13492 = ~n13490 | ~n13489;
  assign n13493 = ~n13492 ^ n13491;
  assign n13504 = ~n13493 | ~n16575;
  assign n13497 = ~n13494 | ~n13871;
  assign n13496 = ~n13495 | ~n13935;
  assign n13502 = ~n13497 | ~n13496;
  assign n13500 = ~n16569 | ~n14102;
  assign n13498 = ~n16624 | ~n13881;
  assign n16830 = ~P2_REG3_REG_15__SCAN_IN | ~P2_U3152;
  assign n13499 = n13498 & n16830;
  assign n13501 = ~n13500 | ~n13499;
  assign n13503 = ~n13502 & ~n13501;
  assign P2_U3243 = ~n13504 | ~n13503;
  assign n13522 = ~n13531 | ~n13505;
  assign n13507 = ~n13522 & ~n13506;
  assign n13944 = ~n13507 ^ n13945;
  assign n13513 = ~n13944;
  assign n13509 = ~n13508 & ~n13948;
  assign n13511 = ~n13510 | ~n13509;
  assign n13512 = ~n12487;
  assign n13521 = ~n13513 | ~n17186;
  assign n13519 = ~n13945 & ~n17068;
  assign n13946 = n13515 | n13514;
  assign n13954 = ~n13946;
  assign n13523 = ~n17087 | ~n13954;
  assign n13516 = ~P2_REG2_REG_31__SCAN_IN;
  assign n13517 = n17087 | n13516;
  assign n13518 = ~n13523 | ~n13517;
  assign n13520 = ~n13519 & ~n13518;
  assign P2_U3265 = ~n13521 | ~n13520;
  assign n13952 = ~n13953 ^ n13522;
  assign n13528 = ~n13952 | ~n17186;
  assign n13526 = ~n13953 & ~n17068;
  assign n13524 = ~n17218 | ~P2_REG2_REG_30__SCAN_IN;
  assign n13525 = ~n13524 | ~n13523;
  assign n13527 = ~n13526 & ~n13525;
  assign P2_U3266 = ~n13528 | ~n13527;
  assign n13536 = ~n13530 | ~n17186;
  assign n13534 = ~n13531 & ~n17068;
  assign n13533 = ~n17209 & ~n13532;
  assign n13535 = ~n13534 & ~n13533;
  assign n13568 = ~n13538 | ~n13537;
  assign n17213 = ~n17173 | ~n13568;
  assign n13677 = n17087 & n17213;
  assign n13540 = ~n13539 | ~n13677;
  assign n13542 = n13555 ^ n13541;
  assign n13544 = ~n13542 | ~n17212;
  assign n13968 = ~n13544 | ~n13543;
  assign n13545 = ~n17087 & ~P2_REG2_REG_28__SCAN_IN;
  assign n13553 = ~n13546 & ~n13545;
  assign n13963 = ~n13569 ^ n9749;
  assign n13552 = ~n13963 | ~n17186;
  assign n13550 = ~n9749 & ~n17068;
  assign n13548 = ~n13547;
  assign n13549 = ~n17209 & ~n13548;
  assign n13551 = ~n13550 & ~n13549;
  assign n13962 = ~n13554 ^ n13555;
  assign n13556 = ~n13962 | ~n13677;
  assign n13565 = ~n13972 & ~n17173;
  assign n13561 = ~n13559 ^ n13560;
  assign n13563 = ~n13561 | ~n17212;
  assign n13564 = ~n13563 | ~n13562;
  assign n13567 = ~n13980 | ~n17087;
  assign n13566 = n17087 | P2_REG2_REG_27__SCAN_IN;
  assign n13582 = ~n13567 | ~n13566;
  assign n17176 = ~n13568;
  assign n13580 = ~n13972 & ~n17130;
  assign n13571 = ~n13569;
  assign n13570 = ~n13572 & ~n9023;
  assign n13973 = ~n13571 & ~n13570;
  assign n13578 = ~n13973 | ~n17186;
  assign n13576 = ~n13572 & ~n17068;
  assign n13574 = ~n13573;
  assign n13575 = ~n17209 & ~n13574;
  assign n13577 = ~n13576 & ~n13575;
  assign n13579 = ~n13578 | ~n13577;
  assign n13581 = ~n13580 & ~n13579;
  assign P2_U3269 = ~n13582 | ~n13581;
  assign n13585 = ~n13583 | ~n13606;
  assign n13586 = ~n13585 | ~n13584;
  assign n13983 = ~n13586 ^ n13587;
  assign n13602 = ~n13983 | ~n17213;
  assign n13589 = ~n13588 ^ n13587;
  assign n13592 = ~n13589 | ~n17212;
  assign n13591 = ~n13590;
  assign n13988 = ~n13592 | ~n13591;
  assign n13594 = ~n13984 | ~n13593;
  assign n13595 = ~n13594 | ~n17502;
  assign n13597 = ~n13596 & ~n17209;
  assign n13598 = ~n17218 & ~n13597;
  assign n13600 = ~n13599 | ~n13598;
  assign n13601 = ~n13988 & ~n13600;
  assign n13603 = n17087 | P2_REG2_REG_26__SCAN_IN;
  assign n13604 = ~n13984 | ~n17206;
  assign P2_U3270 = ~n13605 | ~n13604;
  assign n13993 = ~n13606 ^ n13583;
  assign n13619 = ~n13993 | ~n17213;
  assign n13609 = ~n13607 & ~n13608;
  assign n13611 = ~n13609 & ~n17362;
  assign n13614 = ~n13611 | ~n13610;
  assign n13613 = ~n13612;
  assign n13999 = ~n13614 | ~n13613;
  assign n13994 = ~n13615 ^ n13995;
  assign n13616 = ~n13994 | ~n13512;
  assign n13617 = ~n13616 | ~n17087;
  assign n13618 = ~n13999 & ~n13617;
  assign n13621 = ~n13619 | ~n13618;
  assign n13620 = n17087 | P2_REG2_REG_25__SCAN_IN;
  assign n13628 = ~n13621 | ~n13620;
  assign n13626 = ~n13622 & ~n17068;
  assign n13624 = ~n13623;
  assign n13625 = ~n13624 & ~n17209;
  assign n13627 = ~n13626 & ~n13625;
  assign P2_U3271 = ~n13628 | ~n13627;
  assign n14004 = ~n13629 ^ n13631;
  assign n13640 = ~n14004 & ~n17173;
  assign n13632 = ~n13630 & ~n13631;
  assign n13633 = ~n13632 & ~n17362;
  assign n13638 = n13634 & n13633;
  assign n13636 = ~n17576 | ~n16628;
  assign n13635 = ~n17570 | ~n16626;
  assign n13637 = ~n13636 | ~n13635;
  assign n13642 = n14012 & n17087;
  assign n13641 = ~n17087 & ~P2_REG2_REG_24__SCAN_IN;
  assign n13653 = ~n13642 & ~n13641;
  assign n13651 = n14004 | n17130;
  assign n14005 = ~n13644 ^ n13643;
  assign n13649 = ~n14005 | ~n17186;
  assign n13647 = ~n14006 | ~n17206;
  assign n17190 = ~n17209;
  assign n13646 = ~n13645 | ~n17190;
  assign n13648 = n13647 & n13646;
  assign n13650 = n13649 & n13648;
  assign n13652 = ~n13651 | ~n13650;
  assign P2_U3272 = n13653 | n13652;
  assign n14015 = ~n9135 ^ n9947;
  assign n13662 = ~n14015 & ~n17173;
  assign n13660 = ~n13654 | ~n17212;
  assign n13658 = ~n13655 & ~n16604;
  assign n13657 = ~n13656 & ~n16605;
  assign n13659 = ~n13658 & ~n13657;
  assign n13661 = ~n13660 | ~n13659;
  assign n14023 = ~n13662 & ~n13661;
  assign n13664 = ~n14023 | ~n17087;
  assign n13663 = n17087 | P2_REG2_REG_23__SCAN_IN;
  assign n13676 = ~n13664 | ~n13663;
  assign n13674 = ~n14015 & ~n17130;
  assign n14016 = ~n13665 ^ n14017;
  assign n13672 = ~n14016 | ~n17186;
  assign n13670 = ~n13666 & ~n17068;
  assign n13668 = ~n13667;
  assign n13669 = ~n13668 & ~n17209;
  assign n13671 = ~n13670 & ~n13669;
  assign n13673 = ~n13672 | ~n13671;
  assign n13675 = ~n13674 & ~n13673;
  assign P2_U3273 = ~n13676 | ~n13675;
  assign n14026 = ~n9116 ^ n13680;
  assign n13700 = ~n14026 | ~n13677;
  assign n13683 = ~n13678;
  assign n13681 = ~n13679 | ~n13680;
  assign n13682 = ~n13681 | ~n17212;
  assign n13687 = ~n13683 & ~n13682;
  assign n13685 = ~n17570 | ~n16628;
  assign n13684 = ~n16626 | ~n17564;
  assign n13686 = ~n13685 | ~n13684;
  assign n14031 = n13687 | n13686;
  assign n13689 = ~n14031 & ~n17218;
  assign n13688 = ~n17087 & ~P2_REG2_REG_22__SCAN_IN;
  assign n13698 = ~n13689 & ~n13688;
  assign n14027 = ~n9143 ^ n11008;
  assign n13696 = ~n14027 | ~n17186;
  assign n13694 = ~n13690 & ~n17068;
  assign n13692 = ~n13691;
  assign n13693 = ~n13692 & ~n17209;
  assign n13695 = ~n13694 & ~n13693;
  assign n13697 = ~n13696 | ~n13695;
  assign n13699 = ~n13698 & ~n13697;
  assign P2_U3274 = ~n13700 | ~n13699;
  assign n14036 = ~n13701 ^ n13703;
  assign n13710 = ~n14036 & ~n17173;
  assign n13704 = n13702 ^ n13703;
  assign n13708 = ~n13704 & ~n17362;
  assign n13706 = ~n17567 | ~n16628;
  assign n13705 = ~n16626 | ~n17561;
  assign n13707 = ~n13706 | ~n13705;
  assign n13709 = n13708 | n13707;
  assign n14044 = ~n13710 & ~n13709;
  assign n13712 = ~n14044 | ~n17087;
  assign n13711 = n17087 | P2_REG2_REG_21__SCAN_IN;
  assign n13724 = ~n13712 | ~n13711;
  assign n13722 = ~n14036 & ~n17130;
  assign n14037 = ~n13713 ^ n14038;
  assign n13720 = ~n14037 | ~n17186;
  assign n13718 = ~n13714 & ~n17068;
  assign n13716 = ~n13715;
  assign n13717 = ~n17209 & ~n13716;
  assign n13719 = ~n13718 & ~n13717;
  assign n13721 = ~n13720 | ~n13719;
  assign n13723 = ~n13722 & ~n13721;
  assign P2_U3275 = ~n13724 | ~n13723;
  assign n14047 = ~n13725 ^ n13727;
  assign n13735 = ~n14047 & ~n17173;
  assign n13728 = ~n13726 ^ n13727;
  assign n13733 = ~n13728 | ~n17212;
  assign n13731 = ~n16604 & ~n13729;
  assign n13730 = ~n13777 & ~n16605;
  assign n13732 = ~n13731 & ~n13730;
  assign n13734 = ~n13733 | ~n13732;
  assign n14055 = ~n13735 & ~n13734;
  assign n13737 = ~n14055 | ~n17087;
  assign n13736 = n17087 | P2_REG2_REG_20__SCAN_IN;
  assign n13747 = ~n13737 | ~n13736;
  assign n13745 = ~n14047 & ~n17130;
  assign n14048 = n14049 ^ n9100;
  assign n13743 = ~n14048 | ~n17186;
  assign n13741 = ~n9765 & ~n17068;
  assign n13739 = ~n13738;
  assign n13740 = ~n17209 & ~n13739;
  assign n13742 = ~n13741 & ~n13740;
  assign n13744 = ~n13743 | ~n13742;
  assign n13746 = ~n13745 & ~n13744;
  assign P2_U3276 = ~n13747 | ~n13746;
  assign n14058 = ~n13748 ^ n13750;
  assign n13762 = ~n14058 | ~n17150;
  assign n13751 = n13749 ^ n13750;
  assign n13756 = ~n13751 | ~n17212;
  assign n13754 = ~n16604 & ~n13752;
  assign n13753 = ~n16605 & ~n13805;
  assign n13755 = ~n13754 & ~n13753;
  assign n14064 = ~n13756 | ~n13755;
  assign n13758 = ~n13757 | ~n14060;
  assign n14059 = n9100 & n13758;
  assign n13759 = ~n14059 | ~n13512;
  assign n13760 = ~n13759 | ~n17087;
  assign n13761 = ~n14064 & ~n13760;
  assign n13765 = ~n13762 | ~n13761;
  assign n13763 = ~P2_REG2_REG_19__SCAN_IN;
  assign n13764 = ~n17218 | ~n13763;
  assign n13772 = ~n13765 | ~n13764;
  assign n17144 = ~n17130;
  assign n13770 = ~n14058 | ~n17144;
  assign n13768 = ~n14060 | ~n17206;
  assign n13767 = n17209 | n13766;
  assign n13769 = n13768 & n13767;
  assign n13771 = n13770 & n13769;
  assign P2_U3277 = ~n13772 | ~n13771;
  assign n14069 = n13773 ^ n13775;
  assign n13784 = ~n14069 & ~n17173;
  assign n13776 = n13774 ^ n13775;
  assign n13782 = ~n13776 | ~n17212;
  assign n13780 = ~n16604 & ~n13777;
  assign n13779 = ~n16605 & ~n13778;
  assign n13781 = ~n13780 & ~n13779;
  assign n13783 = ~n13782 | ~n13781;
  assign n14077 = ~n13784 & ~n13783;
  assign n13786 = ~n14077 | ~n17087;
  assign n16896 = ~P2_REG2_REG_18__SCAN_IN;
  assign n13785 = ~n17218 | ~n16896;
  assign n13798 = ~n13786 | ~n13785;
  assign n13796 = ~n14069 & ~n17130;
  assign n14070 = ~n13787 ^ n14071;
  assign n13794 = ~n14070 | ~n17186;
  assign n13792 = ~n13788 & ~n17068;
  assign n13790 = ~n13789;
  assign n13791 = ~n17209 & ~n13790;
  assign n13793 = ~n13792 & ~n13791;
  assign n13795 = ~n13794 | ~n13793;
  assign n13797 = ~n13796 & ~n13795;
  assign P2_U3278 = ~n13798 | ~n13797;
  assign n14080 = n13799 ^ n13801;
  assign n13812 = ~n14080 & ~n17173;
  assign n13802 = ~n13800 & ~n13801;
  assign n13804 = ~n13802 & ~n17362;
  assign n13810 = ~n13804 | ~n13803;
  assign n13808 = ~n16604 & ~n13805;
  assign n13807 = ~n16605 & ~n13806;
  assign n13809 = ~n13808 & ~n13807;
  assign n13811 = ~n13810 | ~n13809;
  assign n14087 = ~n13812 & ~n13811;
  assign n14081 = ~n13847 ^ n13813;
  assign n13814 = ~n14081 | ~n13512;
  assign n13815 = n13814 & n17087;
  assign n13817 = ~n14087 | ~n13815;
  assign n16877 = ~P2_REG2_REG_17__SCAN_IN;
  assign n13816 = ~n17218 | ~n16877;
  assign n13824 = ~n13817 | ~n13816;
  assign n13822 = ~n14080 & ~n17130;
  assign n13820 = ~n13279 | ~n17206;
  assign n13819 = ~n17190 | ~n13818;
  assign n13821 = ~n13820 | ~n13819;
  assign n13823 = ~n13822 & ~n13821;
  assign P2_U3279 = ~n13824 | ~n13823;
  assign n13863 = ~n13825 | ~n13826;
  assign n13828 = ~n13863 | ~n13832;
  assign n13829 = n13828 & n13827;
  assign n13855 = ~n13829 ^ n9512;
  assign n13844 = ~n13855 | ~n17150;
  assign n13831 = ~n13830;
  assign n13867 = ~n13895 | ~n13831;
  assign n13866 = ~n13832;
  assign n13865 = ~n13867 | ~n13866;
  assign n13834 = ~n13865 | ~n13833;
  assign n13836 = n13835 ^ n13834;
  assign n13842 = ~n13836 & ~n17362;
  assign n13840 = ~n16626 | ~n13837;
  assign n13839 = ~n16628 | ~n13838;
  assign n13841 = ~n13840 | ~n13839;
  assign n13843 = ~n13842 & ~n13841;
  assign n14096 = ~n13844 | ~n13843;
  assign n13851 = ~n14096;
  assign n13846 = ~n13845 | ~n14091;
  assign n13848 = n13846 & n17502;
  assign n14093 = ~n13848 | ~n13847;
  assign n13849 = ~n14093 & ~n17098;
  assign n13850 = ~n13849 & ~n17218;
  assign n13854 = ~n13851 | ~n13850;
  assign n13852 = ~P2_REG2_REG_16__SCAN_IN;
  assign n13853 = ~n17218 | ~n13852;
  assign n13862 = ~n13854 | ~n13853;
  assign n14090 = ~n13855;
  assign n13860 = ~n14090 & ~n17130;
  assign n13858 = ~n17206 | ~n14091;
  assign n13857 = ~n17190 | ~n13856;
  assign n13859 = ~n13858 | ~n13857;
  assign n13861 = ~n13860 & ~n13859;
  assign P2_U3280 = ~n13862 | ~n13861;
  assign n14100 = ~n13863 ^ n13866;
  assign n13864 = ~n14100;
  assign n13877 = ~n13864 | ~n17150;
  assign n13870 = ~n13865;
  assign n13868 = n13867 | n13866;
  assign n13869 = ~n13868 | ~n17212;
  assign n13875 = ~n13870 & ~n13869;
  assign n13873 = ~n16626 | ~n13935;
  assign n13872 = ~n16628 | ~n13871;
  assign n13874 = ~n13873 | ~n13872;
  assign n13876 = ~n13875 & ~n13874;
  assign n13880 = ~n14107 | ~n17087;
  assign n13878 = ~P2_REG2_REG_15__SCAN_IN;
  assign n13879 = ~n17218 | ~n13878;
  assign n13890 = ~n13880 | ~n13879;
  assign n13888 = ~n14100 & ~n17130;
  assign n14101 = n14102 ^ n9159;
  assign n13886 = ~n14101 | ~n17186;
  assign n13884 = ~n17068 & ~n9214;
  assign n13882 = ~n13881;
  assign n13883 = ~n17209 & ~n13882;
  assign n13885 = ~n13884 & ~n13883;
  assign n13887 = ~n13886 | ~n13885;
  assign n13889 = ~n13888 & ~n13887;
  assign P2_U3281 = ~n13890 | ~n13889;
  assign n14111 = ~n13891 ^ n9952;
  assign n13904 = ~n14111 & ~n17173;
  assign n13894 = ~n13892 | ~n13893;
  assign n13896 = n13894 & n17212;
  assign n13902 = ~n13896 | ~n13895;
  assign n13900 = ~n16604 & ~n13897;
  assign n13899 = ~n16605 & ~n13898;
  assign n13901 = ~n13900 & ~n13899;
  assign n13903 = ~n13902 | ~n13901;
  assign n14120 = ~n13904 & ~n13903;
  assign n13907 = ~n14120 | ~n17087;
  assign n13905 = ~P2_REG2_REG_14__SCAN_IN;
  assign n13906 = ~n17218 | ~n13905;
  assign n13919 = ~n13907 | ~n13906;
  assign n13917 = ~n14111 & ~n17130;
  assign n14112 = ~n13908 ^ n14114;
  assign n13915 = ~n14112 | ~n17186;
  assign n13913 = ~n17068 & ~n13909;
  assign n13911 = ~n13910;
  assign n13912 = ~n17209 & ~n13911;
  assign n13914 = ~n13913 & ~n13912;
  assign n13916 = ~n13915 | ~n13914;
  assign n13918 = ~n13917 & ~n13916;
  assign P2_U3282 = ~n13919 | ~n13918;
  assign n13922 = ~n17206 | ~n13920;
  assign n13921 = ~n17218 | ~P2_REG2_REG_13__SCAN_IN;
  assign n13925 = n13922 & n13921;
  assign n13924 = ~n13923 | ~n17190;
  assign n13931 = ~n13925 | ~n13924;
  assign n14123 = ~n9042 ^ n9577;
  assign n13929 = ~n14123 | ~n17144;
  assign n14124 = ~n13926 ^ n14125;
  assign n13927 = ~n14124;
  assign n13928 = ~n13927 | ~n17186;
  assign n13930 = ~n13929 | ~n13928;
  assign n13943 = ~n13931 & ~n13930;
  assign n13941 = ~n14123 | ~n17150;
  assign n13934 = ~n13932 ^ n13933;
  assign n13939 = ~n13934 & ~n17362;
  assign n13937 = ~n16626 | ~n16592;
  assign n13936 = ~n16628 | ~n13935;
  assign n13938 = ~n13937 | ~n13936;
  assign n13940 = ~n13939 & ~n13938;
  assign n14131 = ~n13941 | ~n13940;
  assign n13942 = ~n14131 | ~n17087;
  assign P2_U3283 = ~n13943 | ~n13942;
  assign n13947 = n13945 | n17487;
  assign n13950 = ~n17553 | ~P2_REG1_REG_31__SCAN_IN;
  assign P2_U3551 = ~n13951 | ~n13950;
  assign n13957 = ~n13952 | ~n17502;
  assign n13955 = ~n13953 & ~n17487;
  assign n13956 = ~n13955 & ~n13954;
  assign n14136 = ~n13957 | ~n13956;
  assign n13959 = ~n14136 | ~n17555;
  assign n13958 = ~n17553 | ~P2_REG1_REG_30__SCAN_IN;
  assign P2_U3550 = ~n13959 | ~n13958;
  assign n13960 = ~n17553 | ~P2_REG1_REG_29__SCAN_IN;
  assign P2_U3549 = ~n13961 | ~n13960;
  assign n13966 = ~n13963 | ~n17502;
  assign n13965 = ~n13964 | ~n17504;
  assign n13967 = ~n13966 | ~n13965;
  assign n13969 = ~n13968 & ~n13967;
  assign n13971 = ~n14139 | ~n17555;
  assign n13970 = ~n17553 | ~P2_REG1_REG_28__SCAN_IN;
  assign P2_U3548 = ~n13971 | ~n13970;
  assign n13978 = ~n13972 & ~n17493;
  assign n13976 = ~n13973 | ~n17502;
  assign n13975 = ~n13974 | ~n17504;
  assign n13977 = ~n13976 | ~n13975;
  assign n13979 = ~n13978 & ~n13977;
  assign n14142 = ~n13980 | ~n13979;
  assign n13982 = ~n14142 | ~n17555;
  assign n13981 = ~n17553 | ~P2_REG1_REG_27__SCAN_IN;
  assign P2_U3547 = ~n13982 | ~n13981;
  assign n13990 = ~n13983 | ~n17446;
  assign n13985 = ~n13984 | ~n14113;
  assign n13987 = ~n13986 | ~n13985;
  assign n13989 = ~n13988 & ~n13987;
  assign n14145 = ~n13990 | ~n13989;
  assign n13992 = ~n14145 | ~n17555;
  assign n13991 = ~n17553 | ~P2_REG1_REG_26__SCAN_IN;
  assign P2_U3546 = ~n13992 | ~n13991;
  assign n14001 = ~n13993 | ~n17446;
  assign n13997 = ~n13994 | ~n17502;
  assign n13996 = ~n13995 | ~n17504;
  assign n13998 = ~n13997 | ~n13996;
  assign n14000 = ~n13999 & ~n13998;
  assign n14148 = ~n14001 | ~n14000;
  assign n14003 = ~n14148 | ~n17555;
  assign n14002 = ~n17553 | ~P2_REG1_REG_25__SCAN_IN;
  assign P2_U3545 = ~n14003 | ~n14002;
  assign n14010 = ~n14004 & ~n17493;
  assign n14008 = ~n14005 | ~n17502;
  assign n14007 = ~n14006 | ~n17504;
  assign n14009 = ~n14008 | ~n14007;
  assign n14011 = ~n14010 & ~n14009;
  assign n14151 = ~n14012 | ~n14011;
  assign n14014 = ~n14151 | ~n17555;
  assign n14013 = ~n17553 | ~P2_REG1_REG_24__SCAN_IN;
  assign P2_U3544 = ~n14014 | ~n14013;
  assign n14021 = ~n14015 & ~n17493;
  assign n14019 = ~n14016 | ~n17502;
  assign n14018 = ~n14017 | ~n14113;
  assign n14020 = ~n14019 | ~n14018;
  assign n14022 = ~n14021 & ~n14020;
  assign n14154 = ~n14023 | ~n14022;
  assign n14025 = ~n14154 | ~n17555;
  assign n14024 = ~n17553 | ~P2_REG1_REG_23__SCAN_IN;
  assign P2_U3543 = ~n14025 | ~n14024;
  assign n14033 = ~n14026 | ~n17446;
  assign n14029 = ~n14027 | ~n17502;
  assign n14028 = ~n11008 | ~n17504;
  assign n14030 = ~n14029 | ~n14028;
  assign n14032 = ~n14031 & ~n14030;
  assign n14157 = ~n14033 | ~n14032;
  assign n14035 = ~n14157 | ~n17555;
  assign n14034 = ~n17553 | ~P2_REG1_REG_22__SCAN_IN;
  assign P2_U3542 = ~n14035 | ~n14034;
  assign n14042 = ~n14036 & ~n17493;
  assign n14040 = ~n14037 | ~n17502;
  assign n14039 = ~n14038 | ~n17504;
  assign n14041 = ~n14040 | ~n14039;
  assign n14043 = ~n14042 & ~n14041;
  assign n14160 = ~n14044 | ~n14043;
  assign n14046 = ~n14160 | ~n17555;
  assign n14045 = ~n17553 | ~P2_REG1_REG_21__SCAN_IN;
  assign P2_U3541 = ~n14046 | ~n14045;
  assign n14053 = ~n14047 & ~n17493;
  assign n14051 = ~n14048 | ~n17502;
  assign n14050 = ~n14049 | ~n14113;
  assign n14052 = ~n14051 | ~n14050;
  assign n14054 = ~n14053 & ~n14052;
  assign n14163 = ~n14055 | ~n14054;
  assign n14057 = ~n14163 | ~n17555;
  assign n14056 = ~n17553 | ~P2_REG1_REG_20__SCAN_IN;
  assign P2_U3540 = ~n14057 | ~n14056;
  assign n14066 = ~n14058 | ~n17446;
  assign n14062 = ~n14059 | ~n17502;
  assign n14061 = ~n14060 | ~n17504;
  assign n14063 = ~n14062 | ~n14061;
  assign n14065 = ~n14064 & ~n14063;
  assign n14166 = ~n14066 | ~n14065;
  assign n14068 = ~n14166 | ~n17555;
  assign n14067 = ~n17553 | ~P2_REG1_REG_19__SCAN_IN;
  assign P2_U3539 = ~n14068 | ~n14067;
  assign n14075 = ~n14069 & ~n17493;
  assign n14073 = ~n14070 | ~n17502;
  assign n14072 = ~n14071 | ~n17504;
  assign n14074 = ~n14073 | ~n14072;
  assign n14076 = ~n14075 & ~n14074;
  assign n14169 = ~n14077 | ~n14076;
  assign n14079 = ~n14169 | ~n17555;
  assign n14078 = ~n17553 | ~P2_REG1_REG_18__SCAN_IN;
  assign P2_U3538 = ~n14079 | ~n14078;
  assign n14085 = ~n14080 & ~n17493;
  assign n14083 = ~n14081 | ~n17502;
  assign n14082 = ~n13279 | ~n17504;
  assign n14084 = ~n14083 | ~n14082;
  assign n14086 = ~n14085 & ~n14084;
  assign n14172 = ~n14087 | ~n14086;
  assign n14089 = ~n14172 | ~n17555;
  assign n14088 = ~n17553 | ~P2_REG1_REG_17__SCAN_IN;
  assign P2_U3537 = ~n14089 | ~n14088;
  assign n14095 = n14090 | n17493;
  assign n14092 = ~n14091 | ~n14113;
  assign n14094 = n14093 & n14092;
  assign n14097 = ~n14095 | ~n14094;
  assign n14099 = ~n14175 | ~n17555;
  assign n14098 = ~n17553 | ~P2_REG1_REG_16__SCAN_IN;
  assign P2_U3536 = ~n14099 | ~n14098;
  assign n14106 = ~n14100 & ~n17493;
  assign n14104 = ~n14101 | ~n17502;
  assign n14103 = ~n14102 | ~n17504;
  assign n14105 = ~n14104 | ~n14103;
  assign n14108 = ~n14106 & ~n14105;
  assign n14178 = ~n14108 | ~n14107;
  assign n14110 = ~n14178 | ~n17555;
  assign n14109 = ~n17553 | ~P2_REG1_REG_15__SCAN_IN;
  assign P2_U3535 = ~n14110 | ~n14109;
  assign n14118 = ~n14111 & ~n17493;
  assign n14116 = ~n14112 | ~n17502;
  assign n14115 = ~n14114 | ~n14113;
  assign n14117 = ~n14116 | ~n14115;
  assign n14119 = ~n14118 & ~n14117;
  assign n14181 = ~n14120 | ~n14119;
  assign n14122 = ~n14181 | ~n17555;
  assign n14121 = ~n17553 | ~P2_REG1_REG_14__SCAN_IN;
  assign P2_U3534 = ~n14122 | ~n14121;
  assign n17481 = ~n17493;
  assign n14129 = ~n14123 | ~n17481;
  assign n14127 = ~n14124 & ~n12581;
  assign n14126 = ~n14125 & ~n17487;
  assign n14128 = ~n14127 & ~n14126;
  assign n14130 = ~n14129 | ~n14128;
  assign n14133 = ~n14184 | ~n17555;
  assign n14132 = ~n17553 | ~P2_REG1_REG_13__SCAN_IN;
  assign P2_U3533 = ~n14133 | ~n14132;
  assign n14134 = ~n17501 | ~P2_REG0_REG_31__SCAN_IN;
  assign P2_U3519 = ~n14135 | ~n14134;
  assign n14138 = ~n14136 | ~n17514;
  assign n14137 = ~n17501 | ~P2_REG0_REG_30__SCAN_IN;
  assign P2_U3518 = ~n14138 | ~n14137;
  assign n14140 = ~n17501 | ~P2_REG0_REG_28__SCAN_IN;
  assign P2_U3516 = ~n14141 | ~n14140;
  assign n14144 = ~n14142 | ~n17514;
  assign n14143 = ~n17501 | ~P2_REG0_REG_27__SCAN_IN;
  assign P2_U3515 = ~n14144 | ~n14143;
  assign n14147 = ~n14145 | ~n17514;
  assign n14146 = ~n17501 | ~P2_REG0_REG_26__SCAN_IN;
  assign P2_U3514 = ~n14147 | ~n14146;
  assign n14150 = ~n14148 | ~n17514;
  assign n14149 = ~n17501 | ~P2_REG0_REG_25__SCAN_IN;
  assign P2_U3513 = ~n14150 | ~n14149;
  assign n14153 = ~n14151 | ~n17514;
  assign n14152 = ~n17501 | ~P2_REG0_REG_24__SCAN_IN;
  assign P2_U3512 = ~n14153 | ~n14152;
  assign n14156 = ~n14154 | ~n17514;
  assign n14155 = ~n17501 | ~P2_REG0_REG_23__SCAN_IN;
  assign P2_U3511 = ~n14156 | ~n14155;
  assign n14159 = ~n14157 | ~n17514;
  assign n14158 = ~n17501 | ~P2_REG0_REG_22__SCAN_IN;
  assign P2_U3510 = ~n14159 | ~n14158;
  assign n14162 = ~n14160 | ~n17514;
  assign n14161 = ~n17501 | ~P2_REG0_REG_21__SCAN_IN;
  assign P2_U3509 = ~n14162 | ~n14161;
  assign n14165 = ~n14163 | ~n17514;
  assign n14164 = ~n17501 | ~P2_REG0_REG_20__SCAN_IN;
  assign P2_U3508 = ~n14165 | ~n14164;
  assign n14168 = ~n14166 | ~n17514;
  assign n14167 = ~n17501 | ~P2_REG0_REG_19__SCAN_IN;
  assign P2_U3507 = ~n14168 | ~n14167;
  assign n14171 = ~n14169 | ~n17514;
  assign n14170 = ~n17501 | ~P2_REG0_REG_18__SCAN_IN;
  assign P2_U3505 = ~n14171 | ~n14170;
  assign n14174 = ~n14172 | ~n17514;
  assign n14173 = ~n17501 | ~P2_REG0_REG_17__SCAN_IN;
  assign P2_U3502 = ~n14174 | ~n14173;
  assign n14177 = ~n14175 | ~n17514;
  assign n14176 = ~n17501 | ~P2_REG0_REG_16__SCAN_IN;
  assign P2_U3499 = ~n14177 | ~n14176;
  assign n14180 = ~n14178 | ~n17514;
  assign n14179 = ~n17501 | ~P2_REG0_REG_15__SCAN_IN;
  assign P2_U3496 = ~n14180 | ~n14179;
  assign n14183 = ~n14181 | ~n17514;
  assign n14182 = ~n17501 | ~P2_REG0_REG_14__SCAN_IN;
  assign P2_U3493 = ~n14183 | ~n14182;
  assign n14186 = ~n14184 | ~n17514;
  assign n14185 = ~n17501 | ~P2_REG0_REG_13__SCAN_IN;
  assign P2_U3490 = ~n14186 | ~n14185;
  assign n14194 = ~n15275 | ~n14227;
  assign n14188 = ~n10523 & ~P2_IR_REG_30__SCAN_IN;
  assign n14189 = ~n14188 | ~P2_STATE_REG_SCAN_IN;
  assign n14192 = ~n14187 & ~n14189;
  assign n14190 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n14191 = ~n14229 & ~n14190;
  assign n14193 = ~n14192 & ~n14191;
  assign P2_U3327 = ~n14194 | ~n14193;
  assign n15285 = ~n14195;
  assign n14201 = ~n15285 | ~n14227;
  assign n14199 = ~n14196 & ~P2_U3152;
  assign n14198 = ~n14229 & ~n14197;
  assign n14200 = ~n14199 & ~n14198;
  assign P2_U3328 = ~n14201 | ~n14200;
  assign n15292 = ~n14202;
  assign n14207 = ~n15292 | ~n14227;
  assign n14205 = ~n9996 & ~P2_U3152;
  assign n14204 = ~n14229 & ~n14203;
  assign n14206 = ~n14205 & ~n14204;
  assign P2_U3329 = ~n14207 | ~n14206;
  assign n15298 = ~n14208;
  assign n14212 = ~n15298 & ~n17340;
  assign n14209 = ~n17347 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n14211 = ~n14210 | ~n14209;
  assign P2_U3330 = n14212 | n14211;
  assign n15304 = ~n14213;
  assign n14219 = ~n15304 | ~n14227;
  assign n14217 = ~n14214 & ~P2_U3152;
  assign n14216 = ~n14229 & ~n14215;
  assign n14218 = ~n14217 & ~n14216;
  assign P2_U3331 = ~n14219 | ~n14218;
  assign n14225 = ~n15309 | ~n14227;
  assign n14223 = ~n14220 & ~P2_U3152;
  assign n14222 = ~n14229 & ~n14221;
  assign n14224 = ~n14223 & ~n14222;
  assign P2_U3332 = ~n14225 | ~n14224;
  assign n15318 = ~n14226;
  assign n14234 = ~n15318 | ~n14227;
  assign n14232 = ~n14229 & ~n14228;
  assign n14230 = ~n17352;
  assign n14231 = ~P2_U3152 & ~n14230;
  assign n14233 = ~n14232 & ~n14231;
  assign P2_U3334 = ~n14234 | ~n14233;
  assign n14236 = ~n14235;
  assign n14238 = ~n14237 & ~n14236;
  assign n14240 = ~n14239 ^ n14238;
  assign n14250 = ~n14240 | ~n15457;
  assign n14248 = ~n15035 | ~n15421;
  assign n14246 = ~n14586 & ~n15441;
  assign n14244 = ~n15402 | ~n14597;
  assign n14242 = ~n15419 | ~n16416;
  assign n14241 = ~P1_REG3_REG_27__SCAN_IN | ~P1_U3084;
  assign n14243 = n14242 & n14241;
  assign n14245 = ~n14244 | ~n14243;
  assign n14247 = ~n14246 & ~n14245;
  assign n14249 = n14248 & n14247;
  assign P1_U3212 = ~n14250 | ~n14249;
  assign n14253 = ~n14252 ^ n14251;
  assign n14255 = ~n14254 ^ n14253;
  assign n14264 = ~n14255 | ~n15457;
  assign n14262 = ~n14919 & ~n15442;
  assign n14260 = ~n15402 | ~n14924;
  assign n14256 = ~n15429 | ~n14907;
  assign n15722 = ~P1_REG3_REG_14__SCAN_IN | ~P1_U3084;
  assign n14258 = ~n14256 | ~n15722;
  assign n14257 = ~n15438 & ~n14364;
  assign n14259 = ~n14258 & ~n14257;
  assign n14261 = ~n14260 | ~n14259;
  assign n14263 = ~n14262 & ~n14261;
  assign P1_U3213 = ~n14264 | ~n14263;
  assign n14268 = n14266 | n14265;
  assign n14392 = ~n14268 | ~n14269;
  assign n14267 = ~n14392;
  assign n14391 = ~n14266 | ~n14265;
  assign n14273 = ~n14267 | ~n14391;
  assign n14271 = ~n14268 | ~n14391;
  assign n14270 = ~n14269;
  assign n14272 = ~n14271 | ~n14270;
  assign n14274 = ~n14273 | ~n14272;
  assign n14285 = ~n14274 | ~n15457;
  assign n14691 = ~n15080;
  assign n14283 = ~n14691 & ~n15442;
  assign n14275 = ~n14692;
  assign n14281 = ~n15402 | ~n14275;
  assign n14279 = ~n16398 | ~n15429;
  assign n14277 = ~n15419 | ~n16404;
  assign n14276 = ~P1_REG3_REG_23__SCAN_IN | ~P1_U3084;
  assign n14278 = n14277 & n14276;
  assign n14280 = n14279 & n14278;
  assign n14282 = ~n14281 | ~n14280;
  assign n14284 = ~n14283 & ~n14282;
  assign P1_U3214 = ~n14285 | ~n14284;
  assign n14286 = ~n14289;
  assign n14486 = ~n14286 | ~n14287;
  assign n14288 = ~n14287;
  assign n14484 = ~n14289 | ~n14288;
  assign n14290 = ~n14486 | ~n14484;
  assign n14291 = n14483 ^ n14290;
  assign n14302 = ~n14291 & ~n15414;
  assign n14300 = ~n15402 | ~n14292;
  assign n14293 = ~n15429 | ~n15881;
  assign n15646 = ~P1_REG3_REG_10__SCAN_IN | ~P1_U3084;
  assign n14295 = ~n14293 | ~n15646;
  assign n14294 = ~n15438 & ~n14964;
  assign n14298 = ~n14295 & ~n14294;
  assign n14297 = ~n14296 | ~n15421;
  assign n14299 = n14298 & n14297;
  assign n14301 = ~n14300 | ~n14299;
  assign P1_U3215 = n14302 | n14301;
  assign n14305 = ~n14303;
  assign n14304 = ~n14504;
  assign n14502 = ~n14306 | ~n14305;
  assign n14319 = n14500 & n14502;
  assign n14307 = ~n14318 | ~n14320;
  assign n14308 = ~n14319 ^ n14307;
  assign n14317 = ~n14308 | ~n15457;
  assign n14315 = ~n9684 & ~n15442;
  assign n14313 = ~n15402 | ~n14780;
  assign n14309 = ~n15419 | ~n14774;
  assign n15808 = ~P1_REG3_REG_19__SCAN_IN | ~P1_U3084;
  assign n14311 = ~n14309 | ~n15808;
  assign n14310 = n15429 & n14775;
  assign n14312 = ~n14311 & ~n14310;
  assign n14314 = ~n14313 | ~n14312;
  assign n14316 = ~n14315 & ~n14314;
  assign P1_U3217 = ~n14317 | ~n14316;
  assign n14321 = ~n14319 | ~n14318;
  assign n14430 = ~n14321 | ~n14320;
  assign n14429 = ~n14323 | ~n14322;
  assign n14325 = ~n14430 & ~n14429;
  assign n14324 = ~n14323;
  assign n14328 = ~n14327 | ~n14326;
  assign n14330 = ~n14329 ^ n14328;
  assign n14342 = ~n14330 | ~n15457;
  assign n14340 = ~n14737 & ~n15442;
  assign n14335 = ~n14331 & ~n15438;
  assign n14333 = ~n15429 | ~n14774;
  assign n14332 = ~P1_REG3_REG_21__SCAN_IN | ~P1_U3084;
  assign n14334 = ~n14333 | ~n14332;
  assign n14338 = ~n14335 & ~n14334;
  assign n14336 = ~n14738;
  assign n14337 = ~n15402 | ~n14336;
  assign n14339 = ~n14338 | ~n14337;
  assign n14341 = ~n14340 & ~n14339;
  assign P1_U3221 = ~n14342 | ~n14341;
  assign n14346 = ~n14344 | ~n14343;
  assign n14347 = n14346 ^ n14345;
  assign n14357 = ~n14347 | ~n15457;
  assign n14644 = ~n15059;
  assign n14355 = ~n14644 & ~n15442;
  assign n14351 = ~n15447 & ~n14645;
  assign n14349 = ~n15429 | ~n16404;
  assign n14348 = ~P1_REG3_REG_25__SCAN_IN | ~P1_U3084;
  assign n14350 = ~n14349 | ~n14348;
  assign n14353 = ~n14351 & ~n14350;
  assign n14352 = ~n16410 | ~n15419;
  assign n14354 = ~n14353 | ~n14352;
  assign n14356 = ~n14355 & ~n14354;
  assign P1_U3223 = ~n14357 | ~n14356;
  assign n14360 = ~n14359 | ~n14358;
  assign n14362 = ~n14361 ^ n14360;
  assign n14373 = ~n14362 | ~n15457;
  assign n14371 = ~n14363 & ~n15442;
  assign n14369 = ~n15402 | ~n14872;
  assign n14367 = ~n15441 & ~n14364;
  assign n14365 = ~n15419 | ~n14859;
  assign n15755 = ~P1_REG3_REG_16__SCAN_IN | ~P1_U3084;
  assign n14366 = ~n14365 | ~n15755;
  assign n14368 = ~n14367 & ~n14366;
  assign n14370 = ~n14369 | ~n14368;
  assign n14372 = ~n14371 & ~n14370;
  assign P1_U3224 = ~n14373 | ~n14372;
  assign n14380 = ~n9074 | ~n14375;
  assign n14376 = ~n14374;
  assign n14377 = ~n14376 | ~n14375;
  assign n14379 = ~n14378 | ~n14377;
  assign n14381 = ~n14380 | ~n14379;
  assign n14390 = ~n14381 | ~n15457;
  assign n14388 = ~n14843 & ~n15442;
  assign n14386 = ~n15402 | ~n14844;
  assign n14382 = ~n15429 | ~n14533;
  assign n15774 = ~P1_REG3_REG_17__SCAN_IN | ~P1_U3084;
  assign n14384 = ~n14382 | ~n15774;
  assign n14383 = ~n15438 & ~n14828;
  assign n14385 = ~n14384 & ~n14383;
  assign n14387 = ~n14386 | ~n14385;
  assign n14389 = ~n14388 & ~n14387;
  assign P1_U3226 = ~n14390 | ~n14389;
  assign n14396 = ~n14392 | ~n14391;
  assign n14395 = ~n14394 & ~n14393;
  assign n14397 = ~n14396 ^ n14395;
  assign n14409 = ~n14397 | ~n15457;
  assign n14407 = ~n15069 | ~n15421;
  assign n14405 = ~n14608 & ~n15438;
  assign n14398 = ~n14669;
  assign n14401 = ~n15447 & ~n14398;
  assign n14400 = ~P1_STATE_REG_SCAN_IN & ~n14399;
  assign n14403 = ~n14401 & ~n14400;
  assign n14402 = ~n16401 | ~n15429;
  assign n14404 = ~n14403 | ~n14402;
  assign n14406 = ~n14405 & ~n14404;
  assign n14408 = n14407 & n14406;
  assign P1_U3227 = ~n14409 | ~n14408;
  assign n14413 = n14411 & n14410;
  assign n14412 = ~n14411 & ~n14410;
  assign n15364 = ~n14413 & ~n14412;
  assign n14415 = ~n15364 | ~n15365;
  assign n14414 = ~n14413;
  assign n14416 = ~n14415 | ~n14414;
  assign n14418 = n14417 ^ n14416;
  assign n14428 = ~n14418 & ~n15414;
  assign n14426 = ~n15402 | ~n14419;
  assign n14420 = ~n15429 | ~n15903;
  assign n15635 = ~P1_REG3_REG_9__SCAN_IN | ~P1_U3084;
  assign n14422 = ~n14420 | ~n15635;
  assign n14421 = ~n15438 & ~n15847;
  assign n14424 = ~n14422 & ~n14421;
  assign n14423 = ~n15421 | ~n16353;
  assign n14425 = n14424 & n14423;
  assign n14427 = ~n14426 | ~n14425;
  assign P1_U3229 = n14428 | n14427;
  assign n14431 = ~n14430 ^ n14429;
  assign n14443 = ~n14431 | ~n15457;
  assign n14441 = ~n14762 & ~n15442;
  assign n14432 = ~n14763;
  assign n14439 = ~n15402 | ~n14432;
  assign n14435 = ~n15438 & ~n14751;
  assign n14433 = ~P1_REG3_REG_20__SCAN_IN;
  assign n14434 = ~P1_STATE_REG_SCAN_IN & ~n14433;
  assign n14437 = n14435 | n14434;
  assign n14436 = n15429 & n14509;
  assign n14438 = ~n14437 & ~n14436;
  assign n14440 = ~n14439 | ~n14438;
  assign n14442 = ~n14441 & ~n14440;
  assign P1_U3231 = ~n14443 | ~n14442;
  assign n14446 = ~n14445;
  assign n14451 = ~n14447 & ~n14446;
  assign n14450 = ~n14449 | ~n14448;
  assign n14452 = ~n14451 ^ n14450;
  assign n14462 = ~n14452 | ~n15457;
  assign n14460 = ~n9692 & ~n15442;
  assign n14458 = ~n15402 | ~n14948;
  assign n14454 = ~n15429 | ~n14453;
  assign n15702 = ~P1_REG3_REG_13__SCAN_IN | ~P1_U3084;
  assign n14456 = ~n14454 | ~n15702;
  assign n14455 = ~n15438 & ~n14937;
  assign n14457 = ~n14456 & ~n14455;
  assign n14459 = ~n14458 | ~n14457;
  assign n14461 = ~n14460 & ~n14459;
  assign P1_U3232 = ~n14462 | ~n14461;
  assign n14465 = ~n14464 ^ n14463;
  assign n14467 = ~n14466 ^ n14465;
  assign n14480 = ~n14467 | ~n15457;
  assign n14478 = ~n15091 | ~n15421;
  assign n14476 = ~n14468 & ~n15438;
  assign n14474 = ~n15402 | ~n14469;
  assign n14472 = ~n15441 & ~n14751;
  assign n14471 = ~P1_STATE_REG_SCAN_IN & ~n14470;
  assign n14473 = ~n14472 & ~n14471;
  assign n14475 = ~n14474 | ~n14473;
  assign n14477 = ~n14476 & ~n14475;
  assign n14479 = n14478 & n14477;
  assign P1_U3233 = ~n14480 | ~n14479;
  assign n14488 = ~n14482 | ~n14481;
  assign n14485 = ~n14484 | ~n14483;
  assign n14487 = ~n14486 | ~n14485;
  assign n14489 = n14488 ^ n14487;
  assign n14499 = ~n14489 & ~n15414;
  assign n14497 = ~n15402 | ~n15005;
  assign n14495 = ~n15209 | ~n15421;
  assign n14491 = ~n15429 | ~n14490;
  assign n15677 = ~P1_REG3_REG_11__SCAN_IN | ~P1_U3084;
  assign n14493 = ~n14491 | ~n15677;
  assign n14492 = ~n15438 & ~n14993;
  assign n14494 = ~n14493 & ~n14492;
  assign n14496 = n14495 & n14494;
  assign n14498 = ~n14497 | ~n14496;
  assign P1_U3234 = n14499 | n14498;
  assign n14501 = ~n14500;
  assign n14507 = ~n14501 | ~n14502;
  assign n14505 = ~n14503 | ~n14502;
  assign n14506 = ~n14505 | ~n14504;
  assign n14508 = ~n14507 | ~n14506;
  assign n14518 = ~n14508 | ~n15457;
  assign n14816 = ~n15134;
  assign n14516 = ~n14816 & ~n15442;
  assign n14514 = ~n15402 | ~n14817;
  assign n14510 = ~n15419 | ~n14509;
  assign n15791 = ~P1_REG3_REG_18__SCAN_IN | ~P1_U3084;
  assign n14512 = ~n14510 | ~n15791;
  assign n14511 = n15429 & n14859;
  assign n14513 = ~n14512 & ~n14511;
  assign n14515 = ~n14514 | ~n14513;
  assign n14517 = ~n14516 & ~n14515;
  assign P1_U3236 = ~n14518 | ~n14517;
  assign n14528 = ~n15047 | ~n15421;
  assign n14526 = ~n14608 & ~n15441;
  assign n14524 = ~n15402 | ~n14623;
  assign n14522 = ~n15419 | ~n16413;
  assign n14521 = ~P1_REG3_REG_26__SCAN_IN | ~P1_U3084;
  assign n14523 = n14522 & n14521;
  assign n14525 = ~n14524 | ~n14523;
  assign n14527 = ~n14526 & ~n14525;
  assign n14532 = ~n14531 ^ n14530;
  assign n14543 = ~n14532 | ~n15457;
  assign n14541 = ~n9689 & ~n15442;
  assign n14539 = ~n15402 | ~n14895;
  assign n14534 = ~n15419 | ~n14533;
  assign n15736 = ~P1_REG3_REG_15__SCAN_IN | ~P1_U3084;
  assign n14537 = ~n14534 | ~n15736;
  assign n14536 = n15429 & n14535;
  assign n14538 = ~n14537 & ~n14536;
  assign n14540 = ~n14539 | ~n14538;
  assign n14542 = ~n14541 & ~n14540;
  assign P1_U3239 = ~n14543 | ~n14542;
  assign n14551 = n14544 | n16040;
  assign n14549 = ~n14545 & ~n15996;
  assign n15017 = ~n14546;
  assign n14554 = ~n16119 | ~n15017;
  assign n14547 = ~n16104 | ~P1_REG2_REG_31__SCAN_IN;
  assign n14548 = ~n14554 | ~n14547;
  assign n14550 = ~n14549 & ~n14548;
  assign P1_U3261 = ~n14551 | ~n14550;
  assign n15015 = n14552 ^ n15016;
  assign n14558 = ~n15015 | ~n16109;
  assign n14556 = ~n15016 & ~n15996;
  assign n14553 = ~n16104 | ~P1_REG2_REG_30__SCAN_IN;
  assign n14555 = ~n14554 | ~n14553;
  assign n14557 = ~n14556 & ~n14555;
  assign P1_U3262 = ~n14558 | ~n14557;
  assign n14561 = ~n14560 ^ n14559;
  assign n14566 = ~n14561 | ~n16055;
  assign n14564 = ~n14562 & ~n16025;
  assign n14563 = ~n14609 & ~n16023;
  assign n14565 = ~n14564 & ~n14563;
  assign n14570 = ~n14566 | ~n14565;
  assign n14569 = ~n15023 & ~n16045;
  assign n14572 = ~n15031 | ~n16119;
  assign n14571 = n16119 | P1_REG2_REG_28__SCAN_IN;
  assign n14583 = ~n14572 | ~n14571;
  assign n14581 = ~n15023 & ~n16003;
  assign n14579 = ~n15024 | ~n16109;
  assign n14577 = ~n15025 & ~n15996;
  assign n14575 = ~n14574;
  assign n14576 = ~n16011 & ~n14575;
  assign n14578 = ~n14577 & ~n14576;
  assign n14580 = ~n14579 | ~n14578;
  assign n14582 = ~n14581 & ~n14580;
  assign P1_U3263 = ~n14583 | ~n14582;
  assign n14585 = ~n14584 ^ n9616;
  assign n14591 = ~n14585 | ~n16055;
  assign n14589 = ~n14586 & ~n16023;
  assign n14588 = ~n14587 & ~n16025;
  assign n14590 = ~n14589 & ~n14588;
  assign n15039 = ~n14591 | ~n14590;
  assign n14593 = ~n15039 & ~n16104;
  assign n14592 = ~n16119 & ~P1_REG2_REG_27__SCAN_IN;
  assign n14603 = ~n14593 & ~n14592;
  assign n15040 = ~n14594 ^ n9616;
  assign n14595 = ~n16119 | ~n16084;
  assign n14643 = ~n16003 | ~n14595;
  assign n14601 = n15034 & n16109;
  assign n14599 = ~n15035 | ~n16108;
  assign n14598 = ~n16105 | ~n14597;
  assign n14600 = ~n14599 | ~n14598;
  assign n14602 = ~n14601 & ~n14600;
  assign n14606 = ~n14604 | ~n14605;
  assign n14607 = ~n14606 ^ n14614;
  assign n14613 = ~n14607 | ~n16055;
  assign n14611 = ~n14608 & ~n16023;
  assign n14610 = ~n14609 & ~n16025;
  assign n14612 = ~n14611 & ~n14610;
  assign n14618 = ~n14613 | ~n14612;
  assign n14615 = ~n14614;
  assign n15045 = ~n14616 ^ n14615;
  assign n14617 = ~n15045 & ~n16045;
  assign n15053 = ~n14618 & ~n14617;
  assign n14620 = ~n15053 | ~n16119;
  assign n14619 = n16119 | P1_REG2_REG_26__SCAN_IN;
  assign n14632 = ~n14620 | ~n14619;
  assign n14630 = ~n15045 & ~n16003;
  assign n15046 = ~n14621 ^ n15047;
  assign n14628 = ~n15046 | ~n16109;
  assign n14626 = ~n14622 & ~n15996;
  assign n14624 = ~n14623;
  assign n14625 = ~n14624 & ~n16011;
  assign n14627 = ~n14626 & ~n14625;
  assign n14629 = ~n14628 | ~n14627;
  assign n14631 = ~n14630 & ~n14629;
  assign P1_U3265 = ~n14632 | ~n14631;
  assign n14634 = n14641 ^ n14633;
  assign n14638 = ~n14634 & ~n16074;
  assign n14636 = ~n16410 | ~n16116;
  assign n14635 = ~n16404 | ~n16077;
  assign n14637 = ~n14636 | ~n14635;
  assign n14640 = ~n15065 | ~n16119;
  assign n14639 = n16119 | P1_REG2_REG_25__SCAN_IN;
  assign n14653 = ~n14640 | ~n14639;
  assign n15057 = n14642 ^ n14641;
  assign n14651 = ~n15057 & ~n14918;
  assign n15058 = n15059 ^ n14666;
  assign n14649 = ~n15058 | ~n16109;
  assign n14647 = ~n14644 & ~n15996;
  assign n14646 = ~n14645 & ~n16011;
  assign n14648 = ~n14647 & ~n14646;
  assign n14650 = ~n14649 | ~n14648;
  assign n14652 = ~n14651 & ~n14650;
  assign P1_U3266 = ~n14653 | ~n14652;
  assign n14655 = n14660 ^ n14654;
  assign n14659 = ~n14655 & ~n16074;
  assign n14657 = ~n16407 | ~n16116;
  assign n14656 = ~n16401 | ~n16077;
  assign n14658 = ~n14657 | ~n14656;
  assign n15075 = ~n14659 & ~n14658;
  assign n15068 = ~n14661 ^ n14660;
  assign n14662 = ~n16095;
  assign n14732 = ~n16084 & ~n14662;
  assign n14675 = ~n15068 & ~n14732;
  assign n14664 = ~n14663;
  assign n14665 = ~n15069 | ~n14664;
  assign n14668 = ~n14665 | ~n16350;
  assign n14667 = ~n14666;
  assign n15071 = n14668 | n14667;
  assign n14673 = ~n15071 & ~n16090;
  assign n16092 = ~n16059;
  assign n14671 = ~n15069 | ~n16092;
  assign n14670 = ~n16105 | ~n14669;
  assign n14672 = ~n14671 | ~n14670;
  assign n14674 = n14673 | n14672;
  assign n14676 = ~n14675 & ~n14674;
  assign n14677 = ~n15075 | ~n14676;
  assign n14679 = ~n14677 | ~n16119;
  assign n14678 = ~n16104 | ~P1_REG2_REG_24__SCAN_IN;
  assign P1_U3267 = ~n14679 | ~n14678;
  assign n14682 = ~n14681 ^ n14680;
  assign n14686 = ~n14682 & ~n16074;
  assign n14684 = ~n16398 | ~n16077;
  assign n14683 = ~n16404 | ~n16116;
  assign n14685 = ~n14684 | ~n14683;
  assign n15086 = ~n14686 & ~n14685;
  assign n14688 = ~n15086 | ~n16119;
  assign n14687 = n16119 | P1_REG2_REG_23__SCAN_IN;
  assign n14700 = ~n14688 | ~n14687;
  assign n15078 = ~n14689 ^ n14690;
  assign n14698 = ~n15078 & ~n14918;
  assign n15079 = ~n14713 ^ n14691;
  assign n14696 = ~n15079 | ~n16109;
  assign n14694 = ~n14691 & ~n15996;
  assign n14693 = ~n14692 & ~n16011;
  assign n14695 = ~n14694 & ~n14693;
  assign n14697 = ~n14696 | ~n14695;
  assign n14699 = ~n14698 & ~n14697;
  assign P1_U3268 = ~n14700 | ~n14699;
  assign n14702 = ~n14701 ^ n14710;
  assign n14707 = ~n14702 & ~n16074;
  assign n14705 = ~n16401 | ~n16116;
  assign n14704 = ~n14703 | ~n16077;
  assign n14706 = ~n14705 | ~n14704;
  assign n15097 = ~n14707 & ~n14706;
  assign n14709 = ~n15097 | ~n16119;
  assign n14708 = n16119 | P1_REG2_REG_22__SCAN_IN;
  assign n14723 = ~n14709 | ~n14708;
  assign n15089 = ~n14711 ^ n14710;
  assign n14721 = ~n15089 & ~n14918;
  assign n14712 = ~n14735 | ~n15091;
  assign n15090 = n14713 & n14712;
  assign n14719 = ~n15090 | ~n16109;
  assign n14717 = ~n14714 & ~n15996;
  assign n14716 = ~n14715 & ~n16011;
  assign n14718 = ~n14717 & ~n14716;
  assign n14720 = ~n14719 | ~n14718;
  assign n14722 = ~n14721 & ~n14720;
  assign P1_U3269 = ~n14723 | ~n14722;
  assign n14725 = n14724 ^ n14730;
  assign n14729 = ~n14725 & ~n16074;
  assign n14727 = ~n16398 | ~n16116;
  assign n14726 = ~n14774 | ~n16077;
  assign n14728 = ~n14727 | ~n14726;
  assign n15107 = ~n14729 & ~n14728;
  assign n15100 = ~n14731 ^ n14730;
  assign n14744 = ~n15100 & ~n14732;
  assign n14734 = n14733 | n14737;
  assign n14736 = n14734 & n16350;
  assign n15103 = ~n14736 | ~n14735;
  assign n14742 = n15103 | n16090;
  assign n14740 = ~n14737 & ~n16059;
  assign n14739 = ~n14738 & ~n16011;
  assign n14741 = ~n14740 & ~n14739;
  assign n14743 = ~n14742 | ~n14741;
  assign n14745 = ~n14744 & ~n14743;
  assign n14746 = ~n15107 | ~n14745;
  assign n14748 = ~n14746 | ~n16119;
  assign n14747 = ~n16104 | ~P1_REG2_REG_21__SCAN_IN;
  assign P1_U3270 = ~n14748 | ~n14747;
  assign n14750 = ~n14749 ^ n14756;
  assign n14755 = ~n14750 | ~n16055;
  assign n14753 = ~n14751 & ~n16025;
  assign n14752 = ~n14803 & ~n16023;
  assign n14754 = ~n14753 & ~n14752;
  assign n14759 = ~n14755 | ~n14754;
  assign n15110 = ~n14757 ^ n14756;
  assign n14758 = ~n15110 & ~n16045;
  assign n15118 = ~n14759 & ~n14758;
  assign n14761 = ~n15118 | ~n16119;
  assign n14760 = n16119 | P1_REG2_REG_20__SCAN_IN;
  assign n14771 = ~n14761 | ~n14760;
  assign n14769 = ~n15110 & ~n16003;
  assign n15111 = ~n14792 ^ n15112;
  assign n14767 = ~n15111 | ~n16109;
  assign n14765 = ~n14762 & ~n15996;
  assign n14764 = ~n16011 & ~n14763;
  assign n14766 = ~n14765 & ~n14764;
  assign n14768 = ~n14767 | ~n14766;
  assign n14770 = ~n14769 & ~n14768;
  assign P1_U3271 = ~n14771 | ~n14770;
  assign n14773 = n14772 ^ n14789;
  assign n14779 = ~n14773 & ~n16074;
  assign n14777 = ~n14774 | ~n16116;
  assign n14776 = ~n14775 | ~n16077;
  assign n14778 = ~n14777 | ~n14776;
  assign n15129 = ~n14779 & ~n14778;
  assign n14781 = ~n14780;
  assign n14782 = ~n16011 & ~n14781;
  assign n14783 = ~n16104 & ~n14782;
  assign n14785 = ~n15129 | ~n14783;
  assign n15827 = ~P1_REG2_REG_19__SCAN_IN;
  assign n14784 = ~n16104 | ~n15827;
  assign n14798 = ~n14785 | ~n14784;
  assign n14787 = ~n9045 | ~n14809;
  assign n14788 = ~n14787 | ~n14786;
  assign n15121 = n14789 ^ n14788;
  assign n14796 = ~n15121 & ~n14918;
  assign n14791 = n14790 & n15123;
  assign n15122 = ~n14792 & ~n14791;
  assign n14794 = ~n15122 | ~n16109;
  assign n14793 = ~n15123 | ~n16108;
  assign n14795 = ~n14794 | ~n14793;
  assign n14797 = ~n14796 & ~n14795;
  assign P1_U3272 = ~n14798 | ~n14797;
  assign n14801 = ~n14799 | ~n14800;
  assign n14802 = ~n14801 ^ n14809;
  assign n14808 = ~n14802 | ~n16055;
  assign n14806 = ~n14803 & ~n16025;
  assign n14805 = ~n14804 & ~n16023;
  assign n14807 = ~n14806 & ~n14805;
  assign n14811 = ~n14808 | ~n14807;
  assign n15132 = ~n9045 ^ n14809;
  assign n14810 = ~n15132 & ~n16045;
  assign n15140 = ~n14811 & ~n14810;
  assign n14814 = ~n15140 | ~n16119;
  assign n14812 = ~P1_REG2_REG_18__SCAN_IN;
  assign n14813 = ~n16104 | ~n14812;
  assign n14826 = ~n14814 | ~n14813;
  assign n14824 = ~n15132 & ~n16003;
  assign n15133 = ~n14815 ^ n14816;
  assign n14822 = ~n15133 | ~n16109;
  assign n14820 = ~n14816 & ~n15996;
  assign n14818 = ~n14817;
  assign n14819 = ~n16011 & ~n14818;
  assign n14821 = ~n14820 & ~n14819;
  assign n14823 = ~n14822 | ~n14821;
  assign n14825 = ~n14824 & ~n14823;
  assign P1_U3273 = ~n14826 | ~n14825;
  assign n14827 = n9139 ^ n14835;
  assign n14832 = ~n14827 | ~n16055;
  assign n14830 = ~n14885 & ~n16023;
  assign n14829 = ~n14828 & ~n16025;
  assign n14831 = ~n14830 & ~n14829;
  assign n14839 = ~n14832 | ~n14831;
  assign n14837 = ~n14834 | ~n14833;
  assign n14836 = ~n14835;
  assign n15143 = ~n14837 ^ n14836;
  assign n14838 = ~n15143 & ~n16045;
  assign n15151 = ~n14839 & ~n14838;
  assign n14842 = ~n15151 | ~n16119;
  assign n14840 = ~P1_REG2_REG_17__SCAN_IN;
  assign n14841 = ~n16104 | ~n14840;
  assign n14853 = ~n14842 | ~n14841;
  assign n14851 = ~n15143 & ~n16003;
  assign n15144 = ~n14871 ^ n15145;
  assign n14849 = ~n15144 | ~n16109;
  assign n14847 = ~n14843 & ~n15996;
  assign n14845 = ~n14844;
  assign n14846 = ~n16011 & ~n14845;
  assign n14848 = ~n14847 & ~n14846;
  assign n14850 = ~n14849 | ~n14848;
  assign n14852 = ~n14851 & ~n14850;
  assign P1_U3274 = ~n14853 | ~n14852;
  assign n14855 = ~n14854;
  assign n14857 = ~n14856 & ~n14855;
  assign n14858 = ~n14857 ^ n14867;
  assign n14863 = ~n14858 & ~n16074;
  assign n14861 = ~n14859 | ~n16116;
  assign n14860 = ~n14908 | ~n16077;
  assign n14862 = ~n14861 | ~n14860;
  assign n15161 = ~n14863 & ~n14862;
  assign n14866 = ~n15161 | ~n16119;
  assign n14864 = ~P1_REG2_REG_16__SCAN_IN;
  assign n14865 = ~n16104 | ~n14864;
  assign n14880 = ~n14866 | ~n14865;
  assign n15154 = ~n14868 ^ n14867;
  assign n14878 = ~n15154 & ~n14918;
  assign n14869 = ~n9147 | ~n15155;
  assign n14870 = ~n14869 | ~n16350;
  assign n15157 = n14871 | n14870;
  assign n14876 = ~n15157 & ~n14979;
  assign n14874 = ~n15155 | ~n16108;
  assign n14873 = ~n16105 | ~n14872;
  assign n14875 = ~n14874 | ~n14873;
  assign n14877 = n14876 | n14875;
  assign n14879 = ~n14878 & ~n14877;
  assign P1_U3275 = ~n14880 | ~n14879;
  assign n14882 = ~n14881 ^ n14883;
  assign n14891 = ~n14882 & ~n16074;
  assign n14894 = n14884 ^ n14883;
  assign n14889 = ~n14894 | ~n16084;
  assign n14887 = ~n14885 & ~n16025;
  assign n14886 = ~n14937 & ~n16023;
  assign n14888 = ~n14887 & ~n14886;
  assign n14890 = ~n14889 | ~n14888;
  assign n15172 = ~n14891 & ~n14890;
  assign n14893 = ~n15172 | ~n16119;
  assign n15741 = ~P1_REG2_REG_15__SCAN_IN;
  assign n14892 = ~n16104 | ~n15741;
  assign n14904 = ~n14893 | ~n14892;
  assign n15164 = ~n14894;
  assign n14902 = ~n15164 & ~n16003;
  assign n15165 = ~n14922 ^ n9689;
  assign n14900 = ~n15165 | ~n16109;
  assign n14898 = ~n9689 & ~n15996;
  assign n14896 = ~n14895;
  assign n14897 = ~n16011 & ~n14896;
  assign n14899 = ~n14898 & ~n14897;
  assign n14901 = ~n14900 | ~n14899;
  assign n14903 = ~n14902 & ~n14901;
  assign P1_U3276 = ~n14904 | ~n14903;
  assign n14906 = ~n14905 ^ n14916;
  assign n14912 = ~n14906 & ~n16074;
  assign n14910 = ~n14907 | ~n16077;
  assign n14909 = ~n14908 | ~n16116;
  assign n14911 = ~n14910 | ~n14909;
  assign n15183 = ~n14912 & ~n14911;
  assign n14915 = ~n15183 | ~n16119;
  assign n14913 = ~P1_REG2_REG_14__SCAN_IN;
  assign n14914 = ~n16104 | ~n14913;
  assign n14932 = ~n14915 | ~n14914;
  assign n15176 = ~n14917 ^ n14916;
  assign n14930 = ~n15176 & ~n14918;
  assign n14921 = n14920 | n14919;
  assign n14923 = ~n14921 | ~n16350;
  assign n15179 = n14923 | n9687;
  assign n14928 = ~n15179 & ~n14979;
  assign n14926 = ~n15177 | ~n16108;
  assign n14925 = ~n16105 | ~n14924;
  assign n14927 = ~n14926 | ~n14925;
  assign n14929 = n14928 | n14927;
  assign n14931 = ~n14930 & ~n14929;
  assign P1_U3277 = ~n14932 | ~n14931;
  assign n14934 = n14933 ^ n14935;
  assign n14943 = ~n14934 & ~n16074;
  assign n14947 = ~n14936 ^ n14935;
  assign n14941 = ~n14947 | ~n16084;
  assign n14939 = ~n14937 & ~n16025;
  assign n14938 = ~n14993 & ~n16023;
  assign n14940 = ~n14939 & ~n14938;
  assign n14942 = ~n14941 | ~n14940;
  assign n15194 = ~n14943 & ~n14942;
  assign n14946 = ~n15194 | ~n16119;
  assign n14944 = ~P1_REG2_REG_13__SCAN_IN;
  assign n14945 = ~n16104 | ~n14944;
  assign n14957 = ~n14946 | ~n14945;
  assign n15186 = ~n14947;
  assign n14955 = ~n15186 & ~n16003;
  assign n15187 = n15188 ^ n14977;
  assign n14953 = ~n15187 | ~n16109;
  assign n14951 = ~n9692 & ~n15996;
  assign n14949 = ~n14948;
  assign n14950 = ~n16011 & ~n14949;
  assign n14952 = ~n14951 & ~n14950;
  assign n14954 = ~n14953 | ~n14952;
  assign n14956 = ~n14955 & ~n14954;
  assign P1_U3278 = ~n14957 | ~n14956;
  assign n14960 = ~n14959 | ~n14958;
  assign n14961 = n14962 ^ n14960;
  assign n14971 = ~n14961 & ~n16074;
  assign n15197 = ~n14963 ^ n14962;
  assign n14969 = n15197 | n16045;
  assign n14967 = n14964 | n16023;
  assign n14966 = n14965 | n16025;
  assign n14968 = n14967 & n14966;
  assign n14970 = ~n14969 | ~n14968;
  assign n15204 = ~n14971 & ~n14970;
  assign n14974 = ~n15204 | ~n16119;
  assign n14972 = ~P1_REG2_REG_12__SCAN_IN;
  assign n14973 = ~n16104 | ~n14972;
  assign n14988 = ~n14974 | ~n14973;
  assign n14986 = ~n15197 & ~n16003;
  assign n14976 = ~n14975 | ~n15198;
  assign n14978 = n14976 & n16350;
  assign n15200 = ~n14978 | ~n14977;
  assign n14984 = ~n15200 & ~n14979;
  assign n14982 = ~n15198 | ~n16108;
  assign n14981 = ~n16105 | ~n14980;
  assign n14983 = ~n14982 | ~n14981;
  assign n14985 = n14984 | n14983;
  assign n14987 = ~n14986 & ~n14985;
  assign P1_U3279 = ~n14988 | ~n14987;
  assign n14990 = n14989 ^ n14991;
  assign n14999 = ~n14990 & ~n16074;
  assign n15002 = n14992 ^ n14991;
  assign n14997 = ~n15002 | ~n16084;
  assign n14995 = ~n14993 & ~n16025;
  assign n14994 = ~n15847 & ~n16023;
  assign n14996 = ~n14995 & ~n14994;
  assign n14998 = ~n14997 | ~n14996;
  assign n15215 = ~n14999 & ~n14998;
  assign n15001 = ~n15215 | ~n16119;
  assign n15675 = ~P1_REG2_REG_11__SCAN_IN;
  assign n15000 = ~n16104 | ~n15675;
  assign n15014 = ~n15001 | ~n15000;
  assign n15207 = ~n15002;
  assign n15012 = ~n15207 & ~n16003;
  assign n15208 = n15003 ^ n15209;
  assign n15010 = ~n15208 | ~n16109;
  assign n15004 = ~n15209;
  assign n15008 = ~n15004 & ~n15996;
  assign n15006 = ~n15005;
  assign n15007 = ~n16011 & ~n15006;
  assign n15009 = ~n15008 & ~n15007;
  assign n15011 = ~n15010 | ~n15009;
  assign n15013 = ~n15012 & ~n15011;
  assign P1_U3280 = ~n15014 | ~n15013;
  assign n15020 = ~n15015 | ~n16350;
  assign n15018 = ~n15016 & ~n16309;
  assign n15019 = ~n15018 & ~n15017;
  assign n15218 = ~n15020 | ~n15019;
  assign n15022 = ~n15218 | ~n16395;
  assign n15021 = ~n16393 | ~P1_REG1_REG_30__SCAN_IN;
  assign P1_U3553 = ~n15022 | ~n15021;
  assign n15029 = ~n15023 & ~n16357;
  assign n15027 = ~n15024 | ~n16350;
  assign n15026 = ~n9698 | ~n16352;
  assign n15028 = ~n15027 | ~n15026;
  assign n15030 = ~n15029 & ~n15028;
  assign n15221 = ~n15031 | ~n15030;
  assign n15033 = ~n15221 | ~n16395;
  assign n15032 = ~n16393 | ~P1_REG1_REG_28__SCAN_IN;
  assign P1_U3551 = ~n15033 | ~n15032;
  assign n15037 = ~n15034 | ~n16350;
  assign n15036 = ~n15035 | ~n16352;
  assign n15038 = ~n15037 | ~n15036;
  assign n15042 = ~n15039 & ~n15038;
  assign n15056 = ~n16045 | ~n16357;
  assign n15041 = ~n15040 | ~n15056;
  assign n15224 = ~n15042 | ~n15041;
  assign n15044 = ~n15224 | ~n16395;
  assign n15043 = ~n16393 | ~P1_REG1_REG_27__SCAN_IN;
  assign P1_U3550 = ~n15044 | ~n15043;
  assign n15051 = ~n15045 & ~n16357;
  assign n15049 = ~n15046 | ~n16350;
  assign n15048 = ~n15047 | ~n16352;
  assign n15050 = ~n15049 | ~n15048;
  assign n15052 = ~n15051 & ~n15050;
  assign n15227 = ~n15053 | ~n15052;
  assign n15055 = ~n15227 | ~n16395;
  assign n15054 = ~n16393 | ~P1_REG1_REG_26__SCAN_IN;
  assign P1_U3549 = ~n15055 | ~n15054;
  assign n15063 = ~n15057 & ~n15175;
  assign n15061 = ~n15058 | ~n16350;
  assign n15060 = ~n15059 | ~n16352;
  assign n15062 = ~n15061 | ~n15060;
  assign n15064 = ~n15063 & ~n15062;
  assign n15230 = ~n15065 | ~n15064;
  assign n15067 = ~n15230 | ~n16395;
  assign n15066 = ~n16393 | ~P1_REG1_REG_25__SCAN_IN;
  assign P1_U3548 = ~n15067 | ~n15066;
  assign n15073 = ~n15068 & ~n15175;
  assign n15070 = ~n15069 | ~n16352;
  assign n15072 = ~n15071 | ~n15070;
  assign n15074 = ~n15073 & ~n15072;
  assign n15233 = ~n15075 | ~n15074;
  assign n15077 = ~n15233 | ~n16395;
  assign n15076 = ~n16393 | ~P1_REG1_REG_24__SCAN_IN;
  assign P1_U3547 = ~n15077 | ~n15076;
  assign n15084 = ~n15078 & ~n15175;
  assign n15082 = ~n15079 | ~n16350;
  assign n15081 = ~n15080 | ~n16352;
  assign n15083 = ~n15082 | ~n15081;
  assign n15085 = ~n15084 & ~n15083;
  assign n15236 = ~n15086 | ~n15085;
  assign n15088 = ~n15236 | ~n16395;
  assign n15087 = ~n16393 | ~P1_REG1_REG_23__SCAN_IN;
  assign P1_U3546 = ~n15088 | ~n15087;
  assign n15095 = ~n15089 & ~n15175;
  assign n15093 = ~n15090 | ~n16350;
  assign n15092 = ~n15091 | ~n16352;
  assign n15094 = ~n15093 | ~n15092;
  assign n15096 = ~n15095 & ~n15094;
  assign n15239 = ~n15097 | ~n15096;
  assign n15099 = ~n15239 | ~n16395;
  assign n15098 = ~n16393 | ~P1_REG1_REG_22__SCAN_IN;
  assign P1_U3545 = ~n15099 | ~n15098;
  assign n15105 = ~n15100 & ~n15175;
  assign n15102 = ~n15101 | ~n16352;
  assign n15104 = ~n15103 | ~n15102;
  assign n15106 = ~n15105 & ~n15104;
  assign n15242 = ~n15107 | ~n15106;
  assign n15109 = ~n15242 | ~n16395;
  assign n15108 = ~n16393 | ~P1_REG1_REG_21__SCAN_IN;
  assign P1_U3544 = ~n15109 | ~n15108;
  assign n15116 = ~n15110 & ~n16357;
  assign n15114 = ~n15111 | ~n16350;
  assign n15113 = ~n15112 | ~n16352;
  assign n15115 = ~n15114 | ~n15113;
  assign n15117 = ~n15116 & ~n15115;
  assign n15245 = ~n15118 | ~n15117;
  assign n15120 = ~n15245 | ~n16395;
  assign n15119 = ~n16393 | ~P1_REG1_REG_20__SCAN_IN;
  assign P1_U3543 = ~n15120 | ~n15119;
  assign n15127 = ~n15121 & ~n15175;
  assign n15125 = ~n15122 | ~n16350;
  assign n15124 = ~n15123 | ~n16352;
  assign n15126 = ~n15125 | ~n15124;
  assign n15128 = ~n15127 & ~n15126;
  assign n15248 = ~n15129 | ~n15128;
  assign n15131 = ~n15248 | ~n16395;
  assign n15130 = ~n16393 | ~P1_REG1_REG_19__SCAN_IN;
  assign P1_U3542 = ~n15131 | ~n15130;
  assign n15138 = ~n15132 & ~n16357;
  assign n15136 = ~n15133 | ~n16350;
  assign n15135 = ~n15134 | ~n16352;
  assign n15137 = ~n15136 | ~n15135;
  assign n15139 = ~n15138 & ~n15137;
  assign n15251 = ~n15140 | ~n15139;
  assign n15142 = ~n15251 | ~n16395;
  assign n15141 = ~n16393 | ~P1_REG1_REG_18__SCAN_IN;
  assign P1_U3541 = ~n15142 | ~n15141;
  assign n15149 = ~n15143 & ~n16357;
  assign n15147 = ~n15144 | ~n16350;
  assign n15146 = ~n15145 | ~n16352;
  assign n15148 = ~n15147 | ~n15146;
  assign n15150 = ~n15149 & ~n15148;
  assign n15254 = ~n15151 | ~n15150;
  assign n15153 = ~n15254 | ~n16395;
  assign n15152 = ~n16393 | ~P1_REG1_REG_17__SCAN_IN;
  assign P1_U3540 = ~n15153 | ~n15152;
  assign n15159 = ~n15154 & ~n15175;
  assign n15156 = ~n15155 | ~n16352;
  assign n15158 = ~n15157 | ~n15156;
  assign n15160 = ~n15159 & ~n15158;
  assign n15257 = ~n15161 | ~n15160;
  assign n15163 = ~n15257 | ~n16395;
  assign n15162 = ~n16393 | ~P1_REG1_REG_16__SCAN_IN;
  assign P1_U3539 = ~n15163 | ~n15162;
  assign n15170 = ~n15164 & ~n16357;
  assign n15168 = ~n15165 | ~n16350;
  assign n15167 = ~n15166 | ~n16352;
  assign n15169 = ~n15168 | ~n15167;
  assign n15171 = ~n15170 & ~n15169;
  assign n15260 = ~n15172 | ~n15171;
  assign n15174 = ~n15260 | ~n16395;
  assign n15173 = ~n16393 | ~P1_REG1_REG_15__SCAN_IN;
  assign P1_U3538 = ~n15174 | ~n15173;
  assign n15181 = ~n15176 & ~n15175;
  assign n15178 = ~n15177 | ~n16352;
  assign n15180 = ~n15179 | ~n15178;
  assign n15182 = ~n15181 & ~n15180;
  assign n15263 = ~n15183 | ~n15182;
  assign n15185 = ~n15263 | ~n16395;
  assign n15184 = ~n16393 | ~P1_REG1_REG_14__SCAN_IN;
  assign P1_U3537 = ~n15185 | ~n15184;
  assign n15192 = ~n15186 & ~n16357;
  assign n15190 = ~n15187 | ~n16350;
  assign n15189 = ~n15188 | ~n16352;
  assign n15191 = ~n15190 | ~n15189;
  assign n15193 = ~n15192 & ~n15191;
  assign n15266 = ~n15194 | ~n15193;
  assign n15196 = ~n15266 | ~n16395;
  assign n15195 = ~n16393 | ~P1_REG1_REG_13__SCAN_IN;
  assign P1_U3536 = ~n15196 | ~n15195;
  assign n15202 = ~n15197 & ~n16357;
  assign n15199 = ~n15198 | ~n16352;
  assign n15201 = ~n15200 | ~n15199;
  assign n15203 = ~n15202 & ~n15201;
  assign n15269 = ~n15204 | ~n15203;
  assign n15206 = ~n15269 | ~n16395;
  assign n15205 = ~n16393 | ~P1_REG1_REG_12__SCAN_IN;
  assign P1_U3535 = ~n15206 | ~n15205;
  assign n15213 = ~n15207 & ~n16357;
  assign n15211 = ~n15208 | ~n16350;
  assign n15210 = ~n15209 | ~n16352;
  assign n15212 = ~n15211 | ~n15210;
  assign n15214 = ~n15213 & ~n15212;
  assign n15272 = ~n15215 | ~n15214;
  assign n15217 = ~n15272 | ~n16395;
  assign n15216 = ~n16393 | ~P1_REG1_REG_11__SCAN_IN;
  assign P1_U3534 = ~n15217 | ~n15216;
  assign n15220 = ~n15218 | ~n16363;
  assign n15219 = ~n16349 | ~P1_REG0_REG_30__SCAN_IN;
  assign P1_U3521 = ~n15220 | ~n15219;
  assign n15223 = ~n15221 | ~n16363;
  assign n15222 = ~n16349 | ~P1_REG0_REG_28__SCAN_IN;
  assign P1_U3519 = ~n15223 | ~n15222;
  assign n15226 = ~n15224 | ~n16363;
  assign n15225 = ~n16349 | ~P1_REG0_REG_27__SCAN_IN;
  assign P1_U3518 = ~n15226 | ~n15225;
  assign n15229 = ~n15227 | ~n16363;
  assign n15228 = ~n16349 | ~P1_REG0_REG_26__SCAN_IN;
  assign P1_U3517 = ~n15229 | ~n15228;
  assign n15232 = ~n15230 | ~n16363;
  assign n15231 = ~n16349 | ~P1_REG0_REG_25__SCAN_IN;
  assign P1_U3516 = ~n15232 | ~n15231;
  assign n15235 = ~n15233 | ~n16363;
  assign n15234 = ~n16349 | ~P1_REG0_REG_24__SCAN_IN;
  assign P1_U3515 = ~n15235 | ~n15234;
  assign n15238 = ~n15236 | ~n16363;
  assign n15237 = ~n16349 | ~P1_REG0_REG_23__SCAN_IN;
  assign P1_U3514 = ~n15238 | ~n15237;
  assign n15241 = ~n15239 | ~n16363;
  assign n15240 = ~n16349 | ~P1_REG0_REG_22__SCAN_IN;
  assign P1_U3513 = ~n15241 | ~n15240;
  assign n15244 = ~n15242 | ~n16363;
  assign n15243 = ~n16349 | ~P1_REG0_REG_21__SCAN_IN;
  assign P1_U3512 = ~n15244 | ~n15243;
  assign n15247 = ~n15245 | ~n16363;
  assign n15246 = ~n16349 | ~P1_REG0_REG_20__SCAN_IN;
  assign P1_U3511 = ~n15247 | ~n15246;
  assign n15250 = ~n15248 | ~n16363;
  assign n15249 = ~n16349 | ~P1_REG0_REG_19__SCAN_IN;
  assign P1_U3510 = ~n15250 | ~n15249;
  assign n15253 = ~n15251 | ~n16363;
  assign n15252 = ~n16349 | ~P1_REG0_REG_18__SCAN_IN;
  assign P1_U3508 = ~n15253 | ~n15252;
  assign n15256 = ~n15254 | ~n16363;
  assign n15255 = ~n16349 | ~P1_REG0_REG_17__SCAN_IN;
  assign P1_U3505 = ~n15256 | ~n15255;
  assign n15259 = ~n15257 | ~n16363;
  assign n15258 = ~n16349 | ~P1_REG0_REG_16__SCAN_IN;
  assign P1_U3502 = ~n15259 | ~n15258;
  assign n15262 = ~n15260 | ~n16363;
  assign n15261 = ~n16349 | ~P1_REG0_REG_15__SCAN_IN;
  assign P1_U3499 = ~n15262 | ~n15261;
  assign n15265 = ~n15263 | ~n16363;
  assign n15264 = ~n16349 | ~P1_REG0_REG_14__SCAN_IN;
  assign P1_U3496 = ~n15265 | ~n15264;
  assign n15268 = ~n15266 | ~n16363;
  assign n15267 = ~n16349 | ~P1_REG0_REG_13__SCAN_IN;
  assign P1_U3493 = ~n15268 | ~n15267;
  assign n15271 = ~n15269 | ~n16363;
  assign n15270 = ~n16349 | ~P1_REG0_REG_12__SCAN_IN;
  assign P1_U3490 = ~n15271 | ~n15270;
  assign n15274 = ~n15272 | ~n16363;
  assign n15273 = ~n16349 | ~P1_REG0_REG_11__SCAN_IN;
  assign P1_U3487 = ~n15274 | ~n15273;
  assign n15284 = ~n15275 | ~n15317;
  assign n15278 = ~P1_U3084 & ~n11228;
  assign n15279 = ~n15278 | ~n15277;
  assign n15282 = ~n15276 & ~n15279;
  assign n15280 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n15281 = ~n16128 & ~n15280;
  assign n15283 = ~n15282 & ~n15281;
  assign P1_U3322 = ~n15284 | ~n15283;
  assign n15291 = ~n15285 | ~n15317;
  assign n15289 = ~n15286 & ~P1_U3084;
  assign n15288 = ~n16128 & ~n15287;
  assign n15290 = ~n15289 & ~n15288;
  assign P1_U3323 = ~n15291 | ~n15290;
  assign n15297 = ~n15292 | ~n15317;
  assign n15295 = ~n11232 & ~P1_U3084;
  assign n15294 = ~n16128 & ~n15293;
  assign n15296 = ~n15295 & ~n15294;
  assign P1_U3324 = ~n15297 | ~n15296;
  assign n15303 = ~n15298 & ~n16225;
  assign n15301 = n11945 | P1_U3084;
  assign n15299 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n15300 = n16128 | n15299;
  assign n15302 = ~n15301 | ~n15300;
  assign P1_U3325 = n15303 | n15302;
  assign n15308 = ~n15304 | ~n15317;
  assign n15306 = ~n16128 & ~n15305;
  assign n15307 = ~n9160 & ~n15306;
  assign P1_U3326 = ~n15308 | ~n15307;
  assign n15316 = ~n15309 | ~n15317;
  assign n15311 = ~n15310;
  assign n15314 = ~n15311 & ~P1_U3084;
  assign n15313 = ~n16128 & ~n15312;
  assign n15315 = ~n15314 & ~n15313;
  assign P1_U3327 = ~n15316 | ~n15315;
  assign n15325 = ~n15318 | ~n15317;
  assign n15320 = ~n15319;
  assign n15323 = ~n15320 & ~P1_U3084;
  assign n15322 = ~n16128 & ~n15321;
  assign n15324 = ~n15323 & ~n15322;
  assign P1_U3329 = ~n15325 | ~n15324;
  assign U123 = ~P1_WR_REG_SCAN_IN ^ P2_WR_REG_SCAN_IN;
  assign U126 = ~P2_RD_REG_SCAN_IN ^ P1_RD_REG_SCAN_IN;
  assign n15329 = ~n15441 & ~n15326;
  assign n15327 = ~n16320;
  assign n15328 = ~n15442 & ~n15327;
  assign n15340 = ~n15329 & ~n15328;
  assign n15330 = ~n15419 | ~n15903;
  assign n15595 = ~P1_REG3_REG_7__SCAN_IN | ~P1_U3084;
  assign n15338 = ~n15330 | ~n15595;
  assign n15332 = ~n9021 | ~n15331;
  assign n15334 = ~n15333 ^ n15332;
  assign n15336 = ~n15334 | ~n15457;
  assign n15335 = ~n15914 | ~n15402;
  assign n15337 = ~n15336 | ~n15335;
  assign n15339 = ~n15338 & ~n15337;
  assign P1_U3211 = ~n15340 | ~n15339;
  assign n15342 = ~n15419 | ~n15972;
  assign n15346 = ~n15342 | ~n15341;
  assign n15344 = ~n15421 | ~n16274;
  assign n15343 = ~n15429 | ~n16076;
  assign n15345 = ~n15344 | ~n15343;
  assign n15358 = ~n15346 & ~n15345;
  assign n15350 = ~n15347;
  assign n15353 = ~n15348 & ~n15350;
  assign n15351 = ~n15350 & ~n15349;
  assign n15354 = ~n15353 & ~n15352;
  assign n15356 = ~n15354 & ~n15414;
  assign n15355 = ~P1_REG3_REG_3__SCAN_IN & ~n15447;
  assign n15357 = ~n15356 & ~n15355;
  assign P1_U3216 = ~n15358 | ~n15357;
  assign n15359 = ~n15419 | ~n15881;
  assign n15611 = ~P1_REG3_REG_8__SCAN_IN | ~P1_U3084;
  assign n15363 = ~n15359 | ~n15611;
  assign n15361 = ~n15421 | ~n16334;
  assign n15360 = ~n15429 | ~n15929;
  assign n15362 = ~n15361 | ~n15360;
  assign n15370 = ~n15363 & ~n15362;
  assign n15366 = n15365 ^ n15364;
  assign n15368 = ~n15366 & ~n15414;
  assign n15367 = ~n15447 & ~n15878;
  assign n15369 = ~n15368 & ~n15367;
  assign P1_U3219 = ~n15370 | ~n15369;
  assign n15371 = ~n16078;
  assign n15373 = ~n15441 & ~n15371;
  assign n15372 = ~n15442 & ~n16088;
  assign n15387 = ~n15373 & ~n15372;
  assign n15377 = n15376 ^ n15375;
  assign n15385 = ~n15377 & ~n15414;
  assign n15381 = ~n15379 & ~n15378;
  assign n15434 = ~n15381 | ~n15380;
  assign n15383 = ~P1_REG3_REG_1__SCAN_IN | ~n15434;
  assign n15382 = ~n15419 | ~n16076;
  assign n15384 = ~n15383 | ~n15382;
  assign n15386 = ~n15385 & ~n15384;
  assign P1_U3220 = ~n15387 | ~n15386;
  assign n15390 = ~n15441 & ~n15388;
  assign n15389 = ~n15442 & ~n16283;
  assign n15408 = ~n15390 & ~n15389;
  assign n15391 = ~n15419 | ~n15930;
  assign n15523 = ~P1_REG3_REG_4__SCAN_IN | ~P1_U3084;
  assign n15406 = ~n15391 | ~n15523;
  assign n15393 = ~n15392;
  assign n15400 = ~n15393 | ~n15396;
  assign n15398 = ~n15394;
  assign n15397 = ~n15396 | ~n15395;
  assign n15399 = ~n15398 | ~n15397;
  assign n15401 = ~n15400 | ~n15399;
  assign n15404 = ~n15401 | ~n15457;
  assign n15403 = ~n15402 | ~n15982;
  assign n15405 = ~n15404 | ~n15403;
  assign n15407 = ~n15406 & ~n15405;
  assign P1_U3228 = ~n15408 | ~n15407;
  assign n15410 = ~n15419 | ~n11249;
  assign n15409 = ~n15421 | ~n9487;
  assign n15416 = ~n15410 | ~n15409;
  assign n15413 = ~n15411;
  assign n15495 = ~n15412 ^ n15413;
  assign n15415 = ~n15495 & ~n15414;
  assign n15418 = ~n15416 & ~n15415;
  assign n15417 = ~P1_REG3_REG_0__SCAN_IN | ~n15434;
  assign P1_U3230 = ~n15418 | ~n15417;
  assign n15423 = ~n15419 | ~n16046;
  assign n15422 = ~n15421 | ~n15420;
  assign n15433 = ~n15423 | ~n15422;
  assign n15426 = ~n15425 | ~n15424;
  assign n15428 = ~n15427 ^ n15426;
  assign n15431 = ~n15428 | ~n15457;
  assign n15430 = ~n15429 | ~n11249;
  assign n15432 = ~n15431 | ~n15430;
  assign n15436 = ~n15433 & ~n15432;
  assign n15435 = ~P1_REG3_REG_2__SCAN_IN | ~n15434;
  assign P1_U3235 = ~n15436 | ~n15435;
  assign n15440 = ~n15438 & ~n15437;
  assign n15439 = ~P1_REG3_REG_6__SCAN_IN;
  assign n15556 = ~P1_STATE_REG_SCAN_IN & ~n15439;
  assign n15446 = ~n15440 & ~n15556;
  assign n15981 = ~n15930;
  assign n15444 = ~n15441 & ~n15981;
  assign n15443 = ~n15442 & ~n16310;
  assign n15445 = ~n15444 & ~n15443;
  assign n15449 = ~n15446 | ~n15445;
  assign n15448 = ~n15447 & ~n15943;
  assign n15460 = ~n15449 & ~n15448;
  assign n15456 = ~n15451 | ~n15450;
  assign n15453 = ~n15452;
  assign n15455 = ~n15454 | ~n15453;
  assign n15458 = n15456 ^ n15455;
  assign n15459 = ~n15458 | ~n15457;
  assign P1_U3237 = ~n15460 | ~n15459;
  assign n15461 = ~n15494 & ~P1_REG2_REG_0__SCAN_IN;
  assign n15499 = n15461 | n11945;
  assign n15462 = ~n15496 & ~P1_REG1_REG_0__SCAN_IN;
  assign n15463 = ~n15499 & ~n15462;
  assign n15464 = ~n15463 ^ n15502;
  assign n15467 = ~n15465 & ~n15464;
  assign n15466 = P1_U3084 & P1_REG3_REG_0__SCAN_IN;
  assign n15469 = ~n15467 & ~n15466;
  assign n15468 = ~n15818 | ~P1_ADDR_REG_0__SCAN_IN;
  assign P1_U3241 = ~n15469 | ~n15468;
  assign n15471 = ~P1_ADDR_REG_1__SCAN_IN | ~n15818;
  assign n15470 = ~P1_REG3_REG_1__SCAN_IN | ~P1_U3084;
  assign n15478 = ~n15471 | ~n15470;
  assign n15474 = n15473 ^ n15472;
  assign n15476 = ~n15816 | ~n15474;
  assign n15475 = ~n12098 | ~n16226;
  assign n15477 = ~n15476 | ~n15475;
  assign n15483 = ~n15478 & ~n15477;
  assign n15481 = ~n15480 ^ n15479;
  assign n15482 = ~n15830 | ~n15481;
  assign P1_U3242 = ~n15483 | ~n15482;
  assign n15486 = n15485 ^ n15484;
  assign n15488 = ~n15830 | ~n15486;
  assign n15487 = ~P1_REG3_REG_2__SCAN_IN | ~P1_U3084;
  assign n15493 = ~n15488 | ~n15487;
  assign n15491 = ~n15818 | ~P1_ADDR_REG_2__SCAN_IN;
  assign n15490 = ~n12098 | ~n15489;
  assign n15492 = ~n15491 | ~n15490;
  assign n15513 = ~n15493 & ~n15492;
  assign n15498 = ~n15495 | ~n15494;
  assign n15497 = ~n15496 | ~n15502;
  assign n15500 = ~n15498 | ~n15497;
  assign n15503 = ~n15499;
  assign n15501 = ~n15500 | ~n15503;
  assign n15505 = ~P1_U4006 | ~n15501;
  assign n15504 = ~n15503 & ~n15502;
  assign n15535 = ~n15505 & ~n15504;
  assign n15510 = ~n15816 | ~n15506;
  assign n15509 = ~n15508 & ~n15507;
  assign n15511 = ~n15510 & ~n15509;
  assign n15512 = ~n15535 & ~n15511;
  assign P1_U3243 = ~n15513 | ~n15512;
  assign n15517 = ~n15515 | ~n15514;
  assign n15516 = ~n16219 | ~P1_REG2_REG_3__SCAN_IN;
  assign n15520 = ~n15517 | ~n15516;
  assign n15550 = n16213 | P1_REG2_REG_4__SCAN_IN;
  assign n15518 = ~n16213 | ~P1_REG2_REG_4__SCAN_IN;
  assign n15519 = ~n15550 | ~n15518;
  assign n15551 = n15520 | n15519;
  assign n15521 = ~n15520 | ~n15519;
  assign n15522 = ~n15551 | ~n15521;
  assign n15524 = ~n15830 | ~n15522;
  assign n15528 = ~n15524 | ~n15523;
  assign n15526 = ~n15818 | ~P1_ADDR_REG_4__SCAN_IN;
  assign n15525 = ~n12098 | ~n16213;
  assign n15527 = ~n15526 | ~n15525;
  assign n15537 = ~n15528 & ~n15527;
  assign n15542 = n16213 | P1_REG1_REG_4__SCAN_IN;
  assign n15529 = ~n16213 | ~P1_REG1_REG_4__SCAN_IN;
  assign n15540 = ~n15542 | ~n15529;
  assign n15532 = ~n16219 | ~P1_REG1_REG_3__SCAN_IN;
  assign n15533 = n15540 ^ n15541;
  assign n15534 = ~n15653 & ~n15533;
  assign n15536 = ~n15535 & ~n15534;
  assign P1_U3245 = ~n15537 | ~n15536;
  assign n15538 = ~n15818 | ~P1_ADDR_REG_5__SCAN_IN;
  assign n15549 = ~n15539 | ~n15538;
  assign n15559 = n15543 & n15542;
  assign n15544 = ~P1_REG1_REG_5__SCAN_IN;
  assign n15558 = ~n16207 ^ n15544;
  assign n15545 = n15559 ^ n15558;
  assign n15547 = ~n15816 | ~n15545;
  assign n15546 = ~n12098 | ~n16207;
  assign n15548 = ~n15547 | ~n15546;
  assign n15555 = ~n15549 & ~n15548;
  assign n15570 = ~n15551 | ~n15550;
  assign n15552 = ~P1_REG2_REG_5__SCAN_IN;
  assign n15569 = ~n16207 ^ n15552;
  assign n15553 = ~n15570 ^ n15569;
  assign n15554 = ~n15830 | ~n15553;
  assign P1_U3246 = ~n15555 | ~n15554;
  assign n15647 = ~n12098;
  assign n16202 = ~n15588;
  assign n15557 = ~n15647 & ~n16202;
  assign n15580 = ~n15557 & ~n15556;
  assign n15561 = ~n15559 | ~n15558;
  assign n15560 = ~n16207 | ~P1_REG1_REG_5__SCAN_IN;
  assign n15564 = ~n15561 | ~n15560;
  assign n15581 = n15588 | P1_REG1_REG_6__SCAN_IN;
  assign n15562 = ~n15588 | ~P1_REG1_REG_6__SCAN_IN;
  assign n15563 = ~n15581 | ~n15562;
  assign n15565 = ~n15564 | ~n15563;
  assign n15566 = ~n15582 | ~n15565;
  assign n15568 = ~n15816 | ~n15566;
  assign n15567 = ~n15818 | ~P1_ADDR_REG_6__SCAN_IN;
  assign n15578 = ~n15568 | ~n15567;
  assign n15572 = ~n15570 | ~n15569;
  assign n15571 = n16207 | P1_REG2_REG_5__SCAN_IN;
  assign n15574 = ~n15572 | ~n15571;
  assign n15573 = ~n15588 ^ P1_REG2_REG_6__SCAN_IN;
  assign n15576 = n15574 & n15573;
  assign n15590 = n15574 | n15573;
  assign n15575 = ~n15830 | ~n15590;
  assign n15577 = ~n15576 & ~n15575;
  assign n15579 = ~n15578 & ~n15577;
  assign P1_U3247 = ~n15580 | ~n15579;
  assign n15603 = n16196 | P1_REG1_REG_7__SCAN_IN;
  assign n15583 = ~n16196 | ~P1_REG1_REG_7__SCAN_IN;
  assign n15584 = n15603 & n15583;
  assign n15586 = n15585 | n15584;
  assign n15587 = ~n15586 | ~n15604;
  assign n15602 = ~n15816 | ~n15587;
  assign n15589 = ~n15588 | ~P1_REG2_REG_6__SCAN_IN;
  assign n15592 = n15590 & n15589;
  assign n15911 = ~P1_REG2_REG_7__SCAN_IN;
  assign n15591 = ~n16196 ^ n15911;
  assign n15593 = n15592 | n15591;
  assign n15613 = ~n15592 | ~n15591;
  assign n15594 = ~n15593 | ~n15613;
  assign n15596 = ~n15830 | ~n15594;
  assign n15600 = ~n15596 | ~n15595;
  assign n15598 = ~n15818 | ~P1_ADDR_REG_7__SCAN_IN;
  assign n15597 = ~n12098 | ~n16196;
  assign n15599 = ~n15598 | ~n15597;
  assign n15601 = ~n15600 & ~n15599;
  assign P1_U3248 = ~n15602 | ~n15601;
  assign n15625 = n16190 | P1_REG1_REG_8__SCAN_IN;
  assign n15605 = ~n16190 | ~P1_REG1_REG_8__SCAN_IN;
  assign n15606 = n15625 & n15605;
  assign n15608 = n15607 | n15606;
  assign n15626 = ~n15607 | ~n15606;
  assign n15609 = ~n15608 | ~n15626;
  assign n15624 = ~n15816 | ~n15609;
  assign n15610 = ~n15818 | ~P1_ADDR_REG_8__SCAN_IN;
  assign n15622 = ~n15611 | ~n15610;
  assign n15612 = n16196 | P1_REG2_REG_7__SCAN_IN;
  assign n15616 = ~n15613 | ~n15612;
  assign n15636 = n16190 | P1_REG2_REG_8__SCAN_IN;
  assign n15614 = ~n16190 | ~P1_REG2_REG_8__SCAN_IN;
  assign n15615 = n15636 & n15614;
  assign n15637 = ~n15616 | ~n15615;
  assign n15617 = n15616 | n15615;
  assign n15618 = ~n15637 | ~n15617;
  assign n15620 = ~n15618 | ~n15830;
  assign n15619 = ~n12098 | ~n16190;
  assign n15621 = ~n15620 | ~n15619;
  assign n15623 = ~n15622 & ~n15621;
  assign P1_U3249 = ~n15624 | ~n15623;
  assign n15630 = n15626 & n15625;
  assign n16185 = ~n15657;
  assign n15627 = ~P1_REG1_REG_9__SCAN_IN;
  assign n15650 = ~n16185 | ~n15627;
  assign n15628 = ~n15657 | ~P1_REG1_REG_9__SCAN_IN;
  assign n15629 = ~n15650 | ~n15628;
  assign n15652 = ~n15630 & ~n15629;
  assign n15632 = ~n15652;
  assign n15631 = ~n15630 | ~n15629;
  assign n15633 = ~n15632 | ~n15631;
  assign n15644 = ~n15633 | ~n15816;
  assign n15634 = ~n15818 | ~P1_ADDR_REG_9__SCAN_IN;
  assign n15642 = ~n15635 | ~n15634;
  assign n15655 = ~n15657 ^ P1_REG2_REG_9__SCAN_IN;
  assign n15656 = ~n15637 | ~n15636;
  assign n15638 = n15655 ^ n15656;
  assign n15640 = ~n15638 | ~n15830;
  assign n15639 = ~n12098 | ~n15657;
  assign n15641 = ~n15640 | ~n15639;
  assign n15643 = ~n15642 & ~n15641;
  assign P1_U3250 = ~n15644 | ~n15643;
  assign n15645 = ~n15818 | ~P1_ADDR_REG_10__SCAN_IN;
  assign n15649 = ~n15646 | ~n15645;
  assign n16179 = ~n15672;
  assign n15648 = ~n15647 & ~n16179;
  assign n15667 = ~n15649 & ~n15648;
  assign n15668 = ~P1_REG1_REG_10__SCAN_IN ^ n15672;
  assign n15651 = ~n15650;
  assign n15669 = ~n15652 & ~n15651;
  assign n15654 = n15668 ^ n15669;
  assign n15665 = ~n15654 & ~n15653;
  assign n15660 = P1_REG2_REG_10__SCAN_IN ^ n15672;
  assign n15659 = n15656 | n15655;
  assign n15658 = ~n15657 | ~P1_REG2_REG_9__SCAN_IN;
  assign n15661 = ~n15659 | ~n15658;
  assign n15663 = ~n15660 & ~n15661;
  assign n15673 = ~n15661 | ~n15660;
  assign n15662 = ~n15673 | ~n15830;
  assign n15664 = ~n15663 & ~n15662;
  assign n15666 = ~n15665 & ~n15664;
  assign P1_U3251 = ~n15667 | ~n15666;
  assign n15685 = ~P1_REG1_REG_11__SCAN_IN ^ n16173;
  assign n15670 = ~n15672 & ~P1_REG1_REG_10__SCAN_IN;
  assign n15671 = ~n15685 ^ n15686;
  assign n15684 = ~n15671 | ~n15816;
  assign n15674 = ~n15672 | ~P1_REG2_REG_10__SCAN_IN;
  assign n15690 = ~n15674 | ~n15673;
  assign n15691 = n16173 ^ n15675;
  assign n15676 = ~n15690 ^ n15691;
  assign n15678 = ~n15676 | ~n15830;
  assign n15682 = ~n15678 | ~n15677;
  assign n15680 = ~P1_ADDR_REG_11__SCAN_IN | ~n15818;
  assign n15679 = ~n12098 | ~n16173;
  assign n15681 = ~n15680 | ~n15679;
  assign n15683 = ~n15682 & ~n15681;
  assign P1_U3252 = ~n15684 | ~n15683;
  assign n15703 = ~P1_REG1_REG_12__SCAN_IN ^ n16167;
  assign n15687 = ~n15703 ^ n9011;
  assign n15700 = ~n15687 | ~n15816;
  assign n15688 = ~n15818 | ~P1_ADDR_REG_12__SCAN_IN;
  assign n15698 = ~n15689 | ~n15688;
  assign n15693 = ~n16173 & ~P1_REG2_REG_11__SCAN_IN;
  assign n15692 = ~n15691 & ~n15690;
  assign n15712 = ~n15693 & ~n15692;
  assign n15711 = P1_REG2_REG_12__SCAN_IN ^ n16167;
  assign n15694 = n15712 ^ n15711;
  assign n15696 = ~n15694 | ~n15830;
  assign n15695 = ~n12098 | ~n16167;
  assign n15697 = ~n15696 | ~n15695;
  assign n15699 = ~n15698 & ~n15697;
  assign P1_U3253 = ~n15700 | ~n15699;
  assign n15701 = ~n12098 | ~n16161;
  assign n15710 = ~n15702 | ~n15701;
  assign n15718 = ~P1_REG1_REG_13__SCAN_IN ^ n16161;
  assign n15705 = ~n16167 & ~P1_REG1_REG_12__SCAN_IN;
  assign n15704 = ~n9011 & ~n15703;
  assign n15706 = ~n15718 ^ n15719;
  assign n15708 = ~n15706 | ~n15816;
  assign n15707 = ~n15818 | ~P1_ADDR_REG_13__SCAN_IN;
  assign n15709 = ~n15708 | ~n15707;
  assign n15717 = ~n15710 & ~n15709;
  assign n15724 = P1_REG2_REG_13__SCAN_IN ^ n16161;
  assign n15714 = ~n16167 | ~P1_REG2_REG_12__SCAN_IN;
  assign n15713 = ~n15712 | ~n15711;
  assign n15723 = ~n15714 | ~n15713;
  assign n15715 = n15724 ^ n15723;
  assign n15716 = ~n15715 | ~n15830;
  assign P1_U3254 = ~n15717 | ~n15716;
  assign n15747 = ~P1_REG1_REG_14__SCAN_IN ^ n16155;
  assign n15720 = ~n15747 ^ n15748;
  assign n15734 = ~n15720 | ~n15816;
  assign n15721 = ~n15818 | ~P1_ADDR_REG_14__SCAN_IN;
  assign n15732 = ~n15722 | ~n15721;
  assign n15726 = ~n16161 | ~P1_REG2_REG_13__SCAN_IN;
  assign n15725 = ~n15724 | ~n15723;
  assign n15737 = ~n15726 | ~n15725;
  assign n15740 = ~n16155 | ~P1_REG2_REG_14__SCAN_IN;
  assign n15738 = n16155 | P1_REG2_REG_14__SCAN_IN;
  assign n15727 = ~n15740 | ~n15738;
  assign n15728 = ~n15737 ^ n15727;
  assign n15730 = ~n15728 | ~n15830;
  assign n15729 = ~n12098 | ~n16155;
  assign n15731 = ~n15730 | ~n15729;
  assign n15733 = ~n15732 & ~n15731;
  assign P1_U3255 = ~n15734 | ~n15733;
  assign n15735 = ~n15818 | ~P1_ADDR_REG_15__SCAN_IN;
  assign n15746 = ~n15736 | ~n15735;
  assign n15739 = ~n15738 | ~n15737;
  assign n15756 = ~n15740 | ~n15739;
  assign n15757 = ~n15756 ^ n16150;
  assign n15742 = ~n15757 ^ n15741;
  assign n15744 = ~n15742 | ~n15830;
  assign n15761 = ~n16150;
  assign n15743 = ~n12098 | ~n15761;
  assign n15745 = ~n15744 | ~n15743;
  assign n15753 = ~n15746 & ~n15745;
  assign n15750 = ~n16155 & ~P1_REG1_REG_14__SCAN_IN;
  assign n15762 = ~n15750 & ~n15749;
  assign n15763 = ~n15762 ^ n16150;
  assign n15751 = P1_REG1_REG_15__SCAN_IN ^ n15763;
  assign n15752 = ~n15751 | ~n15816;
  assign P1_U3256 = ~n15753 | ~n15752;
  assign n15754 = ~n12098 | ~n16144;
  assign n15770 = ~n15755 | ~n15754;
  assign n15776 = P1_REG2_REG_16__SCAN_IN ^ n16144;
  assign n15759 = ~n15756 | ~n15761;
  assign n15758 = ~P1_REG2_REG_15__SCAN_IN | ~n15757;
  assign n15775 = ~n15759 | ~n15758;
  assign n15760 = n15776 ^ n15775;
  assign n15768 = ~n15760 | ~n15830;
  assign n15781 = P1_REG1_REG_16__SCAN_IN ^ n16144;
  assign n15765 = ~n15762 | ~n15761;
  assign n15764 = ~P1_REG1_REG_15__SCAN_IN | ~n15763;
  assign n15766 = n15781 ^ n15780;
  assign n15767 = ~n15766 | ~n15816;
  assign n15769 = ~n15768 | ~n15767;
  assign n15772 = ~n15770 & ~n15769;
  assign n15771 = ~n15818 | ~P1_ADDR_REG_16__SCAN_IN;
  assign P1_U3257 = ~n15772 | ~n15771;
  assign n15773 = ~n15818 | ~P1_ADDR_REG_17__SCAN_IN;
  assign n15787 = ~n15774 | ~n15773;
  assign n15802 = P1_REG2_REG_17__SCAN_IN ^ n16138;
  assign n15778 = ~n16144 | ~P1_REG2_REG_16__SCAN_IN;
  assign n15777 = ~n15776 | ~n15775;
  assign n15801 = ~n15778 | ~n15777;
  assign n15779 = n15802 ^ n15801;
  assign n15785 = ~n15779 | ~n15830;
  assign n15793 = P1_REG1_REG_17__SCAN_IN ^ n16138;
  assign n15782 = ~n16144 | ~P1_REG1_REG_16__SCAN_IN;
  assign n15783 = n15793 ^ n15792;
  assign n15784 = ~n15783 | ~n15816;
  assign n15786 = ~n15785 | ~n15784;
  assign n15789 = ~n15787 & ~n15786;
  assign n15788 = ~n12098 | ~n16138;
  assign P1_U3258 = ~n15789 | ~n15788;
  assign n15790 = ~n12098 | ~n16132;
  assign n15800 = ~n15791 | ~n15790;
  assign n15795 = ~n16138 | ~P1_REG1_REG_17__SCAN_IN;
  assign n15811 = ~n15795 | ~n15794;
  assign n15810 = ~P1_REG1_REG_18__SCAN_IN ^ n16132;
  assign n15796 = ~n15811 ^ n15810;
  assign n15798 = ~n15796 | ~n15816;
  assign n15797 = ~n15818 | ~P1_ADDR_REG_18__SCAN_IN;
  assign n15799 = ~n15798 | ~n15797;
  assign n15807 = ~n15800 & ~n15799;
  assign n15824 = P1_REG2_REG_18__SCAN_IN ^ n16132;
  assign n15804 = ~n16138 | ~P1_REG2_REG_17__SCAN_IN;
  assign n15803 = ~n15802 | ~n15801;
  assign n15823 = ~n15804 | ~n15803;
  assign n15805 = n15824 ^ n15823;
  assign n15806 = ~n15805 | ~n15830;
  assign P1_U3259 = ~n15807 | ~n15806;
  assign n15809 = ~n12098 | ~n16090;
  assign n15822 = ~n15809 | ~n15808;
  assign n15813 = ~n16132 & ~P1_REG1_REG_18__SCAN_IN;
  assign n15812 = ~n15811 & ~n15810;
  assign n15815 = ~n15813 & ~n15812;
  assign n15814 = P1_REG1_REG_19__SCAN_IN ^ n16125;
  assign n15817 = ~n15815 ^ n15814;
  assign n15820 = ~n15817 | ~n15816;
  assign n15819 = ~n15818 | ~P1_ADDR_REG_19__SCAN_IN;
  assign n15821 = ~n15820 | ~n15819;
  assign n15833 = ~n15822 & ~n15821;
  assign n15826 = ~n16132 | ~P1_REG2_REG_18__SCAN_IN;
  assign n15825 = ~n15824 | ~n15823;
  assign n15829 = ~n15826 | ~n15825;
  assign n15828 = ~n16125 ^ n15827;
  assign n15831 = ~n15829 ^ n15828;
  assign n15832 = ~n15831 | ~n15830;
  assign P1_U3260 = ~n15833 | ~n15832;
  assign n15835 = ~n16108 | ~n16353;
  assign n15834 = ~n16104 | ~P1_REG2_REG_9__SCAN_IN;
  assign n15838 = ~n15835 | ~n15834;
  assign n15837 = ~n16011 & ~n15836;
  assign n15858 = ~n15838 & ~n15837;
  assign n16351 = ~n15874 ^ n16353;
  assign n15843 = ~n16351 | ~n16109;
  assign n15844 = ~n15840 & ~n15839;
  assign n16356 = ~n15841 ^ n15844;
  assign n16017 = ~n16003;
  assign n15842 = ~n16356 | ~n16017;
  assign n15856 = ~n15843 | ~n15842;
  assign n15846 = ~n15845 ^ n15844;
  assign n15854 = ~n15846 & ~n16074;
  assign n15852 = ~n16356 | ~n16084;
  assign n15850 = ~n15847 & ~n16025;
  assign n15849 = ~n15848 & ~n16023;
  assign n15851 = ~n15850 & ~n15849;
  assign n15853 = ~n15852 | ~n15851;
  assign n16362 = ~n15854 & ~n15853;
  assign n15855 = ~n16104 & ~n16362;
  assign n15857 = ~n15856 & ~n15855;
  assign P1_U3282 = ~n15858 | ~n15857;
  assign n15860 = ~n16108 | ~n16334;
  assign n15859 = ~n16104 | ~P1_REG2_REG_8__SCAN_IN;
  assign n15887 = ~n15860 | ~n15859;
  assign n15862 = ~n15896 | ~n15861;
  assign n15863 = ~n15862 ^ n15869;
  assign n15873 = ~n15863 & ~n16074;
  assign n15866 = ~n15865;
  assign n15868 = ~n15867 & ~n15866;
  assign n16341 = n15869 ^ n15868;
  assign n15871 = ~n16341 | ~n16084;
  assign n15870 = ~n15929 | ~n16077;
  assign n15872 = ~n15871 | ~n15870;
  assign n16346 = ~n15873 & ~n15872;
  assign n15884 = ~n16346;
  assign n15877 = ~n15874;
  assign n15876 = ~n15875 | ~n16334;
  assign n16338 = ~n15877 | ~n15876;
  assign n15880 = ~n16338 & ~n15940;
  assign n15879 = ~n15878 & ~n16011;
  assign n15882 = ~n15880 & ~n15879;
  assign n16335 = ~n15881 | ~n16116;
  assign n15883 = ~n15882 | ~n16335;
  assign n15885 = ~n15884 & ~n15883;
  assign n15886 = ~n16104 & ~n15885;
  assign n15889 = ~n15887 & ~n15886;
  assign n15888 = ~n16341 | ~n16017;
  assign P1_U3283 = ~n15889 | ~n15888;
  assign n15892 = ~n15927 & ~n15890;
  assign n16323 = ~n15892 ^ n15891;
  assign n15909 = ~n16323 & ~n16095;
  assign n15895 = n15894 | n15893;
  assign n15897 = ~n15896 | ~n15895;
  assign n15899 = ~n15897 | ~n16055;
  assign n15898 = ~n15958 | ~n16077;
  assign n15901 = ~n15899 | ~n15898;
  assign n15900 = ~n16323 & ~n16045;
  assign n16331 = ~n15901 & ~n15900;
  assign n15902 = n16320 ^ n15938;
  assign n16327 = ~n15902 | ~n16350;
  assign n15906 = ~n16327 & ~n16090;
  assign n15904 = ~n16320 | ~n16092;
  assign n16321 = ~n15903 | ~n16116;
  assign n15905 = ~n15904 | ~n16321;
  assign n15907 = ~n15906 & ~n15905;
  assign n15908 = ~n16331 | ~n15907;
  assign n15910 = ~n15909 & ~n15908;
  assign n15913 = ~n16104 & ~n15910;
  assign n15912 = ~n16119 & ~n15911;
  assign n15916 = ~n15913 & ~n15912;
  assign n15915 = ~n16105 | ~n15914;
  assign P1_U3284 = ~n15916 | ~n15915;
  assign n15919 = ~n9155 & ~n15917;
  assign n15970 = ~n15919 & ~n15918;
  assign n15922 = ~n15970 & ~n15920;
  assign n15923 = ~n15922 & ~n15921;
  assign n15924 = ~n15923 ^ n15925;
  assign n15936 = ~n15924 | ~n16055;
  assign n15928 = ~n15926 & ~n15925;
  assign n16313 = ~n15928 & ~n15927;
  assign n15934 = ~n16313 & ~n16045;
  assign n15932 = ~n15929 | ~n16116;
  assign n15931 = ~n15930 | ~n16077;
  assign n15933 = ~n15932 | ~n15931;
  assign n15935 = ~n15934 & ~n15933;
  assign n16315 = ~n15936 | ~n15935;
  assign n15937 = ~n15956;
  assign n15939 = ~n15937 | ~n15946;
  assign n16308 = ~n15939 | ~n15938;
  assign n15941 = ~n16308 & ~n15940;
  assign n15942 = ~n16315 & ~n15941;
  assign n15950 = ~n16104 & ~n15942;
  assign n15945 = P1_REG2_REG_6__SCAN_IN & n16104;
  assign n15944 = ~n15943 & ~n16011;
  assign n15948 = ~n15945 & ~n15944;
  assign n15947 = ~n16108 | ~n15946;
  assign n15949 = ~n15948 | ~n15947;
  assign n15953 = ~n15950 & ~n15949;
  assign n15951 = ~n16313;
  assign n15952 = ~n15951 | ~n16017;
  assign P1_U3285 = ~n15953 | ~n15952;
  assign n15955 = n15954 | n15961;
  assign n15957 = ~n15955 | ~n16350;
  assign n16303 = ~n15957 & ~n15956;
  assign n15965 = ~n16303 | ~n16125;
  assign n16298 = ~n15958 | ~n16116;
  assign n15960 = ~n16105 | ~n15959;
  assign n15963 = ~n16298 | ~n15960;
  assign n15962 = ~n15961 & ~n16059;
  assign n15964 = ~n15963 & ~n15962;
  assign n15968 = ~n15965 | ~n15964;
  assign n15966 = ~n16299;
  assign n15967 = ~n15966 & ~n16095;
  assign n15977 = ~n15968 & ~n15967;
  assign n15971 = ~n15970 ^ n15969;
  assign n15976 = ~n15971 & ~n16074;
  assign n15974 = ~n16299 | ~n16084;
  assign n15973 = ~n15972 | ~n16077;
  assign n15975 = ~n15974 | ~n15973;
  assign n16305 = ~n15976 & ~n15975;
  assign n15978 = ~n15977 | ~n16305;
  assign n15980 = ~n16119 | ~n15978;
  assign n15979 = ~n16104 | ~P1_REG2_REG_5__SCAN_IN;
  assign P1_U3286 = ~n15980 | ~n15979;
  assign n16285 = ~n15981 & ~n16025;
  assign n15983 = ~n15982;
  assign n15984 = ~n16011 & ~n15983;
  assign n15994 = ~n16285 & ~n15984;
  assign n15985 = ~n9013 ^ n15989;
  assign n15993 = ~n15985 & ~n16074;
  assign n16016 = n15986 & n16020;
  assign n15988 = ~n16016 & ~n15987;
  assign n16002 = n15989 ^ n15988;
  assign n15991 = ~n16002 | ~n16084;
  assign n15990 = ~n16046 | ~n16077;
  assign n15992 = ~n15991 | ~n15990;
  assign n16293 = ~n15993 & ~n15992;
  assign n15995 = ~n15994 | ~n16293;
  assign n16001 = ~n15995 | ~n16119;
  assign n15999 = ~n15996 & ~n16283;
  assign n15997 = ~P1_REG2_REG_4__SCAN_IN;
  assign n15998 = ~n16119 & ~n15997;
  assign n16000 = ~n15999 & ~n15998;
  assign n16005 = ~n16001 | ~n16000;
  assign n16289 = ~n16002;
  assign n16004 = ~n16289 & ~n16003;
  assign n16008 = ~n16005 & ~n16004;
  assign n16286 = ~n16006 ^ n16283;
  assign n16007 = ~n16286 | ~n16109;
  assign P1_U3287 = ~n16008 | ~n16007;
  assign n16010 = ~n16108 | ~n16274;
  assign n16009 = ~n16104 | ~P1_REG2_REG_3__SCAN_IN;
  assign n16013 = ~n16010 | ~n16009;
  assign n16012 = ~P1_REG3_REG_3__SCAN_IN & ~n16011;
  assign n16036 = ~n16013 & ~n16012;
  assign n16273 = ~n16039 ^ n16014;
  assign n16019 = ~n16109 | ~n16273;
  assign n16015 = ~n15986 & ~n16020;
  assign n16271 = n16016 | n16015;
  assign n16018 = ~n16271 | ~n16017;
  assign n16034 = ~n16019 | ~n16018;
  assign n16022 = ~n16021 ^ n16020;
  assign n16032 = ~n16022 & ~n16074;
  assign n16030 = ~n16271 | ~n16084;
  assign n16024 = ~n16076;
  assign n16028 = ~n16024 & ~n16023;
  assign n16027 = ~n16026 & ~n16025;
  assign n16029 = ~n16028 & ~n16027;
  assign n16031 = ~n16030 | ~n16029;
  assign n16280 = ~n16032 & ~n16031;
  assign n16033 = ~n16104 & ~n16280;
  assign n16035 = ~n16034 & ~n16033;
  assign P1_U3288 = ~n16036 | ~n16035;
  assign n16038 = n16037 | n16261;
  assign n16260 = ~n16039 | ~n16038;
  assign n16067 = ~n16040 & ~n16260;
  assign n16044 = ~n16041;
  assign n16043 = ~n16042 & ~n16051;
  assign n16264 = ~n16044 & ~n16043;
  assign n16050 = ~n16264 & ~n16045;
  assign n16048 = ~n16046 | ~n16116;
  assign n16047 = ~n11249 | ~n16077;
  assign n16049 = ~n16048 | ~n16047;
  assign n16058 = ~n16050 & ~n16049;
  assign n16052 = ~n13133;
  assign n16054 = ~n16052 | ~n16051;
  assign n16056 = ~n16054 | ~n16053;
  assign n16057 = ~n16056 | ~n16055;
  assign n16266 = ~n16058 | ~n16057;
  assign n16060 = ~n16261 & ~n16059;
  assign n16062 = ~n16266 & ~n16060;
  assign n16061 = ~n16105 | ~P1_REG3_REG_2__SCAN_IN;
  assign n16064 = ~n16062 | ~n16061;
  assign n16063 = ~n16264 & ~n16095;
  assign n16065 = ~n16064 & ~n16063;
  assign n16066 = ~n16104 & ~n16065;
  assign n16069 = ~n16067 & ~n16066;
  assign n16068 = ~P1_REG2_REG_2__SCAN_IN | ~n16104;
  assign P1_U3289 = ~n16069 | ~n16068;
  assign n16073 = ~n16070;
  assign n16072 = ~n12800 & ~n16071;
  assign n16075 = ~n16073 & ~n16072;
  assign n16082 = ~n16075 & ~n16074;
  assign n16080 = ~n16076 | ~n16116;
  assign n16079 = ~n16078 | ~n16077;
  assign n16081 = ~n16080 | ~n16079;
  assign n16086 = ~n16082 & ~n16081;
  assign n16250 = n12800 ^ n16083;
  assign n16085 = ~n16250 | ~n16084;
  assign n16255 = ~n16086 | ~n16085;
  assign n16089 = ~n16088 ^ n9487;
  assign n16256 = ~n16089 | ~n16350;
  assign n16091 = ~n16256 & ~n16090;
  assign n16100 = ~n16255 & ~n16091;
  assign n16094 = ~n16105 | ~P1_REG3_REG_1__SCAN_IN;
  assign n16093 = ~n16251 | ~n16092;
  assign n16098 = ~n16094 | ~n16093;
  assign n16096 = ~n16250;
  assign n16097 = ~n16096 & ~n16095;
  assign n16099 = ~n16098 & ~n16097;
  assign n16101 = ~n16100 | ~n16099;
  assign n16103 = ~n16119 | ~n16101;
  assign n16102 = ~n16104 | ~P1_REG2_REG_1__SCAN_IN;
  assign P1_U3290 = ~n16103 | ~n16102;
  assign n16107 = ~n16104 | ~P1_REG2_REG_0__SCAN_IN;
  assign n16106 = ~P1_REG3_REG_0__SCAN_IN | ~n16105;
  assign n16112 = ~n16107 | ~n16106;
  assign n16110 = ~n16109 & ~n16108;
  assign n16111 = ~n16110 & ~n16244;
  assign n16121 = ~n16112 & ~n16111;
  assign n16114 = ~n16113 | ~n16245;
  assign n16118 = n16115 | n16114;
  assign n16117 = ~n11249 | ~n16116;
  assign n16247 = ~n16118 | ~n16117;
  assign n16120 = ~n16119 | ~n16247;
  assign P1_U3291 = ~n16121 | ~n16120;
  assign n16123 = ~n16122;
  assign P1_U3292 = P1_D_REG_31__SCAN_IN & n16233;
  assign P1_U3293 = P1_D_REG_30__SCAN_IN & n16233;
  assign P1_U3294 = P1_D_REG_29__SCAN_IN & n16233;
  assign P1_U3295 = P1_D_REG_28__SCAN_IN & n16233;
  assign P1_U3296 = P1_D_REG_27__SCAN_IN & n16233;
  assign P1_U3297 = P1_D_REG_26__SCAN_IN & n16233;
  assign P1_U3298 = P1_D_REG_25__SCAN_IN & n16233;
  assign P1_U3299 = P1_D_REG_24__SCAN_IN & n16233;
  assign P1_U3300 = P1_D_REG_23__SCAN_IN & n16233;
  assign P1_U3301 = P1_D_REG_22__SCAN_IN & n16233;
  assign P1_U3302 = P1_D_REG_21__SCAN_IN & n16233;
  assign P1_U3303 = P1_D_REG_20__SCAN_IN & n16233;
  assign P1_U3304 = P1_D_REG_19__SCAN_IN & n16233;
  assign P1_U3305 = P1_D_REG_18__SCAN_IN & n16233;
  assign P1_U3306 = P1_D_REG_17__SCAN_IN & n16233;
  assign P1_U3307 = P1_D_REG_16__SCAN_IN & n16233;
  assign P1_U3308 = P1_D_REG_15__SCAN_IN & n16233;
  assign P1_U3309 = P1_D_REG_14__SCAN_IN & n16233;
  assign P1_U3310 = P1_D_REG_13__SCAN_IN & n16233;
  assign P1_U3311 = P1_D_REG_12__SCAN_IN & n16233;
  assign P1_U3312 = P1_D_REG_11__SCAN_IN & n16233;
  assign P1_U3313 = P1_D_REG_10__SCAN_IN & n16233;
  assign P1_U3314 = P1_D_REG_9__SCAN_IN & n16233;
  assign P1_U3315 = P1_D_REG_8__SCAN_IN & n16233;
  assign P1_U3316 = P1_D_REG_7__SCAN_IN & n16233;
  assign P1_U3317 = P1_D_REG_6__SCAN_IN & n16233;
  assign P1_U3318 = P1_D_REG_5__SCAN_IN & n16233;
  assign P1_U3319 = P1_D_REG_4__SCAN_IN & n16233;
  assign P1_U3320 = P1_D_REG_3__SCAN_IN & n16233;
  assign P1_U3321 = P1_D_REG_2__SCAN_IN & n16233;
  assign n17226 = ~n16124;
  assign n16127 = ~n17226 & ~n16225;
  assign n16126 = ~n16125 & ~P1_U3084;
  assign n16130 = ~n16127 & ~n16126;
  assign n16230 = ~n16128;
  assign n16129 = ~n16230 | ~P2_DATAO_REG_19__SCAN_IN;
  assign P1_U3334 = ~n16130 | ~n16129;
  assign n17232 = ~n16131;
  assign n16135 = ~n17232 & ~n16225;
  assign n16133 = ~n16132;
  assign n16134 = ~n16133 & ~P1_U3084;
  assign n16137 = ~n16135 & ~n16134;
  assign n16136 = ~n16230 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P1_U3335 = ~n16137 | ~n16136;
  assign n16141 = ~n17238 & ~n16225;
  assign n16139 = ~n16138;
  assign n16140 = ~n16139 & ~P1_U3084;
  assign n16143 = ~n16141 & ~n16140;
  assign n16142 = ~n16230 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P1_U3336 = ~n16143 | ~n16142;
  assign n16147 = ~n17245 & ~n16225;
  assign n16145 = ~n16144;
  assign n16146 = ~n16145 & ~P1_U3084;
  assign n16149 = ~n16147 & ~n16146;
  assign n16148 = ~n16230 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P1_U3337 = ~n16149 | ~n16148;
  assign n16152 = ~n17252 & ~n16225;
  assign n16151 = ~n16150 & ~P1_U3084;
  assign n16154 = ~n16152 & ~n16151;
  assign n16153 = ~n16230 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P1_U3338 = ~n16154 | ~n16153;
  assign n16158 = ~n17258 & ~n16225;
  assign n16156 = ~n16155;
  assign n16157 = ~n16156 & ~P1_U3084;
  assign n16160 = ~n16158 & ~n16157;
  assign n16159 = ~n16230 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P1_U3339 = ~n16160 | ~n16159;
  assign n16164 = ~n17265 & ~n16225;
  assign n16162 = ~n16161;
  assign n16163 = ~n16162 & ~P1_U3084;
  assign n16166 = ~n16164 & ~n16163;
  assign n16165 = ~n16230 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P1_U3340 = ~n16166 | ~n16165;
  assign n16170 = ~n17271 & ~n16225;
  assign n16168 = ~n16167;
  assign n16169 = ~n16168 & ~P1_U3084;
  assign n16172 = ~n16170 & ~n16169;
  assign n16171 = ~n16230 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P1_U3341 = ~n16172 | ~n16171;
  assign n16176 = ~n17278 & ~n16225;
  assign n16174 = ~n16173;
  assign n16175 = ~n16174 & ~P1_U3084;
  assign n16178 = ~n16176 & ~n16175;
  assign n16177 = ~n16230 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P1_U3342 = ~n16178 | ~n16177;
  assign n16181 = ~n17284 & ~n16225;
  assign n16180 = ~n16179 & ~P1_U3084;
  assign n16183 = ~n16181 & ~n16180;
  assign n16182 = ~n16230 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P1_U3343 = ~n16183 | ~n16182;
  assign n16187 = ~n17291 & ~n16225;
  assign n16186 = ~n16185 & ~P1_U3084;
  assign n16189 = ~n16187 & ~n16186;
  assign n16188 = ~n16230 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P1_U3344 = ~n16189 | ~n16188;
  assign n16193 = ~n17298 & ~n16225;
  assign n16191 = ~n16190;
  assign n16192 = ~n16191 & ~P1_U3084;
  assign n16195 = ~n16193 & ~n16192;
  assign n16194 = ~n16230 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P1_U3345 = ~n16195 | ~n16194;
  assign n16199 = ~n17305 & ~n16225;
  assign n16197 = ~n16196;
  assign n16198 = ~n16197 & ~P1_U3084;
  assign n16201 = ~n16199 & ~n16198;
  assign n16200 = ~n16230 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P1_U3346 = ~n16201 | ~n16200;
  assign n16204 = ~n17312 & ~n16225;
  assign n16203 = ~n16202 & ~P1_U3084;
  assign n16206 = ~n16204 & ~n16203;
  assign n16205 = ~n16230 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P1_U3347 = ~n16206 | ~n16205;
  assign n16210 = ~n17319 & ~n16225;
  assign n16208 = ~n16207;
  assign n16209 = ~n16208 & ~P1_U3084;
  assign n16212 = ~n16210 & ~n16209;
  assign n16211 = ~n16230 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P1_U3348 = ~n16212 | ~n16211;
  assign n16216 = ~n17326 & ~n16225;
  assign n16214 = ~n16213;
  assign n16215 = ~n16214 & ~P1_U3084;
  assign n16218 = ~n16216 & ~n16215;
  assign n16217 = ~n16230 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P1_U3349 = ~n16218 | ~n16217;
  assign n16222 = ~n17333 & ~n16225;
  assign n16220 = ~n16219;
  assign n16221 = ~n16220 & ~P1_U3084;
  assign n16224 = ~n16222 & ~n16221;
  assign n16223 = ~n16230 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P1_U3350 = ~n16224 | ~n16223;
  assign n16229 = ~n17341 & ~n16225;
  assign n16227 = ~n16226;
  assign n16228 = ~n16227 & ~P1_U3084;
  assign n16232 = ~n16229 & ~n16228;
  assign n16231 = ~n16230 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P1_U3352 = ~n16232 | ~n16231;
  assign n16237 = ~P1_D_REG_0__SCAN_IN | ~n16233;
  assign n16235 = ~n16233;
  assign n16236 = ~n16235 | ~n16234;
  assign P1_U3440 = ~n16237 | ~n16236;
  assign n16243 = ~P1_D_REG_1__SCAN_IN | ~n16238;
  assign n16240 = ~n16239;
  assign n16242 = ~n16241 | ~n16240;
  assign P1_U3441 = ~n16243 | ~n16242;
  assign n16249 = ~P1_REG0_REG_0__SCAN_IN | ~n16349;
  assign n16246 = ~n16245 & ~n16244;
  assign n16366 = n16247 | n16246;
  assign n16248 = ~n16363 | ~n16366;
  assign P1_U3454 = ~n16249 | ~n16248;
  assign n16259 = ~P1_REG0_REG_1__SCAN_IN | ~n16349;
  assign n16324 = ~n16357;
  assign n16253 = ~n16250 | ~n16324;
  assign n16252 = ~n16251 | ~n16352;
  assign n16254 = ~n16253 | ~n16252;
  assign n16257 = ~n16255 & ~n16254;
  assign n16369 = ~n16257 | ~n16256;
  assign n16258 = ~n16363 | ~n16369;
  assign P1_U3457 = ~n16259 | ~n16258;
  assign n16270 = ~P1_REG0_REG_2__SCAN_IN | ~n16349;
  assign n16263 = ~n16260 & ~n16337;
  assign n16262 = ~n16261 & ~n16309;
  assign n16268 = ~n16263 & ~n16262;
  assign n16265 = ~n16264 & ~n16357;
  assign n16267 = ~n16266 & ~n16265;
  assign n16372 = ~n16268 | ~n16267;
  assign n16269 = ~n16363 | ~n16372;
  assign P1_U3460 = ~n16270 | ~n16269;
  assign n16282 = ~P1_REG0_REG_3__SCAN_IN | ~n16349;
  assign n16272 = ~n16271;
  assign n16278 = ~n16272 & ~n16357;
  assign n16276 = ~n16273 | ~n16350;
  assign n16275 = ~n16274 | ~n16352;
  assign n16277 = ~n16276 | ~n16275;
  assign n16279 = ~n16278 & ~n16277;
  assign n16375 = ~n16280 | ~n16279;
  assign n16281 = ~n16363 | ~n16375;
  assign P1_U3463 = ~n16282 | ~n16281;
  assign n16295 = ~P1_REG0_REG_4__SCAN_IN | ~n16349;
  assign n16284 = ~n16283 & ~n16309;
  assign n16288 = ~n16285 & ~n16284;
  assign n16287 = ~n16286 | ~n16350;
  assign n16291 = ~n16288 | ~n16287;
  assign n16290 = ~n16289 & ~n16357;
  assign n16292 = ~n16291 & ~n16290;
  assign n16378 = ~n16293 | ~n16292;
  assign n16294 = ~n16363 | ~n16378;
  assign P1_U3466 = ~n16295 | ~n16294;
  assign n16307 = ~P1_REG0_REG_5__SCAN_IN | ~n16349;
  assign n16297 = ~n16296 | ~n16352;
  assign n16301 = n16298 & n16297;
  assign n16300 = ~n16299 | ~n16324;
  assign n16302 = ~n16301 | ~n16300;
  assign n16304 = ~n16303 & ~n16302;
  assign n16381 = ~n16305 | ~n16304;
  assign n16306 = ~n16363 | ~n16381;
  assign P1_U3469 = ~n16307 | ~n16306;
  assign n16319 = ~P1_REG0_REG_6__SCAN_IN | ~n16349;
  assign n16312 = ~n16308 & ~n16337;
  assign n16311 = ~n16310 & ~n16309;
  assign n16317 = ~n16312 & ~n16311;
  assign n16314 = ~n16313 & ~n16357;
  assign n16316 = ~n16315 & ~n16314;
  assign n16384 = ~n16317 | ~n16316;
  assign n16318 = ~n16363 | ~n16384;
  assign P1_U3472 = ~n16319 | ~n16318;
  assign n16333 = ~P1_REG0_REG_7__SCAN_IN | ~n16349;
  assign n16322 = ~n16320 | ~n16352;
  assign n16329 = ~n16322 | ~n16321;
  assign n16325 = ~n16323;
  assign n16326 = ~n16325 | ~n16324;
  assign n16328 = ~n16327 | ~n16326;
  assign n16330 = ~n16329 & ~n16328;
  assign n16387 = ~n16331 | ~n16330;
  assign n16332 = ~n16363 | ~n16387;
  assign P1_U3475 = ~n16333 | ~n16332;
  assign n16348 = ~P1_REG0_REG_8__SCAN_IN | ~n16349;
  assign n16336 = ~n16334 | ~n16352;
  assign n16340 = n16336 & n16335;
  assign n16339 = n16338 | n16337;
  assign n16344 = ~n16340 | ~n16339;
  assign n16342 = ~n16341;
  assign n16343 = ~n16342 & ~n16357;
  assign n16345 = ~n16344 & ~n16343;
  assign n16390 = ~n16346 | ~n16345;
  assign n16347 = ~n16363 | ~n16390;
  assign P1_U3478 = ~n16348 | ~n16347;
  assign n16365 = ~P1_REG0_REG_9__SCAN_IN | ~n16349;
  assign n16355 = ~n16351 | ~n16350;
  assign n16354 = ~n16353 | ~n16352;
  assign n16360 = ~n16355 | ~n16354;
  assign n16358 = ~n16356;
  assign n16359 = ~n16358 & ~n16357;
  assign n16361 = ~n16360 & ~n16359;
  assign n16394 = ~n16362 | ~n16361;
  assign n16364 = ~n16363 | ~n16394;
  assign P1_U3481 = ~n16365 | ~n16364;
  assign n16368 = ~P1_REG1_REG_0__SCAN_IN | ~n16393;
  assign n16367 = ~n16395 | ~n16366;
  assign P1_U3523 = ~n16368 | ~n16367;
  assign n16371 = ~P1_REG1_REG_1__SCAN_IN | ~n16393;
  assign n16370 = ~n16395 | ~n16369;
  assign P1_U3524 = ~n16371 | ~n16370;
  assign n16374 = ~P1_REG1_REG_2__SCAN_IN | ~n16393;
  assign n16373 = ~n16395 | ~n16372;
  assign P1_U3525 = ~n16374 | ~n16373;
  assign n16377 = ~P1_REG1_REG_3__SCAN_IN | ~n16393;
  assign n16376 = ~n16395 | ~n16375;
  assign P1_U3526 = ~n16377 | ~n16376;
  assign n16380 = ~P1_REG1_REG_4__SCAN_IN | ~n16393;
  assign n16379 = ~n16395 | ~n16378;
  assign P1_U3527 = ~n16380 | ~n16379;
  assign n16383 = ~P1_REG1_REG_5__SCAN_IN | ~n16393;
  assign n16382 = ~n16395 | ~n16381;
  assign P1_U3528 = ~n16383 | ~n16382;
  assign n16386 = ~P1_REG1_REG_6__SCAN_IN | ~n16393;
  assign n16385 = ~n16395 | ~n16384;
  assign P1_U3529 = ~n16386 | ~n16385;
  assign n16389 = ~P1_REG1_REG_7__SCAN_IN | ~n16393;
  assign n16388 = ~n16395 | ~n16387;
  assign P1_U3530 = ~n16389 | ~n16388;
  assign n16392 = ~P1_REG1_REG_8__SCAN_IN | ~n16393;
  assign n16391 = ~n16395 | ~n16390;
  assign P1_U3531 = ~n16392 | ~n16391;
  assign n16397 = ~P1_REG1_REG_9__SCAN_IN | ~n16393;
  assign n16396 = ~n16395 | ~n16394;
  assign P1_U3532 = ~n16397 | ~n16396;
  assign n16400 = ~P1_DATAO_REG_22__SCAN_IN | ~n16425;
  assign n16399 = ~P1_U4006 | ~n16398;
  assign P1_U3577 = ~n16400 | ~n16399;
  assign n16403 = ~P1_DATAO_REG_23__SCAN_IN | ~n16425;
  assign n16402 = ~P1_U4006 | ~n16401;
  assign P1_U3578 = ~n16403 | ~n16402;
  assign n16406 = ~P1_DATAO_REG_24__SCAN_IN | ~n16425;
  assign n16405 = ~P1_U4006 | ~n16404;
  assign P1_U3579 = ~n16406 | ~n16405;
  assign n16409 = ~P1_DATAO_REG_25__SCAN_IN | ~n16425;
  assign n16408 = ~P1_U4006 | ~n16407;
  assign P1_U3580 = ~n16409 | ~n16408;
  assign n16412 = ~P1_DATAO_REG_26__SCAN_IN | ~n16425;
  assign n16411 = ~P1_U4006 | ~n16410;
  assign P1_U3581 = ~n16412 | ~n16411;
  assign n16415 = ~P1_DATAO_REG_27__SCAN_IN | ~n16425;
  assign n16414 = ~P1_U4006 | ~n16413;
  assign P1_U3582 = ~n16415 | ~n16414;
  assign n16418 = ~P1_DATAO_REG_28__SCAN_IN | ~n16425;
  assign n16417 = ~P1_U4006 | ~n16416;
  assign P1_U3583 = ~n16418 | ~n16417;
  assign n16421 = ~P1_DATAO_REG_29__SCAN_IN | ~n16425;
  assign n16420 = ~P1_U4006 | ~n16419;
  assign P1_U3584 = ~n16421 | ~n16420;
  assign n16424 = ~P1_DATAO_REG_30__SCAN_IN | ~n16425;
  assign n16423 = ~P1_U4006 | ~n16422;
  assign P1_U3585 = ~n16424 | ~n16423;
  assign n16428 = ~P1_DATAO_REG_31__SCAN_IN | ~n16425;
  assign n16427 = ~P1_U4006 | ~n16426;
  assign P1_U3586 = ~n16428 | ~n16427;
  assign P2_U3151 = ~P2_U3966 & ~n16913;
  assign n17052 = ~n17443;
  assign n16429 = ~n16617 & ~n17052;
  assign n16703 = P2_U3152 & P2_REG3_REG_7__SCAN_IN;
  assign n16441 = ~n16429 & ~n16703;
  assign n16432 = n16430 ^ n16431;
  assign n16434 = ~n16432 | ~n16575;
  assign n16433 = ~n17054 | ~n16624;
  assign n16439 = ~n16434 | ~n16433;
  assign n16437 = ~n16604 & ~n16435;
  assign n16436 = ~n16605 & ~n16516;
  assign n17050 = ~n16437 & ~n16436;
  assign n16438 = ~n17050 & ~n16608;
  assign n16440 = ~n16439 & ~n16438;
  assign P2_U3215 = ~n16441 | ~n16440;
  assign n16444 = ~n16617 & ~n16442;
  assign n16734 = ~P2_STATE_REG_SCAN_IN & ~n16443;
  assign n16455 = ~n16444 & ~n16734;
  assign n16447 = ~n16445 ^ n16446;
  assign n16453 = ~n16447 & ~n16622;
  assign n16451 = ~n16980 | ~n16624;
  assign n16449 = ~n16626 | ~n16477;
  assign n16448 = ~n16628 | ~n16505;
  assign n16995 = ~n16449 | ~n16448;
  assign n16450 = ~n16631 | ~n16995;
  assign n16452 = ~n16451 | ~n16450;
  assign n16454 = ~n16453 & ~n16452;
  assign P2_U3219 = ~n16455 | ~n16454;
  assign n16457 = ~n16617 & ~n17141;
  assign n16654 = ~P2_STATE_REG_SCAN_IN & ~n16456;
  assign n16471 = ~n16457 & ~n16654;
  assign n16461 = ~n16459 | ~n16458;
  assign n16462 = n16461 ^ n16460;
  assign n16467 = ~n16575 | ~n16462;
  assign n16465 = ~n16626 | ~n16463;
  assign n16464 = ~n16628 | ~n16517;
  assign n17154 = ~n16465 | ~n16464;
  assign n16466 = ~n16631 | ~n17154;
  assign n16469 = ~n16467 | ~n16466;
  assign n16588 = ~n16624;
  assign n16468 = ~P2_REG3_REG_3__SCAN_IN & ~n16588;
  assign n16470 = ~n16469 & ~n16468;
  assign P2_U3220 = ~n16471 | ~n16470;
  assign n17454 = ~n17041;
  assign n16473 = ~n16617 & ~n17454;
  assign n16718 = ~P2_STATE_REG_SCAN_IN & ~n16472;
  assign n16485 = ~n16473 & ~n16718;
  assign n16476 = ~n16474 ^ n16475;
  assign n16483 = ~n16476 & ~n16622;
  assign n16481 = ~n17023 | ~n16624;
  assign n16479 = ~n16626 | ~n16627;
  assign n16478 = ~n16628 | ~n16477;
  assign n17035 = ~n16479 | ~n16478;
  assign n16480 = ~n16631 | ~n17035;
  assign n16482 = ~n16481 | ~n16480;
  assign n16484 = ~n16483 & ~n16482;
  assign P2_U3223 = ~n16485 | ~n16484;
  assign n16488 = n16486 ^ n16487;
  assign n16494 = ~n16622 & ~n16488;
  assign n16492 = ~n16604 & ~n16489;
  assign n16491 = ~n16605 & ~n16490;
  assign n17378 = ~n16492 & ~n16491;
  assign n16493 = ~n17378 & ~n16608;
  assign n16499 = ~n16494 & ~n16493;
  assign n16612 = ~n16624 & ~P2_U3152;
  assign n16495 = ~P2_REG3_REG_1__SCAN_IN;
  assign n16497 = ~n16612 & ~n16495;
  assign n16496 = ~n16617 & ~n12429;
  assign n16498 = ~n16497 & ~n16496;
  assign P2_U3224 = ~n16499 | ~n16498;
  assign n16502 = ~n16501 | ~n16500;
  assign n16504 = ~n16503 ^ n16502;
  assign n16515 = ~n16504 | ~n16575;
  assign n16778 = ~P2_REG3_REG_12__SCAN_IN | ~P2_U3152;
  assign n16508 = ~n16626 | ~n16505;
  assign n16507 = ~n16628 | ~n16506;
  assign n16936 = ~n16508 | ~n16507;
  assign n16509 = ~n16631 | ~n16936;
  assign n16513 = ~n16778 | ~n16509;
  assign n16511 = ~n16569 | ~n17505;
  assign n16510 = ~n16624 | ~n16940;
  assign n16512 = ~n16511 | ~n16510;
  assign n16514 = ~n16513 & ~n16512;
  assign P2_U3226 = ~n16515 | ~n16514;
  assign n17421 = ~n16604 & ~n16516;
  assign n16518 = ~n17421;
  assign n17093 = ~n16626 | ~n16517;
  assign n16519 = ~n16518 | ~n17093;
  assign n16533 = ~n16519 | ~n16631;
  assign n16521 = ~n16569 | ~n17095;
  assign n16531 = ~n16521 | ~n16520;
  assign n16524 = ~n16522;
  assign n16525 = ~n16524 | ~n16523;
  assign n16527 = ~n16526 ^ n16525;
  assign n16529 = ~n16575 | ~n16527;
  assign n16528 = ~n17102 | ~n16624;
  assign n16530 = ~n16529 | ~n16528;
  assign n16532 = ~n16531 & ~n16530;
  assign P2_U3229 = ~n16533 | ~n16532;
  assign n16535 = ~n16617 & ~n17133;
  assign n16670 = ~P2_STATE_REG_SCAN_IN & ~n16534;
  assign n16549 = ~n16535 & ~n16670;
  assign n16539 = ~n16538 | ~n16537;
  assign n16540 = ~n16536 ^ n16539;
  assign n16545 = ~n16575 | ~n16540;
  assign n16543 = ~n16626 | ~n16541;
  assign n16542 = ~n16628 | ~n16625;
  assign n17119 = ~n16543 | ~n16542;
  assign n16544 = ~n16631 | ~n17119;
  assign n16547 = ~n16545 | ~n16544;
  assign n16546 = ~n16588 & ~n17125;
  assign n16548 = ~n16547 & ~n16546;
  assign P2_U3232 = ~n16549 | ~n16548;
  assign n16553 = ~n16552 | ~n16551;
  assign n16555 = ~n16554 ^ n16553;
  assign n16567 = ~n16555 | ~n16575;
  assign n16557 = ~n16569 | ~n17465;
  assign n16565 = ~n16557 | ~n16556;
  assign n16563 = ~n17005 | ~n16624;
  assign n16561 = ~n16626 | ~n16558;
  assign n16560 = ~n16628 | ~n16559;
  assign n17017 = ~n16561 | ~n16560;
  assign n16562 = ~n16631 | ~n17017;
  assign n16564 = ~n16563 | ~n16562;
  assign n16566 = ~n16565 & ~n16564;
  assign P2_U3233 = ~n16567 | ~n16566;
  assign n16577 = ~n16569 | ~n16568;
  assign n16572 = ~n13512 | ~n17365;
  assign n16571 = ~n12487 | ~n16570;
  assign n16573 = ~n16572 | ~n16571;
  assign n16576 = ~n16575 | ~n16574;
  assign n16579 = ~n16577 | ~n16576;
  assign n17208 = ~P2_REG3_REG_0__SCAN_IN;
  assign n16578 = ~n16612 & ~n17208;
  assign n16581 = ~n16579 & ~n16578;
  assign n17367 = n16628 & n12430;
  assign n16580 = ~n16631 | ~n17367;
  assign P2_U3234 = ~n16581 | ~n16580;
  assign n16586 = ~n16583 | ~n16582;
  assign n16585 = n16584;
  assign n16587 = n16586 ^ n16585;
  assign n16590 = ~n16587 & ~n16622;
  assign n16589 = ~n16588 & ~n16950;
  assign n16597 = ~n16590 & ~n16589;
  assign n17488 = ~n16955;
  assign n16595 = ~n16617 & ~n17488;
  assign n16760 = ~P2_REG3_REG_11__SCAN_IN | ~P2_U3152;
  assign n16970 = n16605 | n16591;
  assign n16956 = ~n16628 | ~n16592;
  assign n17489 = ~n16970 | ~n16956;
  assign n16593 = ~n16631 | ~n17489;
  assign n16594 = ~n16760 | ~n16593;
  assign n16596 = ~n16595 & ~n16594;
  assign P2_U3238 = ~n16597 | ~n16596;
  assign n16601 = ~n16600 | ~n16599;
  assign n16602 = n16598 ^ n16601;
  assign n16610 = ~n16622 & ~n16602;
  assign n16607 = ~n16604 & ~n16603;
  assign n16606 = ~n16605 & ~n10027;
  assign n17167 = ~n16607 & ~n16606;
  assign n16609 = ~n17167 & ~n16608;
  assign n16616 = ~n16610 & ~n16609;
  assign n16611 = ~P2_REG3_REG_2__SCAN_IN;
  assign n16614 = ~n16612 & ~n16611;
  assign n16613 = ~n16617 & ~n12439;
  assign n16615 = ~n16614 & ~n16613;
  assign P2_U3239 = ~n16616 | ~n16615;
  assign n16619 = ~n16617 & ~n17067;
  assign n16686 = ~P2_STATE_REG_SCAN_IN & ~n16618;
  assign n16637 = ~n16619 & ~n16686;
  assign n16623 = n16620 ^ n16621;
  assign n16635 = ~n16623 & ~n16622;
  assign n16633 = ~n17069 | ~n16624;
  assign n16630 = ~n16626 | ~n16625;
  assign n16629 = ~n16628 | ~n16627;
  assign n17084 = ~n16630 | ~n16629;
  assign n16632 = ~n16631 | ~n17084;
  assign n16634 = ~n16633 | ~n16632;
  assign n16636 = ~n16635 & ~n16634;
  assign P2_U3241 = ~n16637 | ~n16636;
  assign n16639 = n16921 & n16638;
  assign n16641 = ~n16922 & ~n16639;
  assign n16640 = ~n16911 | ~n17219;
  assign n16642 = n16641 & n16640;
  assign n16646 = ~n16642 & ~n16650;
  assign n16644 = ~P2_ADDR_REG_0__SCAN_IN | ~n16913;
  assign n16643 = ~P2_REG3_REG_0__SCAN_IN | ~P2_U3152;
  assign n16645 = ~n16644 | ~n16643;
  assign n16652 = ~n16646 & ~n16645;
  assign n16648 = ~n16921 | ~P2_REG1_REG_0__SCAN_IN;
  assign n16647 = ~n16911 | ~P2_REG2_REG_0__SCAN_IN;
  assign n16649 = ~n16648 | ~n16647;
  assign n16651 = ~n16650 | ~n16649;
  assign P2_U3245 = ~n16652 | ~n16651;
  assign n16653 = n16913 & P2_ADDR_REG_3__SCAN_IN;
  assign n16668 = ~n16654 & ~n16653;
  assign n16659 = ~n16922 | ~n17334;
  assign n16657 = n16656 ^ n16655;
  assign n16658 = ~n16921 | ~n16657;
  assign n16666 = ~n16659 | ~n16658;
  assign n16664 = ~n16661 & ~n16660;
  assign n16663 = ~n16911 | ~n16662;
  assign n16665 = ~n16664 & ~n16663;
  assign n16667 = ~n16666 & ~n16665;
  assign P2_U3248 = ~n16668 | ~n16667;
  assign n16669 = n16913 & P2_ADDR_REG_4__SCAN_IN;
  assign n16684 = ~n16670 & ~n16669;
  assign n16675 = ~n16922 | ~n17327;
  assign n16673 = n16672 ^ n16671;
  assign n16674 = ~n16921 | ~n16673;
  assign n16682 = ~n16675 | ~n16674;
  assign n16680 = ~n16677 & ~n16676;
  assign n16679 = ~n16911 | ~n16678;
  assign n16681 = ~n16680 & ~n16679;
  assign n16683 = ~n16682 & ~n16681;
  assign P2_U3249 = ~n16684 | ~n16683;
  assign n16685 = n16913 & P2_ADDR_REG_6__SCAN_IN;
  assign n16701 = ~n16686 & ~n16685;
  assign n16689 = ~n9025 & ~n16687;
  assign n16690 = n16689 ^ n16688;
  assign n16692 = ~n16911 | ~n16690;
  assign n16691 = ~n16872 | ~n17313;
  assign n16699 = ~n16692 | ~n16691;
  assign n16697 = ~n16921 | ~n16693;
  assign n16696 = ~n16695 & ~n16694;
  assign n16698 = ~n16697 & ~n16696;
  assign n16700 = ~n16699 & ~n16698;
  assign P2_U3251 = ~n16701 | ~n16700;
  assign n16702 = n16913 & P2_ADDR_REG_7__SCAN_IN;
  assign n16716 = ~n16703 & ~n16702;
  assign n16707 = ~n16922 | ~n17306;
  assign n16705 = n16704 ^ n9162;
  assign n16706 = ~n16921 | ~n16705;
  assign n16714 = ~n16707 | ~n16706;
  assign n16712 = ~n16709 & ~n16708;
  assign n16711 = ~n16911 | ~n16710;
  assign n16713 = ~n16712 & ~n16711;
  assign n16715 = ~n16714 & ~n16713;
  assign P2_U3252 = ~n16716 | ~n16715;
  assign n16717 = n16913 & P2_ADDR_REG_8__SCAN_IN;
  assign n16732 = ~n16718 & ~n16717;
  assign n16723 = ~n16922 | ~n17299;
  assign n16721 = ~n16720 ^ n16719;
  assign n16722 = ~n16921 | ~n16721;
  assign n16730 = ~n16723 | ~n16722;
  assign n16728 = ~n16725 & ~n16724;
  assign n16727 = ~n16911 | ~n16726;
  assign n16729 = ~n16728 & ~n16727;
  assign n16731 = ~n16730 & ~n16729;
  assign P2_U3253 = ~n16732 | ~n16731;
  assign n16733 = n16913 & P2_ADDR_REG_10__SCAN_IN;
  assign n16753 = ~n16734 & ~n16733;
  assign n16755 = P2_REG2_REG_10__SCAN_IN ^ n17285;
  assign n16736 = ~n16735;
  assign n16739 = ~n16737 | ~n16736;
  assign n16738 = ~n17292 | ~P2_REG2_REG_9__SCAN_IN;
  assign n16754 = ~n16739 | ~n16738;
  assign n16740 = n16755 ^ n16754;
  assign n16742 = ~n16740 | ~n16911;
  assign n16741 = ~n16872 | ~n17285;
  assign n16751 = ~n16742 | ~n16741;
  assign n16745 = ~n17292 | ~P2_REG1_REG_9__SCAN_IN;
  assign n16747 = P2_REG1_REG_10__SCAN_IN ^ n17285;
  assign n16761 = ~n16746 | ~n16747;
  assign n16749 = ~n16921 | ~n16761;
  assign n16748 = ~n16747 & ~n16746;
  assign n16750 = ~n16749 & ~n16748;
  assign n16752 = ~n16751 & ~n16750;
  assign P2_U3255 = ~n16753 | ~n16752;
  assign n16757 = ~P2_REG2_REG_10__SCAN_IN | ~n17285;
  assign n16756 = ~n16755 | ~n16754;
  assign n16781 = ~n16757 | ~n16756;
  assign n17279 = ~n16779;
  assign n16780 = P2_REG2_REG_11__SCAN_IN ^ n17279;
  assign n16758 = ~n16781 ^ n16780;
  assign n16769 = ~n16758 | ~n16911;
  assign n16759 = ~n16913 | ~P2_ADDR_REG_11__SCAN_IN;
  assign n16767 = ~n16760 | ~n16759;
  assign n16771 = ~P2_REG1_REG_11__SCAN_IN ^ n17279;
  assign n16762 = ~P2_REG1_REG_10__SCAN_IN | ~n17285;
  assign n16770 = ~n16762 | ~n16761;
  assign n16763 = n16771 ^ n16770;
  assign n16765 = ~n16763 | ~n16921;
  assign n16764 = ~n16922 | ~n16779;
  assign n16766 = ~n16765 | ~n16764;
  assign n16768 = ~n16767 & ~n16766;
  assign P2_U3256 = ~n16769 | ~n16768;
  assign n16773 = ~P2_REG1_REG_11__SCAN_IN | ~n16779;
  assign n16772 = ~n16771 | ~n16770;
  assign n16795 = ~n17272 & ~P2_REG1_REG_12__SCAN_IN;
  assign n16775 = ~n16795;
  assign n16774 = ~n17272 | ~P2_REG1_REG_12__SCAN_IN;
  assign n16793 = ~n16775 | ~n16774;
  assign n16776 = ~n16794 ^ n16793;
  assign n16792 = ~n16776 | ~n16921;
  assign n16777 = ~n16913 | ~P2_ADDR_REG_12__SCAN_IN;
  assign n16790 = ~n16778 | ~n16777;
  assign n16788 = ~n16922 | ~n17272;
  assign n16783 = ~P2_REG2_REG_11__SCAN_IN & ~n16779;
  assign n16782 = ~n16781 & ~n16780;
  assign n16800 = ~n16783 & ~n16782;
  assign n16802 = ~n17272 & ~P2_REG2_REG_12__SCAN_IN;
  assign n16785 = ~n16802;
  assign n16784 = ~n17272 | ~P2_REG2_REG_12__SCAN_IN;
  assign n16799 = ~n16785 | ~n16784;
  assign n16786 = ~n16800 ^ n16799;
  assign n16787 = ~n16911 | ~n16786;
  assign n16789 = ~n16788 | ~n16787;
  assign n16791 = ~n16790 & ~n16789;
  assign P2_U3257 = ~n16792 | ~n16791;
  assign n16810 = ~P2_REG1_REG_13__SCAN_IN ^ n16817;
  assign n16796 = ~n16810 ^ n16811;
  assign n16809 = ~n16796 | ~n16921;
  assign n16797 = ~n16913 | ~P2_ADDR_REG_13__SCAN_IN;
  assign n16807 = ~n16798 | ~n16797;
  assign n16805 = ~n16872 | ~n16817;
  assign n16801 = ~n16800 & ~n16799;
  assign n16819 = ~n16802 & ~n16801;
  assign n17266 = ~n16817;
  assign n16818 = P2_REG2_REG_13__SCAN_IN ^ n17266;
  assign n16803 = ~n16819 ^ n16818;
  assign n16804 = ~n16911 | ~n16803;
  assign n16806 = ~n16805 | ~n16804;
  assign n16808 = ~n16807 & ~n16806;
  assign P2_U3258 = ~n16809 | ~n16808;
  assign n16831 = ~P2_REG1_REG_14__SCAN_IN ^ n17259;
  assign n16813 = ~P2_REG1_REG_13__SCAN_IN & ~n16817;
  assign n16832 = ~n16813 & ~n16812;
  assign n16814 = ~n16831 ^ n16832;
  assign n16828 = ~n16814 | ~n16921;
  assign n16815 = ~n16913 | ~P2_ADDR_REG_14__SCAN_IN;
  assign n16826 = ~n16816 | ~n16815;
  assign n16824 = ~n16922 | ~n17259;
  assign n16821 = ~P2_REG2_REG_13__SCAN_IN & ~n16817;
  assign n16820 = ~n16819 & ~n16818;
  assign n16841 = ~n16821 & ~n16820;
  assign n16840 = ~P2_REG2_REG_14__SCAN_IN ^ n17259;
  assign n16822 = ~n16841 ^ n16840;
  assign n16823 = ~n16911 | ~n16822;
  assign n16825 = ~n16824 | ~n16823;
  assign n16827 = ~n16826 & ~n16825;
  assign P2_U3259 = ~n16828 | ~n16827;
  assign n16829 = ~n16913 | ~P2_ADDR_REG_15__SCAN_IN;
  assign n16839 = ~n16830 | ~n16829;
  assign n16834 = ~P2_REG1_REG_14__SCAN_IN & ~n17259;
  assign n16833 = ~n16832 & ~n16831;
  assign n16847 = ~n16834 & ~n16833;
  assign n16835 = P2_REG1_REG_15__SCAN_IN ^ n16848;
  assign n16837 = ~n16835 | ~n16921;
  assign n16836 = ~n16922 | ~n17253;
  assign n16838 = ~n16837 | ~n16836;
  assign n16846 = ~n16839 & ~n16838;
  assign n16843 = ~P2_REG2_REG_14__SCAN_IN & ~n17259;
  assign n16842 = ~n16841 & ~n16840;
  assign n16853 = ~n16843 & ~n16842;
  assign n16854 = ~n16853 ^ n17253;
  assign n16844 = ~P2_REG2_REG_15__SCAN_IN ^ n16854;
  assign n16845 = ~n16844 | ~n16911;
  assign P2_U3260 = ~n16846 | ~n16845;
  assign n16867 = ~P2_REG1_REG_16__SCAN_IN ^ n17246;
  assign n16849 = ~n17253 | ~n16847;
  assign n16850 = ~n16867 ^ n16868;
  assign n16863 = ~n16850 | ~n16921;
  assign n16851 = ~n16913 | ~P2_ADDR_REG_16__SCAN_IN;
  assign n16861 = ~n16852 | ~n16851;
  assign n16879 = P2_REG2_REG_16__SCAN_IN ^ n17246;
  assign n16856 = ~n17253 & ~n16853;
  assign n16855 = ~P2_REG2_REG_15__SCAN_IN & ~n16854;
  assign n16878 = ~n16856 & ~n16855;
  assign n16857 = n16879 ^ n16878;
  assign n16859 = ~n16857 | ~n16911;
  assign n16858 = ~n16872 | ~n17246;
  assign n16860 = ~n16859 | ~n16858;
  assign n16862 = ~n16861 & ~n16860;
  assign P2_U3261 = ~n16863 | ~n16862;
  assign n16864 = ~n16913 | ~P2_ADDR_REG_17__SCAN_IN;
  assign n16876 = ~n16865 | ~n16864;
  assign n16866 = ~P2_REG1_REG_17__SCAN_IN;
  assign n16885 = ~n17239 ^ n16866;
  assign n16870 = ~P2_REG1_REG_16__SCAN_IN & ~n17246;
  assign n16886 = ~n16870 & ~n16869;
  assign n16871 = n16885 ^ n16886;
  assign n16874 = ~n16871 | ~n16921;
  assign n16873 = ~n16872 | ~n17239;
  assign n16875 = ~n16874 | ~n16873;
  assign n16884 = ~n16876 & ~n16875;
  assign n16893 = ~n17239 ^ n16877;
  assign n16881 = ~P2_REG2_REG_16__SCAN_IN | ~n17246;
  assign n16880 = ~n16879 | ~n16878;
  assign n16892 = ~n16881 | ~n16880;
  assign n16882 = n16893 ^ n16892;
  assign n16883 = ~n16911 | ~n16882;
  assign P2_U3262 = ~n16884 | ~n16883;
  assign n16888 = ~n17239 | ~P2_REG1_REG_17__SCAN_IN;
  assign n16887 = ~n16886 | ~n16885;
  assign n16917 = ~n16888 | ~n16887;
  assign n16918 = ~P2_REG1_REG_18__SCAN_IN ^ n16916;
  assign n16889 = ~n16917 ^ n16918;
  assign n16904 = ~n16889 | ~n16921;
  assign n16890 = ~n16913 | ~P2_ADDR_REG_18__SCAN_IN;
  assign n16902 = ~n16891 | ~n16890;
  assign n16895 = ~n17239 | ~P2_REG2_REG_17__SCAN_IN;
  assign n16894 = ~n16893 | ~n16892;
  assign n16905 = ~n16895 | ~n16894;
  assign n16907 = ~P2_REG2_REG_18__SCAN_IN | ~n16916;
  assign n17233 = ~n16916;
  assign n16906 = ~n16896 | ~n17233;
  assign n16897 = ~n16907 | ~n16906;
  assign n16898 = ~n16905 ^ n16897;
  assign n16900 = ~n16898 | ~n16911;
  assign n16899 = ~n16922 | ~n16916;
  assign n16901 = ~n16900 | ~n16899;
  assign n16903 = ~n16902 & ~n16901;
  assign P2_U3263 = ~n16904 | ~n16903;
  assign n16908 = ~n16906 | ~n16905;
  assign n16909 = ~n16908 | ~n16907;
  assign n16910 = ~n16909 ^ P2_REG2_REG_19__SCAN_IN;
  assign n16912 = ~n16910 ^ n17098;
  assign n16928 = ~n16912 | ~n16911;
  assign n16914 = ~P2_ADDR_REG_19__SCAN_IN | ~n16913;
  assign n16926 = ~n16915 | ~n16914;
  assign n16920 = ~P2_REG1_REG_18__SCAN_IN & ~n16916;
  assign n16919 = ~n16918 & ~n16917;
  assign n16923 = ~n16922 | ~n17098;
  assign n16925 = ~n16924 | ~n16923;
  assign n16927 = ~n16926 & ~n16925;
  assign P2_U3264 = ~n16928 | ~n16927;
  assign n17509 = n16934 ^ n16929;
  assign n16930 = ~n17509;
  assign n16938 = ~n16930 | ~n17213;
  assign n16967 = ~n16964 & ~n16963;
  assign n16932 = ~n16931;
  assign n16933 = ~n16967 & ~n16932;
  assign n16935 = n16934 ^ n16933;
  assign n16937 = ~n16935 & ~n17362;
  assign n17513 = ~n16937 & ~n16936;
  assign n16939 = ~n16938 | ~n17513;
  assign n16949 = ~n16939 | ~n17087;
  assign n16942 = ~n17218 | ~P2_REG2_REG_12__SCAN_IN;
  assign n16941 = ~n17190 | ~n16940;
  assign n16947 = ~n16942 | ~n16941;
  assign n17503 = n16943 ^ n17505;
  assign n16945 = ~n17503 | ~n17186;
  assign n16944 = ~n17206 | ~n17505;
  assign n16946 = ~n16945 | ~n16944;
  assign n16948 = ~n16947 & ~n16946;
  assign P2_U3284 = ~n16949 | ~n16948;
  assign n16952 = ~n16950 & ~n17209;
  assign n16951 = n17218 & P2_REG2_REG_11__SCAN_IN;
  assign n16977 = ~n16952 & ~n16951;
  assign n16954 = ~n16953 ^ n17488;
  assign n17497 = ~n16954 | ~n17502;
  assign n16959 = ~n17497 & ~n17098;
  assign n16957 = ~n16955 | ~n17191;
  assign n16958 = ~n16957 | ~n16956;
  assign n16972 = n16959 | n16958;
  assign n16962 = n16960 | n16963;
  assign n17494 = ~n16962 | ~n16961;
  assign n16969 = ~n17494 & ~n17173;
  assign n16965 = ~n16964 | ~n16963;
  assign n16966 = ~n16965 | ~n17212;
  assign n16968 = ~n16967 & ~n16966;
  assign n17492 = ~n16969 & ~n16968;
  assign n16971 = ~n17492 | ~n16970;
  assign n16973 = ~n16972 & ~n16971;
  assign n16975 = ~n17218 & ~n16973;
  assign n16974 = ~n17494 & ~n17130;
  assign n16976 = ~n16975 & ~n16974;
  assign P2_U3285 = ~n16977 | ~n16976;
  assign n16979 = ~n17206 | ~n17476;
  assign n16978 = ~n17218 | ~P2_REG2_REG_10__SCAN_IN;
  assign n16982 = n16979 & n16978;
  assign n16981 = ~n16980 | ~n17190;
  assign n16988 = ~n16982 | ~n16981;
  assign n17482 = ~n16983 ^ n9059;
  assign n16986 = ~n17482 | ~n17144;
  assign n17475 = ~n16984 ^ n17476;
  assign n16985 = ~n17186 | ~n17475;
  assign n16987 = ~n16986 | ~n16985;
  assign n17000 = ~n16988 & ~n16987;
  assign n17014 = ~n16989 | ~n16990;
  assign n16992 = ~n17014 | ~n17015;
  assign n16993 = ~n16992 | ~n16991;
  assign n16994 = ~n16993 ^ n9059;
  assign n16996 = ~n16994 & ~n17362;
  assign n16998 = ~n16996 & ~n16995;
  assign n16997 = ~n17482 | ~n17150;
  assign n17480 = ~n16998 | ~n16997;
  assign n16999 = ~n17087 | ~n17480;
  assign P2_U3286 = ~n17000 | ~n16999;
  assign n17004 = ~n17068 & ~n17001;
  assign n17002 = ~P2_REG2_REG_9__SCAN_IN;
  assign n17003 = ~n17087 & ~n17002;
  assign n17007 = ~n17004 & ~n17003;
  assign n17006 = ~n17005 | ~n17190;
  assign n17013 = ~n17007 | ~n17006;
  assign n17464 = ~n17008 ^ n17465;
  assign n17011 = ~n17186 | ~n17464;
  assign n17470 = ~n17009 ^ n17015;
  assign n17010 = ~n17470 | ~n17144;
  assign n17012 = ~n17011 | ~n17010;
  assign n17022 = ~n17013 & ~n17012;
  assign n17016 = n17015 ^ n17014;
  assign n17018 = ~n17016 & ~n17362;
  assign n17020 = ~n17018 & ~n17017;
  assign n17019 = ~n17470 | ~n17150;
  assign n17469 = ~n17020 | ~n17019;
  assign n17021 = ~n17087 | ~n17469;
  assign P2_U3287 = ~n17022 | ~n17021;
  assign n17025 = ~n17218 | ~P2_REG2_REG_8__SCAN_IN;
  assign n17024 = ~n17190 | ~n17023;
  assign n17030 = ~n17025 | ~n17024;
  assign n17027 = ~n17026 | ~n17033;
  assign n17031 = n17028 & n17027;
  assign n17457 = ~n17031;
  assign n17029 = ~n17457 & ~n17130;
  assign n17047 = ~n17030 & ~n17029;
  assign n17038 = ~n17031 | ~n17150;
  assign n17034 = n17032 ^ n17033;
  assign n17036 = ~n17362 & ~n17034;
  assign n17037 = ~n17036 & ~n17035;
  assign n17459 = ~n17038 | ~n17037;
  assign n17040 = ~n17039 ^ n17041;
  assign n17456 = ~n17040 & ~n12581;
  assign n17043 = ~n17456 | ~n17227;
  assign n17042 = ~n17041 | ~n17191;
  assign n17044 = ~n17043 | ~n17042;
  assign n17045 = n17459 | n17044;
  assign n17046 = ~n17045 | ~n17087;
  assign P2_U3288 = ~n17047 | ~n17046;
  assign n17049 = n17048 ^ n17058;
  assign n17051 = ~n17049 | ~n17212;
  assign n17449 = ~n17051 | ~n17050;
  assign n17100 = ~n17191;
  assign n17053 = ~n17052 & ~n17100;
  assign n17056 = ~n17449 & ~n17053;
  assign n17055 = ~n17054 | ~n17190;
  assign n17063 = ~n17056 | ~n17055;
  assign n17447 = ~n17057 ^ n17058;
  assign n17061 = ~n17447 | ~n17213;
  assign n17442 = n17443 ^ n17059;
  assign n17060 = ~n17442 | ~n13512;
  assign n17062 = ~n17061 | ~n17060;
  assign n17064 = n17063 | n17062;
  assign n17066 = ~n17064 | ~n17087;
  assign n17065 = ~P2_REG2_REG_7__SCAN_IN | ~n17218;
  assign P2_U3289 = ~n17066 | ~n17065;
  assign n17073 = ~n17068 & ~n17067;
  assign n17071 = ~n17190 | ~n17069;
  assign n17070 = ~n17218 | ~P2_REG2_REG_6__SCAN_IN;
  assign n17072 = ~n17071 | ~n17070;
  assign n17076 = ~n17073 & ~n17072;
  assign n17431 = ~n17074 ^ n17432;
  assign n17075 = ~n17186 | ~n17431;
  assign n17079 = ~n17076 | ~n17075;
  assign n17435 = n17077 ^ n17081;
  assign n17078 = ~n17130 & ~n17435;
  assign n17090 = ~n17079 & ~n17078;
  assign n17080 = ~n17435;
  assign n17086 = ~n17080 | ~n17150;
  assign n17083 = n17082 ^ n17081;
  assign n17085 = ~n17083 & ~n17362;
  assign n17439 = ~n17085 & ~n17084;
  assign n17088 = ~n17086 | ~n17439;
  assign n17089 = ~n17088 | ~n17087;
  assign P2_U3290 = ~n17090 | ~n17089;
  assign n17092 = ~n17091 ^ n17106;
  assign n17094 = ~n17092 | ~n17212;
  assign n17424 = ~n17094 | ~n17093;
  assign n17097 = ~n17096 ^ n17095;
  assign n17427 = ~n17097 | ~n17502;
  assign n17099 = ~n17427 & ~n17098;
  assign n17110 = ~n17424 & ~n17099;
  assign n17101 = ~n17100 & ~n17419;
  assign n17104 = ~n17421 & ~n17101;
  assign n17103 = ~n17102 | ~n17190;
  assign n17108 = ~n17104 | ~n17103;
  assign n17422 = n17105 ^ n17106;
  assign n17199 = ~n17213;
  assign n17107 = ~n17422 & ~n17199;
  assign n17109 = ~n17108 & ~n17107;
  assign n17111 = ~n17110 | ~n17109;
  assign n17113 = ~n17087 | ~n17111;
  assign n17112 = ~n17218 | ~P2_REG2_REG_5__SCAN_IN;
  assign P2_U3291 = ~n17113 | ~n17112;
  assign n17412 = ~n17114 ^ n17117;
  assign n17115 = ~n17412;
  assign n17121 = ~n17115 | ~n17150;
  assign n17118 = ~n17116 ^ n17117;
  assign n17120 = ~n17118 & ~n17362;
  assign n17416 = ~n17120 & ~n17119;
  assign n17122 = ~n17121 | ~n17416;
  assign n17129 = ~n17122 | ~n17087;
  assign n17124 = ~n17206 | ~n17409;
  assign n17123 = ~n17218 | ~P2_REG2_REG_4__SCAN_IN;
  assign n17127 = ~n17124 | ~n17123;
  assign n17126 = ~n17125 & ~n17209;
  assign n17128 = ~n17127 & ~n17126;
  assign n17132 = ~n17129 | ~n17128;
  assign n17131 = ~n17130 & ~n17412;
  assign n17136 = ~n17132 & ~n17131;
  assign n17408 = ~n17134 ^ n17133;
  assign n17135 = ~n17186 | ~n17408;
  assign P2_U3292 = ~n17136 | ~n17135;
  assign n17138 = ~n17206 | ~n17399;
  assign n17137 = ~n17218 | ~P2_REG2_REG_3__SCAN_IN;
  assign n17140 = ~n17138 | ~n17137;
  assign n17139 = ~P2_REG3_REG_3__SCAN_IN & ~n17209;
  assign n17158 = ~n17140 & ~n17139;
  assign n17398 = ~n17142 ^ n17141;
  assign n17146 = ~n17186 | ~n17398;
  assign n17396 = ~n17143 ^ n17148;
  assign n17145 = ~n17144 | ~n17396;
  assign n17156 = ~n17146 | ~n17145;
  assign n17149 = n17147 ^ n17148;
  assign n17152 = ~n17149 | ~n17212;
  assign n17151 = ~n17396 | ~n17150;
  assign n17153 = ~n17152 | ~n17151;
  assign n17405 = ~n17154 & ~n17153;
  assign n17155 = ~n17218 & ~n17405;
  assign n17157 = ~n17156 & ~n17155;
  assign P2_U3293 = ~n17158 | ~n17157;
  assign n17160 = ~n17218 | ~P2_REG2_REG_2__SCAN_IN;
  assign n17159 = ~n17190 | ~P2_REG3_REG_2__SCAN_IN;
  assign n17184 = ~n17160 | ~n17159;
  assign n17162 = ~n17198;
  assign n17164 = ~n17162 | ~n17161;
  assign n17165 = ~n17164 | ~n17163;
  assign n17166 = n13204 ^ n17165;
  assign n17168 = ~n17166 | ~n17212;
  assign n17175 = ~n17168 | ~n17167;
  assign n17171 = ~n17198 | ~n17169;
  assign n17172 = ~n17171 | ~n17170;
  assign n17177 = ~n13204 ^ n17172;
  assign n17385 = ~n17177;
  assign n17174 = ~n17385 & ~n17173;
  assign n17393 = ~n17175 & ~n17174;
  assign n17181 = ~n17393;
  assign n17179 = ~n17177 | ~n17176;
  assign n17178 = ~n17191 | ~n17387;
  assign n17180 = ~n17179 | ~n17178;
  assign n17182 = ~n17181 & ~n17180;
  assign n17183 = ~n17218 & ~n17182;
  assign n17188 = ~n17184 & ~n17183;
  assign n17386 = ~n17185 ^ n17387;
  assign n17187 = ~n17186 | ~n17386;
  assign P2_U3294 = ~n17188 | ~n17187;
  assign n17381 = ~n17189 | ~n17212;
  assign n17195 = n17190 & P2_REG3_REG_1__SCAN_IN;
  assign n17372 = ~n17373 ^ n17365;
  assign n17193 = ~n13512 | ~n17372;
  assign n17192 = ~n17191 | ~n17373;
  assign n17194 = ~n17193 | ~n17192;
  assign n17196 = ~n17195 & ~n17194;
  assign n17201 = ~n17378 | ~n17196;
  assign n17376 = ~n17198 ^ n17197;
  assign n17200 = ~n17376 & ~n17199;
  assign n17202 = ~n17201 & ~n17200;
  assign n17203 = ~n17381 | ~n17202;
  assign n17205 = ~n17087 | ~n17203;
  assign n17204 = ~n17218 | ~P2_REG2_REG_1__SCAN_IN;
  assign P2_U3295 = ~n17205 | ~n17204;
  assign n17207 = ~n17206 & ~n17186;
  assign n17211 = ~n17207 & ~n17365;
  assign n17210 = ~n17209 & ~n17208;
  assign n17223 = ~n17211 & ~n17210;
  assign n17215 = ~n17213 & ~n17212;
  assign n17214 = ~n17363;
  assign n17216 = ~n17215 & ~n17214;
  assign n17217 = ~n17216 & ~n17367;
  assign n17221 = ~n17218 & ~n17217;
  assign n17220 = ~n17219 & ~n17087;
  assign n17222 = ~n17221 & ~n17220;
  assign P2_U3296 = ~n17223 | ~n17222;
  assign P2_U3297 = P2_D_REG_31__SCAN_IN & n17350;
  assign P2_U3298 = P2_D_REG_30__SCAN_IN & n17350;
  assign P2_U3299 = P2_D_REG_29__SCAN_IN & n17350;
  assign P2_U3300 = P2_D_REG_28__SCAN_IN & n17350;
  assign P2_U3301 = P2_D_REG_27__SCAN_IN & n17350;
  assign P2_U3302 = P2_D_REG_26__SCAN_IN & n17350;
  assign P2_U3303 = P2_D_REG_25__SCAN_IN & n17350;
  assign P2_U3304 = P2_D_REG_24__SCAN_IN & n17350;
  assign P2_U3305 = P2_D_REG_23__SCAN_IN & n17350;
  assign P2_U3306 = P2_D_REG_22__SCAN_IN & n17350;
  assign P2_U3307 = P2_D_REG_21__SCAN_IN & n17350;
  assign P2_U3308 = P2_D_REG_20__SCAN_IN & n17350;
  assign P2_U3309 = P2_D_REG_19__SCAN_IN & n17350;
  assign P2_U3310 = P2_D_REG_18__SCAN_IN & n17350;
  assign P2_U3311 = P2_D_REG_17__SCAN_IN & n17350;
  assign P2_U3312 = P2_D_REG_16__SCAN_IN & n17350;
  assign n17359 = ~n17350;
  assign n17353 = ~n17359;
  assign P2_U3313 = P2_D_REG_15__SCAN_IN & n17353;
  assign P2_U3314 = P2_D_REG_14__SCAN_IN & n17350;
  assign P2_U3315 = P2_D_REG_13__SCAN_IN & n17350;
  assign P2_U3316 = P2_D_REG_12__SCAN_IN & n17350;
  assign P2_U3317 = P2_D_REG_11__SCAN_IN & n17350;
  assign P2_U3318 = P2_D_REG_10__SCAN_IN & n17350;
  assign P2_U3319 = P2_D_REG_9__SCAN_IN & n17350;
  assign P2_U3320 = P2_D_REG_8__SCAN_IN & n17350;
  assign P2_U3321 = P2_D_REG_7__SCAN_IN & n17350;
  assign P2_U3322 = P2_D_REG_6__SCAN_IN & n17350;
  assign P2_U3323 = P2_D_REG_5__SCAN_IN & n17350;
  assign P2_U3324 = P2_D_REG_4__SCAN_IN & n17350;
  assign P2_U3325 = P2_D_REG_3__SCAN_IN & n17350;
  assign P2_U3326 = P2_D_REG_2__SCAN_IN & n17350;
  assign n17229 = ~n17226 & ~n17340;
  assign n17228 = ~n17227 & ~P2_U3152;
  assign n17231 = ~n17229 & ~n17228;
  assign n17230 = ~n17347 | ~P1_DATAO_REG_19__SCAN_IN;
  assign P2_U3339 = ~n17231 | ~n17230;
  assign n17235 = ~n17232 & ~n17340;
  assign n17234 = ~n17233 & ~P2_U3152;
  assign n17237 = ~n17235 & ~n17234;
  assign n17236 = ~n17347 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P2_U3340 = ~n17237 | ~n17236;
  assign n17242 = ~n17238 & ~n17340;
  assign n17240 = ~n17239;
  assign n17241 = ~n17240 & ~P2_U3152;
  assign n17244 = ~n17242 & ~n17241;
  assign n17243 = ~n17347 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P2_U3341 = ~n17244 | ~n17243;
  assign n17249 = ~n17245 & ~n17340;
  assign n17247 = ~n17246;
  assign n17248 = ~n17247 & ~P2_U3152;
  assign n17251 = ~n17249 & ~n17248;
  assign n17250 = ~n17347 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P2_U3342 = ~n17251 | ~n17250;
  assign n17255 = ~n17252 & ~n17340;
  assign n17254 = ~n9270 & ~P2_U3152;
  assign n17257 = ~n17255 & ~n17254;
  assign n17256 = ~n17347 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P2_U3343 = ~n17257 | ~n17256;
  assign n17262 = ~n17258 & ~n17340;
  assign n17260 = ~n17259;
  assign n17261 = ~n17260 & ~P2_U3152;
  assign n17264 = ~n17262 & ~n17261;
  assign n17263 = ~n17347 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P2_U3344 = ~n17264 | ~n17263;
  assign n17268 = ~n17265 & ~n17340;
  assign n17267 = ~n17266 & ~P2_U3152;
  assign n17270 = ~n17268 & ~n17267;
  assign n17269 = ~n17347 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P2_U3345 = ~n17270 | ~n17269;
  assign n17275 = ~n17271 & ~n17340;
  assign n17273 = ~n17272;
  assign n17274 = ~n17273 & ~P2_U3152;
  assign n17277 = ~n17275 & ~n17274;
  assign n17276 = ~n17347 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P2_U3346 = ~n17277 | ~n17276;
  assign n17281 = ~n17278 & ~n17340;
  assign n17280 = ~n17279 & ~P2_U3152;
  assign n17283 = ~n17281 & ~n17280;
  assign n17282 = ~n17347 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P2_U3347 = ~n17283 | ~n17282;
  assign n17288 = ~n17284 & ~n17340;
  assign n17286 = ~n17285;
  assign n17287 = ~n17286 & ~P2_U3152;
  assign n17290 = ~n17288 & ~n17287;
  assign n17289 = ~n17347 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P2_U3348 = ~n17290 | ~n17289;
  assign n17295 = ~n17291 & ~n17340;
  assign n17293 = ~n17292;
  assign n17294 = ~n17293 & ~P2_U3152;
  assign n17297 = ~n17295 & ~n17294;
  assign n17296 = ~n17347 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P2_U3349 = ~n17297 | ~n17296;
  assign n17302 = ~n17298 & ~n17340;
  assign n17300 = ~n17299;
  assign n17301 = ~n17300 & ~P2_U3152;
  assign n17304 = ~n17302 & ~n17301;
  assign n17303 = ~n17347 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P2_U3350 = ~n17304 | ~n17303;
  assign n17309 = ~n17305 & ~n17340;
  assign n17307 = ~n17306;
  assign n17308 = ~n17307 & ~P2_U3152;
  assign n17311 = ~n17309 & ~n17308;
  assign n17310 = ~n17347 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P2_U3351 = ~n17311 | ~n17310;
  assign n17316 = ~n17312 & ~n17340;
  assign n17314 = ~n17313;
  assign n17315 = ~n17314 & ~P2_U3152;
  assign n17318 = ~n17316 & ~n17315;
  assign n17317 = ~n17347 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P2_U3352 = ~n17318 | ~n17317;
  assign n17323 = ~n17319 & ~n17340;
  assign n17321 = ~n17320;
  assign n17322 = ~n17321 & ~P2_U3152;
  assign n17325 = ~n17323 & ~n17322;
  assign n17324 = ~n17347 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P2_U3353 = ~n17325 | ~n17324;
  assign n17330 = ~n17326 & ~n17340;
  assign n17328 = ~n17327;
  assign n17329 = ~n17328 & ~P2_U3152;
  assign n17332 = ~n17330 & ~n17329;
  assign n17331 = ~n17347 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P2_U3354 = ~n17332 | ~n17331;
  assign n17337 = ~n17333 & ~n17340;
  assign n17335 = ~n17334;
  assign n17336 = ~n17335 & ~P2_U3152;
  assign n17339 = ~n17337 & ~n17336;
  assign n17338 = ~n17347 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P2_U3355 = ~n17339 | ~n17338;
  assign n17346 = ~n17341 & ~n17340;
  assign n17344 = ~n17342;
  assign n17345 = ~n17344 & ~P2_U3152;
  assign n17349 = ~n17346 & ~n17345;
  assign n17348 = ~n17347 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P2_U3357 = ~n17349 | ~n17348;
  assign n17356 = ~P2_D_REG_0__SCAN_IN | ~n17350;
  assign n17354 = ~n17352 & ~n17351;
  assign n17355 = n17354 | n17353;
  assign P2_U3437 = ~n17356 | ~n17355;
  assign n17361 = n17358 & n17357;
  assign n17360 = ~P2_D_REG_1__SCAN_IN & ~n17359;
  assign P2_U3438 = ~n17361 & ~n17360;
  assign n17371 = ~P2_REG0_REG_0__SCAN_IN | ~n17501;
  assign n17508 = ~n17446;
  assign n17364 = ~n17508 | ~n17362;
  assign n17369 = ~n17364 | ~n17363;
  assign n17366 = ~n12427 & ~n17365;
  assign n17368 = ~n17367 & ~n17366;
  assign n17517 = ~n17369 | ~n17368;
  assign n17370 = ~n17514 | ~n17517;
  assign P2_U3451 = ~n17371 | ~n17370;
  assign n17384 = ~P2_REG0_REG_1__SCAN_IN | ~n17501;
  assign n17375 = ~n17372 | ~n17502;
  assign n17374 = ~n17504 | ~n17373;
  assign n17380 = ~n17375 | ~n17374;
  assign n17377 = n17376 | n17508;
  assign n17379 = ~n17378 | ~n17377;
  assign n17382 = ~n17380 & ~n17379;
  assign n17520 = ~n17382 | ~n17381;
  assign n17383 = ~n17514 | ~n17520;
  assign P2_U3454 = ~n17384 | ~n17383;
  assign n17395 = ~P2_REG0_REG_2__SCAN_IN | ~n17501;
  assign n17391 = ~n17385 & ~n17493;
  assign n17389 = ~n17386 | ~n17502;
  assign n17388 = ~n17504 | ~n17387;
  assign n17390 = ~n17389 | ~n17388;
  assign n17392 = ~n17391 & ~n17390;
  assign n17523 = ~n17393 | ~n17392;
  assign n17394 = ~n17514 | ~n17523;
  assign P2_U3457 = ~n17395 | ~n17394;
  assign n17407 = ~P2_REG0_REG_3__SCAN_IN | ~n17501;
  assign n17397 = ~n17396;
  assign n17403 = ~n17397 & ~n17493;
  assign n17401 = ~n17398 | ~n17502;
  assign n17400 = ~n17504 | ~n17399;
  assign n17402 = ~n17401 | ~n17400;
  assign n17404 = ~n17403 & ~n17402;
  assign n17526 = ~n17405 | ~n17404;
  assign n17406 = ~n17514 | ~n17526;
  assign P2_U3460 = ~n17407 | ~n17406;
  assign n17418 = ~P2_REG0_REG_4__SCAN_IN | ~n17501;
  assign n17411 = ~n17408 | ~n17502;
  assign n17410 = ~n17504 | ~n17409;
  assign n17414 = ~n17411 | ~n17410;
  assign n17413 = ~n17412 & ~n17508;
  assign n17415 = ~n17414 & ~n17413;
  assign n17529 = ~n17416 | ~n17415;
  assign n17417 = ~n17514 | ~n17529;
  assign P2_U3463 = ~n17418 | ~n17417;
  assign n17430 = ~P2_REG0_REG_5__SCAN_IN | ~n17501;
  assign n17420 = ~n17487 & ~n17419;
  assign n17426 = ~n17421 & ~n17420;
  assign n17423 = ~n17422 & ~n17508;
  assign n17425 = ~n17424 & ~n17423;
  assign n17428 = n17426 & n17425;
  assign n17532 = ~n17428 | ~n17427;
  assign n17429 = ~n17514 | ~n17532;
  assign P2_U3466 = ~n17430 | ~n17429;
  assign n17441 = ~P2_REG0_REG_6__SCAN_IN | ~n17501;
  assign n17434 = ~n17431 | ~n17502;
  assign n17433 = ~n17504 | ~n17432;
  assign n17437 = ~n17434 | ~n17433;
  assign n17436 = ~n17435 & ~n17508;
  assign n17438 = ~n17437 & ~n17436;
  assign n17535 = ~n17439 | ~n17438;
  assign n17440 = ~n17514 | ~n17535;
  assign P2_U3469 = ~n17441 | ~n17440;
  assign n17453 = ~P2_REG0_REG_7__SCAN_IN | ~n17501;
  assign n17445 = ~n17442 | ~n17502;
  assign n17444 = ~n17443 | ~n17504;
  assign n17451 = n17445 & n17444;
  assign n17448 = n17447 & n17446;
  assign n17450 = ~n17449 & ~n17448;
  assign n17538 = ~n17451 | ~n17450;
  assign n17452 = ~n17514 | ~n17538;
  assign P2_U3472 = ~n17453 | ~n17452;
  assign n17463 = ~P2_REG0_REG_8__SCAN_IN | ~n17501;
  assign n17455 = ~n17454 & ~n17487;
  assign n17461 = ~n17456 & ~n17455;
  assign n17458 = ~n17457 & ~n17493;
  assign n17460 = ~n17459 & ~n17458;
  assign n17541 = ~n17461 | ~n17460;
  assign n17462 = ~n17514 | ~n17541;
  assign P2_U3475 = ~n17463 | ~n17462;
  assign n17474 = ~P2_REG0_REG_9__SCAN_IN | ~n17501;
  assign n17467 = ~n17464 | ~n17502;
  assign n17466 = ~n17465 | ~n17504;
  assign n17468 = ~n17467 | ~n17466;
  assign n17472 = ~n17469 & ~n17468;
  assign n17471 = ~n17470 | ~n17481;
  assign n17544 = ~n17472 | ~n17471;
  assign n17473 = ~n17514 | ~n17544;
  assign P2_U3478 = ~n17474 | ~n17473;
  assign n17486 = ~P2_REG0_REG_10__SCAN_IN | ~n17501;
  assign n17478 = ~n17475 | ~n17502;
  assign n17477 = ~n17476 | ~n17504;
  assign n17479 = ~n17478 | ~n17477;
  assign n17484 = ~n17480 & ~n17479;
  assign n17483 = ~n17482 | ~n17481;
  assign n17547 = ~n17484 | ~n17483;
  assign n17485 = ~n17514 | ~n17547;
  assign P2_U3481 = ~n17486 | ~n17485;
  assign n17500 = ~P2_REG0_REG_11__SCAN_IN | ~n17501;
  assign n17490 = ~n17488 & ~n17487;
  assign n17491 = ~n17490 & ~n17489;
  assign n17496 = ~n17492 | ~n17491;
  assign n17495 = ~n17494 & ~n17493;
  assign n17498 = ~n17496 & ~n17495;
  assign n17550 = ~n17498 | ~n17497;
  assign n17499 = ~n17514 | ~n17550;
  assign P2_U3484 = ~n17500 | ~n17499;
  assign n17516 = ~P2_REG0_REG_12__SCAN_IN | ~n17501;
  assign n17507 = ~n17503 | ~n17502;
  assign n17506 = ~n17505 | ~n17504;
  assign n17511 = ~n17507 | ~n17506;
  assign n17510 = ~n17509 & ~n17508;
  assign n17512 = ~n17511 & ~n17510;
  assign n17554 = ~n17513 | ~n17512;
  assign n17515 = ~n17514 | ~n17554;
  assign P2_U3487 = ~n17516 | ~n17515;
  assign n17519 = ~P2_REG1_REG_0__SCAN_IN | ~n17553;
  assign n17518 = ~n17555 | ~n17517;
  assign P2_U3520 = ~n17519 | ~n17518;
  assign n17522 = ~P2_REG1_REG_1__SCAN_IN | ~n17553;
  assign n17521 = ~n17555 | ~n17520;
  assign P2_U3521 = ~n17522 | ~n17521;
  assign n17525 = ~P2_REG1_REG_2__SCAN_IN | ~n17553;
  assign n17524 = ~n17555 | ~n17523;
  assign P2_U3522 = ~n17525 | ~n17524;
  assign n17528 = ~P2_REG1_REG_3__SCAN_IN | ~n17553;
  assign n17527 = ~n17555 | ~n17526;
  assign P2_U3523 = ~n17528 | ~n17527;
  assign n17531 = ~P2_REG1_REG_4__SCAN_IN | ~n17553;
  assign n17530 = ~n17555 | ~n17529;
  assign P2_U3524 = ~n17531 | ~n17530;
  assign n17534 = ~P2_REG1_REG_5__SCAN_IN | ~n17553;
  assign n17533 = ~n17555 | ~n17532;
  assign P2_U3525 = ~n17534 | ~n17533;
  assign n17537 = ~P2_REG1_REG_6__SCAN_IN | ~n17553;
  assign n17536 = ~n17555 | ~n17535;
  assign P2_U3526 = ~n17537 | ~n17536;
  assign n17540 = ~P2_REG1_REG_7__SCAN_IN | ~n17553;
  assign n17539 = ~n17555 | ~n17538;
  assign P2_U3527 = ~n17540 | ~n17539;
  assign n17543 = ~P2_REG1_REG_8__SCAN_IN | ~n17553;
  assign n17542 = ~n17555 | ~n17541;
  assign P2_U3528 = ~n17543 | ~n17542;
  assign n17546 = ~P2_REG1_REG_9__SCAN_IN | ~n17553;
  assign n17545 = ~n17555 | ~n17544;
  assign P2_U3529 = ~n17546 | ~n17545;
  assign n17549 = ~P2_REG1_REG_10__SCAN_IN | ~n17553;
  assign n17548 = ~n17555 | ~n17547;
  assign P2_U3530 = ~n17549 | ~n17548;
  assign n17552 = ~P2_REG1_REG_11__SCAN_IN | ~n17553;
  assign n17551 = ~n17555 | ~n17550;
  assign P2_U3531 = ~n17552 | ~n17551;
  assign n17557 = ~P2_REG1_REG_12__SCAN_IN | ~n17553;
  assign n17556 = ~n17555 | ~n17554;
  assign P2_U3532 = ~n17557 | ~n17556;
  assign n17560 = ~P2_DATAO_REG_19__SCAN_IN | ~n17594;
  assign n17559 = ~P2_U3966 | ~n17558;
  assign P2_U3571 = ~n17560 | ~n17559;
  assign n17563 = ~P2_DATAO_REG_20__SCAN_IN | ~n17594;
  assign n17562 = ~P2_U3966 | ~n17561;
  assign P2_U3572 = ~n17563 | ~n17562;
  assign n17566 = ~P2_DATAO_REG_21__SCAN_IN | ~n17594;
  assign n17565 = ~P2_U3966 | ~n17564;
  assign P2_U3573 = ~n17566 | ~n17565;
  assign n17569 = ~P2_DATAO_REG_22__SCAN_IN | ~n17594;
  assign n17568 = ~P2_U3966 | ~n17567;
  assign P2_U3574 = ~n17569 | ~n17568;
  assign n17572 = ~P2_DATAO_REG_23__SCAN_IN | ~n17594;
  assign n17571 = ~P2_U3966 | ~n17570;
  assign P2_U3575 = ~n17572 | ~n17571;
  assign n17575 = ~P2_DATAO_REG_24__SCAN_IN | ~n17594;
  assign n17574 = ~P2_U3966 | ~n17573;
  assign P2_U3576 = ~n17575 | ~n17574;
  assign n17578 = ~P2_DATAO_REG_25__SCAN_IN | ~n17594;
  assign n17577 = ~P2_U3966 | ~n17576;
  assign P2_U3577 = ~n17578 | ~n17577;
  assign n17581 = ~P2_DATAO_REG_26__SCAN_IN | ~n17594;
  assign n17580 = ~P2_U3966 | ~n17579;
  assign P2_U3578 = ~n17581 | ~n17580;
  assign n17584 = ~P2_DATAO_REG_27__SCAN_IN | ~n17594;
  assign n17583 = ~P2_U3966 | ~n17582;
  assign P2_U3579 = ~n17584 | ~n17583;
  assign n17587 = ~P2_DATAO_REG_28__SCAN_IN | ~n17594;
  assign n17586 = ~P2_U3966 | ~n17585;
  assign P2_U3580 = ~n17587 | ~n17586;
  assign n17590 = ~P2_DATAO_REG_29__SCAN_IN | ~n17594;
  assign n17589 = ~P2_U3966 | ~n17588;
  assign P2_U3581 = ~n17590 | ~n17589;
  assign n17593 = ~P2_DATAO_REG_30__SCAN_IN | ~n17594;
  assign n17592 = ~P2_U3966 | ~n17591;
  assign P2_U3582 = ~n17593 | ~n17592;
  assign n17597 = ~P2_DATAO_REG_31__SCAN_IN | ~n17594;
  assign n17596 = ~P2_U3966 | ~n17595;
  assign P2_U3583 = ~n17597 | ~n17596;
  assign n17600 = ~n17599 & ~n17598;
  assign ADD_1071_U5 = P2_ADDR_REG_1__SCAN_IN ^ n17600;
  assign ADD_1071_U46 = P1_ADDR_REG_0__SCAN_IN ^ P2_ADDR_REG_0__SCAN_IN;
  assign ADD_1071_U47 = ~n17602 ^ n17601;
  assign ADD_1071_U48 = ~n17604 ^ n17603;
  assign ADD_1071_U49 = ~n17606 ^ n17605;
  assign ADD_1071_U50 = ~n17608 ^ n17607;
  assign ADD_1071_U51 = ~n17610 ^ n17609;
  assign ADD_1071_U52 = ~n17612 ^ n17611;
  assign ADD_1071_U53 = n17614 ^ n17613;
  assign ADD_1071_U54 = n17616 ^ n17615;
  assign ADD_1071_U55 = ~n17618 ^ n17617;
  assign n17621 = ~n17620 & ~n17619;
  assign ADD_1071_U56 = n17622 ^ n17621;
  assign n17625 = ~n17624 & ~n17623;
  assign ADD_1071_U57 = n17626 ^ n17625;
  assign n17629 = ~n17628 & ~n17627;
  assign ADD_1071_U58 = n17630 ^ n17629;
  assign n17633 = ~n17632 & ~n17631;
  assign ADD_1071_U59 = n17634 ^ n17633;
  assign n17637 = ~n17636 & ~n17635;
  assign ADD_1071_U60 = n17638 ^ n17637;
  assign n17641 = ~n17640 & ~n17639;
  assign ADD_1071_U61 = n17642 ^ n17641;
  assign n17645 = ~n17644 & ~n17643;
  assign ADD_1071_U62 = n17646 ^ n17645;
  assign n17649 = ~n17648 & ~n17647;
  assign ADD_1071_U63 = n17650 ^ n17649;
  assign n16090 = ~n16125;
endmodule


