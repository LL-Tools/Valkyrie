

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5128, n5130, n5131, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11284;

  OAI21_X1 U5192 ( .B1(n9916), .B2(n6460), .A(n9562), .ZN(n9401) );
  NAND2_X1 U5193 ( .A1(n5511), .A2(n5510), .ZN(n10480) );
  CLKBUF_X2 U5195 ( .A(n6111), .Z(n8250) );
  INV_X1 U5196 ( .A(n10228), .ZN(n10334) );
  NAND4_X1 U5197 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n10335)
         );
  INV_X4 U5198 ( .A(n6625), .ZN(n6954) );
  NOR2_X1 U5200 ( .A1(n5967), .A2(n5968), .ZN(n6092) );
  INV_X2 U5201 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  INV_X1 U5202 ( .A(n11284), .ZN(n5128) );
  INV_X2 U5203 ( .A(n5128), .ZN(P2_U3151) );
  INV_X1 U5204 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n11284) );
  NAND2_X2 U5205 ( .A1(n7574), .A2(n7639), .ZN(n10704) );
  AOI211_X1 U5206 ( .C1(n9910), .C2(n9898), .A(n9403), .B(n9402), .ZN(n9404)
         );
  NAND2_X1 U5207 ( .A1(n7199), .A2(n7579), .ZN(n7208) );
  AND2_X1 U5208 ( .A1(n5960), .A2(n8794), .ZN(n6339) );
  AND2_X1 U5209 ( .A1(n7485), .A2(n9627), .ZN(n9580) );
  NAND2_X1 U5211 ( .A1(n10334), .A2(n11043), .ZN(n7029) );
  OR2_X1 U5212 ( .A1(n6342), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6073) );
  OR2_X1 U5213 ( .A1(n6186), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U5215 ( .A1(n7172), .A2(n7474), .ZN(n7644) );
  OAI21_X1 U5216 ( .B1(n6183), .B2(n6182), .A(n6006), .ZN(n6193) );
  INV_X1 U5217 ( .A(n5988), .ZN(n6525) );
  NAND2_X1 U5218 ( .A1(n6084), .A2(n5588), .ZN(n8390) );
  AOI21_X1 U5219 ( .B1(n5486), .B2(n5488), .A(n5154), .ZN(n10294) );
  BUF_X1 U5220 ( .A(n6924), .Z(n6969) );
  OAI22_X1 U5221 ( .A1(n9225), .A2(n9224), .B1(n9223), .B2(n10284), .ZN(n9307)
         );
  XNOR2_X1 U5222 ( .A(n9314), .B(n9313), .ZN(n10617) );
  XNOR2_X1 U5223 ( .A(n6152), .B(SI_5_), .ZN(n7547) );
  INV_X1 U5224 ( .A(n9944), .ZN(n9789) );
  NOR3_X2 U5225 ( .A1(n10294), .A2(n7445), .A3(n7444), .ZN(n9651) );
  INV_X1 U5226 ( .A(n7196), .ZN(n8381) );
  AND2_X1 U5227 ( .A1(n5967), .A2(n5968), .ZN(n6119) );
  AND2_X1 U5228 ( .A1(n7579), .A2(n7201), .ZN(n7211) );
  NAND2_X2 U5230 ( .A1(n8022), .A2(n8021), .ZN(n8107) );
  NAND2_X2 U5231 ( .A1(n7759), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7830) );
  XNOR2_X2 U5232 ( .A(n6528), .B(n10688), .ZN(n6531) );
  OAI21_X2 U5233 ( .B1(n6096), .B2(n5619), .A(n5980), .ZN(n6106) );
  AOI21_X2 U5234 ( .B1(n10290), .B2(n11238), .A(n9179), .ZN(n9225) );
  OAI21_X2 U5235 ( .B1(n9117), .B2(n5537), .A(n5536), .ZN(n9817) );
  XNOR2_X2 U5236 ( .A(n5860), .B(n9130), .ZN(n9117) );
  BUF_X8 U5237 ( .A(n6119), .Z(n5130) );
  AND2_X1 U5238 ( .A1(n11247), .A2(n11246), .ZN(n5641) );
  NAND2_X1 U5239 ( .A1(n8193), .A2(n9598), .ZN(n8192) );
  NAND3_X1 U5240 ( .A1(n7709), .A2(n7217), .A3(n7687), .ZN(n7685) );
  NAND2_X1 U5241 ( .A1(n10994), .A2(n9438), .ZN(n8233) );
  INV_X1 U5242 ( .A(n9807), .ZN(n5131) );
  INV_X1 U5243 ( .A(n6103), .ZN(n6102) );
  INV_X4 U5244 ( .A(n5138), .ZN(n9633) );
  INV_X1 U5245 ( .A(n7211), .ZN(n7255) );
  INV_X1 U5246 ( .A(n8058), .ZN(n11043) );
  NAND4_X1 U5247 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n9806)
         );
  INV_X2 U5248 ( .A(n7730), .ZN(n11020) );
  CLKBUF_X1 U5249 ( .A(n9621), .Z(n5136) );
  INV_X1 U5250 ( .A(n6630), .ZN(n7581) );
  INV_X1 U5251 ( .A(n6924), .ZN(n6895) );
  INV_X4 U5252 ( .A(n10599), .ZN(n7172) );
  INV_X1 U5253 ( .A(n6531), .ZN(n5625) );
  AND3_X2 U5254 ( .A1(n6543), .A2(n6542), .A3(n6541), .ZN(n10599) );
  INV_X1 U5255 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8873) );
  AOI22_X1 U5256 ( .A1(n10040), .A2(n10039), .B1(n11158), .B2(n10038), .ZN(
        n10047) );
  OAI21_X1 U5257 ( .B1(n10294), .B2(n7445), .A(n7444), .ZN(n7446) );
  INV_X1 U5258 ( .A(n9401), .ZN(n9910) );
  OAI21_X1 U5259 ( .B1(n9714), .B2(n9716), .A(n9715), .ZN(n9771) );
  NAND2_X1 U5260 ( .A1(n6459), .A2(n9560), .ZN(n9916) );
  NAND2_X1 U5261 ( .A1(n7394), .A2(n5472), .ZN(n10197) );
  NAND2_X1 U5262 ( .A1(n5655), .A2(n5654), .ZN(n10528) );
  AND2_X1 U5263 ( .A1(n8264), .A2(n6437), .ZN(n9419) );
  NOR2_X1 U5264 ( .A1(n9826), .A2(n10101), .ZN(n9825) );
  OR2_X1 U5265 ( .A1(n9075), .A2(n5680), .ZN(n5676) );
  OR2_X1 U5266 ( .A1(n6425), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U5267 ( .A1(n7049), .A2(n7048), .ZN(n8453) );
  NAND2_X1 U5268 ( .A1(n5852), .A2(n5851), .ZN(n5857) );
  NAND2_X1 U5269 ( .A1(n5257), .A2(n5256), .ZN(n5852) );
  INV_X1 U5270 ( .A(n10541), .ZN(n10506) );
  NAND2_X1 U5271 ( .A1(n6815), .A2(n6814), .ZN(n11260) );
  OAI21_X1 U5272 ( .B1(n5687), .B2(n5144), .A(n5688), .ZN(n5686) );
  INV_X2 U5273 ( .A(n9355), .ZN(n9373) );
  AND2_X1 U5274 ( .A1(n8177), .A2(n7035), .ZN(n8116) );
  OAI21_X1 U5275 ( .B1(n6225), .B2(n5602), .A(n5599), .ZN(n6248) );
  INV_X1 U5276 ( .A(n7783), .ZN(n9355) );
  NAND2_X1 U5277 ( .A1(n5509), .A2(n6694), .ZN(n8348) );
  AND2_X1 U5278 ( .A1(n6470), .A2(n7543), .ZN(n7985) );
  NAND2_X1 U5279 ( .A1(n5774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U5280 ( .A1(n9637), .A2(n7208), .ZN(n7218) );
  INV_X4 U5281 ( .A(n9637), .ZN(n7232) );
  NOR2_X1 U5282 ( .A1(n10338), .A2(n7651), .ZN(n9254) );
  BUF_X1 U5283 ( .A(n7098), .Z(n10337) );
  NAND4_X1 U5284 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n9805)
         );
  INV_X1 U5285 ( .A(n9621), .ZN(n5135) );
  OAI211_X2 U5286 ( .C1(n7581), .C2(n10363), .A(n6659), .B(n6658), .ZN(n8058)
         );
  AND3_X1 U5287 ( .A1(n6110), .A2(n6109), .A3(n6108), .ZN(n11008) );
  OAI211_X1 U5288 ( .C1(n6100), .C2(n9661), .A(n6099), .B(n6098), .ZN(n8396)
         );
  AND3_X1 U5289 ( .A1(n6129), .A2(n6128), .A3(n6127), .ZN(n11027) );
  CLKBUF_X3 U5290 ( .A(n6092), .Z(n8257) );
  AND2_X1 U5291 ( .A1(n9273), .A2(n5968), .ZN(n6111) );
  NOR2_X1 U5292 ( .A1(n6803), .A2(n10310), .ZN(n6591) );
  NOR2_X1 U5293 ( .A1(n9056), .A2(n9025), .ZN(n7171) );
  NAND2_X1 U5294 ( .A1(n7642), .A2(n7643), .ZN(n11232) );
  AND2_X2 U5295 ( .A1(n10176), .A2(n5967), .ZN(n5160) );
  NAND2_X1 U5296 ( .A1(n7164), .A2(n7167), .ZN(n9056) );
  NAND2_X2 U5297 ( .A1(n9661), .A2(n6525), .ZN(n6104) );
  CLKBUF_X2 U5298 ( .A(n6958), .Z(n5133) );
  INV_X2 U5299 ( .A(n9661), .ZN(n6307) );
  NAND2_X2 U5300 ( .A1(n5872), .A2(n5873), .ZN(n9661) );
  MUX2_X1 U5301 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7162), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n7164) );
  XNOR2_X1 U5302 ( .A(n5762), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U5303 ( .A1(n10599), .A2(n7196), .ZN(n7642) );
  NAND2_X1 U5304 ( .A1(n5758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  AND2_X1 U5305 ( .A1(n7156), .A2(n6551), .ZN(n7196) );
  XNOR2_X1 U5306 ( .A(n7166), .B(n8895), .ZN(n9025) );
  NOR2_X1 U5307 ( .A1(n6013), .A2(n5595), .ZN(n5594) );
  NOR2_X1 U5308 ( .A1(n10936), .A2(n10935), .ZN(n10934) );
  XNOR2_X1 U5309 ( .A(n6988), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7200) );
  BUF_X1 U5310 ( .A(n6531), .Z(n9270) );
  NAND2_X1 U5311 ( .A1(n6522), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7177) );
  OR2_X1 U5312 ( .A1(n6550), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7156) );
  OR2_X1 U5313 ( .A1(n5776), .A2(n5783), .ZN(n5758) );
  NAND2_X1 U5314 ( .A1(n5790), .A2(n5147), .ZN(n5966) );
  INV_X2 U5315 ( .A(n10693), .ZN(n9271) );
  NAND2_X1 U5316 ( .A1(n7160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6987) );
  CLKBUF_X1 U5317 ( .A(n6529), .Z(n10691) );
  NOR2_X1 U5318 ( .A1(n5693), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5848) );
  OR2_X1 U5319 ( .A1(n6156), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6175) );
  NOR2_X1 U5320 ( .A1(n5647), .A2(n5653), .ZN(n6783) );
  AND4_X1 U5321 ( .A1(n6545), .A2(n6544), .A3(n8881), .A4(n8873), .ZN(n6546)
         );
  AND2_X2 U5322 ( .A1(n5597), .A2(n5596), .ZN(n5988) );
  AND3_X1 U5323 ( .A1(n5781), .A2(n5780), .A3(n5779), .ZN(n5786) );
  AND4_X1 U5324 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n5781)
         );
  MUX2_X1 U5325 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5813), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5815) );
  AND2_X1 U5326 ( .A1(n8861), .A2(n5651), .ZN(n5650) );
  AND4_X1 U5327 ( .A1(n5748), .A2(n5771), .A3(n5766), .A4(n5796), .ZN(n5780)
         );
  AND2_X1 U5328 ( .A1(n5645), .A2(n6537), .ZN(n6545) );
  NAND3_X1 U5329 ( .A1(n8173), .A2(n5598), .A3(n5975), .ZN(n5597) );
  NAND3_X1 U5330 ( .A1(n5976), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5331 ( .A1(n5387), .A2(n5386), .ZN(n5814) );
  NOR2_X1 U5332 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6544) );
  INV_X1 U5333 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5386) );
  INV_X1 U5334 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5387) );
  NOR2_X1 U5335 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5753) );
  INV_X1 U5336 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5808) );
  INV_X1 U5337 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5810) );
  INV_X1 U5338 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5833) );
  NOR2_X1 U5339 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5749) );
  NOR2_X1 U5340 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5750) );
  NOR2_X1 U5341 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6631) );
  NOR2_X1 U5342 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5751) );
  NOR2_X1 U5343 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5748) );
  INV_X1 U5344 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5976) );
  INV_X1 U5345 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5975) );
  INV_X1 U5346 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5598) );
  OR2_X1 U5347 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5783) );
  NOR2_X1 U5348 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5754) );
  INV_X1 U5349 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8173) );
  INV_X1 U5350 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8861) );
  INV_X1 U5351 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U5352 ( .B1(n6535), .B2(n6536), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6813) );
  NAND2_X2 U5353 ( .A1(n5625), .A2(n10698), .ZN(n6958) );
  AOI21_X2 U5354 ( .B1(n10445), .B2(n10455), .A(n5197), .ZN(n10446) );
  XNOR2_X2 U5355 ( .A(n5857), .B(n5391), .ZN(n8437) );
  OAI211_X2 U5356 ( .C1(n7581), .C2(n7613), .A(n6633), .B(n6632), .ZN(n8925)
         );
  NAND2_X1 U5357 ( .A1(n9637), .A2(n7208), .ZN(n5134) );
  AOI21_X2 U5358 ( .B1(n7999), .B2(n7262), .A(n7261), .ZN(n8039) );
  BUF_X4 U5359 ( .A(n7208), .Z(n5138) );
  OR2_X1 U5360 ( .A1(n10443), .A2(n6985), .ZN(n5447) );
  OR2_X1 U5361 ( .A1(n9539), .A2(n9988), .ZN(n6334) );
  NOR2_X1 U5362 ( .A1(n6444), .A2(n6443), .ZN(n9591) );
  OR2_X1 U5363 ( .A1(n9864), .A2(n9863), .ZN(n5543) );
  NOR2_X1 U5364 ( .A1(n8142), .A2(n11124), .ZN(n8141) );
  OAI21_X1 U5365 ( .B1(n5463), .B2(n5461), .A(n6825), .ZN(n5460) );
  INV_X1 U5366 ( .A(n6824), .ZN(n5461) );
  NAND2_X1 U5367 ( .A1(n5445), .A2(n5449), .ZN(n5436) );
  INV_X1 U5368 ( .A(n5369), .ZN(n5363) );
  AOI21_X1 U5369 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5366) );
  INV_X1 U5370 ( .A(n6041), .ZN(n5367) );
  INV_X1 U5371 ( .A(n5604), .ZN(n5368) );
  INV_X1 U5372 ( .A(n6006), .ZN(n5384) );
  INV_X1 U5373 ( .A(n5594), .ZN(n5593) );
  INV_X1 U5374 ( .A(n9371), .ZN(n5674) );
  NAND2_X1 U5375 ( .A1(n5340), .A2(n5338), .ZN(n9581) );
  AND2_X1 U5376 ( .A1(n5341), .A2(n5339), .ZN(n5338) );
  OR2_X1 U5377 ( .A1(n5345), .A2(n9577), .ZN(n5341) );
  OR2_X1 U5378 ( .A1(n6461), .A2(n9787), .ZN(n9365) );
  OR2_X1 U5379 ( .A1(n10072), .A2(n9978), .ZN(n9542) );
  INV_X1 U5380 ( .A(n5706), .ZN(n5705) );
  OAI21_X1 U5381 ( .B1(n10024), .B2(n5707), .A(n6302), .ZN(n5706) );
  NOR2_X1 U5382 ( .A1(n5296), .A2(n5295), .ZN(n5294) );
  INV_X1 U5383 ( .A(n5297), .ZN(n5295) );
  INV_X1 U5384 ( .A(n5703), .ZN(n5296) );
  AOI21_X1 U5385 ( .B1(n5312), .B2(n6246), .A(n5310), .ZN(n5309) );
  INV_X1 U5386 ( .A(n9514), .ZN(n5310) );
  INV_X1 U5387 ( .A(n5312), .ZN(n5311) );
  OR2_X1 U5388 ( .A1(n9152), .A2(n9796), .ZN(n5317) );
  NAND2_X1 U5389 ( .A1(n5316), .A2(n5315), .ZN(n5314) );
  INV_X1 U5390 ( .A(n8958), .ZN(n5316) );
  AND2_X1 U5391 ( .A1(n5709), .A2(n8226), .ZN(n5303) );
  NAND2_X1 U5392 ( .A1(n5205), .A2(n10998), .ZN(n5726) );
  NAND2_X1 U5393 ( .A1(n11002), .A2(n11027), .ZN(n5728) );
  INV_X1 U5394 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U5395 ( .A1(n5772), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6432) );
  AOI21_X1 U5396 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n5691), .A(
        P2_IR_REG_19__SCAN_IN), .ZN(n5690) );
  INV_X1 U5397 ( .A(n5477), .ZN(n5476) );
  OAI21_X1 U5398 ( .B1(n5480), .B2(n5478), .A(n7274), .ZN(n5477) );
  XNOR2_X1 U5399 ( .A(n7214), .B(n5138), .ZN(n7215) );
  NOR2_X1 U5400 ( .A1(n6990), .A2(n5442), .ZN(n5441) );
  INV_X1 U5401 ( .A(n7080), .ZN(n5442) );
  NAND2_X1 U5402 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  NOR2_X1 U5403 ( .A1(n10698), .A2(n6611), .ZN(n5626) );
  AND2_X1 U5404 ( .A1(n10632), .A2(n10324), .ZN(n5639) );
  INV_X1 U5405 ( .A(n7070), .ZN(n5623) );
  NAND2_X1 U5406 ( .A1(n5515), .A2(n5513), .ZN(n5372) );
  NAND2_X1 U5407 ( .A1(n10516), .A2(n9293), .ZN(n5350) );
  NOR2_X1 U5408 ( .A1(n10537), .A2(n10538), .ZN(n5518) );
  NAND2_X1 U5409 ( .A1(n10548), .A2(n10547), .ZN(n10536) );
  NOR2_X1 U5410 ( .A1(n7574), .A2(n7459), .ZN(n7737) );
  NOR2_X1 U5411 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5644) );
  NOR2_X1 U5412 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5643) );
  INV_X1 U5413 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8903) );
  OAI21_X1 U5414 ( .B1(n6369), .B2(n5612), .A(n5610), .ZN(n6399) );
  AOI21_X1 U5415 ( .B1(n5613), .B2(n5611), .A(n5254), .ZN(n5610) );
  INV_X1 U5416 ( .A(n5613), .ZN(n5612) );
  INV_X1 U5417 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8899) );
  INV_X1 U5418 ( .A(SI_21_), .ZN(n6055) );
  AND2_X1 U5419 ( .A1(n6041), .A2(n6040), .ZN(n6282) );
  INV_X1 U5420 ( .A(n6248), .ZN(n6029) );
  OAI211_X1 U5421 ( .C1(n6152), .C2(n5618), .A(n5739), .B(n5616), .ZN(n6183)
         );
  NAND2_X1 U5422 ( .A1(n5996), .A2(SI_5_), .ZN(n5618) );
  NAND2_X1 U5423 ( .A1(n5617), .A2(n5996), .ZN(n5616) );
  NOR2_X1 U5424 ( .A1(n7187), .A2(n6486), .ZN(n7523) );
  OR3_X1 U5425 ( .A1(n7485), .A2(n6466), .A3(n8387), .ZN(n7494) );
  NAND2_X1 U5426 ( .A1(n5264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  OAI211_X1 U5427 ( .C1(n7870), .C2(n5409), .A(n5407), .B(n5402), .ZN(n5400)
         );
  NOR2_X1 U5428 ( .A1(n5187), .A2(n5403), .ZN(n5402) );
  NAND2_X1 U5429 ( .A1(n5543), .A2(n5172), .ZN(n5542) );
  AND2_X1 U5430 ( .A1(n5542), .A2(n5541), .ZN(n10969) );
  INV_X1 U5431 ( .A(n10970), .ZN(n5541) );
  NAND2_X1 U5432 ( .A1(n5730), .A2(n5729), .ZN(n6367) );
  NAND2_X1 U5433 ( .A1(n9553), .A2(n9790), .ZN(n5729) );
  NAND2_X1 U5434 ( .A1(n5732), .A2(n5731), .ZN(n5730) );
  NAND2_X1 U5435 ( .A1(n10134), .A2(n9954), .ZN(n5731) );
  XNOR2_X1 U5436 ( .A(n9553), .B(n9790), .ZN(n9940) );
  AOI21_X1 U5437 ( .B1(n9977), .B2(n5570), .A(n5150), .ZN(n5569) );
  NAND2_X1 U5438 ( .A1(n5566), .A2(n5148), .ZN(n10011) );
  NAND2_X1 U5439 ( .A1(n6446), .A2(n9453), .ZN(n9277) );
  NAND2_X1 U5440 ( .A1(n8235), .A2(n5576), .ZN(n6446) );
  NOR2_X1 U5441 ( .A1(n5577), .A2(n6443), .ZN(n5576) );
  NAND2_X1 U5442 ( .A1(n9661), .A2(n7532), .ZN(n6137) );
  OR2_X1 U5443 ( .A1(n9574), .A2(n7183), .ZN(n7515) );
  INV_X1 U5444 ( .A(n6104), .ZN(n6306) );
  NAND2_X1 U5445 ( .A1(n10167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U5446 ( .A(n5320), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U5447 ( .A1(n5966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5320) );
  NOR2_X1 U5448 ( .A1(n10627), .A2(n10484), .ZN(n10461) );
  INV_X1 U5449 ( .A(n10324), .ZN(n10504) );
  OR2_X1 U5450 ( .A1(n10646), .A2(n10549), .ZN(n9308) );
  OR2_X1 U5451 ( .A1(n10664), .A2(n10571), .ZN(n9305) );
  NAND2_X1 U5452 ( .A1(n9140), .A2(n9139), .ZN(n5629) );
  OR2_X1 U5453 ( .A1(n9220), .A2(n7911), .ZN(n10507) );
  XNOR2_X1 U5454 ( .A(n6399), .B(n6398), .ZN(n9109) );
  INV_X1 U5455 ( .A(n6063), .ZN(n5358) );
  INV_X1 U5456 ( .A(n8360), .ZN(n5256) );
  INV_X1 U5457 ( .A(n8361), .ZN(n5257) );
  NAND2_X1 U5458 ( .A1(n5715), .A2(n5719), .ZN(n9653) );
  OAI21_X1 U5459 ( .B1(n5298), .B2(n11000), .A(n5300), .ZN(n10052) );
  AOI21_X1 U5460 ( .B1(n9786), .B2(n10003), .A(n5301), .ZN(n5300) );
  XNOR2_X1 U5461 ( .A(n9907), .B(n9909), .ZN(n5298) );
  NOR2_X1 U5462 ( .A1(n9932), .A2(n11001), .ZN(n5301) );
  OR2_X1 U5463 ( .A1(n6662), .A2(n6949), .ZN(n5454) );
  INV_X1 U5464 ( .A(n7910), .ZN(n6661) );
  OAI21_X1 U5465 ( .B1(n5464), .B2(n6824), .A(n5194), .ZN(n5463) );
  NOR2_X1 U5466 ( .A1(n5733), .A2(n7046), .ZN(n5464) );
  AOI21_X1 U5467 ( .B1(n5322), .B2(n9498), .A(n5321), .ZN(n9513) );
  INV_X1 U5468 ( .A(n9501), .ZN(n5321) );
  NAND2_X1 U5469 ( .A1(n5325), .A2(n5323), .ZN(n5322) );
  NAND2_X1 U5470 ( .A1(n9552), .A2(n9940), .ZN(n5329) );
  NOR2_X1 U5471 ( .A1(n5331), .A2(n5193), .ZN(n5330) );
  INV_X1 U5472 ( .A(n9956), .ZN(n5331) );
  INV_X1 U5473 ( .A(n9575), .ZN(n5345) );
  OR2_X1 U5474 ( .A1(n9803), .A2(n11063), .ZN(n9465) );
  NAND2_X1 U5475 ( .A1(n5789), .A2(n5790), .ZN(n5283) );
  AND2_X1 U5476 ( .A1(n5788), .A2(n5139), .ZN(n5789) );
  NAND2_X1 U5477 ( .A1(n6945), .A2(n6985), .ZN(n6951) );
  AOI22_X1 U5478 ( .A1(n5621), .A2(n5620), .B1(n7138), .B2(n5623), .ZN(n6944)
         );
  NOR2_X1 U5479 ( .A1(n10479), .A2(n5622), .ZN(n5621) );
  NAND2_X1 U5480 ( .A1(n5465), .A2(n6949), .ZN(n6950) );
  OAI21_X1 U5481 ( .B1(n5466), .B2(n10467), .A(n7069), .ZN(n5465) );
  INV_X1 U5482 ( .A(n5467), .ZN(n5466) );
  OAI21_X1 U5483 ( .B1(n6947), .B2(n5469), .A(n5468), .ZN(n5467) );
  INV_X1 U5484 ( .A(n6368), .ZN(n5611) );
  INV_X1 U5485 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5645) );
  INV_X1 U5486 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8881) );
  INV_X1 U5487 ( .A(n5681), .ZN(n5680) );
  AOI21_X1 U5488 ( .B1(n9159), .B2(n9074), .A(n5682), .ZN(n5681) );
  INV_X1 U5489 ( .A(n9159), .ZN(n5679) );
  NOR2_X1 U5490 ( .A1(n7887), .A2(n5819), .ZN(n10936) );
  AND2_X1 U5491 ( .A1(n5883), .A2(n6151), .ZN(n5399) );
  INV_X1 U5492 ( .A(n5883), .ZN(n5394) );
  OR2_X1 U5493 ( .A1(n5399), .A2(n9284), .ZN(n5395) );
  OR2_X1 U5494 ( .A1(n7960), .A2(n5263), .ZN(n5262) );
  NOR2_X1 U5495 ( .A1(n7969), .A2(n5829), .ZN(n5263) );
  INV_X1 U5496 ( .A(n8153), .ZN(n5410) );
  INV_X1 U5497 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U5498 ( .A1(n10004), .A2(n10146), .ZN(n5297) );
  AOI21_X1 U5499 ( .B1(n5705), .B2(n5707), .A(n5191), .ZN(n5703) );
  OR2_X1 U5500 ( .A1(n10086), .A2(n10020), .ZN(n9530) );
  AND2_X1 U5501 ( .A1(n5550), .A2(n9605), .ZN(n5546) );
  INV_X1 U5502 ( .A(n5317), .ZN(n5313) );
  AND2_X1 U5503 ( .A1(n5697), .A2(n5173), .ZN(n5695) );
  NAND2_X1 U5504 ( .A1(n5210), .A2(n5145), .ZN(n5709) );
  INV_X1 U5505 ( .A(n6155), .ZN(n5710) );
  AND2_X1 U5506 ( .A1(n9465), .A2(n9464), .ZN(n8204) );
  NAND2_X1 U5507 ( .A1(n5790), .A2(n5281), .ZN(n5791) );
  AND2_X1 U5508 ( .A1(n5786), .A2(n5139), .ZN(n5281) );
  AND2_X1 U5509 ( .A1(n5780), .A2(n5781), .ZN(n5788) );
  INV_X1 U5510 ( .A(n5484), .ZN(n5483) );
  OAI21_X1 U5511 ( .B1(n8977), .B2(n5485), .A(n9046), .ZN(n5484) );
  INV_X1 U5512 ( .A(n7318), .ZN(n5485) );
  NAND2_X1 U5513 ( .A1(n5488), .A2(n5494), .ZN(n5487) );
  NOR2_X1 U5514 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6547) );
  INV_X1 U5515 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U5516 ( .A1(n10646), .A2(n5421), .ZN(n5420) );
  INV_X1 U5517 ( .A(n5422), .ZN(n5421) );
  NOR2_X1 U5518 ( .A1(n10652), .A2(n10582), .ZN(n5422) );
  NOR2_X1 U5519 ( .A1(n8480), .A2(n8457), .ZN(n5418) );
  AND2_X1 U5520 ( .A1(n7042), .A2(n7041), .ZN(n7113) );
  NAND2_X1 U5521 ( .A1(n8348), .A2(n8318), .ZN(n8179) );
  NAND2_X1 U5522 ( .A1(n10228), .A2(n8058), .ZN(n7003) );
  INV_X1 U5523 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U5524 ( .A1(n6054), .A2(n6053), .ZN(n6336) );
  NAND2_X1 U5525 ( .A1(n5361), .A2(n5362), .ZN(n6054) );
  AOI21_X1 U5526 ( .B1(n5141), .B2(n5363), .A(n5241), .ZN(n5362) );
  INV_X1 U5527 ( .A(SI_19_), .ZN(n8715) );
  OAI21_X1 U5528 ( .B1(n6305), .B2(n6304), .A(n6303), .ZN(n6315) );
  NAND2_X1 U5529 ( .A1(n5364), .A2(n5366), .ZN(n6305) );
  NAND2_X1 U5530 ( .A1(n5365), .A2(n5369), .ZN(n5364) );
  INV_X1 U5531 ( .A(n6259), .ZN(n5365) );
  INV_X1 U5532 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5651) );
  AOI21_X1 U5533 ( .B1(n5601), .B2(n5600), .A(n5244), .ZN(n5599) );
  INV_X1 U5534 ( .A(n6021), .ZN(n5600) );
  AOI21_X1 U5535 ( .B1(n5383), .B2(n6182), .A(n5382), .ZN(n5381) );
  AOI21_X1 U5536 ( .B1(n5594), .B2(n5592), .A(n5203), .ZN(n5591) );
  NAND2_X1 U5537 ( .A1(n6183), .A2(n5383), .ZN(n5380) );
  INV_X1 U5538 ( .A(n5165), .ZN(n5670) );
  AOI21_X1 U5539 ( .B1(n5672), .B2(n5674), .A(n5208), .ZN(n5671) );
  NAND3_X1 U5540 ( .A1(n9359), .A2(n9360), .A3(n9954), .ZN(n9680) );
  AND2_X1 U5541 ( .A1(n8108), .A2(n8106), .ZN(n5687) );
  OR2_X1 U5542 ( .A1(n8995), .A2(n9799), .ZN(n5660) );
  NAND2_X1 U5543 ( .A1(n5692), .A2(n5770), .ZN(n5691) );
  INV_X1 U5544 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5770) );
  INV_X1 U5545 ( .A(n5769), .ZN(n5692) );
  OR4_X1 U5546 ( .A1(n9617), .A2(n9616), .A3(n9658), .A4(n9615), .ZN(n9619) );
  OAI21_X1 U5547 ( .B1(n9583), .B2(n9582), .A(n9586), .ZN(n5349) );
  AND4_X1 U5548 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n8425)
         );
  OR2_X1 U5549 ( .A1(n5879), .A2(n5582), .ZN(n5880) );
  OR2_X1 U5550 ( .A1(n7754), .A2(n7755), .ZN(n5278) );
  NAND2_X1 U5551 ( .A1(n7817), .A2(n5239), .ZN(n7799) );
  NAND2_X1 U5552 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  AND2_X1 U5553 ( .A1(n5837), .A2(n7568), .ZN(n5838) );
  NAND2_X1 U5554 ( .A1(n5891), .A2(n5410), .ZN(n5408) );
  NOR2_X1 U5555 ( .A1(n7869), .A2(n5891), .ZN(n5892) );
  NAND2_X1 U5556 ( .A1(n5848), .A2(n5849), .ZN(n5853) );
  INV_X1 U5557 ( .A(n5806), .ZN(n5855) );
  NAND2_X1 U5558 ( .A1(n5540), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5537) );
  INV_X1 U5559 ( .A(n9818), .ZN(n5540) );
  OR2_X1 U5560 ( .A1(n9851), .A2(n5530), .ZN(n5529) );
  NOR2_X1 U5561 ( .A1(n9857), .A2(n10097), .ZN(n5530) );
  NAND2_X1 U5562 ( .A1(n5556), .A2(n5555), .ZN(n9659) );
  AOI21_X1 U5563 ( .B1(n5558), .B2(n9402), .A(n5581), .ZN(n5555) );
  INV_X1 U5564 ( .A(n5720), .ZN(n5719) );
  OAI21_X1 U5565 ( .B1(n6418), .B2(n5721), .A(n5198), .ZN(n5720) );
  NAND2_X1 U5566 ( .A1(n6396), .A2(n9365), .ZN(n5721) );
  AND2_X1 U5567 ( .A1(n9570), .A2(n9571), .ZN(n9900) );
  AOI21_X1 U5568 ( .B1(n9918), .B2(n9917), .A(n5188), .ZN(n9907) );
  INV_X1 U5569 ( .A(n9788), .ZN(n9932) );
  OAI21_X1 U5570 ( .B1(n9952), .B2(n5318), .A(n5204), .ZN(n5732) );
  NOR2_X1 U5571 ( .A1(n5319), .A2(n9351), .ZN(n5318) );
  NAND2_X1 U5572 ( .A1(n9963), .A2(n9542), .ZN(n9952) );
  INV_X1 U5573 ( .A(n5293), .ZN(n5292) );
  INV_X1 U5574 ( .A(n5291), .ZN(n5290) );
  OAI21_X1 U5575 ( .B1(n5294), .B2(n5292), .A(n9977), .ZN(n5291) );
  NAND2_X1 U5576 ( .A1(n10018), .A2(n5705), .ZN(n5704) );
  NAND2_X1 U5577 ( .A1(n9995), .A2(n5297), .ZN(n5293) );
  NAND2_X1 U5578 ( .A1(n5704), .A2(n5294), .ZN(n5289) );
  NAND2_X1 U5579 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  INV_X1 U5580 ( .A(n6310), .ZN(n5959) );
  AND2_X1 U5581 ( .A1(n9530), .A2(n9531), .ZN(n10010) );
  NOR2_X1 U5582 ( .A1(n10024), .A2(n5568), .ZN(n5567) );
  NAND2_X1 U5583 ( .A1(n10018), .A2(n10024), .ZN(n10017) );
  AND4_X1 U5584 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(n9764)
         );
  NAND2_X1 U5585 ( .A1(n6453), .A2(n6452), .ZN(n9090) );
  AND2_X1 U5586 ( .A1(n9509), .A2(n9507), .ZN(n9607) );
  INV_X1 U5587 ( .A(n5551), .ZN(n5550) );
  OAI21_X1 U5588 ( .B1(n5552), .B2(n8404), .A(n9499), .ZN(n5551) );
  INV_X1 U5589 ( .A(n8405), .ZN(n5549) );
  NAND2_X1 U5590 ( .A1(n6235), .A2(n6234), .ZN(n8958) );
  NAND2_X1 U5591 ( .A1(n8405), .A2(n8404), .ZN(n8403) );
  AND2_X1 U5592 ( .A1(n9492), .A2(n9490), .ZN(n8414) );
  AND2_X1 U5593 ( .A1(n5698), .A2(n8422), .ZN(n5697) );
  NAND2_X1 U5594 ( .A1(n8421), .A2(n5699), .ZN(n5698) );
  INV_X1 U5595 ( .A(n6203), .ZN(n5699) );
  INV_X1 U5596 ( .A(n8421), .ZN(n5700) );
  OR2_X1 U5597 ( .A1(n11123), .A2(n8425), .ZN(n9484) );
  AND2_X1 U5598 ( .A1(n9484), .A2(n9475), .ZN(n9598) );
  AND2_X1 U5599 ( .A1(n5166), .A2(n9474), .ZN(n9597) );
  NAND2_X1 U5600 ( .A1(n5708), .A2(n5709), .ZN(n5712) );
  NOR2_X1 U5601 ( .A1(n9805), .A2(n5727), .ZN(n5725) );
  NAND2_X1 U5602 ( .A1(n5726), .A2(n5724), .ZN(n6142) );
  INV_X1 U5603 ( .A(n5727), .ZN(n5724) );
  NAND2_X1 U5604 ( .A1(n6445), .A2(n9591), .ZN(n8235) );
  NAND2_X1 U5605 ( .A1(n6117), .A2(n6442), .ZN(n10998) );
  NAND2_X1 U5606 ( .A1(n9580), .A2(n7520), .ZN(n11001) );
  INV_X1 U5607 ( .A(n7901), .ZN(n6100) );
  NOR2_X1 U5608 ( .A1(n8390), .A2(n8034), .ZN(n8394) );
  INV_X1 U5609 ( .A(n11001), .ZN(n10001) );
  OR2_X1 U5610 ( .A1(n9580), .A2(n7182), .ZN(n7988) );
  NAND2_X1 U5611 ( .A1(n9411), .A2(n9410), .ZN(n9424) );
  NAND2_X1 U5612 ( .A1(n6354), .A2(n6353), .ZN(n9432) );
  NAND2_X1 U5613 ( .A1(n6071), .A2(n6070), .ZN(n9553) );
  NAND2_X1 U5614 ( .A1(n6325), .A2(n6324), .ZN(n9539) );
  OR2_X1 U5615 ( .A1(n7485), .A2(n9627), .ZN(n11179) );
  NAND2_X1 U5616 ( .A1(n6489), .A2(n6488), .ZN(n6491) );
  INV_X1 U5617 ( .A(n5873), .ZN(n5944) );
  INV_X1 U5618 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5755) );
  AND2_X2 U5619 ( .A1(n5284), .A2(n5753), .ZN(n5584) );
  INV_X1 U5620 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5587) );
  NOR2_X1 U5621 ( .A1(n5178), .A2(n5143), .ZN(n5503) );
  NAND2_X1 U5622 ( .A1(n8039), .A2(n5480), .ZN(n5475) );
  NAND2_X1 U5623 ( .A1(n5476), .A2(n5478), .ZN(n5473) );
  AOI21_X1 U5624 ( .B1(n5503), .B2(n5501), .A(n5500), .ZN(n5499) );
  INV_X1 U5625 ( .A(n10187), .ZN(n5500) );
  INV_X1 U5626 ( .A(n5504), .ZN(n5501) );
  INV_X1 U5627 ( .A(n5503), .ZN(n5502) );
  INV_X1 U5628 ( .A(n7216), .ZN(n5497) );
  AND2_X1 U5629 ( .A1(n7084), .A2(n7018), .ZN(n7019) );
  NAND2_X1 U5630 ( .A1(n5431), .A2(n5184), .ZN(n7089) );
  NAND2_X1 U5631 ( .A1(n5433), .A2(n5432), .ZN(n5431) );
  AOI21_X1 U5632 ( .B1(n5441), .B2(n5443), .A(n5440), .ZN(n5437) );
  OR2_X1 U5633 ( .A1(n10607), .A2(n6986), .ZN(n7153) );
  OR2_X1 U5635 ( .A1(n6958), .A2(n6614), .ZN(n6615) );
  AOI21_X1 U5636 ( .B1(n10694), .B2(n6690), .A(n6526), .ZN(n9325) );
  NOR2_X1 U5637 ( .A1(n10614), .A2(n10618), .ZN(n5425) );
  INV_X1 U5638 ( .A(n5377), .ZN(n5374) );
  NOR2_X1 U5639 ( .A1(n10468), .A2(n5375), .ZN(n5373) );
  OR2_X1 U5640 ( .A1(n10492), .A2(n10632), .ZN(n10484) );
  AOI21_X2 U5641 ( .B1(n9310), .B2(n5169), .A(n5630), .ZN(n10460) );
  INV_X1 U5642 ( .A(n5631), .ZN(n5630) );
  AOI21_X1 U5643 ( .B1(n10479), .B2(n5634), .A(n5639), .ZN(n5631) );
  NAND2_X1 U5644 ( .A1(n5372), .A2(n9295), .ZN(n5510) );
  NAND2_X1 U5645 ( .A1(n10511), .A2(n5636), .ZN(n5635) );
  INV_X1 U5646 ( .A(n9312), .ZN(n5636) );
  NAND2_X1 U5647 ( .A1(n5623), .A2(n9296), .ZN(n10479) );
  INV_X1 U5648 ( .A(n5372), .ZN(n5512) );
  NAND2_X1 U5649 ( .A1(n5261), .A2(n5517), .ZN(n5514) );
  AOI21_X1 U5650 ( .B1(n5517), .B2(n10537), .A(n5516), .ZN(n5515) );
  AOI21_X1 U5651 ( .B1(n5142), .B2(n10575), .A(n5243), .ZN(n5654) );
  OR2_X1 U5652 ( .A1(n10574), .A2(n10575), .ZN(n5656) );
  AND2_X1 U5653 ( .A1(n9143), .A2(n9142), .ZN(n5628) );
  INV_X1 U5654 ( .A(n9143), .ZN(n11208) );
  OR2_X1 U5655 ( .A1(n8053), .A2(n8058), .ZN(n8089) );
  NOR2_X1 U5656 ( .A1(n5182), .A2(n5260), .ZN(n5259) );
  INV_X1 U5657 ( .A(n10507), .ZN(n11236) );
  NAND2_X1 U5658 ( .A1(n6936), .A2(n6935), .ZN(n10627) );
  NOR2_X1 U5659 ( .A1(n7460), .A2(n7576), .ZN(n8930) );
  NOR2_X1 U5660 ( .A1(n7574), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7460) );
  AND2_X1 U5661 ( .A1(n7637), .A2(n7736), .ZN(n8932) );
  AND2_X1 U5662 ( .A1(n7579), .A2(n7481), .ZN(n7639) );
  NOR2_X1 U5663 ( .A1(n6527), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U5664 ( .A1(n6508), .A2(n6507), .ZN(n6981) );
  OR2_X1 U5665 ( .A1(n6965), .A2(n6502), .ZN(n6508) );
  NAND2_X1 U5666 ( .A1(n5458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5457) );
  INV_X1 U5667 ( .A(n6527), .ZN(n5657) );
  INV_X1 U5668 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8904) );
  OAI21_X1 U5669 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6420) );
  MUX2_X1 U5670 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7168), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n7170) );
  NOR2_X1 U5671 ( .A1(n7165), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U5672 ( .A1(n5615), .A2(n6370), .ZN(n6383) );
  NAND2_X1 U5673 ( .A1(n5495), .A2(n5200), .ZN(n7165) );
  INV_X1 U5674 ( .A(n7160), .ZN(n5495) );
  INV_X1 U5675 ( .A(n5357), .ZN(n5356) );
  OAI21_X1 U5676 ( .B1(n5359), .B2(n5358), .A(n6068), .ZN(n5357) );
  NAND2_X1 U5677 ( .A1(n6059), .A2(n6058), .ZN(n6081) );
  XNOR2_X1 U5678 ( .A(n6305), .B(n6293), .ZN(n8065) );
  OAI21_X1 U5679 ( .B1(n6259), .B2(n5371), .A(n5604), .ZN(n6283) );
  INV_X1 U5680 ( .A(n5653), .ZN(n5652) );
  XNOR2_X1 U5681 ( .A(n6171), .B(n6170), .ZN(n7553) );
  OAI21_X1 U5682 ( .B1(n6152), .B2(n5508), .A(n5506), .ZN(n6171) );
  NAND2_X1 U5683 ( .A1(n6167), .A2(SI_5_), .ZN(n5508) );
  INV_X1 U5684 ( .A(n5507), .ZN(n5506) );
  XNOR2_X1 U5685 ( .A(n6168), .B(n6162), .ZN(n7555) );
  OAI21_X1 U5686 ( .B1(n6152), .B2(n5995), .A(n5994), .ZN(n6168) );
  NOR2_X1 U5687 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6516) );
  NAND2_X1 U5688 ( .A1(n8107), .A2(n5687), .ZN(n8268) );
  AND2_X1 U5689 ( .A1(n6185), .A2(n6184), .ZN(n11104) );
  AND2_X1 U5690 ( .A1(n6154), .A2(n6153), .ZN(n11048) );
  AND4_X1 U5691 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n10019)
         );
  INV_X1 U5692 ( .A(n9790), .ZN(n9954) );
  NAND2_X1 U5693 ( .A1(n6347), .A2(n6346), .ZN(n9978) );
  INV_X1 U5694 ( .A(n9744), .ZN(n10004) );
  INV_X1 U5695 ( .A(n9764), .ZN(n10002) );
  AND2_X1 U5696 ( .A1(n6113), .A2(n6114), .ZN(n5285) );
  NOR2_X1 U5697 ( .A1(n7888), .A2(n10982), .ZN(n7887) );
  AND2_X1 U5698 ( .A1(n5280), .A2(n5279), .ZN(n7754) );
  NAND2_X1 U5699 ( .A1(n5922), .A2(n7559), .ZN(n5279) );
  NOR2_X1 U5700 ( .A1(n8141), .A2(n5847), .ZN(n8361) );
  OR2_X1 U5701 ( .A1(n9117), .A2(n11186), .ZN(n5539) );
  NOR2_X1 U5702 ( .A1(n9866), .A2(n9865), .ZN(n9867) );
  AND2_X1 U5703 ( .A1(n9864), .A2(n9863), .ZN(n9865) );
  INV_X1 U5704 ( .A(n5543), .ZN(n9866) );
  NAND2_X1 U5705 ( .A1(n9871), .A2(n5272), .ZN(n9877) );
  XNOR2_X1 U5706 ( .A(n5529), .B(n8064), .ZN(n9861) );
  NOR2_X1 U5707 ( .A1(n9861), .A2(n9862), .ZN(n9860) );
  NOR2_X1 U5708 ( .A1(n10969), .A2(n5904), .ZN(n5905) );
  NAND2_X1 U5709 ( .A1(n5869), .A2(n5868), .ZN(n5527) );
  OAI21_X1 U5710 ( .B1(n5270), .B2(n5269), .A(n5266), .ZN(n5265) );
  OR4_X1 U5711 ( .A1(n5275), .A2(n5274), .A3(n5276), .A4(n5235), .ZN(n5271) );
  NOR2_X1 U5712 ( .A1(n5276), .A2(n5267), .ZN(n5266) );
  NOR2_X1 U5713 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  OR2_X1 U5714 ( .A1(n9396), .A2(n11181), .ZN(n6464) );
  AND2_X1 U5715 ( .A1(n6389), .A2(n6388), .ZN(n10122) );
  AND2_X1 U5716 ( .A1(n10053), .A2(n11159), .ZN(n5299) );
  AND2_X1 U5717 ( .A1(n7580), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7481) );
  AND2_X1 U5718 ( .A1(n7393), .A2(n7405), .ZN(n5472) );
  NAND2_X1 U5719 ( .A1(n7470), .A2(n9220), .ZN(n10300) );
  NAND2_X1 U5720 ( .A1(n6922), .A2(n6921), .ZN(n10642) );
  NAND2_X1 U5721 ( .A1(n6864), .A2(n6863), .ZN(n10664) );
  OR2_X1 U5722 ( .A1(n6987), .A2(n8890), .ZN(n7091) );
  INV_X1 U5723 ( .A(n5379), .ZN(n10445) );
  OAI21_X1 U5724 ( .B1(n10470), .B2(n10469), .A(n11232), .ZN(n10474) );
  AND2_X1 U5725 ( .A1(n5166), .A2(n9484), .ZN(n9463) );
  AOI21_X1 U5726 ( .B1(n5453), .B2(n6949), .A(n5452), .ZN(n5451) );
  INV_X1 U5727 ( .A(n7029), .ZN(n5452) );
  OR2_X1 U5728 ( .A1(n7910), .A2(n7027), .ZN(n5453) );
  INV_X1 U5729 ( .A(n8179), .ZN(n7000) );
  NAND2_X1 U5730 ( .A1(n5326), .A2(n5237), .ZN(n5325) );
  NAND2_X1 U5731 ( .A1(n9493), .A2(n9492), .ZN(n5326) );
  AOI21_X1 U5732 ( .B1(n5324), .B2(n9580), .A(n9603), .ZN(n5323) );
  NAND2_X1 U5733 ( .A1(n9481), .A2(n9490), .ZN(n5324) );
  NOR2_X1 U5734 ( .A1(n6826), .A2(n7094), .ZN(n6827) );
  OAI21_X1 U5735 ( .B1(n6737), .B2(n5463), .A(n5459), .ZN(n5462) );
  INV_X1 U5736 ( .A(n5460), .ZN(n5459) );
  OR2_X1 U5737 ( .A1(n9511), .A2(n5333), .ZN(n5332) );
  NAND2_X1 U5738 ( .A1(n5337), .A2(n9580), .ZN(n5333) );
  OR2_X1 U5739 ( .A1(n9512), .A2(n5336), .ZN(n5335) );
  NAND2_X1 U5740 ( .A1(n5337), .A2(n9574), .ZN(n5336) );
  OR2_X1 U5741 ( .A1(n9523), .A2(n9522), .ZN(n5334) );
  AOI21_X1 U5742 ( .B1(n6888), .B2(n6949), .A(n10566), .ZN(n6889) );
  OAI21_X1 U5743 ( .B1(n5328), .B2(n5327), .A(n5201), .ZN(n9565) );
  NAND2_X1 U5744 ( .A1(n9558), .A2(n9929), .ZN(n5327) );
  AOI21_X1 U5745 ( .B1(n9549), .B2(n5330), .A(n5329), .ZN(n5328) );
  NAND2_X1 U5746 ( .A1(n5513), .A2(n9294), .ZN(n5622) );
  INV_X1 U5747 ( .A(n6947), .ZN(n5620) );
  OR2_X1 U5748 ( .A1(n7138), .A2(n7068), .ZN(n5469) );
  AOI21_X1 U5749 ( .B1(n6948), .B2(n9296), .A(n7070), .ZN(n5468) );
  NAND2_X1 U5750 ( .A1(n5450), .A2(n10443), .ZN(n5449) );
  NOR2_X1 U5751 ( .A1(n7337), .A2(n10215), .ZN(n7123) );
  INV_X1 U5752 ( .A(SI_17_), .ZN(n8723) );
  INV_X1 U5753 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8626) );
  INV_X1 U5754 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8841) );
  NOR2_X1 U5755 ( .A1(n5344), .A2(n9577), .ZN(n5343) );
  NAND2_X1 U5756 ( .A1(n9868), .A2(n5252), .ZN(n5938) );
  INV_X1 U5757 ( .A(n6292), .ZN(n5707) );
  NAND2_X1 U5758 ( .A1(n9807), .A2(n11008), .ZN(n9445) );
  AND2_X1 U5759 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n6883), .ZN(n6882) );
  AND2_X1 U5760 ( .A1(n10230), .A2(n8005), .ZN(n7106) );
  NOR2_X1 U5761 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5642) );
  NAND2_X1 U5762 ( .A1(n6501), .A2(n6500), .ZN(n6503) );
  NOR2_X1 U5763 ( .A1(n6382), .A2(n5614), .ZN(n5613) );
  INV_X1 U5764 ( .A(n6370), .ZN(n5614) );
  INV_X1 U5765 ( .A(SI_20_), .ZN(n8716) );
  INV_X1 U5766 ( .A(SI_18_), .ZN(n8721) );
  INV_X1 U5767 ( .A(n6282), .ZN(n5370) );
  INV_X1 U5768 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6037) );
  INV_X1 U5769 ( .A(n6032), .ZN(n5608) );
  INV_X1 U5770 ( .A(SI_15_), .ZN(n8728) );
  INV_X1 U5771 ( .A(SI_14_), .ZN(n8729) );
  NAND2_X1 U5772 ( .A1(n6022), .A2(n6021), .ZN(n5603) );
  INV_X1 U5773 ( .A(SI_12_), .ZN(n8733) );
  INV_X1 U5774 ( .A(n6011), .ZN(n5595) );
  INV_X1 U5775 ( .A(n5742), .ZN(n5592) );
  INV_X1 U5776 ( .A(SI_10_), .ZN(n8739) );
  INV_X1 U5777 ( .A(SI_9_), .ZN(n8738) );
  AND2_X1 U5778 ( .A1(n5740), .A2(n9335), .ZN(n5683) );
  INV_X1 U5779 ( .A(n5581), .ZN(n5580) );
  AND2_X1 U5780 ( .A1(n9422), .A2(n5225), .ZN(n5578) );
  AND2_X1 U5781 ( .A1(n9586), .A2(n9421), .ZN(n9422) );
  NOR2_X1 U5782 ( .A1(n9785), .A2(n9405), .ZN(n5579) );
  INV_X1 U5783 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8585) );
  INV_X1 U5784 ( .A(n5408), .ZN(n5406) );
  NOR2_X1 U5785 ( .A1(n5409), .A2(n7871), .ZN(n5403) );
  INV_X1 U5786 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U5787 ( .A1(n9844), .A2(n5934), .ZN(n9869) );
  NAND2_X1 U5788 ( .A1(n9869), .A2(n9870), .ZN(n9868) );
  AND3_X1 U5789 ( .A1(n5561), .A2(n5560), .A3(n5255), .ZN(n5902) );
  INV_X1 U5790 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5564) );
  INV_X1 U5791 ( .A(n5559), .ZN(n5558) );
  OAI21_X1 U5792 ( .B1(n6462), .B2(n9402), .A(n9655), .ZN(n5559) );
  AND2_X1 U5793 ( .A1(n9677), .A2(n9908), .ZN(n9431) );
  INV_X1 U5794 ( .A(n6418), .ZN(n5722) );
  INV_X1 U5795 ( .A(n10122), .ZN(n6461) );
  INV_X1 U5796 ( .A(n5220), .ZN(n5574) );
  NOR2_X1 U5797 ( .A1(n11002), .A2(n11027), .ZN(n5727) );
  OR2_X1 U5798 ( .A1(n7538), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6483) );
  NOR2_X1 U5799 ( .A1(n5782), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5785) );
  INV_X1 U5800 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U5801 ( .A1(n5283), .A2(n5149), .ZN(n5282) );
  AND2_X1 U5802 ( .A1(n6882), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U5803 ( .A1(n8040), .A2(n8041), .ZN(n5479) );
  INV_X1 U5804 ( .A(n6989), .ZN(n5440) );
  NAND2_X1 U5805 ( .A1(n10443), .A2(n6985), .ZN(n5444) );
  INV_X1 U5806 ( .A(n6979), .ZN(n5433) );
  NAND2_X1 U5807 ( .A1(n5435), .A2(n5438), .ZN(n5432) );
  NAND2_X1 U5808 ( .A1(n5441), .A2(n5189), .ZN(n5438) );
  NAND2_X1 U5809 ( .A1(n5434), .A2(n5446), .ZN(n5430) );
  NAND2_X1 U5810 ( .A1(n5378), .A2(n5376), .ZN(n5375) );
  INV_X1 U5811 ( .A(n10467), .ZN(n5376) );
  INV_X1 U5812 ( .A(n5635), .ZN(n5632) );
  OR2_X1 U5813 ( .A1(n10627), .A2(n10482), .ZN(n7069) );
  AND2_X1 U5814 ( .A1(n10664), .A2(n10199), .ZN(n9291) );
  OR2_X1 U5815 ( .A1(n10664), .A2(n10199), .ZN(n7063) );
  NOR2_X1 U5816 ( .A1(n7061), .A2(n5522), .ZN(n5521) );
  NOR2_X1 U5817 ( .A1(n11234), .A2(n5523), .ZN(n5522) );
  NOR2_X1 U5818 ( .A1(n10290), .A2(n5428), .ZN(n5427) );
  INV_X1 U5819 ( .A(n5429), .ZN(n5428) );
  NOR2_X1 U5820 ( .A1(n10602), .A2(n11260), .ZN(n5429) );
  NAND2_X1 U5821 ( .A1(n5745), .A2(n8940), .ZN(n8942) );
  INV_X1 U5822 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U5823 ( .A1(n6789), .A2(n6788), .ZN(n6804) );
  OR2_X1 U5824 ( .A1(n8005), .A2(n10230), .ZN(n7108) );
  INV_X1 U5825 ( .A(n10335), .ZN(n8051) );
  NAND2_X1 U5826 ( .A1(n10598), .A2(n11224), .ZN(n11249) );
  OAI21_X1 U5827 ( .B1(n7574), .B2(P1_D_REG_1__SCAN_IN), .A(n10687), .ZN(n7736) );
  XNOR2_X1 U5828 ( .A(n6503), .B(n6504), .ZN(n6965) );
  NOR2_X1 U5829 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5646) );
  NAND2_X1 U5830 ( .A1(n6783), .A2(n6546), .ZN(n7160) );
  NAND2_X1 U5831 ( .A1(n5354), .A2(n5352), .ZN(n6369) );
  AOI21_X1 U5832 ( .B1(n5356), .B2(n5358), .A(n5353), .ZN(n5352) );
  INV_X1 U5833 ( .A(n6348), .ZN(n5353) );
  AND2_X1 U5834 ( .A1(n6370), .A2(n6352), .ZN(n6368) );
  NOR2_X1 U5835 ( .A1(n6080), .A2(n5360), .ZN(n5359) );
  INV_X1 U5836 ( .A(n6058), .ZN(n5360) );
  AOI21_X1 U5837 ( .B1(n5606), .B2(n5607), .A(n5605), .ZN(n5604) );
  INV_X1 U5838 ( .A(n6036), .ZN(n5605) );
  INV_X1 U5839 ( .A(n6030), .ZN(n5606) );
  INV_X1 U5840 ( .A(n5607), .ZN(n5371) );
  INV_X1 U5841 ( .A(n6214), .ZN(n5385) );
  OAI21_X1 U5842 ( .B1(n5994), .B2(n6162), .A(n6169), .ZN(n5507) );
  NAND2_X1 U5843 ( .A1(n8996), .A2(n8995), .ZN(n5661) );
  NAND2_X1 U5844 ( .A1(n9332), .A2(n9331), .ZN(n5684) );
  OR2_X1 U5845 ( .A1(n8996), .A2(n8995), .ZN(n9027) );
  XNOR2_X1 U5846 ( .A(n10978), .B(n7783), .ZN(n7489) );
  NAND2_X1 U5847 ( .A1(n5957), .A2(n9727), .ZN(n6296) );
  INV_X1 U5848 ( .A(n6286), .ZN(n5957) );
  INV_X1 U5849 ( .A(n9763), .ZN(n9776) );
  AOI21_X1 U5850 ( .B1(n5681), .B2(n5679), .A(n5678), .ZN(n5677) );
  INV_X1 U5851 ( .A(n9192), .ZN(n5678) );
  NAND2_X1 U5852 ( .A1(n5956), .A2(n9207), .ZN(n6274) );
  INV_X1 U5853 ( .A(n6264), .ZN(n5956) );
  NAND2_X1 U5854 ( .A1(n7509), .A2(n7545), .ZN(n7514) );
  NOR2_X1 U5855 ( .A1(n7892), .A2(n7893), .ZN(n7891) );
  XNOR2_X1 U5856 ( .A(n5919), .B(n7901), .ZN(n7893) );
  NAND2_X1 U5857 ( .A1(n5411), .A2(n5877), .ZN(n7890) );
  OR2_X1 U5858 ( .A1(n7901), .A2(n5876), .ZN(n5411) );
  OR2_X1 U5859 ( .A1(n7965), .A2(n7966), .ZN(n5280) );
  NAND2_X1 U5860 ( .A1(n7954), .A2(n5883), .ZN(n5392) );
  NAND2_X1 U5861 ( .A1(n7954), .A2(n5399), .ZN(n5398) );
  OAI211_X1 U5862 ( .C1(n7954), .C2(n5396), .A(n5395), .B(n5393), .ZN(n5885)
         );
  NOR2_X1 U5863 ( .A1(n5528), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U5864 ( .A1(n5394), .A2(n5528), .ZN(n5393) );
  OR2_X1 U5865 ( .A1(n5397), .A2(n7822), .ZN(n7825) );
  NAND2_X1 U5866 ( .A1(n5398), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5397) );
  INV_X1 U5867 ( .A(n5262), .ZN(n5831) );
  AOI21_X1 U5868 ( .B1(n7830), .B2(n5163), .A(n7829), .ZN(n7828) );
  OR2_X1 U5869 ( .A1(n7801), .A2(n8221), .ZN(n7803) );
  NAND2_X1 U5870 ( .A1(n7797), .A2(n5238), .ZN(n7883) );
  NAND2_X1 U5871 ( .A1(n7883), .A2(n7882), .ZN(n7881) );
  NAND2_X1 U5872 ( .A1(n7875), .A2(n5844), .ZN(n5533) );
  INV_X1 U5873 ( .A(n5838), .ZN(n5535) );
  AND2_X1 U5874 ( .A1(n5213), .A2(n5575), .ZN(n9016) );
  NAND2_X1 U5875 ( .A1(n9845), .A2(n9846), .ZN(n9844) );
  OR2_X1 U5876 ( .A1(n9829), .A2(n5562), .ZN(n5561) );
  NAND2_X1 U5877 ( .A1(n5563), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5562) );
  INV_X1 U5878 ( .A(n9843), .ZN(n5563) );
  OR2_X1 U5879 ( .A1(n5161), .A2(n9843), .ZN(n5560) );
  INV_X1 U5880 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5768) );
  INV_X1 U5881 ( .A(n5529), .ZN(n5865) );
  INV_X1 U5882 ( .A(n5268), .ZN(n5267) );
  AOI21_X1 U5883 ( .B1(n5273), .B2(n5272), .A(n5948), .ZN(n5268) );
  INV_X1 U5884 ( .A(n5940), .ZN(n5273) );
  NOR2_X1 U5885 ( .A1(n10953), .A2(n10956), .ZN(n5275) );
  INV_X1 U5886 ( .A(n10954), .ZN(n5274) );
  INV_X1 U5887 ( .A(n5943), .ZN(n5276) );
  NOR2_X1 U5888 ( .A1(n10953), .A2(n10956), .ZN(n5270) );
  NAND2_X1 U5889 ( .A1(n10954), .A2(n5272), .ZN(n5269) );
  NOR2_X1 U5890 ( .A1(n5719), .A2(n5717), .ZN(n5716) );
  INV_X1 U5891 ( .A(n9652), .ZN(n5717) );
  INV_X1 U5892 ( .A(n9919), .ZN(n9917) );
  AND2_X1 U5893 ( .A1(n9563), .A2(n9562), .ZN(n9919) );
  NOR2_X1 U5894 ( .A1(n10130), .A2(n9944), .ZN(n6366) );
  AND2_X1 U5895 ( .A1(n9551), .A2(n9550), .ZN(n9956) );
  AOI21_X1 U5896 ( .B1(n5290), .B2(n5292), .A(n5288), .ZN(n5287) );
  INV_X1 U5897 ( .A(n6334), .ZN(n5288) );
  NAND2_X1 U5898 ( .A1(n5704), .A2(n5703), .ZN(n9987) );
  NAND2_X1 U5899 ( .A1(n5544), .A2(n5545), .ZN(n9060) );
  AOI21_X1 U5900 ( .B1(n5546), .B2(n5552), .A(n5554), .ZN(n5545) );
  INV_X1 U5901 ( .A(n5309), .ZN(n5308) );
  NAND2_X1 U5902 ( .A1(n5309), .A2(n5311), .ZN(n5307) );
  NAND2_X1 U5903 ( .A1(n5314), .A2(n5317), .ZN(n8964) );
  NAND2_X1 U5904 ( .A1(n5314), .A2(n5312), .ZN(n9062) );
  NAND2_X1 U5905 ( .A1(n5954), .A2(n5953), .ZN(n6240) );
  INV_X1 U5906 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5953) );
  INV_X1 U5907 ( .A(n6228), .ZN(n5954) );
  AOI21_X1 U5908 ( .B1(n5152), .B2(n5697), .A(n5234), .ZN(n5696) );
  INV_X1 U5909 ( .A(n5305), .ZN(n5304) );
  OAI21_X1 U5910 ( .B1(n9595), .B2(n5306), .A(n6192), .ZN(n5305) );
  OAI21_X1 U5911 ( .B1(n9277), .B2(n9276), .A(n9457), .ZN(n8205) );
  INV_X1 U5912 ( .A(n11008), .ZN(n6116) );
  OR2_X1 U5913 ( .A1(n6103), .A2(n10978), .ZN(n10995) );
  CLKBUF_X1 U5914 ( .A(n9438), .Z(n10996) );
  INV_X1 U5915 ( .A(n7484), .ZN(n8191) );
  AND3_X1 U5916 ( .A1(n6140), .A2(n6139), .A3(n6138), .ZN(n11035) );
  AND2_X1 U5917 ( .A1(n9660), .A2(n11135), .ZN(n11181) );
  XNOR2_X1 U5918 ( .A(n5765), .B(n5764), .ZN(n7508) );
  INV_X1 U5919 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5764) );
  OR2_X1 U5920 ( .A1(n5776), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5763) );
  INV_X1 U5921 ( .A(n7514), .ZN(n7539) );
  XNOR2_X1 U5922 ( .A(n5761), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6482) );
  INV_X1 U5923 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5773) );
  INV_X1 U5924 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5767) );
  INV_X1 U5925 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5926 ( .A1(n5482), .A2(n5481), .ZN(n9096) );
  AOI21_X1 U5927 ( .B1(n5483), .B2(n5485), .A(n5206), .ZN(n5481) );
  OR2_X1 U5928 ( .A1(n7361), .A2(n7373), .ZN(n5504) );
  AND2_X1 U5929 ( .A1(n7273), .A2(n7272), .ZN(n8313) );
  INV_X1 U5930 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6773) );
  OR2_X1 U5931 ( .A1(n6774), .A2(n6773), .ZN(n6789) );
  INV_X1 U5932 ( .A(n5491), .ZN(n5489) );
  NAND2_X1 U5933 ( .A1(n5233), .A2(n5492), .ZN(n5491) );
  INV_X1 U5934 ( .A(n10248), .ZN(n5492) );
  NAND2_X1 U5935 ( .A1(n10180), .A2(n5493), .ZN(n5490) );
  AND2_X1 U5936 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6671) );
  NOR2_X1 U5937 ( .A1(n6728), .A2(n7629), .ZN(n6744) );
  NAND2_X1 U5938 ( .A1(n7674), .A2(n7672), .ZN(n7673) );
  INV_X1 U5939 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U5940 ( .A1(n7317), .A2(n8977), .ZN(n8980) );
  INV_X1 U5941 ( .A(n6818), .ZN(n6838) );
  INV_X1 U5942 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8890) );
  AND2_X1 U5943 ( .A1(n10878), .A2(n10424), .ZN(n10892) );
  INV_X1 U5944 ( .A(n10455), .ZN(n5378) );
  NAND2_X1 U5945 ( .A1(n7069), .A2(n7074), .ZN(n10467) );
  INV_X1 U5946 ( .A(n6831), .ZN(n6538) );
  NAND2_X1 U5947 ( .A1(n6813), .A2(n6537), .ZN(n6831) );
  INV_X1 U5948 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8669) );
  INV_X1 U5949 ( .A(n10513), .ZN(n10483) );
  INV_X1 U5950 ( .A(n10323), .ZN(n10482) );
  AND2_X1 U5951 ( .A1(n6570), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6569) );
  AND2_X1 U5952 ( .A1(n10577), .A2(n5216), .ZN(n10520) );
  INV_X1 U5953 ( .A(n10642), .ZN(n5419) );
  AOI21_X1 U5954 ( .B1(n5261), .B2(n10538), .A(n10537), .ZN(n10535) );
  NAND2_X1 U5955 ( .A1(n10577), .A2(n5420), .ZN(n10529) );
  INV_X1 U5956 ( .A(n9291), .ZN(n10565) );
  NAND2_X1 U5957 ( .A1(n10577), .A2(n10658), .ZN(n10576) );
  NOR2_X1 U5958 ( .A1(n10664), .A2(n9226), .ZN(n10577) );
  NAND2_X1 U5959 ( .A1(n10598), .A2(n5426), .ZN(n9226) );
  AND2_X1 U5960 ( .A1(n5427), .A2(n9223), .ZN(n5426) );
  AND2_X1 U5961 ( .A1(n7063), .A2(n10565), .ZN(n9306) );
  AOI21_X1 U5962 ( .B1(n5521), .B2(n5523), .A(n6859), .ZN(n5520) );
  NAND2_X1 U5963 ( .A1(n10598), .A2(n5427), .ZN(n9186) );
  AND2_X1 U5964 ( .A1(n11231), .A2(n7129), .ZN(n9133) );
  AND2_X1 U5965 ( .A1(n11260), .A2(n10595), .ZN(n5640) );
  AND2_X1 U5966 ( .A1(n7060), .A2(n6994), .ZN(n9146) );
  CLKBUF_X1 U5967 ( .A(n11230), .Z(n11233) );
  NAND2_X1 U5968 ( .A1(n11233), .A2(n11234), .ZN(n11231) );
  NAND2_X1 U5969 ( .A1(n7058), .A2(n7126), .ZN(n10592) );
  INV_X1 U5970 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U5971 ( .A1(n7054), .A2(n7053), .ZN(n11207) );
  AND2_X1 U5972 ( .A1(n5151), .A2(n11193), .ZN(n5416) );
  AND2_X1 U5973 ( .A1(n7118), .A2(n6997), .ZN(n8483) );
  NAND2_X1 U5974 ( .A1(n8334), .A2(n5418), .ZN(n8484) );
  AND2_X1 U5975 ( .A1(n7050), .A2(n6996), .ZN(n8458) );
  AND2_X1 U5976 ( .A1(n8334), .A2(n11152), .ZN(n8459) );
  OAI21_X1 U5977 ( .B1(n8178), .B2(n7043), .A(n7113), .ZN(n7045) );
  NAND2_X1 U5978 ( .A1(n8129), .A2(n8130), .ZN(n5505) );
  NOR2_X1 U5979 ( .A1(n8290), .A2(n11112), .ZN(n8293) );
  OR2_X1 U5980 ( .A1(n6717), .A2(n6716), .ZN(n6728) );
  INV_X1 U5981 ( .A(n8124), .ZN(n8181) );
  AND2_X1 U5982 ( .A1(n7038), .A2(n8179), .ZN(n8352) );
  NOR2_X1 U5983 ( .A1(n8090), .A2(n8119), .ZN(n8344) );
  NAND2_X1 U5984 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  AND3_X1 U5985 ( .A1(n7739), .A2(n8929), .A3(n7738), .ZN(n7741) );
  NAND2_X1 U5986 ( .A1(n7907), .A2(n7906), .ZN(n8074) );
  NOR2_X1 U5987 ( .A1(n10609), .A2(n7172), .ZN(n7636) );
  NAND2_X1 U5988 ( .A1(n7910), .A2(n7909), .ZN(n8048) );
  INV_X1 U5989 ( .A(n7911), .ZN(n7649) );
  OR2_X1 U5990 ( .A1(n7652), .A2(n7647), .ZN(n10609) );
  INV_X1 U5991 ( .A(n10609), .ZN(n11250) );
  INV_X1 U5992 ( .A(n11269), .ZN(n11111) );
  AND2_X1 U5993 ( .A1(n8947), .A2(n11069), .ZN(n10671) );
  NAND2_X1 U5994 ( .A1(n6529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6528) );
  INV_X1 U5995 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U5996 ( .A1(n7156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7157) );
  XNOR2_X1 U5997 ( .A(n6315), .B(n6316), .ZN(n8278) );
  XNOR2_X1 U5998 ( .A(n6271), .B(n6270), .ZN(n7971) );
  NAND2_X1 U5999 ( .A1(n5609), .A2(n6032), .ZN(n6271) );
  OR4_X1 U6000 ( .A1(n6766), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .A4(P1_IR_REG_9__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U6001 ( .A1(n5380), .A2(n5381), .ZN(n6215) );
  INV_X1 U6002 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8867) );
  INV_X1 U6003 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8860) );
  INV_X1 U6004 ( .A(n6097), .ZN(n5619) );
  AND2_X1 U6005 ( .A1(n8107), .A2(n8106), .ZN(n8109) );
  NAND2_X1 U6006 ( .A1(n9772), .A2(n9371), .ZN(n9673) );
  AND2_X1 U6007 ( .A1(n9360), .A2(n9359), .ZN(n9681) );
  NAND2_X1 U6008 ( .A1(n9027), .A2(n5661), .ZN(n8997) );
  AND4_X1 U6009 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n10020)
         );
  NOR2_X1 U6010 ( .A1(n5673), .A2(n5670), .ZN(n5668) );
  NAND2_X1 U6011 ( .A1(n5667), .A2(n5666), .ZN(n5665) );
  OR2_X1 U6012 ( .A1(n5671), .A2(n5165), .ZN(n5666) );
  NAND2_X1 U6013 ( .A1(n5671), .A2(n5190), .ZN(n5667) );
  NAND2_X1 U6014 ( .A1(n5671), .A2(n5670), .ZN(n5669) );
  NAND2_X1 U6015 ( .A1(n8268), .A2(n8267), .ZN(n8303) );
  AND4_X1 U6016 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n9153)
         );
  AND4_X1 U6017 ( .A1(n6269), .A2(n6268), .A3(n6267), .A4(n6266), .ZN(n9244)
         );
  NAND2_X1 U6018 ( .A1(n5684), .A2(n9335), .ZN(n9725) );
  INV_X1 U6019 ( .A(n5686), .ZN(n5685) );
  OR2_X1 U6020 ( .A1(n8302), .A2(n8304), .ZN(n5688) );
  NAND2_X1 U6021 ( .A1(n11010), .A2(n7525), .ZN(n9731) );
  NOR2_X1 U6022 ( .A1(n9749), .A2(n5663), .ZN(n5662) );
  INV_X1 U6023 ( .A(n9350), .ZN(n5663) );
  NAND2_X1 U6024 ( .A1(n9705), .A2(n9350), .ZN(n9750) );
  AND2_X1 U6025 ( .A1(n7518), .A2(n7517), .ZN(n9779) );
  INV_X1 U6026 ( .A(n9754), .ZN(n9781) );
  OR2_X1 U6027 ( .A1(n7522), .A2(n7521), .ZN(n9763) );
  INV_X1 U6028 ( .A(n9748), .ZN(n9773) );
  INV_X1 U6029 ( .A(n9731), .ZN(n9784) );
  NAND2_X1 U6030 ( .A1(n5347), .A2(n5186), .ZN(n9622) );
  OAI21_X1 U6031 ( .B1(n9585), .B2(n5349), .A(n5348), .ZN(n5347) );
  AND2_X1 U6032 ( .A1(n9584), .A2(n8387), .ZN(n5348) );
  XNOR2_X1 U6033 ( .A(n5777), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9627) );
  AND2_X1 U6034 ( .A1(n8264), .A2(n8263), .ZN(n9663) );
  NAND2_X1 U6035 ( .A1(n6332), .A2(n6331), .ZN(n9988) );
  INV_X1 U6036 ( .A(n10020), .ZN(n9791) );
  INV_X1 U6037 ( .A(n10019), .ZN(n9793) );
  INV_X1 U6038 ( .A(n9244), .ZN(n9794) );
  INV_X1 U6039 ( .A(P2_U3893), .ZN(n10961) );
  AND3_X1 U6040 ( .A1(n6085), .A2(n6086), .A3(n5589), .ZN(n5588) );
  NAND2_X1 U6041 ( .A1(n5817), .A2(n5818), .ZN(n7888) );
  OAI21_X1 U6042 ( .B1(n7890), .B2(n7889), .A(n5877), .ZN(n10948) );
  NAND2_X1 U6043 ( .A1(n10948), .A2(n10949), .ZN(n10947) );
  XNOR2_X1 U6044 ( .A(n6107), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n10949) );
  INV_X1 U6045 ( .A(n5280), .ZN(n7964) );
  OR2_X1 U6046 ( .A1(P2_U3150), .A2(n5942), .ZN(n9873) );
  INV_X1 U6047 ( .A(n5278), .ZN(n7753) );
  NAND2_X1 U6048 ( .A1(n5923), .A2(n5528), .ZN(n5277) );
  NOR2_X1 U6049 ( .A1(n7795), .A2(n5838), .ZN(n7876) );
  NAND2_X1 U6050 ( .A1(n5401), .A2(n5405), .ZN(n5404) );
  NAND2_X1 U6051 ( .A1(n5388), .A2(n5390), .ZN(n8440) );
  INV_X1 U6052 ( .A(n5575), .ZN(n8438) );
  NOR2_X1 U6053 ( .A1(n8437), .A2(n11147), .ZN(n8436) );
  OAI21_X1 U6054 ( .B1(n5158), .B2(n8437), .A(n5531), .ZN(n9005) );
  NOR2_X1 U6055 ( .A1(n9120), .A2(n9119), .ZN(n9118) );
  INV_X1 U6056 ( .A(n5861), .ZN(n5538) );
  OAI21_X1 U6057 ( .B1(n9120), .B2(n5414), .A(n5412), .ZN(n9808) );
  OR2_X1 U6058 ( .A1(n9809), .A2(n9119), .ZN(n5414) );
  NAND2_X1 U6059 ( .A1(n5898), .A2(n5413), .ZN(n5412) );
  INV_X1 U6060 ( .A(n9809), .ZN(n5413) );
  OR2_X1 U6061 ( .A1(n9829), .A2(n9828), .ZN(n5565) );
  NAND2_X1 U6062 ( .A1(n5561), .A2(n5560), .ZN(n9842) );
  INV_X1 U6063 ( .A(n5542), .ZN(n10971) );
  OAI21_X1 U6064 ( .B1(n9897), .B2(n11000), .A(n9896), .ZN(n10048) );
  NOR2_X1 U6065 ( .A1(n9921), .A2(n11001), .ZN(n9895) );
  INV_X1 U6066 ( .A(n6367), .ZN(n9930) );
  INV_X1 U6067 ( .A(n5732), .ZN(n9941) );
  NAND2_X1 U6068 ( .A1(n6338), .A2(n6337), .ZN(n10072) );
  NAND2_X1 U6069 ( .A1(n9980), .A2(n5570), .ZN(n9970) );
  NAND2_X1 U6070 ( .A1(n5289), .A2(n5293), .ZN(n9976) );
  OAI21_X1 U6071 ( .B1(n5704), .B2(n5292), .A(n5290), .ZN(n9975) );
  NAND2_X1 U6072 ( .A1(n6295), .A2(n6294), .ZN(n10086) );
  NAND2_X1 U6073 ( .A1(n10017), .A2(n6292), .ZN(n10000) );
  NAND2_X1 U6074 ( .A1(n9090), .A2(n9519), .ZN(n10025) );
  NAND2_X1 U6075 ( .A1(n5547), .A2(n5550), .ZN(n8972) );
  NAND2_X1 U6076 ( .A1(n5549), .A2(n5548), .ZN(n5547) );
  NAND2_X1 U6077 ( .A1(n8403), .A2(n9494), .ZN(n8957) );
  OAI21_X1 U6078 ( .B1(n8197), .B2(n5700), .A(n5697), .ZN(n8409) );
  NAND2_X1 U6079 ( .A1(n8192), .A2(n9484), .ZN(n8424) );
  NAND2_X1 U6080 ( .A1(n5346), .A2(n6194), .ZN(n11123) );
  NAND2_X1 U6081 ( .A1(n7588), .A2(n6172), .ZN(n5346) );
  NAND2_X1 U6082 ( .A1(n6174), .A2(n6173), .ZN(n9472) );
  INV_X1 U6083 ( .A(n5712), .ZN(n8216) );
  AND2_X1 U6084 ( .A1(n6165), .A2(n6164), .ZN(n11063) );
  NAND2_X1 U6085 ( .A1(n5711), .A2(n6155), .ZN(n8206) );
  NAND2_X1 U6086 ( .A1(n8235), .A2(n9452), .ZN(n8242) );
  INV_X1 U6087 ( .A(n6142), .ZN(n8243) );
  NAND2_X1 U6088 ( .A1(n11015), .A2(n11014), .ZN(n10012) );
  NAND2_X1 U6089 ( .A1(n10998), .A2(n6118), .ZN(n8237) );
  INV_X1 U6090 ( .A(n10030), .ZN(n10015) );
  OR2_X1 U6091 ( .A1(n11179), .A2(n8191), .ZN(n11007) );
  NAND2_X1 U6092 ( .A1(n7524), .A2(n8191), .ZN(n11010) );
  NAND2_X1 U6093 ( .A1(n7990), .A2(n7989), .ZN(n7994) );
  INV_X1 U6094 ( .A(n11010), .ZN(n10028) );
  OR2_X1 U6095 ( .A1(n7994), .A2(n11007), .ZN(n10030) );
  INV_X1 U6096 ( .A(n9424), .ZN(n9418) );
  AND2_X1 U6097 ( .A1(n6405), .A2(n6404), .ZN(n10118) );
  AOI21_X1 U6098 ( .B1(n9054), .B2(n6172), .A(n6371), .ZN(n10126) );
  INV_X1 U6099 ( .A(n9432), .ZN(n10130) );
  INV_X1 U6100 ( .A(n9553), .ZN(n10134) );
  INV_X1 U6101 ( .A(n9539), .ZN(n10143) );
  NAND2_X1 U6102 ( .A1(n6285), .A2(n6284), .ZN(n10151) );
  INV_X1 U6103 ( .A(n9201), .ZN(n10161) );
  AND2_X2 U6104 ( .A1(n6491), .A2(n7539), .ZN(n11191) );
  INV_X1 U6105 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5963) );
  INV_X1 U6106 ( .A(n5968), .ZN(n10176) );
  XNOR2_X1 U6107 ( .A(n5757), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9112) );
  OR2_X1 U6108 ( .A1(n5783), .A2(n5782), .ZN(n5756) );
  INV_X1 U6109 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8505) );
  INV_X1 U6110 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8379) );
  INV_X1 U6111 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8385) );
  INV_X1 U6112 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8062) );
  INV_X1 U6113 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8010) );
  INV_X1 U6114 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7723) );
  INV_X1 U6115 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7655) );
  NOR2_X1 U6116 ( .A1(n7530), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10169) );
  NAND2_X1 U6117 ( .A1(n5826), .A2(n5586), .ZN(n5585) );
  AOI21_X1 U6118 ( .B1(n5821), .B2(n5587), .A(n5584), .ZN(n5583) );
  NOR2_X1 U6119 ( .A1(n5821), .A2(n5587), .ZN(n5586) );
  AND2_X1 U6120 ( .A1(n7998), .A2(n8001), .ZN(n7262) );
  NAND2_X1 U6121 ( .A1(n7553), .A2(n6690), .ZN(n5509) );
  NAND2_X1 U6122 ( .A1(n5498), .A2(n5503), .ZN(n10188) );
  NAND2_X1 U6123 ( .A1(n10212), .A2(n5504), .ZN(n5498) );
  AND2_X1 U6124 ( .A1(n7709), .A2(n7217), .ZN(n7686) );
  NAND2_X1 U6125 ( .A1(n7394), .A2(n7393), .ZN(n10196) );
  NAND2_X1 U6126 ( .A1(n5490), .A2(n5491), .ZN(n10206) );
  NAND2_X1 U6127 ( .A1(n6567), .A2(n6566), .ZN(n10637) );
  NAND2_X1 U6128 ( .A1(n10180), .A2(n7416), .ZN(n10247) );
  INV_X1 U6129 ( .A(n9222), .ZN(n10284) );
  OAI21_X1 U6130 ( .B1(n10212), .B2(n5502), .A(n5499), .ZN(n7385) );
  INV_X1 U6131 ( .A(n10550), .ZN(n10271) );
  AND2_X1 U6132 ( .A1(n7478), .A2(n10580), .ZN(n10318) );
  AND2_X1 U6133 ( .A1(n7346), .A2(n7348), .ZN(n5471) );
  NOR2_X2 U6134 ( .A1(n7473), .A2(n7462), .ZN(n10308) );
  NAND2_X1 U6135 ( .A1(n7089), .A2(n7019), .ZN(n7088) );
  AOI21_X1 U6136 ( .B1(n5747), .B2(n7474), .A(n8507), .ZN(n7158) );
  OAI21_X1 U6137 ( .B1(n10589), .B2(n6971), .A(n6584), .ZN(n11235) );
  NAND2_X1 U6138 ( .A1(n7626), .A2(n7612), .ZN(n10922) );
  INV_X1 U6139 ( .A(n9325), .ZN(n10607) );
  AND2_X1 U6140 ( .A1(n10461), .A2(n5423), .ZN(n9324) );
  NOR2_X1 U6141 ( .A1(n5424), .A2(n10443), .ZN(n5423) );
  INV_X1 U6142 ( .A(n5425), .ZN(n5424) );
  AOI21_X1 U6143 ( .B1(n9304), .B2(n11232), .A(n9303), .ZN(n10615) );
  INV_X1 U6144 ( .A(n9302), .ZN(n9303) );
  NAND2_X1 U6145 ( .A1(n6557), .A2(n6556), .ZN(n10632) );
  OAI21_X1 U6146 ( .B1(n10517), .B2(n5635), .A(n5633), .ZN(n10477) );
  NAND2_X1 U6147 ( .A1(n5514), .A2(n5515), .ZN(n10500) );
  NOR2_X1 U6148 ( .A1(n5638), .A2(n5637), .ZN(n10491) );
  INV_X1 U6149 ( .A(n9311), .ZN(n5637) );
  NAND2_X1 U6150 ( .A1(n5656), .A2(n5142), .ZN(n10552) );
  AND2_X1 U6151 ( .A1(n5656), .A2(n5229), .ZN(n10554) );
  NAND2_X1 U6152 ( .A1(n6894), .A2(n6893), .ZN(n10652) );
  NAND2_X1 U6153 ( .A1(n5629), .A2(n9142), .ZN(n11200) );
  NOR2_X1 U6154 ( .A1(n7742), .A2(n10599), .ZN(n10560) );
  OR2_X1 U6155 ( .A1(n6657), .A2(n7558), .ZN(n6659) );
  INV_X1 U6156 ( .A(n11254), .ZN(n11218) );
  INV_X1 U6157 ( .A(n10560), .ZN(n11253) );
  NAND2_X1 U6158 ( .A1(n7639), .A2(n7636), .ZN(n10580) );
  INV_X1 U6159 ( .A(n10534), .ZN(n11245) );
  AND2_X2 U6160 ( .A1(n8932), .A2(n8931), .ZN(n11276) );
  AND2_X2 U6161 ( .A1(n8932), .A2(n7641), .ZN(n11280) );
  INV_X1 U6162 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10688) );
  XNOR2_X1 U6163 ( .A(n6515), .B(n6514), .ZN(n10694) );
  OAI21_X1 U6164 ( .B1(n6981), .B2(n6980), .A(n6512), .ZN(n6515) );
  NAND2_X1 U6165 ( .A1(n5456), .A2(n5455), .ZN(n6530) );
  NAND2_X1 U6166 ( .A1(n8908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6167 ( .A1(n5457), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5456) );
  XNOR2_X1 U6168 ( .A(n7175), .B(n8904), .ZN(n9220) );
  INV_X1 U6169 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9111) );
  OR2_X1 U6170 ( .A1(n7163), .A2(n7161), .ZN(n7162) );
  INV_X1 U6171 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U6172 ( .A1(n5351), .A2(n5356), .ZN(n6349) );
  OR2_X1 U6173 ( .A1(n6059), .A2(n5358), .ZN(n5351) );
  INV_X1 U6174 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8383) );
  INV_X1 U6175 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8823) );
  XNOR2_X1 U6176 ( .A(n6323), .B(n6322), .ZN(n8384) );
  NOR2_X1 U6177 ( .A1(n7532), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10693) );
  INV_X1 U6178 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8280) );
  AND2_X1 U6179 ( .A1(n6588), .A2(n6587), .ZN(n10859) );
  NAND2_X1 U6180 ( .A1(n6665), .A2(n5652), .ZN(n6781) );
  AND2_X1 U6181 ( .A1(n6752), .A2(n6741), .ZN(n10928) );
  INV_X1 U6182 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U6183 ( .A1(n7532), .A2(P1_U3086), .ZN(n10696) );
  INV_X1 U6184 ( .A(n5852), .ZN(n8359) );
  INV_X1 U6185 ( .A(n5539), .ZN(n9116) );
  OR2_X1 U6186 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  AOI21_X1 U6187 ( .B1(n5415), .B2(n5906), .A(n5207), .ZN(n5524) );
  XNOR2_X1 U6188 ( .A(n5905), .B(n5939), .ZN(n5415) );
  NOR2_X1 U6189 ( .A1(n11187), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U6190 ( .A1(n7190), .A2(n11187), .ZN(n7195) );
  MUX2_X1 U6191 ( .A(n10054), .B(n10119), .S(n11187), .Z(n10055) );
  NOR2_X1 U6192 ( .A1(n11191), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5702) );
  NOR2_X1 U6193 ( .A1(n5737), .A2(n6492), .ZN(n6493) );
  MUX2_X1 U6194 ( .A(n10120), .B(n10119), .S(n11191), .Z(n10121) );
  INV_X1 U6195 ( .A(n7481), .ZN(n7482) );
  AND2_X1 U6196 ( .A1(n5785), .A2(n5784), .ZN(n5139) );
  AND2_X1 U6197 ( .A1(n5200), .A2(n5168), .ZN(n5140) );
  AND2_X1 U6198 ( .A1(n5366), .A2(n5177), .ZN(n5141) );
  NOR2_X1 U6199 ( .A1(n5518), .A2(n5350), .ZN(n5517) );
  AND2_X1 U6200 ( .A1(n10553), .A2(n5229), .ZN(n5142) );
  INV_X1 U6201 ( .A(n9402), .ZN(n9570) );
  NOR2_X1 U6202 ( .A1(n7375), .A2(n7374), .ZN(n5143) );
  NAND2_X1 U6203 ( .A1(n8267), .A2(n5185), .ZN(n5144) );
  OR2_X1 U6204 ( .A1(n11063), .A2(n9281), .ZN(n5145) );
  NAND2_X1 U6205 ( .A1(n6984), .A2(n6983), .ZN(n10443) );
  INV_X1 U6206 ( .A(n10443), .ZN(n5448) );
  AND3_X1 U6207 ( .A1(n10047), .A2(n10045), .A3(n11187), .ZN(n5146) );
  INV_X1 U6208 ( .A(n10501), .ZN(n5513) );
  INV_X1 U6209 ( .A(n9294), .ZN(n5516) );
  NAND2_X1 U6210 ( .A1(n6431), .A2(n6430), .ZN(n9785) );
  AND3_X1 U6211 ( .A1(n5786), .A2(n5962), .A3(n5139), .ZN(n5147) );
  AND2_X1 U6212 ( .A1(n6079), .A2(n6078), .ZN(n9943) );
  INV_X1 U6213 ( .A(n9943), .ZN(n5319) );
  NAND2_X1 U6214 ( .A1(n9310), .A2(n10511), .ZN(n10515) );
  INV_X1 U6215 ( .A(n5552), .ZN(n5548) );
  OR2_X1 U6216 ( .A1(n5553), .A2(n8956), .ZN(n5552) );
  OR2_X1 U6217 ( .A1(n5567), .A2(n6455), .ZN(n5148) );
  AND2_X1 U6218 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5149) );
  NOR2_X1 U6219 ( .A1(n10072), .A2(n9955), .ZN(n5150) );
  AND2_X1 U6220 ( .A1(n5418), .A2(n5417), .ZN(n5151) );
  AND2_X1 U6221 ( .A1(n5173), .A2(n5700), .ZN(n5152) );
  AND2_X1 U6222 ( .A1(n8995), .A2(n9799), .ZN(n5153) );
  NAND2_X1 U6223 ( .A1(n5487), .A2(n5236), .ZN(n5154) );
  AND2_X1 U6224 ( .A1(n6452), .A2(n6454), .ZN(n5155) );
  OR2_X1 U6225 ( .A1(n9619), .A2(n8387), .ZN(n5156) );
  INV_X2 U6226 ( .A(n6985), .ZN(n6949) );
  AND2_X1 U6227 ( .A1(n7595), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6228 ( .A1(n9006), .A2(n11147), .ZN(n5158) );
  AND2_X1 U6229 ( .A1(n5246), .A2(n9027), .ZN(n5159) );
  NAND2_X1 U6230 ( .A1(n6953), .A2(n6952), .ZN(n10618) );
  INV_X1 U6231 ( .A(n10939), .ZN(n5272) );
  INV_X1 U6232 ( .A(n5470), .ZN(n9110) );
  NAND2_X1 U6233 ( .A1(n5392), .A2(n5528), .ZN(n7820) );
  INV_X2 U6234 ( .A(n6525), .ZN(n7530) );
  OR2_X1 U6235 ( .A1(n9839), .A2(n5900), .ZN(n5161) );
  OR2_X1 U6236 ( .A1(n9805), .A2(n11035), .ZN(n5162) );
  NAND2_X1 U6237 ( .A1(n10306), .A2(n7348), .ZN(n10212) );
  OR2_X1 U6238 ( .A1(n5831), .A2(n6151), .ZN(n5163) );
  NAND2_X1 U6239 ( .A1(n9804), .A2(n9286), .ZN(n5164) );
  XNOR2_X1 U6240 ( .A(n9373), .B(n9655), .ZN(n5165) );
  INV_X1 U6241 ( .A(n5582), .ZN(n6126) );
  NAND2_X1 U6242 ( .A1(n5585), .A2(n5583), .ZN(n5582) );
  NAND2_X1 U6243 ( .A1(n11104), .A2(n9801), .ZN(n5166) );
  NOR2_X1 U6244 ( .A1(n10267), .A2(n10264), .ZN(n10179) );
  NOR2_X1 U6245 ( .A1(n9605), .A2(n5313), .ZN(n5312) );
  AND2_X1 U6246 ( .A1(n5490), .A2(n5488), .ZN(n5167) );
  NOR2_X1 U6247 ( .A1(n6270), .A2(n5608), .ZN(n5607) );
  AND4_X1 U6248 ( .A1(n6545), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n5168)
         );
  AOI21_X1 U6249 ( .B1(n5604), .B2(n5371), .A(n5370), .ZN(n5369) );
  AND2_X1 U6250 ( .A1(n10479), .A2(n5632), .ZN(n5169) );
  OR4_X1 U6251 ( .A1(n6827), .A2(n7123), .A3(n7122), .A4(n6949), .ZN(n5170) );
  INV_X1 U6252 ( .A(n5409), .ZN(n5405) );
  OR2_X1 U6253 ( .A1(n5891), .A2(n5410), .ZN(n5409) );
  AND2_X1 U6254 ( .A1(n6655), .A2(n8861), .ZN(n6665) );
  AND2_X1 U6255 ( .A1(n6613), .A2(n5627), .ZN(n5171) );
  OR2_X1 U6256 ( .A1(n9882), .A2(n5902), .ZN(n5172) );
  AND2_X1 U6257 ( .A1(n8226), .A2(n6181), .ZN(n9595) );
  INV_X1 U6258 ( .A(n9595), .ZN(n8217) );
  BUF_X1 U6259 ( .A(n6958), .Z(n6973) );
  NAND2_X1 U6260 ( .A1(n5557), .A2(n9570), .ZN(n9656) );
  OR2_X1 U6261 ( .A1(n11143), .A2(n9798), .ZN(n5173) );
  AND2_X1 U6262 ( .A1(n9774), .A2(n9770), .ZN(n5174) );
  NAND2_X1 U6263 ( .A1(n6579), .A2(n6578), .ZN(n10602) );
  OR2_X1 U6264 ( .A1(n6737), .A2(n5733), .ZN(n5175) );
  AND2_X1 U6265 ( .A1(n9294), .A2(n6946), .ZN(n10516) );
  INV_X1 U6266 ( .A(n10516), .ZN(n10511) );
  NAND2_X1 U6267 ( .A1(n5675), .A2(n9356), .ZN(n9360) );
  NAND2_X1 U6268 ( .A1(n8051), .A2(n7730), .ZN(n8047) );
  AND3_X1 U6269 ( .A1(n6653), .A2(n6652), .A3(n6651), .ZN(n5176) );
  NOR2_X1 U6270 ( .A1(n6304), .A2(n6052), .ZN(n5177) );
  NOR2_X1 U6271 ( .A1(n7376), .A2(n10278), .ZN(n5178) );
  OR2_X1 U6272 ( .A1(n9806), .A2(n11027), .ZN(n9452) );
  NAND2_X1 U6273 ( .A1(n6906), .A2(n6905), .ZN(n10646) );
  NOR2_X1 U6274 ( .A1(n8369), .A2(n5157), .ZN(n5179) );
  NAND2_X2 U6275 ( .A1(n6530), .A2(n10691), .ZN(n10698) );
  INV_X1 U6276 ( .A(n10698), .ZN(n5624) );
  NAND2_X1 U6277 ( .A1(n6837), .A2(n6836), .ZN(n10290) );
  AND2_X1 U6278 ( .A1(n7532), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5180) );
  AND2_X1 U6279 ( .A1(n5278), .A2(n5277), .ZN(n5181) );
  INV_X1 U6280 ( .A(n5634), .ZN(n5633) );
  OAI21_X1 U6281 ( .B1(n9312), .B2(n9311), .A(n5199), .ZN(n5634) );
  AND2_X1 U6282 ( .A1(n6620), .A2(n5180), .ZN(n5182) );
  INV_X1 U6283 ( .A(n9423), .ZN(n10114) );
  INV_X1 U6284 ( .A(n8480), .ZN(n11168) );
  NAND2_X1 U6285 ( .A1(n6770), .A2(n6769), .ZN(n8480) );
  OAI21_X1 U6286 ( .B1(n6978), .B2(n10443), .A(n5444), .ZN(n5443) );
  INV_X1 U6287 ( .A(n6246), .ZN(n5315) );
  NOR2_X1 U6288 ( .A1(n5593), .A2(n5384), .ZN(n5383) );
  INV_X1 U6289 ( .A(n5673), .ZN(n5672) );
  OAI21_X1 U6290 ( .B1(n5174), .B2(n5674), .A(n9672), .ZN(n5673) );
  INV_X1 U6291 ( .A(n5446), .ZN(n5445) );
  OAI21_X1 U6292 ( .B1(n6978), .B2(n5448), .A(n5447), .ZN(n5446) );
  NAND2_X1 U6293 ( .A1(n8941), .A2(n8940), .ZN(n5183) );
  AND2_X1 U6294 ( .A1(n5430), .A2(n5437), .ZN(n5184) );
  NAND2_X1 U6295 ( .A1(n8302), .A2(n8304), .ZN(n5185) );
  INV_X1 U6296 ( .A(n10582), .ZN(n10658) );
  NAND2_X1 U6297 ( .A1(n6879), .A2(n6878), .ZN(n10582) );
  AND2_X1 U6298 ( .A1(n9620), .A2(n5156), .ZN(n5186) );
  OR2_X1 U6299 ( .A1(n5406), .A2(n8200), .ZN(n5187) );
  AND2_X1 U6300 ( .A1(n9932), .A2(n10126), .ZN(n5188) );
  AND2_X1 U6301 ( .A1(n5450), .A2(n5448), .ZN(n5189) );
  AND2_X1 U6302 ( .A1(n8473), .A2(n8498), .ZN(n7046) );
  OR2_X1 U6303 ( .A1(n5672), .A2(n5165), .ZN(n5190) );
  AND2_X1 U6304 ( .A1(n10086), .A2(n9791), .ZN(n5191) );
  AND3_X1 U6305 ( .A1(n10047), .A2(n11191), .A3(n10045), .ZN(n5192) );
  AND2_X1 U6306 ( .A1(n9548), .A2(n9547), .ZN(n5193) );
  AND2_X1 U6307 ( .A1(n6996), .A2(n6998), .ZN(n5194) );
  AND2_X1 U6308 ( .A1(n5514), .A2(n5512), .ZN(n5195) );
  INV_X1 U6309 ( .A(n10515), .ZN(n5638) );
  OR2_X1 U6310 ( .A1(n5776), .A2(n5756), .ZN(n5196) );
  NOR2_X1 U6311 ( .A1(n9657), .A2(n9893), .ZN(n5581) );
  AND2_X1 U6312 ( .A1(n5379), .A2(n5378), .ZN(n5197) );
  INV_X1 U6313 ( .A(n9519), .ZN(n5568) );
  INV_X1 U6314 ( .A(n9786), .ZN(n9908) );
  NAND2_X1 U6315 ( .A1(n6417), .A2(n6416), .ZN(n9786) );
  OR2_X1 U6316 ( .A1(n10118), .A2(n9908), .ZN(n5198) );
  OR2_X1 U6317 ( .A1(n10495), .A2(n10483), .ZN(n5199) );
  AND2_X1 U6318 ( .A1(n6547), .A2(n5646), .ZN(n5200) );
  AND2_X1 U6319 ( .A1(n9919), .A2(n9561), .ZN(n5201) );
  AND2_X1 U6320 ( .A1(n9515), .A2(n5307), .ZN(n5202) );
  AND2_X1 U6321 ( .A1(n6012), .A2(SI_10_), .ZN(n5203) );
  INV_X1 U6322 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5766) );
  INV_X1 U6323 ( .A(n9977), .ZN(n9981) );
  AND2_X1 U6324 ( .A1(n6334), .A2(n6333), .ZN(n9977) );
  NAND2_X1 U6325 ( .A1(n9351), .A2(n5319), .ZN(n5204) );
  INV_X1 U6326 ( .A(n5571), .ZN(n5570) );
  NAND2_X1 U6327 ( .A1(n6456), .A2(n9971), .ZN(n5571) );
  NAND2_X1 U6328 ( .A1(n9348), .A2(n9702), .ZN(n9705) );
  AND2_X1 U6329 ( .A1(n6118), .A2(n5728), .ZN(n5205) );
  NAND2_X1 U6330 ( .A1(n7329), .A2(n7333), .ZN(n5206) );
  INV_X1 U6331 ( .A(n5602), .ZN(n5601) );
  NAND2_X1 U6332 ( .A1(n5603), .A2(n6023), .ZN(n5602) );
  AND2_X1 U6333 ( .A1(n5271), .A2(n5265), .ZN(n5207) );
  NAND2_X1 U6334 ( .A1(n9740), .A2(n9741), .ZN(n9700) );
  AND2_X1 U6335 ( .A1(n9534), .A2(n9535), .ZN(n9995) );
  NOR2_X1 U6336 ( .A1(n9502), .A2(n9795), .ZN(n5554) );
  AND2_X1 U6337 ( .A1(n9372), .A2(n9786), .ZN(n5208) );
  NAND2_X1 U6338 ( .A1(n6848), .A2(n6847), .ZN(n10669) );
  INV_X1 U6339 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8908) );
  AND2_X1 U6340 ( .A1(n5722), .A2(n9365), .ZN(n5209) );
  OR2_X1 U6341 ( .A1(n6166), .A2(n5710), .ZN(n5210) );
  INV_X1 U6342 ( .A(n5435), .ZN(n5434) );
  NAND2_X1 U6343 ( .A1(n5439), .A2(n5436), .ZN(n5435) );
  INV_X1 U6344 ( .A(n9572), .ZN(n5344) );
  INV_X1 U6345 ( .A(n9658), .ZN(n5339) );
  OR2_X1 U6346 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5211) );
  OR2_X1 U6347 ( .A1(n9325), .A2(n7015), .ZN(n5212) );
  OR2_X1 U6348 ( .A1(n8450), .A2(n5179), .ZN(n5213) );
  AND2_X1 U6349 ( .A1(n5381), .A2(n5385), .ZN(n5214) );
  AND3_X1 U6350 ( .A1(n5810), .A2(n5808), .A3(n5833), .ZN(n5215) );
  AND2_X1 U6351 ( .A1(n5420), .A2(n5419), .ZN(n5216) );
  AND2_X1 U6352 ( .A1(n7871), .A2(n5410), .ZN(n5217) );
  AND2_X1 U6353 ( .A1(n9657), .A2(n9785), .ZN(n5218) );
  NAND2_X1 U6354 ( .A1(n9141), .A2(n11210), .ZN(n5219) );
  OR2_X1 U6355 ( .A1(n11139), .A2(n8410), .ZN(n5220) );
  INV_X1 U6356 ( .A(n8226), .ZN(n5306) );
  AND2_X1 U6357 ( .A1(n5517), .A2(n9295), .ZN(n5221) );
  AND2_X1 U6358 ( .A1(n9514), .A2(n6257), .ZN(n8973) );
  OR2_X1 U6359 ( .A1(n5342), .A2(n5343), .ZN(n5222) );
  AND2_X1 U6360 ( .A1(n9980), .A2(n6456), .ZN(n5223) );
  AND2_X1 U6361 ( .A1(n5355), .A2(n6063), .ZN(n5224) );
  NAND2_X1 U6362 ( .A1(n9576), .A2(n5579), .ZN(n5225) );
  INV_X1 U6363 ( .A(n9522), .ZN(n5337) );
  AND2_X1 U6364 ( .A1(n5565), .A2(n5161), .ZN(n5226) );
  NAND2_X1 U6365 ( .A1(n9576), .A2(n5580), .ZN(n5227) );
  AND2_X1 U6366 ( .A1(n5145), .A2(n5164), .ZN(n5228) );
  INV_X1 U6367 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5962) );
  AOI21_X1 U6368 ( .B1(n5378), .B2(n9298), .A(n9299), .ZN(n5377) );
  NAND2_X1 U6369 ( .A1(n10582), .A2(n10550), .ZN(n5229) );
  INV_X1 U6370 ( .A(n8946), .ZN(n7053) );
  OR2_X1 U6371 ( .A1(n9075), .A2(n9074), .ZN(n9160) );
  AND2_X1 U6372 ( .A1(n9160), .A2(n9159), .ZN(n5230) );
  OAI21_X1 U6373 ( .B1(n8958), .B2(n5308), .A(n5202), .ZN(n9061) );
  AND4_X1 U6374 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n8410)
         );
  NAND2_X1 U6375 ( .A1(n10577), .A2(n5422), .ZN(n5231) );
  AND2_X1 U6376 ( .A1(n10598), .A2(n5429), .ZN(n5232) );
  INV_X1 U6377 ( .A(n8410), .ZN(n9799) );
  NAND2_X1 U6378 ( .A1(n6424), .A2(n6423), .ZN(n9657) );
  OR2_X1 U6379 ( .A1(n7423), .A2(n7422), .ZN(n5233) );
  INV_X1 U6380 ( .A(n9494), .ZN(n5553) );
  AOI21_X1 U6381 ( .B1(n10212), .B2(n7361), .A(n5143), .ZN(n10280) );
  AND2_X1 U6382 ( .A1(n11143), .A2(n9798), .ZN(n5234) );
  NOR2_X1 U6383 ( .A1(n5853), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5806) );
  OR2_X1 U6384 ( .A1(n5948), .A2(n5940), .ZN(n5235) );
  NAND2_X1 U6385 ( .A1(n8980), .A2(n7318), .ZN(n9044) );
  INV_X1 U6386 ( .A(n9006), .ZN(n5532) );
  NOR2_X1 U6387 ( .A1(n10205), .A2(n5489), .ZN(n5488) );
  NOR2_X1 U6388 ( .A1(n10295), .A2(n10296), .ZN(n5236) );
  NOR2_X1 U6389 ( .A1(n11203), .A2(n7337), .ZN(n10598) );
  INV_X1 U6390 ( .A(n9580), .ZN(n9574) );
  NOR2_X1 U6391 ( .A1(n9491), .A2(n9580), .ZN(n5237) );
  OR2_X1 U6392 ( .A1(n5925), .A2(n7568), .ZN(n5238) );
  OR2_X1 U6393 ( .A1(n11260), .A2(n10286), .ZN(n7129) );
  INV_X1 U6394 ( .A(n7129), .ZN(n5523) );
  OR2_X1 U6395 ( .A1(n5924), .A2(n7837), .ZN(n5239) );
  AND2_X1 U6396 ( .A1(n5539), .A2(n5538), .ZN(n5240) );
  NAND2_X1 U6397 ( .A1(n6967), .A2(n6966), .ZN(n10614) );
  OR2_X1 U6398 ( .A1(n10642), .A2(n10506), .ZN(n9294) );
  INV_X1 U6399 ( .A(n9351), .ZN(n10138) );
  NAND2_X1 U6400 ( .A1(n6083), .A2(n6082), .ZN(n9351) );
  INV_X1 U6401 ( .A(n5494), .ZN(n5493) );
  NAND2_X1 U6402 ( .A1(n5233), .A2(n7416), .ZN(n5494) );
  NOR2_X1 U6403 ( .A1(n6052), .A2(n6051), .ZN(n5241) );
  OR2_X1 U6404 ( .A1(n5793), .A2(n5769), .ZN(n5242) );
  NOR2_X1 U6405 ( .A1(n10652), .A2(n10570), .ZN(n5243) );
  AND2_X1 U6406 ( .A1(n6024), .A2(SI_13_), .ZN(n5244) );
  NAND2_X1 U6407 ( .A1(n9090), .A2(n5567), .ZN(n5245) );
  AND2_X1 U6408 ( .A1(n5661), .A2(n8410), .ZN(n5246) );
  INV_X1 U6409 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5771) );
  NOR2_X1 U6410 ( .A1(n9118), .A2(n5898), .ZN(n5247) );
  NAND2_X1 U6411 ( .A1(n6802), .A2(n6801), .ZN(n9141) );
  AND2_X1 U6412 ( .A1(n10010), .A2(n9529), .ZN(n5248) );
  AND2_X1 U6413 ( .A1(n5856), .A2(n5855), .ZN(n8450) );
  INV_X1 U6414 ( .A(n8450), .ZN(n5391) );
  XNOR2_X1 U6415 ( .A(n5870), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U6416 ( .A1(n9580), .A2(n7521), .ZN(n11003) );
  NAND2_X1 U6417 ( .A1(n5712), .A2(n9595), .ZN(n8214) );
  AND2_X1 U6418 ( .A1(n5475), .A2(n5479), .ZN(n5249) );
  INV_X1 U6419 ( .A(n10041), .ZN(n11000) );
  AND2_X1 U6420 ( .A1(n8334), .A2(n5151), .ZN(n5250) );
  AND2_X1 U6421 ( .A1(n7170), .A2(n7169), .ZN(n5470) );
  INV_X1 U6422 ( .A(n9857), .ZN(n8012) );
  OR2_X1 U6423 ( .A1(n9618), .A2(n5135), .ZN(n7484) );
  NAND2_X1 U6424 ( .A1(n8197), .A2(n6203), .ZN(n8420) );
  INV_X1 U6425 ( .A(n9191), .ZN(n5682) );
  NOR2_X1 U6426 ( .A1(n5859), .A2(n8436), .ZN(n5251) );
  OR2_X1 U6427 ( .A1(n8064), .A2(n5935), .ZN(n5252) );
  NOR2_X1 U6428 ( .A1(n7876), .A2(n7875), .ZN(n5253) );
  AND2_X1 U6429 ( .A1(n6381), .A2(SI_25_), .ZN(n5254) );
  NAND3_X1 U6430 ( .A1(n5474), .A2(n7280), .A3(n5473), .ZN(n9384) );
  AND2_X2 U6431 ( .A1(n7189), .A2(n7188), .ZN(n11187) );
  OR2_X1 U6432 ( .A1(n9857), .A2(n5564), .ZN(n5255) );
  AND2_X1 U6433 ( .A1(n10599), .A2(n8381), .ZN(n6985) );
  NAND2_X1 U6434 ( .A1(n6786), .A2(n6785), .ZN(n9043) );
  INV_X1 U6435 ( .A(n9043), .ZN(n5417) );
  XNOR2_X1 U6436 ( .A(n6432), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9618) );
  INV_X1 U6437 ( .A(n9618), .ZN(n8387) );
  NAND2_X1 U6438 ( .A1(n9220), .A2(n7649), .ZN(n10505) );
  INV_X1 U6439 ( .A(n10505), .ZN(n11237) );
  AOI21_X1 U6440 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8088) );
  NAND2_X1 U6441 ( .A1(n5497), .A2(n5496), .ZN(n7709) );
  INV_X1 U6442 ( .A(n7869), .ZN(n5401) );
  INV_X1 U6443 ( .A(n7474), .ZN(n7647) );
  NAND2_X1 U6444 ( .A1(n7092), .A2(n7091), .ZN(n7474) );
  XNOR2_X1 U6445 ( .A(n5897), .B(n9130), .ZN(n9120) );
  NOR2_X1 U6446 ( .A1(n9130), .A2(n5860), .ZN(n5861) );
  NOR2_X2 U6447 ( .A1(n9825), .A2(n5864), .ZN(n9853) );
  NAND2_X1 U6448 ( .A1(n5535), .A2(n5844), .ZN(n5534) );
  NAND2_X1 U6449 ( .A1(n5859), .A2(n5532), .ZN(n5531) );
  INV_X2 U6450 ( .A(n5814), .ZN(n5284) );
  XNOR2_X1 U6451 ( .A(n5262), .B(n6151), .ZN(n7759) );
  XNOR2_X1 U6452 ( .A(n5846), .B(n8153), .ZN(n8142) );
  NAND2_X1 U6453 ( .A1(n5258), .A2(n10624), .ZN(n10677) );
  INV_X1 U6454 ( .A(n10623), .ZN(n5258) );
  NOR2_X1 U6455 ( .A1(n9290), .A2(n9289), .ZN(n10569) );
  XNOR2_X1 U6456 ( .A(n7098), .B(n9260), .ZN(n9253) );
  NAND2_X2 U6457 ( .A1(n6619), .A2(n5259), .ZN(n9260) );
  NOR2_X1 U6458 ( .A1(n6620), .A2(n7614), .ZN(n5260) );
  AOI21_X2 U6459 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7724), .A(n9817), .ZN(
        n5863) );
  NOR2_X1 U6460 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  INV_X1 U6461 ( .A(n5584), .ZN(n5264) );
  NAND3_X1 U6462 ( .A1(n5282), .A2(n5791), .A3(n5211), .ZN(n5873) );
  INV_X2 U6463 ( .A(n5944), .ZN(n9623) );
  MUX2_X1 U6464 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n5944), .Z(n5919) );
  NAND2_X1 U6465 ( .A1(n5284), .A2(n5820), .ZN(n5826) );
  NAND2_X1 U6466 ( .A1(n5284), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6467 ( .A1(n5284), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5877) );
  NAND3_X1 U6468 ( .A1(n6115), .A2(n6112), .A3(n5285), .ZN(n9807) );
  NAND2_X1 U6469 ( .A1(n5704), .A2(n5290), .ZN(n5286) );
  NAND2_X1 U6470 ( .A1(n5286), .A2(n5287), .ZN(n9964) );
  NOR2_X1 U6471 ( .A1(n10052), .A2(n5299), .ZN(n10119) );
  NAND2_X1 U6472 ( .A1(n5708), .A2(n5303), .ZN(n5302) );
  NAND2_X1 U6473 ( .A1(n5304), .A2(n5302), .ZN(n8194) );
  NAND4_X1 U6474 ( .A1(n5332), .A2(n5248), .A3(n5334), .A4(n5335), .ZN(n9533)
         );
  NAND3_X1 U6475 ( .A1(n5332), .A2(n5335), .A3(n5334), .ZN(n9527) );
  NOR2_X1 U6476 ( .A1(n5345), .A2(n5344), .ZN(n5342) );
  NAND2_X1 U6477 ( .A1(n9573), .A2(n5222), .ZN(n5340) );
  NAND2_X1 U6478 ( .A1(n6059), .A2(n5356), .ZN(n5354) );
  NAND2_X1 U6479 ( .A1(n6059), .A2(n5359), .ZN(n5355) );
  NAND2_X1 U6480 ( .A1(n6259), .A2(n5141), .ZN(n5361) );
  NOR2_X1 U6481 ( .A1(n5373), .A2(n5374), .ZN(n9300) );
  NOR2_X1 U6482 ( .A1(n10468), .A2(n10467), .ZN(n10470) );
  OR2_X2 U6483 ( .A1(n10470), .A2(n9298), .ZN(n5379) );
  NAND2_X1 U6484 ( .A1(n5380), .A2(n5214), .ZN(n6019) );
  INV_X1 U6485 ( .A(n5591), .ZN(n5382) );
  NAND3_X1 U6486 ( .A1(n5584), .A2(n5215), .A3(n5754), .ZN(n5693) );
  NAND3_X1 U6487 ( .A1(n5388), .A2(n5390), .A3(P2_REG2_REG_11__SCAN_IN), .ZN(
        n5575) );
  OR2_X1 U6488 ( .A1(n8369), .A2(n5389), .ZN(n5388) );
  OR2_X1 U6489 ( .A1(n5157), .A2(n5391), .ZN(n5389) );
  OAI21_X1 U6490 ( .B1(n8369), .B2(n5157), .A(n5391), .ZN(n5390) );
  NAND2_X1 U6491 ( .A1(n7820), .A2(n5398), .ZN(n7758) );
  NAND2_X1 U6492 ( .A1(n7870), .A2(n5217), .ZN(n5407) );
  AND2_X1 U6493 ( .A1(n7870), .A2(n7871), .ZN(n7869) );
  INV_X1 U6494 ( .A(n5400), .ZN(n8143) );
  NAND3_X1 U6495 ( .A1(n5407), .A2(n5408), .A3(n5404), .ZN(n8144) );
  AND3_X2 U6496 ( .A1(n5826), .A2(n5822), .A3(n5823), .ZN(n6107) );
  NAND2_X2 U6497 ( .A1(n6620), .A2(n7532), .ZN(n6982) );
  NAND2_X2 U6498 ( .A1(n6524), .A2(n6523), .ZN(n6620) );
  NAND2_X1 U6499 ( .A1(n5416), .A2(n8334), .ZN(n11203) );
  NAND2_X1 U6500 ( .A1(n10461), .A2(n5425), .ZN(n10438) );
  NAND2_X1 U6501 ( .A1(n10461), .A2(n10449), .ZN(n10448) );
  NOR2_X1 U6502 ( .A1(n6990), .A2(n5212), .ZN(n5439) );
  INV_X1 U6503 ( .A(n9313), .ZN(n5450) );
  AOI21_X1 U6504 ( .B1(n5454), .B2(n5451), .A(n6664), .ZN(n6687) );
  NAND3_X1 U6505 ( .A1(n6521), .A2(n5657), .A3(n5140), .ZN(n5458) );
  AOI21_X1 U6506 ( .B1(n5462), .B2(n6997), .A(n8946), .ZN(n6826) );
  NAND2_X2 U6507 ( .A1(n7171), .A2(n5470), .ZN(n7579) );
  NAND2_X1 U6508 ( .A1(n7449), .A2(n5470), .ZN(n7574) );
  NAND3_X1 U6509 ( .A1(n7346), .A2(n10307), .A3(n7348), .ZN(n10306) );
  OAI21_X1 U6510 ( .B1(n10307), .B2(n5471), .A(n10306), .ZN(n10309) );
  AND2_X2 U6511 ( .A1(n10197), .A2(n7409), .ZN(n10263) );
  NAND2_X1 U6512 ( .A1(n8039), .A2(n5476), .ZN(n5474) );
  INV_X1 U6513 ( .A(n5479), .ZN(n5478) );
  OR2_X1 U6514 ( .A1(n8040), .A2(n8041), .ZN(n5480) );
  OAI21_X1 U6515 ( .B1(n7317), .B2(n5485), .A(n5483), .ZN(n9045) );
  NAND2_X1 U6516 ( .A1(n7317), .A2(n5483), .ZN(n5482) );
  INV_X1 U6517 ( .A(n10180), .ZN(n5486) );
  INV_X1 U6518 ( .A(n7215), .ZN(n5496) );
  NAND2_X1 U6519 ( .A1(n5505), .A2(n7047), .ZN(n7049) );
  NAND2_X1 U6520 ( .A1(n5505), .A2(n8327), .ZN(n8328) );
  OAI21_X1 U6521 ( .B1(n8129), .B2(n8130), .A(n5505), .ZN(n8131) );
  XNOR2_X2 U6522 ( .A(n5993), .B(n5992), .ZN(n6152) );
  NOR2_X2 U6523 ( .A1(n10478), .A2(n9297), .ZN(n10468) );
  NAND2_X1 U6524 ( .A1(n10536), .A2(n5221), .ZN(n5511) );
  AND3_X2 U6525 ( .A1(n5519), .A2(n5520), .A3(n9180), .ZN(n9181) );
  NAND2_X1 U6526 ( .A1(n11230), .A2(n5521), .ZN(n5519) );
  NAND2_X1 U6527 ( .A1(n5520), .A2(n5519), .ZN(n9183) );
  NAND2_X1 U6528 ( .A1(n7045), .A2(n7044), .ZN(n8129) );
  NOR2_X1 U6529 ( .A1(n10480), .A2(n10479), .ZN(n10478) );
  NAND2_X1 U6530 ( .A1(n5991), .A2(n5990), .ZN(n5993) );
  OR2_X1 U6531 ( .A1(n6657), .A2(n7563), .ZN(n6619) );
  NAND2_X1 U6532 ( .A1(n6634), .A2(n5744), .ZN(n7910) );
  NOR2_X1 U6533 ( .A1(n8071), .A2(n7027), .ZN(n7028) );
  AND2_X1 U6534 ( .A1(n6517), .A2(n6520), .ZN(n5648) );
  AND3_X1 U6535 ( .A1(n6518), .A2(n6519), .A3(n8873), .ZN(n5649) );
  NAND2_X1 U6536 ( .A1(n5590), .A2(n6011), .ZN(n6205) );
  NAND2_X2 U6537 ( .A1(n6531), .A2(n10698), .ZN(n6625) );
  NAND2_X1 U6538 ( .A1(n5983), .A2(n5982), .ZN(n6124) );
  NAND2_X1 U6539 ( .A1(n7052), .A2(n7118), .ZN(n8945) );
  NAND2_X1 U6540 ( .A1(n5987), .A2(n5986), .ZN(n6135) );
  NAND2_X2 U6541 ( .A1(n7108), .A2(n7033), .ZN(n8096) );
  NAND2_X2 U6542 ( .A1(n6668), .A2(n6667), .ZN(n10230) );
  NAND2_X1 U6543 ( .A1(n6106), .A2(n6105), .ZN(n5983) );
  NAND2_X1 U6544 ( .A1(n7343), .A2(n7342), .ZN(n7346) );
  OAI211_X2 U6545 ( .C1(n7644), .C2(n7196), .A(n7579), .B(n7934), .ZN(n9637)
         );
  NAND2_X1 U6546 ( .A1(n5525), .A2(n5524), .ZN(P2_U3201) );
  NAND2_X1 U6547 ( .A1(n5526), .A2(n5874), .ZN(n5525) );
  XNOR2_X1 U6548 ( .A(n5527), .B(n5871), .ZN(n5526) );
  INV_X1 U6549 ( .A(n6151), .ZN(n5528) );
  OAI21_X2 U6550 ( .B1(n7795), .B2(n5534), .A(n5533), .ZN(n5846) );
  NAND2_X1 U6551 ( .A1(n5861), .A2(n5540), .ZN(n5536) );
  NAND2_X1 U6552 ( .A1(n8405), .A2(n5546), .ZN(n5544) );
  NAND2_X1 U6553 ( .A1(n9899), .A2(n5558), .ZN(n5556) );
  NAND2_X1 U6554 ( .A1(n9899), .A2(n6462), .ZN(n5557) );
  INV_X1 U6555 ( .A(n5565), .ZN(n9827) );
  NAND2_X1 U6556 ( .A1(n6453), .A2(n5155), .ZN(n5566) );
  NAND2_X1 U6557 ( .A1(n7803), .A2(n5888), .ZN(n7870) );
  OAI21_X2 U6558 ( .B1(n9982), .B2(n5571), .A(n5569), .ZN(n9957) );
  NAND2_X1 U6559 ( .A1(n8192), .A2(n5572), .ZN(n6450) );
  NOR2_X1 U6560 ( .A1(n5574), .A2(n5573), .ZN(n5572) );
  INV_X1 U6561 ( .A(n9484), .ZN(n5573) );
  INV_X1 U6562 ( .A(n5162), .ZN(n5577) );
  OAI21_X1 U6563 ( .B1(n9406), .B2(n5227), .A(n5578), .ZN(n9429) );
  XNOR2_X2 U6564 ( .A(n5965), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5967) );
  NAND3_X1 U6565 ( .A1(n10176), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n5967), .ZN(
        n5589) );
  NAND2_X1 U6566 ( .A1(n6193), .A2(n5742), .ZN(n5590) );
  NAND2_X1 U6567 ( .A1(n5988), .A2(n5977), .ZN(n6089) );
  OAI21_X1 U6568 ( .B1(n6225), .B2(n6022), .A(n6021), .ZN(n6237) );
  NAND2_X1 U6569 ( .A1(n6259), .A2(n6030), .ZN(n5609) );
  NAND2_X1 U6570 ( .A1(n6369), .A2(n6368), .ZN(n5615) );
  INV_X1 U6571 ( .A(n5994), .ZN(n5617) );
  NAND2_X2 U6572 ( .A1(n5625), .A2(n5624), .ZN(n6649) );
  NAND2_X1 U6573 ( .A1(n5629), .A2(n5628), .ZN(n11202) );
  NOR2_X2 U6574 ( .A1(n5641), .A2(n5640), .ZN(n9147) );
  OR2_X1 U6575 ( .A1(n5641), .A2(n11248), .ZN(n11259) );
  NAND4_X1 U6576 ( .A1(n6518), .A2(n6520), .A3(n6519), .A4(n6517), .ZN(n5653)
         );
  NAND2_X1 U6577 ( .A1(n6655), .A2(n5650), .ZN(n5647) );
  NAND4_X1 U6578 ( .A1(n5649), .A2(n6655), .A3(n5648), .A4(n5650), .ZN(n6535)
         );
  NAND2_X1 U6579 ( .A1(n10574), .A2(n5142), .ZN(n5655) );
  INV_X1 U6580 ( .A(n5656), .ZN(n10573) );
  NAND2_X1 U6581 ( .A1(n6521), .A2(n5140), .ZN(n7169) );
  NAND3_X1 U6582 ( .A1(n6521), .A2(n5140), .A3(n5658), .ZN(n6529) );
  INV_X1 U6583 ( .A(n9253), .ZN(n7004) );
  NAND2_X1 U6584 ( .A1(n7902), .A2(n7004), .ZN(n9251) );
  OR2_X1 U6585 ( .A1(n8996), .A2(n5153), .ZN(n5659) );
  NAND2_X1 U6586 ( .A1(n5659), .A2(n5660), .ZN(n9029) );
  NAND2_X1 U6587 ( .A1(n9705), .A2(n5662), .ZN(n9751) );
  NAND2_X1 U6588 ( .A1(n9771), .A2(n5668), .ZN(n5664) );
  OAI211_X1 U6589 ( .C1(n9771), .C2(n5669), .A(n5664), .B(n5665), .ZN(n9379)
         );
  NAND2_X1 U6590 ( .A1(n9771), .A2(n5174), .ZN(n9772) );
  INV_X1 U6591 ( .A(n9358), .ZN(n5675) );
  NAND2_X1 U6592 ( .A1(n5676), .A2(n5677), .ZN(n9204) );
  NAND2_X1 U6593 ( .A1(n5684), .A2(n5683), .ZN(n9344) );
  OAI21_X1 U6594 ( .B1(n8107), .B2(n5144), .A(n5685), .ZN(n8990) );
  INV_X1 U6595 ( .A(n5793), .ZN(n5689) );
  OAI21_X1 U6596 ( .B1(n5793), .B2(n5691), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5870) );
  OAI21_X1 U6597 ( .B1(n5689), .B2(n5821), .A(n5690), .ZN(n5772) );
  INV_X2 U6598 ( .A(n5693), .ZN(n5790) );
  NAND2_X1 U6599 ( .A1(n8197), .A2(n5695), .ZN(n5694) );
  NAND2_X1 U6600 ( .A1(n5694), .A2(n5696), .ZN(n8400) );
  AOI21_X1 U6601 ( .B1(n5146), .B2(n10046), .A(n5701), .ZN(P2_U3488) );
  AOI21_X1 U6602 ( .B1(n5192), .B2(n10046), .A(n5702), .ZN(P2_U3456) );
  NAND3_X1 U6603 ( .A1(n6144), .A2(n6143), .A3(n5228), .ZN(n5708) );
  NAND3_X1 U6604 ( .A1(n6144), .A2(n6143), .A3(n5164), .ZN(n5711) );
  NAND2_X1 U6605 ( .A1(n6144), .A2(n6143), .ZN(n9278) );
  OAI21_X1 U6606 ( .B1(n9907), .B2(n6396), .A(n9365), .ZN(n9892) );
  NAND2_X1 U6607 ( .A1(n5714), .A2(n5713), .ZN(n9654) );
  NOR2_X1 U6608 ( .A1(n5716), .A2(n5218), .ZN(n5713) );
  NAND2_X1 U6609 ( .A1(n9907), .A2(n5718), .ZN(n5714) );
  NAND2_X1 U6610 ( .A1(n9907), .A2(n5209), .ZN(n5715) );
  AND2_X1 U6611 ( .A1(n5209), .A2(n9652), .ZN(n5718) );
  NAND2_X1 U6612 ( .A1(n5791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  NAND3_X1 U6613 ( .A1(n10176), .A2(P2_REG2_REG_1__SCAN_IN), .A3(n5967), .ZN(
        n5723) );
  NAND4_X2 U6614 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n5723), .ZN(n6103)
         );
  NAND2_X1 U6615 ( .A1(n5726), .A2(n5725), .ZN(n6141) );
  NAND2_X1 U6616 ( .A1(n5788), .A2(n5790), .ZN(n5776) );
  NAND2_X1 U6617 ( .A1(n6432), .A2(n5773), .ZN(n5774) );
  XNOR2_X1 U6618 ( .A(n5979), .B(SI_1_), .ZN(n6096) );
  OAI21_X1 U6619 ( .B1(n5988), .B2(n5978), .A(n6089), .ZN(n5979) );
  NAND2_X1 U6620 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  OAI222_X1 U6621 ( .A1(P2_U3151), .A2(n10176), .B1(n10175), .B2(n10699), .C1(
        n10174), .C2(n10173), .ZN(P2_U3266) );
  NOR2_X2 U6622 ( .A1(n9181), .A2(n7135), .ZN(n9290) );
  OR2_X1 U6623 ( .A1(n6736), .A2(n6999), .ZN(n5733) );
  INV_X1 U6624 ( .A(n9384), .ZN(n9385) );
  XOR2_X1 U6625 ( .A(n5136), .B(P2_REG1_REG_19__SCAN_IN), .Z(n5734) );
  NOR2_X1 U6626 ( .A1(n9405), .A2(n10103), .ZN(n7192) );
  INV_X1 U6627 ( .A(n11003), .ZN(n10003) );
  OR2_X1 U6628 ( .A1(n7179), .A2(n7178), .ZN(n5735) );
  INV_X2 U6629 ( .A(n11244), .ZN(n10600) );
  OR2_X1 U6630 ( .A1(n9318), .A2(n10272), .ZN(n5736) );
  NOR2_X1 U6631 ( .A1(n11191), .A2(n6490), .ZN(n5737) );
  INV_X1 U6632 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7161) );
  AND2_X1 U6633 ( .A1(n7295), .A2(n7293), .ZN(n5738) );
  AND2_X1 U6634 ( .A1(n6001), .A2(n6000), .ZN(n5739) );
  INV_X1 U6635 ( .A(n10967), .ZN(n5874) );
  AND3_X1 U6636 ( .A1(n9692), .A2(n9336), .A3(n9691), .ZN(n5740) );
  OR2_X1 U6637 ( .A1(n10462), .A2(n10318), .ZN(n5741) );
  AND2_X1 U6638 ( .A1(n6011), .A2(n6010), .ZN(n5742) );
  NAND2_X1 U6639 ( .A1(n10038), .A2(n9419), .ZN(n5743) );
  INV_X1 U6640 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5820) );
  INV_X2 U6641 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U6642 ( .A1(n10336), .A2(n7936), .ZN(n5744) );
  INV_X1 U6643 ( .A(n9456), .ZN(n6444) );
  NAND2_X1 U6644 ( .A1(n8936), .A2(n8935), .ZN(n5745) );
  AND3_X1 U6645 ( .A1(n7247), .A2(n7246), .A3(n7975), .ZN(n5746) );
  NAND2_X1 U6646 ( .A1(n6422), .A2(n6421), .ZN(n6496) );
  XOR2_X1 U6647 ( .A(n7155), .B(n7172), .Z(n5747) );
  INV_X1 U6648 ( .A(n9465), .ZN(n6447) );
  MUX2_X1 U6649 ( .A(P2_U3893), .B(n5946), .S(n5872), .Z(n9881) );
  INV_X1 U6650 ( .A(n9881), .ZN(n5947) );
  NAND2_X2 U6651 ( .A1(n7994), .A2(n11010), .ZN(n11015) );
  NOR2_X1 U6652 ( .A1(n9405), .A2(n10160), .ZN(n6492) );
  INV_X1 U6653 ( .A(n10646), .ZN(n9318) );
  AND2_X1 U6654 ( .A1(n7003), .A2(n8047), .ZN(n6660) );
  AND2_X1 U6655 ( .A1(n7103), .A2(n6949), .ZN(n6664) );
  AOI211_X1 U6656 ( .C1(n6704), .C2(n7108), .A(n7000), .B(n7034), .ZN(n6706)
         );
  AND2_X1 U6657 ( .A1(n7118), .A2(n7050), .ZN(n6825) );
  OAI211_X1 U6658 ( .C1(n6829), .C2(n6828), .A(n11234), .B(n5170), .ZN(n6830)
         );
  NOR3_X1 U6659 ( .A1(n6934), .A2(n6933), .A3(n10511), .ZN(n6947) );
  OR2_X1 U6660 ( .A1(n9043), .A2(n10325), .ZN(n8936) );
  INV_X1 U6661 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6662 ( .B1(n6964), .B2(n10455), .A(n6963), .ZN(n6979) );
  INV_X1 U6663 ( .A(n7034), .ZN(n7035) );
  OR4_X1 U6664 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n7455) );
  INV_X1 U6665 ( .A(n7485), .ZN(n7483) );
  AND2_X1 U6666 ( .A1(n9420), .A2(n5743), .ZN(n9421) );
  INV_X1 U6667 ( .A(n5890), .ZN(n5891) );
  OR2_X1 U6668 ( .A1(n9432), .A2(n9789), .ZN(n6365) );
  OR2_X1 U6669 ( .A1(n8314), .A2(n8313), .ZN(n7279) );
  NOR2_X1 U6670 ( .A1(n10602), .A2(n10242), .ZN(n7122) );
  NOR2_X1 U6671 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  INV_X1 U6672 ( .A(n9357), .ZN(n9356) );
  INV_X1 U6673 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8794) );
  INV_X1 U6674 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9727) );
  INV_X1 U6675 ( .A(n9425), .ZN(n9426) );
  AND2_X1 U6676 ( .A1(n10945), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5825) );
  NOR2_X1 U6677 ( .A1(n9873), .A2(n9872), .ZN(n9875) );
  AND2_X1 U6678 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  OR2_X1 U6679 ( .A1(n6274), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6286) );
  OR2_X1 U6680 ( .A1(n7538), .A2(n6481), .ZN(n7185) );
  NAND2_X1 U6681 ( .A1(n9439), .A2(n9445), .ZN(n6442) );
  AND2_X1 U6682 ( .A1(n9382), .A2(n7279), .ZN(n7280) );
  AND2_X1 U6683 ( .A1(n6897), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6909) );
  OR2_X1 U6684 ( .A1(n10396), .A2(n10395), .ZN(n10855) );
  OR2_X1 U6685 ( .A1(n10409), .A2(n10408), .ZN(n10874) );
  AND2_X1 U6686 ( .A1(n6909), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6570) );
  INV_X1 U6687 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6716) );
  XNOR2_X1 U6688 ( .A(n10336), .B(n8925), .ZN(n7922) );
  NAND2_X1 U6689 ( .A1(n8904), .A2(n8903), .ZN(n6527) );
  INV_X1 U6690 ( .A(SI_22_), .ZN(n8711) );
  INV_X1 U6691 ( .A(SI_16_), .ZN(n8722) );
  INV_X1 U6692 ( .A(SI_11_), .ZN(n8737) );
  INV_X1 U6693 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U6694 ( .A1(n7501), .A2(n7500), .ZN(n7786) );
  INV_X1 U6695 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9124) );
  OR2_X1 U6696 ( .A1(n6208), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U6697 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  NOR2_X1 U6698 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U6699 ( .A1(n6372), .A2(n8779), .ZN(n6406) );
  INV_X1 U6700 ( .A(n5160), .ZN(n8260) );
  NOR2_X1 U6701 ( .A1(n9875), .A2(n9874), .ZN(n9876) );
  NAND2_X1 U6702 ( .A1(n6409), .A2(n8764), .ZN(n6425) );
  NOR2_X1 U6703 ( .A1(n9893), .A2(n11003), .ZN(n9894) );
  AND2_X1 U6704 ( .A1(n6483), .A2(n7540), .ZN(n6485) );
  INV_X1 U6705 ( .A(n6454), .ZN(n6455) );
  INV_X1 U6706 ( .A(n8392), .ZN(n9589) );
  NAND2_X1 U6707 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U6708 ( .A1(n7414), .A2(n7415), .ZN(n7416) );
  NAND2_X1 U6709 ( .A1(n7345), .A2(n7344), .ZN(n7348) );
  NOR2_X1 U6710 ( .A1(n6849), .A2(n10257), .ZN(n6883) );
  AND2_X1 U6711 ( .A1(n6744), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6757) );
  INV_X1 U6712 ( .A(n6620), .ZN(n6630) );
  OR2_X1 U6713 ( .A1(n10839), .A2(n10838), .ZN(n10841) );
  OR2_X1 U6714 ( .A1(n10874), .A2(n10873), .ZN(n10876) );
  OR2_X1 U6715 ( .A1(n10893), .A2(n10414), .ZN(n10894) );
  NOR2_X1 U6716 ( .A1(n10504), .A2(n10507), .ZN(n10472) );
  NOR2_X1 U6717 ( .A1(n9260), .A2(n9259), .ZN(n9263) );
  AOI22_X1 U6718 ( .A1(n10322), .A2(n11236), .B1(n9327), .B2(n10320), .ZN(
        n9302) );
  INV_X1 U6719 ( .A(n10618), .ZN(n10449) );
  INV_X1 U6720 ( .A(n6859), .ZN(n7060) );
  INV_X1 U6721 ( .A(n7046), .ZN(n8327) );
  NAND2_X1 U6722 ( .A1(n7200), .A2(n7196), .ZN(n7911) );
  INV_X1 U6723 ( .A(SI_25_), .ZN(n8518) );
  NAND2_X1 U6724 ( .A1(n7092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U6725 ( .A1(n6318), .A2(n6317), .ZN(n6320) );
  OR2_X1 U6726 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6536) );
  INV_X1 U6727 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8872) );
  OR2_X1 U6728 ( .A1(n6251), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U6729 ( .A1(n6339), .A2(n8778), .ZN(n6342) );
  NAND2_X1 U6730 ( .A1(n6356), .A2(n6355), .ZN(n6373) );
  AND2_X1 U6731 ( .A1(n6484), .A2(n7983), .ZN(n7519) );
  NAND2_X1 U6732 ( .A1(n5959), .A2(n5958), .ZN(n6326) );
  OR2_X1 U6733 ( .A1(n6218), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6228) );
  OR2_X1 U6734 ( .A1(n6296), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U6735 ( .A1(n6092), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U6736 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  NOR2_X1 U6737 ( .A1(n5866), .A2(n9860), .ZN(n10966) );
  INV_X1 U6738 ( .A(n9785), .ZN(n9893) );
  NOR2_X1 U6739 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  INV_X1 U6740 ( .A(n9474), .ZN(n6448) );
  INV_X1 U6741 ( .A(n6485), .ZN(n7983) );
  OR2_X1 U6742 ( .A1(n9887), .A2(n9886), .ZN(n10110) );
  INV_X1 U6743 ( .A(n9797), .ZN(n9495) );
  INV_X1 U6744 ( .A(n9801), .ZN(n8304) );
  NAND2_X1 U6745 ( .A1(n9384), .A2(n5738), .ZN(n8465) );
  INV_X1 U6746 ( .A(n10195), .ZN(n7405) );
  INV_X1 U6747 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7629) );
  AND2_X1 U6748 ( .A1(n7228), .A2(n7226), .ZN(n7710) );
  OR2_X1 U6749 ( .A1(n6649), .A2(n10451), .ZN(n6960) );
  NAND2_X1 U6750 ( .A1(n6838), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6851) );
  AOI21_X1 U6751 ( .B1(n10322), .B2(n11237), .A(n10472), .ZN(n10473) );
  NAND2_X1 U6752 ( .A1(n10642), .A2(n10541), .ZN(n9311) );
  INV_X1 U6753 ( .A(n10566), .ZN(n10575) );
  NAND2_X1 U6754 ( .A1(n7971), .A2(n6690), .ZN(n6579) );
  AND2_X1 U6755 ( .A1(n7639), .A2(n7638), .ZN(n8929) );
  INV_X1 U6756 ( .A(n11232), .ZN(n10503) );
  AND2_X1 U6757 ( .A1(n6421), .A2(n6403), .ZN(n6419) );
  INV_X1 U6758 ( .A(n9779), .ZN(n9766) );
  AND2_X1 U6759 ( .A1(n6364), .A2(n6363), .ZN(n9944) );
  AND3_X1 U6760 ( .A1(n6314), .A2(n6313), .A3(n6312), .ZN(n9744) );
  AND4_X1 U6761 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9070)
         );
  INV_X1 U6762 ( .A(n9873), .ZN(n10959) );
  OR2_X1 U6763 ( .A1(n9425), .A2(n6465), .ZN(n10041) );
  AOI21_X1 U6764 ( .B1(n8205), .B2(n8204), .A(n6447), .ZN(n8213) );
  INV_X1 U6765 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8763) );
  INV_X1 U6766 ( .A(n10012), .ZN(n10033) );
  NOR2_X1 U6767 ( .A1(n11179), .A2(n7514), .ZN(n7524) );
  INV_X1 U6768 ( .A(n11179), .ZN(n11158) );
  INV_X1 U6769 ( .A(n11181), .ZN(n11159) );
  NAND2_X1 U6770 ( .A1(n6469), .A2(n9112), .ZN(n7538) );
  INV_X1 U6771 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5802) );
  INV_X1 U6772 ( .A(n10318), .ZN(n10289) );
  INV_X1 U6773 ( .A(n10300), .ZN(n10315) );
  AND4_X1 U6774 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n10471)
         );
  INV_X1 U6775 ( .A(n10922), .ZN(n10895) );
  INV_X1 U6776 ( .A(n10918), .ZN(n10846) );
  AND2_X1 U6777 ( .A1(n6993), .A2(n6992), .ZN(n9180) );
  OR2_X1 U6778 ( .A1(n11244), .A2(n7743), .ZN(n10534) );
  AND2_X1 U6779 ( .A1(n8930), .A2(n8929), .ZN(n8931) );
  NAND2_X1 U6780 ( .A1(n7644), .A2(n7744), .ZN(n11269) );
  AND2_X1 U6781 ( .A1(n11202), .A2(n11201), .ZN(n11219) );
  INV_X1 U6782 ( .A(n10671), .ZN(n11273) );
  NOR2_X1 U6783 ( .A1(n7640), .A2(n8930), .ZN(n7641) );
  XNOR2_X1 U6784 ( .A(n7157), .B(n8677), .ZN(n7580) );
  AND2_X1 U6785 ( .A1(n6712), .A2(n6766), .ZN(n10813) );
  OR2_X1 U6786 ( .A1(n7509), .A2(n8503), .ZN(n5941) );
  OR2_X1 U6787 ( .A1(n7522), .A2(n7520), .ZN(n9754) );
  NAND2_X1 U6788 ( .A1(n7497), .A2(n7496), .ZN(n9748) );
  AND2_X1 U6789 ( .A1(n8264), .A2(n8255), .ZN(n9887) );
  INV_X1 U6790 ( .A(n10961), .ZN(n9792) );
  INV_X1 U6791 ( .A(n8425), .ZN(n9800) );
  OR2_X1 U6792 ( .A1(n7701), .A2(n9623), .ZN(n10972) );
  OR2_X1 U6793 ( .A1(n7701), .A2(n5944), .ZN(n10967) );
  AOI21_X1 U6794 ( .B1(n6440), .B2(n10041), .A(n6439), .ZN(n9400) );
  NOR2_X1 U6795 ( .A1(n7193), .A2(n7192), .ZN(n7194) );
  NAND2_X1 U6796 ( .A1(n11187), .A2(n11158), .ZN(n10103) );
  INV_X1 U6797 ( .A(n11187), .ZN(n11185) );
  NAND2_X1 U6798 ( .A1(n6491), .A2(n7524), .ZN(n10160) );
  INV_X1 U6799 ( .A(n11191), .ZN(n11188) );
  AND2_X1 U6800 ( .A1(n7508), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7545) );
  NAND2_X1 U6801 ( .A1(n7539), .A2(n7538), .ZN(n7549) );
  INV_X1 U6802 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9040) );
  INV_X1 U6803 ( .A(n10962), .ZN(n10956) );
  NAND2_X1 U6804 ( .A1(n7532), .A2(P2_U3151), .ZN(n10175) );
  INV_X2 U6805 ( .A(n10169), .ZN(n10173) );
  INV_X1 U6806 ( .A(n10602), .ZN(n11224) );
  INV_X1 U6807 ( .A(n10308), .ZN(n10292) );
  OR2_X1 U6808 ( .A1(n6823), .A2(n6822), .ZN(n10595) );
  OR2_X1 U6809 ( .A1(n7585), .A2(n7584), .ZN(n10933) );
  INV_X1 U6810 ( .A(n10600), .ZN(n11258) );
  NAND2_X1 U6811 ( .A1(n10600), .A2(n7935), .ZN(n11254) );
  AND2_X1 U6812 ( .A1(n7742), .A2(n10580), .ZN(n11244) );
  INV_X1 U6813 ( .A(n11276), .ZN(n11275) );
  INV_X1 U6814 ( .A(n11280), .ZN(n11277) );
  AND2_X1 U6815 ( .A1(n9110), .A2(n9025), .ZN(n7576) );
  INV_X1 U6816 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8630) );
  NOR2_X2 U6817 ( .A1(n5941), .A2(P2_U3151), .ZN(P2_U3893) );
  NAND2_X1 U6818 ( .A1(n7195), .A2(n7194), .ZN(P2_U3487) );
  NAND2_X1 U6819 ( .A1(n6494), .A2(n6493), .ZN(P2_U3455) );
  NOR2_X1 U6820 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5752) );
  NAND2_X1 U6821 ( .A1(n5759), .A2(n5755), .ZN(n5782) );
  NAND2_X1 U6822 ( .A1(n5196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6823 ( .A1(n5762), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U6824 ( .A1(n5760), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5761) );
  NAND3_X1 U6825 ( .A1(n9112), .A2(n6482), .A3(n9039), .ZN(n7509) );
  NAND2_X1 U6826 ( .A1(n5763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  INV_X1 U6827 ( .A(n7508), .ZN(n8503) );
  NAND2_X1 U6828 ( .A1(n5806), .A2(n5767), .ZN(n5804) );
  NOR2_X2 U6829 ( .A1(n5804), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6830 ( .A1(n5801), .A2(n5802), .ZN(n5793) );
  NAND3_X1 U6831 ( .A1(n5796), .A2(n5794), .A3(n5768), .ZN(n5769) );
  XNOR2_X2 U6832 ( .A(n5775), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U6833 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U6834 ( .A1(n9580), .A2(n7508), .ZN(n5778) );
  NAND2_X1 U6835 ( .A1(n5778), .A2(n5941), .ZN(n5945) );
  XNOR2_X2 U6836 ( .A(n5787), .B(n5962), .ZN(n5872) );
  OR2_X1 U6837 ( .A1(n5945), .A2(n6307), .ZN(n5792) );
  NAND2_X1 U6838 ( .A1(n5792), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U6839 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6840 ( .A1(n5800), .A2(n5794), .ZN(n5795) );
  NAND2_X1 U6841 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U6842 ( .A1(n5799), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U6843 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U6844 ( .A(n5798), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U6845 ( .A(n5799), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9857) );
  XNOR2_X1 U6846 ( .A(n5800), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9839) );
  OR2_X1 U6847 ( .A1(n5801), .A2(n5821), .ZN(n5803) );
  XNOR2_X1 U6848 ( .A(n5803), .B(n5802), .ZN(n7724) );
  NAND2_X1 U6849 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5805) );
  XNOR2_X1 U6850 ( .A(n5805), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U6851 ( .A1(n5855), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U6852 ( .A(n5807), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9020) );
  INV_X1 U6853 ( .A(n9020), .ZN(n7696) );
  NAND2_X1 U6854 ( .A1(n5812), .A2(n5808), .ZN(n5809) );
  NAND2_X1 U6855 ( .A1(n5809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U6856 ( .A1(n5830), .A2(n5810), .ZN(n5811) );
  NAND2_X1 U6857 ( .A1(n5811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5834) );
  XNOR2_X1 U6858 ( .A(n5834), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6163) );
  INV_X1 U6859 ( .A(n6163), .ZN(n7837) );
  XNOR2_X1 U6860 ( .A(n5812), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7969) );
  INV_X1 U6861 ( .A(n7969), .ZN(n7559) );
  INV_X1 U6862 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6863 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5813) );
  NAND2_X2 U6864 ( .A1(n5815), .A2(n5814), .ZN(n7901) );
  OAI21_X1 U6865 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n5816), .A(n6100), .ZN(n5817) );
  INV_X1 U6866 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10982) );
  INV_X1 U6867 ( .A(n5818), .ZN(n5819) );
  INV_X1 U6868 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5824) );
  NAND3_X1 U6869 ( .A1(n5814), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  MUX2_X1 U6870 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5824), .S(n6107), .Z(n10935)
         );
  INV_X1 U6871 ( .A(n6107), .ZN(n10945) );
  NOR2_X1 U6872 ( .A1(n10934), .A2(n5825), .ZN(n5827) );
  NOR2_X1 U6873 ( .A1(n5827), .A2(n6126), .ZN(n5828) );
  AOI21_X1 U6874 ( .B1(n5827), .B2(n6126), .A(n5828), .ZN(n7767) );
  NAND2_X1 U6875 ( .A1(n7767), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7766) );
  INV_X1 U6876 ( .A(n5828), .ZN(n7957) );
  INV_X1 U6877 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U6878 ( .A(n7969), .B(n5829), .ZN(n7958) );
  AOI21_X1 U6879 ( .B1(n7766), .B2(n7957), .A(n7958), .ZN(n7960) );
  XNOR2_X1 U6880 ( .A(n5830), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6151) );
  INV_X1 U6881 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5832) );
  MUX2_X1 U6882 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n5832), .S(n6163), .Z(n7829)
         );
  AOI21_X1 U6883 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7837), .A(n7828), .ZN(
        n5836) );
  NAND2_X1 U6884 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  NAND2_X1 U6885 ( .A1(n5835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U6886 ( .A(n5840), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7807) );
  XNOR2_X1 U6887 ( .A(n5836), .B(n7807), .ZN(n7796) );
  INV_X1 U6888 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11091) );
  NOR2_X2 U6889 ( .A1(n7796), .A2(n11091), .ZN(n7795) );
  INV_X1 U6890 ( .A(n5836), .ZN(n5837) );
  INV_X1 U6891 ( .A(n7807), .ZN(n7568) );
  INV_X1 U6892 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6893 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  NAND2_X1 U6894 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  INV_X1 U6895 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5842) );
  XNOR2_X1 U6896 ( .A(n5843), .B(n5842), .ZN(n7573) );
  NAND2_X1 U6897 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7573), .ZN(n5844) );
  OAI21_X1 U6898 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7573), .A(n5844), .ZN(
        n7875) );
  OR2_X1 U6899 ( .A1(n5790), .A2(n5821), .ZN(n5845) );
  XNOR2_X1 U6900 ( .A(n5845), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8153) );
  INV_X1 U6901 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11124) );
  NOR2_X1 U6902 ( .A1(n8153), .A2(n5846), .ZN(n5847) );
  OR2_X1 U6903 ( .A1(n5848), .A2(n5821), .ZN(n5850) );
  XNOR2_X1 U6904 ( .A(n5850), .B(n5849), .ZN(n7595) );
  NAND2_X1 U6905 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7595), .ZN(n5851) );
  OAI21_X1 U6906 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7595), .A(n5851), .ZN(
        n8360) );
  NAND2_X1 U6907 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  MUX2_X1 U6908 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5854), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5856) );
  INV_X1 U6909 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11147) );
  INV_X1 U6910 ( .A(n5857), .ZN(n5858) );
  NOR2_X1 U6911 ( .A1(n8450), .A2(n5858), .ZN(n5859) );
  INV_X1 U6912 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U6913 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9020), .B1(n7696), .B2(
        n11163), .ZN(n9006) );
  AOI21_X2 U6914 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7696), .A(n9005), .ZN(
        n5860) );
  INV_X1 U6915 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U6916 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7724), .ZN(n5862) );
  OAI21_X1 U6917 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7724), .A(n5862), .ZN(
        n9818) );
  NOR2_X1 U6918 ( .A1(n9839), .A2(n5863), .ZN(n5864) );
  INV_X1 U6919 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10101) );
  XNOR2_X1 U6920 ( .A(n5863), .B(n9839), .ZN(n9826) );
  INV_X1 U6921 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10097) );
  AOI22_X1 U6922 ( .A1(n9857), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10097), .B2(
        n8012), .ZN(n9852) );
  NOR2_X1 U6923 ( .A1(n9882), .A2(n5865), .ZN(n5866) );
  INV_X1 U6924 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9862) );
  INV_X1 U6925 ( .A(n9882), .ZN(n8064) );
  NAND2_X1 U6926 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U6927 ( .A(n5867), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U6928 ( .A1(n10956), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U6929 ( .B1(n10956), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5868), .ZN(
        n10965) );
  NOR2_X1 U6930 ( .A1(n10966), .A2(n10965), .ZN(n10964) );
  INV_X1 U6931 ( .A(n10964), .ZN(n5869) );
  INV_X1 U6932 ( .A(n5734), .ZN(n5871) );
  OR2_X1 U6933 ( .A1(n5872), .A2(P2_U3151), .ZN(n9215) );
  OR2_X1 U6934 ( .A1(n5945), .A2(n9215), .ZN(n7701) );
  INV_X1 U6935 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5875) );
  MUX2_X1 U6936 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5875), .S(n5136), .Z(n5939)
         );
  INV_X1 U6937 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11017) );
  INV_X1 U6938 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6091) );
  AND2_X1 U6939 ( .A1(n6091), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5876) );
  INV_X1 U6940 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7889) );
  OR2_X1 U6941 ( .A1(n6107), .A2(n11017), .ZN(n5878) );
  NAND2_X1 U6942 ( .A1(n10947), .A2(n5878), .ZN(n5879) );
  NAND2_X1 U6943 ( .A1(n5879), .A2(n5582), .ZN(n7950) );
  NAND2_X1 U6944 ( .A1(n7950), .A2(n5880), .ZN(n7769) );
  INV_X1 U6945 ( .A(n7769), .ZN(n5881) );
  INV_X1 U6946 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U6947 ( .A1(n5881), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U6948 ( .A1(n7952), .A2(n7950), .ZN(n5882) );
  XNOR2_X1 U6949 ( .A(n7969), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U6950 ( .A1(n5882), .A2(n7949), .ZN(n7954) );
  INV_X1 U6951 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8245) );
  OR2_X1 U6952 ( .A1(n7969), .A2(n8245), .ZN(n5883) );
  INV_X1 U6953 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9284) );
  INV_X1 U6954 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5884) );
  MUX2_X1 U6955 ( .A(n5884), .B(P2_REG2_REG_6__SCAN_IN), .S(n6163), .Z(n7821)
         );
  NAND2_X1 U6956 ( .A1(n5885), .A2(n7821), .ZN(n7823) );
  OR2_X1 U6957 ( .A1(n6163), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U6958 ( .A1(n7823), .A2(n5886), .ZN(n5887) );
  NAND2_X1 U6959 ( .A1(n5887), .A2(n7568), .ZN(n5888) );
  OAI21_X1 U6960 ( .B1(n5887), .B2(n7568), .A(n5888), .ZN(n7801) );
  INV_X1 U6961 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8221) );
  OR2_X1 U6962 ( .A1(n7573), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U6963 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7573), .ZN(n5890) );
  AND2_X1 U6964 ( .A1(n5889), .A2(n5890), .ZN(n7871) );
  NOR2_X1 U6965 ( .A1(n8153), .A2(n5892), .ZN(n5893) );
  INV_X1 U6966 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8200) );
  NOR2_X1 U6967 ( .A1(n5893), .A2(n8143), .ZN(n8371) );
  NAND2_X1 U6968 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7595), .ZN(n5894) );
  OAI21_X1 U6969 ( .B1(n7595), .B2(P2_REG2_REG_10__SCAN_IN), .A(n5894), .ZN(
        n8370) );
  NOR2_X1 U6970 ( .A1(n8371), .A2(n8370), .ZN(n8369) );
  INV_X1 U6971 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8439) );
  INV_X1 U6972 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5895) );
  MUX2_X1 U6973 ( .A(n5895), .B(P2_REG2_REG_12__SCAN_IN), .S(n9020), .Z(n5896)
         );
  INV_X1 U6974 ( .A(n5896), .ZN(n9015) );
  NOR2_X1 U6975 ( .A1(n9016), .A2(n9015), .ZN(n9014) );
  AOI21_X1 U6976 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7696), .A(n9014), .ZN(
        n5897) );
  NOR2_X1 U6977 ( .A1(n9130), .A2(n5897), .ZN(n5898) );
  INV_X1 U6978 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U6979 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7724), .ZN(n5899) );
  OAI21_X1 U6980 ( .B1(n7724), .B2(P2_REG2_REG_14__SCAN_IN), .A(n5899), .ZN(
        n9809) );
  AOI21_X1 U6981 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7724), .A(n9808), .ZN(
        n5900) );
  INV_X1 U6982 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9828) );
  XNOR2_X1 U6983 ( .A(n9839), .B(n5900), .ZN(n9829) );
  NAND2_X1 U6984 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8012), .ZN(n5901) );
  OAI21_X1 U6985 ( .B1(n8012), .B2(P2_REG2_REG_16__SCAN_IN), .A(n5901), .ZN(
        n9843) );
  INV_X1 U6986 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9863) );
  XNOR2_X1 U6987 ( .A(n9882), .B(n5902), .ZN(n9864) );
  NAND2_X1 U6988 ( .A1(n10956), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6989 ( .B1(n10956), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5903), .ZN(
        n10970) );
  INV_X1 U6990 ( .A(n5903), .ZN(n5904) );
  INV_X1 U6991 ( .A(n10972), .ZN(n5906) );
  MUX2_X1 U6992 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9623), .Z(n5935) );
  XNOR2_X1 U6993 ( .A(n9882), .B(n5935), .ZN(n9870) );
  MUX2_X1 U6994 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9623), .Z(n5907) );
  OR2_X1 U6995 ( .A1(n5907), .A2(n8012), .ZN(n5934) );
  XNOR2_X1 U6996 ( .A(n9857), .B(n5907), .ZN(n9846) );
  MUX2_X1 U6997 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9623), .Z(n5909) );
  INV_X1 U6998 ( .A(n5909), .ZN(n5908) );
  NAND2_X1 U6999 ( .A1(n9839), .A2(n5908), .ZN(n5933) );
  XNOR2_X1 U7000 ( .A(n5909), .B(n9839), .ZN(n9832) );
  MUX2_X1 U7001 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9623), .Z(n5910) );
  OR2_X1 U7002 ( .A1(n5910), .A2(n7724), .ZN(n5932) );
  INV_X1 U7003 ( .A(n7724), .ZN(n9822) );
  XNOR2_X1 U7004 ( .A(n5910), .B(n9822), .ZN(n9812) );
  MUX2_X1 U7005 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9623), .Z(n5912) );
  INV_X1 U7006 ( .A(n5912), .ZN(n5911) );
  NAND2_X1 U7007 ( .A1(n9130), .A2(n5911), .ZN(n5931) );
  XNOR2_X1 U7008 ( .A(n5912), .B(n9130), .ZN(n9123) );
  MUX2_X1 U7009 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9623), .Z(n5913) );
  OR2_X1 U7010 ( .A1(n5913), .A2(n7696), .ZN(n5930) );
  XNOR2_X1 U7011 ( .A(n5913), .B(n9020), .ZN(n9009) );
  MUX2_X1 U7012 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9623), .Z(n5914) );
  OR2_X1 U7013 ( .A1(n5914), .A2(n5391), .ZN(n5929) );
  XNOR2_X1 U7014 ( .A(n5914), .B(n8450), .ZN(n8443) );
  MUX2_X1 U7015 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9623), .Z(n5915) );
  OR2_X1 U7016 ( .A1(n5915), .A2(n7595), .ZN(n5928) );
  INV_X1 U7017 ( .A(n7595), .ZN(n8375) );
  XNOR2_X1 U7018 ( .A(n5915), .B(n8375), .ZN(n8364) );
  MUX2_X1 U7019 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9623), .Z(n5917) );
  INV_X1 U7020 ( .A(n5917), .ZN(n5916) );
  NAND2_X1 U7021 ( .A1(n8153), .A2(n5916), .ZN(n5927) );
  XNOR2_X1 U7022 ( .A(n5917), .B(n8153), .ZN(n8147) );
  MUX2_X1 U7023 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9623), .Z(n5918) );
  OR2_X1 U7024 ( .A1(n5918), .A2(n7573), .ZN(n5926) );
  INV_X1 U7025 ( .A(n7573), .ZN(n7872) );
  XNOR2_X1 U7026 ( .A(n5918), .B(n7872), .ZN(n7882) );
  MUX2_X1 U7027 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9623), .Z(n5925) );
  MUX2_X1 U7028 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9623), .Z(n5924) );
  MUX2_X1 U7029 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9623), .Z(n5923) );
  MUX2_X1 U7030 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9623), .Z(n5922) );
  MUX2_X1 U7031 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9623), .Z(n5921) );
  MUX2_X1 U7032 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9623), .Z(n5920) );
  INV_X1 U7033 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7991) );
  MUX2_X1 U7034 ( .A(n7991), .B(n5816), .S(n9623), .Z(n7703) );
  AND2_X1 U7035 ( .A1(n7703), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7892) );
  AOI21_X1 U7036 ( .B1(n5919), .B2(n7901), .A(n7891), .ZN(n10940) );
  XOR2_X1 U7037 ( .A(n6107), .B(n5920), .Z(n10941) );
  NOR2_X1 U7038 ( .A1(n10940), .A2(n10941), .ZN(n10938) );
  AOI21_X1 U7039 ( .B1(n5920), .B2(n10945), .A(n10938), .ZN(n7778) );
  XNOR2_X1 U7040 ( .A(n5921), .B(n6126), .ZN(n7777) );
  NAND2_X1 U7041 ( .A1(n7778), .A2(n7777), .ZN(n7776) );
  OAI21_X1 U7042 ( .B1(n5921), .B2(n5582), .A(n7776), .ZN(n7965) );
  XOR2_X1 U7043 ( .A(n7969), .B(n5922), .Z(n7966) );
  XOR2_X1 U7044 ( .A(n6151), .B(n5923), .Z(n7755) );
  XNOR2_X1 U7045 ( .A(n5924), .B(n6163), .ZN(n7818) );
  NAND2_X1 U7046 ( .A1(n5181), .A2(n7818), .ZN(n7817) );
  XNOR2_X1 U7047 ( .A(n5925), .B(n7807), .ZN(n7798) );
  NAND2_X1 U7048 ( .A1(n5926), .A2(n7881), .ZN(n8146) );
  NAND2_X1 U7049 ( .A1(n8147), .A2(n8146), .ZN(n8145) );
  NAND2_X1 U7050 ( .A1(n5927), .A2(n8145), .ZN(n8363) );
  NAND2_X1 U7051 ( .A1(n8364), .A2(n8363), .ZN(n8362) );
  NAND2_X1 U7052 ( .A1(n5928), .A2(n8362), .ZN(n8442) );
  NAND2_X1 U7053 ( .A1(n8443), .A2(n8442), .ZN(n8441) );
  NAND2_X1 U7054 ( .A1(n5929), .A2(n8441), .ZN(n9008) );
  NAND2_X1 U7055 ( .A1(n9009), .A2(n9008), .ZN(n9007) );
  NAND2_X1 U7056 ( .A1(n5930), .A2(n9007), .ZN(n9122) );
  NAND2_X1 U7057 ( .A1(n9123), .A2(n9122), .ZN(n9121) );
  NAND2_X1 U7058 ( .A1(n5931), .A2(n9121), .ZN(n9811) );
  NAND2_X1 U7059 ( .A1(n9812), .A2(n9811), .ZN(n9810) );
  NAND2_X1 U7060 ( .A1(n5932), .A2(n9810), .ZN(n9831) );
  NAND2_X1 U7061 ( .A1(n9832), .A2(n9831), .ZN(n9830) );
  NAND2_X1 U7062 ( .A1(n5933), .A2(n9830), .ZN(n9845) );
  INV_X1 U7063 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10008) );
  INV_X1 U7064 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5936) );
  MUX2_X1 U7065 ( .A(n10008), .B(n5936), .S(n9623), .Z(n5937) );
  NOR2_X1 U7066 ( .A1(n5938), .A2(n5937), .ZN(n10953) );
  NAND2_X1 U7067 ( .A1(n5938), .A2(n5937), .ZN(n10954) );
  MUX2_X1 U7068 ( .A(n5939), .B(n5734), .S(n9623), .Z(n5940) );
  NAND2_X1 U7069 ( .A1(P2_U3893), .A2(n5872), .ZN(n10939) );
  INV_X1 U7070 ( .A(n5941), .ZN(n5942) );
  INV_X1 U7071 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5958) );
  NOR2_X1 U7072 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5958), .ZN(n9694) );
  AOI21_X1 U7073 ( .B1(n10959), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9694), .ZN(
        n5943) );
  NAND2_X1 U7074 ( .A1(n5944), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9172) );
  NOR2_X1 U7075 ( .A1(n5945), .A2(n9172), .ZN(n5946) );
  NOR2_X1 U7076 ( .A1(n5947), .A2(n5135), .ZN(n5948) );
  INV_X1 U7077 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U7078 ( .A1(n8790), .A2(n8763), .ZN(n6145) );
  INV_X1 U7079 ( .A(n6145), .ZN(n5950) );
  INV_X1 U7080 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7081 ( .A1(n5950), .A2(n5949), .ZN(n6156) );
  INV_X1 U7082 ( .A(n6175), .ZN(n5951) );
  NAND2_X1 U7083 ( .A1(n5951), .A2(n8760), .ZN(n6186) );
  INV_X1 U7084 ( .A(n6195), .ZN(n5952) );
  NAND2_X1 U7085 ( .A1(n5952), .A2(n8585), .ZN(n6208) );
  INV_X1 U7086 ( .A(n6240), .ZN(n5955) );
  NAND2_X1 U7087 ( .A1(n5955), .A2(n9124), .ZN(n6251) );
  INV_X1 U7088 ( .A(n6326), .ZN(n5960) );
  INV_X1 U7089 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8778) );
  OR2_X2 U7090 ( .A1(n6073), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7091 ( .A1(n6073), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7092 ( .A1(n6357), .A2(n5961), .ZN(n9947) );
  INV_X1 U7093 ( .A(n5966), .ZN(n5964) );
  NAND2_X1 U7094 ( .A1(n5964), .A2(n5963), .ZN(n10167) );
  NAND2_X1 U7095 ( .A1(n9947), .A2(n5130), .ZN(n5974) );
  INV_X1 U7096 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7097 ( .A1(n8257), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5970) );
  INV_X1 U7098 ( .A(n5967), .ZN(n9273) );
  NAND2_X1 U7099 ( .A1(n8250), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5969) );
  OAI211_X1 U7100 ( .C1(n5971), .C2(n8260), .A(n5970), .B(n5969), .ZN(n5972)
         );
  INV_X1 U7101 ( .A(n5972), .ZN(n5973) );
  NAND2_X1 U7102 ( .A1(n5974), .A2(n5973), .ZN(n9790) );
  NAND2_X1 U7103 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5978) );
  AND2_X1 U7104 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5977) );
  MUX2_X1 U7105 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5988), .Z(n6097) );
  NAND2_X1 U7106 ( .A1(n5979), .A2(SI_1_), .ZN(n5980) );
  MUX2_X1 U7107 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5988), .Z(n5981) );
  INV_X1 U7108 ( .A(SI_2_), .ZN(n8552) );
  XNOR2_X1 U7109 ( .A(n5981), .B(n8552), .ZN(n6105) );
  NAND2_X1 U7110 ( .A1(n5981), .A2(SI_2_), .ZN(n5982) );
  MUX2_X1 U7111 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5988), .Z(n5985) );
  INV_X1 U7112 ( .A(SI_3_), .ZN(n5984) );
  XNOR2_X1 U7113 ( .A(n5985), .B(n5984), .ZN(n6125) );
  NAND2_X1 U7114 ( .A1(n6124), .A2(n6125), .ZN(n5987) );
  NAND2_X1 U7115 ( .A1(n5985), .A2(SI_3_), .ZN(n5986) );
  MUX2_X1 U7116 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7530), .Z(n5989) );
  INV_X1 U7117 ( .A(SI_4_), .ZN(n8748) );
  XNOR2_X1 U7118 ( .A(n5989), .B(n8748), .ZN(n6136) );
  NAND2_X1 U7119 ( .A1(n6135), .A2(n6136), .ZN(n5991) );
  NAND2_X1 U7120 ( .A1(n5989), .A2(SI_4_), .ZN(n5990) );
  MUX2_X1 U7121 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7530), .Z(n5992) );
  INV_X1 U7122 ( .A(SI_5_), .ZN(n5995) );
  NAND2_X1 U7123 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  MUX2_X1 U7124 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7530), .Z(n5998) );
  XNOR2_X1 U7125 ( .A(n5998), .B(SI_6_), .ZN(n6162) );
  INV_X1 U7126 ( .A(n6162), .ZN(n6167) );
  MUX2_X1 U7127 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7532), .Z(n5999) );
  XNOR2_X1 U7128 ( .A(n5999), .B(SI_7_), .ZN(n6170) );
  INV_X1 U7129 ( .A(n6170), .ZN(n5997) );
  AND2_X1 U7130 ( .A1(n6167), .A2(n5997), .ZN(n5996) );
  NAND2_X1 U7131 ( .A1(n5998), .A2(SI_6_), .ZN(n6169) );
  OR2_X1 U7132 ( .A1(n6170), .A2(n6169), .ZN(n6001) );
  NAND2_X1 U7133 ( .A1(n5999), .A2(SI_7_), .ZN(n6000) );
  INV_X1 U7134 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7571) );
  INV_X4 U7135 ( .A(n6525), .ZN(n7532) );
  MUX2_X1 U7136 ( .A(n8841), .B(n7571), .S(n7532), .Z(n6003) );
  INV_X1 U7137 ( .A(SI_8_), .ZN(n6002) );
  NAND2_X1 U7138 ( .A1(n6003), .A2(n6002), .ZN(n6006) );
  INV_X1 U7139 ( .A(n6003), .ZN(n6004) );
  NAND2_X1 U7140 ( .A1(n6004), .A2(SI_8_), .ZN(n6005) );
  NAND2_X1 U7141 ( .A1(n6006), .A2(n6005), .ZN(n6182) );
  INV_X1 U7142 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6007) );
  MUX2_X1 U7143 ( .A(n8842), .B(n6007), .S(n7532), .Z(n6008) );
  NAND2_X1 U7144 ( .A1(n6008), .A2(n8738), .ZN(n6011) );
  INV_X1 U7145 ( .A(n6008), .ZN(n6009) );
  NAND2_X1 U7146 ( .A1(n6009), .A2(SI_9_), .ZN(n6010) );
  MUX2_X1 U7147 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7532), .Z(n6012) );
  XNOR2_X1 U7148 ( .A(n6012), .B(n8739), .ZN(n6204) );
  INV_X1 U7149 ( .A(n6204), .ZN(n6013) );
  INV_X1 U7150 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6014) );
  MUX2_X1 U7151 ( .A(n6014), .B(n7655), .S(n7532), .Z(n6015) );
  NAND2_X1 U7152 ( .A1(n6015), .A2(n8737), .ZN(n6018) );
  INV_X1 U7153 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7154 ( .A1(n6016), .A2(SI_11_), .ZN(n6017) );
  NAND2_X1 U7155 ( .A1(n6018), .A2(n6017), .ZN(n6214) );
  NAND2_X1 U7156 ( .A1(n6019), .A2(n6018), .ZN(n6225) );
  MUX2_X1 U7157 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n7532), .Z(n6020) );
  XNOR2_X1 U7158 ( .A(n6020), .B(n8733), .ZN(n6224) );
  INV_X1 U7159 ( .A(n6224), .ZN(n6022) );
  NAND2_X1 U7160 ( .A1(n6020), .A2(SI_12_), .ZN(n6021) );
  MUX2_X1 U7161 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n7530), .Z(n6024) );
  XNOR2_X1 U7162 ( .A(n6024), .B(SI_13_), .ZN(n6236) );
  INV_X1 U7163 ( .A(n6236), .ZN(n6023) );
  MUX2_X1 U7164 ( .A(n8630), .B(n7723), .S(n7532), .Z(n6025) );
  NAND2_X1 U7165 ( .A1(n6025), .A2(n8729), .ZN(n6258) );
  INV_X1 U7166 ( .A(n6025), .ZN(n6026) );
  NAND2_X1 U7167 ( .A1(n6026), .A2(SI_14_), .ZN(n6027) );
  NAND2_X1 U7168 ( .A1(n6258), .A2(n6027), .ZN(n6247) );
  INV_X1 U7169 ( .A(n6247), .ZN(n6028) );
  NAND2_X1 U7170 ( .A1(n6029), .A2(n6028), .ZN(n6259) );
  MUX2_X1 U7171 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7532), .Z(n6031) );
  XNOR2_X1 U7172 ( .A(n6031), .B(n8728), .ZN(n6260) );
  AND2_X1 U7173 ( .A1(n6258), .A2(n6260), .ZN(n6030) );
  NAND2_X1 U7174 ( .A1(n6031), .A2(SI_15_), .ZN(n6032) );
  MUX2_X1 U7175 ( .A(n8626), .B(n8010), .S(n7530), .Z(n6033) );
  NAND2_X1 U7176 ( .A1(n6033), .A2(n8722), .ZN(n6036) );
  INV_X1 U7177 ( .A(n6033), .ZN(n6034) );
  NAND2_X1 U7178 ( .A1(n6034), .A2(SI_16_), .ZN(n6035) );
  NAND2_X1 U7179 ( .A1(n6036), .A2(n6035), .ZN(n6270) );
  MUX2_X1 U7180 ( .A(n6037), .B(n8062), .S(n7530), .Z(n6038) );
  NAND2_X1 U7181 ( .A1(n6038), .A2(n8723), .ZN(n6041) );
  INV_X1 U7182 ( .A(n6038), .ZN(n6039) );
  NAND2_X1 U7183 ( .A1(n6039), .A2(SI_17_), .ZN(n6040) );
  MUX2_X1 U7184 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7532), .Z(n6049) );
  XNOR2_X1 U7185 ( .A(n6049), .B(n8721), .ZN(n6293) );
  INV_X1 U7186 ( .A(n6293), .ZN(n6304) );
  MUX2_X1 U7187 ( .A(n8823), .B(n8385), .S(n7530), .Z(n6042) );
  NAND2_X1 U7188 ( .A1(n6042), .A2(n8716), .ZN(n6053) );
  INV_X1 U7189 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U7190 ( .A1(n6043), .A2(SI_20_), .ZN(n6044) );
  NAND2_X1 U7191 ( .A1(n6053), .A2(n6044), .ZN(n6321) );
  INV_X1 U7192 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6045) );
  MUX2_X1 U7193 ( .A(n8280), .B(n6045), .S(n7532), .Z(n6046) );
  NAND2_X1 U7194 ( .A1(n6046), .A2(n8715), .ZN(n6319) );
  NOR2_X1 U7195 ( .A1(n6321), .A2(n6319), .ZN(n6052) );
  INV_X1 U7196 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7197 ( .A1(n6047), .A2(SI_19_), .ZN(n6048) );
  NAND2_X1 U7198 ( .A1(n6319), .A2(n6048), .ZN(n6316) );
  NOR2_X1 U7199 ( .A1(n6316), .A2(n6321), .ZN(n6050) );
  NAND2_X1 U7200 ( .A1(n6049), .A2(SI_18_), .ZN(n6303) );
  AND2_X1 U7201 ( .A1(n6050), .A2(n6303), .ZN(n6051) );
  INV_X1 U7202 ( .A(n6336), .ZN(n6056) );
  MUX2_X1 U7203 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7532), .Z(n6057) );
  XNOR2_X1 U7204 ( .A(n6057), .B(n6055), .ZN(n6335) );
  NAND2_X1 U7205 ( .A1(n6056), .A2(n6335), .ZN(n6059) );
  NAND2_X1 U7206 ( .A1(n6057), .A2(SI_21_), .ZN(n6058) );
  MUX2_X1 U7207 ( .A(n8383), .B(n8379), .S(n7532), .Z(n6060) );
  NAND2_X1 U7208 ( .A1(n6060), .A2(n8711), .ZN(n6063) );
  INV_X1 U7209 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7210 ( .A1(n6061), .A2(SI_22_), .ZN(n6062) );
  NAND2_X1 U7211 ( .A1(n6063), .A2(n6062), .ZN(n6080) );
  MUX2_X1 U7212 ( .A(n8824), .B(n8505), .S(n7530), .Z(n6064) );
  INV_X1 U7213 ( .A(SI_23_), .ZN(n8710) );
  NAND2_X1 U7214 ( .A1(n6064), .A2(n8710), .ZN(n6348) );
  INV_X1 U7215 ( .A(n6064), .ZN(n6065) );
  NAND2_X1 U7216 ( .A1(n6065), .A2(SI_23_), .ZN(n6066) );
  NAND2_X1 U7217 ( .A1(n6348), .A2(n6066), .ZN(n6067) );
  NAND2_X1 U7218 ( .A1(n5224), .A2(n6067), .ZN(n6069) );
  INV_X1 U7219 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7220 ( .A1(n6069), .A2(n6349), .ZN(n8506) );
  INV_X2 U7221 ( .A(n6137), .ZN(n6172) );
  NAND2_X1 U7222 ( .A1(n8506), .A2(n6172), .ZN(n6071) );
  OR2_X1 U7223 ( .A1(n6104), .A2(n8505), .ZN(n6070) );
  NAND2_X1 U7224 ( .A1(n6342), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7225 ( .A1(n6073), .A2(n6072), .ZN(n9958) );
  NAND2_X1 U7226 ( .A1(n9958), .A2(n5130), .ZN(n6079) );
  INV_X1 U7227 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7228 ( .A1(n8257), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7229 ( .A1(n8250), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7230 ( .C1(n6076), .C2(n8260), .A(n6075), .B(n6074), .ZN(n6077)
         );
  INV_X1 U7231 ( .A(n6077), .ZN(n6078) );
  XNOR2_X1 U7232 ( .A(n6081), .B(n6080), .ZN(n8378) );
  NAND2_X1 U7233 ( .A1(n8378), .A2(n6172), .ZN(n6083) );
  OR2_X1 U7234 ( .A1(n6104), .A2(n8379), .ZN(n6082) );
  NAND2_X1 U7235 ( .A1(n6111), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7236 ( .A1(n5130), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7237 ( .A1(n7532), .A2(SI_0_), .ZN(n6088) );
  INV_X1 U7238 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7239 ( .A1(n6088), .A2(n6087), .ZN(n6090) );
  NAND2_X1 U7240 ( .A1(n6090), .A2(n6089), .ZN(n10177) );
  MUX2_X1 U7241 ( .A(n6091), .B(n10177), .S(n9661), .Z(n8034) );
  INV_X1 U7242 ( .A(n8034), .ZN(n7719) );
  NAND2_X1 U7243 ( .A1(n8390), .A2(n7719), .ZN(n8389) );
  NAND2_X1 U7244 ( .A1(n6111), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7245 ( .A1(n6119), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7246 ( .A1(n6092), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7247 ( .A(n6096), .B(n6097), .ZN(n6618) );
  OR2_X1 U7248 ( .A1(n6137), .A2(n6618), .ZN(n6099) );
  OR2_X1 U7249 ( .A1(n6104), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6098) );
  INV_X1 U7250 ( .A(n8396), .ZN(n6101) );
  NAND2_X1 U7251 ( .A1(n6102), .A2(n6101), .ZN(n6441) );
  NAND2_X1 U7252 ( .A1(n6103), .A2(n8396), .ZN(n9435) );
  AND2_X1 U7253 ( .A1(n6441), .A2(n9435), .ZN(n8392) );
  NAND2_X1 U7254 ( .A1(n8389), .A2(n9589), .ZN(n8388) );
  INV_X1 U7255 ( .A(n8396), .ZN(n10978) );
  NAND2_X1 U7256 ( .A1(n8388), .A2(n10995), .ZN(n6117) );
  INV_X1 U7257 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7565) );
  OR2_X1 U7258 ( .A1(n6104), .A2(n7565), .ZN(n6110) );
  XNOR2_X1 U7259 ( .A(n6106), .B(n6105), .ZN(n7564) );
  OR2_X1 U7260 ( .A1(n6137), .A2(n7564), .ZN(n6109) );
  NAND2_X1 U7261 ( .A1(n6307), .A2(n6107), .ZN(n6108) );
  NAND2_X1 U7262 ( .A1(n5130), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7263 ( .A1(n6111), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7264 ( .A1(n6092), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7265 ( .A1(n5160), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7266 ( .A1(n6116), .A2(n5131), .ZN(n9439) );
  NAND2_X1 U7267 ( .A1(n5131), .A2(n11008), .ZN(n6118) );
  NAND2_X1 U7268 ( .A1(n5130), .A2(n8763), .ZN(n6123) );
  NAND2_X1 U7269 ( .A1(n6111), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7270 ( .A1(n5160), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7271 ( .A1(n6092), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6120) );
  INV_X1 U7272 ( .A(n9806), .ZN(n11002) );
  XNOR2_X1 U7273 ( .A(n6125), .B(n6124), .ZN(n7533) );
  OR2_X1 U7274 ( .A1(n6137), .A2(n7533), .ZN(n6129) );
  INV_X1 U7275 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7531) );
  OR2_X1 U7276 ( .A1(n6104), .A2(n7531), .ZN(n6128) );
  NAND2_X1 U7277 ( .A1(n6307), .A2(n6126), .ZN(n6127) );
  NAND2_X1 U7278 ( .A1(n6111), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7279 ( .A1(n5160), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7280 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6130) );
  NAND2_X1 U7281 ( .A1(n6145), .A2(n6130), .ZN(n8246) );
  NAND2_X1 U7282 ( .A1(n5130), .A2(n8246), .ZN(n6132) );
  NAND2_X1 U7283 ( .A1(n8257), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6131) );
  INV_X1 U7284 ( .A(n9805), .ZN(n9280) );
  XNOR2_X1 U7285 ( .A(n6135), .B(n6136), .ZN(n7558) );
  OR2_X1 U7286 ( .A1(n6137), .A2(n7558), .ZN(n6140) );
  INV_X1 U7287 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7557) );
  OR2_X1 U7288 ( .A1(n6104), .A2(n7557), .ZN(n6139) );
  NAND2_X1 U7289 ( .A1(n6307), .A2(n7969), .ZN(n6138) );
  INV_X1 U7290 ( .A(n11035), .ZN(n8247) );
  NAND2_X1 U7291 ( .A1(n6141), .A2(n8247), .ZN(n6144) );
  NAND2_X1 U7292 ( .A1(n6142), .A2(n9805), .ZN(n6143) );
  NAND2_X1 U7293 ( .A1(n8250), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7294 ( .A1(n5160), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7295 ( .A1(n6145), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7296 ( .A1(n6156), .A2(n6146), .ZN(n9282) );
  NAND2_X1 U7297 ( .A1(n5130), .A2(n9282), .ZN(n6148) );
  NAND2_X1 U7298 ( .A1(n8257), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6147) );
  NAND4_X1 U7299 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n9804)
         );
  AOI22_X1 U7300 ( .A1(n6306), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6307), .B2(
        n6151), .ZN(n6154) );
  NAND2_X1 U7301 ( .A1(n7547), .A2(n6172), .ZN(n6153) );
  INV_X1 U7302 ( .A(n11048), .ZN(n9286) );
  INV_X1 U7303 ( .A(n9804), .ZN(n8025) );
  NAND2_X1 U7304 ( .A1(n8025), .A2(n11048), .ZN(n6155) );
  NAND2_X1 U7305 ( .A1(n8257), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7306 ( .A1(n8250), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7307 ( .A1(n6156), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7308 ( .A1(n6175), .A2(n6157), .ZN(n8208) );
  NAND2_X1 U7309 ( .A1(n5130), .A2(n8208), .ZN(n6159) );
  NAND2_X1 U7310 ( .A1(n5160), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6158) );
  NAND4_X1 U7311 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n9803)
         );
  INV_X1 U7312 ( .A(n9803), .ZN(n9281) );
  NAND2_X1 U7313 ( .A1(n7555), .A2(n6172), .ZN(n6165) );
  AOI22_X1 U7314 ( .A1(n6306), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6307), .B2(
        n6163), .ZN(n6164) );
  AND2_X1 U7315 ( .A1(n9281), .A2(n11063), .ZN(n6166) );
  NAND2_X1 U7316 ( .A1(n7553), .A2(n6172), .ZN(n6174) );
  AOI22_X1 U7317 ( .A1(n6306), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6307), .B2(
        n7807), .ZN(n6173) );
  NAND2_X1 U7318 ( .A1(n8257), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7319 ( .A1(n8250), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7320 ( .A1(n6175), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7321 ( .A1(n6186), .A2(n6176), .ZN(n8219) );
  NAND2_X1 U7322 ( .A1(n5130), .A2(n8219), .ZN(n6178) );
  NAND2_X1 U7323 ( .A1(n5160), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7324 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n9802)
         );
  OR2_X1 U7325 ( .A1(n9472), .A2(n9802), .ZN(n8226) );
  NAND2_X1 U7326 ( .A1(n9472), .A2(n9802), .ZN(n6181) );
  XNOR2_X1 U7327 ( .A(n6183), .B(n6182), .ZN(n7569) );
  NAND2_X1 U7328 ( .A1(n7569), .A2(n6172), .ZN(n6185) );
  AOI22_X1 U7329 ( .A1(n6306), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6307), .B2(
        n7872), .ZN(n6184) );
  NAND2_X1 U7330 ( .A1(n8250), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7331 ( .A1(n8257), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7332 ( .A1(n6186), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7333 ( .A1(n6195), .A2(n6187), .ZN(n8274) );
  NAND2_X1 U7334 ( .A1(n5130), .A2(n8274), .ZN(n6189) );
  NAND2_X1 U7335 ( .A1(n5160), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6188) );
  NAND4_X1 U7336 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n9801)
         );
  INV_X1 U7337 ( .A(n11104), .ZN(n8230) );
  NAND2_X1 U7338 ( .A1(n8230), .A2(n8304), .ZN(n9474) );
  INV_X1 U7339 ( .A(n9597), .ZN(n6192) );
  NAND2_X1 U7340 ( .A1(n11104), .A2(n8304), .ZN(n8195) );
  NAND2_X1 U7341 ( .A1(n8194), .A2(n8195), .ZN(n6202) );
  XNOR2_X1 U7342 ( .A(n6193), .B(n5742), .ZN(n7588) );
  AOI22_X1 U7343 ( .A1(n6306), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6307), .B2(
        n8153), .ZN(n6194) );
  NAND2_X1 U7344 ( .A1(n8250), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7345 ( .A1(n8257), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7346 ( .A1(n6195), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7347 ( .A1(n6208), .A2(n6196), .ZN(n8309) );
  NAND2_X1 U7348 ( .A1(n5130), .A2(n8309), .ZN(n6198) );
  NAND2_X1 U7349 ( .A1(n5160), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7350 ( .A1(n11123), .A2(n8425), .ZN(n9475) );
  INV_X1 U7351 ( .A(n9598), .ZN(n6201) );
  NAND2_X1 U7352 ( .A1(n6202), .A2(n6201), .ZN(n8197) );
  OR2_X1 U7353 ( .A1(n11123), .A2(n9800), .ZN(n6203) );
  XNOR2_X1 U7354 ( .A(n6205), .B(n6204), .ZN(n7591) );
  NAND2_X1 U7355 ( .A1(n7591), .A2(n6172), .ZN(n6207) );
  AOI22_X1 U7356 ( .A1(n6306), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6307), .B2(
        n8375), .ZN(n6206) );
  NAND2_X1 U7357 ( .A1(n6207), .A2(n6206), .ZN(n11139) );
  NAND2_X1 U7358 ( .A1(n8250), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7359 ( .A1(n8257), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7360 ( .A1(n6208), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7361 ( .A1(n6218), .A2(n6209), .ZN(n8998) );
  NAND2_X1 U7362 ( .A1(n5130), .A2(n8998), .ZN(n6211) );
  NAND2_X1 U7363 ( .A1(n5160), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7364 ( .A1(n11139), .A2(n9799), .ZN(n8421) );
  OR2_X1 U7365 ( .A1(n11139), .A2(n9799), .ZN(n8422) );
  XNOR2_X1 U7366 ( .A(n6215), .B(n6214), .ZN(n7596) );
  NAND2_X1 U7367 ( .A1(n7596), .A2(n6172), .ZN(n6217) );
  AOI22_X1 U7368 ( .A1(n6306), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6307), .B2(
        n8450), .ZN(n6216) );
  NAND2_X1 U7369 ( .A1(n6217), .A2(n6216), .ZN(n11143) );
  NAND2_X1 U7370 ( .A1(n8257), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7371 ( .A1(n8250), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7372 ( .A1(n6218), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7373 ( .A1(n6228), .A2(n6219), .ZN(n9035) );
  NAND2_X1 U7374 ( .A1(n5130), .A2(n9035), .ZN(n6221) );
  NAND2_X1 U7375 ( .A1(n5160), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6220) );
  INV_X1 U7376 ( .A(n9070), .ZN(n9798) );
  XNOR2_X1 U7377 ( .A(n6225), .B(n6224), .ZN(n7683) );
  NAND2_X1 U7378 ( .A1(n7683), .A2(n6172), .ZN(n6227) );
  AOI22_X1 U7379 ( .A1(n6306), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6307), .B2(
        n9020), .ZN(n6226) );
  NAND2_X1 U7380 ( .A1(n6227), .A2(n6226), .ZN(n11157) );
  NAND2_X1 U7381 ( .A1(n8257), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7382 ( .A1(n8250), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7383 ( .A1(n6228), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7384 ( .A1(n6240), .A2(n6229), .ZN(n9080) );
  NAND2_X1 U7385 ( .A1(n5130), .A2(n9080), .ZN(n6231) );
  NAND2_X1 U7386 ( .A1(n5160), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6230) );
  NAND4_X1 U7387 ( .A1(n6233), .A2(n6232), .A3(n6231), .A4(n6230), .ZN(n9797)
         );
  XNOR2_X1 U7388 ( .A(n11157), .B(n9797), .ZN(n8404) );
  INV_X1 U7389 ( .A(n8404), .ZN(n9603) );
  NAND2_X1 U7390 ( .A1(n8400), .A2(n9603), .ZN(n6235) );
  NAND2_X1 U7391 ( .A1(n11157), .A2(n9797), .ZN(n6234) );
  XNOR2_X1 U7392 ( .A(n6237), .B(n6236), .ZN(n7697) );
  NAND2_X1 U7393 ( .A1(n7697), .A2(n6172), .ZN(n6239) );
  AOI22_X1 U7394 ( .A1(n6306), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6307), .B2(
        n9130), .ZN(n6238) );
  NAND2_X1 U7395 ( .A1(n6239), .A2(n6238), .ZN(n9152) );
  NAND2_X1 U7396 ( .A1(n8250), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7397 ( .A1(n8257), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7398 ( .A1(n6240), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7399 ( .A1(n6251), .A2(n6241), .ZN(n9169) );
  NAND2_X1 U7400 ( .A1(n5130), .A2(n9169), .ZN(n6243) );
  NAND2_X1 U7401 ( .A1(n5160), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6242) );
  INV_X1 U7402 ( .A(n9153), .ZN(n9796) );
  AND2_X1 U7403 ( .A1(n9152), .A2(n9796), .ZN(n6246) );
  XNOR2_X1 U7404 ( .A(n6248), .B(n6247), .ZN(n7722) );
  NAND2_X1 U7405 ( .A1(n7722), .A2(n6172), .ZN(n6250) );
  AOI22_X1 U7406 ( .A1(n6306), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6307), .B2(
        n9822), .ZN(n6249) );
  NAND2_X1 U7407 ( .A1(n6250), .A2(n6249), .ZN(n10164) );
  NAND2_X1 U7408 ( .A1(n8250), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7409 ( .A1(n8257), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7410 ( .A1(n6251), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7411 ( .A1(n6264), .A2(n6252), .ZN(n9197) );
  NAND2_X1 U7412 ( .A1(n5130), .A2(n9197), .ZN(n6254) );
  NAND2_X1 U7413 ( .A1(n5160), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6253) );
  NAND4_X1 U7414 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n9795)
         );
  NAND2_X1 U7415 ( .A1(n10164), .A2(n9795), .ZN(n9514) );
  OR2_X1 U7416 ( .A1(n10164), .A2(n9795), .ZN(n6257) );
  INV_X1 U7417 ( .A(n8973), .ZN(n9605) );
  NAND2_X1 U7418 ( .A1(n6259), .A2(n6258), .ZN(n6261) );
  XNOR2_X1 U7419 ( .A(n6261), .B(n6260), .ZN(n6585) );
  NAND2_X1 U7420 ( .A1(n6585), .A2(n6172), .ZN(n6263) );
  AOI22_X1 U7421 ( .A1(n6306), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6307), .B2(
        n9839), .ZN(n6262) );
  NAND2_X1 U7422 ( .A1(n6263), .A2(n6262), .ZN(n9201) );
  NAND2_X1 U7423 ( .A1(n8250), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7424 ( .A1(n5160), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7425 ( .A1(n6264), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7426 ( .A1(n6274), .A2(n6265), .ZN(n9211) );
  NAND2_X1 U7427 ( .A1(n5130), .A2(n9211), .ZN(n6267) );
  NAND2_X1 U7428 ( .A1(n8257), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7429 ( .A1(n9201), .A2(n9244), .ZN(n9509) );
  NAND2_X1 U7430 ( .A1(n9201), .A2(n9244), .ZN(n9507) );
  INV_X1 U7431 ( .A(n9607), .ZN(n9515) );
  NAND2_X1 U7432 ( .A1(n9201), .A2(n9794), .ZN(n9084) );
  NAND2_X1 U7433 ( .A1(n9061), .A2(n9084), .ZN(n6280) );
  NAND2_X1 U7434 ( .A1(n7971), .A2(n6172), .ZN(n6273) );
  AOI22_X1 U7435 ( .A1(n6306), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9857), .B2(
        n6307), .ZN(n6272) );
  NAND2_X1 U7436 ( .A1(n6273), .A2(n6272), .ZN(n9246) );
  NAND2_X1 U7437 ( .A1(n8257), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7438 ( .A1(n8250), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7439 ( .A1(n6274), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7440 ( .A1(n6286), .A2(n6275), .ZN(n9240) );
  NAND2_X1 U7441 ( .A1(n5130), .A2(n9240), .ZN(n6277) );
  NAND2_X1 U7442 ( .A1(n5160), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6276) );
  OR2_X1 U7443 ( .A1(n9246), .A2(n10019), .ZN(n9519) );
  NAND2_X1 U7444 ( .A1(n9246), .A2(n10019), .ZN(n9520) );
  NAND2_X1 U7445 ( .A1(n9519), .A2(n9520), .ZN(n9516) );
  NAND2_X1 U7446 ( .A1(n6280), .A2(n9516), .ZN(n9086) );
  NAND2_X1 U7447 ( .A1(n9246), .A2(n9793), .ZN(n6281) );
  NAND2_X1 U7448 ( .A1(n9086), .A2(n6281), .ZN(n10018) );
  XNOR2_X1 U7449 ( .A(n6283), .B(n6282), .ZN(n8030) );
  NAND2_X1 U7450 ( .A1(n8030), .A2(n6172), .ZN(n6285) );
  AOI22_X1 U7451 ( .A1(n9882), .A2(n6307), .B1(n6306), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7452 ( .A1(n8257), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7453 ( .A1(n8250), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7454 ( .A1(n6286), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7455 ( .A1(n6296), .A2(n6287), .ZN(n10027) );
  NAND2_X1 U7456 ( .A1(n5130), .A2(n10027), .ZN(n6289) );
  NAND2_X1 U7457 ( .A1(n5160), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6288) );
  XNOR2_X1 U7458 ( .A(n10151), .B(n9764), .ZN(n10024) );
  NAND2_X1 U7459 ( .A1(n10151), .A2(n10002), .ZN(n6292) );
  NAND2_X1 U7460 ( .A1(n8065), .A2(n6172), .ZN(n6295) );
  AOI22_X1 U7461 ( .A1(n6306), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6307), .B2(
        n10962), .ZN(n6294) );
  NAND2_X1 U7462 ( .A1(n6296), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7463 ( .A1(n6310), .A2(n6297), .ZN(n10006) );
  NAND2_X1 U7464 ( .A1(n10006), .A2(n5130), .ZN(n6301) );
  NAND2_X1 U7465 ( .A1(n8257), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7466 ( .A1(n8250), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7467 ( .A1(n5160), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6298) );
  OR2_X1 U7468 ( .A1(n10086), .A2(n9791), .ZN(n6302) );
  NAND2_X1 U7469 ( .A1(n8278), .A2(n6172), .ZN(n6309) );
  AOI22_X1 U7470 ( .A1(n5136), .A2(n6307), .B1(n6306), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7471 ( .A1(n6309), .A2(n6308), .ZN(n10146) );
  NAND2_X1 U7472 ( .A1(n6310), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7473 ( .A1(n6326), .A2(n6311), .ZN(n9992) );
  NAND2_X1 U7474 ( .A1(n9992), .A2(n5130), .ZN(n6314) );
  AOI22_X1 U7475 ( .A1(n8250), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8257), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7476 ( .A1(n5160), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6312) );
  OR2_X1 U7477 ( .A1(n10146), .A2(n9744), .ZN(n9534) );
  NAND2_X1 U7478 ( .A1(n10146), .A2(n9744), .ZN(n9535) );
  INV_X1 U7479 ( .A(n9995), .ZN(n9610) );
  INV_X1 U7480 ( .A(n6315), .ZN(n6318) );
  INV_X1 U7481 ( .A(n6316), .ZN(n6317) );
  NAND2_X1 U7482 ( .A1(n6320), .A2(n6319), .ZN(n6323) );
  INV_X1 U7483 ( .A(n6321), .ZN(n6322) );
  NAND2_X1 U7484 ( .A1(n8384), .A2(n6172), .ZN(n6325) );
  OR2_X1 U7485 ( .A1(n6104), .A2(n8385), .ZN(n6324) );
  XNOR2_X1 U7486 ( .A(n6326), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U7487 ( .A1(n9983), .A2(n5130), .ZN(n6332) );
  INV_X1 U7488 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7489 ( .A1(n8257), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7490 ( .A1(n8250), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6327) );
  OAI211_X1 U7491 ( .C1(n6329), .C2(n8260), .A(n6328), .B(n6327), .ZN(n6330)
         );
  INV_X1 U7492 ( .A(n6330), .ZN(n6331) );
  NAND2_X1 U7493 ( .A1(n9539), .A2(n9988), .ZN(n6333) );
  XNOR2_X1 U7494 ( .A(n6336), .B(n6335), .ZN(n8300) );
  NAND2_X1 U7495 ( .A1(n8300), .A2(n6172), .ZN(n6338) );
  INV_X1 U7496 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8325) );
  OR2_X1 U7497 ( .A1(n6104), .A2(n8325), .ZN(n6337) );
  INV_X1 U7498 ( .A(n6339), .ZN(n6340) );
  NAND2_X1 U7499 ( .A1(n6340), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7500 ( .A1(n6342), .A2(n6341), .ZN(n9967) );
  NAND2_X1 U7501 ( .A1(n9967), .A2(n5130), .ZN(n6347) );
  INV_X1 U7502 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U7503 ( .A1(n8257), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7504 ( .A1(n8250), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6343) );
  OAI211_X1 U7505 ( .C1(n9969), .C2(n8260), .A(n6344), .B(n6343), .ZN(n6345)
         );
  INV_X1 U7506 ( .A(n6345), .ZN(n6346) );
  NAND2_X1 U7507 ( .A1(n10072), .A2(n9978), .ZN(n9547) );
  NAND2_X1 U7508 ( .A1(n9542), .A2(n9547), .ZN(n9971) );
  INV_X1 U7509 ( .A(n9971), .ZN(n9965) );
  NAND2_X1 U7510 ( .A1(n9964), .A2(n9965), .ZN(n9963) );
  INV_X1 U7511 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9024) );
  MUX2_X1 U7512 ( .A(n9024), .B(n9040), .S(n7530), .Z(n6350) );
  INV_X1 U7513 ( .A(SI_24_), .ZN(n8517) );
  NAND2_X1 U7514 ( .A1(n6350), .A2(n8517), .ZN(n6370) );
  INV_X1 U7515 ( .A(n6350), .ZN(n6351) );
  NAND2_X1 U7516 ( .A1(n6351), .A2(SI_24_), .ZN(n6352) );
  XNOR2_X1 U7517 ( .A(n6369), .B(n6368), .ZN(n9023) );
  NAND2_X1 U7518 ( .A1(n9023), .A2(n6172), .ZN(n6354) );
  OR2_X1 U7519 ( .A1(n6104), .A2(n9040), .ZN(n6353) );
  INV_X1 U7520 ( .A(n6357), .ZN(n6356) );
  INV_X1 U7521 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U7522 ( .A1(n6357), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7523 ( .A1(n6373), .A2(n6358), .ZN(n9935) );
  NAND2_X1 U7524 ( .A1(n9935), .A2(n5130), .ZN(n6364) );
  INV_X1 U7525 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7526 ( .A1(n8257), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7527 ( .A1(n8250), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6359) );
  OAI211_X1 U7528 ( .C1(n6361), .C2(n8260), .A(n6360), .B(n6359), .ZN(n6362)
         );
  INV_X1 U7529 ( .A(n6362), .ZN(n6363) );
  OAI21_X1 U7530 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n9918) );
  MUX2_X1 U7531 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n7532), .Z(n6381) );
  XNOR2_X1 U7532 ( .A(n6381), .B(n8518), .ZN(n6380) );
  XNOR2_X1 U7533 ( .A(n6383), .B(n6380), .ZN(n9054) );
  INV_X1 U7534 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9057) );
  NOR2_X1 U7535 ( .A1(n6104), .A2(n9057), .ZN(n6371) );
  INV_X1 U7536 ( .A(n6373), .ZN(n6372) );
  INV_X1 U7537 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U7538 ( .A1(n6373), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7539 ( .A1(n6406), .A2(n6374), .ZN(n9719) );
  NAND2_X1 U7540 ( .A1(n9719), .A2(n5130), .ZN(n6379) );
  INV_X1 U7541 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U7542 ( .A1(n8257), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7543 ( .A1(n8250), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U7544 ( .C1(n9922), .C2(n8260), .A(n6376), .B(n6375), .ZN(n6377)
         );
  INV_X1 U7545 ( .A(n6377), .ZN(n6378) );
  NAND2_X1 U7546 ( .A1(n6379), .A2(n6378), .ZN(n9788) );
  AND2_X1 U7547 ( .A1(n10126), .A2(n9788), .ZN(n6460) );
  INV_X1 U7548 ( .A(n6460), .ZN(n9563) );
  INV_X1 U7549 ( .A(n10126), .ZN(n9925) );
  NAND2_X1 U7550 ( .A1(n9925), .A2(n9932), .ZN(n9562) );
  INV_X1 U7551 ( .A(n6380), .ZN(n6382) );
  INV_X1 U7552 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9113) );
  MUX2_X1 U7553 ( .A(n9111), .B(n9113), .S(n7532), .Z(n6385) );
  INV_X1 U7554 ( .A(SI_26_), .ZN(n6384) );
  NAND2_X1 U7555 ( .A1(n6385), .A2(n6384), .ZN(n6397) );
  INV_X1 U7556 ( .A(n6385), .ZN(n6386) );
  NAND2_X1 U7557 ( .A1(n6386), .A2(SI_26_), .ZN(n6387) );
  NAND2_X1 U7558 ( .A1(n6397), .A2(n6387), .ZN(n6398) );
  NAND2_X1 U7559 ( .A1(n9109), .A2(n6172), .ZN(n6389) );
  OR2_X1 U7560 ( .A1(n6104), .A2(n9113), .ZN(n6388) );
  XNOR2_X1 U7561 ( .A(n6406), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U7562 ( .A1(n9911), .A2(n5130), .ZN(n6395) );
  INV_X1 U7563 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7564 ( .A1(n8257), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7565 ( .A1(n8250), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6390) );
  OAI211_X1 U7566 ( .C1(n6392), .C2(n8260), .A(n6391), .B(n6390), .ZN(n6393)
         );
  INV_X1 U7567 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U7568 ( .A1(n6395), .A2(n6394), .ZN(n9787) );
  NAND2_X1 U7569 ( .A1(n6461), .A2(n9787), .ZN(n9370) );
  INV_X1 U7570 ( .A(n9370), .ZN(n6396) );
  INV_X1 U7571 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9176) );
  INV_X1 U7572 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9174) );
  MUX2_X1 U7573 ( .A(n9176), .B(n9174), .S(n7532), .Z(n6401) );
  INV_X1 U7574 ( .A(SI_27_), .ZN(n6400) );
  NAND2_X1 U7575 ( .A1(n6401), .A2(n6400), .ZN(n6421) );
  INV_X1 U7576 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U7577 ( .A1(n6402), .A2(SI_27_), .ZN(n6403) );
  XNOR2_X1 U7578 ( .A(n6420), .B(n6419), .ZN(n9175) );
  NAND2_X1 U7579 ( .A1(n9175), .A2(n6172), .ZN(n6405) );
  OR2_X1 U7580 ( .A1(n6104), .A2(n9174), .ZN(n6404) );
  INV_X1 U7581 ( .A(n10118), .ZN(n9677) );
  INV_X1 U7582 ( .A(n6406), .ZN(n6408) );
  INV_X1 U7583 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6407) );
  INV_X1 U7584 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8764) );
  INV_X1 U7585 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U7586 ( .A1(n6410), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U7587 ( .A1(n6425), .A2(n6411), .ZN(n9902) );
  NAND2_X1 U7588 ( .A1(n9902), .A2(n5130), .ZN(n6417) );
  INV_X1 U7589 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7590 ( .A1(n8257), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7591 ( .A1(n8250), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6412) );
  OAI211_X1 U7592 ( .C1(n6414), .C2(n8260), .A(n6413), .B(n6412), .ZN(n6415)
         );
  INV_X1 U7593 ( .A(n6415), .ZN(n6416) );
  NOR2_X1 U7594 ( .A1(n9677), .A2(n9786), .ZN(n6418) );
  NAND2_X1 U7595 ( .A1(n6420), .A2(n6419), .ZN(n6422) );
  MUX2_X1 U7596 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n7530), .Z(n6497) );
  INV_X1 U7597 ( .A(SI_28_), .ZN(n6498) );
  XNOR2_X1 U7598 ( .A(n6497), .B(n6498), .ZN(n6495) );
  XNOR2_X1 U7599 ( .A(n6496), .B(n6495), .ZN(n9218) );
  NAND2_X1 U7600 ( .A1(n9218), .A2(n6172), .ZN(n6424) );
  INV_X1 U7601 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9217) );
  OR2_X1 U7602 ( .A1(n6104), .A2(n9217), .ZN(n6423) );
  NAND2_X1 U7603 ( .A1(n6425), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7604 ( .A1(n9665), .A2(n6426), .ZN(n9374) );
  NAND2_X1 U7605 ( .A1(n9374), .A2(n5130), .ZN(n6431) );
  INV_X1 U7606 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U7607 ( .A1(n8257), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U7608 ( .A1(n8250), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6427) );
  OAI211_X1 U7609 ( .C1(n9394), .C2(n8260), .A(n6428), .B(n6427), .ZN(n6429)
         );
  INV_X1 U7610 ( .A(n6429), .ZN(n6430) );
  XNOR2_X1 U7611 ( .A(n9657), .B(n9785), .ZN(n9655) );
  XNOR2_X1 U7612 ( .A(n9653), .B(n9655), .ZN(n6440) );
  AND2_X1 U7613 ( .A1(n7485), .A2(n9618), .ZN(n9425) );
  AND2_X1 U7614 ( .A1(n5136), .A2(n9627), .ZN(n6465) );
  INV_X1 U7615 ( .A(n9665), .ZN(n6433) );
  NAND2_X1 U7616 ( .A1(n6433), .A2(n5130), .ZN(n8264) );
  INV_X1 U7617 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U7618 ( .A1(n8257), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7619 ( .A1(n8250), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6434) );
  OAI211_X1 U7620 ( .C1(n9664), .C2(n8260), .A(n6435), .B(n6434), .ZN(n6436)
         );
  INV_X1 U7621 ( .A(n6436), .ZN(n6437) );
  OR2_X1 U7622 ( .A1(n5872), .A2(n9623), .ZN(n6438) );
  NAND2_X1 U7623 ( .A1(n9661), .A2(n6438), .ZN(n7521) );
  INV_X1 U7624 ( .A(n7521), .ZN(n7520) );
  OAI22_X1 U7625 ( .A1(n9419), .A2(n11003), .B1(n9908), .B2(n11001), .ZN(n6439) );
  NAND2_X1 U7626 ( .A1(n8394), .A2(n8392), .ZN(n8393) );
  NAND2_X1 U7627 ( .A1(n8393), .A2(n6441), .ZN(n10994) );
  INV_X1 U7628 ( .A(n6442), .ZN(n9438) );
  NAND2_X1 U7629 ( .A1(n8233), .A2(n9439), .ZN(n6445) );
  NAND2_X1 U7630 ( .A1(n9806), .A2(n11027), .ZN(n9456) );
  INV_X1 U7631 ( .A(n9452), .ZN(n6443) );
  NAND2_X1 U7632 ( .A1(n9805), .A2(n11035), .ZN(n9453) );
  AND2_X1 U7633 ( .A1(n9804), .A2(n11048), .ZN(n9276) );
  OR2_X1 U7634 ( .A1(n9804), .A2(n11048), .ZN(n9457) );
  NAND2_X1 U7635 ( .A1(n11063), .A2(n9803), .ZN(n9464) );
  NAND2_X1 U7636 ( .A1(n8213), .A2(n8217), .ZN(n8212) );
  INV_X1 U7637 ( .A(n9802), .ZN(n9471) );
  OR2_X1 U7638 ( .A1(n9472), .A2(n9471), .ZN(n9483) );
  NAND2_X1 U7639 ( .A1(n8212), .A2(n9483), .ZN(n8225) );
  INV_X1 U7640 ( .A(n8225), .ZN(n6449) );
  AOI21_X2 U7641 ( .B1(n6449), .B2(n5166), .A(n6448), .ZN(n8193) );
  NAND2_X1 U7642 ( .A1(n11139), .A2(n8410), .ZN(n9487) );
  NAND2_X1 U7643 ( .A1(n6450), .A2(n9487), .ZN(n8415) );
  OR2_X1 U7644 ( .A1(n11143), .A2(n9070), .ZN(n9492) );
  NAND2_X1 U7645 ( .A1(n11143), .A2(n9070), .ZN(n9490) );
  NAND2_X1 U7646 ( .A1(n8415), .A2(n8414), .ZN(n8413) );
  NAND2_X1 U7647 ( .A1(n8413), .A2(n9490), .ZN(n8405) );
  NAND2_X1 U7648 ( .A1(n11157), .A2(n9495), .ZN(n9494) );
  AND2_X1 U7649 ( .A1(n9152), .A2(n9153), .ZN(n8956) );
  OR2_X1 U7650 ( .A1(n9152), .A2(n9153), .ZN(n9499) );
  INV_X1 U7651 ( .A(n10164), .ZN(n9502) );
  NAND2_X1 U7652 ( .A1(n9060), .A2(n9607), .ZN(n6451) );
  NAND2_X1 U7653 ( .A1(n6451), .A2(n9507), .ZN(n9089) );
  INV_X1 U7654 ( .A(n9089), .ZN(n6453) );
  INV_X1 U7655 ( .A(n9516), .ZN(n6452) );
  NAND2_X1 U7656 ( .A1(n10151), .A2(n9764), .ZN(n6454) );
  NAND2_X1 U7657 ( .A1(n10086), .A2(n10020), .ZN(n9531) );
  NAND2_X1 U7658 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  NAND2_X1 U7659 ( .A1(n10009), .A2(n9530), .ZN(n9996) );
  NAND2_X1 U7660 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  AND2_X2 U7661 ( .A1(n9994), .A2(n9534), .ZN(n9982) );
  INV_X1 U7662 ( .A(n9988), .ZN(n9709) );
  NAND2_X1 U7663 ( .A1(n9539), .A2(n9709), .ZN(n6456) );
  INV_X1 U7664 ( .A(n9978), .ZN(n9955) );
  NAND2_X1 U7665 ( .A1(n9351), .A2(n9943), .ZN(n9550) );
  NAND2_X1 U7666 ( .A1(n9957), .A2(n9550), .ZN(n6457) );
  OR2_X1 U7667 ( .A1(n9351), .A2(n9943), .ZN(n9551) );
  NAND2_X1 U7668 ( .A1(n6457), .A2(n9551), .ZN(n9945) );
  NAND2_X1 U7669 ( .A1(n9945), .A2(n9940), .ZN(n6458) );
  OR2_X1 U7670 ( .A1(n9553), .A2(n9954), .ZN(n9554) );
  NAND2_X1 U7671 ( .A1(n6458), .A2(n9554), .ZN(n9933) );
  NAND2_X1 U7672 ( .A1(n9432), .A2(n9944), .ZN(n9559) );
  NAND2_X1 U7673 ( .A1(n9933), .A2(n9559), .ZN(n6459) );
  OR2_X1 U7674 ( .A1(n9432), .A2(n9944), .ZN(n9560) );
  AND2_X1 U7675 ( .A1(n10122), .A2(n9787), .ZN(n9403) );
  INV_X1 U7676 ( .A(n9403), .ZN(n9567) );
  NAND2_X1 U7677 ( .A1(n9401), .A2(n9567), .ZN(n9899) );
  INV_X1 U7678 ( .A(n9787), .ZN(n9921) );
  NAND2_X1 U7679 ( .A1(n6461), .A2(n9921), .ZN(n9898) );
  INV_X1 U7680 ( .A(n9898), .ZN(n9366) );
  NOR2_X1 U7681 ( .A1(n9431), .A2(n9366), .ZN(n6462) );
  AND2_X1 U7682 ( .A1(n10118), .A2(n9786), .ZN(n9402) );
  XNOR2_X1 U7683 ( .A(n9656), .B(n9655), .ZN(n9396) );
  NAND2_X1 U7684 ( .A1(n8387), .A2(n5135), .ZN(n7183) );
  NAND2_X1 U7685 ( .A1(n7515), .A2(n11179), .ZN(n7992) );
  INV_X1 U7686 ( .A(n9627), .ZN(n8380) );
  AND2_X1 U7687 ( .A1(n9618), .A2(n8380), .ZN(n6463) );
  OR3_X1 U7688 ( .A1(n7992), .A2(n5136), .A3(n6463), .ZN(n9660) );
  NOR2_X1 U7689 ( .A1(n7484), .A2(n9627), .ZN(n10039) );
  INV_X1 U7690 ( .A(n10039), .ZN(n11135) );
  NAND2_X1 U7691 ( .A1(n9400), .A2(n6464), .ZN(n7190) );
  INV_X1 U7692 ( .A(n6465), .ZN(n6466) );
  NAND3_X1 U7693 ( .A1(n9574), .A2(n11179), .A3(n7494), .ZN(n6467) );
  NAND2_X1 U7694 ( .A1(n6467), .A2(n11007), .ZN(n7506) );
  INV_X1 U7695 ( .A(n6482), .ZN(n9059) );
  INV_X1 U7696 ( .A(P2_B_REG_SCAN_IN), .ZN(n8809) );
  XNOR2_X1 U7697 ( .A(n9039), .B(n8809), .ZN(n6468) );
  NAND2_X1 U7698 ( .A1(n9059), .A2(n6468), .ZN(n6469) );
  OR2_X1 U7699 ( .A1(n7538), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6470) );
  OR2_X1 U7700 ( .A1(n9112), .A2(n9039), .ZN(n7543) );
  NOR2_X1 U7701 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6474) );
  NOR4_X1 U7702 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6473) );
  NOR4_X1 U7703 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6472) );
  NOR4_X1 U7704 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6471) );
  NAND4_X1 U7705 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6480)
         );
  NOR4_X1 U7706 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6478) );
  NOR4_X1 U7707 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6477) );
  NOR4_X1 U7708 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6476) );
  NOR4_X1 U7709 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6475) );
  NAND4_X1 U7710 ( .A1(n6478), .A2(n6477), .A3(n6476), .A4(n6475), .ZN(n6479)
         );
  NOR2_X1 U7711 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  INV_X1 U7712 ( .A(n7185), .ZN(n6486) );
  NOR2_X1 U7713 ( .A1(n7985), .A2(n6486), .ZN(n6484) );
  OR2_X1 U7714 ( .A1(n6482), .A2(n9112), .ZN(n7540) );
  NAND2_X1 U7715 ( .A1(n7506), .A2(n7519), .ZN(n6489) );
  NAND2_X1 U7716 ( .A1(n7515), .A2(n7494), .ZN(n6487) );
  NAND2_X1 U7717 ( .A1(n7985), .A2(n6485), .ZN(n7187) );
  NAND2_X1 U7718 ( .A1(n6487), .A2(n7523), .ZN(n6488) );
  NAND2_X1 U7719 ( .A1(n7190), .A2(n11191), .ZN(n6494) );
  INV_X1 U7720 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U7721 ( .A1(n6496), .A2(n6495), .ZN(n6501) );
  INV_X1 U7722 ( .A(n6497), .ZN(n6499) );
  NAND2_X1 U7723 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  INV_X1 U7724 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10697) );
  INV_X1 U7725 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10174) );
  MUX2_X1 U7726 ( .A(n10697), .B(n10174), .S(n7530), .Z(n6504) );
  INV_X1 U7727 ( .A(SI_29_), .ZN(n6502) );
  INV_X1 U7728 ( .A(n6503), .ZN(n6506) );
  INV_X1 U7729 ( .A(n6504), .ZN(n6505) );
  NAND2_X1 U7730 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  INV_X1 U7731 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9272) );
  INV_X1 U7732 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9413) );
  MUX2_X1 U7733 ( .A(n9272), .B(n9413), .S(n7532), .Z(n6509) );
  INV_X1 U7734 ( .A(SI_30_), .ZN(n8509) );
  NAND2_X1 U7735 ( .A1(n6509), .A2(n8509), .ZN(n6512) );
  INV_X1 U7736 ( .A(n6509), .ZN(n6510) );
  NAND2_X1 U7737 ( .A1(n6510), .A2(SI_30_), .ZN(n6511) );
  NAND2_X1 U7738 ( .A1(n6512), .A2(n6511), .ZN(n6980) );
  MUX2_X1 U7739 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7532), .Z(n6513) );
  INV_X1 U7740 ( .A(SI_31_), .ZN(n8698) );
  XNOR2_X1 U7741 ( .A(n6513), .B(n8698), .ZN(n6514) );
  AND2_X2 U7742 ( .A1(n6631), .A2(n6516), .ZN(n6655) );
  NOR2_X1 U7743 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6520) );
  NOR2_X1 U7744 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6519) );
  NOR2_X1 U7745 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6518) );
  NOR2_X1 U7746 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6517) );
  INV_X1 U7747 ( .A(n6535), .ZN(n6521) );
  NAND2_X1 U7748 ( .A1(n7169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7174) );
  INV_X1 U7749 ( .A(n7174), .ZN(n6522) );
  NAND2_X1 U7750 ( .A1(n7177), .A2(n6527), .ZN(n6524) );
  NAND2_X1 U7751 ( .A1(n6522), .A2(n8904), .ZN(n6523) );
  NAND2_X2 U7752 ( .A1(n6620), .A2(n6525), .ZN(n6657) );
  INV_X2 U7753 ( .A(n6657), .ZN(n6690) );
  INV_X1 U7754 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10689) );
  NOR2_X1 U7755 ( .A1(n6982), .A2(n10689), .ZN(n6526) );
  NAND2_X2 U7756 ( .A1(n9270), .A2(n5624), .ZN(n6924) );
  INV_X1 U7757 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7758 ( .A1(n6954), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6533) );
  INV_X1 U7759 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9326) );
  OR2_X1 U7760 ( .A1(n6958), .A2(n9326), .ZN(n6532) );
  OAI211_X1 U7761 ( .C1(n6969), .C2(n6534), .A(n6533), .B(n6532), .ZN(n10319)
         );
  INV_X1 U7762 ( .A(n10319), .ZN(n6986) );
  NAND3_X1 U7763 ( .A1(n6831), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7764 ( .A1(n6538), .A2(n6544), .ZN(n6542) );
  NAND2_X1 U7765 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n6539) );
  NAND2_X1 U7766 ( .A1(n6539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6540) );
  OAI21_X1 U7767 ( .B1(n8669), .B2(P1_IR_REG_31__SCAN_IN), .A(n6540), .ZN(
        n6541) );
  INV_X1 U7768 ( .A(n6547), .ZN(n6548) );
  NAND2_X1 U7769 ( .A1(n6548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7770 ( .A1(n6987), .A2(n6549), .ZN(n6550) );
  NAND2_X1 U7771 ( .A1(n6550), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U7772 ( .B1(n7153), .B2(n7172), .A(n8381), .ZN(n7090) );
  NAND2_X1 U7773 ( .A1(n6954), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6555) );
  INV_X1 U7774 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6552) );
  OR2_X1 U7775 ( .A1(n6969), .A2(n6552), .ZN(n6554) );
  INV_X1 U7776 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10440) );
  OR2_X1 U7777 ( .A1(n6958), .A2(n10440), .ZN(n6553) );
  AND3_X1 U7778 ( .A1(n6555), .A2(n6554), .A3(n6553), .ZN(n7015) );
  INV_X1 U7779 ( .A(n7015), .ZN(n10320) );
  NAND2_X1 U7780 ( .A1(n10319), .A2(n10320), .ZN(n7080) );
  NAND2_X1 U7781 ( .A1(n9109), .A2(n6690), .ZN(n6557) );
  OR2_X1 U7782 ( .A1(n6982), .A2(n9111), .ZN(n6556) );
  NAND2_X1 U7783 ( .A1(n6954), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6565) );
  INV_X1 U7784 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6558) );
  OR2_X1 U7785 ( .A1(n6969), .A2(n6558), .ZN(n6564) );
  INV_X1 U7786 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6559) );
  OR2_X1 U7787 ( .A1(n6958), .A2(n6559), .ZN(n6563) );
  NAND2_X1 U7788 ( .A1(n6671), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6681) );
  INV_X1 U7789 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6680) );
  NOR2_X1 U7790 ( .A1(n6681), .A2(n6680), .ZN(n6697) );
  NAND2_X1 U7791 ( .A1(n6697), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U7792 ( .A1(n6757), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U7793 ( .A1(n6804), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U7794 ( .A1(n6591), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6817) );
  INV_X1 U7795 ( .A(n6817), .ZN(n6560) );
  NAND2_X1 U7796 ( .A1(n6560), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6818) );
  INV_X1 U7797 ( .A(n6851), .ZN(n6561) );
  NAND2_X1 U7798 ( .A1(n6561), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U7799 ( .A1(n6569), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U7800 ( .B1(n6569), .B2(P1_REG3_REG_26__SCAN_IN), .A(n6938), .ZN(
        n10486) );
  OR2_X1 U7801 ( .A1(n6649), .A2(n10486), .ZN(n6562) );
  NAND4_X1 U7802 ( .A1(n6565), .A2(n6564), .A3(n6563), .A4(n6562), .ZN(n10324)
         );
  NAND2_X1 U7803 ( .A1(n10632), .A2(n10504), .ZN(n9296) );
  NAND2_X1 U7804 ( .A1(n9054), .A2(n6690), .ZN(n6567) );
  INV_X1 U7805 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9055) );
  OR2_X1 U7806 ( .A1(n6982), .A2(n9055), .ZN(n6566) );
  NAND2_X1 U7807 ( .A1(n6954), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6576) );
  INV_X1 U7808 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7809 ( .A1(n6969), .A2(n6568), .ZN(n6575) );
  INV_X1 U7810 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10497) );
  OR2_X1 U7811 ( .A1(n6958), .A2(n10497), .ZN(n6574) );
  INV_X1 U7812 ( .A(n6569), .ZN(n6572) );
  INV_X1 U7813 ( .A(n6570), .ZN(n6928) );
  INV_X1 U7814 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U7815 ( .A1(n6928), .A2(n10207), .ZN(n6571) );
  NAND2_X1 U7816 ( .A1(n6572), .A2(n6571), .ZN(n10496) );
  OR2_X1 U7817 ( .A1(n6971), .A2(n10496), .ZN(n6573) );
  NAND4_X1 U7818 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .ZN(n10513)
         );
  NAND2_X1 U7819 ( .A1(n10637), .A2(n10483), .ZN(n9295) );
  NAND2_X1 U7820 ( .A1(n9296), .A2(n9295), .ZN(n7138) );
  NOR2_X1 U7821 ( .A1(n10632), .A2(n10504), .ZN(n7070) );
  INV_X2 U7822 ( .A(n6982), .ZN(n6846) );
  OR2_X1 U7823 ( .A1(n6535), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U7824 ( .A1(n6587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6577) );
  XNOR2_X1 U7825 ( .A(n6577), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U7826 ( .A1(n6846), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6845), .B2(
        n10407), .ZN(n6578) );
  OAI21_X1 U7827 ( .B1(n6591), .B2(P1_REG3_REG_16__SCAN_IN), .A(n6817), .ZN(
        n10589) );
  INV_X1 U7828 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7829 ( .A1(n6954), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6581) );
  INV_X1 U7830 ( .A(n6958), .ZN(n6622) );
  NAND2_X1 U7831 ( .A1(n6622), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U7832 ( .C1(n6969), .C2(n6582), .A(n6581), .B(n6580), .ZN(n6583)
         );
  INV_X1 U7833 ( .A(n6583), .ZN(n6584) );
  INV_X1 U7834 ( .A(n11235), .ZN(n10242) );
  NAND2_X1 U7835 ( .A1(n10602), .A2(n10242), .ZN(n7126) );
  NAND2_X1 U7836 ( .A1(n6585), .A2(n6690), .ZN(n6590) );
  NAND2_X1 U7837 ( .A1(n6535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6586) );
  MUX2_X1 U7838 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6586), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6588) );
  AOI22_X1 U7839 ( .A1(n6846), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6845), .B2(
        n10859), .ZN(n6589) );
  NAND2_X1 U7840 ( .A1(n6590), .A2(n6589), .ZN(n7337) );
  INV_X1 U7841 ( .A(n6649), .ZN(n6852) );
  AOI21_X1 U7842 ( .B1(n6803), .B2(n10310), .A(n6591), .ZN(n11215) );
  NAND2_X1 U7843 ( .A1(n6852), .A2(n11215), .ZN(n6598) );
  INV_X1 U7844 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6592) );
  OR2_X1 U7845 ( .A1(n6924), .A2(n6592), .ZN(n6597) );
  INV_X1 U7846 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6593) );
  OR2_X1 U7847 ( .A1(n5133), .A2(n6593), .ZN(n6596) );
  INV_X1 U7848 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6594) );
  OR2_X1 U7849 ( .A1(n6625), .A2(n6594), .ZN(n6595) );
  NAND4_X1 U7850 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n10594)
         );
  INV_X1 U7851 ( .A(n10594), .ZN(n10215) );
  NAND2_X1 U7852 ( .A1(n7337), .A2(n10215), .ZN(n6995) );
  OAI211_X1 U7853 ( .C1(n11235), .C2(n6995), .A(n11224), .B(n6949), .ZN(n6600)
         );
  NAND3_X1 U7854 ( .A1(n6995), .A2(n11235), .A3(n6949), .ZN(n6599) );
  OAI211_X1 U7855 ( .C1(n6949), .C2(n7126), .A(n6600), .B(n6599), .ZN(n6601)
         );
  INV_X1 U7856 ( .A(n6601), .ZN(n6829) );
  NAND2_X1 U7857 ( .A1(n6954), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6607) );
  INV_X1 U7858 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6602) );
  OR2_X1 U7859 ( .A1(n6924), .A2(n6602), .ZN(n6606) );
  INV_X1 U7860 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7748) );
  OR2_X1 U7861 ( .A1(n6649), .A2(n7748), .ZN(n6605) );
  INV_X1 U7862 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6603) );
  OR2_X1 U7863 ( .A1(n6958), .A2(n6603), .ZN(n6604) );
  NAND4_X2 U7864 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n10338)
         );
  INV_X1 U7865 ( .A(SI_0_), .ZN(n6608) );
  NOR2_X1 U7866 ( .A1(n7532), .A2(n6608), .ZN(n6610) );
  INV_X1 U7867 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6609) );
  XNOR2_X1 U7868 ( .A(n6610), .B(n6609), .ZN(n10700) );
  MUX2_X1 U7869 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10700), .S(n6620), .Z(n9259)
         );
  INV_X1 U7870 ( .A(n9259), .ZN(n7651) );
  INV_X1 U7871 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6611) );
  INV_X1 U7872 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6612) );
  OR2_X1 U7873 ( .A1(n6625), .A2(n6612), .ZN(n6613) );
  NAND2_X1 U7874 ( .A1(n6895), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6616) );
  INV_X1 U7875 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6614) );
  NAND3_X1 U7876 ( .A1(n5171), .A2(n6616), .A3(n6615), .ZN(n7098) );
  INV_X1 U7877 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U7878 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6617) );
  XNOR2_X1 U7879 ( .A(n8851), .B(n6617), .ZN(n7614) );
  INV_X1 U7880 ( .A(n6618), .ZN(n7563) );
  NAND2_X1 U7881 ( .A1(n9254), .A2(n9253), .ZN(n9252) );
  INV_X1 U7882 ( .A(n7098), .ZN(n7903) );
  NAND2_X1 U7883 ( .A1(n7903), .A2(n9260), .ZN(n6621) );
  NAND2_X1 U7884 ( .A1(n9252), .A2(n6621), .ZN(n7921) );
  NAND2_X1 U7885 ( .A1(n6622), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6629) );
  INV_X1 U7886 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6623) );
  OR2_X1 U7887 ( .A1(n6924), .A2(n6623), .ZN(n6628) );
  INV_X1 U7888 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6624) );
  OR2_X1 U7889 ( .A1(n6625), .A2(n6624), .ZN(n6627) );
  INV_X1 U7890 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7658) );
  OR2_X1 U7891 ( .A1(n6649), .A2(n7658), .ZN(n6626) );
  NAND4_X2 U7892 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n10336)
         );
  OR2_X1 U7893 ( .A1(n6631), .A2(n7161), .ZN(n6641) );
  INV_X1 U7894 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8850) );
  XNOR2_X1 U7895 ( .A(n6641), .B(n8850), .ZN(n7613) );
  OR2_X1 U7896 ( .A1(n6657), .A2(n7564), .ZN(n6633) );
  INV_X1 U7897 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7535) );
  OR2_X1 U7898 ( .A1(n6982), .A2(n7535), .ZN(n6632) );
  NAND2_X1 U7899 ( .A1(n7921), .A2(n7922), .ZN(n6634) );
  INV_X1 U7900 ( .A(n8925), .ZN(n7936) );
  NAND2_X1 U7901 ( .A1(n6954), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6640) );
  OR2_X1 U7902 ( .A1(n6649), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6639) );
  INV_X1 U7903 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6635) );
  OR2_X1 U7904 ( .A1(n6958), .A2(n6635), .ZN(n6638) );
  INV_X1 U7905 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6636) );
  OR2_X1 U7906 ( .A1(n6924), .A2(n6636), .ZN(n6637) );
  NAND2_X1 U7907 ( .A1(n6641), .A2(n8850), .ZN(n6642) );
  NAND2_X1 U7908 ( .A1(n6642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6643) );
  INV_X1 U7909 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8856) );
  XNOR2_X1 U7910 ( .A(n6643), .B(n8856), .ZN(n7617) );
  OR2_X1 U7911 ( .A1(n6657), .A2(n7533), .ZN(n6645) );
  INV_X1 U7912 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7534) );
  OR2_X1 U7913 ( .A1(n6982), .A2(n7534), .ZN(n6644) );
  OAI211_X1 U7914 ( .C1(n7581), .C2(n7617), .A(n6645), .B(n6644), .ZN(n7730)
         );
  AND2_X1 U7915 ( .A1(n10335), .A2(n11020), .ZN(n6663) );
  NAND2_X1 U7916 ( .A1(n6954), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6653) );
  INV_X1 U7917 ( .A(n6671), .ZN(n6648) );
  INV_X1 U7918 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6646) );
  INV_X1 U7919 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U7920 ( .A1(n6646), .A2(n7978), .ZN(n6647) );
  NAND2_X1 U7921 ( .A1(n6648), .A2(n6647), .ZN(n8055) );
  OR2_X1 U7922 ( .A1(n6649), .A2(n8055), .ZN(n6652) );
  INV_X1 U7923 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6650) );
  OR2_X1 U7924 ( .A1(n6924), .A2(n6650), .ZN(n6651) );
  INV_X1 U7925 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8056) );
  OR2_X1 U7926 ( .A1(n5133), .A2(n8056), .ZN(n6654) );
  AND2_X2 U7927 ( .A1(n5176), .A2(n6654), .ZN(n10228) );
  OR2_X1 U7928 ( .A1(n6655), .A2(n7161), .ZN(n6656) );
  XNOR2_X1 U7929 ( .A(n6656), .B(n8861), .ZN(n10363) );
  INV_X1 U7930 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7537) );
  OR2_X1 U7931 ( .A1(n6982), .A2(n7537), .ZN(n6658) );
  OAI21_X1 U7932 ( .B1(n6661), .B2(n6663), .A(n6660), .ZN(n6662) );
  INV_X1 U7933 ( .A(n6663), .ZN(n7002) );
  NAND2_X1 U7934 ( .A1(n7029), .A2(n7002), .ZN(n7103) );
  NAND2_X1 U7935 ( .A1(n7547), .A2(n6690), .ZN(n6668) );
  OR2_X1 U7936 ( .A1(n6665), .A2(n7161), .ZN(n6666) );
  XNOR2_X1 U7937 ( .A(n6666), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U7938 ( .A1(n6846), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6845), .B2(
        n10764), .ZN(n6667) );
  NAND2_X1 U7939 ( .A1(n6954), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6675) );
  INV_X1 U7940 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6669) );
  OR2_X1 U7941 ( .A1(n6924), .A2(n6669), .ZN(n6674) );
  INV_X1 U7942 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6670) );
  OR2_X1 U7943 ( .A1(n6973), .A2(n6670), .ZN(n6673) );
  OAI21_X1 U7944 ( .B1(n6671), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6681), .ZN(
        n10227) );
  OR2_X1 U7945 ( .A1(n6649), .A2(n10227), .ZN(n6672) );
  NAND4_X1 U7946 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n10333)
         );
  INV_X1 U7947 ( .A(n10333), .ZN(n8005) );
  INV_X1 U7948 ( .A(n7106), .ZN(n7033) );
  NAND2_X1 U7949 ( .A1(n7555), .A2(n6690), .ZN(n6677) );
  INV_X1 U7950 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7951 ( .A1(n6665), .A2(n8648), .ZN(n6709) );
  NAND2_X1 U7952 ( .A1(n6709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6691) );
  XNOR2_X1 U7953 ( .A(n6691), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U7954 ( .A1(n6846), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6845), .B2(
        n10785), .ZN(n6676) );
  NAND2_X1 U7955 ( .A1(n6677), .A2(n6676), .ZN(n8119) );
  NAND2_X1 U7956 ( .A1(n6954), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6686) );
  INV_X1 U7957 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6678) );
  OR2_X1 U7958 ( .A1(n6969), .A2(n6678), .ZN(n6685) );
  INV_X1 U7959 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6679) );
  OR2_X1 U7960 ( .A1(n5133), .A2(n6679), .ZN(n6684) );
  AND2_X1 U7961 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  OR2_X1 U7962 ( .A1(n6682), .A2(n6697), .ZN(n8082) );
  OR2_X1 U7963 ( .A1(n6649), .A2(n8082), .ZN(n6683) );
  NAND4_X1 U7964 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n10332)
         );
  INV_X1 U7965 ( .A(n10332), .ZN(n8099) );
  NOR2_X1 U7966 ( .A1(n8119), .A2(n8099), .ZN(n7001) );
  AOI21_X1 U7967 ( .B1(n6687), .B2(n7033), .A(n7001), .ZN(n6689) );
  OAI21_X1 U7968 ( .B1(n6687), .B2(n7106), .A(n7108), .ZN(n6688) );
  MUX2_X1 U7969 ( .A(n6689), .B(n6688), .S(n6949), .Z(n6704) );
  NAND2_X1 U7970 ( .A1(n6691), .A2(n8860), .ZN(n6692) );
  NAND2_X1 U7971 ( .A1(n6692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U7972 ( .A(n6693), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U7973 ( .A1(n6846), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6845), .B2(
        n10800), .ZN(n6694) );
  NAND2_X1 U7974 ( .A1(n6954), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6702) );
  INV_X1 U7975 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6695) );
  OR2_X1 U7976 ( .A1(n6969), .A2(n6695), .ZN(n6701) );
  INV_X1 U7977 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6696) );
  OR2_X1 U7978 ( .A1(n5133), .A2(n6696), .ZN(n6700) );
  OR2_X1 U7979 ( .A1(n6697), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U7980 ( .A1(n6717), .A2(n6698), .ZN(n8346) );
  OR2_X1 U7981 ( .A1(n6649), .A2(n8346), .ZN(n6699) );
  NAND4_X1 U7982 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n10331)
         );
  INV_X1 U7983 ( .A(n10331), .ZN(n8318) );
  AND2_X1 U7984 ( .A1(n8119), .A2(n8099), .ZN(n7034) );
  INV_X1 U7985 ( .A(n7003), .ZN(n7105) );
  AOI21_X1 U7986 ( .B1(n7105), .B2(n7108), .A(n7034), .ZN(n6703) );
  AOI21_X1 U7987 ( .B1(n6704), .B2(n6703), .A(n7001), .ZN(n6705) );
  MUX2_X1 U7988 ( .A(n6706), .B(n6705), .S(n6949), .Z(n6724) );
  NOR2_X1 U7989 ( .A1(n8348), .A2(n8318), .ZN(n6707) );
  INV_X1 U7990 ( .A(n6707), .ZN(n7038) );
  MUX2_X1 U7991 ( .A(n6707), .B(n7000), .S(n6949), .Z(n6723) );
  NAND2_X1 U7992 ( .A1(n7569), .A2(n6690), .ZN(n6714) );
  INV_X1 U7993 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U7994 ( .A1(n8860), .A2(n8653), .ZN(n6708) );
  NOR2_X1 U7995 ( .A1(n6709), .A2(n6708), .ZN(n6711) );
  OR2_X1 U7996 ( .A1(n6711), .A2(n7161), .ZN(n6710) );
  MUX2_X1 U7997 ( .A(n6710), .B(P1_IR_REG_31__SCAN_IN), .S(n8867), .Z(n6712)
         );
  NAND2_X1 U7998 ( .A1(n6711), .A2(n8867), .ZN(n6766) );
  AOI22_X1 U7999 ( .A1(n6846), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6845), .B2(
        n10813), .ZN(n6713) );
  NAND2_X1 U8000 ( .A1(n6714), .A2(n6713), .ZN(n8321) );
  NAND2_X1 U8001 ( .A1(n6954), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6722) );
  INV_X1 U8002 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6715) );
  OR2_X1 U8003 ( .A1(n6969), .A2(n6715), .ZN(n6721) );
  NAND2_X1 U8004 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  NAND2_X1 U8005 ( .A1(n6728), .A2(n6718), .ZN(n8317) );
  OR2_X1 U8006 ( .A1(n6971), .A2(n8317), .ZN(n6720) );
  INV_X1 U8007 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8185) );
  OR2_X1 U8008 ( .A1(n5133), .A2(n8185), .ZN(n6719) );
  NAND4_X1 U8009 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n10330)
         );
  INV_X1 U8010 ( .A(n10330), .ZN(n9388) );
  OR2_X1 U8011 ( .A1(n8321), .A2(n9388), .ZN(n7039) );
  NAND2_X1 U8012 ( .A1(n8321), .A2(n9388), .ZN(n7037) );
  NAND2_X1 U8013 ( .A1(n7039), .A2(n7037), .ZN(n8124) );
  AOI211_X1 U8014 ( .C1(n6724), .C2(n7038), .A(n6723), .B(n8124), .ZN(n6737)
         );
  INV_X1 U8015 ( .A(n7037), .ZN(n6735) );
  NAND2_X1 U8016 ( .A1(n7588), .A2(n6690), .ZN(n6726) );
  NAND2_X1 U8017 ( .A1(n6766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U8018 ( .A(n6738), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7859) );
  AOI22_X1 U8019 ( .A1(n6846), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6845), .B2(
        n7859), .ZN(n6725) );
  NAND2_X1 U8020 ( .A1(n6726), .A2(n6725), .ZN(n11112) );
  NAND2_X1 U8021 ( .A1(n6954), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6733) );
  INV_X1 U8022 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8023 ( .A1(n6969), .A2(n6727), .ZN(n6732) );
  INV_X1 U8024 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8294) );
  OR2_X1 U8025 ( .A1(n6973), .A2(n8294), .ZN(n6731) );
  AND2_X1 U8026 ( .A1(n6728), .A2(n7629), .ZN(n6729) );
  OR2_X1 U8027 ( .A1(n6729), .A2(n6744), .ZN(n9387) );
  OR2_X1 U8028 ( .A1(n6971), .A2(n9387), .ZN(n6730) );
  NAND4_X1 U8029 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n10329)
         );
  INV_X1 U8030 ( .A(n10329), .ZN(n8470) );
  OR2_X1 U8031 ( .A1(n11112), .A2(n8470), .ZN(n7041) );
  NAND2_X1 U8032 ( .A1(n7041), .A2(n7039), .ZN(n6734) );
  MUX2_X1 U8033 ( .A(n6735), .B(n6734), .S(n6949), .Z(n6736) );
  AND2_X1 U8034 ( .A1(n11112), .A2(n8470), .ZN(n6999) );
  NAND2_X1 U8035 ( .A1(n7591), .A2(n6690), .ZN(n6743) );
  INV_X1 U8036 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U8037 ( .A1(n6738), .A2(n8866), .ZN(n6739) );
  NAND2_X1 U8038 ( .A1(n6739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8039 ( .A1(n6740), .A2(n8872), .ZN(n6752) );
  OR2_X1 U8040 ( .A1(n6740), .A2(n8872), .ZN(n6741) );
  AOI22_X1 U8041 ( .A1(n6846), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6845), .B2(
        n10928), .ZN(n6742) );
  NAND2_X2 U8042 ( .A1(n6743), .A2(n6742), .ZN(n8473) );
  NAND2_X1 U8043 ( .A1(n6895), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6750) );
  INV_X1 U8044 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8135) );
  OR2_X1 U8045 ( .A1(n5133), .A2(n8135), .ZN(n6749) );
  NOR2_X1 U8046 ( .A1(n6744), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6745) );
  OR2_X1 U8047 ( .A1(n6757), .A2(n6745), .ZN(n8469) );
  OR2_X1 U8048 ( .A1(n6971), .A2(n8469), .ZN(n6748) );
  INV_X1 U8049 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6746) );
  OR2_X1 U8050 ( .A1(n6625), .A2(n6746), .ZN(n6747) );
  NAND4_X1 U8051 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n10328)
         );
  INV_X1 U8052 ( .A(n10328), .ZN(n8498) );
  OR2_X1 U8053 ( .A1(n8473), .A2(n8498), .ZN(n7111) );
  INV_X1 U8054 ( .A(n7111), .ZN(n6751) );
  NOR2_X1 U8055 ( .A1(n5175), .A2(n6751), .ZN(n6780) );
  NAND2_X1 U8056 ( .A1(n7596), .A2(n6690), .ZN(n6755) );
  NAND2_X1 U8057 ( .A1(n6752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6753) );
  XNOR2_X1 U8058 ( .A(n6753), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U8059 ( .A1(n6846), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6845), .B2(
        n10826), .ZN(n6754) );
  NAND2_X1 U8060 ( .A1(n6755), .A2(n6754), .ZN(n8457) );
  NAND2_X1 U8061 ( .A1(n6954), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6762) );
  INV_X1 U8062 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7860) );
  OR2_X1 U8063 ( .A1(n6924), .A2(n7860), .ZN(n6761) );
  INV_X1 U8064 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6756) );
  OR2_X1 U8065 ( .A1(n6973), .A2(n6756), .ZN(n6760) );
  OR2_X1 U8066 ( .A1(n6757), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8067 ( .A1(n6774), .A2(n6758), .ZN(n8497) );
  OR2_X1 U8068 ( .A1(n6971), .A2(n8497), .ZN(n6759) );
  NAND4_X1 U8069 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n10327)
         );
  INV_X1 U8070 ( .A(n10327), .ZN(n8983) );
  OR2_X1 U8071 ( .A1(n8457), .A2(n8983), .ZN(n7048) );
  OAI211_X1 U8072 ( .C1(n7046), .C2(n7041), .A(n7048), .B(n7111), .ZN(n6765)
         );
  NAND2_X1 U8073 ( .A1(n7111), .A2(n6999), .ZN(n6763) );
  AND2_X1 U8074 ( .A1(n6763), .A2(n8327), .ZN(n6764) );
  NAND2_X1 U8075 ( .A1(n8457), .A2(n8983), .ZN(n6998) );
  NAND2_X1 U8076 ( .A1(n6764), .A2(n6998), .ZN(n7115) );
  MUX2_X1 U8077 ( .A(n6765), .B(n7115), .S(n6949), .Z(n6824) );
  NAND2_X1 U8078 ( .A1(n7683), .A2(n6690), .ZN(n6770) );
  NAND2_X1 U8079 ( .A1(n6767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6768) );
  XNOR2_X1 U8080 ( .A(n6768), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U8081 ( .A1(n6846), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6845), .B2(
        n10390), .ZN(n6769) );
  NAND2_X1 U8082 ( .A1(n6954), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6779) );
  INV_X1 U8083 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6771) );
  OR2_X1 U8084 ( .A1(n6969), .A2(n6771), .ZN(n6778) );
  INV_X1 U8085 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6772) );
  OR2_X1 U8086 ( .A1(n5133), .A2(n6772), .ZN(n6777) );
  NAND2_X1 U8087 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NAND2_X1 U8088 ( .A1(n6789), .A2(n6775), .ZN(n8984) );
  OR2_X1 U8089 ( .A1(n6971), .A2(n8984), .ZN(n6776) );
  NAND4_X1 U8090 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n10326)
         );
  INV_X1 U8091 ( .A(n10326), .ZN(n9049) );
  OR2_X1 U8092 ( .A1(n8480), .A2(n9049), .ZN(n7050) );
  AND2_X1 U8093 ( .A1(n7050), .A2(n7048), .ZN(n7096) );
  OAI21_X1 U8094 ( .B1(n6780), .B2(n6824), .A(n7096), .ZN(n6797) );
  NAND2_X1 U8095 ( .A1(n7697), .A2(n6690), .ZN(n6786) );
  NAND2_X1 U8096 ( .A1(n6781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6782) );
  MUX2_X1 U8097 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6782), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6784) );
  INV_X1 U8098 ( .A(n6783), .ZN(n6798) );
  AND2_X1 U8099 ( .A1(n6784), .A2(n6798), .ZN(n10914) );
  AOI22_X1 U8100 ( .A1(n6846), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6845), .B2(
        n10914), .ZN(n6785) );
  NAND2_X1 U8101 ( .A1(n6954), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6795) );
  INV_X1 U8102 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10377) );
  OR2_X1 U8103 ( .A1(n6969), .A2(n10377), .ZN(n6794) );
  INV_X1 U8104 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6787) );
  OR2_X1 U8105 ( .A1(n6973), .A2(n6787), .ZN(n6793) );
  NAND2_X1 U8106 ( .A1(n6789), .A2(n6788), .ZN(n6791) );
  INV_X1 U8107 ( .A(n6804), .ZN(n6790) );
  NAND2_X1 U8108 ( .A1(n6791), .A2(n6790), .ZN(n9048) );
  OR2_X1 U8109 ( .A1(n6971), .A2(n9048), .ZN(n6792) );
  NAND4_X1 U8110 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n10325)
         );
  INV_X1 U8111 ( .A(n10325), .ZN(n9103) );
  NAND2_X1 U8112 ( .A1(n9043), .A2(n9103), .ZN(n6997) );
  NAND2_X1 U8113 ( .A1(n8480), .A2(n9049), .ZN(n6996) );
  AND2_X1 U8114 ( .A1(n6997), .A2(n6996), .ZN(n7095) );
  OR2_X1 U8115 ( .A1(n9043), .A2(n9103), .ZN(n7118) );
  INV_X1 U8116 ( .A(n7118), .ZN(n6796) );
  AOI21_X1 U8117 ( .B1(n6797), .B2(n7095), .A(n6796), .ZN(n6811) );
  NAND2_X1 U8118 ( .A1(n7722), .A2(n6690), .ZN(n6802) );
  NAND2_X1 U8119 ( .A1(n6798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6799) );
  MUX2_X1 U8120 ( .A(n6799), .B(P1_IR_REG_31__SCAN_IN), .S(n8873), .Z(n6800)
         );
  NAND2_X1 U8121 ( .A1(n6800), .A2(n6535), .ZN(n10393) );
  INV_X1 U8122 ( .A(n10393), .ZN(n10847) );
  AOI22_X1 U8123 ( .A1(n6846), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6845), .B2(
        n10847), .ZN(n6801) );
  OAI21_X1 U8124 ( .B1(n6804), .B2(P1_REG3_REG_14__SCAN_IN), .A(n6803), .ZN(
        n9102) );
  OR2_X1 U8125 ( .A1(n9102), .A2(n6971), .ZN(n6808) );
  NAND2_X1 U8126 ( .A1(n6954), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6807) );
  INV_X1 U8127 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10392) );
  OR2_X1 U8128 ( .A1(n6973), .A2(n10392), .ZN(n6806) );
  INV_X1 U8129 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10383) );
  OR2_X1 U8130 ( .A1(n6969), .A2(n10383), .ZN(n6805) );
  NAND4_X1 U8131 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n11210)
         );
  INV_X1 U8132 ( .A(n11210), .ZN(n10312) );
  OR2_X1 U8133 ( .A1(n9141), .A2(n10312), .ZN(n7119) );
  NAND2_X1 U8134 ( .A1(n9141), .A2(n10312), .ZN(n11206) );
  NAND2_X1 U8135 ( .A1(n7119), .A2(n11206), .ZN(n8946) );
  INV_X1 U8136 ( .A(n7119), .ZN(n6809) );
  NOR4_X1 U8137 ( .A1(n7122), .A2(n7123), .A3(n6809), .A4(n6985), .ZN(n6810)
         );
  OAI21_X1 U8138 ( .B1(n6811), .B2(n8946), .A(n6810), .ZN(n6812) );
  INV_X1 U8139 ( .A(n6812), .ZN(n6828) );
  NAND2_X1 U8140 ( .A1(n8030), .A2(n6690), .ZN(n6815) );
  XNOR2_X1 U8141 ( .A(n6813), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U8142 ( .A1(n6846), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6845), .B2(
        n10877), .ZN(n6814) );
  INV_X1 U8143 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8144 ( .A1(n6817), .A2(n6816), .ZN(n6819) );
  NAND2_X1 U8145 ( .A1(n6819), .A2(n6818), .ZN(n11241) );
  NOR2_X1 U8146 ( .A1(n11241), .A2(n6971), .ZN(n6823) );
  INV_X1 U8147 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U8148 ( .A1(n6622), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8149 ( .A1(n6954), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6820) );
  OAI211_X1 U8150 ( .C1(n6969), .C2(n10422), .A(n6821), .B(n6820), .ZN(n6822)
         );
  INV_X1 U8151 ( .A(n10595), .ZN(n10286) );
  NAND2_X1 U8152 ( .A1(n11260), .A2(n10286), .ZN(n6843) );
  NAND2_X1 U8153 ( .A1(n7129), .A2(n6843), .ZN(n11246) );
  NAND2_X1 U8154 ( .A1(n6995), .A2(n11206), .ZN(n7094) );
  INV_X1 U8155 ( .A(n6830), .ZN(n6862) );
  NAND2_X1 U8156 ( .A1(n8065), .A2(n6690), .ZN(n6837) );
  AND2_X1 U8157 ( .A1(n6831), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8158 ( .A1(n6832), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6835) );
  INV_X1 U8159 ( .A(n6832), .ZN(n6833) );
  INV_X1 U8160 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U8161 ( .A1(n6833), .A2(n8886), .ZN(n6834) );
  AND2_X1 U8162 ( .A1(n6835), .A2(n6834), .ZN(n10898) );
  AOI22_X1 U8163 ( .A1(n6846), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10898), 
        .B2(n6845), .ZN(n6836) );
  OAI21_X1 U8164 ( .B1(n6838), .B2(P1_REG3_REG_18__SCAN_IN), .A(n6851), .ZN(
        n10285) );
  INV_X1 U8165 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U8166 ( .A1(n6954), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8167 ( .A1(n6622), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6839) );
  OAI211_X1 U8168 ( .C1(n10427), .C2(n6969), .A(n6840), .B(n6839), .ZN(n6841)
         );
  INV_X1 U8169 ( .A(n6841), .ZN(n6842) );
  OAI21_X1 U8170 ( .B1(n10285), .B2(n6971), .A(n6842), .ZN(n11238) );
  INV_X1 U8171 ( .A(n11238), .ZN(n10241) );
  NOR2_X1 U8172 ( .A1(n10290), .A2(n10241), .ZN(n6859) );
  NAND2_X1 U8173 ( .A1(n7060), .A2(n7129), .ZN(n6844) );
  NAND2_X1 U8174 ( .A1(n10290), .A2(n10241), .ZN(n6994) );
  NAND2_X1 U8175 ( .A1(n6994), .A2(n6843), .ZN(n7130) );
  MUX2_X1 U8176 ( .A(n6844), .B(n7130), .S(n6949), .Z(n6861) );
  NAND2_X1 U8177 ( .A1(n8278), .A2(n6690), .ZN(n6848) );
  AOI22_X1 U8178 ( .A1(n6846), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10599), 
        .B2(n6845), .ZN(n6847) );
  INV_X1 U8179 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6850) );
  INV_X1 U8180 ( .A(n6849), .ZN(n6867) );
  AOI21_X1 U8181 ( .B1(n6851), .B2(n6850), .A(n6867), .ZN(n10189) );
  NAND2_X1 U8182 ( .A1(n10189), .A2(n6852), .ZN(n6858) );
  INV_X1 U8183 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8184 ( .A1(n6954), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8185 ( .A1(n6895), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6853) );
  OAI211_X1 U8186 ( .C1(n6855), .C2(n5133), .A(n6854), .B(n6853), .ZN(n6856)
         );
  INV_X1 U8187 ( .A(n6856), .ZN(n6857) );
  NAND2_X1 U8188 ( .A1(n6858), .A2(n6857), .ZN(n9222) );
  NAND2_X1 U8189 ( .A1(n10669), .A2(n10284), .ZN(n6992) );
  NOR2_X1 U8190 ( .A1(n10669), .A2(n10284), .ZN(n6874) );
  NOR2_X1 U8191 ( .A1(n6874), .A2(n6859), .ZN(n7137) );
  MUX2_X1 U8192 ( .A(n6994), .B(n7137), .S(n6949), .Z(n6860) );
  OAI211_X1 U8193 ( .C1(n6862), .C2(n6861), .A(n6992), .B(n6860), .ZN(n6873)
         );
  NAND2_X1 U8194 ( .A1(n8384), .A2(n6690), .ZN(n6864) );
  OR2_X1 U8195 ( .A1(n6982), .A2(n8823), .ZN(n6863) );
  NAND2_X1 U8196 ( .A1(n6895), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6871) );
  INV_X1 U8197 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6865) );
  OR2_X1 U8198 ( .A1(n6625), .A2(n6865), .ZN(n6870) );
  INV_X1 U8199 ( .A(n6883), .ZN(n6866) );
  OAI21_X1 U8200 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n6867), .A(n6866), .ZN(
        n10258) );
  OR2_X1 U8201 ( .A1(n6649), .A2(n10258), .ZN(n6869) );
  INV_X1 U8202 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9229) );
  OR2_X1 U8203 ( .A1(n5133), .A2(n9229), .ZN(n6868) );
  NAND4_X1 U8204 ( .A1(n6871), .A2(n6870), .A3(n6869), .A4(n6868), .ZN(n10571)
         );
  INV_X1 U8205 ( .A(n10571), .ZN(n10199) );
  INV_X1 U8206 ( .A(n6992), .ZN(n7135) );
  OAI21_X1 U8207 ( .B1(n9291), .B2(n7135), .A(n6949), .ZN(n6872) );
  NAND2_X1 U8208 ( .A1(n6873), .A2(n6872), .ZN(n6877) );
  INV_X1 U8209 ( .A(n6874), .ZN(n6993) );
  NAND2_X1 U8210 ( .A1(n7063), .A2(n6993), .ZN(n6875) );
  OAI21_X1 U8211 ( .B1(n6877), .B2(n6875), .A(n10565), .ZN(n6876) );
  NAND2_X1 U8212 ( .A1(n6876), .A2(n6985), .ZN(n6890) );
  NAND2_X1 U8213 ( .A1(n6877), .A2(n7063), .ZN(n6888) );
  NAND2_X1 U8214 ( .A1(n8300), .A2(n6690), .ZN(n6879) );
  INV_X1 U8215 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8301) );
  OR2_X1 U8216 ( .A1(n6982), .A2(n8301), .ZN(n6878) );
  NAND2_X1 U8217 ( .A1(n6954), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6887) );
  INV_X1 U8218 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6880) );
  OR2_X1 U8219 ( .A1(n6924), .A2(n6880), .ZN(n6886) );
  INV_X1 U8220 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6881) );
  OR2_X1 U8221 ( .A1(n6973), .A2(n6881), .ZN(n6885) );
  INV_X1 U8222 ( .A(n6882), .ZN(n6898) );
  OAI21_X1 U8223 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n6883), .A(n6898), .ZN(
        n10579) );
  OR2_X1 U8224 ( .A1(n6649), .A2(n10579), .ZN(n6884) );
  NAND4_X1 U8225 ( .A1(n6887), .A2(n6886), .A3(n6885), .A4(n6884), .ZN(n10550)
         );
  OR2_X1 U8226 ( .A1(n10582), .A2(n10271), .ZN(n7024) );
  NAND2_X1 U8227 ( .A1(n10582), .A2(n10271), .ZN(n9292) );
  NAND2_X1 U8228 ( .A1(n7024), .A2(n9292), .ZN(n10566) );
  NAND2_X1 U8229 ( .A1(n6890), .A2(n6889), .ZN(n6892) );
  MUX2_X1 U8230 ( .A(n7024), .B(n9292), .S(n6949), .Z(n6891) );
  NAND2_X1 U8231 ( .A1(n6892), .A2(n6891), .ZN(n6919) );
  NAND2_X1 U8232 ( .A1(n8378), .A2(n6690), .ZN(n6894) );
  OR2_X1 U8233 ( .A1(n6982), .A2(n8383), .ZN(n6893) );
  NAND2_X1 U8234 ( .A1(n6895), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6904) );
  INV_X1 U8235 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6896) );
  OR2_X1 U8236 ( .A1(n6625), .A2(n6896), .ZN(n6903) );
  INV_X1 U8237 ( .A(n6897), .ZN(n6911) );
  INV_X1 U8238 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U8239 ( .A1(n6898), .A2(n10270), .ZN(n6899) );
  NAND2_X1 U8240 ( .A1(n6911), .A2(n6899), .ZN(n10557) );
  OR2_X1 U8241 ( .A1(n6971), .A2(n10557), .ZN(n6902) );
  INV_X1 U8242 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6900) );
  OR2_X1 U8243 ( .A1(n5133), .A2(n6900), .ZN(n6901) );
  NAND4_X1 U8244 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n10570)
         );
  XNOR2_X1 U8245 ( .A(n10652), .B(n10570), .ZN(n10547) );
  NAND2_X1 U8246 ( .A1(n8506), .A2(n6690), .ZN(n6906) );
  OR2_X1 U8247 ( .A1(n6982), .A2(n8824), .ZN(n6905) );
  NAND2_X1 U8248 ( .A1(n6954), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6916) );
  INV_X1 U8249 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6907) );
  OR2_X1 U8250 ( .A1(n6969), .A2(n6907), .ZN(n6915) );
  INV_X1 U8251 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6908) );
  OR2_X1 U8252 ( .A1(n6973), .A2(n6908), .ZN(n6914) );
  INV_X1 U8253 ( .A(n6909), .ZN(n6926) );
  INV_X1 U8254 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8255 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8256 ( .A1(n6926), .A2(n6912), .ZN(n10531) );
  OR2_X1 U8257 ( .A1(n6649), .A2(n10531), .ZN(n6913) );
  NAND4_X1 U8258 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n10549)
         );
  INV_X1 U8259 ( .A(n10549), .ZN(n10272) );
  OR2_X1 U8260 ( .A1(n10646), .A2(n10272), .ZN(n6991) );
  INV_X1 U8261 ( .A(n10570), .ZN(n10200) );
  OR2_X1 U8262 ( .A1(n10652), .A2(n10200), .ZN(n6917) );
  NAND2_X1 U8263 ( .A1(n6991), .A2(n6917), .ZN(n7062) );
  NAND2_X1 U8264 ( .A1(n10646), .A2(n10272), .ZN(n9293) );
  NAND2_X1 U8265 ( .A1(n10652), .A2(n10200), .ZN(n10538) );
  NAND2_X1 U8266 ( .A1(n9293), .A2(n10538), .ZN(n7025) );
  MUX2_X1 U8267 ( .A(n7062), .B(n7025), .S(n6949), .Z(n6918) );
  AOI21_X1 U8268 ( .B1(n6919), .B2(n10547), .A(n6918), .ZN(n6934) );
  INV_X1 U8269 ( .A(n9293), .ZN(n10510) );
  INV_X1 U8270 ( .A(n6991), .ZN(n6920) );
  MUX2_X1 U8271 ( .A(n10510), .B(n6920), .S(n6949), .Z(n6933) );
  NAND2_X1 U8272 ( .A1(n9023), .A2(n6690), .ZN(n6922) );
  OR2_X1 U8273 ( .A1(n6982), .A2(n9024), .ZN(n6921) );
  NAND2_X1 U8274 ( .A1(n6954), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6932) );
  INV_X1 U8275 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6923) );
  OR2_X1 U8276 ( .A1(n6924), .A2(n6923), .ZN(n6931) );
  INV_X1 U8277 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6925) );
  OR2_X1 U8278 ( .A1(n5133), .A2(n6925), .ZN(n6930) );
  INV_X1 U8279 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U8280 ( .A1(n6926), .A2(n10250), .ZN(n6927) );
  NAND2_X1 U8281 ( .A1(n6928), .A2(n6927), .ZN(n10521) );
  OR2_X1 U8282 ( .A1(n6649), .A2(n10521), .ZN(n6929) );
  NAND4_X1 U8283 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n10541)
         );
  NAND2_X1 U8284 ( .A1(n10642), .A2(n10506), .ZN(n6946) );
  NOR2_X1 U8285 ( .A1(n10637), .A2(n10483), .ZN(n6948) );
  INV_X1 U8286 ( .A(n6948), .ZN(n7065) );
  NAND2_X1 U8287 ( .A1(n7065), .A2(n9295), .ZN(n10501) );
  NAND2_X1 U8288 ( .A1(n9175), .A2(n6690), .ZN(n6936) );
  OR2_X1 U8289 ( .A1(n6982), .A2(n9176), .ZN(n6935) );
  NAND2_X1 U8290 ( .A1(n6954), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6943) );
  INV_X1 U8291 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6937) );
  OR2_X1 U8292 ( .A1(n6969), .A2(n6937), .ZN(n6942) );
  INV_X1 U8293 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10464) );
  OR2_X1 U8294 ( .A1(n6958), .A2(n10464), .ZN(n6941) );
  INV_X1 U8295 ( .A(n6938), .ZN(n6939) );
  NAND2_X1 U8296 ( .A1(n6939), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6956) );
  OAI21_X1 U8297 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n6939), .A(n6956), .ZN(
        n10463) );
  OR2_X1 U8298 ( .A1(n6649), .A2(n10463), .ZN(n6940) );
  NAND4_X1 U8299 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n10323)
         );
  NAND2_X1 U8300 ( .A1(n10627), .A2(n10482), .ZN(n7074) );
  OAI21_X1 U8301 ( .B1(n6944), .B2(n10467), .A(n7074), .ZN(n6945) );
  INV_X1 U8302 ( .A(n6946), .ZN(n7068) );
  NAND2_X1 U8303 ( .A1(n6951), .A2(n6950), .ZN(n6964) );
  NAND2_X1 U8304 ( .A1(n9218), .A2(n6690), .ZN(n6953) );
  INV_X1 U8305 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9219) );
  OR2_X1 U8306 ( .A1(n6982), .A2(n9219), .ZN(n6952) );
  NAND2_X1 U8307 ( .A1(n6954), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6962) );
  INV_X1 U8308 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6955) );
  OR2_X1 U8309 ( .A1(n6969), .A2(n6955), .ZN(n6961) );
  INV_X1 U8310 ( .A(n6956), .ZN(n6970) );
  XNOR2_X1 U8311 ( .A(P1_REG3_REG_28__SCAN_IN), .B(n6970), .ZN(n10451) );
  INV_X1 U8312 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6957) );
  OR2_X1 U8313 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  OR2_X1 U8314 ( .A1(n10618), .A2(n10471), .ZN(n7021) );
  NAND2_X1 U8315 ( .A1(n10618), .A2(n10471), .ZN(n7073) );
  NAND2_X1 U8316 ( .A1(n7021), .A2(n7073), .ZN(n10455) );
  MUX2_X1 U8317 ( .A(n7021), .B(n7073), .S(n6949), .Z(n6963) );
  XNOR2_X1 U8318 ( .A(n6965), .B(SI_29_), .ZN(n10172) );
  NAND2_X1 U8319 ( .A1(n10172), .A2(n6690), .ZN(n6967) );
  OR2_X1 U8320 ( .A1(n6982), .A2(n10697), .ZN(n6966) );
  NAND2_X1 U8321 ( .A1(n6954), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6977) );
  INV_X1 U8322 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6968) );
  OR2_X1 U8323 ( .A1(n6969), .A2(n6968), .ZN(n6976) );
  NAND2_X1 U8324 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n6970), .ZN(n9316) );
  OR2_X1 U8325 ( .A1(n6971), .A2(n9316), .ZN(n6975) );
  INV_X1 U8326 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6972) );
  OR2_X1 U8327 ( .A1(n6958), .A2(n6972), .ZN(n6974) );
  NAND4_X1 U8328 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n10321)
         );
  INV_X1 U8329 ( .A(n10321), .ZN(n10447) );
  OR2_X1 U8330 ( .A1(n10614), .A2(n10447), .ZN(n7020) );
  NAND2_X1 U8331 ( .A1(n10614), .A2(n10447), .ZN(n7147) );
  NAND2_X1 U8332 ( .A1(n7020), .A2(n7147), .ZN(n9313) );
  MUX2_X1 U8333 ( .A(n7147), .B(n7020), .S(n6949), .Z(n6978) );
  XNOR2_X1 U8334 ( .A(n6981), .B(n6980), .ZN(n9412) );
  NAND2_X1 U8335 ( .A1(n9412), .A2(n6690), .ZN(n6984) );
  OR2_X1 U8336 ( .A1(n6982), .A2(n9272), .ZN(n6983) );
  AND2_X1 U8337 ( .A1(n10607), .A2(n6986), .ZN(n7082) );
  INV_X1 U8338 ( .A(n7082), .ZN(n7152) );
  NAND2_X1 U8339 ( .A1(n7153), .A2(n7152), .ZN(n6990) );
  NAND2_X1 U8340 ( .A1(n6987), .A2(n8890), .ZN(n7092) );
  AOI21_X1 U8341 ( .B1(n7082), .B2(n6949), .A(n7197), .ZN(n6989) );
  INV_X1 U8342 ( .A(n6990), .ZN(n7017) );
  INV_X1 U8343 ( .A(n10479), .ZN(n7013) );
  NAND2_X1 U8344 ( .A1(n6991), .A2(n9293), .ZN(n10537) );
  INV_X1 U8345 ( .A(n10547), .ZN(n10553) );
  INV_X1 U8346 ( .A(n7123), .ZN(n7055) );
  NAND2_X1 U8347 ( .A1(n7055), .A2(n6995), .ZN(n9143) );
  INV_X1 U8348 ( .A(n7122), .ZN(n7058) );
  NAND2_X1 U8349 ( .A1(n7048), .A2(n6998), .ZN(n8455) );
  NAND2_X2 U8350 ( .A1(n7111), .A2(n8327), .ZN(n8330) );
  INV_X1 U8351 ( .A(n6999), .ZN(n7044) );
  NAND2_X1 U8352 ( .A1(n7041), .A2(n7044), .ZN(n8284) );
  INV_X1 U8353 ( .A(n7001), .ZN(n8177) );
  AND2_X2 U8354 ( .A1(n8047), .A2(n7002), .ZN(n7909) );
  AND2_X1 U8355 ( .A1(n10338), .A2(n7651), .ZN(n7097) );
  NOR2_X1 U8356 ( .A1(n9254), .A2(n7097), .ZN(n7746) );
  NAND4_X1 U8357 ( .A1(n7909), .A2(n7746), .A3(n7197), .A4(n7922), .ZN(n7005)
         );
  NAND2_X2 U8358 ( .A1(n7003), .A2(n7029), .ZN(n8071) );
  NOR4_X1 U8359 ( .A1(n7005), .A2(n7004), .A3(n8071), .A4(n8096), .ZN(n7006)
         );
  NAND4_X1 U8360 ( .A1(n8181), .A2(n8352), .A3(n8116), .A4(n7006), .ZN(n7007)
         );
  NOR4_X1 U8361 ( .A1(n8455), .A2(n8330), .A3(n8284), .A4(n7007), .ZN(n7008)
         );
  NAND4_X1 U8362 ( .A1(n7053), .A2(n8458), .A3(n8483), .A4(n7008), .ZN(n7009)
         );
  NOR4_X1 U8363 ( .A1(n11246), .A2(n9143), .A3(n10592), .A4(n7009), .ZN(n7010)
         );
  NAND4_X1 U8364 ( .A1(n9180), .A2(n9146), .A3(n9306), .A4(n7010), .ZN(n7011)
         );
  NOR4_X1 U8365 ( .A1(n10537), .A2(n10553), .A3(n10566), .A4(n7011), .ZN(n7012) );
  NAND4_X1 U8366 ( .A1(n7013), .A2(n10516), .A3(n5513), .A4(n7012), .ZN(n7014)
         );
  NOR4_X1 U8367 ( .A1(n9313), .A2(n10455), .A3(n10467), .A4(n7014), .ZN(n7016)
         );
  NAND2_X1 U8368 ( .A1(n5448), .A2(n10320), .ZN(n7151) );
  NAND2_X1 U8369 ( .A1(n10443), .A2(n7015), .ZN(n7146) );
  NAND4_X1 U8370 ( .A1(n7017), .A2(n7016), .A3(n7151), .A4(n7146), .ZN(n7084)
         );
  NAND2_X1 U8371 ( .A1(n10599), .A2(n7197), .ZN(n7198) );
  NAND2_X1 U8372 ( .A1(n7198), .A2(n7642), .ZN(n7018) );
  INV_X1 U8373 ( .A(n7020), .ZN(n7023) );
  INV_X1 U8374 ( .A(n7021), .ZN(n7022) );
  NOR2_X1 U8375 ( .A1(n7023), .A2(n7022), .ZN(n7093) );
  INV_X1 U8376 ( .A(n7024), .ZN(n7064) );
  AOI21_X1 U8377 ( .B1(n10565), .B2(n9292), .A(n7064), .ZN(n7026) );
  NOR3_X1 U8378 ( .A1(n7068), .A2(n7026), .A3(n7025), .ZN(n7133) );
  INV_X1 U8379 ( .A(n8047), .ZN(n7027) );
  NAND2_X1 U8380 ( .A1(n8048), .A2(n7028), .ZN(n7030) );
  NAND2_X1 U8381 ( .A1(n7030), .A2(n7029), .ZN(n8097) );
  INV_X1 U8382 ( .A(n8097), .ZN(n7032) );
  INV_X1 U8383 ( .A(n8096), .ZN(n7031) );
  NAND2_X1 U8384 ( .A1(n7032), .A2(n7031), .ZN(n8094) );
  NAND2_X1 U8385 ( .A1(n8094), .A2(n7033), .ZN(n8077) );
  INV_X1 U8386 ( .A(n8077), .ZN(n7036) );
  NAND2_X1 U8387 ( .A1(n7036), .A2(n7035), .ZN(n8178) );
  NAND2_X1 U8388 ( .A1(n7037), .A2(n8179), .ZN(n7043) );
  NAND2_X1 U8389 ( .A1(n7043), .A2(n7039), .ZN(n8282) );
  NAND3_X1 U8390 ( .A1(n7039), .A2(n8177), .A3(n7038), .ZN(n7040) );
  NAND2_X1 U8391 ( .A1(n8282), .A2(n7040), .ZN(n7042) );
  INV_X1 U8392 ( .A(n8330), .ZN(n8130) );
  NOR2_X1 U8393 ( .A1(n8455), .A2(n7046), .ZN(n7047) );
  NAND2_X1 U8394 ( .A1(n8453), .A2(n8458), .ZN(n7051) );
  NAND2_X1 U8395 ( .A1(n7051), .A2(n7050), .ZN(n8477) );
  NAND2_X1 U8396 ( .A1(n8477), .A2(n8483), .ZN(n7052) );
  INV_X1 U8397 ( .A(n8945), .ZN(n7054) );
  NAND3_X1 U8398 ( .A1(n11207), .A2(n11208), .A3(n11206), .ZN(n7056) );
  NAND2_X1 U8399 ( .A1(n7056), .A2(n7055), .ZN(n10591) );
  INV_X1 U8400 ( .A(n10592), .ZN(n7057) );
  NAND2_X1 U8401 ( .A1(n10591), .A2(n7057), .ZN(n7059) );
  NAND2_X1 U8402 ( .A1(n7059), .A2(n7058), .ZN(n11230) );
  INV_X1 U8403 ( .A(n11246), .ZN(n11234) );
  INV_X1 U8404 ( .A(n9146), .ZN(n7061) );
  INV_X1 U8405 ( .A(n9180), .ZN(n9182) );
  AOI21_X1 U8406 ( .B1(n9293), .B2(n7062), .A(n5516), .ZN(n7067) );
  INV_X1 U8407 ( .A(n7063), .ZN(n9289) );
  OAI21_X1 U8408 ( .B1(n7064), .B2(n9289), .A(n7133), .ZN(n7066) );
  OAI211_X1 U8409 ( .C1(n7068), .C2(n7067), .A(n7066), .B(n7065), .ZN(n7141)
         );
  AOI21_X1 U8410 ( .B1(n7133), .B2(n9290), .A(n7141), .ZN(n7072) );
  INV_X1 U8411 ( .A(n7069), .ZN(n7071) );
  NOR2_X1 U8412 ( .A1(n7071), .A2(n7070), .ZN(n7145) );
  OAI21_X1 U8413 ( .B1(n7072), .B2(n7138), .A(n7145), .ZN(n7075) );
  INV_X1 U8414 ( .A(n7073), .ZN(n9299) );
  INV_X1 U8415 ( .A(n7074), .ZN(n9298) );
  NOR2_X1 U8416 ( .A1(n9299), .A2(n9298), .ZN(n7142) );
  NAND2_X1 U8417 ( .A1(n7075), .A2(n7142), .ZN(n7077) );
  INV_X1 U8418 ( .A(n7147), .ZN(n7076) );
  AOI21_X1 U8419 ( .B1(n7093), .B2(n7077), .A(n7076), .ZN(n7078) );
  NOR2_X1 U8420 ( .A1(n7078), .A2(n5448), .ZN(n7081) );
  INV_X1 U8421 ( .A(n7078), .ZN(n7079) );
  OAI22_X1 U8422 ( .A1(n7081), .A2(n7080), .B1(n10443), .B2(n7079), .ZN(n7083)
         );
  AOI211_X1 U8423 ( .C1(n7083), .C2(n7153), .A(n7082), .B(n7911), .ZN(n7086)
         );
  INV_X1 U8424 ( .A(n7084), .ZN(n7085) );
  OAI21_X1 U8425 ( .B1(n7086), .B2(n7085), .A(n7172), .ZN(n7087) );
  OAI211_X1 U8426 ( .C1(n7090), .C2(n7089), .A(n7088), .B(n7087), .ZN(n7159)
         );
  INV_X1 U8427 ( .A(n7093), .ZN(n7149) );
  INV_X1 U8428 ( .A(n7094), .ZN(n7125) );
  INV_X1 U8429 ( .A(n7095), .ZN(n7121) );
  INV_X1 U8430 ( .A(n7096), .ZN(n7117) );
  INV_X1 U8431 ( .A(n7097), .ZN(n7100) );
  INV_X1 U8432 ( .A(n9260), .ZN(n10987) );
  NAND2_X1 U8433 ( .A1(n10337), .A2(n10987), .ZN(n7099) );
  NAND3_X1 U8434 ( .A1(n7100), .A2(n7200), .A3(n7099), .ZN(n7101) );
  NAND2_X1 U8435 ( .A1(n5744), .A2(n7101), .ZN(n7102) );
  INV_X1 U8436 ( .A(n10336), .ZN(n7912) );
  OAI22_X1 U8437 ( .A1(n7921), .A2(n7102), .B1(n7912), .B2(n8925), .ZN(n7104)
         );
  AOI21_X1 U8438 ( .B1(n7104), .B2(n8047), .A(n7103), .ZN(n7107) );
  OR3_X1 U8439 ( .A1(n7107), .A2(n7106), .A3(n7105), .ZN(n7109) );
  NAND2_X1 U8440 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  NAND3_X1 U8441 ( .A1(n7110), .A2(n8282), .A3(n7035), .ZN(n7112) );
  AND3_X1 U8442 ( .A1(n7113), .A2(n7112), .A3(n7111), .ZN(n7114) );
  NOR2_X1 U8443 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  NOR2_X1 U8444 ( .A1(n7117), .A2(n7116), .ZN(n7120) );
  OAI211_X1 U8445 ( .C1(n7121), .C2(n7120), .A(n7119), .B(n7118), .ZN(n7124)
         );
  AOI211_X1 U8446 ( .C1(n7125), .C2(n7124), .A(n7123), .B(n7122), .ZN(n7128)
         );
  INV_X1 U8447 ( .A(n7126), .ZN(n7127) );
  NOR2_X1 U8448 ( .A1(n7128), .A2(n7127), .ZN(n7132) );
  INV_X1 U8449 ( .A(n7130), .ZN(n7131) );
  OAI21_X1 U8450 ( .B1(n7132), .B2(n5523), .A(n7131), .ZN(n7136) );
  INV_X1 U8451 ( .A(n7133), .ZN(n7134) );
  AOI211_X1 U8452 ( .C1(n7137), .C2(n7136), .A(n7135), .B(n7134), .ZN(n7140)
         );
  INV_X1 U8453 ( .A(n7138), .ZN(n7139) );
  OAI21_X1 U8454 ( .B1(n7141), .B2(n7140), .A(n7139), .ZN(n7144) );
  INV_X1 U8455 ( .A(n7142), .ZN(n7143) );
  AOI21_X1 U8456 ( .B1(n7145), .B2(n7144), .A(n7143), .ZN(n7148) );
  OAI211_X1 U8457 ( .C1(n7149), .C2(n7148), .A(n7147), .B(n7146), .ZN(n7150)
         );
  NAND3_X1 U8458 ( .A1(n7152), .A2(n7151), .A3(n7150), .ZN(n7154) );
  NAND2_X1 U8459 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  OR2_X1 U8460 ( .A1(n7580), .A2(P1_U3086), .ZN(n8507) );
  OAI21_X1 U8461 ( .B1(n7159), .B2(n7474), .A(n7158), .ZN(n7180) );
  NAND2_X1 U8462 ( .A1(n7163), .A2(n8899), .ZN(n7167) );
  NAND2_X1 U8463 ( .A1(n7165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U8464 ( .A1(n7167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7168) );
  INV_X1 U8465 ( .A(n7644), .ZN(n7173) );
  AND2_X1 U8466 ( .A1(n7173), .A2(n7649), .ZN(n7745) );
  NAND2_X1 U8467 ( .A1(n7639), .A2(n7745), .ZN(n7466) );
  NAND2_X1 U8468 ( .A1(n7174), .A2(n8903), .ZN(n7176) );
  NAND2_X1 U8469 ( .A1(n7176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8470 ( .A1(n7177), .A2(n7176), .ZN(n9177) );
  OR2_X1 U8471 ( .A1(n9220), .A2(n9177), .ZN(n7611) );
  NOR2_X1 U8472 ( .A1(n7466), .A2(n7611), .ZN(n7179) );
  OAI21_X1 U8473 ( .B1(n8507), .B2(n7196), .A(P1_B_REG_SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8474 ( .A1(n7180), .A2(n5735), .ZN(P1_U3242) );
  NOR2_X1 U8475 ( .A1(n5136), .A2(n8380), .ZN(n7181) );
  AND2_X1 U8476 ( .A1(n9618), .A2(n7181), .ZN(n7182) );
  NAND2_X1 U8477 ( .A1(n9580), .A2(n7183), .ZN(n7507) );
  NAND2_X1 U8478 ( .A1(n7988), .A2(n7507), .ZN(n7984) );
  OAI21_X1 U8479 ( .B1(n11179), .B2(n7484), .A(n7985), .ZN(n7184) );
  NAND2_X1 U8480 ( .A1(n7984), .A2(n7184), .ZN(n7189) );
  AND2_X1 U8481 ( .A1(n7185), .A2(n7539), .ZN(n7186) );
  NAND2_X1 U8482 ( .A1(n7187), .A2(n7186), .ZN(n7986) );
  AOI21_X1 U8483 ( .B1(n7988), .B2(n7983), .A(n7986), .ZN(n7188) );
  INV_X1 U8484 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7191) );
  NOR2_X1 U8485 ( .A1(n11187), .A2(n7191), .ZN(n7193) );
  NAND3_X1 U8486 ( .A1(n10599), .A2(n7200), .A3(n7474), .ZN(n7934) );
  NAND2_X2 U8487 ( .A1(n7197), .A2(n8381), .ZN(n7652) );
  NAND2_X1 U8488 ( .A1(n7200), .A2(n7647), .ZN(n7643) );
  NAND3_X1 U8489 ( .A1(n7198), .A2(n7652), .A3(n7643), .ZN(n7199) );
  NAND2_X1 U8490 ( .A1(n5134), .A2(n9259), .ZN(n7203) );
  AND2_X1 U8491 ( .A1(n7200), .A2(n7474), .ZN(n7201) );
  NAND2_X1 U8492 ( .A1(n10338), .A2(n7211), .ZN(n7202) );
  AND2_X1 U8493 ( .A1(n7203), .A2(n7202), .ZN(n7209) );
  INV_X1 U8494 ( .A(n7579), .ZN(n7205) );
  NAND2_X1 U8495 ( .A1(n7205), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U8496 ( .A1(n7209), .A2(n7204), .ZN(n7674) );
  NAND2_X1 U8497 ( .A1(n10338), .A2(n7232), .ZN(n7207) );
  AOI22_X1 U8498 ( .A1(n7211), .A2(n9259), .B1(n7205), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U8499 ( .A1(n7207), .A2(n7206), .ZN(n7672) );
  NAND2_X1 U8500 ( .A1(n7209), .A2(n9633), .ZN(n7210) );
  NAND2_X1 U8501 ( .A1(n7673), .A2(n7210), .ZN(n7216) );
  INV_X2 U8502 ( .A(n7255), .ZN(n7265) );
  NAND2_X1 U8503 ( .A1(n10337), .A2(n7265), .ZN(n7213) );
  NAND2_X1 U8504 ( .A1(n7218), .A2(n9260), .ZN(n7212) );
  NAND2_X1 U8505 ( .A1(n7213), .A2(n7212), .ZN(n7214) );
  NAND2_X1 U8506 ( .A1(n7216), .A2(n7215), .ZN(n7217) );
  AOI22_X1 U8507 ( .A1(n10337), .A2(n7232), .B1(n9635), .B2(n9260), .ZN(n7687)
         );
  NAND2_X1 U8508 ( .A1(n7685), .A2(n7709), .ZN(n7227) );
  NAND2_X1 U8509 ( .A1(n10336), .A2(n7265), .ZN(n7220) );
  NAND2_X1 U8510 ( .A1(n7218), .A2(n8925), .ZN(n7219) );
  NAND2_X1 U8511 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  XNOR2_X1 U8512 ( .A(n7221), .B(n9633), .ZN(n7222) );
  AOI22_X1 U8513 ( .A1(n10336), .A2(n7232), .B1(n9635), .B2(n8925), .ZN(n7223)
         );
  NAND2_X1 U8514 ( .A1(n7222), .A2(n7223), .ZN(n7228) );
  INV_X1 U8515 ( .A(n7222), .ZN(n7225) );
  INV_X1 U8516 ( .A(n7223), .ZN(n7224) );
  NAND2_X1 U8517 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  NAND2_X1 U8518 ( .A1(n7227), .A2(n7710), .ZN(n7712) );
  NAND2_X1 U8519 ( .A1(n7712), .A2(n7228), .ZN(n7727) );
  NAND2_X1 U8520 ( .A1(n10335), .A2(n7265), .ZN(n7230) );
  NAND2_X1 U8521 ( .A1(n7218), .A2(n7730), .ZN(n7229) );
  NAND2_X1 U8522 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  XNOR2_X1 U8523 ( .A(n7231), .B(n5138), .ZN(n7243) );
  AOI22_X1 U8524 ( .A1(n10335), .A2(n7232), .B1(n9635), .B2(n7730), .ZN(n7244)
         );
  XNOR2_X1 U8525 ( .A(n7243), .B(n7244), .ZN(n7728) );
  NAND2_X1 U8526 ( .A1(n7727), .A2(n7728), .ZN(n7726) );
  NAND2_X1 U8527 ( .A1(n10230), .A2(n7218), .ZN(n7234) );
  NAND2_X1 U8528 ( .A1(n10333), .A2(n7265), .ZN(n7233) );
  NAND2_X1 U8529 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  XNOR2_X1 U8530 ( .A(n7235), .B(n9633), .ZN(n10222) );
  NAND2_X1 U8531 ( .A1(n10230), .A2(n7265), .ZN(n7237) );
  NAND2_X1 U8532 ( .A1(n10333), .A2(n7232), .ZN(n7236) );
  AND2_X1 U8533 ( .A1(n7237), .A2(n7236), .ZN(n7249) );
  NAND2_X1 U8534 ( .A1(n10222), .A2(n7249), .ZN(n7247) );
  NAND2_X1 U8535 ( .A1(n10334), .A2(n7265), .ZN(n7239) );
  NAND2_X1 U8536 ( .A1(n7218), .A2(n8058), .ZN(n7238) );
  NAND2_X1 U8537 ( .A1(n7239), .A2(n7238), .ZN(n7240) );
  XNOR2_X1 U8538 ( .A(n7240), .B(n9633), .ZN(n7974) );
  NAND2_X1 U8539 ( .A1(n10334), .A2(n7232), .ZN(n7242) );
  NAND2_X1 U8540 ( .A1(n9635), .A2(n8058), .ZN(n7241) );
  AND2_X1 U8541 ( .A1(n7242), .A2(n7241), .ZN(n7973) );
  NAND2_X1 U8542 ( .A1(n7974), .A2(n7973), .ZN(n7246) );
  INV_X1 U8543 ( .A(n7243), .ZN(n7245) );
  NAND2_X1 U8544 ( .A1(n7245), .A2(n7244), .ZN(n7975) );
  NAND2_X1 U8545 ( .A1(n7726), .A2(n5746), .ZN(n7999) );
  INV_X1 U8546 ( .A(n10222), .ZN(n7251) );
  OR2_X1 U8547 ( .A1(n7974), .A2(n7973), .ZN(n7248) );
  NAND2_X1 U8548 ( .A1(n7248), .A2(n7249), .ZN(n7250) );
  INV_X1 U8549 ( .A(n7248), .ZN(n10219) );
  INV_X1 U8550 ( .A(n7249), .ZN(n10221) );
  AOI22_X1 U8551 ( .A1(n7251), .A2(n7250), .B1(n10219), .B2(n10221), .ZN(n7998) );
  NAND2_X1 U8552 ( .A1(n8119), .A2(n7218), .ZN(n7253) );
  NAND2_X1 U8553 ( .A1(n10332), .A2(n7265), .ZN(n7252) );
  NAND2_X1 U8554 ( .A1(n7253), .A2(n7252), .ZN(n7254) );
  XNOR2_X1 U8555 ( .A(n7254), .B(n9633), .ZN(n7260) );
  INV_X1 U8556 ( .A(n7260), .ZN(n7258) );
  INV_X2 U8557 ( .A(n7255), .ZN(n9635) );
  AND2_X1 U8558 ( .A1(n10332), .A2(n7232), .ZN(n7256) );
  AOI21_X1 U8559 ( .B1(n8119), .B2(n9635), .A(n7256), .ZN(n7259) );
  INV_X1 U8560 ( .A(n7259), .ZN(n7257) );
  NAND2_X1 U8561 ( .A1(n7258), .A2(n7257), .ZN(n8001) );
  NAND2_X1 U8562 ( .A1(n7260), .A2(n7259), .ZN(n8000) );
  INV_X1 U8563 ( .A(n8000), .ZN(n7261) );
  NAND2_X1 U8564 ( .A1(n8348), .A2(n7265), .ZN(n7264) );
  NAND2_X1 U8565 ( .A1(n10331), .A2(n7232), .ZN(n7263) );
  NAND2_X1 U8566 ( .A1(n7264), .A2(n7263), .ZN(n8041) );
  NAND2_X1 U8567 ( .A1(n8348), .A2(n7412), .ZN(n7267) );
  NAND2_X1 U8568 ( .A1(n10331), .A2(n7265), .ZN(n7266) );
  NAND2_X1 U8569 ( .A1(n7267), .A2(n7266), .ZN(n7268) );
  XNOR2_X1 U8570 ( .A(n7268), .B(n5138), .ZN(n8040) );
  NAND2_X1 U8571 ( .A1(n8321), .A2(n7412), .ZN(n7270) );
  NAND2_X1 U8572 ( .A1(n10330), .A2(n9635), .ZN(n7269) );
  NAND2_X1 U8573 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  XNOR2_X1 U8574 ( .A(n7271), .B(n9633), .ZN(n8314) );
  NAND2_X1 U8575 ( .A1(n8321), .A2(n9635), .ZN(n7273) );
  NAND2_X1 U8576 ( .A1(n10330), .A2(n7232), .ZN(n7272) );
  NAND2_X1 U8577 ( .A1(n8314), .A2(n8313), .ZN(n7274) );
  NAND2_X1 U8578 ( .A1(n11112), .A2(n7412), .ZN(n7276) );
  NAND2_X1 U8579 ( .A1(n10329), .A2(n9635), .ZN(n7275) );
  NAND2_X1 U8580 ( .A1(n7276), .A2(n7275), .ZN(n7277) );
  XNOR2_X1 U8581 ( .A(n7277), .B(n5138), .ZN(n7281) );
  AND2_X1 U8582 ( .A1(n10329), .A2(n7232), .ZN(n7278) );
  AOI21_X1 U8583 ( .B1(n11112), .B2(n9635), .A(n7278), .ZN(n7282) );
  XNOR2_X1 U8584 ( .A(n7281), .B(n7282), .ZN(n9382) );
  INV_X1 U8585 ( .A(n7281), .ZN(n7283) );
  NAND2_X1 U8586 ( .A1(n7283), .A2(n7282), .ZN(n7295) );
  NAND2_X1 U8587 ( .A1(n8473), .A2(n9635), .ZN(n7285) );
  NAND2_X1 U8588 ( .A1(n10328), .A2(n7232), .ZN(n7284) );
  NAND2_X1 U8589 ( .A1(n7285), .A2(n7284), .ZN(n8468) );
  INV_X1 U8590 ( .A(n8468), .ZN(n7286) );
  AND2_X1 U8591 ( .A1(n7295), .A2(n7286), .ZN(n7287) );
  NAND2_X1 U8592 ( .A1(n9384), .A2(n7287), .ZN(n7292) );
  NAND2_X1 U8593 ( .A1(n8473), .A2(n7412), .ZN(n7289) );
  NAND2_X1 U8594 ( .A1(n10328), .A2(n9635), .ZN(n7288) );
  NAND2_X1 U8595 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  XNOR2_X1 U8596 ( .A(n7290), .B(n9633), .ZN(n7296) );
  OR2_X1 U8597 ( .A1(n8468), .A2(n7296), .ZN(n7291) );
  NAND2_X1 U8598 ( .A1(n7292), .A2(n7291), .ZN(n7294) );
  INV_X1 U8599 ( .A(n7296), .ZN(n7293) );
  NAND2_X1 U8600 ( .A1(n7294), .A2(n8465), .ZN(n8466) );
  NAND2_X1 U8601 ( .A1(n9384), .A2(n7295), .ZN(n7297) );
  NAND2_X1 U8602 ( .A1(n7297), .A2(n7296), .ZN(n8491) );
  NAND2_X1 U8603 ( .A1(n8466), .A2(n8491), .ZN(n7307) );
  NAND2_X1 U8604 ( .A1(n8457), .A2(n7412), .ZN(n7299) );
  NAND2_X1 U8605 ( .A1(n10327), .A2(n9635), .ZN(n7298) );
  NAND2_X1 U8606 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  XNOR2_X1 U8607 ( .A(n7300), .B(n9633), .ZN(n7302) );
  AND2_X1 U8608 ( .A1(n10327), .A2(n7232), .ZN(n7301) );
  AOI21_X1 U8609 ( .B1(n8457), .B2(n9635), .A(n7301), .ZN(n7303) );
  NAND2_X1 U8610 ( .A1(n7302), .A2(n7303), .ZN(n8976) );
  INV_X1 U8611 ( .A(n7302), .ZN(n7305) );
  INV_X1 U8612 ( .A(n7303), .ZN(n7304) );
  NAND2_X1 U8613 ( .A1(n7305), .A2(n7304), .ZN(n7306) );
  AND2_X1 U8614 ( .A1(n8976), .A2(n7306), .ZN(n8492) );
  NAND2_X1 U8615 ( .A1(n7307), .A2(n8492), .ZN(n8495) );
  NAND2_X1 U8616 ( .A1(n8495), .A2(n8976), .ZN(n7317) );
  NAND2_X1 U8617 ( .A1(n8480), .A2(n7412), .ZN(n7309) );
  NAND2_X1 U8618 ( .A1(n10326), .A2(n9635), .ZN(n7308) );
  NAND2_X1 U8619 ( .A1(n7309), .A2(n7308), .ZN(n7310) );
  XNOR2_X1 U8620 ( .A(n7310), .B(n9633), .ZN(n7312) );
  AND2_X1 U8621 ( .A1(n10326), .A2(n7232), .ZN(n7311) );
  AOI21_X1 U8622 ( .B1(n8480), .B2(n9635), .A(n7311), .ZN(n7313) );
  NAND2_X1 U8623 ( .A1(n7312), .A2(n7313), .ZN(n7318) );
  INV_X1 U8624 ( .A(n7312), .ZN(n7315) );
  INV_X1 U8625 ( .A(n7313), .ZN(n7314) );
  NAND2_X1 U8626 ( .A1(n7315), .A2(n7314), .ZN(n7316) );
  AND2_X1 U8627 ( .A1(n7318), .A2(n7316), .ZN(n8977) );
  NAND2_X1 U8628 ( .A1(n9043), .A2(n7412), .ZN(n7320) );
  NAND2_X1 U8629 ( .A1(n10325), .A2(n9635), .ZN(n7319) );
  NAND2_X1 U8630 ( .A1(n7320), .A2(n7319), .ZN(n7321) );
  XNOR2_X1 U8631 ( .A(n7321), .B(n5138), .ZN(n7326) );
  AND2_X1 U8632 ( .A1(n10325), .A2(n7232), .ZN(n7322) );
  AOI21_X1 U8633 ( .B1(n9043), .B2(n9635), .A(n7322), .ZN(n7327) );
  XNOR2_X1 U8634 ( .A(n7326), .B(n7327), .ZN(n9046) );
  NAND2_X1 U8635 ( .A1(n9141), .A2(n7412), .ZN(n7324) );
  NAND2_X1 U8636 ( .A1(n11210), .A2(n9635), .ZN(n7323) );
  NAND2_X1 U8637 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  XNOR2_X1 U8638 ( .A(n7325), .B(n9633), .ZN(n7334) );
  INV_X1 U8639 ( .A(n7334), .ZN(n7329) );
  INV_X1 U8640 ( .A(n7326), .ZN(n7328) );
  NAND2_X1 U8641 ( .A1(n7328), .A2(n7327), .ZN(n7333) );
  NAND2_X1 U8642 ( .A1(n9141), .A2(n7265), .ZN(n7331) );
  NAND2_X1 U8643 ( .A1(n11210), .A2(n7232), .ZN(n7330) );
  NAND2_X1 U8644 ( .A1(n7331), .A2(n7330), .ZN(n9101) );
  INV_X1 U8645 ( .A(n9101), .ZN(n7332) );
  AND2_X1 U8646 ( .A1(n9096), .A2(n7332), .ZN(n7336) );
  NAND2_X1 U8647 ( .A1(n9045), .A2(n7333), .ZN(n7335) );
  NAND2_X1 U8648 ( .A1(n7335), .A2(n7334), .ZN(n9097) );
  NAND2_X1 U8649 ( .A1(n7336), .A2(n9097), .ZN(n9098) );
  NAND2_X1 U8650 ( .A1(n9098), .A2(n9097), .ZN(n7345) );
  INV_X1 U8651 ( .A(n7345), .ZN(n7343) );
  INV_X1 U8652 ( .A(n7337), .ZN(n7338) );
  NAND2_X1 U8653 ( .A1(n7337), .A2(n7412), .ZN(n7340) );
  NAND2_X1 U8654 ( .A1(n10594), .A2(n7265), .ZN(n7339) );
  NAND2_X1 U8655 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  XNOR2_X1 U8656 ( .A(n7341), .B(n9633), .ZN(n7344) );
  INV_X1 U8657 ( .A(n7344), .ZN(n7342) );
  AND2_X1 U8658 ( .A1(n10594), .A2(n7232), .ZN(n7347) );
  AOI21_X1 U8659 ( .B1(n7337), .B2(n9635), .A(n7347), .ZN(n10307) );
  NAND2_X1 U8660 ( .A1(n10602), .A2(n7412), .ZN(n7350) );
  NAND2_X1 U8661 ( .A1(n11235), .A2(n9635), .ZN(n7349) );
  NAND2_X1 U8662 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  XNOR2_X1 U8663 ( .A(n7351), .B(n5138), .ZN(n7363) );
  AND2_X1 U8664 ( .A1(n11235), .A2(n7232), .ZN(n7352) );
  AOI21_X1 U8665 ( .B1(n10602), .B2(n9635), .A(n7352), .ZN(n7364) );
  XNOR2_X1 U8666 ( .A(n7363), .B(n7364), .ZN(n10213) );
  NAND2_X1 U8667 ( .A1(n11260), .A2(n7412), .ZN(n7354) );
  NAND2_X1 U8668 ( .A1(n10595), .A2(n9635), .ZN(n7353) );
  NAND2_X1 U8669 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
  XNOR2_X1 U8670 ( .A(n7355), .B(n5138), .ZN(n7366) );
  NAND2_X1 U8671 ( .A1(n11260), .A2(n9635), .ZN(n7357) );
  NAND2_X1 U8672 ( .A1(n10595), .A2(n7232), .ZN(n7356) );
  NAND2_X1 U8673 ( .A1(n7357), .A2(n7356), .ZN(n7367) );
  NAND2_X1 U8674 ( .A1(n7366), .A2(n7367), .ZN(n10238) );
  AND2_X1 U8675 ( .A1(n10213), .A2(n10238), .ZN(n10277) );
  NAND2_X1 U8676 ( .A1(n10290), .A2(n7412), .ZN(n7359) );
  NAND2_X1 U8677 ( .A1(n11238), .A2(n7265), .ZN(n7358) );
  NAND2_X1 U8678 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  XNOR2_X1 U8679 ( .A(n7360), .B(n9633), .ZN(n7362) );
  AND2_X1 U8680 ( .A1(n10277), .A2(n7362), .ZN(n7361) );
  INV_X1 U8681 ( .A(n7362), .ZN(n7375) );
  INV_X1 U8682 ( .A(n10238), .ZN(n7371) );
  INV_X1 U8683 ( .A(n7363), .ZN(n7365) );
  NAND2_X1 U8684 ( .A1(n7365), .A2(n7364), .ZN(n10235) );
  INV_X1 U8685 ( .A(n7366), .ZN(n7369) );
  INV_X1 U8686 ( .A(n7367), .ZN(n7368) );
  NAND2_X1 U8687 ( .A1(n7369), .A2(n7368), .ZN(n10237) );
  AND2_X1 U8688 ( .A1(n10235), .A2(n10237), .ZN(n7370) );
  OR2_X1 U8689 ( .A1(n7371), .A2(n7370), .ZN(n7374) );
  AND2_X1 U8690 ( .A1(n11238), .A2(n7232), .ZN(n7372) );
  AOI21_X1 U8691 ( .B1(n10290), .B2(n5137), .A(n7372), .ZN(n10282) );
  AND2_X1 U8692 ( .A1(n10277), .A2(n10282), .ZN(n7373) );
  INV_X1 U8693 ( .A(n10282), .ZN(n7376) );
  AND2_X1 U8694 ( .A1(n7375), .A2(n7374), .ZN(n10278) );
  NAND2_X1 U8695 ( .A1(n10669), .A2(n7412), .ZN(n7378) );
  NAND2_X1 U8696 ( .A1(n9222), .A2(n5137), .ZN(n7377) );
  NAND2_X1 U8697 ( .A1(n7378), .A2(n7377), .ZN(n7379) );
  XNOR2_X1 U8698 ( .A(n7379), .B(n5138), .ZN(n7381) );
  AND2_X1 U8699 ( .A1(n9222), .A2(n7232), .ZN(n7380) );
  AOI21_X1 U8700 ( .B1(n10669), .B2(n5137), .A(n7380), .ZN(n7382) );
  XNOR2_X1 U8701 ( .A(n7381), .B(n7382), .ZN(n10187) );
  INV_X1 U8702 ( .A(n7381), .ZN(n7383) );
  NAND2_X1 U8703 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  NAND2_X1 U8704 ( .A1(n7385), .A2(n7384), .ZN(n10255) );
  NAND2_X1 U8705 ( .A1(n10664), .A2(n7412), .ZN(n7387) );
  NAND2_X1 U8706 ( .A1(n10571), .A2(n5137), .ZN(n7386) );
  NAND2_X1 U8707 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  XNOR2_X1 U8708 ( .A(n7388), .B(n5138), .ZN(n7390) );
  AND2_X1 U8709 ( .A1(n10571), .A2(n7232), .ZN(n7389) );
  AOI21_X1 U8710 ( .B1(n10664), .B2(n5137), .A(n7389), .ZN(n7391) );
  XNOR2_X1 U8711 ( .A(n7390), .B(n7391), .ZN(n10256) );
  NAND2_X1 U8712 ( .A1(n10255), .A2(n10256), .ZN(n7394) );
  INV_X1 U8713 ( .A(n7390), .ZN(n7392) );
  NAND2_X1 U8714 ( .A1(n7392), .A2(n7391), .ZN(n7393) );
  NAND2_X1 U8715 ( .A1(n10582), .A2(n7412), .ZN(n7396) );
  NAND2_X1 U8716 ( .A1(n10550), .A2(n5137), .ZN(n7395) );
  NAND2_X1 U8717 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  XNOR2_X1 U8718 ( .A(n7397), .B(n5138), .ZN(n7400) );
  NAND2_X1 U8719 ( .A1(n10582), .A2(n5137), .ZN(n7399) );
  NAND2_X1 U8720 ( .A1(n10550), .A2(n7232), .ZN(n7398) );
  NAND2_X1 U8721 ( .A1(n7399), .A2(n7398), .ZN(n7401) );
  NAND2_X1 U8722 ( .A1(n7400), .A2(n7401), .ZN(n7411) );
  INV_X1 U8723 ( .A(n7400), .ZN(n7403) );
  INV_X1 U8724 ( .A(n7401), .ZN(n7402) );
  NAND2_X1 U8725 ( .A1(n7403), .A2(n7402), .ZN(n7404) );
  NAND2_X1 U8726 ( .A1(n7411), .A2(n7404), .ZN(n10195) );
  NAND2_X1 U8727 ( .A1(n10652), .A2(n7412), .ZN(n7407) );
  NAND2_X1 U8728 ( .A1(n10570), .A2(n5137), .ZN(n7406) );
  NAND2_X1 U8729 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  XNOR2_X1 U8730 ( .A(n7408), .B(n9633), .ZN(n7410) );
  AND2_X1 U8731 ( .A1(n7410), .A2(n7411), .ZN(n7409) );
  AOI22_X1 U8732 ( .A1(n10652), .A2(n9635), .B1(n7232), .B2(n10570), .ZN(
        n10265) );
  NOR2_X1 U8733 ( .A1(n10263), .A2(n10265), .ZN(n10267) );
  AOI21_X1 U8734 ( .B1(n10197), .B2(n7411), .A(n7410), .ZN(n10264) );
  AOI22_X1 U8735 ( .A1(n10646), .A2(n9635), .B1(n7232), .B2(n10549), .ZN(n7415) );
  AOI22_X1 U8736 ( .A1(n10646), .A2(n7412), .B1(n5137), .B2(n10549), .ZN(n7413) );
  XNOR2_X1 U8737 ( .A(n7413), .B(n5138), .ZN(n7414) );
  XOR2_X1 U8738 ( .A(n7415), .B(n7414), .Z(n10181) );
  NAND2_X1 U8739 ( .A1(n10179), .A2(n10181), .ZN(n10180) );
  NAND2_X1 U8740 ( .A1(n10642), .A2(n7412), .ZN(n7418) );
  NAND2_X1 U8741 ( .A1(n10541), .A2(n5137), .ZN(n7417) );
  NAND2_X1 U8742 ( .A1(n7418), .A2(n7417), .ZN(n7419) );
  XNOR2_X1 U8743 ( .A(n7419), .B(n5138), .ZN(n7423) );
  NAND2_X1 U8744 ( .A1(n10642), .A2(n5137), .ZN(n7421) );
  NAND2_X1 U8745 ( .A1(n10541), .A2(n7232), .ZN(n7420) );
  NAND2_X1 U8746 ( .A1(n7421), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U8747 ( .A1(n7423), .A2(n7422), .ZN(n10248) );
  AOI22_X1 U8748 ( .A1(n10637), .A2(n9635), .B1(n7232), .B2(n10513), .ZN(n7431) );
  NAND2_X1 U8749 ( .A1(n10637), .A2(n7412), .ZN(n7425) );
  NAND2_X1 U8750 ( .A1(n10513), .A2(n5137), .ZN(n7424) );
  NAND2_X1 U8751 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  XNOR2_X1 U8752 ( .A(n7426), .B(n5138), .ZN(n7433) );
  XOR2_X1 U8753 ( .A(n7431), .B(n7433), .Z(n10205) );
  NAND2_X1 U8754 ( .A1(n10632), .A2(n7412), .ZN(n7428) );
  NAND2_X1 U8755 ( .A1(n10324), .A2(n5137), .ZN(n7427) );
  NAND2_X1 U8756 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  XNOR2_X1 U8757 ( .A(n7429), .B(n9633), .ZN(n7434) );
  AND2_X1 U8758 ( .A1(n10324), .A2(n7232), .ZN(n7430) );
  AOI21_X1 U8759 ( .B1(n10632), .B2(n5137), .A(n7430), .ZN(n7435) );
  XNOR2_X1 U8760 ( .A(n7434), .B(n7435), .ZN(n10295) );
  INV_X1 U8761 ( .A(n7431), .ZN(n7432) );
  NOR2_X1 U8762 ( .A1(n7433), .A2(n7432), .ZN(n10296) );
  INV_X1 U8763 ( .A(n7434), .ZN(n7437) );
  INV_X1 U8764 ( .A(n7435), .ZN(n7436) );
  AND2_X1 U8765 ( .A1(n7437), .A2(n7436), .ZN(n7445) );
  NAND2_X1 U8766 ( .A1(n10627), .A2(n7412), .ZN(n7439) );
  NAND2_X1 U8767 ( .A1(n10323), .A2(n5137), .ZN(n7438) );
  NAND2_X1 U8768 ( .A1(n7439), .A2(n7438), .ZN(n7440) );
  XNOR2_X1 U8769 ( .A(n7440), .B(n9633), .ZN(n7443) );
  AND2_X1 U8770 ( .A1(n10323), .A2(n7232), .ZN(n7441) );
  AOI21_X1 U8771 ( .B1(n10627), .B2(n5137), .A(n7441), .ZN(n7442) );
  NAND2_X1 U8772 ( .A1(n7443), .A2(n7442), .ZN(n9644) );
  OAI21_X1 U8773 ( .B1(n7443), .B2(n7442), .A(n9644), .ZN(n7444) );
  INV_X1 U8774 ( .A(n7446), .ZN(n7463) );
  NAND2_X1 U8775 ( .A1(n9056), .A2(P1_B_REG_SCAN_IN), .ZN(n7448) );
  INV_X1 U8776 ( .A(n9025), .ZN(n7447) );
  MUX2_X1 U8777 ( .A(n7448), .B(P1_B_REG_SCAN_IN), .S(n7447), .Z(n7449) );
  NAND2_X1 U8778 ( .A1(n9110), .A2(n9056), .ZN(n10687) );
  NOR4_X1 U8779 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n7458) );
  NOR4_X1 U8780 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n7457) );
  NOR4_X1 U8781 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n7453) );
  NOR4_X1 U8782 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n7452) );
  NOR4_X1 U8783 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7451) );
  NOR4_X1 U8784 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n7450) );
  NAND4_X1 U8785 ( .A1(n7453), .A2(n7452), .A3(n7451), .A4(n7450), .ZN(n7454)
         );
  NOR4_X1 U8786 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        n7455), .A4(n7454), .ZN(n7456) );
  AND3_X1 U8787 ( .A1(n7458), .A2(n7457), .A3(n7456), .ZN(n7459) );
  NOR2_X1 U8788 ( .A1(n7736), .A2(n7737), .ZN(n7461) );
  NAND2_X1 U8789 ( .A1(n7461), .A2(n8930), .ZN(n7473) );
  INV_X1 U8790 ( .A(n7652), .ZN(n7744) );
  AND2_X1 U8791 ( .A1(n11269), .A2(n7911), .ZN(n7464) );
  NAND2_X1 U8792 ( .A1(n7639), .A2(n7464), .ZN(n7462) );
  OAI21_X1 U8793 ( .B1(n9651), .B2(n7463), .A(n10308), .ZN(n7480) );
  NOR2_X1 U8794 ( .A1(n7473), .A2(n7466), .ZN(n7470) );
  INV_X1 U8795 ( .A(n9220), .ZN(n7627) );
  NAND2_X2 U8796 ( .A1(n7470), .A2(n7627), .ZN(n10313) );
  NOR2_X1 U8797 ( .A1(n10313), .A2(n10504), .ZN(n7472) );
  INV_X1 U8798 ( .A(n7464), .ZN(n7465) );
  OR2_X1 U8799 ( .A1(n7474), .A2(P1_U3086), .ZN(n8357) );
  NAND3_X1 U8800 ( .A1(n7466), .A2(n7465), .A3(n8357), .ZN(n7467) );
  NAND2_X1 U8801 ( .A1(n7473), .A2(n7467), .ZN(n7679) );
  NAND2_X1 U8802 ( .A1(n7644), .A2(n7649), .ZN(n7638) );
  AND3_X1 U8803 ( .A1(n7579), .A2(n7580), .A3(n7638), .ZN(n7468) );
  NAND2_X1 U8804 ( .A1(n7679), .A2(n7468), .ZN(n7469) );
  NAND2_X2 U8805 ( .A1(n7469), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10299) );
  OAI22_X1 U8806 ( .A1(n10299), .A2(n10463), .B1(n10471), .B2(n10300), .ZN(
        n7471) );
  AOI211_X1 U8807 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n7472), 
        .B(n7471), .ZN(n7479) );
  INV_X1 U8808 ( .A(n10627), .ZN(n10462) );
  INV_X1 U8809 ( .A(n7473), .ZN(n7477) );
  INV_X1 U8810 ( .A(n7639), .ZN(n7475) );
  OR2_X1 U8811 ( .A1(n7652), .A2(n7474), .ZN(n7743) );
  NOR2_X1 U8812 ( .A1(n7475), .A2(n7743), .ZN(n7476) );
  NAND2_X1 U8813 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  NAND3_X1 U8814 ( .A1(n7480), .A2(n7479), .A3(n5741), .ZN(P1_U3214) );
  NOR2_X4 U8815 ( .A1(n7579), .A2(n7482), .ZN(P1_U3973) );
  NAND3_X1 U8816 ( .A1(n7484), .A2(n7985), .A3(n7483), .ZN(n7487) );
  NAND2_X1 U8817 ( .A1(n7485), .A2(n8387), .ZN(n7486) );
  NAND2_X2 U8818 ( .A1(n7487), .A2(n7486), .ZN(n7783) );
  XNOR2_X1 U8819 ( .A(n7783), .B(n11027), .ZN(n7782) );
  XNOR2_X1 U8820 ( .A(n7782), .B(n9806), .ZN(n7504) );
  XNOR2_X1 U8821 ( .A(n7489), .B(n6103), .ZN(n7845) );
  MUX2_X1 U8822 ( .A(n7783), .B(n8390), .S(n7719), .Z(n7488) );
  INV_X1 U8823 ( .A(n7488), .ZN(n7846) );
  NAND2_X1 U8824 ( .A1(n7845), .A2(n7846), .ZN(n7844) );
  NAND2_X1 U8825 ( .A1(n7489), .A2(n6102), .ZN(n7490) );
  NAND2_X1 U8826 ( .A1(n7844), .A2(n7490), .ZN(n7811) );
  XNOR2_X1 U8827 ( .A(n7783), .B(n11008), .ZN(n7491) );
  XNOR2_X1 U8828 ( .A(n7491), .B(n5131), .ZN(n7812) );
  NAND2_X1 U8829 ( .A1(n7811), .A2(n7812), .ZN(n7501) );
  INV_X1 U8830 ( .A(n7491), .ZN(n7492) );
  NAND2_X1 U8831 ( .A1(n7492), .A2(n5131), .ZN(n7498) );
  NAND2_X1 U8832 ( .A1(n7501), .A2(n7498), .ZN(n7503) );
  INV_X1 U8833 ( .A(n7494), .ZN(n7493) );
  INV_X1 U8834 ( .A(n7519), .ZN(n7516) );
  NAND2_X1 U8835 ( .A1(n7493), .A2(n7516), .ZN(n7510) );
  AND2_X1 U8836 ( .A1(n7510), .A2(n7539), .ZN(n7497) );
  NAND3_X1 U8837 ( .A1(n9574), .A2(n7523), .A3(n11179), .ZN(n7495) );
  NAND2_X1 U8838 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  INV_X1 U8839 ( .A(n7504), .ZN(n7499) );
  AND2_X1 U8840 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  INV_X1 U8841 ( .A(n7786), .ZN(n7502) );
  AOI211_X1 U8842 ( .C1(n7504), .C2(n7503), .A(n9748), .B(n7502), .ZN(n7529)
         );
  INV_X1 U8843 ( .A(n7523), .ZN(n7505) );
  NAND2_X1 U8844 ( .A1(n7506), .A2(n7505), .ZN(n7512) );
  AND4_X1 U8845 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n7511)
         );
  NAND2_X1 U8846 ( .A1(n7512), .A2(n7511), .ZN(n7513) );
  NAND2_X1 U8847 ( .A1(n7513), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7518) );
  NOR2_X1 U8848 ( .A1(n7515), .A2(n7514), .ZN(n9625) );
  NAND2_X1 U8849 ( .A1(n9625), .A2(n7516), .ZN(n7517) );
  MUX2_X1 U8850 ( .A(n9766), .B(P2_U3151), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7528) );
  NAND2_X1 U8851 ( .A1(n9625), .A2(n7519), .ZN(n7522) );
  NOR2_X1 U8852 ( .A1(n9754), .A2(n9280), .ZN(n7527) );
  NAND2_X1 U8853 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  OAI22_X1 U8854 ( .A1(n5131), .A2(n9763), .B1(n9784), .B2(n11027), .ZN(n7526)
         );
  OR4_X1 U8855 ( .A1(n7529), .A2(n7528), .A3(n7527), .A4(n7526), .ZN(P2_U3158)
         );
  XNOR2_X1 U8856 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI222_X1 U8857 ( .A1(n5582), .A2(P2_U3151), .B1(n10175), .B2(n7533), .C1(
        n7531), .C2(n10173), .ZN(P2_U3292) );
  OAI222_X1 U8858 ( .A1(n10696), .A2(n7534), .B1(n9271), .B2(n7533), .C1(
        P1_U3086), .C2(n7617), .ZN(P1_U3352) );
  OAI222_X1 U8859 ( .A1(n10696), .A2(n7535), .B1(n9271), .B2(n7564), .C1(
        P1_U3086), .C2(n7613), .ZN(P1_U3353) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7536) );
  OAI222_X1 U8861 ( .A1(n10696), .A2(n7536), .B1(n9271), .B2(n7563), .C1(
        P1_U3086), .C2(n7614), .ZN(P1_U3354) );
  OAI222_X1 U8862 ( .A1(n10696), .A2(n7537), .B1(n9271), .B2(n7558), .C1(
        P1_U3086), .C2(n10363), .ZN(P1_U3351) );
  INV_X1 U8863 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7542) );
  INV_X1 U8864 ( .A(n7540), .ZN(n7541) );
  AOI22_X1 U8865 ( .A1(n7549), .A2(n7542), .B1(n7545), .B2(n7541), .ZN(
        P2_U3377) );
  INV_X1 U8866 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7546) );
  INV_X1 U8867 ( .A(n7543), .ZN(n7544) );
  AOI22_X1 U8868 ( .A1(n7549), .A2(n7546), .B1(n7545), .B2(n7544), .ZN(
        P2_U3376) );
  INV_X1 U8869 ( .A(n7547), .ZN(n7552) );
  INV_X1 U8870 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7548) );
  OAI222_X1 U8871 ( .A1(n5528), .A2(P2_U3151), .B1(n10175), .B2(n7552), .C1(
        n7548), .C2(n10173), .ZN(P2_U3290) );
  AND2_X1 U8872 ( .A1(n7549), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8873 ( .A1(n7549), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8874 ( .A1(n7549), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8875 ( .A1(n7549), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8876 ( .A1(n7549), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8877 ( .A1(n7549), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8878 ( .A1(n7549), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8879 ( .A1(n7549), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8880 ( .A1(n7549), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8881 ( .A1(n7549), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8882 ( .A1(n7549), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8883 ( .A1(n7549), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8884 ( .A1(n7549), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8885 ( .A1(n7549), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8886 ( .A1(n7549), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8887 ( .A1(n7549), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8888 ( .A1(n7549), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8889 ( .A1(n7549), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8890 ( .A1(n7549), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8891 ( .A1(n7549), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8892 ( .A1(n7549), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8893 ( .A1(n7549), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8894 ( .A1(n7549), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8895 ( .A1(n7549), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8896 ( .A1(n7549), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8897 ( .A1(n7549), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8898 ( .A1(n7549), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8899 ( .A1(n7549), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8900 ( .A1(n7549), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8901 ( .A1(n7549), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  NAND2_X1 U8902 ( .A1(n8390), .A2(P2_U3893), .ZN(n7550) );
  OAI21_X1 U8903 ( .B1(P2_U3893), .B2(n6609), .A(n7550), .ZN(P2_U3491) );
  INV_X1 U8904 ( .A(n10696), .ZN(n8066) );
  AOI22_X1 U8905 ( .A1(n10764), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n8066), .ZN(n7551) );
  OAI21_X1 U8906 ( .B1(n7552), .B2(n9271), .A(n7551), .ZN(P1_U3350) );
  INV_X1 U8907 ( .A(n7553), .ZN(n7567) );
  AOI22_X1 U8908 ( .A1(n10800), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n8066), .ZN(n7554) );
  OAI21_X1 U8909 ( .B1(n7567), .B2(n9271), .A(n7554), .ZN(P1_U3348) );
  INV_X1 U8910 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7556) );
  INV_X1 U8911 ( .A(n7555), .ZN(n7561) );
  INV_X1 U8912 ( .A(n10785), .ZN(n7605) );
  OAI222_X1 U8913 ( .A1(n10696), .A2(n7556), .B1(n9271), .B2(n7561), .C1(
        P1_U3086), .C2(n7605), .ZN(P1_U3349) );
  INV_X1 U8914 ( .A(n10175), .ZN(n9214) );
  INV_X1 U8915 ( .A(n9214), .ZN(n9275) );
  OAI222_X1 U8916 ( .A1(n7559), .A2(P2_U3151), .B1(n9275), .B2(n7558), .C1(
        n7557), .C2(n10173), .ZN(P2_U3291) );
  INV_X1 U8917 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7560) );
  OAI222_X1 U8918 ( .A1(n7837), .A2(P2_U3151), .B1(n9275), .B2(n7561), .C1(
        n7560), .C2(n10173), .ZN(P2_U3289) );
  INV_X1 U8919 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7562) );
  OAI222_X1 U8920 ( .A1(P2_U3151), .A2(n7901), .B1(n9275), .B2(n7563), .C1(
        n7562), .C2(n10173), .ZN(P2_U3294) );
  OAI222_X1 U8921 ( .A1(n10173), .A2(n7565), .B1(n9275), .B2(n7564), .C1(
        n10945), .C2(P2_U3151), .ZN(P2_U3293) );
  INV_X1 U8922 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7566) );
  OAI222_X1 U8923 ( .A1(n7568), .A2(P2_U3151), .B1(n9275), .B2(n7567), .C1(
        n7566), .C2(n10173), .ZN(P2_U3288) );
  INV_X1 U8924 ( .A(n7569), .ZN(n7572) );
  AOI22_X1 U8925 ( .A1(n10813), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n8066), .ZN(n7570) );
  OAI21_X1 U8926 ( .B1(n7572), .B2(n9271), .A(n7570), .ZN(P1_U3347) );
  OAI222_X1 U8927 ( .A1(n7573), .A2(P2_U3151), .B1(n9275), .B2(n7572), .C1(
        n7571), .C2(n10173), .ZN(P2_U3287) );
  NAND2_X1 U8928 ( .A1(n10704), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7575) );
  OAI21_X1 U8929 ( .B1(n10704), .B2(n7576), .A(n7575), .ZN(P1_U3439) );
  INV_X1 U8930 ( .A(n9177), .ZN(n9301) );
  NOR2_X1 U8931 ( .A1(n9220), .A2(n9301), .ZN(n7677) );
  NOR2_X1 U8932 ( .A1(n9220), .A2(n6603), .ZN(n7671) );
  AOI22_X1 U8933 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n7677), .B1(n7671), .B2(
        n9301), .ZN(n7577) );
  XOR2_X1 U8934 ( .A(P1_IR_REG_0__SCAN_IN), .B(n7577), .Z(n7587) );
  INV_X1 U8935 ( .A(n7580), .ZN(n7578) );
  OAI21_X1 U8936 ( .B1(n7579), .B2(n7578), .A(P1_STATE_REG_SCAN_IN), .ZN(n7585) );
  NAND2_X1 U8937 ( .A1(n7649), .A2(n7580), .ZN(n7582) );
  NAND2_X1 U8938 ( .A1(n7582), .A2(n7581), .ZN(n7583) );
  OR2_X1 U8939 ( .A1(n7585), .A2(n7583), .ZN(n7628) );
  INV_X1 U8940 ( .A(n7583), .ZN(n7584) );
  INV_X1 U8941 ( .A(n10933), .ZN(n10430) );
  AOI22_X1 U8942 ( .A1(n10430), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n7586) );
  OAI21_X1 U8943 ( .B1(n7587), .B2(n7628), .A(n7586), .ZN(P1_U3243) );
  INV_X1 U8944 ( .A(n7588), .ZN(n7590) );
  AOI22_X1 U8945 ( .A1(n8153), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n10169), .ZN(n7589) );
  OAI21_X1 U8946 ( .B1(n7590), .B2(n10175), .A(n7589), .ZN(P2_U3286) );
  INV_X1 U8947 ( .A(n7859), .ZN(n7631) );
  OAI222_X1 U8948 ( .A1(n9271), .A2(n7590), .B1(n7631), .B2(P1_U3086), .C1(
        n8842), .C2(n10696), .ZN(P1_U3346) );
  INV_X1 U8949 ( .A(n7591), .ZN(n7594) );
  AOI22_X1 U8950 ( .A1(n10928), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n8066), .ZN(n7592) );
  OAI21_X1 U8951 ( .B1(n7594), .B2(n9271), .A(n7592), .ZN(P1_U3345) );
  INV_X1 U8952 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7593) );
  OAI222_X1 U8953 ( .A1(P2_U3151), .A2(n7595), .B1(n9275), .B2(n7594), .C1(
        n7593), .C2(n10173), .ZN(P2_U3285) );
  NOR2_X1 U8954 ( .A1(n10430), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8955 ( .A(n7596), .ZN(n7656) );
  AOI22_X1 U8956 ( .A1(n10826), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n8066), .ZN(n7597) );
  OAI21_X1 U8957 ( .B1(n7656), .B2(n9271), .A(n7597), .ZN(P1_U3344) );
  NOR2_X1 U8958 ( .A1(n7859), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7598) );
  AOI21_X1 U8959 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7859), .A(n7598), .ZN(
        n7609) );
  INV_X1 U8960 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7599) );
  MUX2_X1 U8961 ( .A(n7599), .B(P1_REG2_REG_2__SCAN_IN), .S(n7613), .Z(n7662)
         );
  MUX2_X1 U8962 ( .A(n6614), .B(P1_REG2_REG_1__SCAN_IN), .S(n7614), .Z(n10341)
         );
  AND2_X1 U8963 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U8964 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  INV_X1 U8965 ( .A(n7614), .ZN(n10345) );
  NAND2_X1 U8966 ( .A1(n10345), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7600) );
  NAND2_X1 U8967 ( .A1(n10339), .A2(n7600), .ZN(n7661) );
  NAND2_X1 U8968 ( .A1(n7662), .A2(n7661), .ZN(n7660) );
  INV_X1 U8969 ( .A(n7613), .ZN(n7670) );
  NAND2_X1 U8970 ( .A1(n7670), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U8971 ( .A1(n7660), .A2(n7601), .ZN(n10351) );
  XNOR2_X1 U8972 ( .A(n7617), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U8973 ( .A1(n10351), .A2(n10352), .ZN(n10350) );
  INV_X1 U8974 ( .A(n7617), .ZN(n10359) );
  NAND2_X1 U8975 ( .A1(n10359), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U8976 ( .A1(n10350), .A2(n7602), .ZN(n10370) );
  XNOR2_X1 U8977 ( .A(n10363), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U8978 ( .A1(n10370), .A2(n10371), .ZN(n10369) );
  INV_X1 U8979 ( .A(n10363), .ZN(n7619) );
  NAND2_X1 U8980 ( .A1(n7619), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U8981 ( .A1(n10369), .A2(n7603), .ZN(n10762) );
  MUX2_X1 U8982 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6670), .S(n10764), .Z(n10763) );
  NAND2_X1 U8983 ( .A1(n10762), .A2(n10763), .ZN(n10761) );
  NAND2_X1 U8984 ( .A1(n10764), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7604) );
  AND2_X1 U8985 ( .A1(n10761), .A2(n7604), .ZN(n10777) );
  AOI22_X1 U8986 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n7605), .B1(n10785), .B2(
        n6679), .ZN(n10776) );
  NOR2_X1 U8987 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  AOI21_X1 U8988 ( .B1(n10785), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10778), .ZN(
        n10797) );
  NAND2_X1 U8989 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n10800), .ZN(n7606) );
  OAI21_X1 U8990 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n10800), .A(n7606), .ZN(
        n10796) );
  NOR2_X1 U8991 ( .A1(n10797), .A2(n10796), .ZN(n10795) );
  AOI21_X1 U8992 ( .B1(n10800), .B2(P1_REG2_REG_7__SCAN_IN), .A(n10795), .ZN(
        n10804) );
  NAND2_X1 U8993 ( .A1(n10813), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U8994 ( .B1(n10813), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7607), .ZN(
        n10805) );
  NOR2_X1 U8995 ( .A1(n10804), .A2(n10805), .ZN(n10806) );
  AOI21_X1 U8996 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10813), .A(n10806), .ZN(
        n7608) );
  NAND2_X1 U8997 ( .A1(n7609), .A2(n7608), .ZN(n7853) );
  OAI21_X1 U8998 ( .B1(n7609), .B2(n7608), .A(n7853), .ZN(n7610) );
  INV_X1 U8999 ( .A(n7610), .ZN(n7635) );
  INV_X1 U9000 ( .A(n7628), .ZN(n7626) );
  INV_X1 U9001 ( .A(n7611), .ZN(n7612) );
  AOI22_X1 U9002 ( .A1(n7859), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n6727), .B2(
        n7631), .ZN(n7625) );
  MUX2_X1 U9003 ( .A(n6623), .B(P1_REG1_REG_2__SCAN_IN), .S(n7613), .Z(n7665)
         );
  INV_X1 U9004 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10991) );
  MUX2_X1 U9005 ( .A(n10991), .B(P1_REG1_REG_1__SCAN_IN), .S(n7614), .Z(n10344) );
  AND2_X1 U9006 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10343) );
  NAND2_X1 U9007 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  NAND2_X1 U9008 ( .A1(n10345), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9009 ( .A1(n10342), .A2(n7615), .ZN(n7664) );
  NAND2_X1 U9010 ( .A1(n7665), .A2(n7664), .ZN(n7663) );
  NAND2_X1 U9011 ( .A1(n7670), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U9012 ( .A1(n7663), .A2(n7616), .ZN(n10354) );
  XNOR2_X1 U9013 ( .A(n7617), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U9014 ( .A1(n10354), .A2(n10355), .ZN(n10353) );
  NAND2_X1 U9015 ( .A1(n10359), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U9016 ( .A1(n10353), .A2(n7618), .ZN(n10367) );
  XNOR2_X1 U9017 ( .A(n10363), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U9018 ( .A1(n10367), .A2(n10368), .ZN(n10366) );
  NAND2_X1 U9019 ( .A1(n7619), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9020 ( .A1(n10366), .A2(n7620), .ZN(n10766) );
  MUX2_X1 U9021 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6669), .S(n10764), .Z(n10767) );
  NAND2_X1 U9022 ( .A1(n10766), .A2(n10767), .ZN(n10765) );
  NAND2_X1 U9023 ( .A1(n10764), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U9024 ( .A1(n10765), .A2(n7621), .ZN(n10783) );
  MUX2_X1 U9025 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6678), .S(n10785), .Z(n10784) );
  AND2_X1 U9026 ( .A1(n10783), .A2(n10784), .ZN(n10781) );
  AOI21_X1 U9027 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10785), .A(n10781), .ZN(
        n10794) );
  NAND2_X1 U9028 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n10800), .ZN(n7622) );
  OAI21_X1 U9029 ( .B1(n10800), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7622), .ZN(
        n10793) );
  NOR2_X1 U9030 ( .A1(n10794), .A2(n10793), .ZN(n10792) );
  AOI21_X1 U9031 ( .B1(n10800), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10792), .ZN(
        n10810) );
  NAND2_X1 U9032 ( .A1(n10813), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7623) );
  OAI21_X1 U9033 ( .B1(n10813), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7623), .ZN(
        n10811) );
  NOR2_X1 U9034 ( .A1(n10810), .A2(n10811), .ZN(n10809) );
  AOI21_X1 U9035 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10813), .A(n10809), .ZN(
        n7624) );
  NAND2_X1 U9036 ( .A1(n7625), .A2(n7624), .ZN(n7858) );
  OAI21_X1 U9037 ( .B1(n7625), .B2(n7624), .A(n7858), .ZN(n7633) );
  NAND2_X1 U9038 ( .A1(n7626), .A2(n9177), .ZN(n10918) );
  NOR2_X2 U9039 ( .A1(n7628), .A2(n7627), .ZN(n10929) );
  INV_X1 U9040 ( .A(n10929), .ZN(n10433) );
  NOR2_X1 U9041 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7629), .ZN(n9390) );
  AOI21_X1 U9042 ( .B1(n10430), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9390), .ZN(
        n7630) );
  OAI21_X1 U9043 ( .B1(n10433), .B2(n7631), .A(n7630), .ZN(n7632) );
  AOI21_X1 U9044 ( .B1(n7633), .B2(n10846), .A(n7632), .ZN(n7634) );
  OAI21_X1 U9045 ( .B1(n7635), .B2(n10922), .A(n7634), .ZN(P1_U3252) );
  NOR2_X1 U9046 ( .A1(n7737), .A2(n7636), .ZN(n7637) );
  INV_X1 U9047 ( .A(n8929), .ZN(n7640) );
  INV_X1 U9048 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7654) );
  INV_X1 U9049 ( .A(n7745), .ZN(n7646) );
  OAI22_X1 U9050 ( .A1(n7197), .A2(n7644), .B1(n10599), .B2(n8381), .ZN(n7645)
         );
  NAND2_X1 U9051 ( .A1(n7646), .A2(n7645), .ZN(n8947) );
  OR2_X1 U9052 ( .A1(n6949), .A2(n7647), .ZN(n11069) );
  INV_X1 U9053 ( .A(n7746), .ZN(n7648) );
  OAI21_X1 U9054 ( .B1(n11232), .B2(n11273), .A(n7648), .ZN(n7650) );
  NAND2_X1 U9055 ( .A1(n10337), .A2(n11237), .ZN(n7747) );
  OAI211_X1 U9056 ( .C1(n7652), .C2(n7651), .A(n7650), .B(n7747), .ZN(n10673)
         );
  NAND2_X1 U9057 ( .A1(n10673), .A2(n11280), .ZN(n7653) );
  OAI21_X1 U9058 ( .B1(n11280), .B2(n7654), .A(n7653), .ZN(P1_U3453) );
  OAI222_X1 U9059 ( .A1(n5391), .A2(P2_U3151), .B1(n9275), .B2(n7656), .C1(
        n7655), .C2(n10173), .ZN(P2_U3284) );
  NAND2_X1 U9060 ( .A1(n9222), .A2(P1_U3973), .ZN(n7657) );
  OAI21_X1 U9061 ( .B1(n6045), .B2(P1_U3973), .A(n7657), .ZN(P1_U3573) );
  INV_X1 U9062 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7659) );
  OAI22_X1 U9063 ( .A1(n10933), .A2(n7659), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7658), .ZN(n7669) );
  OAI21_X1 U9064 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7667) );
  OAI21_X1 U9065 ( .B1(n7665), .B2(n7664), .A(n7663), .ZN(n7666) );
  OAI22_X1 U9066 ( .A1(n10922), .A2(n7667), .B1(n10918), .B2(n7666), .ZN(n7668) );
  AOI211_X1 U9067 ( .C1(n7670), .C2(n10929), .A(n7669), .B(n7668), .ZN(n7678)
         );
  XOR2_X1 U9068 ( .A(P1_IR_REG_0__SCAN_IN), .B(n7671), .Z(n7676) );
  OAI21_X1 U9069 ( .B1(n7674), .B2(n7672), .A(n7673), .ZN(n7682) );
  NAND2_X1 U9070 ( .A1(n7682), .A2(n7677), .ZN(n7675) );
  OAI211_X1 U9071 ( .C1(n7677), .C2(n7676), .A(n7675), .B(P1_U3973), .ZN(
        n10374) );
  NAND2_X1 U9072 ( .A1(n7678), .A2(n10374), .ZN(P1_U3245) );
  NAND2_X1 U9073 ( .A1(n7679), .A2(n8929), .ZN(n7715) );
  AOI22_X1 U9074 ( .A1(n10315), .A2(n10337), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7715), .ZN(n7681) );
  NAND2_X1 U9075 ( .A1(n10289), .A2(n9259), .ZN(n7680) );
  OAI211_X1 U9076 ( .C1(n10292), .C2(n7682), .A(n7681), .B(n7680), .ZN(
        P1_U3232) );
  INV_X1 U9077 ( .A(n7683), .ZN(n7695) );
  INV_X1 U9078 ( .A(n10390), .ZN(n7864) );
  INV_X1 U9079 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7684) );
  OAI222_X1 U9080 ( .A1(n9271), .A2(n7695), .B1(n7864), .B2(P1_U3086), .C1(
        n7684), .C2(n10696), .ZN(P1_U3343) );
  OAI21_X1 U9081 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n7692) );
  INV_X1 U9082 ( .A(n7715), .ZN(n7688) );
  OAI22_X1 U9083 ( .A1(n7688), .A2(n6611), .B1(n10318), .B2(n10987), .ZN(n7691) );
  INV_X1 U9084 ( .A(n10338), .ZN(n7689) );
  OAI22_X1 U9085 ( .A1(n7689), .A2(n10313), .B1(n10300), .B2(n7912), .ZN(n7690) );
  AOI211_X1 U9086 ( .C1(n7692), .C2(n10308), .A(n7691), .B(n7690), .ZN(n7693)
         );
  INV_X1 U9087 ( .A(n7693), .ZN(P1_U3222) );
  INV_X1 U9088 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7694) );
  OAI222_X1 U9089 ( .A1(P2_U3151), .A2(n7696), .B1(n9275), .B2(n7695), .C1(
        n7694), .C2(n10173), .ZN(P2_U3283) );
  INV_X1 U9090 ( .A(n7697), .ZN(n7700) );
  AOI22_X1 U9091 ( .A1(n9130), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n10169), .ZN(n7698) );
  OAI21_X1 U9092 ( .B1(n7700), .B2(n9275), .A(n7698), .ZN(P2_U3282) );
  AOI22_X1 U9093 ( .A1(n10914), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n8066), .ZN(n7699) );
  OAI21_X1 U9094 ( .B1(n7700), .B2(n9271), .A(n7699), .ZN(P1_U3342) );
  INV_X1 U9095 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U9096 ( .A1(n9881), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9097 ( .A1(n7701), .A2(n10939), .ZN(n7705) );
  INV_X1 U9098 ( .A(n7892), .ZN(n7702) );
  OAI21_X1 U9099 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7703), .A(n7702), .ZN(n7704) );
  AOI22_X1 U9100 ( .A1(n7705), .A2(n7704), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7706) );
  OAI211_X1 U9101 ( .C1(n9873), .C2(n7708), .A(n7707), .B(n7706), .ZN(P2_U3182) );
  INV_X1 U9102 ( .A(n7709), .ZN(n7711) );
  NOR2_X1 U9103 ( .A1(n7711), .A2(n7710), .ZN(n7714) );
  INV_X1 U9104 ( .A(n7712), .ZN(n7713) );
  AOI21_X1 U9105 ( .B1(n7714), .B2(n7685), .A(n7713), .ZN(n7718) );
  AOI22_X1 U9106 ( .A1(n10289), .A2(n8925), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7715), .ZN(n7717) );
  INV_X1 U9107 ( .A(n10313), .ZN(n9641) );
  AOI22_X1 U9108 ( .A1(n9641), .A2(n10337), .B1(n10315), .B2(n10335), .ZN(
        n7716) );
  OAI211_X1 U9109 ( .C1(n7718), .C2(n10292), .A(n7717), .B(n7716), .ZN(
        P1_U3237) );
  NAND2_X1 U9110 ( .A1(n9779), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7841) );
  NAND2_X1 U9111 ( .A1(n7841), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7721) );
  INV_X1 U9112 ( .A(n8394), .ZN(n9433) );
  NAND2_X1 U9113 ( .A1(n8390), .A2(n8034), .ZN(n9442) );
  NAND2_X1 U9114 ( .A1(n9433), .A2(n9442), .ZN(n9588) );
  AOI22_X1 U9115 ( .A1(n9773), .A2(n9588), .B1(n9731), .B2(n7719), .ZN(n7720)
         );
  OAI211_X1 U9116 ( .C1(n6102), .C2(n9754), .A(n7721), .B(n7720), .ZN(P2_U3172) );
  INV_X1 U9117 ( .A(n7722), .ZN(n7725) );
  OAI222_X1 U9118 ( .A1(n7724), .A2(P2_U3151), .B1(n9275), .B2(n7725), .C1(
        n7723), .C2(n10173), .ZN(P2_U3281) );
  OAI222_X1 U9119 ( .A1(n10696), .A2(n8630), .B1(n9271), .B2(n7725), .C1(
        P1_U3086), .C2(n10393), .ZN(P1_U3341) );
  OAI21_X1 U9120 ( .B1(n7728), .B2(n7727), .A(n7726), .ZN(n7734) );
  AOI22_X1 U9121 ( .A1(n10315), .A2(n10334), .B1(n9641), .B2(n10336), .ZN(
        n7732) );
  NAND2_X1 U9122 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10356) );
  INV_X1 U9123 ( .A(n10356), .ZN(n7729) );
  AOI21_X1 U9124 ( .B1(n10289), .B2(n7730), .A(n7729), .ZN(n7731) );
  OAI211_X1 U9125 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10299), .A(n7732), .B(
        n7731), .ZN(n7733) );
  AOI21_X1 U9126 ( .B1(n7734), .B2(n10308), .A(n7733), .ZN(n7735) );
  INV_X1 U9127 ( .A(n7735), .ZN(P1_U3218) );
  INV_X1 U9128 ( .A(n7736), .ZN(n7739) );
  INV_X1 U9129 ( .A(n7737), .ZN(n7738) );
  INV_X1 U9130 ( .A(n8930), .ZN(n7740) );
  NAND2_X1 U9131 ( .A1(n10560), .A2(n11250), .ZN(n9330) );
  INV_X1 U9132 ( .A(n9330), .ZN(n10545) );
  OAI21_X1 U9133 ( .B1(n10545), .B2(n11245), .A(n9259), .ZN(n7752) );
  NOR3_X1 U9134 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(n7750) );
  OAI21_X1 U9135 ( .B1(n10580), .B2(n7748), .A(n7747), .ZN(n7749) );
  OAI21_X1 U9136 ( .B1(n7750), .B2(n7749), .A(n10600), .ZN(n7751) );
  OAI211_X1 U9137 ( .C1(n6603), .C2(n10600), .A(n7752), .B(n7751), .ZN(
        P1_U3293) );
  AOI211_X1 U9138 ( .C1(n7755), .C2(n7754), .A(n10939), .B(n7753), .ZN(n7756)
         );
  INV_X1 U9139 ( .A(n7756), .ZN(n7765) );
  INV_X1 U9140 ( .A(n7825), .ZN(n7757) );
  AOI21_X1 U9141 ( .B1(n9284), .B2(n7758), .A(n7757), .ZN(n7762) );
  OAI21_X1 U9142 ( .B1(n7759), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7830), .ZN(
        n7760) );
  NAND2_X1 U9143 ( .A1(n7760), .A2(n5874), .ZN(n7761) );
  NAND2_X1 U9144 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7944) );
  OAI211_X1 U9145 ( .C1(n7762), .C2(n10972), .A(n7761), .B(n7944), .ZN(n7763)
         );
  AOI21_X1 U9146 ( .B1(n10959), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7763), .ZN(
        n7764) );
  OAI211_X1 U9147 ( .C1(n5947), .C2(n5528), .A(n7765), .B(n7764), .ZN(P2_U3187) );
  OAI21_X1 U9148 ( .B1(n7767), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7766), .ZN(
        n7775) );
  INV_X1 U9149 ( .A(n7952), .ZN(n7768) );
  AOI21_X1 U9150 ( .B1(n7770), .B2(n7769), .A(n7768), .ZN(n7771) );
  OAI22_X1 U9151 ( .A1(n10972), .A2(n7771), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8763), .ZN(n7774) );
  INV_X1 U9152 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7772) );
  NOR2_X1 U9153 ( .A1(n9873), .A2(n7772), .ZN(n7773) );
  AOI211_X1 U9154 ( .C1(n5874), .C2(n7775), .A(n7774), .B(n7773), .ZN(n7781)
         );
  OAI21_X1 U9155 ( .B1(n7778), .B2(n7777), .A(n7776), .ZN(n7779) );
  NAND2_X1 U9156 ( .A1(n7779), .A2(n5272), .ZN(n7780) );
  OAI211_X1 U9157 ( .C1(n5947), .C2(n5582), .A(n7781), .B(n7780), .ZN(P2_U3185) );
  NAND2_X1 U9158 ( .A1(n7782), .A2(n9806), .ZN(n7784) );
  AND2_X1 U9159 ( .A1(n7786), .A2(n7784), .ZN(n7788) );
  XNOR2_X1 U9160 ( .A(n7783), .B(n11035), .ZN(n7939) );
  XNOR2_X1 U9161 ( .A(n7939), .B(n9280), .ZN(n7787) );
  AND2_X1 U9162 ( .A1(n7787), .A2(n7784), .ZN(n7785) );
  NAND2_X1 U9163 ( .A1(n7786), .A2(n7785), .ZN(n7942) );
  OAI21_X1 U9164 ( .B1(n7788), .B2(n7787), .A(n7942), .ZN(n7789) );
  NAND2_X1 U9165 ( .A1(n7789), .A2(n9773), .ZN(n7794) );
  NOR2_X1 U9166 ( .A1(n9754), .A2(n8025), .ZN(n7792) );
  AND2_X1 U9167 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7955) );
  AOI21_X1 U9168 ( .B1(n9731), .B2(n8247), .A(n7955), .ZN(n7790) );
  OAI21_X1 U9169 ( .B1(n9763), .B2(n11002), .A(n7790), .ZN(n7791) );
  AOI211_X1 U9170 ( .C1(n8246), .C2(n9766), .A(n7792), .B(n7791), .ZN(n7793)
         );
  NAND2_X1 U9171 ( .A1(n7794), .A2(n7793), .ZN(P2_U3170) );
  AOI21_X1 U9172 ( .B1(n11091), .B2(n7796), .A(n7795), .ZN(n7810) );
  OAI21_X1 U9173 ( .B1(n7799), .B2(n7798), .A(n7797), .ZN(n7800) );
  NAND2_X1 U9174 ( .A1(n7800), .A2(n5272), .ZN(n7809) );
  NAND2_X1 U9175 ( .A1(n7801), .A2(n8221), .ZN(n7802) );
  AOI21_X1 U9176 ( .B1(n7803), .B2(n7802), .A(n10972), .ZN(n7806) );
  INV_X1 U9177 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U9178 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8111) );
  OAI21_X1 U9179 ( .B1(n9873), .B2(n7804), .A(n8111), .ZN(n7805) );
  AOI211_X1 U9180 ( .C1(n9881), .C2(n7807), .A(n7806), .B(n7805), .ZN(n7808)
         );
  OAI211_X1 U9181 ( .C1(n7810), .C2(n10967), .A(n7809), .B(n7808), .ZN(
        P2_U3189) );
  XOR2_X1 U9182 ( .A(n7812), .B(n7811), .Z(n7816) );
  NOR2_X1 U9183 ( .A1(n9754), .A2(n11002), .ZN(n7814) );
  OAI22_X1 U9184 ( .A1(n6102), .A2(n9763), .B1(n9784), .B2(n11008), .ZN(n7813)
         );
  AOI211_X1 U9185 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7841), .A(n7814), .B(
        n7813), .ZN(n7815) );
  OAI21_X1 U9186 ( .B1(n7816), .B2(n9748), .A(n7815), .ZN(P2_U3177) );
  OAI21_X1 U9187 ( .B1(n5181), .B2(n7818), .A(n7817), .ZN(n7819) );
  NAND2_X1 U9188 ( .A1(n7819), .A2(n5272), .ZN(n7836) );
  INV_X1 U9189 ( .A(n7820), .ZN(n7822) );
  NOR2_X1 U9190 ( .A1(n7822), .A2(n7821), .ZN(n7826) );
  INV_X1 U9191 ( .A(n7823), .ZN(n7824) );
  AOI21_X1 U9192 ( .B1(n7826), .B2(n7825), .A(n7824), .ZN(n7827) );
  NAND2_X1 U9193 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8024) );
  OAI21_X1 U9194 ( .B1(n10972), .B2(n7827), .A(n8024), .ZN(n7834) );
  INV_X1 U9195 ( .A(n7828), .ZN(n7832) );
  NAND3_X1 U9196 ( .A1(n7830), .A2(n7829), .A3(n5163), .ZN(n7831) );
  AOI21_X1 U9197 ( .B1(n7832), .B2(n7831), .A(n10967), .ZN(n7833) );
  AOI211_X1 U9198 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10959), .A(n7834), .B(
        n7833), .ZN(n7835) );
  OAI211_X1 U9199 ( .C1(n5947), .C2(n7837), .A(n7836), .B(n7835), .ZN(P2_U3188) );
  INV_X1 U9200 ( .A(n6585), .ZN(n7840) );
  AOI22_X1 U9201 ( .A1(n10859), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n8066), .ZN(n7838) );
  OAI21_X1 U9202 ( .B1(n7840), .B2(n9271), .A(n7838), .ZN(P1_U3340) );
  AOI22_X1 U9203 ( .A1(n9839), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n10169), .ZN(n7839) );
  OAI21_X1 U9204 ( .B1(n7840), .B2(n9275), .A(n7839), .ZN(P2_U3280) );
  INV_X1 U9205 ( .A(n7841), .ZN(n7850) );
  INV_X1 U9206 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8395) );
  INV_X1 U9207 ( .A(n8390), .ZN(n7842) );
  OAI22_X1 U9208 ( .A1(n7842), .A2(n9763), .B1(n9784), .B2(n8396), .ZN(n7843)
         );
  AOI21_X1 U9209 ( .B1(n9781), .B2(n9807), .A(n7843), .ZN(n7849) );
  OAI21_X1 U9210 ( .B1(n7846), .B2(n7845), .A(n7844), .ZN(n7847) );
  NAND2_X1 U9211 ( .A1(n7847), .A2(n9773), .ZN(n7848) );
  OAI211_X1 U9212 ( .C1(n7850), .C2(n8395), .A(n7849), .B(n7848), .ZN(P2_U3162) );
  NOR2_X1 U9213 ( .A1(n10390), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7851) );
  AOI21_X1 U9214 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10390), .A(n7851), .ZN(
        n7856) );
  NAND2_X1 U9215 ( .A1(n10928), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7852) );
  OAI21_X1 U9216 ( .B1(n10928), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7852), .ZN(
        n10924) );
  OAI21_X1 U9217 ( .B1(n7859), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7853), .ZN(
        n10925) );
  NOR2_X1 U9218 ( .A1(n10924), .A2(n10925), .ZN(n10923) );
  AOI21_X1 U9219 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10928), .A(n10923), .ZN(
        n10821) );
  NAND2_X1 U9220 ( .A1(n10826), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7854) );
  OAI21_X1 U9221 ( .B1(n10826), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7854), .ZN(
        n10822) );
  NOR2_X1 U9222 ( .A1(n10821), .A2(n10822), .ZN(n10823) );
  AOI21_X1 U9223 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10826), .A(n10823), .ZN(
        n7855) );
  NAND2_X1 U9224 ( .A1(n7856), .A2(n7855), .ZN(n10389) );
  OAI21_X1 U9225 ( .B1(n7856), .B2(n7855), .A(n10389), .ZN(n7857) );
  INV_X1 U9226 ( .A(n7857), .ZN(n7868) );
  AOI22_X1 U9227 ( .A1(n10390), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n6771), .B2(
        n7864), .ZN(n7862) );
  OAI21_X1 U9228 ( .B1(n7859), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7858), .ZN(
        n10921) );
  MUX2_X1 U9229 ( .A(n11132), .B(P1_REG1_REG_10__SCAN_IN), .S(n10928), .Z(
        n10920) );
  NOR2_X1 U9230 ( .A1(n10921), .A2(n10920), .ZN(n10919) );
  AOI21_X1 U9231 ( .B1(n10928), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10919), .ZN(
        n10827) );
  MUX2_X1 U9232 ( .A(n7860), .B(P1_REG1_REG_11__SCAN_IN), .S(n10826), .Z(
        n10828) );
  NOR2_X1 U9233 ( .A1(n10827), .A2(n10828), .ZN(n10829) );
  AOI21_X1 U9234 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10826), .A(n10829), .ZN(
        n7861) );
  NAND2_X1 U9235 ( .A1(n7862), .A2(n7861), .ZN(n10379) );
  OAI21_X1 U9236 ( .B1(n7862), .B2(n7861), .A(n10379), .ZN(n7866) );
  AND2_X1 U9237 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8986) );
  AOI21_X1 U9238 ( .B1(n10430), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8986), .ZN(
        n7863) );
  OAI21_X1 U9239 ( .B1(n10433), .B2(n7864), .A(n7863), .ZN(n7865) );
  AOI21_X1 U9240 ( .B1(n7866), .B2(n10846), .A(n7865), .ZN(n7867) );
  OAI21_X1 U9241 ( .B1(n7868), .B2(n10922), .A(n7867), .ZN(P1_U3255) );
  OAI21_X1 U9242 ( .B1(n7871), .B2(n7870), .A(n5401), .ZN(n7880) );
  INV_X1 U9243 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9244 ( .A1(n9881), .A2(n7872), .ZN(n7873) );
  NAND2_X1 U9245 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8271) );
  OAI211_X1 U9246 ( .C1(n9873), .C2(n7874), .A(n7873), .B(n8271), .ZN(n7879)
         );
  AOI21_X1 U9247 ( .B1(n7876), .B2(n7875), .A(n5253), .ZN(n7877) );
  NOR2_X1 U9248 ( .A1(n7877), .A2(n10967), .ZN(n7878) );
  AOI211_X1 U9249 ( .C1(n5906), .C2(n7880), .A(n7879), .B(n7878), .ZN(n7886)
         );
  OAI21_X1 U9250 ( .B1(n7883), .B2(n7882), .A(n7881), .ZN(n7884) );
  NAND2_X1 U9251 ( .A1(n7884), .A2(n5272), .ZN(n7885) );
  NAND2_X1 U9252 ( .A1(n7886), .A2(n7885), .ZN(P2_U3190) );
  AOI21_X1 U9253 ( .B1(n10982), .B2(n7888), .A(n7887), .ZN(n7898) );
  XNOR2_X1 U9254 ( .A(n7890), .B(n7889), .ZN(n7896) );
  NOR2_X1 U9255 ( .A1(n8395), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7895) );
  AOI211_X1 U9256 ( .C1(n7893), .C2(n7892), .A(n10939), .B(n7891), .ZN(n7894)
         );
  AOI211_X1 U9257 ( .C1(n5906), .C2(n7896), .A(n7895), .B(n7894), .ZN(n7897)
         );
  OAI21_X1 U9258 ( .B1(n7898), .B2(n10967), .A(n7897), .ZN(n7899) );
  AOI21_X1 U9259 ( .B1(n10959), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n7899), .ZN(
        n7900) );
  OAI21_X1 U9260 ( .B1(n7901), .B2(n5947), .A(n7900), .ZN(P2_U3183) );
  INV_X1 U9261 ( .A(n7922), .ZN(n7931) );
  AND2_X1 U9262 ( .A1(n10338), .A2(n9259), .ZN(n9249) );
  INV_X1 U9263 ( .A(n9249), .ZN(n7902) );
  NAND2_X1 U9264 ( .A1(n7903), .A2(n10987), .ZN(n7904) );
  NAND2_X1 U9265 ( .A1(n9251), .A2(n7904), .ZN(n7932) );
  NAND2_X1 U9266 ( .A1(n7931), .A2(n7932), .ZN(n7930) );
  NAND2_X1 U9267 ( .A1(n7912), .A2(n7936), .ZN(n7905) );
  NAND2_X1 U9268 ( .A1(n7930), .A2(n7905), .ZN(n7907) );
  INV_X1 U9269 ( .A(n7909), .ZN(n7906) );
  OAI21_X1 U9270 ( .B1(n7907), .B2(n7906), .A(n8074), .ZN(n11023) );
  INV_X1 U9271 ( .A(n11023), .ZN(n7920) );
  INV_X1 U9272 ( .A(n7934), .ZN(n7908) );
  NAND2_X1 U9273 ( .A1(n10600), .A2(n7908), .ZN(n9267) );
  OAI21_X1 U9274 ( .B1(n7910), .B2(n7909), .A(n8048), .ZN(n7914) );
  OAI22_X1 U9275 ( .A1(n10228), .A2(n10505), .B1(n7912), .B2(n10507), .ZN(
        n7913) );
  AOI21_X1 U9276 ( .B1(n7914), .B2(n11232), .A(n7913), .ZN(n7915) );
  OAI21_X1 U9277 ( .B1(n7920), .B2(n8947), .A(n7915), .ZN(n11021) );
  NAND2_X1 U9278 ( .A1(n11021), .A2(n10600), .ZN(n7919) );
  AND2_X1 U9279 ( .A1(n9263), .A2(n7936), .ZN(n7926) );
  NAND2_X1 U9280 ( .A1(n7926), .A2(n11020), .ZN(n8053) );
  OAI211_X1 U9281 ( .C1(n7926), .C2(n11020), .A(n11250), .B(n8053), .ZN(n11019) );
  OAI22_X1 U9282 ( .A1(n11253), .A2(n11019), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10580), .ZN(n7917) );
  NOR2_X1 U9283 ( .A1(n10534), .A2(n11020), .ZN(n7916) );
  AOI211_X1 U9284 ( .C1(n11258), .C2(P1_REG2_REG_3__SCAN_IN), .A(n7917), .B(
        n7916), .ZN(n7918) );
  OAI211_X1 U9285 ( .C1(n7920), .C2(n9267), .A(n7919), .B(n7918), .ZN(P1_U3290) );
  XNOR2_X1 U9286 ( .A(n7921), .B(n7922), .ZN(n7923) );
  NAND2_X1 U9287 ( .A1(n7923), .A2(n11232), .ZN(n7925) );
  AOI22_X1 U9288 ( .A1(n11236), .A2(n10337), .B1(n10335), .B2(n11237), .ZN(
        n7924) );
  AND2_X1 U9289 ( .A1(n7925), .A2(n7924), .ZN(n8927) );
  OAI21_X1 U9290 ( .B1(n9263), .B2(n7936), .A(n11250), .ZN(n7927) );
  NOR2_X1 U9291 ( .A1(n7927), .A2(n7926), .ZN(n8924) );
  INV_X1 U9292 ( .A(n10580), .ZN(n11243) );
  AOI22_X1 U9293 ( .A1(n8924), .A2(n7172), .B1(n11243), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U9294 ( .A1(n8927), .A2(n7928), .ZN(n7929) );
  MUX2_X1 U9295 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7929), .S(n10600), .Z(n7938)
         );
  OAI21_X1 U9296 ( .B1(n7932), .B2(n7931), .A(n7930), .ZN(n7933) );
  INV_X1 U9297 ( .A(n7933), .ZN(n8928) );
  NAND2_X1 U9298 ( .A1(n8947), .A2(n7934), .ZN(n7935) );
  OAI22_X1 U9299 ( .A1(n8928), .A2(n11254), .B1(n10534), .B2(n7936), .ZN(n7937) );
  OR2_X1 U9300 ( .A1(n7938), .A2(n7937), .ZN(P1_U3291) );
  INV_X1 U9301 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U9302 ( .A1(n7940), .A2(n9280), .ZN(n7941) );
  NAND2_X1 U9303 ( .A1(n7942), .A2(n7941), .ZN(n8014) );
  XNOR2_X1 U9304 ( .A(n7783), .B(n11048), .ZN(n8015) );
  XNOR2_X1 U9305 ( .A(n8015), .B(n8025), .ZN(n8013) );
  XNOR2_X1 U9306 ( .A(n8014), .B(n8013), .ZN(n7943) );
  NAND2_X1 U9307 ( .A1(n7943), .A2(n9773), .ZN(n7948) );
  NOR2_X1 U9308 ( .A1(n9754), .A2(n9281), .ZN(n7946) );
  OAI21_X1 U9309 ( .B1(n9763), .B2(n9280), .A(n7944), .ZN(n7945) );
  AOI211_X1 U9310 ( .C1(n9282), .C2(n9766), .A(n7946), .B(n7945), .ZN(n7947)
         );
  OAI211_X1 U9311 ( .C1(n11048), .C2(n9784), .A(n7948), .B(n7947), .ZN(
        P2_U3167) );
  INV_X1 U9312 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7963) );
  INV_X1 U9313 ( .A(n7949), .ZN(n7951) );
  NAND3_X1 U9314 ( .A1(n7952), .A2(n7951), .A3(n7950), .ZN(n7953) );
  AOI21_X1 U9315 ( .B1(n7954), .B2(n7953), .A(n10972), .ZN(n7956) );
  NOR2_X1 U9316 ( .A1(n7956), .A2(n7955), .ZN(n7962) );
  AND3_X1 U9317 ( .A1(n7766), .A2(n7958), .A3(n7957), .ZN(n7959) );
  OAI21_X1 U9318 ( .B1(n7960), .B2(n7959), .A(n5874), .ZN(n7961) );
  OAI211_X1 U9319 ( .C1(n7963), .C2(n9873), .A(n7962), .B(n7961), .ZN(n7968)
         );
  AOI211_X1 U9320 ( .C1(n7966), .C2(n7965), .A(n10939), .B(n7964), .ZN(n7967)
         );
  AOI211_X1 U9321 ( .C1(n9881), .C2(n7969), .A(n7968), .B(n7967), .ZN(n7970)
         );
  INV_X1 U9322 ( .A(n7970), .ZN(P2_U3186) );
  INV_X1 U9323 ( .A(n7971), .ZN(n8011) );
  AOI22_X1 U9324 ( .A1(n10407), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n8066), .ZN(n7972) );
  OAI21_X1 U9325 ( .B1(n8011), .B2(n9271), .A(n7972), .ZN(P1_U3339) );
  XNOR2_X1 U9326 ( .A(n7974), .B(n7973), .ZN(n7977) );
  NAND2_X1 U9327 ( .A1(n7726), .A2(n7975), .ZN(n7976) );
  NOR2_X1 U9328 ( .A1(n7976), .A2(n7977), .ZN(n10220) );
  AOI211_X1 U9329 ( .C1(n7977), .C2(n7976), .A(n10292), .B(n10220), .ZN(n7982)
         );
  AOI22_X1 U9330 ( .A1(n9641), .A2(n10335), .B1(n10315), .B2(n10333), .ZN(
        n7980) );
  NOR2_X1 U9331 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7978), .ZN(n10365) );
  AOI21_X1 U9332 ( .B1(n10289), .B2(n8058), .A(n10365), .ZN(n7979) );
  OAI211_X1 U9333 ( .C1(n8055), .C2(n10299), .A(n7980), .B(n7979), .ZN(n7981)
         );
  OR2_X1 U9334 ( .A1(n7982), .A2(n7981), .ZN(P1_U3230) );
  NAND2_X1 U9335 ( .A1(n7984), .A2(n7983), .ZN(n7990) );
  INV_X1 U9336 ( .A(n7985), .ZN(n7987) );
  AOI21_X1 U9337 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  OR2_X1 U9338 ( .A1(n11003), .A2(n6102), .ZN(n8032) );
  MUX2_X1 U9339 ( .A(n7991), .B(n8032), .S(n11015), .Z(n7997) );
  INV_X1 U9340 ( .A(n9588), .ZN(n7993) );
  NOR3_X1 U9341 ( .A1(n7994), .A2(n7993), .A3(n7992), .ZN(n7995) );
  AOI21_X1 U9342 ( .B1(n10028), .B2(P2_REG3_REG_0__SCAN_IN), .A(n7995), .ZN(
        n7996) );
  OAI211_X1 U9343 ( .C1(n8034), .C2(n10030), .A(n7997), .B(n7996), .ZN(
        P2_U3233) );
  INV_X1 U9344 ( .A(n8119), .ZN(n11073) );
  NAND2_X1 U9345 ( .A1(n7999), .A2(n7998), .ZN(n8003) );
  NAND2_X1 U9346 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  XNOR2_X1 U9347 ( .A(n8003), .B(n8002), .ZN(n8004) );
  NAND2_X1 U9348 ( .A1(n8004), .A2(n10308), .ZN(n8009) );
  NAND2_X1 U9349 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10789) );
  INV_X1 U9350 ( .A(n10789), .ZN(n8007) );
  OAI22_X1 U9351 ( .A1(n10313), .A2(n8005), .B1(n10299), .B2(n8082), .ZN(n8006) );
  AOI211_X1 U9352 ( .C1(n10315), .C2(n10331), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI211_X1 U9353 ( .C1(n11073), .C2(n10318), .A(n8009), .B(n8008), .ZN(
        P1_U3239) );
  OAI222_X1 U9354 ( .A1(n8012), .A2(P2_U3151), .B1(n9275), .B2(n8011), .C1(
        n8010), .C2(n10173), .ZN(P2_U3279) );
  NAND2_X1 U9355 ( .A1(n8014), .A2(n8013), .ZN(n8018) );
  INV_X1 U9356 ( .A(n8015), .ZN(n8016) );
  NAND2_X1 U9357 ( .A1(n8016), .A2(n8025), .ZN(n8017) );
  XNOR2_X1 U9358 ( .A(n9373), .B(n11063), .ZN(n8105) );
  XNOR2_X1 U9359 ( .A(n8105), .B(n9803), .ZN(n8020) );
  AOI21_X1 U9360 ( .B1(n8019), .B2(n8020), .A(n9748), .ZN(n8023) );
  INV_X1 U9361 ( .A(n8019), .ZN(n8022) );
  INV_X1 U9362 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U9363 ( .A1(n8023), .A2(n8107), .ZN(n8029) );
  NOR2_X1 U9364 ( .A1(n9754), .A2(n9471), .ZN(n8027) );
  OAI21_X1 U9365 ( .B1(n9763), .B2(n8025), .A(n8024), .ZN(n8026) );
  AOI211_X1 U9366 ( .C1(n8208), .C2(n9766), .A(n8027), .B(n8026), .ZN(n8028)
         );
  OAI211_X1 U9367 ( .C1(n11063), .C2(n9784), .A(n8029), .B(n8028), .ZN(
        P2_U3179) );
  INV_X1 U9368 ( .A(n8030), .ZN(n8063) );
  AOI22_X1 U9369 ( .A1(n10877), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n8066), .ZN(n8031) );
  OAI21_X1 U9370 ( .B1(n8063), .B2(n9271), .A(n8031), .ZN(P1_U3338) );
  INV_X1 U9371 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8036) );
  OAI21_X1 U9372 ( .B1(n11159), .B2(n10041), .A(n9588), .ZN(n8033) );
  OAI211_X1 U9373 ( .C1(n11179), .C2(n8034), .A(n8033), .B(n8032), .ZN(n8037)
         );
  NAND2_X1 U9374 ( .A1(n8037), .A2(n11191), .ZN(n8035) );
  OAI21_X1 U9375 ( .B1(n11191), .B2(n8036), .A(n8035), .ZN(P2_U3390) );
  NAND2_X1 U9376 ( .A1(n8037), .A2(n11187), .ZN(n8038) );
  OAI21_X1 U9377 ( .B1(n11187), .B2(n5816), .A(n8038), .ZN(P2_U3459) );
  XOR2_X1 U9378 ( .A(n8041), .B(n8040), .Z(n8042) );
  XNOR2_X1 U9379 ( .A(n8039), .B(n8042), .ZN(n8046) );
  NAND2_X1 U9380 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10801) );
  OAI21_X1 U9381 ( .B1(n10300), .B2(n9388), .A(n10801), .ZN(n8044) );
  OAI22_X1 U9382 ( .A1(n10313), .A2(n8099), .B1(n10299), .B2(n8346), .ZN(n8043) );
  AOI211_X1 U9383 ( .C1(n8348), .C2(n10289), .A(n8044), .B(n8043), .ZN(n8045)
         );
  OAI21_X1 U9384 ( .B1(n8046), .B2(n10292), .A(n8045), .ZN(P1_U3213) );
  NAND2_X1 U9385 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  XOR2_X1 U9386 ( .A(n8071), .B(n8049), .Z(n8050) );
  AOI222_X1 U9387 ( .A1(n11232), .A2(n8050), .B1(n10333), .B2(n11237), .C1(
        n10335), .C2(n11236), .ZN(n11042) );
  NAND2_X1 U9388 ( .A1(n8051), .A2(n11020), .ZN(n8068) );
  NAND2_X1 U9389 ( .A1(n8074), .A2(n8068), .ZN(n8052) );
  XNOR2_X1 U9390 ( .A(n8052), .B(n8071), .ZN(n11045) );
  INV_X1 U9391 ( .A(n8053), .ZN(n8054) );
  OAI211_X1 U9392 ( .C1(n8054), .C2(n11043), .A(n11250), .B(n8089), .ZN(n11041) );
  OAI22_X1 U9393 ( .A1(n10600), .A2(n8056), .B1(n8055), .B2(n10580), .ZN(n8057) );
  AOI21_X1 U9394 ( .B1(n11245), .B2(n8058), .A(n8057), .ZN(n8059) );
  OAI21_X1 U9395 ( .B1(n11253), .B2(n11041), .A(n8059), .ZN(n8060) );
  AOI21_X1 U9396 ( .B1(n11045), .B2(n11218), .A(n8060), .ZN(n8061) );
  OAI21_X1 U9397 ( .B1(n11042), .B2(n11244), .A(n8061), .ZN(P1_U3289) );
  OAI222_X1 U9398 ( .A1(P2_U3151), .A2(n8064), .B1(n9275), .B2(n8063), .C1(
        n8062), .C2(n10173), .ZN(P2_U3278) );
  INV_X1 U9399 ( .A(n8065), .ZN(n8104) );
  AOI22_X1 U9400 ( .A1(n10898), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n8066), .ZN(n8067) );
  OAI21_X1 U9401 ( .B1(n8104), .B2(n9271), .A(n8067), .ZN(P1_U3337) );
  NAND2_X1 U9402 ( .A1(n10228), .A2(n11043), .ZN(n8069) );
  AND2_X1 U9403 ( .A1(n8068), .A2(n8069), .ZN(n8073) );
  INV_X1 U9404 ( .A(n8069), .ZN(n8070) );
  NAND2_X1 U9405 ( .A1(n8088), .A2(n8096), .ZN(n8076) );
  OR2_X1 U9406 ( .A1(n10333), .A2(n10230), .ZN(n8075) );
  NAND2_X1 U9407 ( .A1(n8076), .A2(n8075), .ZN(n8118) );
  XNOR2_X1 U9408 ( .A(n8118), .B(n8116), .ZN(n11070) );
  XNOR2_X1 U9409 ( .A(n8077), .B(n8116), .ZN(n8078) );
  AOI222_X1 U9410 ( .A1(n11232), .A2(n8078), .B1(n10331), .B2(n11237), .C1(
        n10333), .C2(n11236), .ZN(n11072) );
  INV_X1 U9411 ( .A(n11072), .ZN(n8086) );
  OR2_X1 U9412 ( .A1(n8089), .A2(n10230), .ZN(n8090) );
  INV_X1 U9413 ( .A(n8344), .ZN(n8080) );
  AOI21_X1 U9414 ( .B1(n8090), .B2(n8119), .A(n10609), .ZN(n8079) );
  NAND2_X1 U9415 ( .A1(n8080), .A2(n8079), .ZN(n11071) );
  NAND2_X1 U9416 ( .A1(n11258), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8081) );
  OAI21_X1 U9417 ( .B1(n10580), .B2(n8082), .A(n8081), .ZN(n8083) );
  AOI21_X1 U9418 ( .B1(n11245), .B2(n8119), .A(n8083), .ZN(n8084) );
  OAI21_X1 U9419 ( .B1(n11071), .B2(n11253), .A(n8084), .ZN(n8085) );
  AOI21_X1 U9420 ( .B1(n8086), .B2(n10600), .A(n8085), .ZN(n8087) );
  OAI21_X1 U9421 ( .B1(n11070), .B2(n11254), .A(n8087), .ZN(P1_U3287) );
  XNOR2_X1 U9422 ( .A(n8088), .B(n8096), .ZN(n11059) );
  INV_X1 U9423 ( .A(n8089), .ZN(n8091) );
  INV_X1 U9424 ( .A(n10230), .ZN(n11056) );
  OAI211_X1 U9425 ( .C1(n8091), .C2(n11056), .A(n11250), .B(n8090), .ZN(n11055) );
  INV_X1 U9426 ( .A(n10227), .ZN(n8092) );
  AOI22_X1 U9427 ( .A1(n11245), .A2(n10230), .B1(n11243), .B2(n8092), .ZN(
        n8093) );
  OAI21_X1 U9428 ( .B1(n11253), .B2(n11055), .A(n8093), .ZN(n8101) );
  INV_X1 U9429 ( .A(n8094), .ZN(n8095) );
  AOI21_X1 U9430 ( .B1(n8097), .B2(n8096), .A(n8095), .ZN(n8098) );
  OAI222_X1 U9431 ( .A1(n10505), .A2(n8099), .B1(n10507), .B2(n10228), .C1(
        n10503), .C2(n8098), .ZN(n11057) );
  MUX2_X1 U9432 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11057), .S(n10600), .Z(n8100) );
  AOI211_X1 U9433 ( .C1(n11218), .C2(n11059), .A(n8101), .B(n8100), .ZN(n8102)
         );
  INV_X1 U9434 ( .A(n8102), .ZN(P1_U3288) );
  INV_X1 U9435 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8103) );
  OAI222_X1 U9436 ( .A1(P2_U3151), .A2(n10956), .B1(n10175), .B2(n8104), .C1(
        n8103), .C2(n10173), .ZN(P2_U3277) );
  INV_X1 U9437 ( .A(n9472), .ZN(n11087) );
  NAND2_X1 U9438 ( .A1(n8105), .A2(n9803), .ZN(n8106) );
  XNOR2_X1 U9439 ( .A(n9472), .B(n9373), .ZN(n8266) );
  XNOR2_X1 U9440 ( .A(n8266), .B(n9802), .ZN(n8108) );
  OAI21_X1 U9441 ( .B1(n8109), .B2(n8108), .A(n8268), .ZN(n8110) );
  NAND2_X1 U9442 ( .A1(n8110), .A2(n9773), .ZN(n8115) );
  NOR2_X1 U9443 ( .A1(n9754), .A2(n8304), .ZN(n8113) );
  OAI21_X1 U9444 ( .B1(n9763), .B2(n9281), .A(n8111), .ZN(n8112) );
  AOI211_X1 U9445 ( .C1(n8219), .C2(n9766), .A(n8113), .B(n8112), .ZN(n8114)
         );
  OAI211_X1 U9446 ( .C1(n11087), .C2(n9784), .A(n8115), .B(n8114), .ZN(
        P2_U3153) );
  INV_X1 U9447 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U9448 ( .A1(n8118), .A2(n8117), .ZN(n8121) );
  OR2_X1 U9449 ( .A1(n8119), .A2(n10332), .ZN(n8120) );
  NAND2_X1 U9450 ( .A1(n8121), .A2(n8120), .ZN(n8342) );
  INV_X1 U9451 ( .A(n8352), .ZN(n8341) );
  NAND2_X1 U9452 ( .A1(n8342), .A2(n8341), .ZN(n8123) );
  OR2_X1 U9453 ( .A1(n8348), .A2(n10331), .ZN(n8122) );
  NAND2_X1 U9454 ( .A1(n8123), .A2(n8122), .ZN(n8176) );
  NAND2_X1 U9455 ( .A1(n8176), .A2(n8124), .ZN(n8126) );
  OR2_X1 U9456 ( .A1(n8321), .A2(n10330), .ZN(n8125) );
  NAND2_X1 U9457 ( .A1(n8126), .A2(n8125), .ZN(n8281) );
  NAND2_X1 U9458 ( .A1(n8281), .A2(n8284), .ZN(n8128) );
  OR2_X1 U9459 ( .A1(n11112), .A2(n10329), .ZN(n8127) );
  NAND2_X1 U9460 ( .A1(n8128), .A2(n8127), .ZN(n8331) );
  XNOR2_X1 U9461 ( .A(n8331), .B(n8330), .ZN(n11131) );
  INV_X1 U9462 ( .A(n11131), .ZN(n8140) );
  NAND2_X1 U9463 ( .A1(n8131), .A2(n11232), .ZN(n8133) );
  AOI22_X1 U9464 ( .A1(n11237), .A2(n10327), .B1(n10329), .B2(n11236), .ZN(
        n8132) );
  NAND2_X1 U9465 ( .A1(n8133), .A2(n8132), .ZN(n11130) );
  INV_X1 U9466 ( .A(n8473), .ZN(n11128) );
  INV_X1 U9467 ( .A(n8348), .ZN(n11082) );
  NAND2_X1 U9468 ( .A1(n8344), .A2(n11082), .ZN(n8343) );
  OR2_X1 U9469 ( .A1(n8343), .A2(n8321), .ZN(n8290) );
  AND2_X1 U9470 ( .A1(n8293), .A2(n11128), .ZN(n8334) );
  INV_X1 U9471 ( .A(n8334), .ZN(n8134) );
  OAI211_X1 U9472 ( .C1(n11128), .C2(n8293), .A(n8134), .B(n11250), .ZN(n11127) );
  OAI22_X1 U9473 ( .A1(n10600), .A2(n8135), .B1(n8469), .B2(n10580), .ZN(n8136) );
  AOI21_X1 U9474 ( .B1(n8473), .B2(n11245), .A(n8136), .ZN(n8137) );
  OAI21_X1 U9475 ( .B1(n11127), .B2(n11253), .A(n8137), .ZN(n8138) );
  AOI21_X1 U9476 ( .B1(n11130), .B2(n10600), .A(n8138), .ZN(n8139) );
  OAI21_X1 U9477 ( .B1(n8140), .B2(n11254), .A(n8139), .ZN(P1_U3283) );
  AOI21_X1 U9478 ( .B1(n11124), .B2(n8142), .A(n8141), .ZN(n8155) );
  AOI21_X1 U9479 ( .B1(n8144), .B2(n8200), .A(n8143), .ZN(n8151) );
  NAND2_X1 U9480 ( .A1(n10959), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n8150) );
  OAI21_X1 U9481 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8148) );
  NOR2_X1 U9482 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8585), .ZN(n8305) );
  AOI21_X1 U9483 ( .B1(n8148), .B2(n5272), .A(n8305), .ZN(n8149) );
  OAI211_X1 U9484 ( .C1(n8151), .C2(n10972), .A(n8150), .B(n8149), .ZN(n8152)
         );
  AOI21_X1 U9485 ( .B1(n8153), .B2(n9881), .A(n8152), .ZN(n8154) );
  OAI21_X1 U9486 ( .B1(n8155), .B2(n10967), .A(n8154), .ZN(P2_U3191) );
  NOR2_X1 U9487 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n8156) );
  AOI21_X1 U9488 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n8156), .ZN(n10760) );
  INV_X1 U9489 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10889) );
  INV_X1 U9490 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U9491 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10889), .B2(n9872), .ZN(n10757) );
  NOR2_X1 U9492 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8157) );
  AOI21_X1 U9493 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8157), .ZN(n10754) );
  NOR2_X1 U9494 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8158) );
  AOI21_X1 U9495 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8158), .ZN(n10751) );
  NOR2_X1 U9496 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8159) );
  AOI21_X1 U9497 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8159), .ZN(n10748) );
  NOR2_X1 U9498 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8160) );
  AOI21_X1 U9499 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8160), .ZN(n10745) );
  NOR2_X1 U9500 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8161) );
  AOI21_X1 U9501 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8161), .ZN(n10742) );
  NOR2_X1 U9502 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8162) );
  AOI21_X1 U9503 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8162), .ZN(n10739) );
  NOR2_X1 U9504 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8163) );
  AOI21_X1 U9505 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8163), .ZN(n10736) );
  NOR2_X1 U9506 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8164) );
  AOI21_X1 U9507 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8164), .ZN(n10733) );
  NOR2_X1 U9508 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8165) );
  AOI21_X1 U9509 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n8165), .ZN(n10730) );
  NOR2_X1 U9510 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8166) );
  AOI21_X1 U9511 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8166), .ZN(n10727) );
  NOR2_X1 U9512 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8167) );
  AOI21_X1 U9513 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n8167), .ZN(n10724) );
  NOR2_X1 U9514 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8168) );
  AOI21_X1 U9515 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8168), .ZN(n10721) );
  NAND2_X1 U9516 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10707) );
  INV_X1 U9517 ( .A(n10707), .ZN(n8169) );
  INV_X1 U9518 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U9519 ( .A1(n10708), .A2(n10707), .ZN(n10706) );
  AOI22_X1 U9520 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n8169), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10706), .ZN(n10712) );
  NAND2_X1 U9521 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8170) );
  OAI21_X1 U9522 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n8170), .ZN(n10711) );
  NOR2_X1 U9523 ( .A1(n10712), .A2(n10711), .ZN(n10710) );
  AOI21_X1 U9524 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10710), .ZN(n10715) );
  NAND2_X1 U9525 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8171) );
  OAI21_X1 U9526 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n8171), .ZN(n10714) );
  NOR2_X1 U9527 ( .A1(n10715), .A2(n10714), .ZN(n10713) );
  AOI21_X1 U9528 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10713), .ZN(n10718) );
  NOR2_X1 U9529 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8172) );
  AOI21_X1 U9530 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n8172), .ZN(n10717) );
  NAND2_X1 U9531 ( .A1(n10718), .A2(n10717), .ZN(n10716) );
  OAI21_X1 U9532 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10716), .ZN(n10720) );
  NAND2_X1 U9533 ( .A1(n10721), .A2(n10720), .ZN(n10719) );
  OAI21_X1 U9534 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10719), .ZN(n10723) );
  NAND2_X1 U9535 ( .A1(n10724), .A2(n10723), .ZN(n10722) );
  OAI21_X1 U9536 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10722), .ZN(n10726) );
  NAND2_X1 U9537 ( .A1(n10727), .A2(n10726), .ZN(n10725) );
  OAI21_X1 U9538 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10725), .ZN(n10729) );
  NAND2_X1 U9539 ( .A1(n10730), .A2(n10729), .ZN(n10728) );
  OAI21_X1 U9540 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10728), .ZN(n10732) );
  NAND2_X1 U9541 ( .A1(n10733), .A2(n10732), .ZN(n10731) );
  OAI21_X1 U9542 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10731), .ZN(n10735) );
  NAND2_X1 U9543 ( .A1(n10736), .A2(n10735), .ZN(n10734) );
  OAI21_X1 U9544 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10734), .ZN(n10738) );
  NAND2_X1 U9545 ( .A1(n10739), .A2(n10738), .ZN(n10737) );
  OAI21_X1 U9546 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10737), .ZN(n10741) );
  NAND2_X1 U9547 ( .A1(n10742), .A2(n10741), .ZN(n10740) );
  OAI21_X1 U9548 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10740), .ZN(n10744) );
  NAND2_X1 U9549 ( .A1(n10745), .A2(n10744), .ZN(n10743) );
  OAI21_X1 U9550 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10743), .ZN(n10747) );
  NAND2_X1 U9551 ( .A1(n10748), .A2(n10747), .ZN(n10746) );
  OAI21_X1 U9552 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10746), .ZN(n10750) );
  NAND2_X1 U9553 ( .A1(n10751), .A2(n10750), .ZN(n10749) );
  OAI21_X1 U9554 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10749), .ZN(n10753) );
  NAND2_X1 U9555 ( .A1(n10754), .A2(n10753), .ZN(n10752) );
  OAI21_X1 U9556 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10752), .ZN(n10756) );
  NAND2_X1 U9557 ( .A1(n10757), .A2(n10756), .ZN(n10755) );
  OAI21_X1 U9558 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10755), .ZN(n10759) );
  NAND2_X1 U9559 ( .A1(n10760), .A2(n10759), .ZN(n10758) );
  OAI21_X1 U9560 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10758), .ZN(n8175) );
  XNOR2_X1 U9561 ( .A(n8173), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8174) );
  XNOR2_X1 U9562 ( .A(n8175), .B(n8174), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9563 ( .A(n8176), .B(n8181), .ZN(n11094) );
  AOI22_X1 U9564 ( .A1(n11236), .A2(n10331), .B1(n10329), .B2(n11237), .ZN(
        n8184) );
  AND2_X1 U9565 ( .A1(n8178), .A2(n8177), .ZN(n8351) );
  NAND2_X1 U9566 ( .A1(n8351), .A2(n8352), .ZN(n8350) );
  NAND2_X1 U9567 ( .A1(n8350), .A2(n8179), .ZN(n8180) );
  NAND2_X1 U9568 ( .A1(n8180), .A2(n8181), .ZN(n8283) );
  OAI21_X1 U9569 ( .B1(n8181), .B2(n8180), .A(n8283), .ZN(n8182) );
  NAND2_X1 U9570 ( .A1(n8182), .A2(n11232), .ZN(n8183) );
  OAI211_X1 U9571 ( .C1(n11094), .C2(n8947), .A(n8184), .B(n8183), .ZN(n11097)
         );
  NAND2_X1 U9572 ( .A1(n11097), .A2(n10600), .ZN(n8190) );
  OAI22_X1 U9573 ( .A1(n10600), .A2(n8185), .B1(n8317), .B2(n10580), .ZN(n8188) );
  INV_X1 U9574 ( .A(n8343), .ZN(n8186) );
  INV_X1 U9575 ( .A(n8321), .ZN(n11096) );
  OAI211_X1 U9576 ( .C1(n8186), .C2(n11096), .A(n11250), .B(n8290), .ZN(n11095) );
  NOR2_X1 U9577 ( .A1(n11095), .A2(n11253), .ZN(n8187) );
  AOI211_X1 U9578 ( .C1(n11245), .C2(n8321), .A(n8188), .B(n8187), .ZN(n8189)
         );
  OAI211_X1 U9579 ( .C1(n11094), .C2(n9267), .A(n8190), .B(n8189), .ZN(
        P1_U3285) );
  NAND2_X1 U9580 ( .A1(n8191), .A2(n7485), .ZN(n8430) );
  NAND2_X1 U9581 ( .A1(n9660), .A2(n8430), .ZN(n11014) );
  OAI21_X1 U9582 ( .B1(n8193), .B2(n9598), .A(n8192), .ZN(n11120) );
  NAND3_X1 U9583 ( .A1(n8194), .A2(n9598), .A3(n8195), .ZN(n8196) );
  AND2_X1 U9584 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  OAI222_X1 U9585 ( .A1(n11003), .A2(n8410), .B1(n11001), .B2(n8304), .C1(
        n11000), .C2(n8198), .ZN(n11121) );
  NAND2_X1 U9586 ( .A1(n11121), .A2(n11015), .ZN(n8203) );
  INV_X1 U9587 ( .A(n8309), .ZN(n8199) );
  OAI22_X1 U9588 ( .A1(n11015), .A2(n8200), .B1(n8199), .B2(n11010), .ZN(n8201) );
  AOI21_X1 U9589 ( .B1(n10015), .B2(n11123), .A(n8201), .ZN(n8202) );
  OAI211_X1 U9590 ( .C1(n10012), .C2(n11120), .A(n8203), .B(n8202), .ZN(
        P2_U3224) );
  INV_X1 U9591 ( .A(n8204), .ZN(n9594) );
  XNOR2_X1 U9592 ( .A(n8205), .B(n9594), .ZN(n11064) );
  XNOR2_X1 U9593 ( .A(n8206), .B(n9594), .ZN(n8207) );
  AOI222_X1 U9594 ( .A1(n10041), .A2(n8207), .B1(n9802), .B2(n10003), .C1(
        n9804), .C2(n10001), .ZN(n11062) );
  MUX2_X1 U9595 ( .A(n5884), .B(n11062), .S(n11015), .Z(n8211) );
  INV_X1 U9596 ( .A(n11063), .ZN(n8209) );
  AOI22_X1 U9597 ( .A1(n10015), .A2(n8209), .B1(n10028), .B2(n8208), .ZN(n8210) );
  OAI211_X1 U9598 ( .C1(n10012), .C2(n11064), .A(n8211), .B(n8210), .ZN(
        P2_U3227) );
  OAI21_X1 U9599 ( .B1(n8213), .B2(n8217), .A(n8212), .ZN(n11088) );
  INV_X1 U9600 ( .A(n8214), .ZN(n8215) );
  AOI21_X1 U9601 ( .B1(n8217), .B2(n8216), .A(n8215), .ZN(n8218) );
  OAI222_X1 U9602 ( .A1(n11003), .A2(n8304), .B1(n11001), .B2(n9281), .C1(
        n11000), .C2(n8218), .ZN(n11090) );
  NAND2_X1 U9603 ( .A1(n11090), .A2(n11015), .ZN(n8224) );
  INV_X1 U9604 ( .A(n8219), .ZN(n8220) );
  OAI22_X1 U9605 ( .A1(n11015), .A2(n8221), .B1(n8220), .B2(n11010), .ZN(n8222) );
  AOI21_X1 U9606 ( .B1(n10015), .B2(n9472), .A(n8222), .ZN(n8223) );
  OAI211_X1 U9607 ( .C1(n10012), .C2(n11088), .A(n8224), .B(n8223), .ZN(
        P2_U3226) );
  XNOR2_X1 U9608 ( .A(n8225), .B(n9597), .ZN(n11102) );
  INV_X1 U9609 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8229) );
  NAND3_X1 U9610 ( .A1(n8214), .A2(n9597), .A3(n8226), .ZN(n8227) );
  NAND2_X1 U9611 ( .A1(n8194), .A2(n8227), .ZN(n8228) );
  AOI222_X1 U9612 ( .A1(n10041), .A2(n8228), .B1(n9800), .B2(n10003), .C1(
        n9802), .C2(n10001), .ZN(n11103) );
  MUX2_X1 U9613 ( .A(n8229), .B(n11103), .S(n11015), .Z(n8232) );
  AOI22_X1 U9614 ( .A1(n10015), .A2(n8230), .B1(n10028), .B2(n8274), .ZN(n8231) );
  OAI211_X1 U9615 ( .C1(n11102), .C2(n10012), .A(n8232), .B(n8231), .ZN(
        P2_U3225) );
  INV_X1 U9616 ( .A(n9591), .ZN(n8236) );
  NAND3_X1 U9617 ( .A1(n8233), .A2(n9439), .A3(n8236), .ZN(n8234) );
  AND2_X1 U9618 ( .A1(n8235), .A2(n8234), .ZN(n11028) );
  XNOR2_X1 U9619 ( .A(n8237), .B(n8236), .ZN(n8238) );
  AOI222_X1 U9620 ( .A1(n10041), .A2(n8238), .B1(n9805), .B2(n10003), .C1(
        n9807), .C2(n10001), .ZN(n11026) );
  MUX2_X1 U9621 ( .A(n7770), .B(n11026), .S(n11015), .Z(n8241) );
  INV_X1 U9622 ( .A(n11027), .ZN(n8239) );
  AOI22_X1 U9623 ( .A1(n10015), .A2(n8239), .B1(n10028), .B2(n8763), .ZN(n8240) );
  OAI211_X1 U9624 ( .C1(n11028), .C2(n10012), .A(n8241), .B(n8240), .ZN(
        P2_U3230) );
  XNOR2_X1 U9625 ( .A(n9805), .B(n8247), .ZN(n9590) );
  XOR2_X1 U9626 ( .A(n8242), .B(n9590), .Z(n11036) );
  XOR2_X1 U9627 ( .A(n8243), .B(n9590), .Z(n8244) );
  AOI222_X1 U9628 ( .A1(n10041), .A2(n8244), .B1(n9804), .B2(n10003), .C1(
        n9806), .C2(n10001), .ZN(n11034) );
  MUX2_X1 U9629 ( .A(n8245), .B(n11034), .S(n11015), .Z(n8249) );
  AOI22_X1 U9630 ( .A1(n10015), .A2(n8247), .B1(n10028), .B2(n8246), .ZN(n8248) );
  OAI211_X1 U9631 ( .C1(n11036), .C2(n10012), .A(n8249), .B(n8248), .ZN(
        P2_U3229) );
  INV_X1 U9632 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U9633 ( .A1(n8257), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9634 ( .A1(n8250), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8251) );
  OAI211_X1 U9635 ( .C1(n8253), .C2(n8260), .A(n8252), .B(n8251), .ZN(n8254)
         );
  INV_X1 U9636 ( .A(n8254), .ZN(n8255) );
  NAND2_X1 U9637 ( .A1(n10961), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8256) );
  OAI21_X1 U9638 ( .B1(n9887), .B2(n10961), .A(n8256), .ZN(P2_U3522) );
  INV_X1 U9639 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U9640 ( .A1(n8250), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U9641 ( .A1(n8257), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8258) );
  OAI211_X1 U9642 ( .C1(n8261), .C2(n8260), .A(n8259), .B(n8258), .ZN(n8262)
         );
  INV_X1 U9643 ( .A(n8262), .ZN(n8263) );
  NAND2_X1 U9644 ( .A1(n10961), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8265) );
  OAI21_X1 U9645 ( .B1(n9663), .B2(n10961), .A(n8265), .ZN(P2_U3521) );
  NAND2_X1 U9646 ( .A1(n8266), .A2(n9471), .ZN(n8267) );
  XNOR2_X1 U9647 ( .A(n11104), .B(n9355), .ZN(n8302) );
  XNOR2_X1 U9648 ( .A(n8302), .B(n9801), .ZN(n8269) );
  XNOR2_X1 U9649 ( .A(n8303), .B(n8269), .ZN(n8270) );
  NAND2_X1 U9650 ( .A1(n8270), .A2(n9773), .ZN(n8276) );
  NOR2_X1 U9651 ( .A1(n9754), .A2(n8425), .ZN(n8273) );
  OAI21_X1 U9652 ( .B1(n9763), .B2(n9471), .A(n8271), .ZN(n8272) );
  AOI211_X1 U9653 ( .C1(n8274), .C2(n9766), .A(n8273), .B(n8272), .ZN(n8275)
         );
  OAI211_X1 U9654 ( .C1(n11104), .C2(n9784), .A(n8276), .B(n8275), .ZN(
        P2_U3161) );
  NAND2_X1 U9655 ( .A1(n10961), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8277) );
  OAI21_X1 U9656 ( .B1(n9419), .B2(n10961), .A(n8277), .ZN(P2_U3520) );
  INV_X1 U9657 ( .A(n8278), .ZN(n8279) );
  OAI222_X1 U9658 ( .A1(n5135), .A2(P2_U3151), .B1(n10175), .B2(n8279), .C1(
        n10173), .C2(n6045), .ZN(P2_U3276) );
  OAI222_X1 U9659 ( .A1(n10696), .A2(n8280), .B1(n9271), .B2(n8279), .C1(
        P1_U3086), .C2(n7172), .ZN(P1_U3336) );
  XNOR2_X1 U9660 ( .A(n8281), .B(n8284), .ZN(n11110) );
  INV_X1 U9661 ( .A(n11110), .ZN(n8299) );
  NAND2_X1 U9662 ( .A1(n8283), .A2(n8282), .ZN(n8286) );
  INV_X1 U9663 ( .A(n8284), .ZN(n8285) );
  XNOR2_X1 U9664 ( .A(n8286), .B(n8285), .ZN(n8287) );
  NAND2_X1 U9665 ( .A1(n8287), .A2(n11232), .ZN(n8289) );
  NAND2_X1 U9666 ( .A1(n10330), .A2(n11236), .ZN(n8288) );
  NAND2_X1 U9667 ( .A1(n8289), .A2(n8288), .ZN(n11117) );
  NAND2_X1 U9668 ( .A1(n11117), .A2(n10600), .ZN(n8298) );
  NAND2_X1 U9669 ( .A1(n8290), .A2(n11112), .ZN(n8291) );
  NAND2_X1 U9670 ( .A1(n8291), .A2(n11250), .ZN(n8292) );
  OAI22_X1 U9671 ( .A1(n8293), .A2(n8292), .B1(n8498), .B2(n10505), .ZN(n11114) );
  INV_X1 U9672 ( .A(n11112), .ZN(n9393) );
  NOR2_X1 U9673 ( .A1(n9393), .A2(n10534), .ZN(n8296) );
  OAI22_X1 U9674 ( .A1(n10600), .A2(n8294), .B1(n9387), .B2(n10580), .ZN(n8295) );
  AOI211_X1 U9675 ( .C1(n11114), .C2(n10560), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI211_X1 U9676 ( .C1(n8299), .C2(n11254), .A(n8298), .B(n8297), .ZN(
        P1_U3284) );
  INV_X1 U9677 ( .A(n8300), .ZN(n8326) );
  OAI222_X1 U9678 ( .A1(n9271), .A2(n8326), .B1(n7197), .B2(P1_U3086), .C1(
        n8301), .C2(n10696), .ZN(P1_U3334) );
  XNOR2_X1 U9679 ( .A(n11123), .B(n9373), .ZN(n8991) );
  XNOR2_X1 U9680 ( .A(n8991), .B(n9800), .ZN(n8989) );
  XNOR2_X1 U9681 ( .A(n8990), .B(n8989), .ZN(n8312) );
  OR2_X1 U9682 ( .A1(n9763), .A2(n8304), .ZN(n8307) );
  INV_X1 U9683 ( .A(n8305), .ZN(n8306) );
  OAI211_X1 U9684 ( .C1(n9754), .C2(n8410), .A(n8307), .B(n8306), .ZN(n8308)
         );
  AOI21_X1 U9685 ( .B1(n8309), .B2(n9766), .A(n8308), .ZN(n8311) );
  NAND2_X1 U9686 ( .A1(n11123), .A2(n9731), .ZN(n8310) );
  OAI211_X1 U9687 ( .C1(n8312), .C2(n9748), .A(n8311), .B(n8310), .ZN(P2_U3171) );
  INV_X1 U9688 ( .A(n8313), .ZN(n8316) );
  NAND2_X1 U9689 ( .A1(n5249), .A2(n8314), .ZN(n9380) );
  OAI21_X1 U9690 ( .B1(n5249), .B2(n8314), .A(n9380), .ZN(n8315) );
  NOR2_X1 U9691 ( .A1(n8315), .A2(n8316), .ZN(n9383) );
  AOI21_X1 U9692 ( .B1(n8316), .B2(n8315), .A(n9383), .ZN(n8324) );
  NAND2_X1 U9693 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10818) );
  INV_X1 U9694 ( .A(n10818), .ZN(n8320) );
  OAI22_X1 U9695 ( .A1(n10313), .A2(n8318), .B1(n10299), .B2(n8317), .ZN(n8319) );
  AOI211_X1 U9696 ( .C1(n10315), .C2(n10329), .A(n8320), .B(n8319), .ZN(n8323)
         );
  NAND2_X1 U9697 ( .A1(n8321), .A2(n10289), .ZN(n8322) );
  OAI211_X1 U9698 ( .C1(n8324), .C2(n10292), .A(n8323), .B(n8322), .ZN(
        P1_U3221) );
  OAI222_X1 U9699 ( .A1(P2_U3151), .A2(n7483), .B1(n10175), .B2(n8326), .C1(
        n8325), .C2(n10173), .ZN(P2_U3274) );
  XOR2_X1 U9700 ( .A(n8455), .B(n8328), .Z(n8329) );
  AOI222_X1 U9701 ( .A1(n11232), .A2(n8329), .B1(n10328), .B2(n11236), .C1(
        n10326), .C2(n11237), .ZN(n11151) );
  NAND2_X1 U9702 ( .A1(n8331), .A2(n8330), .ZN(n8333) );
  OR2_X1 U9703 ( .A1(n8473), .A2(n10328), .ZN(n8332) );
  NAND2_X1 U9704 ( .A1(n8333), .A2(n8332), .ZN(n8456) );
  XNOR2_X1 U9705 ( .A(n8456), .B(n8455), .ZN(n11154) );
  INV_X1 U9706 ( .A(n8457), .ZN(n11152) );
  OAI21_X1 U9707 ( .B1(n8334), .B2(n11152), .A(n11250), .ZN(n8335) );
  OR2_X1 U9708 ( .A1(n8459), .A2(n8335), .ZN(n11150) );
  NAND2_X1 U9709 ( .A1(n11258), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8336) );
  OAI21_X1 U9710 ( .B1(n10580), .B2(n8497), .A(n8336), .ZN(n8337) );
  AOI21_X1 U9711 ( .B1(n8457), .B2(n11245), .A(n8337), .ZN(n8338) );
  OAI21_X1 U9712 ( .B1(n11150), .B2(n11253), .A(n8338), .ZN(n8339) );
  AOI21_X1 U9713 ( .B1(n11154), .B2(n11218), .A(n8339), .ZN(n8340) );
  OAI21_X1 U9714 ( .B1(n11151), .B2(n11244), .A(n8340), .ZN(P1_U3282) );
  XNOR2_X1 U9715 ( .A(n8342), .B(n8341), .ZN(n11084) );
  OAI211_X1 U9716 ( .C1(n8344), .C2(n11082), .A(n11250), .B(n8343), .ZN(n11080) );
  NAND2_X1 U9717 ( .A1(n11258), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8345) );
  OAI21_X1 U9718 ( .B1(n10580), .B2(n8346), .A(n8345), .ZN(n8347) );
  AOI21_X1 U9719 ( .B1(n11245), .B2(n8348), .A(n8347), .ZN(n8349) );
  OAI21_X1 U9720 ( .B1(n11080), .B2(n11253), .A(n8349), .ZN(n8355) );
  OAI21_X1 U9721 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8353) );
  AOI222_X1 U9722 ( .A1(n11232), .A2(n8353), .B1(n10330), .B2(n11237), .C1(
        n10332), .C2(n11236), .ZN(n11081) );
  NOR2_X1 U9723 ( .A1(n11081), .A2(n11244), .ZN(n8354) );
  AOI211_X1 U9724 ( .C1(n11218), .C2(n11084), .A(n8355), .B(n8354), .ZN(n8356)
         );
  INV_X1 U9725 ( .A(n8356), .ZN(P1_U3286) );
  NAND2_X1 U9726 ( .A1(n8384), .A2(n10693), .ZN(n8358) );
  OAI211_X1 U9727 ( .C1(n8823), .C2(n10696), .A(n8358), .B(n8357), .ZN(
        P1_U3335) );
  AOI21_X1 U9728 ( .B1(n8361), .B2(n8360), .A(n8359), .ZN(n8377) );
  INV_X1 U9729 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8368) );
  OAI21_X1 U9730 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(n8366) );
  INV_X1 U9731 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8365) );
  NOR2_X1 U9732 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8365), .ZN(n8999) );
  AOI21_X1 U9733 ( .B1(n8366), .B2(n5272), .A(n8999), .ZN(n8367) );
  OAI21_X1 U9734 ( .B1(n9873), .B2(n8368), .A(n8367), .ZN(n8374) );
  AOI21_X1 U9735 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8372) );
  NOR2_X1 U9736 ( .A1(n8372), .A2(n10972), .ZN(n8373) );
  AOI211_X1 U9737 ( .C1(n9881), .C2(n8375), .A(n8374), .B(n8373), .ZN(n8376)
         );
  OAI21_X1 U9738 ( .B1(n8377), .B2(n10967), .A(n8376), .ZN(P2_U3192) );
  INV_X1 U9739 ( .A(n8378), .ZN(n8382) );
  OAI222_X1 U9740 ( .A1(n8380), .A2(P2_U3151), .B1(n10175), .B2(n8382), .C1(
        n8379), .C2(n10173), .ZN(P2_U3273) );
  OAI222_X1 U9741 ( .A1(n10696), .A2(n8383), .B1(n9271), .B2(n8382), .C1(
        P1_U3086), .C2(n8381), .ZN(P1_U3333) );
  INV_X1 U9742 ( .A(n8384), .ZN(n8386) );
  OAI222_X1 U9743 ( .A1(P2_U3151), .A2(n8387), .B1(n10175), .B2(n8386), .C1(
        n8385), .C2(n10173), .ZN(P2_U3275) );
  OAI21_X1 U9744 ( .B1(n8389), .B2(n9589), .A(n8388), .ZN(n8391) );
  AOI222_X1 U9745 ( .A1(n10041), .A2(n8391), .B1(n9807), .B2(n10003), .C1(
        n8390), .C2(n10001), .ZN(n10981) );
  MUX2_X1 U9746 ( .A(n7889), .B(n10981), .S(n11015), .Z(n8399) );
  OAI21_X1 U9747 ( .B1(n8392), .B2(n8394), .A(n8393), .ZN(n10979) );
  OAI22_X1 U9748 ( .A1(n10030), .A2(n8396), .B1(n8395), .B2(n11010), .ZN(n8397) );
  AOI21_X1 U9749 ( .B1(n10033), .B2(n10979), .A(n8397), .ZN(n8398) );
  NAND2_X1 U9750 ( .A1(n8399), .A2(n8398), .ZN(P2_U3232) );
  XNOR2_X1 U9751 ( .A(n8400), .B(n8404), .ZN(n8402) );
  OAI22_X1 U9752 ( .A1(n9070), .A2(n11001), .B1(n11003), .B2(n9153), .ZN(n8401) );
  AOI21_X1 U9753 ( .B1(n8402), .B2(n10041), .A(n8401), .ZN(n11161) );
  INV_X2 U9754 ( .A(n11015), .ZN(n11018) );
  OAI21_X1 U9755 ( .B1(n8405), .B2(n8404), .A(n8403), .ZN(n11160) );
  INV_X1 U9756 ( .A(n11157), .ZN(n9083) );
  AOI22_X1 U9757 ( .A1(n11018), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10028), 
        .B2(n9080), .ZN(n8406) );
  OAI21_X1 U9758 ( .B1(n9083), .B2(n10030), .A(n8406), .ZN(n8407) );
  AOI21_X1 U9759 ( .B1(n11160), .B2(n10033), .A(n8407), .ZN(n8408) );
  OAI21_X1 U9760 ( .B1(n11161), .B2(n11018), .A(n8408), .ZN(P2_U3221) );
  INV_X1 U9761 ( .A(n8414), .ZN(n9602) );
  XNOR2_X1 U9762 ( .A(n8409), .B(n9602), .ZN(n8412) );
  OAI22_X1 U9763 ( .A1(n9495), .A2(n11003), .B1(n11001), .B2(n8410), .ZN(n8411) );
  AOI21_X1 U9764 ( .B1(n8412), .B2(n10041), .A(n8411), .ZN(n11145) );
  OAI21_X1 U9765 ( .B1(n8415), .B2(n8414), .A(n8413), .ZN(n11144) );
  INV_X1 U9766 ( .A(n11143), .ZN(n9038) );
  NOR2_X1 U9767 ( .A1(n9038), .A2(n10030), .ZN(n8418) );
  INV_X1 U9768 ( .A(n9035), .ZN(n8416) );
  OAI22_X1 U9769 ( .A1(n11015), .A2(n8439), .B1(n8416), .B2(n11010), .ZN(n8417) );
  AOI211_X1 U9770 ( .C1(n11144), .C2(n10033), .A(n8418), .B(n8417), .ZN(n8419)
         );
  OAI21_X1 U9771 ( .B1(n11018), .B2(n11145), .A(n8419), .ZN(P2_U3222) );
  NAND2_X1 U9772 ( .A1(n8422), .A2(n8421), .ZN(n9600) );
  XNOR2_X1 U9773 ( .A(n8420), .B(n9600), .ZN(n8429) );
  INV_X1 U9774 ( .A(n9600), .ZN(n8423) );
  XNOR2_X1 U9775 ( .A(n8424), .B(n8423), .ZN(n11134) );
  INV_X1 U9776 ( .A(n9660), .ZN(n8427) );
  OAI22_X1 U9777 ( .A1(n8425), .A2(n11001), .B1(n11003), .B2(n9070), .ZN(n8426) );
  AOI21_X1 U9778 ( .B1(n11134), .B2(n8427), .A(n8426), .ZN(n8428) );
  OAI21_X1 U9779 ( .B1(n11000), .B2(n8429), .A(n8428), .ZN(n11137) );
  INV_X1 U9780 ( .A(n11137), .ZN(n8435) );
  NOR2_X1 U9781 ( .A1(n11018), .A2(n8430), .ZN(n9668) );
  INV_X1 U9782 ( .A(n11139), .ZN(n8432) );
  AOI22_X1 U9783 ( .A1(n11018), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10028), 
        .B2(n8998), .ZN(n8431) );
  OAI21_X1 U9784 ( .B1(n8432), .B2(n10030), .A(n8431), .ZN(n8433) );
  AOI21_X1 U9785 ( .B1(n11134), .B2(n9668), .A(n8433), .ZN(n8434) );
  OAI21_X1 U9786 ( .B1(n8435), .B2(n11018), .A(n8434), .ZN(P2_U3223) );
  AOI21_X1 U9787 ( .B1(n11147), .B2(n8437), .A(n8436), .ZN(n8452) );
  AOI21_X1 U9788 ( .B1(n8440), .B2(n8439), .A(n8438), .ZN(n8448) );
  NAND2_X1 U9789 ( .A1(n10959), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8447) );
  OAI21_X1 U9790 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8445) );
  INV_X1 U9791 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8444) );
  NOR2_X1 U9792 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8444), .ZN(n9032) );
  AOI21_X1 U9793 ( .B1(n8445), .B2(n5272), .A(n9032), .ZN(n8446) );
  OAI211_X1 U9794 ( .C1(n8448), .C2(n10972), .A(n8447), .B(n8446), .ZN(n8449)
         );
  AOI21_X1 U9795 ( .B1(n8450), .B2(n9881), .A(n8449), .ZN(n8451) );
  OAI21_X1 U9796 ( .B1(n8452), .B2(n10967), .A(n8451), .ZN(P2_U3193) );
  XOR2_X1 U9797 ( .A(n8453), .B(n8458), .Z(n8454) );
  AOI222_X1 U9798 ( .A1(n11232), .A2(n8454), .B1(n10327), .B2(n11236), .C1(
        n10325), .C2(n11237), .ZN(n11167) );
  NAND2_X1 U9799 ( .A1(n8456), .A2(n8455), .ZN(n8939) );
  OR2_X1 U9800 ( .A1(n8457), .A2(n10327), .ZN(n8937) );
  NAND2_X1 U9801 ( .A1(n8939), .A2(n8937), .ZN(n8479) );
  XOR2_X1 U9802 ( .A(n8458), .B(n8479), .Z(n11170) );
  OAI211_X1 U9803 ( .C1(n8459), .C2(n11168), .A(n11250), .B(n8484), .ZN(n11166) );
  NAND2_X1 U9804 ( .A1(n11258), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8460) );
  OAI21_X1 U9805 ( .B1(n10580), .B2(n8984), .A(n8460), .ZN(n8461) );
  AOI21_X1 U9806 ( .B1(n8480), .B2(n11245), .A(n8461), .ZN(n8462) );
  OAI21_X1 U9807 ( .B1(n11166), .B2(n11253), .A(n8462), .ZN(n8463) );
  AOI21_X1 U9808 ( .B1(n11170), .B2(n11218), .A(n8463), .ZN(n8464) );
  OAI21_X1 U9809 ( .B1(n11258), .B2(n11167), .A(n8464), .ZN(P1_U3281) );
  NAND2_X1 U9810 ( .A1(n8491), .A2(n8465), .ZN(n8467) );
  INV_X1 U9811 ( .A(n8466), .ZN(n8494) );
  AOI21_X1 U9812 ( .B1(n8468), .B2(n8467), .A(n8494), .ZN(n8476) );
  NAND2_X1 U9813 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10930) );
  INV_X1 U9814 ( .A(n10930), .ZN(n8472) );
  OAI22_X1 U9815 ( .A1(n10313), .A2(n8470), .B1(n10299), .B2(n8469), .ZN(n8471) );
  AOI211_X1 U9816 ( .C1(n10315), .C2(n10327), .A(n8472), .B(n8471), .ZN(n8475)
         );
  NAND2_X1 U9817 ( .A1(n8473), .A2(n10289), .ZN(n8474) );
  OAI211_X1 U9818 ( .C1(n8476), .C2(n10292), .A(n8475), .B(n8474), .ZN(
        P1_U3217) );
  XOR2_X1 U9819 ( .A(n8477), .B(n8483), .Z(n8478) );
  AOI222_X1 U9820 ( .A1(n11232), .A2(n8478), .B1(n11210), .B2(n11237), .C1(
        n10326), .C2(n11236), .ZN(n11174) );
  NAND2_X1 U9821 ( .A1(n8480), .A2(n10326), .ZN(n8941) );
  NAND2_X1 U9822 ( .A1(n8479), .A2(n8941), .ZN(n8481) );
  OR2_X1 U9823 ( .A1(n8480), .A2(n10326), .ZN(n8935) );
  NAND2_X1 U9824 ( .A1(n8481), .A2(n8935), .ZN(n8482) );
  XOR2_X1 U9825 ( .A(n8483), .B(n8482), .Z(n11176) );
  AND2_X1 U9826 ( .A1(n9043), .A2(n8484), .ZN(n8485) );
  OR3_X1 U9827 ( .A1(n8485), .A2(n5250), .A3(n10609), .ZN(n11173) );
  NAND2_X1 U9828 ( .A1(n11258), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8486) );
  OAI21_X1 U9829 ( .B1(n10580), .B2(n9048), .A(n8486), .ZN(n8487) );
  AOI21_X1 U9830 ( .B1(n9043), .B2(n11245), .A(n8487), .ZN(n8488) );
  OAI21_X1 U9831 ( .B1(n11173), .B2(n11253), .A(n8488), .ZN(n8489) );
  AOI21_X1 U9832 ( .B1(n11176), .B2(n11218), .A(n8489), .ZN(n8490) );
  OAI21_X1 U9833 ( .B1(n11258), .B2(n11174), .A(n8490), .ZN(P1_U3280) );
  INV_X1 U9834 ( .A(n8491), .ZN(n8493) );
  NOR3_X1 U9835 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8496) );
  INV_X1 U9836 ( .A(n8495), .ZN(n8979) );
  OAI21_X1 U9837 ( .B1(n8496), .B2(n8979), .A(n10308), .ZN(n8502) );
  NAND2_X1 U9838 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10835) );
  INV_X1 U9839 ( .A(n10835), .ZN(n8500) );
  OAI22_X1 U9840 ( .A1(n10313), .A2(n8498), .B1(n10299), .B2(n8497), .ZN(n8499) );
  AOI211_X1 U9841 ( .C1(n10315), .C2(n10326), .A(n8500), .B(n8499), .ZN(n8501)
         );
  OAI211_X1 U9842 ( .C1(n11152), .C2(n10318), .A(n8502), .B(n8501), .ZN(
        P1_U3236) );
  NAND2_X1 U9843 ( .A1(n8506), .A2(n9214), .ZN(n8504) );
  NAND2_X1 U9844 ( .A1(n8503), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9629) );
  OAI211_X1 U9845 ( .C1(n8505), .C2(n10173), .A(n8504), .B(n9629), .ZN(
        P2_U3272) );
  NAND2_X1 U9846 ( .A1(n8506), .A2(n10693), .ZN(n8508) );
  OAI211_X1 U9847 ( .C1(n8824), .C2(n10696), .A(n8508), .B(n8507), .ZN(
        P1_U3332) );
  XOR2_X1 U9848 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n8512) );
  XNOR2_X1 U9849 ( .A(n8509), .B(keyinput_130), .ZN(n8511) );
  XNOR2_X1 U9850 ( .A(n8698), .B(keyinput_129), .ZN(n8510) );
  NAND3_X1 U9851 ( .A1(n8512), .A2(n8511), .A3(n8510), .ZN(n8516) );
  XOR2_X1 U9852 ( .A(SI_29_), .B(keyinput_131), .Z(n8515) );
  XNOR2_X1 U9853 ( .A(SI_27_), .B(keyinput_133), .ZN(n8514) );
  XNOR2_X1 U9854 ( .A(SI_28_), .B(keyinput_132), .ZN(n8513) );
  AOI211_X1 U9855 ( .C1(n8516), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8522)
         );
  XNOR2_X1 U9856 ( .A(SI_26_), .B(keyinput_134), .ZN(n8521) );
  XNOR2_X1 U9857 ( .A(n8517), .B(keyinput_136), .ZN(n8520) );
  XNOR2_X1 U9858 ( .A(n8518), .B(keyinput_135), .ZN(n8519) );
  OAI211_X1 U9859 ( .C1(n8522), .C2(n8521), .A(n8520), .B(n8519), .ZN(n8525)
         );
  XNOR2_X1 U9860 ( .A(n8710), .B(keyinput_137), .ZN(n8524) );
  XNOR2_X1 U9861 ( .A(n8711), .B(keyinput_138), .ZN(n8523) );
  AOI21_X1 U9862 ( .B1(n8525), .B2(n8524), .A(n8523), .ZN(n8529) );
  XNOR2_X1 U9863 ( .A(SI_21_), .B(keyinput_139), .ZN(n8528) );
  XNOR2_X1 U9864 ( .A(n8716), .B(keyinput_140), .ZN(n8527) );
  XNOR2_X1 U9865 ( .A(SI_19_), .B(keyinput_141), .ZN(n8526) );
  OAI211_X1 U9866 ( .C1(n8529), .C2(n8528), .A(n8527), .B(n8526), .ZN(n8533)
         );
  XNOR2_X1 U9867 ( .A(SI_17_), .B(keyinput_143), .ZN(n8532) );
  XNOR2_X1 U9868 ( .A(SI_18_), .B(keyinput_142), .ZN(n8531) );
  XNOR2_X1 U9869 ( .A(SI_16_), .B(keyinput_144), .ZN(n8530) );
  NAND4_X1 U9870 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n8536)
         );
  XNOR2_X1 U9871 ( .A(n8728), .B(keyinput_145), .ZN(n8535) );
  XNOR2_X1 U9872 ( .A(n8729), .B(keyinput_146), .ZN(n8534) );
  NAND3_X1 U9873 ( .A1(n8536), .A2(n8535), .A3(n8534), .ZN(n8539) );
  XNOR2_X1 U9874 ( .A(n8733), .B(keyinput_148), .ZN(n8538) );
  XNOR2_X1 U9875 ( .A(SI_13_), .B(keyinput_147), .ZN(n8537) );
  NAND3_X1 U9876 ( .A1(n8539), .A2(n8538), .A3(n8537), .ZN(n8543) );
  XNOR2_X1 U9877 ( .A(SI_11_), .B(keyinput_149), .ZN(n8542) );
  XNOR2_X1 U9878 ( .A(n8739), .B(keyinput_150), .ZN(n8541) );
  XNOR2_X1 U9879 ( .A(n8738), .B(keyinput_151), .ZN(n8540) );
  AOI211_X1 U9880 ( .C1(n8543), .C2(n8542), .A(n8541), .B(n8540), .ZN(n8547)
         );
  XNOR2_X1 U9881 ( .A(SI_8_), .B(keyinput_152), .ZN(n8546) );
  XNOR2_X1 U9882 ( .A(SI_7_), .B(keyinput_153), .ZN(n8545) );
  XNOR2_X1 U9883 ( .A(SI_6_), .B(keyinput_154), .ZN(n8544) );
  OAI211_X1 U9884 ( .C1(n8547), .C2(n8546), .A(n8545), .B(n8544), .ZN(n8551)
         );
  XNOR2_X1 U9885 ( .A(SI_5_), .B(keyinput_155), .ZN(n8550) );
  XNOR2_X1 U9886 ( .A(n8748), .B(keyinput_156), .ZN(n8549) );
  XNOR2_X1 U9887 ( .A(SI_3_), .B(keyinput_157), .ZN(n8548) );
  AOI211_X1 U9888 ( .C1(n8551), .C2(n8550), .A(n8549), .B(n8548), .ZN(n8559)
         );
  XNOR2_X1 U9889 ( .A(n8552), .B(keyinput_158), .ZN(n8556) );
  XNOR2_X1 U9890 ( .A(SI_0_), .B(keyinput_160), .ZN(n8555) );
  XNOR2_X1 U9891 ( .A(SI_1_), .B(keyinput_159), .ZN(n8554) );
  XNOR2_X1 U9892 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n8553) );
  NAND4_X1 U9893 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n8558)
         );
  XNOR2_X1 U9894 ( .A(P2_U3151), .B(keyinput_162), .ZN(n8557) );
  OAI21_X1 U9895 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8561) );
  XNOR2_X1 U9896 ( .A(n8760), .B(keyinput_163), .ZN(n8560) );
  NAND2_X1 U9897 ( .A1(n8561), .A2(n8560), .ZN(n8571) );
  XNOR2_X1 U9898 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n8567) );
  XNOR2_X1 U9899 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n8563)
         );
  XNOR2_X1 U9900 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n8562)
         );
  NAND2_X1 U9901 ( .A1(n8563), .A2(n8562), .ZN(n8566) );
  XNOR2_X1 U9902 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n8565)
         );
  XNOR2_X1 U9903 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n8564)
         );
  NOR4_X1 U9904 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n8570)
         );
  XNOR2_X1 U9905 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n8569)
         );
  XNOR2_X1 U9906 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n8568)
         );
  AOI211_X1 U9907 ( .C1(n8571), .C2(n8570), .A(n8569), .B(n8568), .ZN(n8581)
         );
  XNOR2_X1 U9908 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n8580) );
  XNOR2_X1 U9909 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n8573) );
  XNOR2_X1 U9910 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n8572)
         );
  NAND2_X1 U9911 ( .A1(n8573), .A2(n8572), .ZN(n8579) );
  XOR2_X1 U9912 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n8577) );
  XNOR2_X1 U9913 ( .A(n8778), .B(keyinput_173), .ZN(n8576) );
  XNOR2_X1 U9914 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n8575) );
  XNOR2_X1 U9915 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n8574)
         );
  NAND4_X1 U9916 ( .A1(n8577), .A2(n8576), .A3(n8575), .A4(n8574), .ZN(n8578)
         );
  NOR4_X1 U9917 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n8584)
         );
  XNOR2_X1 U9918 ( .A(n9727), .B(keyinput_178), .ZN(n8583) );
  XNOR2_X1 U9919 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n8582)
         );
  OAI21_X1 U9920 ( .B1(n8584), .B2(n8583), .A(n8582), .ZN(n8588) );
  XNOR2_X1 U9921 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n8587) );
  XNOR2_X1 U9922 ( .A(n8585), .B(keyinput_181), .ZN(n8586) );
  AOI21_X1 U9923 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8592) );
  XNOR2_X1 U9924 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n8591) );
  XNOR2_X1 U9925 ( .A(n9124), .B(keyinput_184), .ZN(n8590) );
  XNOR2_X1 U9926 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n8589)
         );
  OAI211_X1 U9927 ( .C1(n8592), .C2(n8591), .A(n8590), .B(n8589), .ZN(n8595)
         );
  XOR2_X1 U9928 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .Z(n8594) );
  XNOR2_X1 U9929 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n8593)
         );
  AOI21_X1 U9930 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8598) );
  XOR2_X1 U9931 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n8597) );
  XOR2_X1 U9932 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .Z(n8596) );
  OAI21_X1 U9933 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8602) );
  XNOR2_X1 U9934 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n8601) );
  XNOR2_X1 U9935 ( .A(n9207), .B(keyinput_191), .ZN(n8600) );
  XNOR2_X1 U9936 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n8599)
         );
  AOI211_X1 U9937 ( .C1(n8602), .C2(n8601), .A(n8600), .B(n8599), .ZN(n8605)
         );
  XNOR2_X1 U9938 ( .A(n8809), .B(keyinput_192), .ZN(n8604) );
  XOR2_X1 U9939 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n8603) );
  NOR3_X1 U9940 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8612) );
  XNOR2_X1 U9941 ( .A(n9272), .B(keyinput_194), .ZN(n8611) );
  XNOR2_X1 U9942 ( .A(n9176), .B(keyinput_197), .ZN(n8609) );
  XNOR2_X1 U9943 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n8608)
         );
  XNOR2_X1 U9944 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n8607)
         );
  XNOR2_X1 U9945 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n8606)
         );
  NOR4_X1 U9946 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n8610)
         );
  OAI21_X1 U9947 ( .B1(n8612), .B2(n8611), .A(n8610), .ZN(n8615) );
  XNOR2_X1 U9948 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n8614)
         );
  XNOR2_X1 U9949 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n8613)
         );
  AOI21_X1 U9950 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8622) );
  XNOR2_X1 U9951 ( .A(n8824), .B(keyinput_201), .ZN(n8619) );
  XNOR2_X1 U9952 ( .A(n8823), .B(keyinput_204), .ZN(n8618) );
  XNOR2_X1 U9953 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n8617)
         );
  XNOR2_X1 U9954 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n8616)
         );
  NAND4_X1 U9955 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n8621)
         );
  XNOR2_X1 U9956 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n8620)
         );
  OAI21_X1 U9957 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8625) );
  XNOR2_X1 U9958 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n8624)
         );
  XNOR2_X1 U9959 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n8623)
         );
  NAND3_X1 U9960 ( .A1(n8625), .A2(n8624), .A3(n8623), .ZN(n8629) );
  XNOR2_X1 U9961 ( .A(n8626), .B(keyinput_208), .ZN(n8628) );
  XOR2_X1 U9962 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n8627) );
  NAND3_X1 U9963 ( .A1(n8629), .A2(n8628), .A3(n8627), .ZN(n8633) );
  XNOR2_X1 U9964 ( .A(n8630), .B(keyinput_210), .ZN(n8632) );
  XOR2_X1 U9965 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n8631) );
  AOI21_X1 U9966 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(n8640) );
  XNOR2_X1 U9967 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n8639)
         );
  XNOR2_X1 U9968 ( .A(n8842), .B(keyinput_215), .ZN(n8637) );
  XNOR2_X1 U9969 ( .A(n8841), .B(keyinput_216), .ZN(n8636) );
  XNOR2_X1 U9970 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n8635)
         );
  XNOR2_X1 U9971 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n8634)
         );
  NOR4_X1 U9972 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n8638)
         );
  OAI21_X1 U9973 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8647) );
  XOR2_X1 U9974 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n8644) );
  XNOR2_X1 U9975 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_220), .ZN(n8643) );
  XNOR2_X1 U9976 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .ZN(n8642) );
  XNOR2_X1 U9977 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .ZN(n8641) );
  NOR4_X1 U9978 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n8646)
         );
  XNOR2_X1 U9979 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n8645) );
  AOI21_X1 U9980 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8652) );
  XNOR2_X1 U9981 ( .A(n8648), .B(keyinput_223), .ZN(n8651) );
  XNOR2_X1 U9982 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n8650) );
  XNOR2_X1 U9983 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .ZN(n8649) );
  NOR4_X1 U9984 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n8657)
         );
  XNOR2_X1 U9985 ( .A(n8653), .B(keyinput_225), .ZN(n8656) );
  XNOR2_X1 U9986 ( .A(n8867), .B(keyinput_226), .ZN(n8655) );
  XNOR2_X1 U9987 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_227), .ZN(n8654) );
  NOR4_X1 U9988 ( .A1(n8657), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n8664)
         );
  XNOR2_X1 U9989 ( .A(n8872), .B(keyinput_228), .ZN(n8663) );
  XOR2_X1 U9990 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_229), .Z(n8661) );
  XNOR2_X1 U9991 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .ZN(n8660) );
  XNOR2_X1 U9992 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n8659) );
  XNOR2_X1 U9993 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n8658) );
  NOR4_X1 U9994 ( .A1(n8661), .A2(n8660), .A3(n8659), .A4(n8658), .ZN(n8662)
         );
  OAI21_X1 U9995 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8668) );
  XNOR2_X1 U9996 ( .A(n8881), .B(keyinput_233), .ZN(n8667) );
  XOR2_X1 U9997 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .Z(n8666) );
  XNOR2_X1 U9998 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n8665) );
  NAND4_X1 U9999 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n8672)
         );
  XNOR2_X1 U10000 ( .A(n8886), .B(keyinput_236), .ZN(n8671) );
  XNOR2_X1 U10001 ( .A(n8669), .B(keyinput_237), .ZN(n8670) );
  NAND3_X1 U10002 ( .A1(n8672), .A2(n8671), .A3(n8670), .ZN(n8676) );
  XNOR2_X1 U10003 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n8675) );
  XOR2_X1 U10004 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .Z(n8674) );
  XOR2_X1 U10005 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_239), .Z(n8673) );
  AOI211_X1 U10006 ( .C1(n8676), .C2(n8675), .A(n8674), .B(n8673), .ZN(n8680)
         );
  XNOR2_X1 U10007 ( .A(n8677), .B(keyinput_241), .ZN(n8679) );
  XNOR2_X1 U10008 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .ZN(n8678) );
  OAI21_X1 U10009 ( .B1(n8680), .B2(n8679), .A(n8678), .ZN(n8683) );
  XNOR2_X1 U10010 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n8682) );
  XNOR2_X1 U10011 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .ZN(n8681) );
  AOI21_X1 U10012 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(n8686) );
  XNOR2_X1 U10013 ( .A(n8903), .B(keyinput_245), .ZN(n8685) );
  XNOR2_X1 U10014 ( .A(n8904), .B(keyinput_246), .ZN(n8684) );
  OAI21_X1 U10015 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n8693) );
  XOR2_X1 U10016 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .Z(n8690) );
  XOR2_X1 U10017 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .Z(n8689) );
  XNOR2_X1 U10018 ( .A(n8908), .B(keyinput_247), .ZN(n8688) );
  XNOR2_X1 U10019 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n8687) );
  NOR4_X1 U10020 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n8692)
         );
  XOR2_X1 U10021 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .Z(n8691) );
  AOI21_X1 U10022 ( .B1(n8693), .B2(n8692), .A(n8691), .ZN(n8697) );
  INV_X1 U10023 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10701) );
  XNOR2_X1 U10024 ( .A(n10701), .B(keyinput_253), .ZN(n8696) );
  XNOR2_X1 U10025 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_254), .ZN(n8695) );
  XNOR2_X1 U10026 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_252), .ZN(n8694) );
  NOR4_X1 U10027 ( .A1(n8697), .A2(n8696), .A3(n8695), .A4(n8694), .ZN(n8923)
         );
  XNOR2_X1 U10028 ( .A(keyinput_127), .B(keyinput_255), .ZN(n8922) );
  XNOR2_X1 U10029 ( .A(keyinput_127), .B(P1_D_REG_5__SCAN_IN), .ZN(n8921) );
  XOR2_X1 U10030 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n8701) );
  XNOR2_X1 U10031 ( .A(n8698), .B(keyinput_1), .ZN(n8700) );
  XNOR2_X1 U10032 ( .A(SI_30_), .B(keyinput_2), .ZN(n8699) );
  NAND3_X1 U10033 ( .A1(n8701), .A2(n8700), .A3(n8699), .ZN(n8705) );
  XOR2_X1 U10034 ( .A(SI_29_), .B(keyinput_3), .Z(n8704) );
  XNOR2_X1 U10035 ( .A(SI_28_), .B(keyinput_4), .ZN(n8703) );
  XNOR2_X1 U10036 ( .A(SI_27_), .B(keyinput_5), .ZN(n8702) );
  AOI211_X1 U10037 ( .C1(n8705), .C2(n8704), .A(n8703), .B(n8702), .ZN(n8709)
         );
  XNOR2_X1 U10038 ( .A(SI_26_), .B(keyinput_6), .ZN(n8708) );
  XNOR2_X1 U10039 ( .A(SI_25_), .B(keyinput_7), .ZN(n8707) );
  XNOR2_X1 U10040 ( .A(SI_24_), .B(keyinput_8), .ZN(n8706) );
  OAI211_X1 U10041 ( .C1(n8709), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8714)
         );
  XNOR2_X1 U10042 ( .A(n8710), .B(keyinput_9), .ZN(n8713) );
  XNOR2_X1 U10043 ( .A(n8711), .B(keyinput_10), .ZN(n8712) );
  AOI21_X1 U10044 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8720) );
  XNOR2_X1 U10045 ( .A(SI_21_), .B(keyinput_11), .ZN(n8719) );
  XNOR2_X1 U10046 ( .A(n8715), .B(keyinput_13), .ZN(n8718) );
  XNOR2_X1 U10047 ( .A(n8716), .B(keyinput_12), .ZN(n8717) );
  OAI211_X1 U10048 ( .C1(n8720), .C2(n8719), .A(n8718), .B(n8717), .ZN(n8727)
         );
  XNOR2_X1 U10049 ( .A(n8721), .B(keyinput_14), .ZN(n8726) );
  XNOR2_X1 U10050 ( .A(n8722), .B(keyinput_16), .ZN(n8725) );
  XNOR2_X1 U10051 ( .A(n8723), .B(keyinput_15), .ZN(n8724) );
  NAND4_X1 U10052 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n8732)
         );
  XNOR2_X1 U10053 ( .A(n8728), .B(keyinput_17), .ZN(n8731) );
  XNOR2_X1 U10054 ( .A(n8729), .B(keyinput_18), .ZN(n8730) );
  NAND3_X1 U10055 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(n8736) );
  XNOR2_X1 U10056 ( .A(n8733), .B(keyinput_20), .ZN(n8735) );
  XOR2_X1 U10057 ( .A(SI_13_), .B(keyinput_19), .Z(n8734) );
  NAND3_X1 U10058 ( .A1(n8736), .A2(n8735), .A3(n8734), .ZN(n8743) );
  XNOR2_X1 U10059 ( .A(n8737), .B(keyinput_21), .ZN(n8742) );
  XNOR2_X1 U10060 ( .A(n8738), .B(keyinput_23), .ZN(n8741) );
  XNOR2_X1 U10061 ( .A(n8739), .B(keyinput_22), .ZN(n8740) );
  AOI211_X1 U10062 ( .C1(n8743), .C2(n8742), .A(n8741), .B(n8740), .ZN(n8747)
         );
  XNOR2_X1 U10063 ( .A(SI_8_), .B(keyinput_24), .ZN(n8746) );
  XOR2_X1 U10064 ( .A(SI_6_), .B(keyinput_26), .Z(n8745) );
  XNOR2_X1 U10065 ( .A(SI_7_), .B(keyinput_25), .ZN(n8744) );
  OAI211_X1 U10066 ( .C1(n8747), .C2(n8746), .A(n8745), .B(n8744), .ZN(n8752)
         );
  XOR2_X1 U10067 ( .A(SI_5_), .B(keyinput_27), .Z(n8751) );
  XNOR2_X1 U10068 ( .A(n8748), .B(keyinput_28), .ZN(n8750) );
  XNOR2_X1 U10069 ( .A(SI_3_), .B(keyinput_29), .ZN(n8749) );
  AOI211_X1 U10070 ( .C1(n8752), .C2(n8751), .A(n8750), .B(n8749), .ZN(n8759)
         );
  XNOR2_X1 U10071 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n8756) );
  XNOR2_X1 U10072 ( .A(SI_1_), .B(keyinput_31), .ZN(n8755) );
  XNOR2_X1 U10073 ( .A(SI_2_), .B(keyinput_30), .ZN(n8754) );
  XNOR2_X1 U10074 ( .A(SI_0_), .B(keyinput_32), .ZN(n8753) );
  NAND4_X1 U10075 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n8758)
         );
  XNOR2_X1 U10076 ( .A(P2_U3151), .B(keyinput_34), .ZN(n8757) );
  OAI21_X1 U10077 ( .B1(n8759), .B2(n8758), .A(n8757), .ZN(n8762) );
  XNOR2_X1 U10078 ( .A(n8760), .B(keyinput_35), .ZN(n8761) );
  NAND2_X1 U10079 ( .A1(n8762), .A2(n8761), .ZN(n8771) );
  XNOR2_X1 U10080 ( .A(n8763), .B(keyinput_40), .ZN(n8770) );
  XOR2_X1 U10081 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n8767) );
  XNOR2_X1 U10082 ( .A(n8764), .B(keyinput_36), .ZN(n8766) );
  XNOR2_X1 U10083 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n8765)
         );
  NOR3_X1 U10084 ( .A1(n8767), .A2(n8766), .A3(n8765), .ZN(n8769) );
  XNOR2_X1 U10085 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n8768)
         );
  NAND4_X1 U10086 ( .A1(n8771), .A2(n8770), .A3(n8769), .A4(n8768), .ZN(n8774)
         );
  XNOR2_X1 U10087 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n8773)
         );
  XNOR2_X1 U10088 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n8772)
         );
  NAND3_X1 U10089 ( .A1(n8774), .A2(n8773), .A3(n8772), .ZN(n8786) );
  INV_X1 U10090 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9241) );
  OAI22_X1 U10091 ( .A1(n9241), .A2(keyinput_48), .B1(keyinput_46), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n8775) );
  AOI221_X1 U10092 ( .B1(n9241), .B2(keyinput_48), .C1(P2_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n8775), .ZN(n8785) );
  OAI22_X1 U10093 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        keyinput_49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n8776) );
  AOI221_X1 U10094 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n8776), .ZN(n8783) );
  INV_X1 U10095 ( .A(keyinput_44), .ZN(n8777) );
  XNOR2_X1 U10096 ( .A(n8777), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n8782) );
  XNOR2_X1 U10097 ( .A(n8778), .B(keyinput_45), .ZN(n8781) );
  XNOR2_X1 U10098 ( .A(n8779), .B(keyinput_47), .ZN(n8780) );
  AND4_X1 U10099 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n8784)
         );
  NAND3_X1 U10100 ( .A1(n8786), .A2(n8785), .A3(n8784), .ZN(n8789) );
  XNOR2_X1 U10101 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n8788)
         );
  XNOR2_X1 U10102 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n8787)
         );
  AOI21_X1 U10103 ( .B1(n8789), .B2(n8788), .A(n8787), .ZN(n8793) );
  XNOR2_X1 U10104 ( .A(n8790), .B(keyinput_52), .ZN(n8792) );
  XNOR2_X1 U10105 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n8791) );
  OAI21_X1 U10106 ( .B1(n8793), .B2(n8792), .A(n8791), .ZN(n8798) );
  XOR2_X1 U10107 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n8797) );
  XNOR2_X1 U10108 ( .A(n8794), .B(keyinput_55), .ZN(n8796) );
  XNOR2_X1 U10109 ( .A(n9124), .B(keyinput_56), .ZN(n8795) );
  AOI211_X1 U10110 ( .C1(n8798), .C2(n8797), .A(n8796), .B(n8795), .ZN(n8801)
         );
  XNOR2_X1 U10111 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n8800)
         );
  XNOR2_X1 U10112 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n8799)
         );
  OAI21_X1 U10113 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8804) );
  XOR2_X1 U10114 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n8803) );
  XNOR2_X1 U10115 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n8802)
         );
  AOI21_X1 U10116 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8808) );
  XNOR2_X1 U10117 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n8807) );
  XNOR2_X1 U10118 ( .A(n9207), .B(keyinput_63), .ZN(n8806) );
  XNOR2_X1 U10119 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n8805)
         );
  OAI211_X1 U10120 ( .C1(n8808), .C2(n8807), .A(n8806), .B(n8805), .ZN(n8812)
         );
  XNOR2_X1 U10121 ( .A(n8809), .B(keyinput_64), .ZN(n8811) );
  XNOR2_X1 U10122 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n8810)
         );
  NAND3_X1 U10123 ( .A1(n8812), .A2(n8811), .A3(n8810), .ZN(n8819) );
  XNOR2_X1 U10124 ( .A(n9272), .B(keyinput_66), .ZN(n8818) );
  XNOR2_X1 U10125 ( .A(n9111), .B(keyinput_70), .ZN(n8816) );
  XOR2_X1 U10126 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n8815) );
  XNOR2_X1 U10127 ( .A(n9176), .B(keyinput_69), .ZN(n8814) );
  XNOR2_X1 U10128 ( .A(n10697), .B(keyinput_67), .ZN(n8813) );
  NAND4_X1 U10129 ( .A1(n8816), .A2(n8815), .A3(n8814), .A4(n8813), .ZN(n8817)
         );
  AOI21_X1 U10130 ( .B1(n8819), .B2(n8818), .A(n8817), .ZN(n8822) );
  XNOR2_X1 U10131 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n8821)
         );
  XNOR2_X1 U10132 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n8820)
         );
  OAI21_X1 U10133 ( .B1(n8822), .B2(n8821), .A(n8820), .ZN(n8831) );
  XNOR2_X1 U10134 ( .A(n8823), .B(keyinput_76), .ZN(n8828) );
  XNOR2_X1 U10135 ( .A(n8824), .B(keyinput_73), .ZN(n8827) );
  XNOR2_X1 U10136 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n8826)
         );
  XNOR2_X1 U10137 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n8825)
         );
  NOR4_X1 U10138 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(n8830)
         );
  XNOR2_X1 U10139 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n8829)
         );
  AOI21_X1 U10140 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8834) );
  XOR2_X1 U10141 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n8833) );
  XNOR2_X1 U10142 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n8832)
         );
  NOR3_X1 U10143 ( .A1(n8834), .A2(n8833), .A3(n8832), .ZN(n8837) );
  XNOR2_X1 U10144 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n8836)
         );
  XNOR2_X1 U10145 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n8835)
         );
  NOR3_X1 U10146 ( .A1(n8837), .A2(n8836), .A3(n8835), .ZN(n8840) );
  XNOR2_X1 U10147 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n8839)
         );
  XNOR2_X1 U10148 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n8838)
         );
  OAI21_X1 U10149 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8849) );
  XNOR2_X1 U10150 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n8848)
         );
  XNOR2_X1 U10151 ( .A(n8841), .B(keyinput_88), .ZN(n8846) );
  XNOR2_X1 U10152 ( .A(n8842), .B(keyinput_87), .ZN(n8845) );
  XNOR2_X1 U10153 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n8844)
         );
  XNOR2_X1 U10154 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n8843)
         );
  NAND4_X1 U10155 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n8847)
         );
  AOI21_X1 U10156 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8859) );
  XOR2_X1 U10157 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n8855) );
  XNOR2_X1 U10158 ( .A(n8850), .B(keyinput_92), .ZN(n8854) );
  XNOR2_X1 U10159 ( .A(n8851), .B(keyinput_91), .ZN(n8853) );
  XNOR2_X1 U10160 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_90), .ZN(n8852) );
  NAND4_X1 U10161 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n8858)
         );
  XNOR2_X1 U10162 ( .A(n8856), .B(keyinput_93), .ZN(n8857) );
  OAI21_X1 U10163 ( .B1(n8859), .B2(n8858), .A(n8857), .ZN(n8865) );
  XNOR2_X1 U10164 ( .A(n8860), .B(keyinput_96), .ZN(n8864) );
  XNOR2_X1 U10165 ( .A(n8861), .B(keyinput_94), .ZN(n8863) );
  XNOR2_X1 U10166 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n8862) );
  NAND4_X1 U10167 ( .A1(n8865), .A2(n8864), .A3(n8863), .A4(n8862), .ZN(n8871)
         );
  XNOR2_X1 U10168 ( .A(n8866), .B(keyinput_99), .ZN(n8870) );
  XNOR2_X1 U10169 ( .A(n8867), .B(keyinput_98), .ZN(n8869) );
  XNOR2_X1 U10170 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .ZN(n8868) );
  NAND4_X1 U10171 ( .A1(n8871), .A2(n8870), .A3(n8869), .A4(n8868), .ZN(n8880)
         );
  XNOR2_X1 U10172 ( .A(n8872), .B(keyinput_100), .ZN(n8879) );
  XOR2_X1 U10173 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .Z(n8877) );
  XOR2_X1 U10174 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .Z(n8876) );
  XOR2_X1 U10175 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .Z(n8875) );
  XNOR2_X1 U10176 ( .A(n8873), .B(keyinput_104), .ZN(n8874) );
  NAND4_X1 U10177 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8878)
         );
  AOI21_X1 U10178 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8885) );
  XOR2_X1 U10179 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .Z(n8884) );
  XNOR2_X1 U10180 ( .A(n8881), .B(keyinput_105), .ZN(n8883) );
  XNOR2_X1 U10181 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n8882) );
  NOR4_X1 U10182 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(n8889)
         );
  XNOR2_X1 U10183 ( .A(n8886), .B(keyinput_108), .ZN(n8888) );
  XNOR2_X1 U10184 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_109), .ZN(n8887) );
  NOR3_X1 U10185 ( .A1(n8889), .A2(n8888), .A3(n8887), .ZN(n8894) );
  XNOR2_X1 U10186 ( .A(n8890), .B(keyinput_110), .ZN(n8893) );
  XOR2_X1 U10187 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_112), .Z(n8892) );
  XNOR2_X1 U10188 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_111), .ZN(n8891) );
  OAI211_X1 U10189 ( .C1(n8894), .C2(n8893), .A(n8892), .B(n8891), .ZN(n8898)
         );
  XNOR2_X1 U10190 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n8897) );
  XNOR2_X1 U10191 ( .A(n8895), .B(keyinput_114), .ZN(n8896) );
  AOI21_X1 U10192 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8902) );
  XNOR2_X1 U10193 ( .A(n8899), .B(keyinput_115), .ZN(n8901) );
  XNOR2_X1 U10194 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n8900) );
  OAI21_X1 U10195 ( .B1(n8902), .B2(n8901), .A(n8900), .ZN(n8907) );
  XNOR2_X1 U10196 ( .A(n8903), .B(keyinput_117), .ZN(n8906) );
  XNOR2_X1 U10197 ( .A(n8904), .B(keyinput_118), .ZN(n8905) );
  AOI21_X1 U10198 ( .B1(n8907), .B2(n8906), .A(n8905), .ZN(n8915) );
  XOR2_X1 U10199 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .Z(n8912) );
  XNOR2_X1 U10200 ( .A(n8908), .B(keyinput_119), .ZN(n8911) );
  XNOR2_X1 U10201 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n8910) );
  XNOR2_X1 U10202 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .ZN(n8909) );
  NAND4_X1 U10203 ( .A1(n8912), .A2(n8911), .A3(n8910), .A4(n8909), .ZN(n8914)
         );
  XOR2_X1 U10204 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .Z(n8913) );
  OAI21_X1 U10205 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8919) );
  XNOR2_X1 U10206 ( .A(n10701), .B(keyinput_125), .ZN(n8918) );
  XOR2_X1 U10207 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_124), .Z(n8917) );
  XOR2_X1 U10208 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_126), .Z(n8916) );
  NAND4_X1 U10209 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n8920)
         );
  OAI211_X1 U10210 ( .C1(n8923), .C2(n8922), .A(n8921), .B(n8920), .ZN(n8934)
         );
  AOI21_X1 U10211 ( .B1(n11111), .B2(n8925), .A(n8924), .ZN(n8926) );
  OAI211_X1 U10212 ( .C1(n8928), .C2(n10671), .A(n8927), .B(n8926), .ZN(n10993) );
  MUX2_X1 U10213 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10993), .S(n11276), .Z(
        n8933) );
  XNOR2_X1 U10214 ( .A(n8934), .B(n8933), .ZN(P1_U3524) );
  NAND2_X1 U10215 ( .A1(n9043), .A2(n10325), .ZN(n8940) );
  AND2_X1 U10216 ( .A1(n8937), .A2(n8942), .ZN(n8938) );
  NAND2_X1 U10217 ( .A1(n8939), .A2(n8938), .ZN(n9140) );
  NAND2_X1 U10218 ( .A1(n8942), .A2(n5183), .ZN(n9138) );
  NAND2_X1 U10219 ( .A1(n9140), .A2(n9138), .ZN(n8943) );
  XNOR2_X1 U10220 ( .A(n8943), .B(n7053), .ZN(n11196) );
  INV_X1 U10221 ( .A(n11196), .ZN(n8955) );
  INV_X1 U10222 ( .A(n11207), .ZN(n8944) );
  AOI21_X1 U10223 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8950) );
  INV_X1 U10224 ( .A(n8947), .ZN(n11077) );
  NAND2_X1 U10225 ( .A1(n11196), .A2(n11077), .ZN(n8949) );
  AOI22_X1 U10226 ( .A1(n11237), .A2(n10594), .B1(n10325), .B2(n11236), .ZN(
        n8948) );
  OAI211_X1 U10227 ( .C1(n10503), .C2(n8950), .A(n8949), .B(n8948), .ZN(n11194) );
  NAND2_X1 U10228 ( .A1(n11194), .A2(n10600), .ZN(n8954) );
  OAI22_X1 U10229 ( .A1(n10600), .A2(n10392), .B1(n9102), .B2(n10580), .ZN(
        n8952) );
  INV_X1 U10230 ( .A(n9141), .ZN(n11193) );
  OAI211_X1 U10231 ( .C1(n11193), .C2(n5250), .A(n11250), .B(n11203), .ZN(
        n11192) );
  NOR2_X1 U10232 ( .A1(n11192), .A2(n11253), .ZN(n8951) );
  AOI211_X1 U10233 ( .C1(n11245), .C2(n9141), .A(n8952), .B(n8951), .ZN(n8953)
         );
  OAI211_X1 U10234 ( .C1(n8955), .C2(n9267), .A(n8954), .B(n8953), .ZN(
        P1_U3279) );
  INV_X1 U10235 ( .A(n8956), .ZN(n9500) );
  NAND2_X1 U10236 ( .A1(n9499), .A2(n9500), .ZN(n9604) );
  XNOR2_X1 U10237 ( .A(n8957), .B(n9604), .ZN(n11182) );
  INV_X1 U10238 ( .A(n9795), .ZN(n9505) );
  XNOR2_X1 U10239 ( .A(n8958), .B(n9604), .ZN(n8959) );
  OAI222_X1 U10240 ( .A1(n11003), .A2(n9505), .B1(n11001), .B2(n9495), .C1(
        n8959), .C2(n11000), .ZN(n11184) );
  NAND2_X1 U10241 ( .A1(n11184), .A2(n11015), .ZN(n8963) );
  INV_X1 U10242 ( .A(n9169), .ZN(n8960) );
  OAI22_X1 U10243 ( .A1(n11015), .A2(n9119), .B1(n8960), .B2(n11010), .ZN(
        n8961) );
  AOI21_X1 U10244 ( .B1(n9152), .B2(n10015), .A(n8961), .ZN(n8962) );
  OAI211_X1 U10245 ( .C1(n11182), .C2(n10012), .A(n8963), .B(n8962), .ZN(
        P2_U3220) );
  NAND2_X1 U10246 ( .A1(n8964), .A2(n9605), .ZN(n8965) );
  NAND3_X1 U10247 ( .A1(n9062), .A2(n10041), .A3(n8965), .ZN(n8968) );
  OAI22_X1 U10248 ( .A1(n9153), .A2(n11001), .B1(n11003), .B2(n9244), .ZN(
        n8966) );
  INV_X1 U10249 ( .A(n8966), .ZN(n8967) );
  AND2_X1 U10250 ( .A1(n8968), .A2(n8967), .ZN(n10105) );
  INV_X1 U10251 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8970) );
  INV_X1 U10252 ( .A(n9197), .ZN(n8969) );
  OAI22_X1 U10253 ( .A1(n11015), .A2(n8970), .B1(n8969), .B2(n11010), .ZN(
        n8971) );
  AOI21_X1 U10254 ( .B1(n10164), .B2(n10015), .A(n8971), .ZN(n8975) );
  XNOR2_X1 U10255 ( .A(n8972), .B(n8973), .ZN(n10104) );
  NAND2_X1 U10256 ( .A1(n10104), .A2(n10033), .ZN(n8974) );
  OAI211_X1 U10257 ( .C1(n10105), .C2(n11018), .A(n8975), .B(n8974), .ZN(
        P2_U3219) );
  INV_X1 U10258 ( .A(n8976), .ZN(n8978) );
  NOR3_X1 U10259 ( .A1(n8979), .A2(n8978), .A3(n8977), .ZN(n8982) );
  INV_X1 U10260 ( .A(n8980), .ZN(n8981) );
  OAI21_X1 U10261 ( .B1(n8982), .B2(n8981), .A(n10308), .ZN(n8988) );
  OAI22_X1 U10262 ( .A1(n10299), .A2(n8984), .B1(n8983), .B2(n10313), .ZN(
        n8985) );
  AOI211_X1 U10263 ( .C1(n10315), .C2(n10325), .A(n8986), .B(n8985), .ZN(n8987) );
  OAI211_X1 U10264 ( .C1(n11168), .C2(n10318), .A(n8988), .B(n8987), .ZN(
        P1_U3224) );
  NAND2_X1 U10265 ( .A1(n8990), .A2(n8989), .ZN(n8994) );
  INV_X1 U10266 ( .A(n8991), .ZN(n8992) );
  NAND2_X1 U10267 ( .A1(n8992), .A2(n9800), .ZN(n8993) );
  NAND2_X1 U10268 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  XNOR2_X1 U10269 ( .A(n11139), .B(n9355), .ZN(n8995) );
  AOI21_X1 U10270 ( .B1(n9799), .B2(n8997), .A(n5159), .ZN(n9004) );
  NAND2_X1 U10271 ( .A1(n9766), .A2(n8998), .ZN(n9001) );
  AOI21_X1 U10272 ( .B1(n9776), .B2(n9800), .A(n8999), .ZN(n9000) );
  OAI211_X1 U10273 ( .C1(n9070), .C2(n9754), .A(n9001), .B(n9000), .ZN(n9002)
         );
  AOI21_X1 U10274 ( .B1(n11139), .B2(n9731), .A(n9002), .ZN(n9003) );
  OAI21_X1 U10275 ( .B1(n9004), .B2(n9748), .A(n9003), .ZN(P2_U3157) );
  AOI21_X1 U10276 ( .B1(n5251), .B2(n9006), .A(n9005), .ZN(n9022) );
  INV_X1 U10277 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9013) );
  OAI21_X1 U10278 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9011) );
  NAND2_X1 U10279 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9077) );
  INV_X1 U10280 ( .A(n9077), .ZN(n9010) );
  AOI21_X1 U10281 ( .B1(n9011), .B2(n5272), .A(n9010), .ZN(n9012) );
  OAI21_X1 U10282 ( .B1(n9873), .B2(n9013), .A(n9012), .ZN(n9019) );
  AOI21_X1 U10283 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9017) );
  NOR2_X1 U10284 ( .A1(n9017), .A2(n10972), .ZN(n9018) );
  AOI211_X1 U10285 ( .C1(n9881), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9021)
         );
  OAI21_X1 U10286 ( .B1(n9022), .B2(n10967), .A(n9021), .ZN(P2_U3194) );
  INV_X1 U10287 ( .A(n9023), .ZN(n9041) );
  OAI222_X1 U10288 ( .A1(n9271), .A2(n9041), .B1(P1_U3086), .B2(n9025), .C1(
        n9024), .C2(n10696), .ZN(P1_U3331) );
  INV_X1 U10289 ( .A(n9027), .ZN(n9026) );
  XNOR2_X1 U10290 ( .A(n11143), .B(n9373), .ZN(n9071) );
  XNOR2_X1 U10291 ( .A(n9071), .B(n9798), .ZN(n9028) );
  NOR3_X1 U10292 ( .A1(n5159), .A2(n9026), .A3(n9028), .ZN(n9031) );
  NAND2_X1 U10293 ( .A1(n9029), .A2(n9028), .ZN(n9073) );
  INV_X1 U10294 ( .A(n9073), .ZN(n9030) );
  OAI21_X1 U10295 ( .B1(n9031), .B2(n9030), .A(n9773), .ZN(n9037) );
  AOI21_X1 U10296 ( .B1(n9776), .B2(n9799), .A(n9032), .ZN(n9033) );
  OAI21_X1 U10297 ( .B1(n9495), .B2(n9754), .A(n9033), .ZN(n9034) );
  AOI21_X1 U10298 ( .B1(n9035), .B2(n9766), .A(n9034), .ZN(n9036) );
  OAI211_X1 U10299 ( .C1(n9038), .C2(n9784), .A(n9037), .B(n9036), .ZN(
        P2_U3176) );
  INV_X1 U10300 ( .A(n9039), .ZN(n9042) );
  OAI222_X1 U10301 ( .A1(n9042), .A2(P2_U3151), .B1(n10175), .B2(n9041), .C1(
        n9040), .C2(n10173), .ZN(P2_U3271) );
  OAI21_X1 U10302 ( .B1(n9046), .B2(n9044), .A(n9045), .ZN(n9047) );
  NAND2_X1 U10303 ( .A1(n9047), .A2(n10308), .ZN(n9053) );
  NAND2_X1 U10304 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10915)
         );
  INV_X1 U10305 ( .A(n10915), .ZN(n9051) );
  OAI22_X1 U10306 ( .A1(n10313), .A2(n9049), .B1(n10299), .B2(n9048), .ZN(
        n9050) );
  AOI211_X1 U10307 ( .C1(n10315), .C2(n11210), .A(n9051), .B(n9050), .ZN(n9052) );
  OAI211_X1 U10308 ( .C1(n5417), .C2(n10318), .A(n9053), .B(n9052), .ZN(
        P1_U3234) );
  INV_X1 U10309 ( .A(n9054), .ZN(n9058) );
  OAI222_X1 U10310 ( .A1(n9271), .A2(n9058), .B1(P1_U3086), .B2(n9056), .C1(
        n9055), .C2(n10696), .ZN(P1_U3330) );
  OAI222_X1 U10311 ( .A1(n9059), .A2(P2_U3151), .B1(n10175), .B2(n9058), .C1(
        n9057), .C2(n10173), .ZN(P2_U3270) );
  XNOR2_X1 U10312 ( .A(n9060), .B(n9607), .ZN(n10100) );
  INV_X1 U10313 ( .A(n10100), .ZN(n9069) );
  NAND3_X1 U10314 ( .A1(n9062), .A2(n9607), .A3(n9514), .ZN(n9063) );
  NAND3_X1 U10315 ( .A1(n9061), .A2(n10041), .A3(n9063), .ZN(n9065) );
  OR2_X1 U10316 ( .A1(n9505), .A2(n11001), .ZN(n9064) );
  OAI211_X1 U10317 ( .C1(n10019), .C2(n11003), .A(n9065), .B(n9064), .ZN(
        n10099) );
  AOI22_X1 U10318 ( .A1(n11018), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10028), 
        .B2(n9211), .ZN(n9066) );
  OAI21_X1 U10319 ( .B1(n10161), .B2(n10030), .A(n9066), .ZN(n9067) );
  AOI21_X1 U10320 ( .B1(n10099), .B2(n11015), .A(n9067), .ZN(n9068) );
  OAI21_X1 U10321 ( .B1(n9069), .B2(n10012), .A(n9068), .ZN(P2_U3218) );
  NAND2_X1 U10322 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U10323 ( .A1(n9073), .A2(n9072), .ZN(n9075) );
  XNOR2_X1 U10324 ( .A(n11157), .B(n9373), .ZN(n9157) );
  XNOR2_X1 U10325 ( .A(n9157), .B(n9495), .ZN(n9074) );
  AOI21_X1 U10326 ( .B1(n9075), .B2(n9074), .A(n9748), .ZN(n9076) );
  NAND2_X1 U10327 ( .A1(n9076), .A2(n9160), .ZN(n9082) );
  NAND2_X1 U10328 ( .A1(n9776), .A2(n9798), .ZN(n9078) );
  OAI211_X1 U10329 ( .C1(n9153), .C2(n9754), .A(n9078), .B(n9077), .ZN(n9079)
         );
  AOI21_X1 U10330 ( .B1(n9080), .B2(n9766), .A(n9079), .ZN(n9081) );
  OAI211_X1 U10331 ( .C1(n9083), .C2(n9784), .A(n9082), .B(n9081), .ZN(
        P2_U3164) );
  NAND3_X1 U10332 ( .A1(n9061), .A2(n6452), .A3(n9084), .ZN(n9085) );
  NAND3_X1 U10333 ( .A1(n9086), .A2(n10041), .A3(n9085), .ZN(n9088) );
  OR2_X1 U10334 ( .A1(n11001), .A2(n9244), .ZN(n9087) );
  OAI211_X1 U10335 ( .C1(n9764), .C2(n11003), .A(n9088), .B(n9087), .ZN(n10095) );
  INV_X1 U10336 ( .A(n10095), .ZN(n9095) );
  INV_X1 U10337 ( .A(n9090), .ZN(n9091) );
  AOI21_X1 U10338 ( .B1(n9516), .B2(n9089), .A(n9091), .ZN(n10096) );
  INV_X1 U10339 ( .A(n9246), .ZN(n10156) );
  AOI22_X1 U10340 ( .A1(n11018), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10028), 
        .B2(n9240), .ZN(n9092) );
  OAI21_X1 U10341 ( .B1(n10156), .B2(n10030), .A(n9092), .ZN(n9093) );
  AOI21_X1 U10342 ( .B1(n10096), .B2(n10033), .A(n9093), .ZN(n9094) );
  OAI21_X1 U10343 ( .B1(n11018), .B2(n9095), .A(n9094), .ZN(P2_U3217) );
  NAND2_X1 U10344 ( .A1(n9096), .A2(n9097), .ZN(n9100) );
  INV_X1 U10345 ( .A(n9098), .ZN(n9099) );
  AOI21_X1 U10346 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9108) );
  NAND2_X1 U10347 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10852)
         );
  INV_X1 U10348 ( .A(n10852), .ZN(n9105) );
  OAI22_X1 U10349 ( .A1(n10313), .A2(n9103), .B1(n10299), .B2(n9102), .ZN(
        n9104) );
  AOI211_X1 U10350 ( .C1(n10315), .C2(n10594), .A(n9105), .B(n9104), .ZN(n9107) );
  NAND2_X1 U10351 ( .A1(n9141), .A2(n10289), .ZN(n9106) );
  OAI211_X1 U10352 ( .C1(n9108), .C2(n10292), .A(n9107), .B(n9106), .ZN(
        P1_U3215) );
  INV_X1 U10353 ( .A(n9109), .ZN(n9114) );
  OAI222_X1 U10354 ( .A1(n10696), .A2(n9111), .B1(n9271), .B2(n9114), .C1(
        n9110), .C2(P1_U3086), .ZN(P1_U3329) );
  INV_X1 U10355 ( .A(n9112), .ZN(n9115) );
  OAI222_X1 U10356 ( .A1(P2_U3151), .A2(n9115), .B1(n10175), .B2(n9114), .C1(
        n9113), .C2(n10173), .ZN(P2_U3269) );
  AOI21_X1 U10357 ( .B1(n11186), .B2(n9117), .A(n9116), .ZN(n9132) );
  AOI21_X1 U10358 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(n9128) );
  NAND2_X1 U10359 ( .A1(n10959), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9127) );
  OAI21_X1 U10360 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9125) );
  NOR2_X1 U10361 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9124), .ZN(n9166) );
  AOI21_X1 U10362 ( .B1(n9125), .B2(n5272), .A(n9166), .ZN(n9126) );
  OAI211_X1 U10363 ( .C1(n9128), .C2(n10972), .A(n9127), .B(n9126), .ZN(n9129)
         );
  AOI21_X1 U10364 ( .B1(n9130), .B2(n9881), .A(n9129), .ZN(n9131) );
  OAI21_X1 U10365 ( .B1(n9132), .B2(n10967), .A(n9131), .ZN(P2_U3195) );
  INV_X1 U10366 ( .A(n10285), .ZN(n9137) );
  XNOR2_X1 U10367 ( .A(n9133), .B(n9146), .ZN(n9134) );
  NAND2_X1 U10368 ( .A1(n9134), .A2(n11232), .ZN(n9136) );
  AOI22_X1 U10369 ( .A1(n9222), .A2(n11237), .B1(n11236), .B2(n10595), .ZN(
        n9135) );
  NAND2_X1 U10370 ( .A1(n9136), .A2(n9135), .ZN(n11272) );
  AOI21_X1 U10371 ( .B1(n11243), .B2(n9137), .A(n11272), .ZN(n9151) );
  AND2_X1 U10372 ( .A1(n5219), .A2(n9138), .ZN(n9139) );
  OR2_X1 U10373 ( .A1(n9141), .A2(n11210), .ZN(n9142) );
  NAND2_X1 U10374 ( .A1(n7337), .A2(n10594), .ZN(n9144) );
  NAND2_X1 U10375 ( .A1(n11202), .A2(n9144), .ZN(n10587) );
  NAND2_X1 U10376 ( .A1(n10587), .A2(n10592), .ZN(n10586) );
  NAND2_X1 U10377 ( .A1(n10602), .A2(n11235), .ZN(n9145) );
  NAND2_X1 U10378 ( .A1(n10586), .A2(n9145), .ZN(n11247) );
  NOR2_X1 U10379 ( .A1(n9147), .A2(n9146), .ZN(n9179) );
  AOI21_X1 U10380 ( .B1(n9147), .B2(n9146), .A(n9179), .ZN(n11274) );
  INV_X1 U10381 ( .A(n10290), .ZN(n11270) );
  OAI211_X1 U10382 ( .C1(n11270), .C2(n5232), .A(n11250), .B(n9186), .ZN(
        n11268) );
  AOI22_X1 U10383 ( .A1(n10290), .A2(n11245), .B1(n11258), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9148) );
  OAI21_X1 U10384 ( .B1(n11268), .B2(n11253), .A(n9148), .ZN(n9149) );
  AOI21_X1 U10385 ( .B1(n11274), .B2(n11218), .A(n9149), .ZN(n9150) );
  OAI21_X1 U10386 ( .B1(n11258), .B2(n9151), .A(n9150), .ZN(P1_U3275) );
  INV_X1 U10387 ( .A(n9152), .ZN(n11180) );
  XNOR2_X1 U10388 ( .A(n9152), .B(n9373), .ZN(n9154) );
  NAND2_X1 U10389 ( .A1(n9154), .A2(n9153), .ZN(n9191) );
  INV_X1 U10390 ( .A(n9154), .ZN(n9155) );
  NAND2_X1 U10391 ( .A1(n9155), .A2(n9796), .ZN(n9156) );
  NAND2_X1 U10392 ( .A1(n9191), .A2(n9156), .ZN(n9162) );
  INV_X1 U10393 ( .A(n9157), .ZN(n9158) );
  AND2_X1 U10394 ( .A1(n9158), .A2(n9797), .ZN(n9161) );
  NOR2_X1 U10395 ( .A1(n9162), .A2(n9161), .ZN(n9159) );
  INV_X1 U10396 ( .A(n9161), .ZN(n9164) );
  INV_X1 U10397 ( .A(n9162), .ZN(n9163) );
  AOI21_X1 U10398 ( .B1(n9160), .B2(n9164), .A(n9163), .ZN(n9165) );
  OAI21_X1 U10399 ( .B1(n5230), .B2(n9165), .A(n9773), .ZN(n9171) );
  AOI21_X1 U10400 ( .B1(n9776), .B2(n9797), .A(n9166), .ZN(n9167) );
  OAI21_X1 U10401 ( .B1(n9505), .B2(n9754), .A(n9167), .ZN(n9168) );
  AOI21_X1 U10402 ( .B1(n9169), .B2(n9766), .A(n9168), .ZN(n9170) );
  OAI211_X1 U10403 ( .C1(n11180), .C2(n9784), .A(n9171), .B(n9170), .ZN(
        P2_U3174) );
  NAND2_X1 U10404 ( .A1(n9175), .A2(n9214), .ZN(n9173) );
  OAI211_X1 U10405 ( .C1(n10173), .C2(n9174), .A(n9173), .B(n9172), .ZN(
        P2_U3268) );
  INV_X1 U10406 ( .A(n9175), .ZN(n9178) );
  OAI222_X1 U10407 ( .A1(n9271), .A2(n9178), .B1(n9177), .B2(P1_U3086), .C1(
        n9176), .C2(n10696), .ZN(P1_U3328) );
  XNOR2_X1 U10408 ( .A(n9225), .B(n9180), .ZN(n10672) );
  AOI21_X1 U10409 ( .B1(n9183), .B2(n9182), .A(n9181), .ZN(n9184) );
  OAI222_X1 U10410 ( .A1(n10505), .A2(n10199), .B1(n10507), .B2(n10241), .C1(
        n10503), .C2(n9184), .ZN(n10667) );
  INV_X1 U10411 ( .A(n10669), .ZN(n9223) );
  INV_X1 U10412 ( .A(n9226), .ZN(n9185) );
  AOI211_X1 U10413 ( .C1(n10669), .C2(n9186), .A(n10609), .B(n9185), .ZN(
        n10668) );
  NAND2_X1 U10414 ( .A1(n10668), .A2(n10560), .ZN(n9188) );
  AOI22_X1 U10415 ( .A1(n11244), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10189), 
        .B2(n11243), .ZN(n9187) );
  OAI211_X1 U10416 ( .C1(n9223), .C2(n10534), .A(n9188), .B(n9187), .ZN(n9189)
         );
  AOI21_X1 U10417 ( .B1(n10667), .B2(n10600), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10418 ( .B1(n10672), .B2(n11254), .A(n9190), .ZN(P1_U3274) );
  XNOR2_X1 U10419 ( .A(n10164), .B(n9373), .ZN(n9200) );
  XNOR2_X1 U10420 ( .A(n9200), .B(n9795), .ZN(n9192) );
  NOR3_X1 U10421 ( .A1(n5230), .A2(n5682), .A3(n9192), .ZN(n9194) );
  INV_X1 U10422 ( .A(n9204), .ZN(n9193) );
  OAI21_X1 U10423 ( .B1(n9194), .B2(n9193), .A(n9773), .ZN(n9199) );
  AND2_X1 U10424 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9813) );
  AOI21_X1 U10425 ( .B1(n9776), .B2(n9796), .A(n9813), .ZN(n9195) );
  OAI21_X1 U10426 ( .B1(n9244), .B2(n9754), .A(n9195), .ZN(n9196) );
  AOI21_X1 U10427 ( .B1(n9197), .B2(n9766), .A(n9196), .ZN(n9198) );
  OAI211_X1 U10428 ( .C1(n9502), .C2(n9784), .A(n9199), .B(n9198), .ZN(
        P2_U3155) );
  NAND2_X1 U10429 ( .A1(n9200), .A2(n9505), .ZN(n9202) );
  AND2_X1 U10430 ( .A1(n9204), .A2(n9202), .ZN(n9206) );
  XNOR2_X1 U10431 ( .A(n9201), .B(n9373), .ZN(n9236) );
  XNOR2_X1 U10432 ( .A(n9236), .B(n9794), .ZN(n9205) );
  AND2_X1 U10433 ( .A1(n9205), .A2(n9202), .ZN(n9203) );
  NAND2_X1 U10434 ( .A1(n9204), .A2(n9203), .ZN(n9239) );
  OAI211_X1 U10435 ( .C1(n9206), .C2(n9205), .A(n9239), .B(n9773), .ZN(n9213)
         );
  NOR2_X1 U10436 ( .A1(n9754), .A2(n10019), .ZN(n9210) );
  NOR2_X1 U10437 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9207), .ZN(n9833) );
  INV_X1 U10438 ( .A(n9833), .ZN(n9208) );
  OAI21_X1 U10439 ( .B1(n9763), .B2(n9505), .A(n9208), .ZN(n9209) );
  AOI211_X1 U10440 ( .C1(n9211), .C2(n9766), .A(n9210), .B(n9209), .ZN(n9212)
         );
  OAI211_X1 U10441 ( .C1(n10161), .C2(n9784), .A(n9213), .B(n9212), .ZN(
        P2_U3181) );
  NAND2_X1 U10442 ( .A1(n9218), .A2(n9214), .ZN(n9216) );
  OAI211_X1 U10443 ( .C1(n10173), .C2(n9217), .A(n9216), .B(n9215), .ZN(
        P2_U3267) );
  INV_X1 U10444 ( .A(n9218), .ZN(n9221) );
  OAI222_X1 U10445 ( .A1(n9271), .A2(n9221), .B1(n9220), .B2(P1_U3086), .C1(
        n9219), .C2(n10696), .ZN(P1_U3327) );
  NOR2_X1 U10446 ( .A1(n10669), .A2(n9222), .ZN(n9224) );
  XOR2_X1 U10447 ( .A(n9306), .B(n9307), .Z(n10666) );
  NAND2_X1 U10448 ( .A1(n10664), .A2(n9226), .ZN(n9227) );
  NAND2_X1 U10449 ( .A1(n9227), .A2(n11250), .ZN(n9228) );
  NOR2_X1 U10450 ( .A1(n10577), .A2(n9228), .ZN(n10663) );
  OAI22_X1 U10451 ( .A1(n10600), .A2(n9229), .B1(n10258), .B2(n10580), .ZN(
        n9232) );
  INV_X1 U10452 ( .A(n10664), .ZN(n9230) );
  NOR2_X1 U10453 ( .A1(n9230), .A2(n10534), .ZN(n9231) );
  AOI211_X1 U10454 ( .C1(n10663), .C2(n10560), .A(n9232), .B(n9231), .ZN(n9235) );
  XNOR2_X1 U10455 ( .A(n9290), .B(n9306), .ZN(n9233) );
  OAI222_X1 U10456 ( .A1(n10505), .A2(n10271), .B1(n10507), .B2(n10284), .C1(
        n9233), .C2(n10503), .ZN(n10662) );
  NAND2_X1 U10457 ( .A1(n10662), .A2(n10600), .ZN(n9234) );
  OAI211_X1 U10458 ( .C1(n10666), .C2(n11254), .A(n9235), .B(n9234), .ZN(
        P1_U3273) );
  INV_X1 U10459 ( .A(n9236), .ZN(n9237) );
  NAND2_X1 U10460 ( .A1(n9237), .A2(n9794), .ZN(n9238) );
  NAND2_X1 U10461 ( .A1(n9239), .A2(n9238), .ZN(n9332) );
  XNOR2_X1 U10462 ( .A(n9246), .B(n9373), .ZN(n9333) );
  XNOR2_X1 U10463 ( .A(n9333), .B(n9793), .ZN(n9331) );
  XNOR2_X1 U10464 ( .A(n9332), .B(n9331), .ZN(n9248) );
  NAND2_X1 U10465 ( .A1(n9766), .A2(n9240), .ZN(n9243) );
  NOR2_X1 U10466 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9241), .ZN(n9847) );
  AOI21_X1 U10467 ( .B1(n9781), .B2(n10002), .A(n9847), .ZN(n9242) );
  OAI211_X1 U10468 ( .C1(n9244), .C2(n9763), .A(n9243), .B(n9242), .ZN(n9245)
         );
  AOI21_X1 U10469 ( .B1(n9246), .B2(n9731), .A(n9245), .ZN(n9247) );
  OAI21_X1 U10470 ( .B1(n9248), .B2(n9748), .A(n9247), .ZN(P2_U3166) );
  NAND2_X1 U10471 ( .A1(n9253), .A2(n9249), .ZN(n9250) );
  NAND2_X1 U10472 ( .A1(n9251), .A2(n9250), .ZN(n10990) );
  NAND2_X1 U10473 ( .A1(n10990), .A2(n11077), .ZN(n9258) );
  OAI21_X1 U10474 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  NAND2_X1 U10475 ( .A1(n9255), .A2(n11232), .ZN(n9257) );
  AOI22_X1 U10476 ( .A1(n11236), .A2(n10338), .B1(n10336), .B2(n11237), .ZN(
        n9256) );
  NAND3_X1 U10477 ( .A1(n9258), .A2(n9257), .A3(n9256), .ZN(n10988) );
  MUX2_X1 U10478 ( .A(n10988), .B(P1_REG2_REG_1__SCAN_IN), .S(n11258), .Z(
        n9269) );
  INV_X1 U10479 ( .A(n10990), .ZN(n9266) );
  NAND2_X1 U10480 ( .A1(n11245), .A2(n9260), .ZN(n9265) );
  NAND2_X1 U10481 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U10482 ( .A1(n9261), .A2(n11250), .ZN(n9262) );
  NOR2_X1 U10483 ( .A1(n9263), .A2(n9262), .ZN(n10985) );
  AOI22_X1 U10484 ( .A1(n10560), .A2(n10985), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n11243), .ZN(n9264) );
  OAI211_X1 U10485 ( .C1(n9267), .C2(n9266), .A(n9265), .B(n9264), .ZN(n9268)
         );
  OR2_X1 U10486 ( .A1(n9269), .A2(n9268), .ZN(P1_U3292) );
  INV_X1 U10487 ( .A(n9412), .ZN(n9274) );
  OAI222_X1 U10488 ( .A1(n10696), .A2(n9272), .B1(n9271), .B2(n9274), .C1(
        P1_U3086), .C2(n9270), .ZN(P1_U3325) );
  OAI222_X1 U10489 ( .A1(n9273), .A2(P2_U3151), .B1(n9275), .B2(n9274), .C1(
        n9413), .C2(n10173), .ZN(P2_U3265) );
  INV_X1 U10490 ( .A(n9276), .ZN(n9459) );
  NAND2_X1 U10491 ( .A1(n9457), .A2(n9459), .ZN(n9593) );
  XOR2_X1 U10492 ( .A(n9593), .B(n9277), .Z(n11049) );
  XNOR2_X1 U10493 ( .A(n9278), .B(n9593), .ZN(n9279) );
  OAI222_X1 U10494 ( .A1(n11003), .A2(n9281), .B1(n11001), .B2(n9280), .C1(
        n9279), .C2(n11000), .ZN(n11051) );
  NAND2_X1 U10495 ( .A1(n11051), .A2(n11015), .ZN(n9288) );
  INV_X1 U10496 ( .A(n9282), .ZN(n9283) );
  OAI22_X1 U10497 ( .A1(n11015), .A2(n9284), .B1(n9283), .B2(n11010), .ZN(
        n9285) );
  AOI21_X1 U10498 ( .B1(n10015), .B2(n9286), .A(n9285), .ZN(n9287) );
  OAI211_X1 U10499 ( .C1(n11049), .C2(n10012), .A(n9288), .B(n9287), .ZN(
        P2_U3228) );
  OAI21_X1 U10500 ( .B1(n10569), .B2(n9291), .A(n10575), .ZN(n10567) );
  NAND2_X1 U10501 ( .A1(n10567), .A2(n9292), .ZN(n10548) );
  INV_X1 U10502 ( .A(n9296), .ZN(n9297) );
  XNOR2_X1 U10503 ( .A(n9300), .B(n9313), .ZN(n9304) );
  INV_X1 U10504 ( .A(n10471), .ZN(n10322) );
  AOI21_X1 U10505 ( .B1(n9301), .B2(P1_B_REG_SCAN_IN), .A(n10505), .ZN(n9327)
         );
  OAI21_X2 U10506 ( .B1(n9307), .B2(n9306), .A(n9305), .ZN(n10574) );
  NAND2_X1 U10507 ( .A1(n10528), .A2(n5736), .ZN(n9309) );
  NAND2_X1 U10508 ( .A1(n9309), .A2(n9308), .ZN(n10517) );
  INV_X1 U10509 ( .A(n10517), .ZN(n9310) );
  NOR2_X1 U10510 ( .A1(n10637), .A2(n10513), .ZN(n9312) );
  INV_X1 U10511 ( .A(n10637), .ZN(n10495) );
  AOI22_X1 U10512 ( .A1(n10460), .A2(n10467), .B1(n10482), .B2(n10462), .ZN(
        n10456) );
  NAND2_X1 U10513 ( .A1(n10456), .A2(n10455), .ZN(n10454) );
  OAI21_X1 U10514 ( .B1(n10449), .B2(n10471), .A(n10454), .ZN(n9314) );
  NAND2_X1 U10515 ( .A1(n11244), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9315) );
  OAI21_X1 U10516 ( .B1(n10580), .B2(n9316), .A(n9315), .ZN(n9317) );
  AOI21_X1 U10517 ( .B1(n10614), .B2(n11245), .A(n9317), .ZN(n9321) );
  NAND2_X1 U10518 ( .A1(n10495), .A2(n10520), .ZN(n10492) );
  AOI21_X1 U10519 ( .B1(n10614), .B2(n10448), .A(n10609), .ZN(n9319) );
  AND2_X1 U10520 ( .A1(n9319), .A2(n10438), .ZN(n10613) );
  NAND2_X1 U10521 ( .A1(n10613), .A2(n10560), .ZN(n9320) );
  OAI211_X1 U10522 ( .C1(n10617), .C2(n11254), .A(n9321), .B(n9320), .ZN(n9322) );
  INV_X1 U10523 ( .A(n9322), .ZN(n9323) );
  OAI21_X1 U10524 ( .B1(n10615), .B2(n11244), .A(n9323), .ZN(P1_U3356) );
  XNOR2_X1 U10525 ( .A(n9325), .B(n9324), .ZN(n10610) );
  NOR2_X1 U10526 ( .A1(n10600), .A2(n9326), .ZN(n9328) );
  NAND2_X1 U10527 ( .A1(n10319), .A2(n9327), .ZN(n10611) );
  NOR2_X1 U10528 ( .A1(n11244), .A2(n10611), .ZN(n10441) );
  AOI211_X1 U10529 ( .C1(n10607), .C2(n11245), .A(n9328), .B(n10441), .ZN(
        n9329) );
  OAI21_X1 U10530 ( .B1(n10610), .B2(n9330), .A(n9329), .ZN(P1_U3263) );
  INV_X1 U10531 ( .A(n9333), .ZN(n9334) );
  NAND2_X1 U10532 ( .A1(n9334), .A2(n9793), .ZN(n9335) );
  XNOR2_X1 U10533 ( .A(n9995), .B(n9373), .ZN(n9692) );
  XNOR2_X1 U10534 ( .A(n10151), .B(n9355), .ZN(n9687) );
  NAND2_X1 U10535 ( .A1(n9687), .A2(n10002), .ZN(n9336) );
  XNOR2_X1 U10536 ( .A(n10086), .B(n9355), .ZN(n9690) );
  NAND2_X1 U10537 ( .A1(n9690), .A2(n9791), .ZN(n9691) );
  INV_X1 U10538 ( .A(n9687), .ZN(n9337) );
  NAND3_X1 U10539 ( .A1(n9337), .A2(n9764), .A3(n10020), .ZN(n9341) );
  NAND2_X1 U10540 ( .A1(n9337), .A2(n9764), .ZN(n9688) );
  NAND2_X1 U10541 ( .A1(n9688), .A2(n9791), .ZN(n9339) );
  INV_X1 U10542 ( .A(n9690), .ZN(n9338) );
  NAND2_X1 U10543 ( .A1(n9339), .A2(n9338), .ZN(n9340) );
  NAND3_X1 U10544 ( .A1(n9692), .A2(n9341), .A3(n9340), .ZN(n9342) );
  OAI21_X1 U10545 ( .B1(n9692), .B2(n9744), .A(n9342), .ZN(n9343) );
  NAND2_X1 U10546 ( .A1(n9344), .A2(n9343), .ZN(n9740) );
  XNOR2_X1 U10547 ( .A(n9539), .B(n9373), .ZN(n9345) );
  NAND2_X1 U10548 ( .A1(n9345), .A2(n9709), .ZN(n9701) );
  INV_X1 U10549 ( .A(n9345), .ZN(n9346) );
  NAND2_X1 U10550 ( .A1(n9346), .A2(n9988), .ZN(n9347) );
  AND2_X1 U10551 ( .A1(n9701), .A2(n9347), .ZN(n9741) );
  NAND2_X1 U10552 ( .A1(n9700), .A2(n9701), .ZN(n9348) );
  XNOR2_X1 U10553 ( .A(n10072), .B(n9373), .ZN(n9349) );
  XNOR2_X1 U10554 ( .A(n9349), .B(n9978), .ZN(n9702) );
  NAND2_X1 U10555 ( .A1(n9349), .A2(n9955), .ZN(n9350) );
  XNOR2_X1 U10556 ( .A(n9351), .B(n9373), .ZN(n9352) );
  XNOR2_X1 U10557 ( .A(n9352), .B(n9943), .ZN(n9749) );
  INV_X1 U10558 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U10559 ( .A1(n9353), .A2(n5319), .ZN(n9354) );
  NAND2_X1 U10560 ( .A1(n9751), .A2(n9354), .ZN(n9358) );
  XNOR2_X1 U10561 ( .A(n9553), .B(n9355), .ZN(n9357) );
  XNOR2_X1 U10562 ( .A(n9432), .B(n9373), .ZN(n9361) );
  NAND2_X1 U10563 ( .A1(n9361), .A2(n9944), .ZN(n9364) );
  INV_X1 U10564 ( .A(n9361), .ZN(n9362) );
  NAND2_X1 U10565 ( .A1(n9362), .A2(n9789), .ZN(n9363) );
  NAND2_X1 U10566 ( .A1(n9364), .A2(n9363), .ZN(n9734) );
  AOI21_X2 U10567 ( .B1(n9680), .B2(n9360), .A(n9734), .ZN(n9714) );
  INV_X1 U10568 ( .A(n9364), .ZN(n9716) );
  XNOR2_X1 U10569 ( .A(n10126), .B(n9373), .ZN(n9368) );
  XNOR2_X1 U10570 ( .A(n9368), .B(n9932), .ZN(n9715) );
  NAND2_X1 U10571 ( .A1(n9365), .A2(n9370), .ZN(n9613) );
  INV_X1 U10572 ( .A(n9613), .ZN(n9909) );
  NOR2_X1 U10573 ( .A1(n9403), .A2(n9366), .ZN(n9367) );
  MUX2_X1 U10574 ( .A(n9909), .B(n9367), .S(n9373), .Z(n9774) );
  INV_X1 U10575 ( .A(n9368), .ZN(n9369) );
  NAND2_X1 U10576 ( .A1(n9369), .A2(n9932), .ZN(n9770) );
  MUX2_X1 U10577 ( .A(n9370), .B(n9567), .S(n9373), .Z(n9371) );
  XNOR2_X1 U10578 ( .A(n10118), .B(n9373), .ZN(n9372) );
  XNOR2_X1 U10579 ( .A(n9372), .B(n9908), .ZN(n9672) );
  INV_X1 U10580 ( .A(n9374), .ZN(n9395) );
  INV_X1 U10581 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9375) );
  OAI22_X1 U10582 ( .A1(n9395), .A2(n9779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9375), .ZN(n9377) );
  OAI22_X1 U10583 ( .A1(n9419), .A2(n9754), .B1(n9908), .B2(n9763), .ZN(n9376)
         );
  AOI211_X1 U10584 ( .C1(n9657), .C2(n9731), .A(n9377), .B(n9376), .ZN(n9378)
         );
  OAI21_X1 U10585 ( .B1(n9379), .B2(n9748), .A(n9378), .ZN(P2_U3160) );
  INV_X1 U10586 ( .A(n9380), .ZN(n9381) );
  NOR3_X1 U10587 ( .A1(n9383), .A2(n9382), .A3(n9381), .ZN(n9386) );
  OAI21_X1 U10588 ( .B1(n9386), .B2(n9385), .A(n10308), .ZN(n9392) );
  OAI22_X1 U10589 ( .A1(n10313), .A2(n9388), .B1(n10299), .B2(n9387), .ZN(
        n9389) );
  AOI211_X1 U10590 ( .C1(n10315), .C2(n10328), .A(n9390), .B(n9389), .ZN(n9391) );
  OAI211_X1 U10591 ( .C1(n9393), .C2(n10318), .A(n9392), .B(n9391), .ZN(
        P1_U3231) );
  OAI22_X1 U10592 ( .A1(n9395), .A2(n11010), .B1(n11015), .B2(n9394), .ZN(
        n9398) );
  NOR2_X1 U10593 ( .A1(n9396), .A2(n10012), .ZN(n9397) );
  AOI211_X1 U10594 ( .C1(n10015), .C2(n9657), .A(n9398), .B(n9397), .ZN(n9399)
         );
  OAI21_X1 U10595 ( .B1(n9400), .B2(n11018), .A(n9399), .ZN(P2_U3205) );
  NOR2_X1 U10596 ( .A1(n9404), .A2(n9431), .ZN(n9406) );
  INV_X1 U10597 ( .A(n9657), .ZN(n9405) );
  NAND2_X1 U10598 ( .A1(n10172), .A2(n6172), .ZN(n9408) );
  OR2_X1 U10599 ( .A1(n6104), .A2(n10174), .ZN(n9407) );
  NAND2_X1 U10600 ( .A1(n9408), .A2(n9407), .ZN(n10038) );
  OR2_X1 U10601 ( .A1(n10038), .A2(n9419), .ZN(n9576) );
  NAND2_X1 U10602 ( .A1(n10694), .A2(n6172), .ZN(n9411) );
  INV_X1 U10603 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9409) );
  OR2_X1 U10604 ( .A1(n6104), .A2(n9409), .ZN(n9410) );
  OR2_X1 U10605 ( .A1(n9424), .A2(n9887), .ZN(n9417) );
  NAND2_X1 U10606 ( .A1(n9412), .A2(n6172), .ZN(n9415) );
  OR2_X1 U10607 ( .A1(n6104), .A2(n9413), .ZN(n9414) );
  NAND2_X1 U10608 ( .A1(n9415), .A2(n9414), .ZN(n9423) );
  NAND2_X1 U10609 ( .A1(n9423), .A2(n9663), .ZN(n9416) );
  AND2_X1 U10610 ( .A1(n9417), .A2(n9416), .ZN(n9586) );
  NAND2_X1 U10611 ( .A1(n9418), .A2(n9423), .ZN(n9420) );
  NAND2_X1 U10612 ( .A1(n9424), .A2(n9887), .ZN(n9584) );
  OR2_X1 U10613 ( .A1(n9423), .A2(n9663), .ZN(n9578) );
  AND2_X1 U10614 ( .A1(n9584), .A2(n9578), .ZN(n9587) );
  NOR2_X1 U10615 ( .A1(n9587), .A2(n9418), .ZN(n9427) );
  NAND2_X1 U10616 ( .A1(n9429), .A2(n9428), .ZN(n9620) );
  AND2_X1 U10617 ( .A1(n9576), .A2(n9580), .ZN(n9430) );
  NAND2_X1 U10618 ( .A1(n9578), .A2(n9430), .ZN(n9582) );
  OAI22_X1 U10619 ( .A1(n9582), .A2(n9405), .B1(n9580), .B2(n9893), .ZN(n9575)
         );
  INV_X1 U10620 ( .A(n9431), .ZN(n9571) );
  XNOR2_X1 U10621 ( .A(n9432), .B(n9789), .ZN(n9929) );
  NAND2_X1 U10622 ( .A1(n9442), .A2(n7485), .ZN(n9434) );
  NAND2_X1 U10623 ( .A1(n9434), .A2(n9433), .ZN(n9436) );
  NAND2_X1 U10624 ( .A1(n9436), .A2(n9435), .ZN(n9437) );
  NAND2_X1 U10625 ( .A1(n9437), .A2(n6441), .ZN(n9441) );
  NAND2_X1 U10626 ( .A1(n9452), .A2(n9439), .ZN(n9440) );
  AOI21_X1 U10627 ( .B1(n9441), .B2(n10996), .A(n9440), .ZN(n9449) );
  INV_X1 U10628 ( .A(n9442), .ZN(n9443) );
  NAND2_X1 U10629 ( .A1(n6441), .A2(n9443), .ZN(n9444) );
  NAND2_X1 U10630 ( .A1(n9444), .A2(n9435), .ZN(n9447) );
  NAND2_X1 U10631 ( .A1(n9456), .A2(n9445), .ZN(n9446) );
  AOI21_X1 U10632 ( .B1(n10996), .B2(n9447), .A(n9446), .ZN(n9448) );
  MUX2_X1 U10633 ( .A(n9449), .B(n9448), .S(n9580), .Z(n9450) );
  INV_X1 U10634 ( .A(n9450), .ZN(n9451) );
  NAND2_X1 U10635 ( .A1(n9451), .A2(n9453), .ZN(n9458) );
  NAND2_X1 U10636 ( .A1(n9452), .A2(n5162), .ZN(n9454) );
  OAI211_X1 U10637 ( .C1(n9458), .C2(n9454), .A(n9459), .B(n9453), .ZN(n9455)
         );
  NAND3_X1 U10638 ( .A1(n9455), .A2(n9465), .A3(n9457), .ZN(n9462) );
  OAI211_X1 U10639 ( .C1(n9458), .C2(n6444), .A(n9457), .B(n5162), .ZN(n9460)
         );
  NAND3_X1 U10640 ( .A1(n9460), .A2(n9459), .A3(n9464), .ZN(n9461) );
  MUX2_X1 U10641 ( .A(n9462), .B(n9461), .S(n9574), .Z(n9469) );
  MUX2_X1 U10642 ( .A(n9474), .B(n9463), .S(n9580), .Z(n9470) );
  AND2_X1 U10643 ( .A1(n9470), .A2(n9475), .ZN(n9482) );
  INV_X1 U10644 ( .A(n9464), .ZN(n9466) );
  MUX2_X1 U10645 ( .A(n9466), .B(n6447), .S(n9574), .Z(n9467) );
  NOR2_X1 U10646 ( .A1(n9595), .A2(n9467), .ZN(n9468) );
  NAND3_X1 U10647 ( .A1(n9469), .A2(n9482), .A3(n9468), .ZN(n9480) );
  INV_X1 U10648 ( .A(n9470), .ZN(n9477) );
  NAND2_X1 U10649 ( .A1(n9472), .A2(n9471), .ZN(n9473) );
  AND2_X1 U10650 ( .A1(n9474), .A2(n9473), .ZN(n9476) );
  OAI211_X1 U10651 ( .C1(n9477), .C2(n9476), .A(n9487), .B(n9475), .ZN(n9478)
         );
  NAND2_X1 U10652 ( .A1(n9478), .A2(n9580), .ZN(n9479) );
  NAND2_X1 U10653 ( .A1(n9480), .A2(n9479), .ZN(n9489) );
  NAND3_X1 U10654 ( .A1(n9489), .A2(n5220), .A3(n9492), .ZN(n9481) );
  INV_X1 U10655 ( .A(n9482), .ZN(n9486) );
  AND2_X1 U10656 ( .A1(n5166), .A2(n9483), .ZN(n9485) );
  OAI211_X1 U10657 ( .C1(n9486), .C2(n9485), .A(n5220), .B(n9484), .ZN(n9488)
         );
  OAI21_X1 U10658 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9493) );
  INV_X1 U10659 ( .A(n9490), .ZN(n9491) );
  NOR2_X1 U10660 ( .A1(n11157), .A2(n9495), .ZN(n9496) );
  MUX2_X1 U10661 ( .A(n5553), .B(n9496), .S(n9580), .Z(n9497) );
  NOR2_X1 U10662 ( .A1(n9604), .A2(n9497), .ZN(n9498) );
  MUX2_X1 U10663 ( .A(n9500), .B(n9499), .S(n9574), .Z(n9501) );
  NAND2_X1 U10664 ( .A1(n9513), .A2(n9605), .ZN(n9506) );
  AND2_X1 U10665 ( .A1(n9507), .A2(n9502), .ZN(n9504) );
  INV_X1 U10666 ( .A(n9509), .ZN(n9503) );
  AOI21_X1 U10667 ( .B1(n9506), .B2(n9504), .A(n9503), .ZN(n9512) );
  NAND2_X1 U10668 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  NAND2_X1 U10669 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  NAND2_X1 U10670 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  INV_X1 U10671 ( .A(n9513), .ZN(n9518) );
  NOR2_X1 U10672 ( .A1(n9515), .A2(n9514), .ZN(n9517) );
  AOI21_X1 U10673 ( .B1(n9518), .B2(n9517), .A(n9516), .ZN(n9523) );
  INV_X1 U10674 ( .A(n9520), .ZN(n9521) );
  MUX2_X1 U10675 ( .A(n5568), .B(n9521), .S(n9574), .Z(n9522) );
  MUX2_X1 U10676 ( .A(n10002), .B(n10151), .S(n9580), .Z(n9528) );
  NAND2_X1 U10677 ( .A1(n9531), .A2(n10002), .ZN(n9525) );
  NAND2_X1 U10678 ( .A1(n9530), .A2(n10151), .ZN(n9524) );
  MUX2_X1 U10679 ( .A(n9525), .B(n9524), .S(n9574), .Z(n9526) );
  AOI21_X1 U10680 ( .B1(n9527), .B2(n9528), .A(n9526), .ZN(n9538) );
  INV_X1 U10681 ( .A(n9528), .ZN(n9529) );
  MUX2_X1 U10682 ( .A(n9531), .B(n9530), .S(n9580), .Z(n9532) );
  NAND3_X1 U10683 ( .A1(n9533), .A2(n9995), .A3(n9532), .ZN(n9537) );
  MUX2_X1 U10684 ( .A(n9535), .B(n9534), .S(n9574), .Z(n9536) );
  OAI211_X1 U10685 ( .C1(n9538), .C2(n9537), .A(n9981), .B(n9536), .ZN(n9545)
         );
  NAND2_X1 U10686 ( .A1(n9539), .A2(n9574), .ZN(n9541) );
  NAND2_X1 U10687 ( .A1(n10143), .A2(n9580), .ZN(n9540) );
  MUX2_X1 U10688 ( .A(n9541), .B(n9540), .S(n9988), .Z(n9544) );
  INV_X1 U10689 ( .A(n10072), .ZN(n9713) );
  MUX2_X1 U10690 ( .A(n9955), .B(n9713), .S(n9580), .Z(n9546) );
  NAND2_X1 U10691 ( .A1(n9546), .A2(n9542), .ZN(n9543) );
  NAND3_X1 U10692 ( .A1(n9545), .A2(n9544), .A3(n9543), .ZN(n9549) );
  INV_X1 U10693 ( .A(n9546), .ZN(n9548) );
  MUX2_X1 U10694 ( .A(n9551), .B(n9550), .S(n9574), .Z(n9552) );
  AND2_X1 U10695 ( .A1(n9553), .A2(n9954), .ZN(n9556) );
  INV_X1 U10696 ( .A(n9554), .ZN(n9555) );
  MUX2_X1 U10697 ( .A(n9556), .B(n9555), .S(n9574), .Z(n9557) );
  INV_X1 U10698 ( .A(n9557), .ZN(n9558) );
  MUX2_X1 U10699 ( .A(n9560), .B(n9559), .S(n9574), .Z(n9561) );
  MUX2_X1 U10700 ( .A(n9563), .B(n9562), .S(n9580), .Z(n9564) );
  NAND2_X1 U10701 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  NAND2_X1 U10702 ( .A1(n9566), .A2(n9613), .ZN(n9569) );
  MUX2_X1 U10703 ( .A(n9898), .B(n9567), .S(n9574), .Z(n9568) );
  NAND3_X1 U10704 ( .A1(n9900), .A2(n9569), .A3(n9568), .ZN(n9573) );
  MUX2_X1 U10705 ( .A(n9571), .B(n9570), .S(n9580), .Z(n9572) );
  MUX2_X1 U10706 ( .A(n9785), .B(n9657), .S(n9574), .Z(n9577) );
  NAND2_X1 U10707 ( .A1(n9576), .A2(n5743), .ZN(n9658) );
  INV_X1 U10708 ( .A(n9578), .ZN(n9579) );
  AOI211_X1 U10709 ( .C1(n9581), .C2(n5743), .A(n9580), .B(n9579), .ZN(n9585)
         );
  INV_X1 U10710 ( .A(n9581), .ZN(n9583) );
  INV_X1 U10711 ( .A(n9586), .ZN(n9617) );
  INV_X1 U10712 ( .A(n9587), .ZN(n9616) );
  INV_X1 U10713 ( .A(n9940), .ZN(n9946) );
  INV_X1 U10714 ( .A(n9929), .ZN(n9934) );
  INV_X1 U10715 ( .A(n10010), .ZN(n9609) );
  NOR3_X1 U10716 ( .A1(n9589), .A2(n9588), .A3(n7485), .ZN(n9592) );
  NAND4_X1 U10717 ( .A1(n9592), .A2(n9591), .A3(n10996), .A4(n9590), .ZN(n9596) );
  NOR4_X1 U10718 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9599)
         );
  NAND4_X1 U10719 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9601)
         );
  NOR4_X1 U10720 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n9606)
         );
  NAND4_X1 U10721 ( .A1(n6452), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9608)
         );
  NOR4_X1 U10722 ( .A1(n9610), .A2(n10024), .A3(n9609), .A4(n9608), .ZN(n9611)
         );
  NAND4_X1 U10723 ( .A1(n9956), .A2(n9611), .A3(n9971), .A4(n9981), .ZN(n9612)
         );
  NOR4_X1 U10724 ( .A1(n9917), .A2(n9946), .A3(n9934), .A4(n9612), .ZN(n9614)
         );
  NAND4_X1 U10725 ( .A1(n9900), .A2(n9614), .A3(n9613), .A4(n9655), .ZN(n9615)
         );
  XNOR2_X1 U10726 ( .A(n9622), .B(n5136), .ZN(n9630) );
  INV_X1 U10727 ( .A(n5872), .ZN(n9624) );
  NAND3_X1 U10728 ( .A1(n9625), .A2(n9624), .A3(n9623), .ZN(n9626) );
  OAI211_X1 U10729 ( .C1(n9627), .C2(n9629), .A(n9626), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9628) );
  OAI21_X1 U10730 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(P2_U3296) );
  NAND2_X1 U10731 ( .A1(n10618), .A2(n7412), .ZN(n9632) );
  OR2_X1 U10732 ( .A1(n10471), .A2(n7255), .ZN(n9631) );
  NAND2_X1 U10733 ( .A1(n9632), .A2(n9631), .ZN(n9634) );
  XNOR2_X1 U10734 ( .A(n9634), .B(n9633), .ZN(n9639) );
  NAND2_X1 U10735 ( .A1(n10618), .A2(n9635), .ZN(n9636) );
  OAI21_X1 U10736 ( .B1(n10471), .B2(n9637), .A(n9636), .ZN(n9638) );
  XNOR2_X1 U10737 ( .A(n9639), .B(n9638), .ZN(n9640) );
  INV_X1 U10738 ( .A(n9640), .ZN(n9645) );
  NAND3_X1 U10739 ( .A1(n9645), .A2(n10308), .A3(n9644), .ZN(n9650) );
  NAND3_X1 U10740 ( .A1(n9651), .A2(n10308), .A3(n9640), .ZN(n9649) );
  AOI22_X1 U10741 ( .A1(n9641), .A2(n10323), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9643) );
  NAND2_X1 U10742 ( .A1(n10315), .A2(n10321), .ZN(n9642) );
  OAI211_X1 U10743 ( .C1(n10451), .C2(n10299), .A(n9643), .B(n9642), .ZN(n9647) );
  NOR3_X1 U10744 ( .A1(n9645), .A2(n10292), .A3(n9644), .ZN(n9646) );
  AOI211_X1 U10745 ( .C1(n10618), .C2(n10289), .A(n9647), .B(n9646), .ZN(n9648) );
  OAI211_X1 U10746 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(
        P1_U3220) );
  NAND2_X1 U10747 ( .A1(n9405), .A2(n9893), .ZN(n9652) );
  XNOR2_X1 U10748 ( .A(n9654), .B(n5339), .ZN(n10042) );
  XNOR2_X1 U10749 ( .A(n9659), .B(n5339), .ZN(n9667) );
  NOR2_X1 U10750 ( .A1(n9667), .A2(n9660), .ZN(n10044) );
  AND2_X1 U10751 ( .A1(n9661), .A2(P2_B_REG_SCAN_IN), .ZN(n9662) );
  OR2_X1 U10752 ( .A1(n11003), .A2(n9662), .ZN(n9886) );
  OAI22_X1 U10753 ( .A1(n9893), .A2(n11001), .B1(n9663), .B2(n9886), .ZN(
        n10043) );
  AOI211_X1 U10754 ( .C1(n10042), .C2(n10041), .A(n10044), .B(n10043), .ZN(
        n9671) );
  NOR2_X1 U10755 ( .A1(n11015), .A2(n9664), .ZN(n9666) );
  NOR2_X1 U10756 ( .A1(n9665), .A2(n11010), .ZN(n9885) );
  AOI211_X1 U10757 ( .C1(n10038), .C2(n10015), .A(n9666), .B(n9885), .ZN(n9670) );
  INV_X1 U10758 ( .A(n9667), .ZN(n10040) );
  NAND2_X1 U10759 ( .A1(n10040), .A2(n9668), .ZN(n9669) );
  OAI211_X1 U10760 ( .C1(n9671), .C2(n11018), .A(n9670), .B(n9669), .ZN(
        P2_U3204) );
  XNOR2_X1 U10761 ( .A(n9673), .B(n9672), .ZN(n9679) );
  NOR2_X1 U10762 ( .A1(n9921), .A2(n9763), .ZN(n9676) );
  AOI22_X1 U10763 ( .A1(n9902), .A2(n9766), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9674) );
  OAI21_X1 U10764 ( .B1(n9893), .B2(n9754), .A(n9674), .ZN(n9675) );
  AOI211_X1 U10765 ( .C1(n9677), .C2(n9731), .A(n9676), .B(n9675), .ZN(n9678)
         );
  OAI21_X1 U10766 ( .B1(n9679), .B2(n9748), .A(n9678), .ZN(P2_U3154) );
  OAI21_X1 U10767 ( .B1(n9954), .B2(n9681), .A(n9680), .ZN(n9682) );
  NAND2_X1 U10768 ( .A1(n9682), .A2(n9773), .ZN(n9686) );
  AOI22_X1 U10769 ( .A1(n9789), .A2(n9781), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9683) );
  OAI21_X1 U10770 ( .B1(n9943), .B2(n9763), .A(n9683), .ZN(n9684) );
  AOI21_X1 U10771 ( .B1(n9947), .B2(n9766), .A(n9684), .ZN(n9685) );
  OAI211_X1 U10772 ( .C1(n10134), .C2(n9784), .A(n9686), .B(n9685), .ZN(
        P2_U3156) );
  XNOR2_X1 U10773 ( .A(n9687), .B(n10002), .ZN(n9726) );
  NOR2_X1 U10774 ( .A1(n9725), .A2(n9726), .ZN(n9724) );
  INV_X1 U10775 ( .A(n9688), .ZN(n9689) );
  NOR2_X1 U10776 ( .A1(n9724), .A2(n9689), .ZN(n9760) );
  XNOR2_X1 U10777 ( .A(n9690), .B(n10020), .ZN(n9759) );
  NAND2_X1 U10778 ( .A1(n9760), .A2(n9759), .ZN(n9758) );
  NAND2_X1 U10779 ( .A1(n9758), .A2(n9691), .ZN(n9693) );
  XNOR2_X1 U10780 ( .A(n9693), .B(n9692), .ZN(n9699) );
  NAND2_X1 U10781 ( .A1(n9766), .A2(n9992), .ZN(n9696) );
  AOI21_X1 U10782 ( .B1(n9781), .B2(n9988), .A(n9694), .ZN(n9695) );
  OAI211_X1 U10783 ( .C1(n10020), .C2(n9763), .A(n9696), .B(n9695), .ZN(n9697)
         );
  AOI21_X1 U10784 ( .B1(n10146), .B2(n9731), .A(n9697), .ZN(n9698) );
  OAI21_X1 U10785 ( .B1(n9699), .B2(n9748), .A(n9698), .ZN(P2_U3159) );
  INV_X1 U10786 ( .A(n9700), .ZN(n9704) );
  INV_X1 U10787 ( .A(n9701), .ZN(n9703) );
  NOR3_X1 U10788 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9707) );
  INV_X1 U10789 ( .A(n9705), .ZN(n9706) );
  OAI21_X1 U10790 ( .B1(n9707), .B2(n9706), .A(n9773), .ZN(n9712) );
  AOI22_X1 U10791 ( .A1(n5319), .A2(n9781), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9708) );
  OAI21_X1 U10792 ( .B1(n9709), .B2(n9763), .A(n9708), .ZN(n9710) );
  AOI21_X1 U10793 ( .B1(n9967), .B2(n9766), .A(n9710), .ZN(n9711) );
  OAI211_X1 U10794 ( .C1(n9713), .C2(n9784), .A(n9712), .B(n9711), .ZN(
        P2_U3163) );
  INV_X1 U10795 ( .A(n9771), .ZN(n9718) );
  NOR3_X1 U10796 ( .A1(n9714), .A2(n9716), .A3(n9715), .ZN(n9717) );
  OAI21_X1 U10797 ( .B1(n9718), .B2(n9717), .A(n9773), .ZN(n9723) );
  INV_X1 U10798 ( .A(n9719), .ZN(n9923) );
  AOI22_X1 U10799 ( .A1(n9789), .A2(n9776), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9720) );
  OAI21_X1 U10800 ( .B1(n9923), .B2(n9779), .A(n9720), .ZN(n9721) );
  AOI21_X1 U10801 ( .B1(n9781), .B2(n9787), .A(n9721), .ZN(n9722) );
  OAI211_X1 U10802 ( .C1(n10126), .C2(n9784), .A(n9723), .B(n9722), .ZN(
        P2_U3165) );
  AOI21_X1 U10803 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9733) );
  NAND2_X1 U10804 ( .A1(n9766), .A2(n10027), .ZN(n9729) );
  NOR2_X1 U10805 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9727), .ZN(n9874) );
  AOI21_X1 U10806 ( .B1(n9781), .B2(n9791), .A(n9874), .ZN(n9728) );
  OAI211_X1 U10807 ( .C1(n10019), .C2(n9763), .A(n9729), .B(n9728), .ZN(n9730)
         );
  AOI21_X1 U10808 ( .B1(n10151), .B2(n9731), .A(n9730), .ZN(n9732) );
  OAI21_X1 U10809 ( .B1(n9733), .B2(n9748), .A(n9732), .ZN(P2_U3168) );
  AND3_X1 U10810 ( .A1(n9680), .A2(n9360), .A3(n9734), .ZN(n9735) );
  OAI21_X1 U10811 ( .B1(n9714), .B2(n9735), .A(n9773), .ZN(n9739) );
  AOI22_X1 U10812 ( .A1(n9788), .A2(n9781), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9736) );
  OAI21_X1 U10813 ( .B1(n9954), .B2(n9763), .A(n9736), .ZN(n9737) );
  AOI21_X1 U10814 ( .B1(n9935), .B2(n9766), .A(n9737), .ZN(n9738) );
  OAI211_X1 U10815 ( .C1(n10130), .C2(n9784), .A(n9739), .B(n9738), .ZN(
        P2_U3169) );
  OAI21_X1 U10816 ( .B1(n9741), .B2(n9740), .A(n9700), .ZN(n9742) );
  NAND2_X1 U10817 ( .A1(n9742), .A2(n9773), .ZN(n9747) );
  AOI22_X1 U10818 ( .A1(n9781), .A2(n9978), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9743) );
  OAI21_X1 U10819 ( .B1(n9744), .B2(n9763), .A(n9743), .ZN(n9745) );
  AOI21_X1 U10820 ( .B1(n9983), .B2(n9766), .A(n9745), .ZN(n9746) );
  OAI211_X1 U10821 ( .C1(n10143), .C2(n9784), .A(n9747), .B(n9746), .ZN(
        P2_U3173) );
  AOI21_X1 U10822 ( .B1(n9750), .B2(n9749), .A(n9748), .ZN(n9752) );
  NAND2_X1 U10823 ( .A1(n9752), .A2(n9751), .ZN(n9757) );
  AOI22_X1 U10824 ( .A1(n9776), .A2(n9978), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9753) );
  OAI21_X1 U10825 ( .B1(n9954), .B2(n9754), .A(n9753), .ZN(n9755) );
  AOI21_X1 U10826 ( .B1(n9958), .B2(n9766), .A(n9755), .ZN(n9756) );
  OAI211_X1 U10827 ( .C1(n10138), .C2(n9784), .A(n9757), .B(n9756), .ZN(
        P2_U3175) );
  INV_X1 U10828 ( .A(n10086), .ZN(n9769) );
  OAI211_X1 U10829 ( .C1(n9760), .C2(n9759), .A(n9758), .B(n9773), .ZN(n9768)
         );
  INV_X1 U10830 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9761) );
  NOR2_X1 U10831 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9761), .ZN(n10958) );
  AOI21_X1 U10832 ( .B1(n9781), .B2(n10004), .A(n10958), .ZN(n9762) );
  OAI21_X1 U10833 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  AOI21_X1 U10834 ( .B1(n10006), .B2(n9766), .A(n9765), .ZN(n9767) );
  OAI211_X1 U10835 ( .C1(n9769), .C2(n9784), .A(n9768), .B(n9767), .ZN(
        P2_U3178) );
  AND2_X1 U10836 ( .A1(n9771), .A2(n9770), .ZN(n9775) );
  OAI211_X1 U10837 ( .C1(n9775), .C2(n9774), .A(n9773), .B(n9772), .ZN(n9783)
         );
  INV_X1 U10838 ( .A(n9911), .ZN(n9778) );
  AOI22_X1 U10839 ( .A1(n9788), .A2(n9776), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9777) );
  OAI21_X1 U10840 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9780) );
  AOI21_X1 U10841 ( .B1(n9781), .B2(n9786), .A(n9780), .ZN(n9782) );
  OAI211_X1 U10842 ( .C1(n10122), .C2(n9784), .A(n9783), .B(n9782), .ZN(
        P2_U3180) );
  MUX2_X1 U10843 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9785), .S(n9792), .Z(
        P2_U3519) );
  MUX2_X1 U10844 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9786), .S(n9792), .Z(
        P2_U3518) );
  MUX2_X1 U10845 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9787), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10846 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9788), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10847 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9789), .S(n9792), .Z(
        P2_U3515) );
  MUX2_X1 U10848 ( .A(n9790), .B(P2_DATAO_REG_23__SCAN_IN), .S(n10961), .Z(
        P2_U3514) );
  MUX2_X1 U10849 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n5319), .S(n9792), .Z(
        P2_U3513) );
  MUX2_X1 U10850 ( .A(n9978), .B(P2_DATAO_REG_21__SCAN_IN), .S(n10961), .Z(
        P2_U3512) );
  MUX2_X1 U10851 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9988), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10852 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n10004), .S(n9792), .Z(
        P2_U3510) );
  MUX2_X1 U10853 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9791), .S(n9792), .Z(
        P2_U3509) );
  MUX2_X1 U10854 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n10002), .S(n9792), .Z(
        P2_U3508) );
  MUX2_X1 U10855 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9793), .S(n9792), .Z(
        P2_U3507) );
  MUX2_X1 U10856 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9794), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10857 ( .A(n9795), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10961), .Z(
        P2_U3505) );
  MUX2_X1 U10858 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9796), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10859 ( .A(n9797), .B(P2_DATAO_REG_12__SCAN_IN), .S(n10961), .Z(
        P2_U3503) );
  MUX2_X1 U10860 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9798), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10861 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9799), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10862 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9800), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10863 ( .A(n9801), .B(P2_DATAO_REG_8__SCAN_IN), .S(n10961), .Z(
        P2_U3499) );
  MUX2_X1 U10864 ( .A(n9802), .B(P2_DATAO_REG_7__SCAN_IN), .S(n10961), .Z(
        P2_U3498) );
  MUX2_X1 U10865 ( .A(n9803), .B(P2_DATAO_REG_6__SCAN_IN), .S(n10961), .Z(
        P2_U3497) );
  MUX2_X1 U10866 ( .A(n9804), .B(P2_DATAO_REG_5__SCAN_IN), .S(n10961), .Z(
        P2_U3496) );
  MUX2_X1 U10867 ( .A(n9805), .B(P2_DATAO_REG_4__SCAN_IN), .S(n10961), .Z(
        P2_U3495) );
  MUX2_X1 U10868 ( .A(n9806), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10961), .Z(
        P2_U3494) );
  MUX2_X1 U10869 ( .A(n9807), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10961), .Z(
        P2_U3493) );
  MUX2_X1 U10870 ( .A(n6103), .B(P2_DATAO_REG_1__SCAN_IN), .S(n10961), .Z(
        P2_U3492) );
  AOI21_X1 U10871 ( .B1(n5247), .B2(n9809), .A(n9808), .ZN(n9824) );
  INV_X1 U10872 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9816) );
  OAI21_X1 U10873 ( .B1(n9812), .B2(n9811), .A(n9810), .ZN(n9814) );
  AOI21_X1 U10874 ( .B1(n9814), .B2(n5272), .A(n9813), .ZN(n9815) );
  OAI21_X1 U10875 ( .B1(n9873), .B2(n9816), .A(n9815), .ZN(n9821) );
  AOI21_X1 U10876 ( .B1(n5240), .B2(n9818), .A(n9817), .ZN(n9819) );
  NOR2_X1 U10877 ( .A1(n9819), .A2(n10967), .ZN(n9820) );
  AOI211_X1 U10878 ( .C1(n9881), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9823)
         );
  OAI21_X1 U10879 ( .B1(n9824), .B2(n10972), .A(n9823), .ZN(P2_U3196) );
  AOI21_X1 U10880 ( .B1(n10101), .B2(n9826), .A(n9825), .ZN(n9841) );
  AOI21_X1 U10881 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(n9837) );
  NAND2_X1 U10882 ( .A1(n10959), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n9836) );
  OAI21_X1 U10883 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9834) );
  AOI21_X1 U10884 ( .B1(n9834), .B2(n5272), .A(n9833), .ZN(n9835) );
  OAI211_X1 U10885 ( .C1(n9837), .C2(n10972), .A(n9836), .B(n9835), .ZN(n9838)
         );
  AOI21_X1 U10886 ( .B1(n9839), .B2(n9881), .A(n9838), .ZN(n9840) );
  OAI21_X1 U10887 ( .B1(n9841), .B2(n10967), .A(n9840), .ZN(P2_U3197) );
  AOI21_X1 U10888 ( .B1(n5226), .B2(n9843), .A(n9842), .ZN(n9859) );
  INV_X1 U10889 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9850) );
  OAI21_X1 U10890 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9848) );
  AOI21_X1 U10891 ( .B1(n9848), .B2(n5272), .A(n9847), .ZN(n9849) );
  OAI21_X1 U10892 ( .B1(n9873), .B2(n9850), .A(n9849), .ZN(n9856) );
  AOI21_X1 U10893 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9854) );
  NOR2_X1 U10894 ( .A1(n9854), .A2(n10967), .ZN(n9855) );
  AOI211_X1 U10895 ( .C1(n9881), .C2(n9857), .A(n9856), .B(n9855), .ZN(n9858)
         );
  OAI21_X1 U10896 ( .B1(n9859), .B2(n10972), .A(n9858), .ZN(P2_U3198) );
  AOI21_X1 U10897 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9884) );
  NOR2_X1 U10898 ( .A1(n10972), .A2(n9867), .ZN(n9879) );
  OAI21_X1 U10899 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9871) );
  AOI21_X1 U10900 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  OAI21_X1 U10901 ( .B1(n9884), .B2(n10967), .A(n9883), .ZN(P2_U3199) );
  NOR2_X1 U10902 ( .A1(n11018), .A2(n9885), .ZN(n9888) );
  NAND2_X1 U10903 ( .A1(n9888), .A2(n10110), .ZN(n9890) );
  OAI21_X1 U10904 ( .B1(n11015), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9890), .ZN(
        n9889) );
  OAI21_X1 U10905 ( .B1(n9418), .B2(n10030), .A(n9889), .ZN(P2_U3202) );
  OAI21_X1 U10906 ( .B1(n11015), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9890), .ZN(
        n9891) );
  OAI21_X1 U10907 ( .B1(n10114), .B2(n10030), .A(n9891), .ZN(P2_U3203) );
  XNOR2_X1 U10908 ( .A(n9892), .B(n9900), .ZN(n9897) );
  INV_X1 U10909 ( .A(n10048), .ZN(n9906) );
  NAND2_X1 U10910 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  XNOR2_X1 U10911 ( .A(n9901), .B(n9900), .ZN(n10049) );
  AOI22_X1 U10912 ( .A1(n9902), .A2(n10028), .B1(n11018), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9903) );
  OAI21_X1 U10913 ( .B1(n10118), .B2(n10030), .A(n9903), .ZN(n9904) );
  AOI21_X1 U10914 ( .B1(n10049), .B2(n10033), .A(n9904), .ZN(n9905) );
  OAI21_X1 U10915 ( .B1(n9906), .B2(n11018), .A(n9905), .ZN(P2_U3206) );
  INV_X1 U10916 ( .A(n10052), .ZN(n9915) );
  XNOR2_X1 U10917 ( .A(n9910), .B(n9909), .ZN(n10053) );
  AOI22_X1 U10918 ( .A1(n9911), .A2(n10028), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n11018), .ZN(n9912) );
  OAI21_X1 U10919 ( .B1(n10122), .B2(n10030), .A(n9912), .ZN(n9913) );
  AOI21_X1 U10920 ( .B1(n10053), .B2(n10033), .A(n9913), .ZN(n9914) );
  OAI21_X1 U10921 ( .B1(n9915), .B2(n11018), .A(n9914), .ZN(P2_U3207) );
  XNOR2_X1 U10922 ( .A(n9916), .B(n9917), .ZN(n10057) );
  INV_X1 U10923 ( .A(n10057), .ZN(n9928) );
  XNOR2_X1 U10924 ( .A(n9918), .B(n9919), .ZN(n9920) );
  OAI222_X1 U10925 ( .A1(n11003), .A2(n9921), .B1(n11001), .B2(n9944), .C1(
        n11000), .C2(n9920), .ZN(n10056) );
  NAND2_X1 U10926 ( .A1(n10056), .A2(n11015), .ZN(n9927) );
  OAI22_X1 U10927 ( .A1(n9923), .A2(n11010), .B1(n11015), .B2(n9922), .ZN(
        n9924) );
  AOI21_X1 U10928 ( .B1(n9925), .B2(n10015), .A(n9924), .ZN(n9926) );
  OAI211_X1 U10929 ( .C1(n9928), .C2(n10012), .A(n9927), .B(n9926), .ZN(
        P2_U3208) );
  XNOR2_X1 U10930 ( .A(n9930), .B(n9929), .ZN(n9931) );
  OAI222_X1 U10931 ( .A1(n11003), .A2(n9932), .B1(n11001), .B2(n9954), .C1(
        n11000), .C2(n9931), .ZN(n10060) );
  INV_X1 U10932 ( .A(n10060), .ZN(n9939) );
  XNOR2_X1 U10933 ( .A(n9933), .B(n9934), .ZN(n10061) );
  AOI22_X1 U10934 ( .A1(n10028), .A2(n9935), .B1(n11018), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9936) );
  OAI21_X1 U10935 ( .B1(n10130), .B2(n10030), .A(n9936), .ZN(n9937) );
  AOI21_X1 U10936 ( .B1(n10061), .B2(n10033), .A(n9937), .ZN(n9938) );
  OAI21_X1 U10937 ( .B1(n9939), .B2(n11018), .A(n9938), .ZN(P2_U3209) );
  XNOR2_X1 U10938 ( .A(n9941), .B(n9940), .ZN(n9942) );
  OAI222_X1 U10939 ( .A1(n11003), .A2(n9944), .B1(n11001), .B2(n9943), .C1(
        n11000), .C2(n9942), .ZN(n10064) );
  INV_X1 U10940 ( .A(n10064), .ZN(n9951) );
  XNOR2_X1 U10941 ( .A(n9945), .B(n9946), .ZN(n10065) );
  AOI22_X1 U10942 ( .A1(n11018), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n10028), 
        .B2(n9947), .ZN(n9948) );
  OAI21_X1 U10943 ( .B1(n10134), .B2(n10030), .A(n9948), .ZN(n9949) );
  AOI21_X1 U10944 ( .B1(n10065), .B2(n10033), .A(n9949), .ZN(n9950) );
  OAI21_X1 U10945 ( .B1(n9951), .B2(n11018), .A(n9950), .ZN(P2_U3210) );
  XNOR2_X1 U10946 ( .A(n9952), .B(n9956), .ZN(n9953) );
  OAI222_X1 U10947 ( .A1(n11001), .A2(n9955), .B1(n11003), .B2(n9954), .C1(
        n11000), .C2(n9953), .ZN(n10068) );
  INV_X1 U10948 ( .A(n10068), .ZN(n9962) );
  XOR2_X1 U10949 ( .A(n9957), .B(n9956), .Z(n10069) );
  AOI22_X1 U10950 ( .A1(n11018), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n10028), 
        .B2(n9958), .ZN(n9959) );
  OAI21_X1 U10951 ( .B1(n10138), .B2(n10030), .A(n9959), .ZN(n9960) );
  AOI21_X1 U10952 ( .B1(n10069), .B2(n10033), .A(n9960), .ZN(n9961) );
  OAI21_X1 U10953 ( .B1(n11018), .B2(n9962), .A(n9961), .ZN(P2_U3211) );
  OAI21_X1 U10954 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9966) );
  AOI222_X1 U10955 ( .A1(n10041), .A2(n9966), .B1(n5319), .B2(n10003), .C1(
        n9988), .C2(n10001), .ZN(n10074) );
  INV_X1 U10956 ( .A(n9967), .ZN(n9968) );
  OAI22_X1 U10957 ( .A1(n11015), .A2(n9969), .B1(n9968), .B2(n11010), .ZN(
        n9973) );
  OAI21_X1 U10958 ( .B1(n5223), .B2(n9971), .A(n9970), .ZN(n10075) );
  NOR2_X1 U10959 ( .A1(n10075), .A2(n10012), .ZN(n9972) );
  AOI211_X1 U10960 ( .C1(n10015), .C2(n10072), .A(n9973), .B(n9972), .ZN(n9974) );
  OAI21_X1 U10961 ( .B1(n11018), .B2(n10074), .A(n9974), .ZN(P2_U3212) );
  OAI21_X1 U10962 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(n9979) );
  AOI222_X1 U10963 ( .A1(n10041), .A2(n9979), .B1(n9978), .B2(n10003), .C1(
        n10004), .C2(n10001), .ZN(n10076) );
  OAI21_X1 U10964 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n10078) );
  AOI22_X1 U10965 ( .A1(n11018), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9983), 
        .B2(n10028), .ZN(n9984) );
  OAI21_X1 U10966 ( .B1(n10143), .B2(n10030), .A(n9984), .ZN(n9985) );
  AOI21_X1 U10967 ( .B1(n10078), .B2(n10033), .A(n9985), .ZN(n9986) );
  OAI21_X1 U10968 ( .B1(n10076), .B2(n11018), .A(n9986), .ZN(P2_U3213) );
  XNOR2_X1 U10969 ( .A(n9987), .B(n9995), .ZN(n9991) );
  NAND2_X1 U10970 ( .A1(n9988), .A2(n10003), .ZN(n9989) );
  OAI21_X1 U10971 ( .B1(n10020), .B2(n11001), .A(n9989), .ZN(n9990) );
  AOI21_X1 U10972 ( .B1(n9991), .B2(n10041), .A(n9990), .ZN(n10082) );
  INV_X1 U10973 ( .A(n9992), .ZN(n9993) );
  OAI22_X1 U10974 ( .A1(n11015), .A2(n5875), .B1(n9993), .B2(n11010), .ZN(
        n9998) );
  OAI21_X1 U10975 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n10081) );
  NOR2_X1 U10976 ( .A1(n10081), .A2(n10012), .ZN(n9997) );
  AOI211_X1 U10977 ( .C1(n10015), .C2(n10146), .A(n9998), .B(n9997), .ZN(n9999) );
  OAI21_X1 U10978 ( .B1(n11018), .B2(n10082), .A(n9999), .ZN(P2_U3214) );
  XNOR2_X1 U10979 ( .A(n10000), .B(n10010), .ZN(n10005) );
  AOI222_X1 U10980 ( .A1(n10041), .A2(n10005), .B1(n10004), .B2(n10003), .C1(
        n10002), .C2(n10001), .ZN(n10088) );
  INV_X1 U10981 ( .A(n10006), .ZN(n10007) );
  OAI22_X1 U10982 ( .A1(n11015), .A2(n10008), .B1(n10007), .B2(n11010), .ZN(
        n10014) );
  OAI21_X1 U10983 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(n10089) );
  NOR2_X1 U10984 ( .A1(n10089), .A2(n10012), .ZN(n10013) );
  AOI211_X1 U10985 ( .C1(n10015), .C2(n10086), .A(n10014), .B(n10013), .ZN(
        n10016) );
  OAI21_X1 U10986 ( .B1(n11018), .B2(n10088), .A(n10016), .ZN(P2_U3215) );
  OAI211_X1 U10987 ( .C1(n10018), .C2(n10024), .A(n10017), .B(n10041), .ZN(
        n10023) );
  OAI22_X1 U10988 ( .A1(n10020), .A2(n11003), .B1(n11001), .B2(n10019), .ZN(
        n10021) );
  INV_X1 U10989 ( .A(n10021), .ZN(n10022) );
  AND2_X1 U10990 ( .A1(n10023), .A2(n10022), .ZN(n10091) );
  NAND2_X1 U10991 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND2_X1 U10992 ( .A1(n5245), .A2(n10026), .ZN(n10090) );
  INV_X1 U10993 ( .A(n10151), .ZN(n10031) );
  AOI22_X1 U10994 ( .A1(n11018), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n10028), 
        .B2(n10027), .ZN(n10029) );
  OAI21_X1 U10995 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10032) );
  AOI21_X1 U10996 ( .B1(n10090), .B2(n10033), .A(n10032), .ZN(n10034) );
  OAI21_X1 U10997 ( .B1(n11018), .B2(n10091), .A(n10034), .ZN(P2_U3216) );
  NOR2_X1 U10998 ( .A1(n10110), .A2(n11185), .ZN(n10036) );
  AOI21_X1 U10999 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n11185), .A(n10036), 
        .ZN(n10035) );
  OAI21_X1 U11000 ( .B1(n9418), .B2(n10103), .A(n10035), .ZN(P2_U3490) );
  AOI21_X1 U11001 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n11185), .A(n10036), 
        .ZN(n10037) );
  OAI21_X1 U11002 ( .B1(n10114), .B2(n10103), .A(n10037), .ZN(P2_U3489) );
  NAND2_X1 U11003 ( .A1(n10042), .A2(n10041), .ZN(n10046) );
  INV_X1 U11004 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10050) );
  AOI21_X1 U11005 ( .B1(n10049), .B2(n11159), .A(n10048), .ZN(n10115) );
  MUX2_X1 U11006 ( .A(n10050), .B(n10115), .S(n11187), .Z(n10051) );
  OAI21_X1 U11007 ( .B1(n10118), .B2(n10103), .A(n10051), .ZN(P2_U3486) );
  INV_X1 U11008 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U11009 ( .B1(n10122), .B2(n10103), .A(n10055), .ZN(P2_U3485) );
  INV_X1 U11010 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10058) );
  AOI21_X1 U11011 ( .B1(n11159), .B2(n10057), .A(n10056), .ZN(n10123) );
  MUX2_X1 U11012 ( .A(n10058), .B(n10123), .S(n11187), .Z(n10059) );
  OAI21_X1 U11013 ( .B1(n10126), .B2(n10103), .A(n10059), .ZN(P2_U3484) );
  INV_X1 U11014 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10062) );
  AOI21_X1 U11015 ( .B1(n10061), .B2(n11159), .A(n10060), .ZN(n10127) );
  MUX2_X1 U11016 ( .A(n10062), .B(n10127), .S(n11187), .Z(n10063) );
  OAI21_X1 U11017 ( .B1(n10130), .B2(n10103), .A(n10063), .ZN(P2_U3483) );
  INV_X1 U11018 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10066) );
  AOI21_X1 U11019 ( .B1(n10065), .B2(n11159), .A(n10064), .ZN(n10131) );
  MUX2_X1 U11020 ( .A(n10066), .B(n10131), .S(n11187), .Z(n10067) );
  OAI21_X1 U11021 ( .B1(n10134), .B2(n10103), .A(n10067), .ZN(P2_U3482) );
  AOI21_X1 U11022 ( .B1(n10069), .B2(n11159), .A(n10068), .ZN(n10136) );
  INV_X1 U11023 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10070) );
  MUX2_X1 U11024 ( .A(n10136), .B(n10070), .S(n11185), .Z(n10071) );
  OAI21_X1 U11025 ( .B1(n10138), .B2(n10103), .A(n10071), .ZN(P2_U3481) );
  NAND2_X1 U11026 ( .A1(n10072), .A2(n11158), .ZN(n10073) );
  OAI211_X1 U11027 ( .C1(n11181), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10139) );
  MUX2_X1 U11028 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n10139), .S(n11187), .Z(
        P2_U3480) );
  INV_X1 U11029 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10079) );
  INV_X1 U11030 ( .A(n10076), .ZN(n10077) );
  AOI21_X1 U11031 ( .B1(n11159), .B2(n10078), .A(n10077), .ZN(n10140) );
  MUX2_X1 U11032 ( .A(n10079), .B(n10140), .S(n11187), .Z(n10080) );
  OAI21_X1 U11033 ( .B1(n10143), .B2(n10103), .A(n10080), .ZN(P2_U3479) );
  INV_X1 U11034 ( .A(n10103), .ZN(n10108) );
  OR2_X1 U11035 ( .A1(n10081), .A2(n11181), .ZN(n10083) );
  NAND2_X1 U11036 ( .A1(n10083), .A2(n10082), .ZN(n10144) );
  MUX2_X1 U11037 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n10144), .S(n11187), .Z(
        n10084) );
  AOI21_X1 U11038 ( .B1(n10108), .B2(n10146), .A(n10084), .ZN(n10085) );
  INV_X1 U11039 ( .A(n10085), .ZN(P2_U3478) );
  NAND2_X1 U11040 ( .A1(n10086), .A2(n11158), .ZN(n10087) );
  OAI211_X1 U11041 ( .C1(n11181), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10148) );
  MUX2_X1 U11042 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n10148), .S(n11187), .Z(
        P2_U3477) );
  NAND2_X1 U11043 ( .A1(n10090), .A2(n11159), .ZN(n10092) );
  NAND2_X1 U11044 ( .A1(n10092), .A2(n10091), .ZN(n10149) );
  MUX2_X1 U11045 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n10149), .S(n11187), .Z(
        n10093) );
  AOI21_X1 U11046 ( .B1(n10108), .B2(n10151), .A(n10093), .ZN(n10094) );
  INV_X1 U11047 ( .A(n10094), .ZN(P2_U3476) );
  AOI21_X1 U11048 ( .B1(n10096), .B2(n11159), .A(n10095), .ZN(n10153) );
  MUX2_X1 U11049 ( .A(n10097), .B(n10153), .S(n11187), .Z(n10098) );
  OAI21_X1 U11050 ( .B1(n10156), .B2(n10103), .A(n10098), .ZN(P2_U3475) );
  AOI21_X1 U11051 ( .B1(n10100), .B2(n11159), .A(n10099), .ZN(n10157) );
  MUX2_X1 U11052 ( .A(n10101), .B(n10157), .S(n11187), .Z(n10102) );
  OAI21_X1 U11053 ( .B1(n10161), .B2(n10103), .A(n10102), .ZN(P2_U3474) );
  NAND2_X1 U11054 ( .A1(n10104), .A2(n11159), .ZN(n10106) );
  NAND2_X1 U11055 ( .A1(n10106), .A2(n10105), .ZN(n10162) );
  MUX2_X1 U11056 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n10162), .S(n11187), .Z(
        n10107) );
  AOI21_X1 U11057 ( .B1(n10108), .B2(n10164), .A(n10107), .ZN(n10109) );
  INV_X1 U11058 ( .A(n10109), .ZN(P2_U3473) );
  NOR2_X1 U11059 ( .A1(n10110), .A2(n11188), .ZN(n10112) );
  AOI21_X1 U11060 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n11188), .A(n10112), 
        .ZN(n10111) );
  OAI21_X1 U11061 ( .B1(n9418), .B2(n10160), .A(n10111), .ZN(P2_U3458) );
  AOI21_X1 U11062 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n11188), .A(n10112), 
        .ZN(n10113) );
  OAI21_X1 U11063 ( .B1(n10114), .B2(n10160), .A(n10113), .ZN(P2_U3457) );
  INV_X1 U11064 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10116) );
  MUX2_X1 U11065 ( .A(n10116), .B(n10115), .S(n11191), .Z(n10117) );
  OAI21_X1 U11066 ( .B1(n10118), .B2(n10160), .A(n10117), .ZN(P2_U3454) );
  INV_X1 U11067 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10120) );
  OAI21_X1 U11068 ( .B1(n10122), .B2(n10160), .A(n10121), .ZN(P2_U3453) );
  INV_X1 U11069 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U11070 ( .A(n10124), .B(n10123), .S(n11191), .Z(n10125) );
  OAI21_X1 U11071 ( .B1(n10126), .B2(n10160), .A(n10125), .ZN(P2_U3452) );
  INV_X1 U11072 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U11073 ( .A(n10128), .B(n10127), .S(n11191), .Z(n10129) );
  OAI21_X1 U11074 ( .B1(n10130), .B2(n10160), .A(n10129), .ZN(P2_U3451) );
  INV_X1 U11075 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U11076 ( .A(n10132), .B(n10131), .S(n11191), .Z(n10133) );
  OAI21_X1 U11077 ( .B1(n10134), .B2(n10160), .A(n10133), .ZN(P2_U3450) );
  INV_X1 U11078 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U11079 ( .A(n10136), .B(n10135), .S(n11188), .Z(n10137) );
  OAI21_X1 U11080 ( .B1(n10138), .B2(n10160), .A(n10137), .ZN(P2_U3449) );
  MUX2_X1 U11081 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n10139), .S(n11191), .Z(
        P2_U3448) );
  INV_X1 U11082 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10141) );
  MUX2_X1 U11083 ( .A(n10141), .B(n10140), .S(n11191), .Z(n10142) );
  OAI21_X1 U11084 ( .B1(n10143), .B2(n10160), .A(n10142), .ZN(P2_U3447) );
  INV_X1 U11085 ( .A(n10160), .ZN(n10165) );
  MUX2_X1 U11086 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n10144), .S(n11191), .Z(
        n10145) );
  AOI21_X1 U11087 ( .B1(n10165), .B2(n10146), .A(n10145), .ZN(n10147) );
  INV_X1 U11088 ( .A(n10147), .ZN(P2_U3446) );
  MUX2_X1 U11089 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n10148), .S(n11191), .Z(
        P2_U3444) );
  MUX2_X1 U11090 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n10149), .S(n11191), .Z(
        n10150) );
  AOI21_X1 U11091 ( .B1(n10165), .B2(n10151), .A(n10150), .ZN(n10152) );
  INV_X1 U11092 ( .A(n10152), .ZN(P2_U3441) );
  INV_X1 U11093 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10154) );
  MUX2_X1 U11094 ( .A(n10154), .B(n10153), .S(n11191), .Z(n10155) );
  OAI21_X1 U11095 ( .B1(n10156), .B2(n10160), .A(n10155), .ZN(P2_U3438) );
  INV_X1 U11096 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10158) );
  MUX2_X1 U11097 ( .A(n10158), .B(n10157), .S(n11191), .Z(n10159) );
  OAI21_X1 U11098 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(P2_U3435) );
  MUX2_X1 U11099 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n10162), .S(n11191), .Z(
        n10163) );
  AOI21_X1 U11100 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(n10166) );
  INV_X1 U11101 ( .A(n10166), .ZN(P2_U3432) );
  INV_X1 U11102 ( .A(n10694), .ZN(n10171) );
  NOR4_X1 U11103 ( .A1(n10167), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), 
        .A4(n5821), .ZN(n10168) );
  AOI21_X1 U11104 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n10169), .A(n10168), 
        .ZN(n10170) );
  OAI21_X1 U11105 ( .B1(n10171), .B2(n10175), .A(n10170), .ZN(P2_U3264) );
  INV_X1 U11106 ( .A(n10172), .ZN(n10699) );
  INV_X1 U11107 ( .A(n10177), .ZN(n10178) );
  MUX2_X1 U11108 ( .A(n10178), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U11109 ( .B1(n10181), .B2(n10179), .A(n10180), .ZN(n10182) );
  NAND2_X1 U11110 ( .A1(n10182), .A2(n10308), .ZN(n10186) );
  NOR2_X1 U11111 ( .A1(n10300), .A2(n10506), .ZN(n10184) );
  OAI22_X1 U11112 ( .A1(n10313), .A2(n10200), .B1(n10299), .B2(n10531), .ZN(
        n10183) );
  AOI211_X1 U11113 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n10184), 
        .B(n10183), .ZN(n10185) );
  OAI211_X1 U11114 ( .C1(n9318), .C2(n10318), .A(n10186), .B(n10185), .ZN(
        P1_U3216) );
  XOR2_X1 U11115 ( .A(n10188), .B(n10187), .Z(n10194) );
  INV_X1 U11116 ( .A(n10299), .ZN(n10190) );
  AOI22_X1 U11117 ( .A1(n10315), .A2(n10571), .B1(n10190), .B2(n10189), .ZN(
        n10191) );
  NAND2_X1 U11118 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10432)
         );
  OAI211_X1 U11119 ( .C1(n10241), .C2(n10313), .A(n10191), .B(n10432), .ZN(
        n10192) );
  AOI21_X1 U11120 ( .B1(n10669), .B2(n10289), .A(n10192), .ZN(n10193) );
  OAI21_X1 U11121 ( .B1(n10194), .B2(n10292), .A(n10193), .ZN(P1_U3219) );
  AOI21_X1 U11122 ( .B1(n10196), .B2(n10195), .A(n10292), .ZN(n10198) );
  NAND2_X1 U11123 ( .A1(n10198), .A2(n10197), .ZN(n10204) );
  NOR2_X1 U11124 ( .A1(n10313), .A2(n10199), .ZN(n10202) );
  OAI22_X1 U11125 ( .A1(n10300), .A2(n10200), .B1(n10299), .B2(n10579), .ZN(
        n10201) );
  AOI211_X1 U11126 ( .C1(P1_REG3_REG_21__SCAN_IN), .C2(P1_U3086), .A(n10202), 
        .B(n10201), .ZN(n10203) );
  OAI211_X1 U11127 ( .C1(n10658), .C2(n10318), .A(n10204), .B(n10203), .ZN(
        P1_U3223) );
  AOI21_X1 U11128 ( .B1(n10206), .B2(n10205), .A(n5167), .ZN(n10211) );
  OAI22_X1 U11129 ( .A1(n10300), .A2(n10504), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10207), .ZN(n10209) );
  OAI22_X1 U11130 ( .A1(n10313), .A2(n10506), .B1(n10299), .B2(n10496), .ZN(
        n10208) );
  AOI211_X1 U11131 ( .C1(n10637), .C2(n10289), .A(n10209), .B(n10208), .ZN(
        n10210) );
  OAI21_X1 U11132 ( .B1(n10211), .B2(n10292), .A(n10210), .ZN(P1_U3225) );
  NAND2_X1 U11133 ( .A1(n10212), .A2(n10213), .ZN(n10236) );
  OAI21_X1 U11134 ( .B1(n10213), .B2(n10212), .A(n10236), .ZN(n10214) );
  NAND2_X1 U11135 ( .A1(n10214), .A2(n10308), .ZN(n10218) );
  AND2_X1 U11136 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10400) );
  OAI22_X1 U11137 ( .A1(n10313), .A2(n10215), .B1(n10299), .B2(n10589), .ZN(
        n10216) );
  AOI211_X1 U11138 ( .C1(n10315), .C2(n10595), .A(n10400), .B(n10216), .ZN(
        n10217) );
  OAI211_X1 U11139 ( .C1(n11224), .C2(n10318), .A(n10218), .B(n10217), .ZN(
        P1_U3226) );
  NOR2_X1 U11140 ( .A1(n10220), .A2(n10219), .ZN(n10224) );
  XNOR2_X1 U11141 ( .A(n10222), .B(n10221), .ZN(n10223) );
  XNOR2_X1 U11142 ( .A(n10224), .B(n10223), .ZN(n10225) );
  NAND2_X1 U11143 ( .A1(n10225), .A2(n10308), .ZN(n10234) );
  NAND2_X1 U11144 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10773) );
  INV_X1 U11145 ( .A(n10773), .ZN(n10226) );
  AOI21_X1 U11146 ( .B1(n10315), .B2(n10332), .A(n10226), .ZN(n10233) );
  OAI22_X1 U11147 ( .A1(n10313), .A2(n10228), .B1(n10299), .B2(n10227), .ZN(
        n10229) );
  INV_X1 U11148 ( .A(n10229), .ZN(n10232) );
  NAND2_X1 U11149 ( .A1(n10289), .A2(n10230), .ZN(n10231) );
  NAND4_X1 U11150 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        P1_U3227) );
  NAND2_X1 U11151 ( .A1(n10236), .A2(n10235), .ZN(n10240) );
  NAND2_X1 U11152 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  XNOR2_X1 U11153 ( .A(n10240), .B(n10239), .ZN(n10246) );
  NAND2_X1 U11154 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10887)
         );
  OAI21_X1 U11155 ( .B1(n10241), .B2(n10300), .A(n10887), .ZN(n10244) );
  OAI22_X1 U11156 ( .A1(n10313), .A2(n10242), .B1(n10299), .B2(n11241), .ZN(
        n10243) );
  AOI211_X1 U11157 ( .C1(n11260), .C2(n10289), .A(n10244), .B(n10243), .ZN(
        n10245) );
  OAI21_X1 U11158 ( .B1(n10246), .B2(n10292), .A(n10245), .ZN(P1_U3228) );
  NAND2_X1 U11159 ( .A1(n5233), .A2(n10248), .ZN(n10249) );
  XNOR2_X1 U11160 ( .A(n10247), .B(n10249), .ZN(n10254) );
  OAI22_X1 U11161 ( .A1(n10300), .A2(n10483), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10250), .ZN(n10252) );
  OAI22_X1 U11162 ( .A1(n10313), .A2(n10272), .B1(n10299), .B2(n10521), .ZN(
        n10251) );
  AOI211_X1 U11163 ( .C1(n10642), .C2(n10289), .A(n10252), .B(n10251), .ZN(
        n10253) );
  OAI21_X1 U11164 ( .B1(n10254), .B2(n10292), .A(n10253), .ZN(P1_U3229) );
  XOR2_X1 U11165 ( .A(n10255), .B(n10256), .Z(n10262) );
  OAI22_X1 U11166 ( .A1(n10300), .A2(n10271), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10257), .ZN(n10260) );
  OAI22_X1 U11167 ( .A1(n10313), .A2(n10284), .B1(n10299), .B2(n10258), .ZN(
        n10259) );
  AOI211_X1 U11168 ( .C1(n10664), .C2(n10289), .A(n10260), .B(n10259), .ZN(
        n10261) );
  OAI21_X1 U11169 ( .B1(n10262), .B2(n10292), .A(n10261), .ZN(P1_U3233) );
  INV_X1 U11170 ( .A(n10263), .ZN(n10269) );
  INV_X1 U11171 ( .A(n10264), .ZN(n10266) );
  AOI21_X1 U11172 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10268) );
  AOI21_X1 U11173 ( .B1(n10179), .B2(n10269), .A(n10268), .ZN(n10276) );
  OAI22_X1 U11174 ( .A1(n10313), .A2(n10271), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10270), .ZN(n10274) );
  OAI22_X1 U11175 ( .A1(n10300), .A2(n10272), .B1(n10299), .B2(n10557), .ZN(
        n10273) );
  AOI211_X1 U11176 ( .C1(n10652), .C2(n10289), .A(n10274), .B(n10273), .ZN(
        n10275) );
  OAI21_X1 U11177 ( .B1(n10276), .B2(n10292), .A(n10275), .ZN(P1_U3235) );
  NAND2_X1 U11178 ( .A1(n10212), .A2(n10277), .ZN(n10279) );
  NAND2_X1 U11179 ( .A1(n10279), .A2(n10278), .ZN(n10281) );
  NAND2_X1 U11180 ( .A1(n10281), .A2(n10280), .ZN(n10283) );
  XNOR2_X1 U11181 ( .A(n10283), .B(n10282), .ZN(n10293) );
  NAND2_X1 U11182 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10903)
         );
  OAI21_X1 U11183 ( .B1(n10300), .B2(n10284), .A(n10903), .ZN(n10288) );
  OAI22_X1 U11184 ( .A1(n10313), .A2(n10286), .B1(n10299), .B2(n10285), .ZN(
        n10287) );
  AOI211_X1 U11185 ( .C1(n10290), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10291) );
  OAI21_X1 U11186 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(P1_U3238) );
  INV_X1 U11187 ( .A(n10632), .ZN(n10305) );
  INV_X1 U11188 ( .A(n10294), .ZN(n10298) );
  OAI21_X1 U11189 ( .B1(n5167), .B2(n10296), .A(n10295), .ZN(n10297) );
  NAND3_X1 U11190 ( .A1(n10298), .A2(n10308), .A3(n10297), .ZN(n10304) );
  NOR2_X1 U11191 ( .A1(n10313), .A2(n10483), .ZN(n10302) );
  OAI22_X1 U11192 ( .A1(n10300), .A2(n10482), .B1(n10299), .B2(n10486), .ZN(
        n10301) );
  AOI211_X1 U11193 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n10302), 
        .B(n10301), .ZN(n10303) );
  OAI211_X1 U11194 ( .C1(n10305), .C2(n10318), .A(n10304), .B(n10303), .ZN(
        P1_U3240) );
  NAND2_X1 U11195 ( .A1(n10309), .A2(n10308), .ZN(n10317) );
  NOR2_X1 U11196 ( .A1(n10310), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10869) );
  INV_X1 U11197 ( .A(n11215), .ZN(n10311) );
  OAI22_X1 U11198 ( .A1(n10313), .A2(n10312), .B1(n10299), .B2(n10311), .ZN(
        n10314) );
  AOI211_X1 U11199 ( .C1(n10315), .C2(n11235), .A(n10869), .B(n10314), .ZN(
        n10316) );
  OAI211_X1 U11200 ( .C1(n7338), .C2(n10318), .A(n10317), .B(n10316), .ZN(
        P1_U3241) );
  MUX2_X1 U11201 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10319), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U11202 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10320), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11203 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10321), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U11204 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10322), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11205 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10323), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11206 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10324), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11207 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10513), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11208 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10541), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11209 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10549), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U11210 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10570), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11211 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10550), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11212 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10571), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11213 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n11238), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11214 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10595), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11215 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n11235), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U11216 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10594), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U11217 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n11210), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11218 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10325), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U11219 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10326), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U11220 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10327), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11221 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10328), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11222 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10329), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U11223 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10330), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11224 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10331), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11225 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10332), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U11226 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10333), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11227 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10334), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U11228 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10335), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11229 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10336), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U11230 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10337), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U11231 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10338), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U11232 ( .C1(n10341), .C2(n10340), .A(n10895), .B(n10339), .ZN(
        n10349) );
  OAI211_X1 U11233 ( .C1(n10344), .C2(n10343), .A(n10846), .B(n10342), .ZN(
        n10348) );
  AOI22_X1 U11234 ( .A1(n10430), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10347) );
  NAND2_X1 U11235 ( .A1(n10929), .A2(n10345), .ZN(n10346) );
  NAND4_X1 U11236 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        P1_U3244) );
  OAI211_X1 U11237 ( .C1(n10352), .C2(n10351), .A(n10895), .B(n10350), .ZN(
        n10362) );
  OAI211_X1 U11238 ( .C1(n10355), .C2(n10354), .A(n10846), .B(n10353), .ZN(
        n10361) );
  INV_X1 U11239 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10357) );
  OAI21_X1 U11240 ( .B1(n10933), .B2(n10357), .A(n10356), .ZN(n10358) );
  AOI21_X1 U11241 ( .B1(n10929), .B2(n10359), .A(n10358), .ZN(n10360) );
  NAND3_X1 U11242 ( .A1(n10362), .A2(n10361), .A3(n10360), .ZN(P1_U3246) );
  NOR2_X1 U11243 ( .A1(n10433), .A2(n10363), .ZN(n10364) );
  AOI211_X1 U11244 ( .C1(n10430), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10365), .B(
        n10364), .ZN(n10375) );
  OAI211_X1 U11245 ( .C1(n10368), .C2(n10367), .A(n10846), .B(n10366), .ZN(
        n10373) );
  OAI211_X1 U11246 ( .C1(n10371), .C2(n10370), .A(n10895), .B(n10369), .ZN(
        n10372) );
  NAND4_X1 U11247 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        P1_U3247) );
  INV_X1 U11248 ( .A(n10407), .ZN(n10406) );
  OR2_X1 U11249 ( .A1(n10407), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U11250 ( .A1(n10407), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10376) );
  AND2_X1 U11251 ( .A1(n10420), .A2(n10376), .ZN(n10388) );
  NOR2_X1 U11252 ( .A1(n10914), .A2(n10377), .ZN(n10378) );
  AOI21_X1 U11253 ( .B1(n10914), .B2(n10377), .A(n10378), .ZN(n10907) );
  OAI21_X1 U11254 ( .B1(n10390), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10379), 
        .ZN(n10908) );
  NOR2_X1 U11255 ( .A1(n10907), .A2(n10908), .ZN(n10906) );
  AOI21_X1 U11256 ( .B1(n10914), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10906), 
        .ZN(n10843) );
  NAND2_X1 U11257 ( .A1(n10847), .A2(n10383), .ZN(n10381) );
  NAND2_X1 U11258 ( .A1(n10393), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10380) );
  AND2_X1 U11259 ( .A1(n10381), .A2(n10380), .ZN(n10844) );
  NOR2_X1 U11260 ( .A1(n10843), .A2(n10844), .ZN(n10842) );
  INV_X1 U11261 ( .A(n10842), .ZN(n10382) );
  OAI21_X1 U11262 ( .B1(n10393), .B2(n10383), .A(n10382), .ZN(n10384) );
  AND2_X1 U11263 ( .A1(n10384), .A2(n10859), .ZN(n10386) );
  NOR2_X1 U11264 ( .A1(n10384), .A2(n10859), .ZN(n10385) );
  OR2_X1 U11265 ( .A1(n10386), .A2(n10385), .ZN(n10861) );
  NOR2_X1 U11266 ( .A1(n10861), .A2(n6592), .ZN(n10860) );
  NOR2_X1 U11267 ( .A1(n10386), .A2(n10860), .ZN(n10387) );
  NAND2_X1 U11268 ( .A1(n10388), .A2(n10387), .ZN(n10421) );
  OAI21_X1 U11269 ( .B1(n10388), .B2(n10387), .A(n10421), .ZN(n10404) );
  INV_X1 U11270 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10402) );
  OAI21_X1 U11271 ( .B1(n10390), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10389), 
        .ZN(n10911) );
  NAND2_X1 U11272 ( .A1(n10914), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10391) );
  OAI21_X1 U11273 ( .B1(n10914), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10391), 
        .ZN(n10910) );
  NOR2_X1 U11274 ( .A1(n10911), .A2(n10910), .ZN(n10909) );
  AOI21_X1 U11275 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10914), .A(n10909), 
        .ZN(n10839) );
  AOI22_X1 U11276 ( .A1(n10847), .A2(n10392), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n10393), .ZN(n10838) );
  OAI21_X1 U11277 ( .B1(n10393), .B2(n10392), .A(n10841), .ZN(n10394) );
  AND2_X1 U11278 ( .A1(n10394), .A2(n10859), .ZN(n10396) );
  NOR2_X1 U11279 ( .A1(n10394), .A2(n10859), .ZN(n10395) );
  NOR2_X1 U11280 ( .A1(n6593), .A2(n10855), .ZN(n10856) );
  NOR2_X1 U11281 ( .A1(n10396), .A2(n10856), .ZN(n10398) );
  XNOR2_X1 U11282 ( .A(n10407), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U11283 ( .A1(n10397), .A2(n10398), .ZN(n10409) );
  AOI211_X1 U11284 ( .C1(n10398), .C2(n10397), .A(n10409), .B(n10922), .ZN(
        n10399) );
  NOR2_X1 U11285 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  OAI21_X1 U11286 ( .B1(n10933), .B2(n10402), .A(n10401), .ZN(n10403) );
  AOI21_X1 U11287 ( .B1(n10846), .B2(n10404), .A(n10403), .ZN(n10405) );
  OAI21_X1 U11288 ( .B1(n10406), .B2(n10433), .A(n10405), .ZN(P1_U3259) );
  AND2_X1 U11289 ( .A1(n10407), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10408) );
  XNOR2_X1 U11290 ( .A(n10877), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n10873) );
  INV_X1 U11291 ( .A(n10877), .ZN(n10423) );
  INV_X1 U11292 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U11293 ( .A1(n10423), .A2(n10410), .ZN(n10411) );
  NAND2_X1 U11294 ( .A1(n10876), .A2(n10411), .ZN(n10893) );
  INV_X1 U11295 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U11296 ( .A1(n10898), .A2(n10413), .ZN(n10412) );
  OAI21_X1 U11297 ( .B1(n10898), .B2(n10413), .A(n10412), .ZN(n10896) );
  INV_X1 U11298 ( .A(n10896), .ZN(n10414) );
  INV_X1 U11299 ( .A(n10894), .ZN(n10415) );
  AOI21_X1 U11300 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n10898), .A(n10415), 
        .ZN(n10417) );
  MUX2_X1 U11301 ( .A(n6855), .B(P1_REG2_REG_19__SCAN_IN), .S(n10599), .Z(
        n10416) );
  XNOR2_X1 U11302 ( .A(n10417), .B(n10416), .ZN(n10437) );
  INV_X1 U11303 ( .A(n10898), .ZN(n10426) );
  NAND2_X1 U11304 ( .A1(n10877), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10418) );
  OAI21_X1 U11305 ( .B1(n10877), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10418), 
        .ZN(n10419) );
  INV_X1 U11306 ( .A(n10419), .ZN(n10880) );
  NAND2_X1 U11307 ( .A1(n10421), .A2(n10420), .ZN(n10879) );
  NAND2_X1 U11308 ( .A1(n10880), .A2(n10879), .ZN(n10878) );
  NAND2_X1 U11309 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  NAND2_X1 U11310 ( .A1(n10898), .A2(n10427), .ZN(n10425) );
  OAI21_X1 U11311 ( .B1(n10898), .B2(n10427), .A(n10425), .ZN(n10891) );
  NAND2_X1 U11312 ( .A1(n10892), .A2(n10891), .ZN(n10890) );
  OAI21_X1 U11313 ( .B1(n10427), .B2(n10426), .A(n10890), .ZN(n10429) );
  XNOR2_X1 U11314 ( .A(n10599), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10428) );
  XNOR2_X1 U11315 ( .A(n10429), .B(n10428), .ZN(n10435) );
  NAND2_X1 U11316 ( .A1(n10430), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n10431) );
  OAI211_X1 U11317 ( .C1(n10433), .C2(n7172), .A(n10432), .B(n10431), .ZN(
        n10434) );
  AOI21_X1 U11318 ( .B1(n10846), .B2(n10435), .A(n10434), .ZN(n10436) );
  OAI21_X1 U11319 ( .B1(n10437), .B2(n10922), .A(n10436), .ZN(P1_U3262) );
  XNOR2_X1 U11320 ( .A(n5448), .B(n10438), .ZN(n10439) );
  NAND2_X1 U11321 ( .A1(n10439), .A2(n11250), .ZN(n10612) );
  NOR2_X1 U11322 ( .A1(n10600), .A2(n10440), .ZN(n10442) );
  AOI211_X1 U11323 ( .C1(n10443), .C2(n11245), .A(n10442), .B(n10441), .ZN(
        n10444) );
  OAI21_X1 U11324 ( .B1(n10612), .B2(n11253), .A(n10444), .ZN(P1_U3264) );
  OAI222_X1 U11325 ( .A1(n10507), .A2(n10482), .B1(n10505), .B2(n10447), .C1(
        n10503), .C2(n10446), .ZN(n10623) );
  OAI211_X1 U11326 ( .C1(n10449), .C2(n10461), .A(n11250), .B(n10448), .ZN(
        n10619) );
  NAND2_X1 U11327 ( .A1(n11258), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n10450) );
  OAI21_X1 U11328 ( .B1(n10451), .B2(n10580), .A(n10450), .ZN(n10452) );
  AOI21_X1 U11329 ( .B1(n10618), .B2(n11245), .A(n10452), .ZN(n10453) );
  OAI21_X1 U11330 ( .B1(n10619), .B2(n11253), .A(n10453), .ZN(n10458) );
  OAI21_X1 U11331 ( .B1(n10456), .B2(n10455), .A(n10454), .ZN(n10621) );
  NOR2_X1 U11332 ( .A1(n10621), .A2(n11254), .ZN(n10457) );
  AOI211_X1 U11333 ( .C1(n10600), .C2(n10623), .A(n10458), .B(n10457), .ZN(
        n10459) );
  INV_X1 U11334 ( .A(n10459), .ZN(P1_U3265) );
  XOR2_X1 U11335 ( .A(n10467), .B(n10460), .Z(n10629) );
  AOI211_X1 U11336 ( .C1(n10627), .C2(n10484), .A(n10609), .B(n10461), .ZN(
        n10626) );
  NOR2_X1 U11337 ( .A1(n10462), .A2(n10534), .ZN(n10466) );
  OAI22_X1 U11338 ( .A1(n10600), .A2(n10464), .B1(n10463), .B2(n10580), .ZN(
        n10465) );
  AOI211_X1 U11339 ( .C1(n10626), .C2(n10560), .A(n10466), .B(n10465), .ZN(
        n10476) );
  AND2_X1 U11340 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  NAND2_X1 U11341 ( .A1(n10474), .A2(n10473), .ZN(n10625) );
  NAND2_X1 U11342 ( .A1(n10625), .A2(n10600), .ZN(n10475) );
  OAI211_X1 U11343 ( .C1(n10629), .C2(n11254), .A(n10476), .B(n10475), .ZN(
        P1_U3266) );
  XNOR2_X1 U11344 ( .A(n10477), .B(n10479), .ZN(n10634) );
  AOI22_X1 U11345 ( .A1(n10632), .A2(n11245), .B1(n11258), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n10490) );
  AOI21_X1 U11346 ( .B1(n10480), .B2(n10479), .A(n10478), .ZN(n10481) );
  OAI222_X1 U11347 ( .A1(n10507), .A2(n10483), .B1(n10505), .B2(n10482), .C1(
        n10503), .C2(n10481), .ZN(n10630) );
  INV_X1 U11348 ( .A(n10484), .ZN(n10485) );
  AOI211_X1 U11349 ( .C1(n10632), .C2(n10492), .A(n10609), .B(n10485), .ZN(
        n10631) );
  INV_X1 U11350 ( .A(n10631), .ZN(n10487) );
  OAI22_X1 U11351 ( .A1(n10487), .A2(n10599), .B1(n10580), .B2(n10486), .ZN(
        n10488) );
  OAI21_X1 U11352 ( .B1(n10630), .B2(n10488), .A(n10600), .ZN(n10489) );
  OAI211_X1 U11353 ( .C1(n10634), .C2(n11254), .A(n10490), .B(n10489), .ZN(
        P1_U3267) );
  XNOR2_X1 U11354 ( .A(n10491), .B(n5513), .ZN(n10639) );
  INV_X1 U11355 ( .A(n10520), .ZN(n10494) );
  INV_X1 U11356 ( .A(n10492), .ZN(n10493) );
  AOI211_X1 U11357 ( .C1(n10637), .C2(n10494), .A(n10609), .B(n10493), .ZN(
        n10636) );
  NOR2_X1 U11358 ( .A1(n10495), .A2(n10534), .ZN(n10499) );
  OAI22_X1 U11359 ( .A1(n10600), .A2(n10497), .B1(n10496), .B2(n10580), .ZN(
        n10498) );
  AOI211_X1 U11360 ( .C1(n10636), .C2(n10560), .A(n10499), .B(n10498), .ZN(
        n10509) );
  AOI21_X1 U11361 ( .B1(n10501), .B2(n10500), .A(n5195), .ZN(n10502) );
  OAI222_X1 U11362 ( .A1(n10507), .A2(n10506), .B1(n10505), .B2(n10504), .C1(
        n10503), .C2(n10502), .ZN(n10635) );
  NAND2_X1 U11363 ( .A1(n10635), .A2(n10600), .ZN(n10508) );
  OAI211_X1 U11364 ( .C1(n10639), .C2(n11254), .A(n10509), .B(n10508), .ZN(
        P1_U3268) );
  NOR2_X1 U11365 ( .A1(n10535), .A2(n10510), .ZN(n10512) );
  XNOR2_X1 U11366 ( .A(n10512), .B(n10511), .ZN(n10514) );
  AOI222_X1 U11367 ( .A1(n11232), .A2(n10514), .B1(n10549), .B2(n11236), .C1(
        n10513), .C2(n11237), .ZN(n10644) );
  NAND2_X1 U11368 ( .A1(n10517), .A2(n10516), .ZN(n10640) );
  NAND3_X1 U11369 ( .A1(n10515), .A2(n11218), .A3(n10640), .ZN(n10527) );
  NAND2_X1 U11370 ( .A1(n10642), .A2(n10529), .ZN(n10518) );
  NAND2_X1 U11371 ( .A1(n10518), .A2(n11250), .ZN(n10519) );
  NOR2_X1 U11372 ( .A1(n10520), .A2(n10519), .ZN(n10641) );
  NAND2_X1 U11373 ( .A1(n10642), .A2(n11245), .ZN(n10524) );
  NOR2_X1 U11374 ( .A1(n10580), .A2(n10521), .ZN(n10522) );
  AOI21_X1 U11375 ( .B1(n11258), .B2(P1_REG2_REG_24__SCAN_IN), .A(n10522), 
        .ZN(n10523) );
  NAND2_X1 U11376 ( .A1(n10524), .A2(n10523), .ZN(n10525) );
  AOI21_X1 U11377 ( .B1(n10641), .B2(n10560), .A(n10525), .ZN(n10526) );
  OAI211_X1 U11378 ( .C1(n11258), .C2(n10644), .A(n10527), .B(n10526), .ZN(
        P1_U3269) );
  XOR2_X1 U11379 ( .A(n10528), .B(n10537), .Z(n10650) );
  INV_X1 U11380 ( .A(n10529), .ZN(n10530) );
  AOI21_X1 U11381 ( .B1(n10646), .B2(n5231), .A(n10530), .ZN(n10647) );
  INV_X1 U11382 ( .A(n10531), .ZN(n10532) );
  AOI22_X1 U11383 ( .A1(n11258), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10532), 
        .B2(n11243), .ZN(n10533) );
  OAI21_X1 U11384 ( .B1(n9318), .B2(n10534), .A(n10533), .ZN(n10544) );
  INV_X1 U11385 ( .A(n10535), .ZN(n10540) );
  NAND3_X1 U11386 ( .A1(n5261), .A2(n10538), .A3(n10537), .ZN(n10539) );
  NAND2_X1 U11387 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  AOI222_X1 U11388 ( .A1(n11232), .A2(n10542), .B1(n10541), .B2(n11237), .C1(
        n10570), .C2(n11236), .ZN(n10649) );
  NOR2_X1 U11389 ( .A1(n10649), .A2(n11244), .ZN(n10543) );
  AOI211_X1 U11390 ( .C1(n10647), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        n10546) );
  OAI21_X1 U11391 ( .B1(n10650), .B2(n11254), .A(n10546), .ZN(P1_U3270) );
  OAI21_X1 U11392 ( .B1(n10548), .B2(n10547), .A(n5261), .ZN(n10551) );
  AOI222_X1 U11393 ( .A1(n11232), .A2(n10551), .B1(n10550), .B2(n11236), .C1(
        n10549), .C2(n11237), .ZN(n10654) );
  OAI21_X1 U11394 ( .B1(n10554), .B2(n10553), .A(n10552), .ZN(n10555) );
  INV_X1 U11395 ( .A(n10555), .ZN(n10655) );
  NAND2_X1 U11396 ( .A1(n11258), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n10556) );
  OAI21_X1 U11397 ( .B1(n10580), .B2(n10557), .A(n10556), .ZN(n10558) );
  AOI21_X1 U11398 ( .B1(n10652), .B2(n11245), .A(n10558), .ZN(n10562) );
  AOI21_X1 U11399 ( .B1(n10652), .B2(n10576), .A(n10609), .ZN(n10559) );
  AND2_X1 U11400 ( .A1(n10559), .A2(n5231), .ZN(n10651) );
  NAND2_X1 U11401 ( .A1(n10651), .A2(n10560), .ZN(n10561) );
  OAI211_X1 U11402 ( .C1(n10655), .C2(n11254), .A(n10562), .B(n10561), .ZN(
        n10563) );
  INV_X1 U11403 ( .A(n10563), .ZN(n10564) );
  OAI21_X1 U11404 ( .B1(n11258), .B2(n10654), .A(n10564), .ZN(P1_U3271) );
  NAND2_X1 U11405 ( .A1(n10566), .A2(n10565), .ZN(n10568) );
  OAI21_X1 U11406 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(n10572) );
  AOI222_X1 U11407 ( .A1(n11232), .A2(n10572), .B1(n10571), .B2(n11236), .C1(
        n10570), .C2(n11237), .ZN(n10657) );
  AOI21_X1 U11408 ( .B1(n10575), .B2(n10574), .A(n10573), .ZN(n10660) );
  OAI211_X1 U11409 ( .C1(n10658), .C2(n10577), .A(n11250), .B(n10576), .ZN(
        n10656) );
  NAND2_X1 U11410 ( .A1(n11258), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n10578) );
  OAI21_X1 U11411 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(n10581) );
  AOI21_X1 U11412 ( .B1(n10582), .B2(n11245), .A(n10581), .ZN(n10583) );
  OAI21_X1 U11413 ( .B1(n10656), .B2(n11253), .A(n10583), .ZN(n10584) );
  AOI21_X1 U11414 ( .B1(n10660), .B2(n11218), .A(n10584), .ZN(n10585) );
  OAI21_X1 U11415 ( .B1(n11258), .B2(n10657), .A(n10585), .ZN(P1_U3272) );
  OAI21_X1 U11416 ( .B1(n10587), .B2(n10592), .A(n10586), .ZN(n10588) );
  INV_X1 U11417 ( .A(n10588), .ZN(n11227) );
  NAND2_X1 U11418 ( .A1(n11227), .A2(n11218), .ZN(n10606) );
  INV_X1 U11419 ( .A(n10589), .ZN(n10590) );
  AOI22_X1 U11420 ( .A1(n11244), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11243), 
        .B2(n10590), .ZN(n10605) );
  XNOR2_X1 U11421 ( .A(n10592), .B(n10591), .ZN(n10593) );
  NAND2_X1 U11422 ( .A1(n10593), .A2(n11232), .ZN(n10597) );
  AOI22_X1 U11423 ( .A1(n10595), .A2(n11237), .B1(n10594), .B2(n11236), .ZN(
        n10596) );
  NAND2_X1 U11424 ( .A1(n10597), .A2(n10596), .ZN(n11226) );
  INV_X1 U11425 ( .A(n10598), .ZN(n11205) );
  OAI211_X1 U11426 ( .C1(n11224), .C2(n10598), .A(n11250), .B(n11249), .ZN(
        n11223) );
  NOR2_X1 U11427 ( .A1(n11223), .A2(n10599), .ZN(n10601) );
  OAI21_X1 U11428 ( .B1(n11226), .B2(n10601), .A(n10600), .ZN(n10604) );
  NAND2_X1 U11429 ( .A1(n10602), .A2(n11245), .ZN(n10603) );
  NAND4_X1 U11430 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        P1_U3277) );
  NAND2_X1 U11431 ( .A1(n10607), .A2(n11111), .ZN(n10608) );
  OAI211_X1 U11432 ( .C1(n10610), .C2(n10609), .A(n10608), .B(n10611), .ZN(
        n10674) );
  MUX2_X1 U11433 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10674), .S(n11276), .Z(
        P1_U3553) );
  OAI211_X1 U11434 ( .C1(n5448), .C2(n11269), .A(n10612), .B(n10611), .ZN(
        n10675) );
  MUX2_X1 U11435 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10675), .S(n11276), .Z(
        P1_U3552) );
  AOI21_X1 U11436 ( .B1(n11111), .B2(n10614), .A(n10613), .ZN(n10616) );
  OAI211_X1 U11437 ( .C1(n10617), .C2(n10671), .A(n10616), .B(n10615), .ZN(
        n10676) );
  MUX2_X1 U11438 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10676), .S(n11276), .Z(
        P1_U3551) );
  NAND2_X1 U11439 ( .A1(n10618), .A2(n11111), .ZN(n10620) );
  OAI211_X1 U11440 ( .C1(n10621), .C2(n10671), .A(n10620), .B(n10619), .ZN(
        n10622) );
  INV_X1 U11441 ( .A(n10622), .ZN(n10624) );
  MUX2_X1 U11442 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10677), .S(n11276), .Z(
        P1_U3550) );
  AOI211_X1 U11443 ( .C1(n11111), .C2(n10627), .A(n10626), .B(n10625), .ZN(
        n10628) );
  OAI21_X1 U11444 ( .B1(n10629), .B2(n10671), .A(n10628), .ZN(n10678) );
  MUX2_X1 U11445 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10678), .S(n11276), .Z(
        P1_U3549) );
  AOI211_X1 U11446 ( .C1(n11111), .C2(n10632), .A(n10631), .B(n10630), .ZN(
        n10633) );
  OAI21_X1 U11447 ( .B1(n10634), .B2(n10671), .A(n10633), .ZN(n10679) );
  MUX2_X1 U11448 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10679), .S(n11276), .Z(
        P1_U3548) );
  AOI211_X1 U11449 ( .C1(n11111), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10638) );
  OAI21_X1 U11450 ( .B1(n10639), .B2(n10671), .A(n10638), .ZN(n10680) );
  MUX2_X1 U11451 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10680), .S(n11276), .Z(
        P1_U3547) );
  NAND2_X1 U11452 ( .A1(n10640), .A2(n11273), .ZN(n10645) );
  AOI21_X1 U11453 ( .B1(n11111), .B2(n10642), .A(n10641), .ZN(n10643) );
  OAI211_X1 U11454 ( .C1(n5638), .C2(n10645), .A(n10644), .B(n10643), .ZN(
        n10681) );
  MUX2_X1 U11455 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10681), .S(n11276), .Z(
        P1_U3546) );
  AOI22_X1 U11456 ( .A1(n10647), .A2(n11250), .B1(n11111), .B2(n10646), .ZN(
        n10648) );
  OAI211_X1 U11457 ( .C1(n10650), .C2(n10671), .A(n10649), .B(n10648), .ZN(
        n10682) );
  MUX2_X1 U11458 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10682), .S(n11276), .Z(
        P1_U3545) );
  AOI21_X1 U11459 ( .B1(n11111), .B2(n10652), .A(n10651), .ZN(n10653) );
  OAI211_X1 U11460 ( .C1(n10655), .C2(n10671), .A(n10654), .B(n10653), .ZN(
        n10683) );
  MUX2_X1 U11461 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10683), .S(n11276), .Z(
        P1_U3544) );
  OAI211_X1 U11462 ( .C1(n10658), .C2(n11269), .A(n10657), .B(n10656), .ZN(
        n10659) );
  AOI21_X1 U11463 ( .B1(n10660), .B2(n11273), .A(n10659), .ZN(n10661) );
  INV_X1 U11464 ( .A(n10661), .ZN(n10684) );
  MUX2_X1 U11465 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10684), .S(n11276), .Z(
        P1_U3543) );
  AOI211_X1 U11466 ( .C1(n11111), .C2(n10664), .A(n10663), .B(n10662), .ZN(
        n10665) );
  OAI21_X1 U11467 ( .B1(n10666), .B2(n10671), .A(n10665), .ZN(n10685) );
  MUX2_X1 U11468 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10685), .S(n11276), .Z(
        P1_U3542) );
  AOI211_X1 U11469 ( .C1(n11111), .C2(n10669), .A(n10668), .B(n10667), .ZN(
        n10670) );
  OAI21_X1 U11470 ( .B1(n10672), .B2(n10671), .A(n10670), .ZN(n10686) );
  MUX2_X1 U11471 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10686), .S(n11276), .Z(
        P1_U3541) );
  MUX2_X1 U11472 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10673), .S(n11276), .Z(
        P1_U3522) );
  MUX2_X1 U11473 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10674), .S(n11280), .Z(
        P1_U3521) );
  MUX2_X1 U11474 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10675), .S(n11280), .Z(
        P1_U3520) );
  MUX2_X1 U11475 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10676), .S(n11280), .Z(
        P1_U3519) );
  MUX2_X1 U11476 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10677), .S(n11280), .Z(
        P1_U3518) );
  MUX2_X1 U11477 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10678), .S(n11280), .Z(
        P1_U3517) );
  MUX2_X1 U11478 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10679), .S(n11280), .Z(
        P1_U3516) );
  MUX2_X1 U11479 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10680), .S(n11280), .Z(
        P1_U3515) );
  MUX2_X1 U11480 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10681), .S(n11280), .Z(
        P1_U3514) );
  MUX2_X1 U11481 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10682), .S(n11280), .Z(
        P1_U3513) );
  MUX2_X1 U11482 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10683), .S(n11280), .Z(
        P1_U3512) );
  MUX2_X1 U11483 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10684), .S(n11280), .Z(
        P1_U3511) );
  MUX2_X1 U11484 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10685), .S(n11280), .Z(
        P1_U3510) );
  MUX2_X1 U11485 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10686), .S(n11280), .Z(
        P1_U3509) );
  MUX2_X1 U11486 ( .A(n10687), .B(P1_D_REG_1__SCAN_IN), .S(n10704), .Z(
        P1_U3440) );
  NAND3_X1 U11487 ( .A1(n10688), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10690) );
  OAI22_X1 U11488 ( .A1(n10691), .A2(n10690), .B1(n10689), .B2(n10696), .ZN(
        n10692) );
  AOI21_X1 U11489 ( .B1(n10694), .B2(n10693), .A(n10692), .ZN(n10695) );
  INV_X1 U11490 ( .A(n10695), .ZN(P1_U3324) );
  OAI222_X1 U11491 ( .A1(n9271), .A2(n10699), .B1(n10698), .B2(P1_U3086), .C1(
        n10697), .C2(n10696), .ZN(P1_U3326) );
  MUX2_X1 U11492 ( .A(n10700), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11493 ( .A1(n10704), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3323) );
  INV_X1 U11494 ( .A(n10704), .ZN(n10703) );
  NOR2_X1 U11495 ( .A1(n10703), .A2(n10701), .ZN(P1_U3322) );
  AND2_X1 U11496 ( .A1(n10704), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U11497 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10702) );
  NOR2_X1 U11498 ( .A1(n10703), .A2(n10702), .ZN(P1_U3320) );
  AND2_X1 U11499 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10704), .ZN(P1_U3319) );
  AND2_X1 U11500 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10704), .ZN(P1_U3318) );
  AND2_X1 U11501 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10704), .ZN(P1_U3317) );
  AND2_X1 U11502 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10704), .ZN(P1_U3316) );
  AND2_X1 U11503 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10704), .ZN(P1_U3315) );
  AND2_X1 U11504 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10704), .ZN(P1_U3314) );
  AND2_X1 U11505 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10704), .ZN(P1_U3313) );
  AND2_X1 U11506 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10704), .ZN(P1_U3312) );
  AND2_X1 U11507 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10704), .ZN(P1_U3311) );
  AND2_X1 U11508 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10704), .ZN(P1_U3310) );
  AND2_X1 U11509 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10704), .ZN(P1_U3309) );
  AND2_X1 U11510 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10704), .ZN(P1_U3308) );
  AND2_X1 U11511 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10704), .ZN(P1_U3307) );
  AND2_X1 U11512 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10704), .ZN(P1_U3306) );
  AND2_X1 U11513 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10704), .ZN(P1_U3305) );
  AND2_X1 U11514 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10704), .ZN(P1_U3304) );
  AND2_X1 U11515 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10704), .ZN(P1_U3303) );
  AND2_X1 U11516 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10704), .ZN(P1_U3302) );
  AND2_X1 U11517 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10704), .ZN(P1_U3301) );
  AND2_X1 U11518 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10704), .ZN(P1_U3300) );
  AND2_X1 U11519 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10704), .ZN(P1_U3299) );
  AND2_X1 U11520 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10704), .ZN(P1_U3298) );
  AND2_X1 U11521 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10704), .ZN(P1_U3297) );
  AND2_X1 U11522 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10704), .ZN(P1_U3296) );
  AND2_X1 U11523 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10704), .ZN(P1_U3295) );
  AND2_X1 U11524 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10704), .ZN(P1_U3294) );
  OAI21_X1 U11525 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10707), .ZN(n10705) );
  INV_X1 U11526 ( .A(n10705), .ZN(ADD_1068_U46) );
  OAI21_X1 U11527 ( .B1(n10708), .B2(n10707), .A(n10706), .ZN(n10709) );
  XNOR2_X1 U11528 ( .A(n10709), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  AOI21_X1 U11529 ( .B1(n10712), .B2(n10711), .A(n10710), .ZN(ADD_1068_U54) );
  AOI21_X1 U11530 ( .B1(n10715), .B2(n10714), .A(n10713), .ZN(ADD_1068_U53) );
  OAI21_X1 U11531 ( .B1(n10718), .B2(n10717), .A(n10716), .ZN(ADD_1068_U52) );
  OAI21_X1 U11532 ( .B1(n10721), .B2(n10720), .A(n10719), .ZN(ADD_1068_U51) );
  OAI21_X1 U11533 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(ADD_1068_U50) );
  OAI21_X1 U11534 ( .B1(n10727), .B2(n10726), .A(n10725), .ZN(ADD_1068_U49) );
  OAI21_X1 U11535 ( .B1(n10730), .B2(n10729), .A(n10728), .ZN(ADD_1068_U48) );
  OAI21_X1 U11536 ( .B1(n10733), .B2(n10732), .A(n10731), .ZN(ADD_1068_U47) );
  OAI21_X1 U11537 ( .B1(n10736), .B2(n10735), .A(n10734), .ZN(ADD_1068_U63) );
  OAI21_X1 U11538 ( .B1(n10739), .B2(n10738), .A(n10737), .ZN(ADD_1068_U62) );
  OAI21_X1 U11539 ( .B1(n10742), .B2(n10741), .A(n10740), .ZN(ADD_1068_U61) );
  OAI21_X1 U11540 ( .B1(n10745), .B2(n10744), .A(n10743), .ZN(ADD_1068_U60) );
  OAI21_X1 U11541 ( .B1(n10748), .B2(n10747), .A(n10746), .ZN(ADD_1068_U59) );
  OAI21_X1 U11542 ( .B1(n10751), .B2(n10750), .A(n10749), .ZN(ADD_1068_U58) );
  OAI21_X1 U11543 ( .B1(n10754), .B2(n10753), .A(n10752), .ZN(ADD_1068_U57) );
  OAI21_X1 U11544 ( .B1(n10757), .B2(n10756), .A(n10755), .ZN(ADD_1068_U56) );
  OAI21_X1 U11545 ( .B1(n10760), .B2(n10759), .A(n10758), .ZN(ADD_1068_U55) );
  INV_X1 U11546 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10775) );
  OAI21_X1 U11547 ( .B1(n10763), .B2(n10762), .A(n10761), .ZN(n10771) );
  NAND2_X1 U11548 ( .A1(n10929), .A2(n10764), .ZN(n10770) );
  OAI21_X1 U11549 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(n10768) );
  OR2_X1 U11550 ( .A1(n10918), .A2(n10768), .ZN(n10769) );
  OAI211_X1 U11551 ( .C1(n10922), .C2(n10771), .A(n10770), .B(n10769), .ZN(
        n10772) );
  INV_X1 U11552 ( .A(n10772), .ZN(n10774) );
  OAI211_X1 U11553 ( .C1(n10933), .C2(n10775), .A(n10774), .B(n10773), .ZN(
        P1_U3248) );
  INV_X1 U11554 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U11555 ( .A1(n10777), .A2(n10776), .ZN(n10780) );
  INV_X1 U11556 ( .A(n10778), .ZN(n10779) );
  NAND3_X1 U11557 ( .A1(n10895), .A2(n10780), .A3(n10779), .ZN(n10788) );
  INV_X1 U11558 ( .A(n10781), .ZN(n10782) );
  OAI211_X1 U11559 ( .C1(n10784), .C2(n10783), .A(n10846), .B(n10782), .ZN(
        n10787) );
  NAND2_X1 U11560 ( .A1(n10929), .A2(n10785), .ZN(n10786) );
  AND3_X1 U11561 ( .A1(n10788), .A2(n10787), .A3(n10786), .ZN(n10790) );
  OAI211_X1 U11562 ( .C1(n10933), .C2(n10791), .A(n10790), .B(n10789), .ZN(
        P1_U3249) );
  INV_X1 U11563 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10803) );
  AOI211_X1 U11564 ( .C1(n10794), .C2(n10793), .A(n10792), .B(n10918), .ZN(
        n10799) );
  AOI211_X1 U11565 ( .C1(n10797), .C2(n10796), .A(n10795), .B(n10922), .ZN(
        n10798) );
  AOI211_X1 U11566 ( .C1(n10929), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10802) );
  OAI211_X1 U11567 ( .C1(n10933), .C2(n10803), .A(n10802), .B(n10801), .ZN(
        P1_U3250) );
  INV_X1 U11568 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U11569 ( .A1(n10805), .A2(n10804), .ZN(n10808) );
  INV_X1 U11570 ( .A(n10806), .ZN(n10807) );
  NAND2_X1 U11571 ( .A1(n10808), .A2(n10807), .ZN(n10816) );
  AOI21_X1 U11572 ( .B1(n10811), .B2(n10810), .A(n10809), .ZN(n10812) );
  NAND2_X1 U11573 ( .A1(n10846), .A2(n10812), .ZN(n10815) );
  NAND2_X1 U11574 ( .A1(n10929), .A2(n10813), .ZN(n10814) );
  OAI211_X1 U11575 ( .C1(n10816), .C2(n10922), .A(n10815), .B(n10814), .ZN(
        n10817) );
  INV_X1 U11576 ( .A(n10817), .ZN(n10819) );
  OAI211_X1 U11577 ( .C1(n10933), .C2(n10820), .A(n10819), .B(n10818), .ZN(
        P1_U3251) );
  INV_X1 U11578 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U11579 ( .A1(n10822), .A2(n10821), .ZN(n10825) );
  INV_X1 U11580 ( .A(n10823), .ZN(n10824) );
  NAND3_X1 U11581 ( .A1(n10895), .A2(n10825), .A3(n10824), .ZN(n10834) );
  NAND2_X1 U11582 ( .A1(n10929), .A2(n10826), .ZN(n10833) );
  NAND2_X1 U11583 ( .A1(n10828), .A2(n10827), .ZN(n10831) );
  INV_X1 U11584 ( .A(n10829), .ZN(n10830) );
  NAND3_X1 U11585 ( .A1(n10846), .A2(n10831), .A3(n10830), .ZN(n10832) );
  AND3_X1 U11586 ( .A1(n10834), .A2(n10833), .A3(n10832), .ZN(n10836) );
  OAI211_X1 U11587 ( .C1(n10933), .C2(n10837), .A(n10836), .B(n10835), .ZN(
        P1_U3254) );
  INV_X1 U11588 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10854) );
  NAND2_X1 U11589 ( .A1(n10839), .A2(n10838), .ZN(n10840) );
  NAND2_X1 U11590 ( .A1(n10841), .A2(n10840), .ZN(n10850) );
  AOI21_X1 U11591 ( .B1(n10844), .B2(n10843), .A(n10842), .ZN(n10845) );
  NAND2_X1 U11592 ( .A1(n10846), .A2(n10845), .ZN(n10849) );
  NAND2_X1 U11593 ( .A1(n10929), .A2(n10847), .ZN(n10848) );
  OAI211_X1 U11594 ( .C1(n10850), .C2(n10922), .A(n10849), .B(n10848), .ZN(
        n10851) );
  INV_X1 U11595 ( .A(n10851), .ZN(n10853) );
  OAI211_X1 U11596 ( .C1(n10933), .C2(n10854), .A(n10853), .B(n10852), .ZN(
        P1_U3257) );
  INV_X1 U11597 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U11598 ( .A1(n10855), .A2(n6593), .ZN(n10858) );
  INV_X1 U11599 ( .A(n10856), .ZN(n10857) );
  NAND2_X1 U11600 ( .A1(n10858), .A2(n10857), .ZN(n10867) );
  NAND2_X1 U11601 ( .A1(n10929), .A2(n10859), .ZN(n10866) );
  INV_X1 U11602 ( .A(n10860), .ZN(n10863) );
  NAND2_X1 U11603 ( .A1(n10861), .A2(n6592), .ZN(n10862) );
  NAND2_X1 U11604 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  OR2_X1 U11605 ( .A1(n10918), .A2(n10864), .ZN(n10865) );
  OAI211_X1 U11606 ( .C1(n10922), .C2(n10867), .A(n10866), .B(n10865), .ZN(
        n10868) );
  INV_X1 U11607 ( .A(n10868), .ZN(n10871) );
  INV_X1 U11608 ( .A(n10869), .ZN(n10870) );
  OAI211_X1 U11609 ( .C1(n10933), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        P1_U3258) );
  NAND2_X1 U11610 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  AND2_X1 U11611 ( .A1(n10876), .A2(n10875), .ZN(n10885) );
  NAND2_X1 U11612 ( .A1(n10929), .A2(n10877), .ZN(n10884) );
  OAI21_X1 U11613 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(n10881) );
  INV_X1 U11614 ( .A(n10881), .ZN(n10882) );
  OR2_X1 U11615 ( .A1(n10918), .A2(n10882), .ZN(n10883) );
  OAI211_X1 U11616 ( .C1(n10922), .C2(n10885), .A(n10884), .B(n10883), .ZN(
        n10886) );
  INV_X1 U11617 ( .A(n10886), .ZN(n10888) );
  OAI211_X1 U11618 ( .C1(n10933), .C2(n10889), .A(n10888), .B(n10887), .ZN(
        P1_U3260) );
  INV_X1 U11619 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10905) );
  OAI21_X1 U11620 ( .B1(n10892), .B2(n10891), .A(n10890), .ZN(n10901) );
  INV_X1 U11621 ( .A(n10893), .ZN(n10897) );
  OAI211_X1 U11622 ( .C1(n10897), .C2(n10896), .A(n10895), .B(n10894), .ZN(
        n10900) );
  NAND2_X1 U11623 ( .A1(n10929), .A2(n10898), .ZN(n10899) );
  OAI211_X1 U11624 ( .C1(n10918), .C2(n10901), .A(n10900), .B(n10899), .ZN(
        n10902) );
  INV_X1 U11625 ( .A(n10902), .ZN(n10904) );
  OAI211_X1 U11626 ( .C1(n10933), .C2(n10905), .A(n10904), .B(n10903), .ZN(
        P1_U3261) );
  INV_X1 U11627 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10917) );
  AOI211_X1 U11628 ( .C1(n10908), .C2(n10907), .A(n10906), .B(n10918), .ZN(
        n10913) );
  AOI211_X1 U11629 ( .C1(n10911), .C2(n10910), .A(n10909), .B(n10922), .ZN(
        n10912) );
  AOI211_X1 U11630 ( .C1(n10914), .C2(n10929), .A(n10913), .B(n10912), .ZN(
        n10916) );
  OAI211_X1 U11631 ( .C1(n10933), .C2(n10917), .A(n10916), .B(n10915), .ZN(
        P1_U3256) );
  INV_X1 U11632 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10932) );
  AOI211_X1 U11633 ( .C1(n10921), .C2(n10920), .A(n10919), .B(n10918), .ZN(
        n10927) );
  AOI211_X1 U11634 ( .C1(n10925), .C2(n10924), .A(n10923), .B(n10922), .ZN(
        n10926) );
  AOI211_X1 U11635 ( .C1(n10929), .C2(n10928), .A(n10927), .B(n10926), .ZN(
        n10931) );
  OAI211_X1 U11636 ( .C1(n10933), .C2(n10932), .A(n10931), .B(n10930), .ZN(
        P1_U3253) );
  INV_X1 U11637 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11009) );
  AOI21_X1 U11638 ( .B1(n10936), .B2(n10935), .A(n10934), .ZN(n10937) );
  NOR2_X1 U11639 ( .A1(n10967), .A2(n10937), .ZN(n10943) );
  AOI211_X1 U11640 ( .C1(n10941), .C2(n10940), .A(n10939), .B(n10938), .ZN(
        n10942) );
  AOI211_X1 U11641 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n10959), .A(n10943), .B(
        n10942), .ZN(n10944) );
  OAI21_X1 U11642 ( .B1(n10945), .B2(n5947), .A(n10944), .ZN(n10946) );
  INV_X1 U11643 ( .A(n10946), .ZN(n10952) );
  OAI21_X1 U11644 ( .B1(n10949), .B2(n10948), .A(n10947), .ZN(n10950) );
  NAND2_X1 U11645 ( .A1(n5906), .A2(n10950), .ZN(n10951) );
  OAI211_X1 U11646 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n11009), .A(n10952), .B(
        n10951), .ZN(P2_U3184) );
  INV_X1 U11647 ( .A(n10953), .ZN(n10955) );
  NAND2_X1 U11648 ( .A1(n10955), .A2(n10954), .ZN(n10960) );
  AND3_X1 U11649 ( .A1(n10960), .A2(n5272), .A3(n10956), .ZN(n10957) );
  AOI211_X1 U11650 ( .C1(n10959), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n10958), 
        .B(n10957), .ZN(n10977) );
  OAI21_X1 U11651 ( .B1(n10961), .B2(n10960), .A(n5947), .ZN(n10963) );
  NAND2_X1 U11652 ( .A1(n10963), .A2(n10962), .ZN(n10976) );
  AOI21_X1 U11653 ( .B1(n10966), .B2(n10965), .A(n10964), .ZN(n10968) );
  OR2_X1 U11654 ( .A1(n10968), .A2(n10967), .ZN(n10975) );
  AOI21_X1 U11655 ( .B1(n10971), .B2(n10970), .A(n10969), .ZN(n10973) );
  OR2_X1 U11656 ( .A1(n10973), .A2(n10972), .ZN(n10974) );
  NAND4_X1 U11657 ( .A1(n10977), .A2(n10976), .A3(n10975), .A4(n10974), .ZN(
        P2_U3200) );
  AOI22_X1 U11658 ( .A1(n11159), .A2(n10979), .B1(n10978), .B2(n11158), .ZN(
        n10980) );
  AND2_X1 U11659 ( .A1(n10981), .A2(n10980), .ZN(n10984) );
  AOI22_X1 U11660 ( .A1(n11187), .A2(n10984), .B1(n10982), .B2(n11185), .ZN(
        P2_U3460) );
  INV_X1 U11661 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U11662 ( .A1(n11191), .A2(n10984), .B1(n10983), .B2(n11188), .ZN(
        P2_U3393) );
  INV_X1 U11663 ( .A(n11069), .ZN(n11197) );
  INV_X1 U11664 ( .A(n10985), .ZN(n10986) );
  OAI21_X1 U11665 ( .B1(n10987), .B2(n11269), .A(n10986), .ZN(n10989) );
  AOI211_X1 U11666 ( .C1(n11197), .C2(n10990), .A(n10989), .B(n10988), .ZN(
        n10992) );
  AOI22_X1 U11667 ( .A1(n11276), .A2(n10992), .B1(n10991), .B2(n11275), .ZN(
        P1_U3523) );
  AOI22_X1 U11668 ( .A1(n11280), .A2(n10992), .B1(n6612), .B2(n11277), .ZN(
        P1_U3456) );
  MUX2_X1 U11669 ( .A(n10993), .B(P1_REG0_REG_2__SCAN_IN), .S(n11277), .Z(
        P1_U3459) );
  OAI21_X1 U11670 ( .B1(n10994), .B2(n10996), .A(n8233), .ZN(n11013) );
  NOR2_X1 U11671 ( .A1(n11179), .A2(n11008), .ZN(n11004) );
  NAND3_X1 U11672 ( .A1(n8388), .A2(n10996), .A3(n10995), .ZN(n10997) );
  AND2_X1 U11673 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  OAI222_X1 U11674 ( .A1(n11003), .A2(n11002), .B1(n11001), .B2(n6102), .C1(
        n11000), .C2(n10999), .ZN(n11011) );
  AOI211_X1 U11675 ( .C1(n11159), .C2(n11013), .A(n11004), .B(n11011), .ZN(
        n11006) );
  AOI22_X1 U11676 ( .A1(n11187), .A2(n11006), .B1(n5824), .B2(n11185), .ZN(
        P2_U3461) );
  INV_X1 U11677 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U11678 ( .A1(n11191), .A2(n11006), .B1(n11005), .B2(n11188), .ZN(
        P2_U3396) );
  OAI22_X1 U11679 ( .A1(n11010), .A2(n11009), .B1(n11008), .B2(n11007), .ZN(
        n11012) );
  AOI211_X1 U11680 ( .C1(n11014), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11016) );
  AOI22_X1 U11681 ( .A1(n11018), .A2(n11017), .B1(n11016), .B2(n11015), .ZN(
        P2_U3231) );
  OAI21_X1 U11682 ( .B1(n11020), .B2(n11269), .A(n11019), .ZN(n11022) );
  AOI211_X1 U11683 ( .C1(n11197), .C2(n11023), .A(n11022), .B(n11021), .ZN(
        n11025) );
  AOI22_X1 U11684 ( .A1(n11276), .A2(n11025), .B1(n6636), .B2(n11275), .ZN(
        P1_U3525) );
  INV_X1 U11685 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U11686 ( .A1(n11280), .A2(n11025), .B1(n11024), .B2(n11277), .ZN(
        P1_U3462) );
  INV_X1 U11687 ( .A(n11026), .ZN(n11030) );
  OAI22_X1 U11688 ( .A1(n11028), .A2(n11181), .B1(n11027), .B2(n11179), .ZN(
        n11029) );
  NOR2_X1 U11689 ( .A1(n11030), .A2(n11029), .ZN(n11033) );
  INV_X1 U11690 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U11691 ( .A1(n11187), .A2(n11033), .B1(n11031), .B2(n11185), .ZN(
        P2_U3462) );
  INV_X1 U11692 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U11693 ( .A1(n11191), .A2(n11033), .B1(n11032), .B2(n11188), .ZN(
        P2_U3399) );
  INV_X1 U11694 ( .A(n11034), .ZN(n11038) );
  OAI22_X1 U11695 ( .A1(n11036), .A2(n11181), .B1(n11035), .B2(n11179), .ZN(
        n11037) );
  NOR2_X1 U11696 ( .A1(n11038), .A2(n11037), .ZN(n11040) );
  AOI22_X1 U11697 ( .A1(n11187), .A2(n11040), .B1(n5829), .B2(n11185), .ZN(
        P2_U3463) );
  INV_X1 U11698 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U11699 ( .A1(n11191), .A2(n11040), .B1(n11039), .B2(n11188), .ZN(
        P2_U3402) );
  OAI211_X1 U11700 ( .C1(n11043), .C2(n11269), .A(n11042), .B(n11041), .ZN(
        n11044) );
  AOI21_X1 U11701 ( .B1(n11273), .B2(n11045), .A(n11044), .ZN(n11047) );
  AOI22_X1 U11702 ( .A1(n11276), .A2(n11047), .B1(n6650), .B2(n11275), .ZN(
        P1_U3526) );
  INV_X1 U11703 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U11704 ( .A1(n11280), .A2(n11047), .B1(n11046), .B2(n11277), .ZN(
        P1_U3465) );
  OAI22_X1 U11705 ( .A1(n11049), .A2(n11181), .B1(n11048), .B2(n11179), .ZN(
        n11050) );
  NOR2_X1 U11706 ( .A1(n11051), .A2(n11050), .ZN(n11054) );
  INV_X1 U11707 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U11708 ( .A1(n11187), .A2(n11054), .B1(n11052), .B2(n11185), .ZN(
        P2_U3464) );
  INV_X1 U11709 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U11710 ( .A1(n11191), .A2(n11054), .B1(n11053), .B2(n11188), .ZN(
        P2_U3405) );
  OAI21_X1 U11711 ( .B1(n11056), .B2(n11269), .A(n11055), .ZN(n11058) );
  AOI211_X1 U11712 ( .C1(n11273), .C2(n11059), .A(n11058), .B(n11057), .ZN(
        n11061) );
  AOI22_X1 U11713 ( .A1(n11276), .A2(n11061), .B1(n6669), .B2(n11275), .ZN(
        P1_U3527) );
  INV_X1 U11714 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U11715 ( .A1(n11280), .A2(n11061), .B1(n11060), .B2(n11277), .ZN(
        P1_U3468) );
  INV_X1 U11716 ( .A(n11062), .ZN(n11066) );
  OAI22_X1 U11717 ( .A1(n11064), .A2(n11181), .B1(n11063), .B2(n11179), .ZN(
        n11065) );
  NOR2_X1 U11718 ( .A1(n11066), .A2(n11065), .ZN(n11068) );
  AOI22_X1 U11719 ( .A1(n11187), .A2(n11068), .B1(n5832), .B2(n11185), .ZN(
        P2_U3465) );
  INV_X1 U11720 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U11721 ( .A1(n11191), .A2(n11068), .B1(n11067), .B2(n11188), .ZN(
        P2_U3408) );
  INV_X1 U11722 ( .A(n11070), .ZN(n11076) );
  NOR2_X1 U11723 ( .A1(n11070), .A2(n11069), .ZN(n11075) );
  OAI211_X1 U11724 ( .C1(n11073), .C2(n11269), .A(n11072), .B(n11071), .ZN(
        n11074) );
  AOI211_X1 U11725 ( .C1(n11077), .C2(n11076), .A(n11075), .B(n11074), .ZN(
        n11079) );
  AOI22_X1 U11726 ( .A1(n11276), .A2(n11079), .B1(n6678), .B2(n11275), .ZN(
        P1_U3528) );
  INV_X1 U11727 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U11728 ( .A1(n11280), .A2(n11079), .B1(n11078), .B2(n11277), .ZN(
        P1_U3471) );
  OAI211_X1 U11729 ( .C1(n11082), .C2(n11269), .A(n11081), .B(n11080), .ZN(
        n11083) );
  AOI21_X1 U11730 ( .B1(n11273), .B2(n11084), .A(n11083), .ZN(n11086) );
  AOI22_X1 U11731 ( .A1(n11276), .A2(n11086), .B1(n6695), .B2(n11275), .ZN(
        P1_U3529) );
  INV_X1 U11732 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U11733 ( .A1(n11280), .A2(n11086), .B1(n11085), .B2(n11277), .ZN(
        P1_U3474) );
  OAI22_X1 U11734 ( .A1(n11088), .A2(n11181), .B1(n11087), .B2(n11179), .ZN(
        n11089) );
  NOR2_X1 U11735 ( .A1(n11090), .A2(n11089), .ZN(n11093) );
  AOI22_X1 U11736 ( .A1(n11187), .A2(n11093), .B1(n11091), .B2(n11185), .ZN(
        P2_U3466) );
  INV_X1 U11737 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U11738 ( .A1(n11191), .A2(n11093), .B1(n11092), .B2(n11188), .ZN(
        P2_U3411) );
  INV_X1 U11739 ( .A(n11094), .ZN(n11099) );
  OAI21_X1 U11740 ( .B1(n11096), .B2(n11269), .A(n11095), .ZN(n11098) );
  AOI211_X1 U11741 ( .C1(n11197), .C2(n11099), .A(n11098), .B(n11097), .ZN(
        n11101) );
  AOI22_X1 U11742 ( .A1(n11276), .A2(n11101), .B1(n6715), .B2(n11275), .ZN(
        P1_U3530) );
  INV_X1 U11743 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11744 ( .A1(n11280), .A2(n11101), .B1(n11100), .B2(n11277), .ZN(
        P1_U3477) );
  INV_X1 U11745 ( .A(n11102), .ZN(n11106) );
  OAI21_X1 U11746 ( .B1(n11104), .B2(n11179), .A(n11103), .ZN(n11105) );
  AOI21_X1 U11747 ( .B1(n11159), .B2(n11106), .A(n11105), .ZN(n11109) );
  INV_X1 U11748 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U11749 ( .A1(n11187), .A2(n11109), .B1(n11107), .B2(n11185), .ZN(
        P2_U3467) );
  INV_X1 U11750 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U11751 ( .A1(n11191), .A2(n11109), .B1(n11108), .B2(n11188), .ZN(
        P2_U3414) );
  AND2_X1 U11752 ( .A1(n11110), .A2(n11273), .ZN(n11116) );
  AND2_X1 U11753 ( .A1(n11112), .A2(n11111), .ZN(n11113) );
  OR2_X1 U11754 ( .A1(n11114), .A2(n11113), .ZN(n11115) );
  NOR3_X1 U11755 ( .A1(n11117), .A2(n11116), .A3(n11115), .ZN(n11119) );
  AOI22_X1 U11756 ( .A1(n11276), .A2(n11119), .B1(n6727), .B2(n11275), .ZN(
        P1_U3531) );
  INV_X1 U11757 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U11758 ( .A1(n11280), .A2(n11119), .B1(n11118), .B2(n11277), .ZN(
        P1_U3480) );
  NOR2_X1 U11759 ( .A1(n11120), .A2(n11181), .ZN(n11122) );
  AOI211_X1 U11760 ( .C1(n11158), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n11126) );
  AOI22_X1 U11761 ( .A1(n11187), .A2(n11126), .B1(n11124), .B2(n11185), .ZN(
        P2_U3468) );
  INV_X1 U11762 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U11763 ( .A1(n11191), .A2(n11126), .B1(n11125), .B2(n11188), .ZN(
        P2_U3417) );
  OAI21_X1 U11764 ( .B1(n11128), .B2(n11269), .A(n11127), .ZN(n11129) );
  AOI211_X1 U11765 ( .C1(n11131), .C2(n11273), .A(n11130), .B(n11129), .ZN(
        n11133) );
  INV_X1 U11766 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U11767 ( .A1(n11276), .A2(n11133), .B1(n11132), .B2(n11275), .ZN(
        P1_U3532) );
  AOI22_X1 U11768 ( .A1(n11280), .A2(n11133), .B1(n6746), .B2(n11277), .ZN(
        P1_U3483) );
  INV_X1 U11769 ( .A(n11134), .ZN(n11136) );
  NOR2_X1 U11770 ( .A1(n11136), .A2(n11135), .ZN(n11138) );
  AOI211_X1 U11771 ( .C1(n11158), .C2(n11139), .A(n11138), .B(n11137), .ZN(
        n11142) );
  INV_X1 U11772 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U11773 ( .A1(n11187), .A2(n11142), .B1(n11140), .B2(n11185), .ZN(
        P2_U3469) );
  INV_X1 U11774 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U11775 ( .A1(n11191), .A2(n11142), .B1(n11141), .B2(n11188), .ZN(
        P2_U3420) );
  AOI22_X1 U11776 ( .A1(n11144), .A2(n11159), .B1(n11158), .B2(n11143), .ZN(
        n11146) );
  AND2_X1 U11777 ( .A1(n11146), .A2(n11145), .ZN(n11149) );
  AOI22_X1 U11778 ( .A1(n11187), .A2(n11149), .B1(n11147), .B2(n11185), .ZN(
        P2_U3470) );
  INV_X1 U11779 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U11780 ( .A1(n11191), .A2(n11149), .B1(n11148), .B2(n11188), .ZN(
        P2_U3423) );
  OAI211_X1 U11781 ( .C1(n11152), .C2(n11269), .A(n11151), .B(n11150), .ZN(
        n11153) );
  AOI21_X1 U11782 ( .B1(n11273), .B2(n11154), .A(n11153), .ZN(n11156) );
  AOI22_X1 U11783 ( .A1(n11276), .A2(n11156), .B1(n7860), .B2(n11275), .ZN(
        P1_U3533) );
  INV_X1 U11784 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11155) );
  AOI22_X1 U11785 ( .A1(n11280), .A2(n11156), .B1(n11155), .B2(n11277), .ZN(
        P1_U3486) );
  AOI22_X1 U11786 ( .A1(n11160), .A2(n11159), .B1(n11158), .B2(n11157), .ZN(
        n11162) );
  AND2_X1 U11787 ( .A1(n11162), .A2(n11161), .ZN(n11165) );
  AOI22_X1 U11788 ( .A1(n11187), .A2(n11165), .B1(n11163), .B2(n11185), .ZN(
        P2_U3471) );
  INV_X1 U11789 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U11790 ( .A1(n11191), .A2(n11165), .B1(n11164), .B2(n11188), .ZN(
        P2_U3426) );
  OAI211_X1 U11791 ( .C1(n11168), .C2(n11269), .A(n11167), .B(n11166), .ZN(
        n11169) );
  AOI21_X1 U11792 ( .B1(n11273), .B2(n11170), .A(n11169), .ZN(n11172) );
  AOI22_X1 U11793 ( .A1(n11276), .A2(n11172), .B1(n6771), .B2(n11275), .ZN(
        P1_U3534) );
  INV_X1 U11794 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U11795 ( .A1(n11280), .A2(n11172), .B1(n11171), .B2(n11277), .ZN(
        P1_U3489) );
  OAI211_X1 U11796 ( .C1(n5417), .C2(n11269), .A(n11174), .B(n11173), .ZN(
        n11175) );
  AOI21_X1 U11797 ( .B1(n11273), .B2(n11176), .A(n11175), .ZN(n11178) );
  AOI22_X1 U11798 ( .A1(n11276), .A2(n11178), .B1(n10377), .B2(n11275), .ZN(
        P1_U3535) );
  INV_X1 U11799 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U11800 ( .A1(n11280), .A2(n11178), .B1(n11177), .B2(n11277), .ZN(
        P1_U3492) );
  OAI22_X1 U11801 ( .A1(n11182), .A2(n11181), .B1(n11180), .B2(n11179), .ZN(
        n11183) );
  NOR2_X1 U11802 ( .A1(n11184), .A2(n11183), .ZN(n11190) );
  AOI22_X1 U11803 ( .A1(n11187), .A2(n11190), .B1(n11186), .B2(n11185), .ZN(
        P2_U3472) );
  INV_X1 U11804 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U11805 ( .A1(n11191), .A2(n11190), .B1(n11189), .B2(n11188), .ZN(
        P2_U3429) );
  OAI21_X1 U11806 ( .B1(n11193), .B2(n11269), .A(n11192), .ZN(n11195) );
  AOI211_X1 U11807 ( .C1(n11197), .C2(n11196), .A(n11195), .B(n11194), .ZN(
        n11199) );
  AOI22_X1 U11808 ( .A1(n11276), .A2(n11199), .B1(n10383), .B2(n11275), .ZN(
        P1_U3536) );
  INV_X1 U11809 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U11810 ( .A1(n11280), .A2(n11199), .B1(n11198), .B2(n11277), .ZN(
        P1_U3495) );
  NAND2_X1 U11811 ( .A1(n11200), .A2(n11208), .ZN(n11201) );
  NAND2_X1 U11812 ( .A1(n11203), .A2(n7337), .ZN(n11204) );
  NAND3_X1 U11813 ( .A1(n11205), .A2(n11250), .A3(n11204), .ZN(n11216) );
  OAI21_X1 U11814 ( .B1(n7338), .B2(n11269), .A(n11216), .ZN(n11213) );
  NAND2_X1 U11815 ( .A1(n11207), .A2(n11206), .ZN(n11209) );
  XNOR2_X1 U11816 ( .A(n11209), .B(n11208), .ZN(n11211) );
  AOI222_X1 U11817 ( .A1(n11232), .A2(n11211), .B1(n11235), .B2(n11237), .C1(
        n11210), .C2(n11236), .ZN(n11222) );
  INV_X1 U11818 ( .A(n11222), .ZN(n11212) );
  AOI211_X1 U11819 ( .C1(n11219), .C2(n11273), .A(n11213), .B(n11212), .ZN(
        n11214) );
  AOI22_X1 U11820 ( .A1(n11276), .A2(n11214), .B1(n6592), .B2(n11275), .ZN(
        P1_U3537) );
  AOI22_X1 U11821 ( .A1(n11280), .A2(n11214), .B1(n6594), .B2(n11277), .ZN(
        P1_U3498) );
  AOI222_X1 U11822 ( .A1(n7337), .A2(n11245), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n11244), .C1(n11243), .C2(n11215), .ZN(n11221) );
  NOR2_X1 U11823 ( .A1(n11216), .A2(n11253), .ZN(n11217) );
  AOI21_X1 U11824 ( .B1(n11219), .B2(n11218), .A(n11217), .ZN(n11220) );
  OAI211_X1 U11825 ( .C1(n11258), .C2(n11222), .A(n11221), .B(n11220), .ZN(
        P1_U3278) );
  OAI21_X1 U11826 ( .B1(n11224), .B2(n11269), .A(n11223), .ZN(n11225) );
  AOI211_X1 U11827 ( .C1(n11227), .C2(n11273), .A(n11226), .B(n11225), .ZN(
        n11229) );
  AOI22_X1 U11828 ( .A1(n11276), .A2(n11229), .B1(n6582), .B2(n11275), .ZN(
        P1_U3538) );
  INV_X1 U11829 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U11830 ( .A1(n11280), .A2(n11229), .B1(n11228), .B2(n11277), .ZN(
        P1_U3501) );
  OAI211_X1 U11831 ( .C1(n11234), .C2(n11233), .A(n11232), .B(n11231), .ZN(
        n11240) );
  AOI22_X1 U11832 ( .A1(n11238), .A2(n11237), .B1(n11236), .B2(n11235), .ZN(
        n11239) );
  AND2_X1 U11833 ( .A1(n11240), .A2(n11239), .ZN(n11262) );
  INV_X1 U11834 ( .A(n11241), .ZN(n11242) );
  AOI222_X1 U11835 ( .A1(n11260), .A2(n11245), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n11244), .C1(n11243), .C2(n11242), .ZN(n11257) );
  NOR2_X1 U11836 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  NAND2_X1 U11837 ( .A1(n11260), .A2(n11249), .ZN(n11251) );
  NAND2_X1 U11838 ( .A1(n11251), .A2(n11250), .ZN(n11252) );
  OR2_X1 U11839 ( .A1(n5232), .A2(n11252), .ZN(n11261) );
  OAI22_X1 U11840 ( .A1(n11259), .A2(n11254), .B1(n11253), .B2(n11261), .ZN(
        n11255) );
  INV_X1 U11841 ( .A(n11255), .ZN(n11256) );
  OAI211_X1 U11842 ( .C1(n11258), .C2(n11262), .A(n11257), .B(n11256), .ZN(
        P1_U3276) );
  INV_X1 U11843 ( .A(n11259), .ZN(n11265) );
  INV_X1 U11844 ( .A(n11260), .ZN(n11263) );
  OAI211_X1 U11845 ( .C1(n11263), .C2(n11269), .A(n11262), .B(n11261), .ZN(
        n11264) );
  AOI21_X1 U11846 ( .B1(n11265), .B2(n11273), .A(n11264), .ZN(n11267) );
  AOI22_X1 U11847 ( .A1(n11276), .A2(n11267), .B1(n10422), .B2(n11275), .ZN(
        P1_U3539) );
  INV_X1 U11848 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U11849 ( .A1(n11280), .A2(n11267), .B1(n11266), .B2(n11277), .ZN(
        P1_U3504) );
  OAI21_X1 U11850 ( .B1(n11270), .B2(n11269), .A(n11268), .ZN(n11271) );
  AOI211_X1 U11851 ( .C1(n11274), .C2(n11273), .A(n11272), .B(n11271), .ZN(
        n11279) );
  AOI22_X1 U11852 ( .A1(n11276), .A2(n11279), .B1(n10427), .B2(n11275), .ZN(
        P1_U3540) );
  INV_X1 U11853 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U11854 ( .A1(n11280), .A2(n11279), .B1(n11278), .B2(n11277), .ZN(
        P1_U3507) );
  XNOR2_X1 U11855 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U5199 ( .A(n7200), .ZN(n7197) );
  CLKBUF_X2 U5194 ( .A(n7218), .Z(n7412) );
  CLKBUF_X1 U5210 ( .A(n6630), .Z(n6845) );
  CLKBUF_X1 U5214 ( .A(n7211), .Z(n5137) );
  CLKBUF_X1 U5229 ( .A(n10536), .Z(n5261) );
  CLKBUF_X1 U5634 ( .A(n6649), .Z(n6971) );
endmodule

