

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7202, n7203, n7204, n7205, n7206, n7207, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981;

  NAND2_X1 U7291 ( .A1(n12762), .A2(n12761), .ZN(n12765) );
  XNOR2_X1 U7292 ( .A(n12408), .B(n12409), .ZN(n12410) );
  INV_X1 U7293 ( .A(n10285), .ZN(n10286) );
  OAI21_X1 U7294 ( .B1(n8485), .B2(n8484), .A(n8209), .ZN(n8501) );
  CLKBUF_X2 U7295 ( .A(n9664), .Z(n10143) );
  INV_X1 U7296 ( .A(n11104), .ZN(n11109) );
  CLKBUF_X3 U7297 ( .A(n12691), .Z(n7192) );
  NAND4_X1 U7298 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n10042)
         );
  CLKBUF_X2 U7299 ( .A(n9103), .Z(n9411) );
  AND2_X1 U7300 ( .A1(n9387), .A2(n15536), .ZN(n11219) );
  INV_X2 U7301 ( .A(n8285), .ZN(n8477) );
  NAND2_X2 U7302 ( .A1(n7244), .A2(n8951), .ZN(n14374) );
  INV_X1 U7303 ( .A(n15527), .ZN(n8941) );
  NAND2_X1 U7304 ( .A1(n8301), .A2(n8293), .ZN(n10423) );
  BUF_X2 U7305 ( .A(n8953), .Z(n7206) );
  NAND2_X2 U7306 ( .A1(n8158), .A2(n8157), .ZN(n8216) );
  AND2_X1 U7307 ( .A1(n8228), .A2(n8225), .ZN(n8035) );
  NOR2_X1 U7308 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8228) );
  NOR2_X1 U7309 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8225) );
  AND2_X1 U7310 ( .A1(n9181), .A2(n8859), .ZN(n8860) );
  NOR2_X1 U7311 ( .A1(n8818), .A2(n7601), .ZN(n7598) );
  AND2_X1 U7312 ( .A1(n8035), .A2(n8033), .ZN(n7616) );
  INV_X1 U7313 ( .A(n8984), .ZN(n9268) );
  AND2_X1 U7314 ( .A1(n10805), .A2(n10397), .ZN(n9675) );
  OR2_X1 U7315 ( .A1(n8572), .A2(n8260), .ZN(n8262) );
  NOR2_X1 U7316 ( .A1(n8753), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8757) );
  AND2_X1 U7317 ( .A1(n8938), .A2(n10398), .ZN(n8953) );
  INV_X1 U7318 ( .A(n10360), .ZN(n8998) );
  INV_X1 U7319 ( .A(n10994), .ZN(n12708) );
  CLKBUF_X2 U7320 ( .A(n9268), .Z(n9419) );
  AOI21_X1 U7321 ( .B1(n12801), .B2(n12800), .A(n7365), .ZN(n12804) );
  INV_X1 U7322 ( .A(n10805), .ZN(n9908) );
  INV_X1 U7323 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U7324 ( .A1(n8040), .A2(n12542), .ZN(n8044) );
  BUF_X1 U7325 ( .A(n10709), .Z(n13521) );
  INV_X1 U7326 ( .A(n8513), .ZN(n8709) );
  OR2_X1 U7327 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  INV_X1 U7328 ( .A(n11709), .ZN(n11712) );
  OAI22_X1 U7329 ( .A1(n12883), .A2(n12884), .B1(n12771), .B2(n12906), .ZN(
        n12801) );
  AOI21_X1 U7330 ( .B1(n11477), .B2(n11476), .A(n11475), .ZN(n11480) );
  AND4_X1 U7331 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n12143)
         );
  AND2_X1 U7333 ( .A1(n8264), .A2(n7302), .ZN(n10709) );
  AOI211_X1 U7334 ( .C1(n15758), .C2(n14151), .A(n14150), .B(n14149), .ZN(
        n14210) );
  AND2_X2 U7335 ( .A1(n10972), .A2(n13780), .ZN(n15758) );
  OR2_X1 U7336 ( .A1(n8237), .A2(n7574), .ZN(n7573) );
  INV_X1 U7337 ( .A(n8216), .ZN(n10398) );
  INV_X1 U7338 ( .A(n10165), .ZN(n11525) );
  NAND2_X1 U7339 ( .A1(n8251), .A2(n8250), .ZN(n14226) );
  AND2_X1 U7340 ( .A1(n10347), .A2(n11219), .ZN(n12691) );
  XOR2_X1 U7341 ( .A(n14146), .B(n12728), .Z(n7190) );
  BUF_X1 U7342 ( .A(n10972), .Z(n7193) );
  XNOR2_X1 U7343 ( .A(n8759), .B(n8758), .ZN(n10972) );
  NAND2_X2 U7344 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  OR2_X2 U7345 ( .A1(n9911), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U7346 ( .A1(n10764), .A2(n10763), .ZN(n7191) );
  NAND2_X1 U7347 ( .A1(n10764), .A2(n10763), .ZN(n11039) );
  CLKBUF_X3 U7348 ( .A(n11039), .Z(n12802) );
  NOR2_X2 U7349 ( .A1(n14727), .A2(n7874), .ZN(n14712) );
  NOR2_X2 U7350 ( .A1(n14728), .A2(n14729), .ZN(n14727) );
  NAND3_X4 U7351 ( .A1(n8934), .A2(n8933), .A3(n8932), .ZN(n14375) );
  XNOR2_X2 U7352 ( .A(n9549), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9818) );
  NAND2_X2 U7353 ( .A1(n7690), .A2(n7689), .ZN(n9549) );
  NAND2_X4 U7354 ( .A1(n13405), .A2(n12201), .ZN(n9641) );
  NAND2_X2 U7355 ( .A1(n8874), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8875) );
  XNOR2_X2 U7356 ( .A(n13089), .B(n13088), .ZN(n13336) );
  OAI21_X2 U7358 ( .B1(n15194), .B2(n7193), .A(n13741), .ZN(n11104) );
  INV_X2 U7359 ( .A(n11109), .ZN(n12728) );
  INV_X1 U7360 ( .A(n11516), .ZN(n15596) );
  OAI211_X4 U7361 ( .C1(n7203), .C2(n10423), .A(n8957), .B(n8956), .ZN(n11516)
         );
  AND2_X4 U7362 ( .A1(n10329), .A2(n10398), .ZN(n13704) );
  AOI22_X2 U7363 ( .A1(n15912), .A2(n15911), .B1(n15944), .B2(n15932), .ZN(
        n14743) );
  NAND2_X2 U7364 ( .A1(n14758), .A2(n12436), .ZN(n15912) );
  INV_X1 U7365 ( .A(n9370), .ZN(n7194) );
  INV_X1 U7366 ( .A(n7194), .ZN(n7195) );
  NAND2_X1 U7367 ( .A1(n12333), .A2(n10224), .ZN(n13246) );
  INV_X1 U7368 ( .A(n12582), .ZN(n12526) );
  NAND2_X1 U7369 ( .A1(n11704), .A2(n11703), .ZN(n15709) );
  NAND2_X1 U7370 ( .A1(n10724), .A2(n10723), .ZN(n12510) );
  NOR2_X1 U7371 ( .A1(n14372), .A2(n11712), .ZN(n11699) );
  AND2_X1 U7372 ( .A1(n7415), .A2(n7308), .ZN(n10993) );
  AOI21_X1 U7373 ( .B1(n11127), .B2(n10715), .A(n11128), .ZN(n11123) );
  OR2_X1 U7374 ( .A1(n10355), .A2(n10913), .ZN(n7415) );
  INV_X4 U7375 ( .A(n12706), .ZN(n11435) );
  AND2_X1 U7376 ( .A1(n11007), .A2(n8297), .ZN(n13747) );
  INV_X2 U7377 ( .A(n12691), .ZN(n12640) );
  INV_X1 U7378 ( .A(n13814), .ZN(n12511) );
  INV_X1 U7379 ( .A(n11634), .ZN(n11198) );
  INV_X1 U7380 ( .A(n13815), .ZN(n11004) );
  INV_X1 U7381 ( .A(n15557), .ZN(n15553) );
  CLKBUF_X2 U7382 ( .A(n9655), .Z(n10011) );
  CLKBUF_X2 U7383 ( .A(n8947), .Z(n9407) );
  CLKBUF_X2 U7384 ( .A(n7206), .Z(n9249) );
  NOR2_X1 U7385 ( .A1(n11229), .A2(n15537), .ZN(n11220) );
  INV_X2 U7386 ( .A(n9015), .ZN(n8947) );
  INV_X1 U7387 ( .A(n8952), .ZN(n7202) );
  BUF_X1 U7388 ( .A(n8953), .Z(n7207) );
  NAND2_X1 U7389 ( .A1(n13779), .A2(n13736), .ZN(n13741) );
  NAND2_X1 U7390 ( .A1(n9496), .A2(n9495), .ZN(n10439) );
  BUF_X1 U7391 ( .A(n9597), .Z(n9598) );
  INV_X2 U7392 ( .A(n8772), .ZN(n13779) );
  CLKBUF_X2 U7393 ( .A(n8938), .Z(n10360) );
  NAND2_X1 U7394 ( .A1(n9485), .A2(n9490), .ZN(n10440) );
  OR2_X1 U7395 ( .A1(n9492), .A2(n9491), .ZN(n9496) );
  NAND2_X1 U7396 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  NAND2_X1 U7397 ( .A1(n8887), .A2(n8868), .ZN(n8870) );
  OAI21_X1 U7398 ( .B1(n8022), .B2(n8021), .A(n8020), .ZN(n9431) );
  MUX2_X1 U7399 ( .A(n13321), .B(n13260), .S(n15970), .Z(n13261) );
  MUX2_X1 U7400 ( .A(n13321), .B(n13320), .S(n15980), .Z(n13322) );
  AND2_X1 U7401 ( .A1(n13259), .A2(n13258), .ZN(n13321) );
  AND2_X1 U7402 ( .A1(n13067), .A2(n13066), .ZN(n13259) );
  AND2_X1 U7403 ( .A1(n13076), .A2(n13075), .ZN(n13327) );
  CLKBUF_X1 U7404 ( .A(n14573), .Z(n14797) );
  NAND2_X1 U7405 ( .A1(n14600), .A2(n14599), .ZN(n14598) );
  NAND2_X1 U7406 ( .A1(n8082), .A2(n8081), .ZN(n14330) );
  NAND2_X1 U7407 ( .A1(n12559), .A2(n12558), .ZN(n12723) );
  NAND2_X1 U7408 ( .A1(n14680), .A2(n12440), .ZN(n14655) );
  OR2_X1 U7409 ( .A1(n13099), .A2(n13136), .ZN(n13140) );
  NAND2_X1 U7410 ( .A1(n14323), .A2(n8086), .ZN(n14264) );
  AND2_X1 U7411 ( .A1(n7870), .A2(n7861), .ZN(n7860) );
  NAND2_X1 U7412 ( .A1(n14695), .A2(n7878), .ZN(n14680) );
  NAND2_X1 U7413 ( .A1(n7465), .A2(n7464), .ZN(n13455) );
  NAND2_X1 U7414 ( .A1(n14274), .A2(n7443), .ZN(n14323) );
  AOI21_X1 U7415 ( .B1(n12547), .B2(n7467), .A(n7466), .ZN(n7464) );
  NAND2_X1 U7416 ( .A1(n9962), .A2(n9961), .ZN(n13333) );
  AOI21_X1 U7417 ( .B1(n7889), .B2(n7893), .A(n7296), .ZN(n7888) );
  NAND2_X1 U7418 ( .A1(n9926), .A2(n8100), .ZN(n13167) );
  NAND2_X1 U7419 ( .A1(n9624), .A2(n9623), .ZN(n13339) );
  NAND3_X1 U7420 ( .A1(n8044), .A2(n8042), .A3(n8041), .ZN(n13488) );
  INV_X1 U7421 ( .A(n14574), .ZN(n14570) );
  OR2_X1 U7422 ( .A1(n12764), .A2(n7762), .ZN(n7755) );
  OR2_X1 U7423 ( .A1(n12763), .A2(n13173), .ZN(n7763) );
  NAND2_X1 U7424 ( .A1(n7585), .A2(n14204), .ZN(n13996) );
  INV_X1 U7425 ( .A(n14008), .ZN(n7585) );
  INV_X1 U7426 ( .A(n14021), .ZN(n7196) );
  XNOR2_X1 U7427 ( .A(n14010), .B(n13796), .ZN(n14006) );
  NAND2_X1 U7428 ( .A1(n12003), .A2(n8808), .ZN(n12054) );
  NAND2_X1 U7429 ( .A1(n7576), .A2(n7575), .ZN(n12191) );
  INV_X1 U7430 ( .A(n12059), .ZN(n7576) );
  OR2_X1 U7431 ( .A1(n10731), .A2(n10732), .ZN(n11023) );
  NAND2_X1 U7432 ( .A1(n8221), .A2(n8543), .ZN(n7954) );
  NAND2_X1 U7433 ( .A1(n8219), .A2(SI_18_), .ZN(n8222) );
  NAND2_X1 U7434 ( .A1(n8453), .A2(n8452), .ZN(n13603) );
  NAND2_X1 U7435 ( .A1(n9149), .A2(n9148), .ZN(n12408) );
  INV_X2 U7436 ( .A(n15818), .ZN(n7197) );
  NAND3_X1 U7437 ( .A1(n12510), .A2(n12513), .A3(n11106), .ZN(n12519) );
  INV_X2 U7438 ( .A(n15688), .ZN(n15690) );
  OR2_X2 U7439 ( .A1(n10332), .A2(P2_U3088), .ZN(n13812) );
  NAND2_X1 U7440 ( .A1(n10043), .A2(n10161), .ZN(n10163) );
  NAND2_X1 U7441 ( .A1(n9034), .A2(n9033), .ZN(n11763) );
  NAND2_X1 U7442 ( .A1(n9544), .A2(n9543), .ZN(n9795) );
  XNOR2_X1 U7443 ( .A(n10911), .B(n11634), .ZN(n10990) );
  AND2_X1 U7444 ( .A1(n10182), .A2(n10183), .ZN(n11679) );
  NAND2_X1 U7445 ( .A1(n8983), .A2(n7905), .ZN(n11709) );
  AND2_X1 U7446 ( .A1(n9949), .A2(n12868), .ZN(n9951) );
  OAI22_X1 U7447 ( .A1(n15529), .A2(n12640), .B1(n15565), .B2(n12708), .ZN(
        n10911) );
  NAND2_X1 U7448 ( .A1(n15553), .A2(n12924), .ZN(n10160) );
  INV_X1 U7449 ( .A(n11666), .ZN(n12920) );
  NOR2_X1 U7450 ( .A1(n10968), .A2(n10708), .ZN(n11174) );
  NAND4_X2 U7451 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n8994), .ZN(n14371)
         );
  NAND2_X1 U7452 ( .A1(n8305), .A2(n8304), .ZN(n13544) );
  NAND4_X1 U7453 ( .A1(n8327), .A2(n8326), .A3(n8325), .A4(n8324), .ZN(n13813)
         );
  NAND4_X1 U7454 ( .A1(n8913), .A2(n8912), .A3(n8911), .A4(n8910), .ZN(n14373)
         );
  NAND3_X1 U7455 ( .A1(n8928), .A2(n8927), .A3(n8144), .ZN(n11503) );
  AND4_X1 U7456 ( .A1(n9716), .A2(n9715), .A3(n9714), .A4(n9713), .ZN(n11666)
         );
  INV_X2 U7457 ( .A(n9759), .ZN(n10012) );
  AND4_X1 U7458 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n11545)
         );
  NAND2_X1 U7459 ( .A1(n7202), .A2(n8270), .ZN(n8927) );
  INV_X4 U7460 ( .A(n10708), .ZN(n14076) );
  AND2_X1 U7461 ( .A1(n7303), .A2(n8280), .ZN(n10973) );
  NAND4_X1 U7462 ( .A1(n8289), .A2(n8288), .A3(n8287), .A4(n8286), .ZN(n13815)
         );
  CLKBUF_X3 U7463 ( .A(n8998), .Z(n7200) );
  OAI211_X1 U7464 ( .C1(n10892), .C2(n10805), .A(n7640), .B(n7639), .ZN(n15580) );
  CLKBUF_X3 U7465 ( .A(n8929), .Z(n9410) );
  AND3_X1 U7466 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(n11045) );
  INV_X2 U7467 ( .A(n9946), .ZN(n10130) );
  OAI21_X1 U7468 ( .B1(n8312), .B2(n7521), .A(n7519), .ZN(n8332) );
  INV_X1 U7469 ( .A(n11219), .ZN(n10909) );
  CLKBUF_X2 U7470 ( .A(n8952), .Z(n7203) );
  NOR2_X1 U7471 ( .A1(n9850), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9866) );
  AND2_X2 U7472 ( .A1(n9598), .A2(n12201), .ZN(n9667) );
  OR2_X1 U7473 ( .A1(n9720), .A2(n9532), .ZN(n9534) );
  MUX2_X1 U7474 ( .A(n8755), .B(n8754), .S(n8783), .Z(n13736) );
  INV_X1 U7475 ( .A(n8877), .ZN(n14881) );
  NAND2_X2 U7476 ( .A1(n8253), .A2(n8252), .ZN(n8285) );
  NAND2_X1 U7477 ( .A1(n9390), .A2(n8898), .ZN(n11229) );
  NAND2_X1 U7478 ( .A1(n9595), .A2(n9594), .ZN(n12201) );
  NAND2_X1 U7479 ( .A1(n8873), .A2(n8874), .ZN(n8877) );
  OAI21_X1 U7480 ( .B1(n9906), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9907) );
  MUX2_X1 U7481 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9593), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9594) );
  INV_X1 U7482 ( .A(n14226), .ZN(n8252) );
  XNOR2_X1 U7483 ( .A(n9596), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U7484 ( .A1(n9583), .A2(n9592), .ZN(n12134) );
  MUX2_X1 U7485 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8869), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8873) );
  CLKBUF_X1 U7486 ( .A(n13036), .Z(n7384) );
  AND2_X1 U7487 ( .A1(n8753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U7488 ( .A1(n9595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U7489 ( .A1(n8249), .A2(n8248), .ZN(n8251) );
  OAI21_X1 U7490 ( .B1(n8173), .B2(n7521), .A(n8329), .ZN(n7520) );
  OR2_X1 U7491 ( .A1(n10030), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U7492 ( .A1(n7567), .A2(n7566), .ZN(n14886) );
  XNOR2_X1 U7493 ( .A(n8907), .B(n8893), .ZN(n15536) );
  MUX2_X1 U7494 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9581), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n9583) );
  AND2_X1 U7495 ( .A1(n8902), .A2(n8906), .ZN(n15537) );
  AND2_X1 U7496 ( .A1(n9862), .A2(n9861), .ZN(n9878) );
  NOR2_X1 U7497 ( .A1(n7572), .A2(n7571), .ZN(n7570) );
  NOR2_X1 U7498 ( .A1(n7231), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U7499 ( .A1(n8244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8236) );
  NAND2_X2 U7500 ( .A1(n10397), .A2(P1_U3086), .ZN(n14893) );
  NAND2_X2 U7501 ( .A1(n10398), .A2(P2_U3088), .ZN(n14239) );
  INV_X4 U7502 ( .A(n10398), .ZN(n10397) );
  AND2_X1 U7503 ( .A1(n8861), .A2(n7992), .ZN(n7991) );
  AND2_X2 U7504 ( .A1(n8980), .A2(n8981), .ZN(n8861) );
  AND2_X1 U7505 ( .A1(n8120), .A2(n9706), .ZN(n8119) );
  AND2_X1 U7506 ( .A1(n7993), .A2(n8088), .ZN(n7992) );
  AND4_X1 U7507 ( .A1(n9572), .A2(n9571), .A3(n9729), .A4(n9783), .ZN(n9573)
         );
  INV_X1 U7508 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9478) );
  NOR2_X1 U7509 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9479) );
  INV_X1 U7510 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9030) );
  INV_X1 U7511 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9059) );
  INV_X1 U7512 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7990) );
  INV_X1 U7513 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9127) );
  INV_X1 U7514 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8154) );
  INV_X1 U7515 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8152) );
  INV_X1 U7516 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8155) );
  INV_X1 U7517 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8153) );
  INV_X1 U7518 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9108) );
  INV_X1 U7519 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9094) );
  NOR2_X1 U7520 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8863) );
  NOR2_X1 U7521 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8120) );
  INV_X1 U7522 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9729) );
  INV_X1 U7523 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U7524 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9571) );
  NOR2_X1 U7525 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9572) );
  INV_X1 U7526 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9833) );
  NOR2_X1 U7527 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7740) );
  NOR2_X1 U7528 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7741) );
  INV_X1 U7529 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n10022) );
  INV_X1 U7530 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8783) );
  INV_X1 U7531 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8776) );
  NOR2_X1 U7532 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7571) );
  INV_X4 U7533 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7534 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8763) );
  NOR2_X1 U7535 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7568) );
  NOR2_X1 U7536 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7569) );
  NOR2_X4 U7537 ( .A1(n9811), .A2(n8142), .ZN(n10069) );
  AND2_X1 U7538 ( .A1(n10972), .A2(n8772), .ZN(n10986) );
  AND2_X1 U7539 ( .A1(n10329), .A2(n10397), .ZN(n7198) );
  AND2_X1 U7540 ( .A1(n10329), .A2(n10397), .ZN(n8420) );
  NOR2_X2 U7541 ( .A1(n14841), .A2(n14715), .ZN(n14704) );
  NAND2_X2 U7543 ( .A1(n13120), .A2(n10262), .ZN(n13110) );
  NAND2_X2 U7544 ( .A1(n7646), .A2(n7315), .ZN(n13120) );
  CLKBUF_X1 U7545 ( .A(n8998), .Z(n7199) );
  NAND4_X1 U7547 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n8961)
         );
  OR2_X1 U7548 ( .A1(n9015), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U7549 ( .A1(n8938), .A2(n10397), .ZN(n8952) );
  NAND2_X2 U7550 ( .A1(n13246), .A2(n13245), .ZN(n13244) );
  AND2_X2 U7551 ( .A1(n14881), .A2(n8882), .ZN(n9103) );
  NAND2_X1 U7552 ( .A1(n8158), .A2(n8157), .ZN(n7204) );
  INV_X1 U7553 ( .A(n12802), .ZN(n7205) );
  AND4_X4 U7554 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(n9652)
         );
  OR2_X1 U7555 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  AOI211_X2 U7556 ( .C1(n14579), .C2(n14578), .A(n14763), .B(n14577), .ZN(
        n14787) );
  OAI21_X2 U7557 ( .B1(n13202), .B2(n10292), .A(n10243), .ZN(n13183) );
  XNOR2_X1 U7558 ( .A(n14371), .B(n11716), .ZN(n15658) );
  NOR2_X4 U7559 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9660) );
  XNOR2_X1 U7561 ( .A(n9907), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13025) );
  NOR2_X4 U7562 ( .A1(n15888), .A2(n14764), .ZN(n15918) );
  OR2_X2 U7563 ( .A1(n12435), .A2(n12421), .ZN(n14764) );
  INV_X1 U7564 ( .A(n9536), .ZN(n7718) );
  NAND2_X1 U7565 ( .A1(n7864), .A2(n7862), .ZN(n7861) );
  INV_X1 U7566 ( .A(n7866), .ZN(n7862) );
  AOI21_X1 U7567 ( .B1(n8112), .B2(n9774), .A(n8111), .ZN(n8110) );
  OR2_X1 U7568 ( .A1(n12738), .A2(n12913), .ZN(n10217) );
  XNOR2_X1 U7569 ( .A(n7501), .B(P3_IR_REG_27__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U7570 ( .A1(n7502), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U7571 ( .A1(n13488), .A2(n12544), .ZN(n12546) );
  NAND2_X1 U7572 ( .A1(n13447), .A2(n7239), .ZN(n12543) );
  INV_X1 U7573 ( .A(n8598), .ZN(n8599) );
  NAND2_X1 U7574 ( .A1(n7955), .A2(n7330), .ZN(n8586) );
  INV_X1 U7575 ( .A(n8565), .ZN(n7952) );
  INV_X1 U7576 ( .A(n9682), .ZN(n9759) );
  AND2_X1 U7577 ( .A1(n9997), .A2(n12806), .ZN(n13055) );
  NAND2_X1 U7578 ( .A1(n8959), .A2(n8958), .ZN(n8967) );
  NAND2_X1 U7579 ( .A1(n8984), .A2(n14374), .ZN(n8959) );
  INV_X1 U7580 ( .A(n13668), .ZN(n7872) );
  INV_X1 U7581 ( .A(n13669), .ZN(n7869) );
  NAND2_X1 U7582 ( .A1(n10270), .A2(n10285), .ZN(n7719) );
  NOR2_X1 U7583 ( .A1(n7369), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U7584 ( .A1(n7899), .A2(n7261), .ZN(n7897) );
  OR2_X1 U7585 ( .A1(n13276), .A2(n13138), .ZN(n10262) );
  AND2_X1 U7586 ( .A1(n7314), .A2(n9955), .ZN(n8124) );
  NAND2_X1 U7587 ( .A1(n8098), .A2(n9666), .ZN(n11533) );
  AND2_X1 U7588 ( .A1(n8099), .A2(n9665), .ZN(n8098) );
  INV_X1 U7589 ( .A(n7700), .ZN(n7698) );
  AOI21_X1 U7590 ( .B1(n7692), .B2(n7694), .A(n7337), .ZN(n7689) );
  NAND2_X1 U7591 ( .A1(n9795), .A2(n7692), .ZN(n7690) );
  NOR2_X1 U7592 ( .A1(n7718), .A2(n7714), .ZN(n7713) );
  INV_X1 U7593 ( .A(n9533), .ZN(n7714) );
  NAND2_X1 U7594 ( .A1(n13670), .A2(n7860), .ZN(n7859) );
  INV_X1 U7595 ( .A(n8254), .ZN(n8253) );
  OR2_X1 U7596 ( .A1(n14104), .A2(n13690), .ZN(n8828) );
  NOR2_X1 U7597 ( .A1(n13920), .A2(n7812), .ZN(n7811) );
  INV_X1 U7598 ( .A(n7813), .ZN(n7812) );
  NOR2_X1 U7599 ( .A1(n14006), .A2(n7801), .ZN(n7800) );
  INV_X1 U7600 ( .A(n7803), .ZN(n7801) );
  INV_X1 U7601 ( .A(n7602), .ZN(n7601) );
  NAND2_X1 U7602 ( .A1(n8802), .A2(n8801), .ZN(n7624) );
  INV_X1 U7603 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8234) );
  NAND4_X1 U7604 ( .A1(n8036), .A2(n8141), .A3(n8233), .A4(n8232), .ZN(n7617)
         );
  NOR2_X1 U7605 ( .A1(n8417), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8435) );
  XNOR2_X1 U7606 ( .A(n9460), .B(n14562), .ZN(n9503) );
  OR2_X1 U7607 ( .A1(n14692), .A2(n14662), .ZN(n12440) );
  INV_X1 U7608 ( .A(n15911), .ZN(n7971) );
  INV_X1 U7609 ( .A(n8905), .ZN(n9387) );
  OR2_X1 U7610 ( .A1(n12079), .A2(n7986), .ZN(n7985) );
  INV_X1 U7611 ( .A(n7988), .ZN(n7986) );
  NAND2_X1 U7612 ( .A1(n7923), .A2(n7922), .ZN(n8669) );
  AOI21_X1 U7613 ( .B1(n7925), .B2(n7927), .A(n7347), .ZN(n7922) );
  OAI21_X1 U7614 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8600) );
  XNOR2_X1 U7615 ( .A(n8564), .B(SI_19_), .ZN(n8565) );
  INV_X1 U7616 ( .A(n8220), .ZN(n8219) );
  INV_X1 U7617 ( .A(n7938), .ZN(n7937) );
  OAI21_X1 U7618 ( .B1(n8366), .B2(n7939), .A(n8188), .ZN(n7938) );
  OAI21_X1 U7619 ( .B1(n8290), .B2(n8170), .A(n8169), .ZN(n8302) );
  NOR2_X1 U7620 ( .A1(n15265), .A2(n15264), .ZN(n15270) );
  NOR2_X1 U7621 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15263), .ZN(n15264) );
  AOI21_X1 U7622 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15292), .A(n15291), .ZN(
        n15299) );
  AND2_X1 U7623 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  NOR2_X1 U7624 ( .A1(n7252), .A2(n7221), .ZN(n7764) );
  INV_X1 U7625 ( .A(n12768), .ZN(n7760) );
  XNOR2_X1 U7626 ( .A(n10816), .B(n10858), .ZN(n10850) );
  NOR2_X1 U7627 ( .A1(n15400), .A2(n7516), .ZN(n7515) );
  INV_X1 U7628 ( .A(n15383), .ZN(n7516) );
  INV_X1 U7629 ( .A(n7513), .ZN(n7512) );
  OAI21_X1 U7630 ( .B1(n15400), .B2(n7514), .A(n7335), .ZN(n7513) );
  NAND2_X1 U7631 ( .A1(n15381), .A2(n15383), .ZN(n7514) );
  NOR2_X1 U7632 ( .A1(n9980), .A2(n9979), .ZN(n9997) );
  NAND2_X1 U7633 ( .A1(n7236), .A2(n13223), .ZN(n13222) );
  OAI21_X1 U7634 ( .B1(n9817), .B2(n8117), .A(n8114), .ZN(n8113) );
  NOR2_X1 U7635 ( .A1(n12738), .A2(n12780), .ZN(n8117) );
  AOI21_X1 U7636 ( .B1(n8118), .B2(n12780), .A(n8115), .ZN(n8114) );
  AOI21_X1 U7637 ( .B1(n8110), .B2(n8107), .A(n7293), .ZN(n8106) );
  INV_X1 U7638 ( .A(n8112), .ZN(n8107) );
  OR2_X1 U7639 ( .A1(n11526), .A2(n15797), .ZN(n10783) );
  INV_X1 U7640 ( .A(n13036), .ZN(n10032) );
  OR2_X1 U7641 ( .A1(n13339), .A2(n13128), .ZN(n10058) );
  NAND2_X1 U7642 ( .A1(n13149), .A2(n10260), .ZN(n7647) );
  INV_X1 U7643 ( .A(n9675), .ZN(n9946) );
  NAND2_X1 U7644 ( .A1(n13167), .A2(n9941), .ZN(n13156) );
  NAND2_X1 U7645 ( .A1(n7656), .A2(n7659), .ZN(n12166) );
  AND2_X1 U7646 ( .A1(n12350), .A2(n7660), .ZN(n7659) );
  NAND2_X1 U7647 ( .A1(n7661), .A2(n10213), .ZN(n7660) );
  NAND2_X1 U7648 ( .A1(n10078), .A2(n10077), .ZN(n10108) );
  AND2_X1 U7649 ( .A1(n10095), .A2(n10076), .ZN(n7747) );
  NAND2_X1 U7650 ( .A1(n7725), .A2(n7723), .ZN(n9990) );
  AOI21_X1 U7651 ( .B1(n7726), .B2(n7728), .A(n7724), .ZN(n7723) );
  INV_X1 U7652 ( .A(n9974), .ZN(n7724) );
  INV_X1 U7653 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9539) );
  XNOR2_X1 U7654 ( .A(n14183), .B(n12730), .ZN(n12731) );
  NOR2_X1 U7655 ( .A1(n12542), .A2(n8047), .ZN(n8045) );
  AND2_X1 U7656 ( .A1(n7584), .A2(n13688), .ZN(n7583) );
  OR2_X1 U7657 ( .A1(n7807), .A2(n13930), .ZN(n7806) );
  NAND2_X1 U7658 ( .A1(n13910), .A2(n8825), .ZN(n13901) );
  OR2_X1 U7659 ( .A1(n13944), .A2(n13792), .ZN(n7813) );
  AND2_X1 U7660 ( .A1(n13962), .A2(n14191), .ZN(n13940) );
  INV_X1 U7661 ( .A(n13933), .ZN(n13930) );
  AOI21_X1 U7662 ( .B1(n7525), .B2(n7528), .A(n7281), .ZN(n7523) );
  AND2_X1 U7663 ( .A1(n13932), .A2(n8666), .ZN(n13966) );
  OAI21_X1 U7664 ( .B1(n8542), .B2(n7792), .A(n7790), .ZN(n14042) );
  INV_X1 U7665 ( .A(n7791), .ZN(n7790) );
  OAI21_X1 U7666 ( .B1(n7241), .B2(n7792), .A(n14044), .ZN(n7791) );
  INV_X1 U7667 ( .A(n8562), .ZN(n7792) );
  NAND2_X1 U7668 ( .A1(n7816), .A2(n7815), .ZN(n12370) );
  AOI21_X1 U7669 ( .B1(n7817), .B2(n12186), .A(n7248), .ZN(n7815) );
  AOI21_X1 U7670 ( .B1(n7787), .B2(n7789), .A(n7271), .ZN(n7785) );
  OAI21_X1 U7671 ( .B1(n8797), .B2(n7608), .A(n7607), .ZN(n11462) );
  INV_X1 U7672 ( .A(n7609), .ZN(n7608) );
  AND2_X1 U7673 ( .A1(n7604), .A2(n13756), .ZN(n7607) );
  NAND2_X1 U7674 ( .A1(n7605), .A2(n7609), .ZN(n7604) );
  INV_X1 U7675 ( .A(n14074), .ZN(n14063) );
  NAND2_X1 U7676 ( .A1(n8550), .A2(n8549), .ZN(n14155) );
  INV_X1 U7677 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8895) );
  OAI21_X1 U7678 ( .B1(n11205), .B2(n7420), .A(n7424), .ZN(n11597) );
  NAND2_X1 U7679 ( .A1(n7427), .A2(n11433), .ZN(n7424) );
  NAND2_X1 U7680 ( .A1(n7425), .A2(n7427), .ZN(n7420) );
  NAND2_X1 U7682 ( .A1(n8876), .A2(n8877), .ZN(n8919) );
  NAND2_X1 U7683 ( .A1(n8892), .A2(n8891), .ZN(n14604) );
  NAND2_X1 U7684 ( .A1(n14633), .A2(n14618), .ZN(n14612) );
  XNOR2_X1 U7685 ( .A(n14817), .B(n14358), .ZN(n14630) );
  NOR2_X1 U7686 ( .A1(n7563), .A2(n14848), .ZN(n7562) );
  INV_X1 U7687 ( .A(n7564), .ZN(n7563) );
  AND2_X1 U7688 ( .A1(n9433), .A2(n12436), .ZN(n14761) );
  AOI21_X1 U7689 ( .B1(n7215), .B2(n7903), .A(n7900), .ZN(n7899) );
  NOR2_X1 U7690 ( .A1(n12408), .A2(n12409), .ZN(n7900) );
  NAND2_X1 U7691 ( .A1(n7873), .A2(n7277), .ZN(n9488) );
  INV_X1 U7692 ( .A(n8899), .ZN(n7873) );
  NAND2_X1 U7693 ( .A1(n15259), .A2(n15258), .ZN(n7406) );
  AND2_X1 U7694 ( .A1(n12799), .A2(n13091), .ZN(n7365) );
  AOI21_X1 U7695 ( .B1(n13070), .B2(n10011), .A(n10001), .ZN(n13077) );
  OR2_X1 U7696 ( .A1(n13895), .A2(n13894), .ZN(n14101) );
  INV_X1 U7697 ( .A(n14183), .ZN(n14104) );
  XNOR2_X1 U7698 ( .A(n15257), .B(n7917), .ZN(n15259) );
  INV_X1 U7699 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7917) );
  INV_X1 U7700 ( .A(n8967), .ZN(n8960) );
  AOI21_X1 U7701 ( .B1(n7840), .B2(n7838), .A(n7837), .ZN(n7836) );
  OR2_X1 U7702 ( .A1(n9115), .A2(n9116), .ZN(n9117) );
  AOI21_X1 U7703 ( .B1(n9100), .B2(n8004), .A(n8002), .ZN(n8001) );
  NAND2_X1 U7704 ( .A1(n13601), .A2(n7823), .ZN(n7822) );
  NOR2_X1 U7705 ( .A1(n7845), .A2(n13613), .ZN(n7846) );
  INV_X1 U7706 ( .A(n13619), .ZN(n7843) );
  NAND2_X1 U7707 ( .A1(n13613), .A2(n7845), .ZN(n7844) );
  NAND2_X1 U7708 ( .A1(n13623), .A2(n13625), .ZN(n7829) );
  NAND2_X1 U7709 ( .A1(n7376), .A2(n7375), .ZN(n9254) );
  NAND2_X1 U7710 ( .A1(n9241), .A2(n9243), .ZN(n7375) );
  INV_X1 U7711 ( .A(n9269), .ZN(n8018) );
  NOR2_X1 U7712 ( .A1(n13650), .A2(n13647), .ZN(n7834) );
  NAND2_X1 U7713 ( .A1(n13650), .A2(n13647), .ZN(n7833) );
  NOR2_X1 U7714 ( .A1(n7872), .A2(n7869), .ZN(n7868) );
  NOR2_X1 U7715 ( .A1(n8012), .A2(n8011), .ZN(n8010) );
  INV_X1 U7716 ( .A(n9304), .ZN(n8011) );
  NOR2_X1 U7717 ( .A1(n9293), .A2(n8013), .ZN(n8012) );
  NOR2_X1 U7718 ( .A1(n8009), .A2(n9305), .ZN(n8008) );
  AND2_X1 U7719 ( .A1(n10309), .A2(n10307), .ZN(n7721) );
  NOR2_X1 U7720 ( .A1(n7850), .A2(n13656), .ZN(n7851) );
  NAND2_X1 U7721 ( .A1(n7850), .A2(n13656), .ZN(n7849) );
  AND2_X1 U7722 ( .A1(n7871), .A2(n7867), .ZN(n7866) );
  NAND2_X1 U7723 ( .A1(n7872), .A2(n7869), .ZN(n7867) );
  AND2_X1 U7724 ( .A1(n13678), .A2(n13666), .ZN(n7871) );
  AND2_X1 U7725 ( .A1(n8776), .A2(n8783), .ZN(n8141) );
  INV_X1 U7726 ( .A(n7926), .ZN(n7925) );
  OAI21_X1 U7727 ( .B1(n7928), .B2(n7927), .A(n8651), .ZN(n7926) );
  AOI21_X1 U7728 ( .B1(n8432), .B2(n8200), .A(n7934), .ZN(n7933) );
  INV_X1 U7729 ( .A(n8446), .ZN(n7934) );
  NOR2_X1 U7730 ( .A1(n15225), .A2(n7921), .ZN(n15231) );
  AND2_X1 U7731 ( .A1(n15226), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7921) );
  INV_X1 U7732 ( .A(n12740), .ZN(n7773) );
  INV_X1 U7733 ( .A(n12351), .ZN(n7770) );
  INV_X1 U7734 ( .A(n12201), .ZN(n9599) );
  NAND2_X1 U7735 ( .A1(n11057), .A2(n11058), .ZN(n11154) );
  NAND2_X1 U7736 ( .A1(n15476), .A2(n12961), .ZN(n12962) );
  NAND2_X1 U7737 ( .A1(n7508), .A2(n15504), .ZN(n7503) );
  INV_X1 U7738 ( .A(n13005), .ZN(n7508) );
  OR2_X1 U7739 ( .A1(n13378), .A2(n12910), .ZN(n10238) );
  NAND2_X1 U7740 ( .A1(n12917), .A2(n11876), .ZN(n8112) );
  NAND2_X1 U7741 ( .A1(n10176), .A2(n10173), .ZN(n8099) );
  INV_X1 U7742 ( .A(n10248), .ZN(n7671) );
  OR2_X1 U7743 ( .A1(n13369), .A2(n13213), .ZN(n10243) );
  AND2_X1 U7744 ( .A1(n13369), .A2(n13213), .ZN(n10292) );
  NAND2_X1 U7745 ( .A1(n11816), .A2(n10074), .ZN(n7748) );
  AND2_X1 U7746 ( .A1(n9578), .A2(n9579), .ZN(n8130) );
  INV_X1 U7747 ( .A(n10020), .ZN(n7739) );
  OAI21_X1 U7748 ( .B1(n9732), .B2(n7718), .A(n9748), .ZN(n7717) );
  AND2_X1 U7749 ( .A1(n10430), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9532) );
  INV_X1 U7750 ( .A(n7239), .ZN(n8047) );
  NOR2_X1 U7751 ( .A1(n12343), .A2(n7462), .ZN(n7461) );
  INV_X1 U7752 ( .A(n8039), .ZN(n7462) );
  AND2_X1 U7753 ( .A1(n7858), .A2(n7313), .ZN(n7857) );
  NAND2_X1 U7754 ( .A1(n7860), .A2(n7863), .ZN(n7858) );
  INV_X1 U7755 ( .A(n14084), .ZN(n7793) );
  INV_X1 U7756 ( .A(n8814), .ZN(n7597) );
  NOR2_X1 U7757 ( .A1(n13767), .A2(n7596), .ZN(n7595) );
  NOR2_X1 U7758 ( .A1(n12186), .A2(n7597), .ZN(n7596) );
  OR2_X1 U7759 ( .A1(n7612), .A2(n7611), .ZN(n7605) );
  INV_X1 U7760 ( .A(n8796), .ZN(n7611) );
  INV_X1 U7761 ( .A(n8798), .ZN(n7612) );
  INV_X1 U7762 ( .A(n8791), .ZN(n7590) );
  NAND2_X1 U7763 ( .A1(n8790), .A2(n8789), .ZN(n11337) );
  OR2_X1 U7764 ( .A1(n8572), .A2(n8276), .ZN(n8278) );
  INV_X1 U7765 ( .A(n14187), .ZN(n13923) );
  AND3_X1 U7766 ( .A1(n8224), .A2(n8227), .A3(n8229), .ZN(n8032) );
  AND2_X1 U7767 ( .A1(n8757), .A2(n8758), .ZN(n8761) );
  NOR2_X1 U7768 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8224) );
  NOR2_X1 U7769 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8226) );
  OAI21_X1 U7770 ( .B1(n12596), .B2(n7419), .A(n7416), .ZN(n12614) );
  INV_X1 U7771 ( .A(n8068), .ZN(n7419) );
  AOI21_X1 U7772 ( .B1(n8068), .B2(n7418), .A(n7417), .ZN(n7416) );
  INV_X1 U7773 ( .A(n12609), .ZN(n7417) );
  NAND2_X1 U7774 ( .A1(n7212), .A2(n7275), .ZN(n14675) );
  NOR2_X1 U7775 ( .A1(n14761), .A2(n12450), .ZN(n7968) );
  INV_X1 U7776 ( .A(n12410), .ZN(n7903) );
  NAND2_X1 U7777 ( .A1(n15565), .A2(n8961), .ZN(n11232) );
  NAND2_X1 U7778 ( .A1(n12103), .A2(n7989), .ZN(n7988) );
  NOR2_X1 U7779 ( .A1(n12095), .A2(n12100), .ZN(n7987) );
  AND2_X1 U7780 ( .A1(n8905), .A2(n11229), .ZN(n15526) );
  INV_X1 U7781 ( .A(n7947), .ZN(n7946) );
  AOI21_X1 U7782 ( .B1(n7947), .B2(n7945), .A(n7944), .ZN(n7943) );
  INV_X1 U7783 ( .A(n9363), .ZN(n7944) );
  INV_X1 U7784 ( .A(n9358), .ZN(n7945) );
  NOR2_X1 U7785 ( .A1(n9374), .A2(n7948), .ZN(n7947) );
  INV_X1 U7786 ( .A(n9361), .ZN(n7948) );
  OAI21_X1 U7787 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n9359) );
  NAND2_X1 U7788 ( .A1(n8894), .A2(n8095), .ZN(n8097) );
  NOR2_X1 U7789 ( .A1(n9480), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U7790 ( .A1(n7438), .A2(n7440), .ZN(n8896) );
  INV_X1 U7791 ( .A(n7441), .ZN(n7440) );
  OAI21_X1 U7792 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7441) );
  INV_X1 U7793 ( .A(n8515), .ZN(n7940) );
  NAND2_X1 U7794 ( .A1(n8416), .A2(n8197), .ZN(n8433) );
  INV_X1 U7795 ( .A(n8186), .ZN(n7939) );
  INV_X1 U7796 ( .A(n8189), .ZN(n7936) );
  INV_X1 U7797 ( .A(n7520), .ZN(n7519) );
  INV_X1 U7798 ( .A(n8174), .ZN(n7521) );
  NAND2_X1 U7799 ( .A1(n8312), .A2(n8173), .ZN(n8315) );
  INV_X1 U7800 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8156) );
  XNOR2_X1 U7801 ( .A(n14384), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n15220) );
  XNOR2_X1 U7802 ( .A(n15231), .B(n7920), .ZN(n15232) );
  AOI21_X1 U7803 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(n15240), .A(n15239), .ZN(
        n15252) );
  INV_X1 U7804 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U7805 ( .A1(n15299), .A2(n15298), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n15297), .ZN(n15304) );
  INV_X1 U7806 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12829) );
  INV_X1 U7807 ( .A(n11040), .ZN(n7752) );
  NAND2_X1 U7808 ( .A1(n11883), .A2(n11882), .ZN(n11981) );
  AOI21_X1 U7809 ( .B1(n7744), .B2(n7746), .A(n7329), .ZN(n7742) );
  INV_X1 U7810 ( .A(n11982), .ZN(n7768) );
  OAI21_X1 U7811 ( .B1(n13076), .B2(n7675), .A(n7673), .ZN(n10149) );
  AOI21_X1 U7812 ( .B1(n7676), .B2(n7674), .A(n7298), .ZN(n7673) );
  INV_X1 U7813 ( .A(n7676), .ZN(n7675) );
  AND4_X1 U7814 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n12838)
         );
  XNOR2_X1 U7815 ( .A(n11154), .B(n9736), .ZN(n11059) );
  NAND2_X1 U7816 ( .A1(n11059), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11156) );
  OR2_X1 U7817 ( .A1(n7512), .A2(n15427), .ZN(n7511) );
  NAND2_X1 U7818 ( .A1(n15451), .A2(n12935), .ZN(n15470) );
  AOI21_X1 U7819 ( .B1(n15470), .B2(n15466), .A(n7491), .ZN(n12937) );
  AND2_X1 U7820 ( .A1(n12970), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7491) );
  OR2_X1 U7821 ( .A1(n15519), .A2(n15518), .ZN(n7493) );
  NOR2_X1 U7822 ( .A1(n12969), .A2(n7505), .ZN(n7504) );
  INV_X1 U7823 ( .A(n15505), .ZN(n7505) );
  OAI21_X1 U7824 ( .B1(n9986), .B2(n8127), .A(n8126), .ZN(n10019) );
  AOI21_X1 U7825 ( .B1(n8128), .B2(n13080), .A(n7225), .ZN(n8126) );
  INV_X1 U7826 ( .A(n8128), .ZN(n8127) );
  NOR2_X1 U7827 ( .A1(n10059), .A2(n7685), .ZN(n7684) );
  INV_X1 U7828 ( .A(n10158), .ZN(n7685) );
  NAND2_X1 U7829 ( .A1(n13068), .A2(n10273), .ZN(n7683) );
  AND2_X1 U7830 ( .A1(n13078), .A2(n9987), .ZN(n13063) );
  NAND2_X1 U7831 ( .A1(n9956), .A2(n9955), .ZN(n13099) );
  INV_X1 U7832 ( .A(n13186), .ZN(n13213) );
  AOI21_X1 U7833 ( .B1(n13229), .B2(n7645), .A(n7644), .ZN(n7643) );
  INV_X1 U7834 ( .A(n10228), .ZN(n7645) );
  INV_X1 U7835 ( .A(n10238), .ZN(n7644) );
  INV_X1 U7836 ( .A(n12910), .ZN(n13242) );
  NAND2_X1 U7837 ( .A1(n12328), .A2(n7274), .ZN(n13236) );
  INV_X1 U7838 ( .A(n13245), .ZN(n9872) );
  AND2_X1 U7839 ( .A1(n10230), .A2(n10228), .ZN(n13245) );
  NAND2_X1 U7840 ( .A1(n12330), .A2(n12329), .ZN(n12328) );
  NAND2_X1 U7841 ( .A1(n8104), .A2(n8102), .ZN(n12155) );
  AOI21_X1 U7842 ( .B1(n7217), .B2(n8108), .A(n8103), .ZN(n8102) );
  INV_X1 U7843 ( .A(n12137), .ZN(n8103) );
  AND2_X1 U7844 ( .A1(n10213), .A2(n10212), .ZN(n12175) );
  NAND2_X1 U7845 ( .A1(n11996), .A2(n10208), .ZN(n12159) );
  INV_X1 U7846 ( .A(n8110), .ZN(n8108) );
  NOR2_X1 U7847 ( .A1(n11897), .A2(n7664), .ZN(n7663) );
  AOI21_X1 U7848 ( .B1(n7652), .B2(n7655), .A(n10153), .ZN(n7650) );
  INV_X1 U7849 ( .A(n10058), .ZN(n7655) );
  NAND2_X1 U7850 ( .A1(n8123), .A2(n8122), .ZN(n13090) );
  NOR2_X1 U7851 ( .A1(n8151), .A2(n7264), .ZN(n8122) );
  AND3_X1 U7852 ( .A1(n9602), .A2(n9601), .A3(n9600), .ZN(n13158) );
  NOR2_X1 U7853 ( .A1(n13169), .A2(n8101), .ZN(n8100) );
  INV_X1 U7854 ( .A(n9925), .ZN(n8101) );
  OR2_X1 U7855 ( .A1(n13183), .A2(n7672), .ZN(n13181) );
  AND2_X1 U7856 ( .A1(n10217), .A2(n10054), .ZN(n12350) );
  NAND2_X1 U7857 ( .A1(n12159), .A2(n12175), .ZN(n12158) );
  AND2_X1 U7858 ( .A1(n9814), .A2(n9813), .ZN(n10053) );
  NAND2_X1 U7859 ( .A1(n9675), .A2(n10405), .ZN(n7640) );
  NAND2_X1 U7860 ( .A1(n9664), .A2(n15075), .ZN(n7639) );
  NAND2_X1 U7861 ( .A1(n10008), .A2(n10007), .ZN(n10120) );
  XNOR2_X1 U7862 ( .A(n10075), .B(P3_IR_REG_26__SCAN_IN), .ZN(n10095) );
  OR2_X1 U7863 ( .A1(n10067), .A2(n9879), .ZN(n10075) );
  OR2_X1 U7864 ( .A1(n10066), .A2(n7776), .ZN(n7775) );
  NAND2_X1 U7865 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n7776) );
  OAI21_X1 U7866 ( .B1(n9613), .B2(n9612), .A(n7736), .ZN(n9617) );
  NOR2_X1 U7867 ( .A1(n7731), .A2(n14243), .ZN(n7730) );
  INV_X1 U7868 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10093) );
  OAI21_X1 U7869 ( .B1(n10092), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10094) );
  INV_X1 U7870 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10021) );
  XNOR2_X1 U7871 ( .A(n9560), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9918) );
  AOI21_X1 U7872 ( .B1(n7700), .B2(n7697), .A(n7348), .ZN(n7696) );
  OR2_X1 U7873 ( .A1(n9876), .A2(n7698), .ZN(n7695) );
  INV_X1 U7874 ( .A(n7702), .ZN(n7701) );
  NOR2_X1 U7875 ( .A1(n7706), .A2(n7707), .ZN(n7704) );
  INV_X1 U7876 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9545) );
  XNOR2_X1 U7877 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9748) );
  INV_X1 U7878 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9535) );
  XNOR2_X1 U7879 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9732) );
  NAND2_X1 U7880 ( .A1(n9534), .A2(n9533), .ZN(n9733) );
  AOI21_X1 U7881 ( .B1(n8060), .B2(n7477), .A(n7476), .ZN(n7475) );
  INV_X1 U7882 ( .A(n12727), .ZN(n7476) );
  INV_X1 U7883 ( .A(n12558), .ZN(n7477) );
  AND2_X1 U7884 ( .A1(n12482), .A2(n11279), .ZN(n11280) );
  NOR2_X1 U7885 ( .A1(n7455), .A2(n7458), .ZN(n7454) );
  INV_X1 U7886 ( .A(n7461), .ZN(n7458) );
  INV_X1 U7887 ( .A(n12359), .ZN(n7455) );
  OR2_X1 U7888 ( .A1(n12309), .A2(n12303), .ZN(n8038) );
  INV_X1 U7889 ( .A(n13468), .ZN(n7466) );
  XNOR2_X1 U7890 ( .A(n12546), .B(n12545), .ZN(n13417) );
  OR2_X1 U7891 ( .A1(n11280), .A2(n8065), .ZN(n8064) );
  INV_X1 U7892 ( .A(n11283), .ZN(n8065) );
  AOI21_X1 U7893 ( .B1(n7479), .B2(n7480), .A(n7478), .ZN(n8051) );
  AND2_X1 U7894 ( .A1(n8052), .A2(n7245), .ZN(n7479) );
  INV_X1 U7895 ( .A(n11850), .ZN(n7478) );
  INV_X1 U7896 ( .A(n12524), .ZN(n8052) );
  NAND2_X1 U7897 ( .A1(n12542), .A2(n8047), .ZN(n8046) );
  AND2_X1 U7898 ( .A1(n8832), .A2(n13779), .ZN(n10720) );
  AND2_X1 U7899 ( .A1(n8715), .A2(n8714), .ZN(n13690) );
  AOI21_X1 U7900 ( .B1(n13924), .B2(n8477), .A(n8693), .ZN(n13693) );
  AND2_X1 U7901 ( .A1(n8435), .A2(n8434), .ZN(n8449) );
  NAND2_X1 U7902 ( .A1(n7814), .A2(n7811), .ZN(n13917) );
  AOI21_X1 U7903 ( .B1(n13971), .B2(n8822), .A(n7620), .ZN(n7619) );
  NAND2_X1 U7904 ( .A1(n7299), .A2(n7220), .ZN(n7602) );
  AND2_X1 U7905 ( .A1(n7255), .A2(n8580), .ZN(n7803) );
  INV_X1 U7906 ( .A(n14028), .ZN(n8817) );
  OAI21_X1 U7907 ( .B1(n7211), .B2(n7266), .A(n7222), .ZN(n7629) );
  NAND2_X1 U7908 ( .A1(n8542), .A2(n7241), .ZN(n14081) );
  AND2_X1 U7909 ( .A1(n13767), .A2(n8514), .ZN(n7817) );
  NAND2_X1 U7910 ( .A1(n12184), .A2(n8514), .ZN(n12383) );
  OR2_X1 U7911 ( .A1(n12182), .A2(n12186), .ZN(n12184) );
  INV_X1 U7912 ( .A(n13766), .ZN(n12186) );
  AND2_X1 U7913 ( .A1(n13762), .A2(n8806), .ZN(n7631) );
  NAND2_X1 U7914 ( .A1(n7622), .A2(n7623), .ZN(n8132) );
  NAND2_X1 U7915 ( .A1(n7624), .A2(n8804), .ZN(n7623) );
  NOR2_X1 U7916 ( .A1(n13759), .A2(n7626), .ZN(n7625) );
  NAND2_X1 U7917 ( .A1(n8132), .A2(n13761), .ZN(n11805) );
  INV_X1 U7918 ( .A(n7624), .ZN(n7627) );
  NAND2_X1 U7919 ( .A1(n11615), .A2(n11614), .ZN(n11613) );
  NAND2_X1 U7920 ( .A1(n8412), .A2(n8411), .ZN(n11612) );
  INV_X1 U7921 ( .A(n7605), .ZN(n7610) );
  NAND2_X1 U7922 ( .A1(n7243), .A2(n8798), .ZN(n7609) );
  NAND2_X1 U7923 ( .A1(n11445), .A2(n7783), .ZN(n11417) );
  AND2_X1 U7924 ( .A1(n13758), .A2(n8381), .ZN(n7783) );
  NAND2_X1 U7925 ( .A1(n11446), .A2(n11448), .ZN(n11445) );
  NAND2_X1 U7926 ( .A1(n11332), .A2(n13750), .ZN(n11334) );
  OR2_X1 U7927 ( .A1(n10973), .A2(n13529), .ZN(n10968) );
  NAND2_X1 U7928 ( .A1(n13976), .A2(n15194), .ZN(n10963) );
  NAND2_X1 U7930 ( .A1(n13707), .A2(n13706), .ZN(n13883) );
  NAND2_X1 U7931 ( .A1(n8674), .A2(n8673), .ZN(n13944) );
  NAND2_X1 U7932 ( .A1(n12477), .A2(n13704), .ZN(n7533) );
  AND3_X1 U7933 ( .A1(n12394), .A2(n12393), .A3(n12392), .ZN(n14172) );
  AND2_X1 U7934 ( .A1(n10326), .A2(n12257), .ZN(n10700) );
  NAND2_X1 U7935 ( .A1(n8741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8744) );
  INV_X1 U7936 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8223) );
  NOR2_X1 U7937 ( .A1(n14267), .A2(n8087), .ZN(n8086) );
  INV_X1 U7938 ( .A(n8133), .ZN(n8087) );
  NAND2_X1 U7939 ( .A1(n14341), .A2(n12616), .ZN(n14294) );
  NAND2_X1 U7940 ( .A1(n7235), .A2(n11206), .ZN(n7422) );
  NAND2_X1 U7941 ( .A1(n11205), .A2(n7235), .ZN(n7423) );
  NOR2_X1 U7942 ( .A1(n11868), .A2(n8091), .ZN(n8090) );
  INV_X1 U7943 ( .A(n8093), .ZN(n8091) );
  NAND2_X1 U7944 ( .A1(n14312), .A2(n8076), .ZN(n14274) );
  NOR2_X1 U7945 ( .A1(n14277), .A2(n8077), .ZN(n8076) );
  INV_X1 U7946 ( .A(n12654), .ZN(n8077) );
  INV_X1 U7947 ( .A(n12681), .ZN(n8085) );
  INV_X1 U7948 ( .A(n8084), .ZN(n8083) );
  OAI21_X1 U7949 ( .B1(n14304), .B2(n8085), .A(n14285), .ZN(n8084) );
  NAND2_X1 U7950 ( .A1(n9357), .A2(n8028), .ZN(n8027) );
  AOI21_X1 U7951 ( .B1(n9357), .B2(n8026), .A(n8025), .ZN(n8024) );
  INV_X1 U7952 ( .A(n9355), .ZN(n8025) );
  NOR2_X1 U7953 ( .A1(n8026), .A2(n9357), .ZN(n8023) );
  AND4_X1 U7954 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n12237)
         );
  AND4_X1 U7955 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n11633)
         );
  NAND2_X1 U7956 ( .A1(n9368), .A2(n9367), .ZN(n9460) );
  NOR3_X1 U7957 ( .A1(n14601), .A2(n14781), .A3(n7551), .ZN(n7550) );
  NAND2_X1 U7958 ( .A1(n9379), .A2(n9378), .ZN(n14558) );
  NAND2_X1 U7959 ( .A1(n7552), .A2(n14784), .ZN(n7551) );
  INV_X1 U7960 ( .A(n7553), .ZN(n7552) );
  NAND2_X1 U7961 ( .A1(n14799), .A2(n14586), .ZN(n14572) );
  XNOR2_X1 U7962 ( .A(n14579), .B(n14355), .ZN(n14574) );
  AND2_X1 U7963 ( .A1(n14619), .A2(n12463), .ZN(n14600) );
  NOR2_X1 U7964 ( .A1(n14683), .A2(n7879), .ZN(n7878) );
  INV_X1 U7965 ( .A(n12439), .ZN(n7879) );
  CLKBUF_X1 U7966 ( .A(n14675), .Z(n14676) );
  INV_X1 U7967 ( .A(n14761), .ZN(n7975) );
  INV_X1 U7968 ( .A(n7974), .ZN(n7973) );
  OAI21_X1 U7969 ( .B1(n14761), .B2(n7977), .A(n7224), .ZN(n7974) );
  NAND2_X1 U7970 ( .A1(n9170), .A2(n9169), .ZN(n12606) );
  NAND2_X1 U7971 ( .A1(n9131), .A2(n9130), .ZN(n12281) );
  OAI21_X1 U7972 ( .B1(n7985), .B2(n7982), .A(n7285), .ZN(n7981) );
  INV_X1 U7973 ( .A(n7985), .ZN(n7983) );
  NAND2_X1 U7974 ( .A1(n7980), .A2(n7979), .ZN(n12205) );
  NOR2_X1 U7975 ( .A1(n7981), .A2(n12202), .ZN(n7979) );
  NAND2_X2 U7976 ( .A1(n15526), .A2(n15536), .ZN(n14763) );
  NOR2_X1 U7977 ( .A1(n11718), .A2(n7886), .ZN(n7883) );
  NAND2_X1 U7978 ( .A1(n7885), .A2(n7233), .ZN(n7884) );
  INV_X1 U7979 ( .A(n15709), .ZN(n7885) );
  INV_X1 U7980 ( .A(n14763), .ZN(n15917) );
  NAND2_X1 U7981 ( .A1(n15917), .A2(n15537), .ZN(n11214) );
  CLKBUF_X2 U7982 ( .A(n8939), .Z(n15529) );
  INV_X1 U7983 ( .A(n14787), .ZN(n14793) );
  NAND2_X1 U7984 ( .A1(n9332), .A2(n9331), .ZN(n14817) );
  NAND2_X1 U7985 ( .A1(n9271), .A2(n9270), .ZN(n14841) );
  INV_X1 U7986 ( .A(n12435), .ZN(n15878) );
  NAND2_X1 U7987 ( .A1(n11231), .A2(n11230), .ZN(n15914) );
  OAI22_X1 U7988 ( .A1(n7203), .A2(n7907), .B1(n10360), .B2(n10461), .ZN(n7906) );
  NAND2_X1 U7989 ( .A1(n7202), .A2(n10418), .ZN(n8143) );
  NAND2_X1 U7990 ( .A1(n15771), .A2(n15744), .ZN(n15923) );
  AND2_X1 U7991 ( .A1(n10444), .A2(n10443), .ZN(n10618) );
  NOR2_X1 U7992 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7993) );
  XNOR2_X1 U7993 ( .A(n8695), .B(n8696), .ZN(n14230) );
  XNOR2_X1 U7994 ( .A(n8684), .B(n8683), .ZN(n14233) );
  INV_X1 U7995 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U7996 ( .A1(n7924), .A2(n8636), .ZN(n8652) );
  NAND2_X1 U7997 ( .A1(n8619), .A2(n7928), .ZN(n7924) );
  NAND2_X1 U7998 ( .A1(n8619), .A2(n8618), .ZN(n8638) );
  NAND2_X1 U7999 ( .A1(n8222), .A2(n7954), .ZN(n8566) );
  NAND2_X1 U8000 ( .A1(n8215), .A2(n7941), .ZN(n8516) );
  OAI21_X1 U8001 ( .B1(n8414), .B2(n7537), .A(n7534), .ZN(n8463) );
  AOI21_X1 U8002 ( .B1(n7538), .B2(n7536), .A(n7535), .ZN(n7534) );
  INV_X1 U8003 ( .A(n7538), .ZN(n7537) );
  INV_X1 U8004 ( .A(n8413), .ZN(n7536) );
  XNOR2_X1 U8005 ( .A(n8433), .B(n8432), .ZN(n10512) );
  NAND2_X1 U8006 ( .A1(n7451), .A2(n7449), .ZN(n8399) );
  AOI21_X1 U8007 ( .B1(n7238), .B2(n7938), .A(n7450), .ZN(n7449) );
  INV_X1 U8008 ( .A(n8396), .ZN(n7450) );
  INV_X1 U8009 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8080) );
  INV_X1 U8010 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8078) );
  INV_X1 U8011 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U8012 ( .A(n15221), .B(n15220), .ZN(n15218) );
  NAND2_X1 U8013 ( .A1(n7389), .A2(n7388), .ZN(n7387) );
  NAND2_X1 U8014 ( .A1(n15230), .A2(n13817), .ZN(n7388) );
  INV_X1 U8015 ( .A(n15229), .ZN(n7389) );
  NAND2_X1 U8016 ( .A1(n7910), .A2(n15245), .ZN(n15246) );
  NAND2_X1 U8017 ( .A1(n15243), .A2(n15244), .ZN(n7910) );
  NAND2_X1 U8018 ( .A1(n7391), .A2(n15366), .ZN(n15257) );
  OAI21_X1 U8019 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15273), .A(n15272), .ZN(
        n15275) );
  OAI21_X1 U8020 ( .B1(n15288), .B2(n15287), .A(n15286), .ZN(n15294) );
  AND3_X1 U8021 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n11987) );
  NAND2_X1 U8022 ( .A1(n7372), .A2(n7371), .ZN(n10919) );
  INV_X1 U8023 ( .A(n10767), .ZN(n7371) );
  INV_X1 U8024 ( .A(n10768), .ZN(n7372) );
  AND4_X1 U8025 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(n13199)
         );
  NAND2_X1 U8026 ( .A1(n12174), .A2(n12173), .ZN(n12349) );
  INV_X1 U8027 ( .A(n11686), .ZN(n15647) );
  NAND2_X1 U8028 ( .A1(n11041), .A2(n11040), .ZN(n11182) );
  NAND2_X1 U8029 ( .A1(n7758), .A2(n7272), .ZN(n7757) );
  AND2_X1 U8030 ( .A1(n10784), .A2(n13143), .ZN(n15128) );
  NAND2_X1 U8031 ( .A1(n10772), .A2(n10771), .ZN(n15131) );
  NAND2_X1 U8032 ( .A1(n11034), .A2(n11357), .ZN(n12900) );
  NAND2_X1 U8033 ( .A1(n10850), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7488) );
  NOR2_X1 U8034 ( .A1(n13028), .A2(n7242), .ZN(n13019) );
  NAND2_X1 U8035 ( .A1(n7497), .A2(n7496), .ZN(n7495) );
  INV_X1 U8036 ( .A(n13043), .ZN(n7496) );
  NAND2_X1 U8037 ( .A1(n7498), .A2(n15515), .ZN(n7497) );
  OR2_X1 U8038 ( .A1(n13055), .A2(n9998), .ZN(n13070) );
  NAND2_X1 U8039 ( .A1(n7648), .A2(n13136), .ZN(n13148) );
  INV_X1 U8040 ( .A(n13150), .ZN(n7648) );
  NAND2_X1 U8041 ( .A1(n9586), .A2(n9585), .ZN(n13147) );
  OR2_X1 U8042 ( .A1(n10783), .A2(n10782), .ZN(n13143) );
  NAND2_X1 U8043 ( .A1(n7651), .A2(n10058), .ZN(n13088) );
  NAND2_X1 U8044 ( .A1(n9836), .A2(n9835), .ZN(n13390) );
  AND2_X1 U8045 ( .A1(n10804), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13393) );
  INV_X1 U8046 ( .A(n13032), .ZN(n13029) );
  OR2_X1 U8047 ( .A1(n12498), .A2(n12294), .ZN(n12295) );
  OAI21_X1 U8048 ( .B1(n11837), .B2(n11836), .A(n12577), .ZN(n12582) );
  NAND2_X1 U8049 ( .A1(n7481), .A2(n7263), .ZN(n13447) );
  NAND2_X1 U8050 ( .A1(n8533), .A2(n8532), .ZN(n13635) );
  NAND2_X1 U8051 ( .A1(n8569), .A2(n8568), .ZN(n14146) );
  NAND2_X1 U8052 ( .A1(n7381), .A2(n13976), .ZN(n14089) );
  XNOR2_X1 U8053 ( .A(n13888), .B(n7382), .ZN(n7381) );
  AOI21_X1 U8054 ( .B1(n8842), .B2(n14074), .A(n8841), .ZN(n14098) );
  NAND2_X1 U8055 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  OR2_X1 U8056 ( .A1(n7810), .A2(n7807), .ZN(n7805) );
  OR2_X1 U8057 ( .A1(n13931), .A2(n7806), .ZN(n7804) );
  AND2_X1 U8058 ( .A1(n13906), .A2(n13905), .ZN(n14102) );
  NAND2_X1 U8059 ( .A1(n7524), .A2(n8649), .ZN(n13967) );
  NAND2_X1 U8060 ( .A1(n13970), .A2(n13971), .ZN(n7524) );
  INV_X1 U8061 ( .A(n14195), .ZN(n13965) );
  AOI21_X1 U8062 ( .B1(n8816), .B2(n7630), .A(n7211), .ZN(n14053) );
  NAND2_X1 U8063 ( .A1(n8523), .A2(n8522), .ZN(n13626) );
  INV_X1 U8064 ( .A(n14200), .ZN(n14126) );
  NAND2_X1 U8065 ( .A1(n14089), .A2(n14091), .ZN(n14173) );
  AND2_X1 U8066 ( .A1(n8705), .A2(n8704), .ZN(n14183) );
  OR2_X1 U8067 ( .A1(n10329), .A2(n10587), .ZN(n8272) );
  AND2_X1 U8068 ( .A1(n7226), .A2(n8245), .ZN(n7796) );
  NOR2_X1 U8069 ( .A1(n10440), .A2(n14889), .ZN(n9498) );
  OAI21_X1 U8070 ( .B1(n14330), .B2(n7437), .A(n7434), .ZN(n14246) );
  NAND2_X1 U8071 ( .A1(n7433), .A2(n14332), .ZN(n14247) );
  NAND2_X1 U8072 ( .A1(n14323), .A2(n8133), .ZN(n14266) );
  NAND2_X1 U8073 ( .A1(n7432), .A2(n7431), .ZN(n12712) );
  AOI21_X1 U8074 ( .B1(n7434), .B2(n7437), .A(n12705), .ZN(n7431) );
  AND4_X1 U8075 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n12409)
         );
  NAND2_X1 U8076 ( .A1(n10360), .A2(n14900), .ZN(n8936) );
  NAND2_X1 U8077 ( .A1(n14314), .A2(n14313), .ZN(n14312) );
  AND4_X1 U8078 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n11764)
         );
  INV_X1 U8079 ( .A(n12667), .ZN(n14359) );
  INV_X1 U8080 ( .A(n9460), .ZN(n14781) );
  NAND2_X1 U8081 ( .A1(n9219), .A2(n9218), .ZN(n15932) );
  AND2_X1 U8082 ( .A1(n9199), .A2(n9198), .ZN(n14775) );
  INV_X1 U8083 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11399) );
  XNOR2_X1 U8084 ( .A(n15218), .B(n7412), .ZN(n15372) );
  XNOR2_X1 U8085 ( .A(n7390), .B(n7387), .ZN(n15235) );
  INV_X1 U8086 ( .A(n15233), .ZN(n7390) );
  XNOR2_X1 U8087 ( .A(n7912), .B(n15246), .ZN(n15248) );
  INV_X1 U8088 ( .A(n15247), .ZN(n7912) );
  OAI211_X1 U8089 ( .C1(n7406), .C2(n15267), .A(n7402), .B(n7405), .ZN(n15268)
         );
  NOR2_X1 U8090 ( .A1(n7404), .A2(n7909), .ZN(n7403) );
  NOR2_X1 U8091 ( .A1(n15303), .A2(n7230), .ZN(n7399) );
  OR2_X1 U8092 ( .A1(n15302), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7400) );
  OR2_X1 U8093 ( .A1(n15302), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U8094 ( .A1(n7230), .A2(n7398), .ZN(n7397) );
  NAND2_X1 U8095 ( .A1(n15303), .A2(n7230), .ZN(n7395) );
  NAND2_X1 U8096 ( .A1(n15347), .A2(n7407), .ZN(n15358) );
  NOR2_X1 U8097 ( .A1(n15355), .A2(n7408), .ZN(n7407) );
  INV_X1 U8098 ( .A(n15348), .ZN(n7408) );
  NAND2_X1 U8099 ( .A1(n8962), .A2(n9268), .ZN(n8963) );
  NAND2_X1 U8100 ( .A1(n13541), .A2(n13543), .ZN(n7819) );
  NAND2_X1 U8101 ( .A1(n13555), .A2(n13558), .ZN(n7855) );
  NOR2_X1 U8102 ( .A1(n13555), .A2(n13558), .ZN(n7856) );
  NAND2_X1 U8103 ( .A1(n13566), .A2(n13565), .ZN(n13570) );
  NOR2_X1 U8104 ( .A1(n7839), .A2(n13577), .ZN(n7840) );
  NAND2_X1 U8105 ( .A1(n7839), .A2(n13577), .ZN(n7838) );
  INV_X1 U8106 ( .A(n13584), .ZN(n7837) );
  NAND2_X1 U8107 ( .A1(n7380), .A2(n7379), .ZN(n9081) );
  NAND2_X1 U8108 ( .A1(n9066), .A2(n9068), .ZN(n7379) );
  INV_X1 U8109 ( .A(n9099), .ZN(n8005) );
  NAND2_X1 U8110 ( .A1(n13588), .A2(n13590), .ZN(n7827) );
  NAND2_X1 U8111 ( .A1(n8003), .A2(n9116), .ZN(n8002) );
  NAND2_X1 U8112 ( .A1(n7219), .A2(n8004), .ZN(n8003) );
  OR2_X1 U8113 ( .A1(n9101), .A2(n8005), .ZN(n8004) );
  OAI22_X1 U8114 ( .A1(n9133), .A2(n7996), .B1(n9134), .B2(n7997), .ZN(n9152)
         );
  AND2_X1 U8115 ( .A1(n9134), .A2(n7997), .ZN(n7996) );
  INV_X1 U8116 ( .A(n9132), .ZN(n7997) );
  NAND2_X1 U8117 ( .A1(n7378), .A2(n7377), .ZN(n9189) );
  NAND2_X1 U8118 ( .A1(n9171), .A2(n9173), .ZN(n7377) );
  AOI21_X1 U8119 ( .B1(n7846), .B2(n7844), .A(n7843), .ZN(n7842) );
  NAND2_X1 U8120 ( .A1(n7374), .A2(n7373), .ZN(n9222) );
  NAND2_X1 U8121 ( .A1(n9207), .A2(n9209), .ZN(n7373) );
  NAND2_X1 U8122 ( .A1(n13636), .A2(n13638), .ZN(n7825) );
  NAND2_X1 U8123 ( .A1(n9278), .A2(n8018), .ZN(n8015) );
  AND2_X1 U8124 ( .A1(n14701), .A2(n8017), .ZN(n8016) );
  NAND2_X1 U8125 ( .A1(n8019), .A2(n9269), .ZN(n8017) );
  INV_X1 U8126 ( .A(n10263), .ZN(n7368) );
  AOI21_X1 U8127 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7831) );
  INV_X1 U8128 ( .A(n13654), .ZN(n7832) );
  AND2_X1 U8129 ( .A1(n7865), .A2(n13682), .ZN(n7864) );
  NAND2_X1 U8130 ( .A1(n7866), .A2(n7868), .ZN(n7865) );
  NAND2_X1 U8131 ( .A1(n8010), .A2(n8013), .ZN(n8007) );
  NAND2_X1 U8132 ( .A1(n7940), .A2(SI_16_), .ZN(n7542) );
  INV_X1 U8133 ( .A(n8529), .ZN(n7544) );
  NAND2_X1 U8134 ( .A1(n10018), .A2(n10275), .ZN(n7722) );
  AOI21_X1 U8135 ( .B1(n7683), .B2(n7681), .A(n7680), .ZN(n7679) );
  INV_X1 U8136 ( .A(n10282), .ZN(n7680) );
  INV_X1 U8137 ( .A(n7684), .ZN(n7681) );
  NAND2_X1 U8138 ( .A1(n12923), .A2(n15613), .ZN(n10176) );
  INV_X1 U8139 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9547) );
  INV_X1 U8140 ( .A(n7693), .ZN(n7692) );
  OAI21_X1 U8141 ( .B1(n9794), .B2(n7694), .A(n9808), .ZN(n7693) );
  INV_X1 U8142 ( .A(n9546), .ZN(n7694) );
  NAND2_X1 U8143 ( .A1(n7851), .A2(n7849), .ZN(n7848) );
  INV_X1 U8144 ( .A(n7864), .ZN(n7863) );
  AND2_X1 U8145 ( .A1(n13724), .A2(n13725), .ZN(n7951) );
  INV_X1 U8146 ( .A(n12595), .ZN(n7418) );
  NAND2_X1 U8147 ( .A1(n10910), .A2(n11223), .ZN(n8908) );
  NAND2_X1 U8148 ( .A1(n9392), .A2(n11230), .ZN(n9380) );
  INV_X1 U8149 ( .A(n8636), .ZN(n7927) );
  NOR2_X1 U8150 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7439) );
  NAND2_X1 U8151 ( .A1(n7541), .A2(n7540), .ZN(n8220) );
  AOI21_X1 U8152 ( .B1(n7214), .B2(n7543), .A(n7336), .ZN(n7540) );
  NAND2_X1 U8153 ( .A1(n8214), .A2(n7214), .ZN(n7541) );
  NOR2_X1 U8154 ( .A1(n7940), .A2(SI_16_), .ZN(n7543) );
  OAI21_X1 U8155 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15329), .A(n15328), .ZN(
        n15340) );
  AND2_X1 U8156 ( .A1(n12875), .A2(n7745), .ZN(n7744) );
  OR2_X1 U8157 ( .A1(n12836), .A2(n7746), .ZN(n7745) );
  INV_X1 U8158 ( .A(n12753), .ZN(n7746) );
  AND2_X1 U8159 ( .A1(n12763), .A2(n13137), .ZN(n7762) );
  AND2_X1 U8160 ( .A1(n7686), .A2(n7677), .ZN(n7676) );
  NAND2_X1 U8161 ( .A1(n7679), .A2(n7682), .ZN(n7677) );
  NOR2_X1 U8162 ( .A1(n10284), .A2(n10146), .ZN(n7686) );
  INV_X1 U8163 ( .A(n7683), .ZN(n7682) );
  INV_X1 U8164 ( .A(n7679), .ZN(n7674) );
  OAI21_X1 U8165 ( .B1(n15405), .B2(n15794), .A(n15407), .ZN(n12979) );
  NAND2_X1 U8166 ( .A1(n15402), .A2(n7328), .ZN(n12932) );
  NAND2_X1 U8167 ( .A1(n15471), .A2(n12985), .ZN(n12986) );
  AOI22_X1 U8168 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12988), .B1(n15508), 
        .B2(n15512), .ZN(n13013) );
  AND2_X1 U8169 ( .A1(n13068), .A2(n9987), .ZN(n8128) );
  NOR2_X1 U8170 ( .A1(n8116), .A2(n9816), .ZN(n8115) );
  NAND2_X1 U8171 ( .A1(n9816), .A2(n8116), .ZN(n8118) );
  AND2_X1 U8172 ( .A1(n13089), .A2(n7653), .ZN(n7652) );
  NAND2_X1 U8173 ( .A1(n7654), .A2(n10058), .ZN(n7653) );
  INV_X1 U8174 ( .A(n10155), .ZN(n7654) );
  INV_X1 U8175 ( .A(n12175), .ZN(n7661) );
  NOR2_X1 U8176 ( .A1(n7662), .A2(n7658), .ZN(n7657) );
  INV_X1 U8177 ( .A(n10208), .ZN(n7658) );
  INV_X1 U8178 ( .A(n10213), .ZN(n7662) );
  AND2_X1 U8179 ( .A1(n8130), .A2(n9580), .ZN(n8129) );
  INV_X1 U8180 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9580) );
  INV_X1 U8181 ( .A(n7727), .ZN(n7726) );
  OAI21_X1 U8182 ( .B1(n9620), .B2(n7728), .A(n9972), .ZN(n7727) );
  INV_X1 U8183 ( .A(n9957), .ZN(n7728) );
  INV_X1 U8184 ( .A(n7734), .ZN(n7731) );
  AND2_X1 U8185 ( .A1(n9611), .A2(n7737), .ZN(n7736) );
  INV_X1 U8186 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9610) );
  AOI21_X1 U8187 ( .B1(n9874), .B2(n9557), .A(n7334), .ZN(n7700) );
  INV_X1 U8188 ( .A(n9557), .ZN(n7697) );
  AND2_X1 U8189 ( .A1(n9878), .A2(n9877), .ZN(n9891) );
  OR2_X1 U8190 ( .A1(n9746), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9766) );
  AND2_X1 U8191 ( .A1(n9524), .A2(n9522), .ZN(n7708) );
  NAND2_X1 U8192 ( .A1(n9649), .A2(n9648), .ZN(n9523) );
  NOR2_X1 U8193 ( .A1(n7190), .A2(n8055), .ZN(n8054) );
  NOR2_X1 U8194 ( .A1(n8536), .A2(n8535), .ZN(n8534) );
  AND2_X1 U8195 ( .A1(n8534), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8241) );
  AND2_X1 U8196 ( .A1(n8675), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8688) );
  AND2_X1 U8197 ( .A1(n7253), .A2(n14183), .ZN(n7584) );
  AND2_X1 U8198 ( .A1(n13951), .A2(n7526), .ZN(n7525) );
  NAND2_X1 U8199 ( .A1(n7527), .A2(n8649), .ZN(n7526) );
  INV_X1 U8200 ( .A(n8649), .ZN(n7528) );
  INV_X1 U8201 ( .A(n13932), .ZN(n7620) );
  NOR2_X1 U8202 ( .A1(n8659), .A2(n13463), .ZN(n8675) );
  NOR2_X1 U8203 ( .A1(n14045), .A2(n14146), .ZN(n7588) );
  NOR2_X1 U8204 ( .A1(n11819), .A2(n13603), .ZN(n7578) );
  AND2_X1 U8205 ( .A1(n7788), .A2(n13760), .ZN(n7787) );
  OR2_X1 U8206 ( .A1(n13759), .A2(n7789), .ZN(n7788) );
  INV_X1 U8207 ( .A(n8431), .ZN(n7789) );
  AND2_X1 U8208 ( .A1(n8404), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8423) );
  INV_X1 U8209 ( .A(n8328), .ZN(n7782) );
  NOR2_X1 U8210 ( .A1(n7782), .A2(n7781), .ZN(n7780) );
  INV_X1 U8211 ( .A(n8311), .ZN(n7781) );
  NAND2_X1 U8212 ( .A1(n7196), .A2(n7586), .ZN(n14008) );
  NAND2_X1 U8213 ( .A1(n12185), .A2(n12186), .ZN(n7594) );
  INV_X1 U8214 ( .A(n7578), .ZN(n12009) );
  INV_X1 U8215 ( .A(n7617), .ZN(n7613) );
  AND2_X1 U8216 ( .A1(n8035), .A2(n8234), .ZN(n7615) );
  OR2_X1 U8217 ( .A1(n8384), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8400) );
  OR2_X1 U8218 ( .A1(n8370), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8384) );
  INV_X1 U8219 ( .A(n11206), .ZN(n7425) );
  INV_X1 U8220 ( .A(n12622), .ZN(n8075) );
  INV_X1 U8221 ( .A(n15898), .ZN(n8072) );
  INV_X1 U8222 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U8223 ( .A1(n14790), .A2(n7554), .ZN(n7553) );
  AOI21_X1 U8224 ( .B1(n7892), .B2(n7210), .A(n7294), .ZN(n7891) );
  NOR2_X1 U8225 ( .A1(n14599), .A2(n7894), .ZN(n7892) );
  NOR2_X1 U8226 ( .A1(n7213), .A2(n12442), .ZN(n7894) );
  NOR2_X1 U8227 ( .A1(n15953), .A2(n15932), .ZN(n7564) );
  NOR2_X1 U8228 ( .A1(n15707), .A2(n7558), .ZN(n7561) );
  NAND2_X1 U8229 ( .A1(n7559), .A2(n12103), .ZN(n7558) );
  INV_X1 U8230 ( .A(n7233), .ZN(n7882) );
  NOR2_X1 U8231 ( .A1(n15781), .A2(n15742), .ZN(n7559) );
  AOI21_X1 U8232 ( .B1(n7896), .B2(n7902), .A(n7227), .ZN(n7895) );
  OR2_X1 U8233 ( .A1(n15706), .A2(n11763), .ZN(n15707) );
  NOR2_X1 U8234 ( .A1(n11503), .A2(n15527), .ZN(n11513) );
  INV_X1 U8235 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U8236 ( .A1(n8684), .A2(n8683), .ZN(n7942) );
  NOR2_X1 U8237 ( .A1(n8637), .A2(n7929), .ZN(n7928) );
  INV_X1 U8238 ( .A(n8618), .ZN(n7929) );
  NAND2_X1 U8239 ( .A1(n8465), .A2(n8206), .ZN(n8485) );
  XNOR2_X1 U8240 ( .A(n8207), .B(SI_14_), .ZN(n8484) );
  NOR2_X1 U8241 ( .A1(n7932), .A2(n7539), .ZN(n7538) );
  INV_X1 U8242 ( .A(n8197), .ZN(n7539) );
  INV_X1 U8243 ( .A(n7933), .ZN(n7932) );
  INV_X1 U8244 ( .A(n7930), .ZN(n7535) );
  AOI21_X1 U8245 ( .B1(n7933), .B2(n7931), .A(n7284), .ZN(n7930) );
  INV_X1 U8246 ( .A(n8200), .ZN(n7931) );
  OR2_X1 U8247 ( .A1(n9062), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9076) );
  INV_X1 U8248 ( .A(n7919), .ZN(n15238) );
  OAI21_X1 U8249 ( .B1(n15232), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7283), .ZN(
        n7919) );
  OAI22_X1 U8250 ( .A1(n15256), .A2(n15255), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n15254), .ZN(n15261) );
  OAI21_X1 U8251 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15307), .A(n15306), .ZN(
        n15309) );
  INV_X1 U8252 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15015) );
  INV_X1 U8253 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15090) );
  INV_X1 U8254 ( .A(n7761), .ZN(n12847) );
  NAND2_X1 U8255 ( .A1(n9951), .A2(n15015), .ZN(n9603) );
  NAND2_X1 U8256 ( .A1(n9757), .A2(n9756), .ZN(n9775) );
  OR2_X1 U8257 ( .A1(n9775), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9788) );
  OR2_X1 U8258 ( .A1(n9788), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U8259 ( .A1(n12750), .A2(n12836), .ZN(n12839) );
  NAND2_X1 U8260 ( .A1(n12819), .A2(n7759), .ZN(n7758) );
  INV_X1 U8261 ( .A(n7764), .ZN(n7759) );
  INV_X1 U8262 ( .A(n7772), .ZN(n7771) );
  AOI21_X1 U8263 ( .B1(n7770), .B2(n7772), .A(n7333), .ZN(n7769) );
  NOR2_X1 U8264 ( .A1(n12777), .A2(n7773), .ZN(n7772) );
  NAND2_X1 U8265 ( .A1(n10881), .A2(n10882), .ZN(n10880) );
  AOI21_X1 U8266 ( .B1(n7487), .B2(n10817), .A(n7489), .ZN(n10866) );
  NAND2_X1 U8267 ( .A1(n10850), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U8268 ( .A1(n11156), .A2(n11157), .ZN(n11158) );
  NAND2_X1 U8269 ( .A1(n15390), .A2(n12930), .ZN(n15404) );
  NAND2_X1 U8270 ( .A1(n15404), .A2(n15403), .ZN(n15402) );
  XNOR2_X1 U8271 ( .A(n12932), .B(n15419), .ZN(n15421) );
  XNOR2_X1 U8272 ( .A(n12934), .B(n15450), .ZN(n15452) );
  NAND2_X1 U8273 ( .A1(n15452), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n15451) );
  XNOR2_X1 U8274 ( .A(n12986), .B(n12936), .ZN(n15487) );
  INV_X1 U8275 ( .A(n12962), .ZN(n12963) );
  NAND2_X1 U8276 ( .A1(n9891), .A2(n9890), .ZN(n9906) );
  INV_X1 U8277 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9890) );
  AND2_X1 U8278 ( .A1(n7493), .A2(n7492), .ZN(n12999) );
  NAND2_X1 U8279 ( .A1(n12988), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7492) );
  XNOR2_X1 U8280 ( .A(n7499), .B(n13039), .ZN(n7498) );
  NAND2_X1 U8281 ( .A1(n13034), .A2(n13033), .ZN(n7499) );
  NAND2_X1 U8282 ( .A1(n13078), .A2(n8128), .ZN(n13062) );
  AND2_X1 U8283 ( .A1(n8123), .A2(n8125), .ZN(n13104) );
  NOR2_X1 U8284 ( .A1(n9932), .A2(n9588), .ZN(n9949) );
  NAND2_X1 U8285 ( .A1(n9896), .A2(n9587), .ZN(n9911) );
  NAND2_X1 U8286 ( .A1(n7643), .A2(n13223), .ZN(n7641) );
  NAND2_X1 U8287 ( .A1(n12263), .A2(n9843), .ZN(n12262) );
  AND2_X1 U8288 ( .A1(n10055), .A2(n10218), .ZN(n12267) );
  AND4_X1 U8289 ( .A1(n9829), .A2(n9828), .A3(n9827), .A4(n9826), .ZN(n12780)
         );
  AND3_X1 U8290 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(n10052) );
  NAND2_X1 U8291 ( .A1(n11997), .A2(n12138), .ZN(n11996) );
  OR2_X1 U8292 ( .A1(n11855), .A2(n9774), .ZN(n8109) );
  NAND2_X1 U8293 ( .A1(n11541), .A2(n8121), .ZN(n11663) );
  AND2_X1 U8294 ( .A1(n7304), .A2(n9695), .ZN(n8121) );
  AND4_X1 U8295 ( .A1(n9745), .A2(n9744), .A3(n9743), .A4(n9742), .ZN(n11879)
         );
  OR2_X1 U8296 ( .A1(n9711), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9723) );
  INV_X1 U8297 ( .A(n7634), .ZN(n10175) );
  AND2_X1 U8298 ( .A1(n11541), .A2(n9695), .ZN(n11682) );
  NAND2_X1 U8299 ( .A1(n10161), .A2(n10160), .ZN(n15549) );
  AND2_X1 U8300 ( .A1(n10152), .A2(n10154), .ZN(n13089) );
  AOI21_X1 U8301 ( .B1(n13085), .B2(n10011), .A(n9984), .ZN(n13091) );
  AOI21_X1 U8302 ( .B1(n13112), .B2(n10011), .A(n9630), .ZN(n13128) );
  NAND2_X1 U8303 ( .A1(n7670), .A2(n7668), .ZN(n13154) );
  AOI21_X1 U8304 ( .B1(n7218), .B2(n7672), .A(n7669), .ZN(n7668) );
  INV_X1 U8305 ( .A(n13155), .ZN(n13153) );
  OR2_X1 U8306 ( .A1(n10257), .A2(n10256), .ZN(n13155) );
  NAND2_X1 U8307 ( .A1(n9926), .A2(n9925), .ZN(n13168) );
  AND2_X1 U8308 ( .A1(n10064), .A2(n10105), .ZN(n15733) );
  NAND2_X1 U8309 ( .A1(n15733), .A2(n15732), .ZN(n15802) );
  NAND2_X1 U8310 ( .A1(n9666), .A2(n9665), .ZN(n11529) );
  NAND2_X1 U8311 ( .A1(n10063), .A2(n11525), .ZN(n15797) );
  NAND2_X1 U8312 ( .A1(n9992), .A2(n9991), .ZN(n10006) );
  AOI21_X1 U8313 ( .B1(n9612), .B2(n7736), .A(n7735), .ZN(n7734) );
  NOR2_X1 U8314 ( .A1(n9611), .A2(n7737), .ZN(n7735) );
  INV_X1 U8315 ( .A(n9612), .ZN(n7738) );
  NAND2_X1 U8316 ( .A1(n9613), .A2(n7736), .ZN(n7729) );
  AND2_X1 U8317 ( .A1(n9567), .A2(n9566), .ZN(n9942) );
  AND2_X1 U8318 ( .A1(n10025), .A2(n10092), .ZN(n10165) );
  INV_X1 U8319 ( .A(n7717), .ZN(n7716) );
  XNOR2_X1 U8320 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9703) );
  XNOR2_X1 U8321 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9690) );
  XNOR2_X1 U8322 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9672) );
  AND2_X2 U8323 ( .A1(n9660), .A2(n9568), .ZN(n9570) );
  INV_X1 U8324 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9568) );
  INV_X1 U8325 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U8326 ( .A1(n9523), .A2(n9522), .ZN(n9663) );
  AND2_X1 U8327 ( .A1(n9521), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9648) );
  INV_X1 U8328 ( .A(n13808), .ZN(n12488) );
  NAND2_X1 U8329 ( .A1(n12536), .A2(n8059), .ZN(n8058) );
  INV_X1 U8330 ( .A(n12537), .ZN(n8059) );
  INV_X1 U8331 ( .A(n7483), .ZN(n7482) );
  OAI21_X1 U8332 ( .B1(n8054), .B2(n7485), .A(n7484), .ZN(n7483) );
  INV_X1 U8333 ( .A(n13474), .ZN(n7485) );
  NAND2_X1 U8334 ( .A1(n7190), .A2(n8055), .ZN(n7484) );
  AND2_X1 U8335 ( .A1(n12556), .A2(n12554), .ZN(n13456) );
  XNOR2_X1 U8336 ( .A(n11109), .B(n13544), .ZN(n12512) );
  NOR2_X1 U8337 ( .A1(n13427), .A2(n8057), .ZN(n8056) );
  INV_X1 U8338 ( .A(n8058), .ZN(n8057) );
  OR2_X1 U8339 ( .A1(n8454), .A2(n11843), .ZN(n8475) );
  OR2_X1 U8340 ( .A1(n12299), .A2(n12300), .ZN(n8039) );
  AOI21_X1 U8341 ( .B1(n7950), .B2(n13733), .A(n13732), .ZN(n13781) );
  AND2_X1 U8342 ( .A1(n8647), .A2(n8646), .ZN(n13665) );
  AND2_X1 U8343 ( .A1(n8253), .A2(n14226), .ZN(n8323) );
  AOI21_X1 U8344 ( .B1(n13822), .B2(n13820), .A(n13821), .ZN(n13819) );
  AND2_X1 U8345 ( .A1(n8449), .A2(n8448), .ZN(n8467) );
  OR2_X1 U8346 ( .A1(n8778), .A2(n8756), .ZN(n8547) );
  OR2_X1 U8347 ( .A1(n15175), .A2(n15169), .ZN(n15189) );
  AND2_X1 U8348 ( .A1(n8721), .A2(n8720), .ZN(n13688) );
  NAND2_X1 U8349 ( .A1(n7808), .A2(n7286), .ZN(n7807) );
  NAND2_X1 U8350 ( .A1(n13900), .A2(n7809), .ZN(n7808) );
  INV_X1 U8351 ( .A(n8694), .ZN(n7809) );
  AND2_X1 U8352 ( .A1(n7811), .A2(n13900), .ZN(n7810) );
  AND2_X1 U8353 ( .A1(n13962), .A2(n7584), .ZN(n13895) );
  AND2_X1 U8354 ( .A1(n13962), .A2(n7253), .ZN(n13921) );
  OR2_X1 U8355 ( .A1(n13965), .A2(n13664), .ZN(n13932) );
  OR2_X1 U8356 ( .A1(n8641), .A2(n13469), .ZN(n8659) );
  NAND2_X1 U8357 ( .A1(n13949), .A2(n8822), .ZN(n13953) );
  NAND2_X1 U8358 ( .A1(n7621), .A2(n7527), .ZN(n13949) );
  INV_X1 U8359 ( .A(n13972), .ZN(n7621) );
  INV_X1 U8360 ( .A(n7799), .ZN(n7798) );
  OAI21_X1 U8361 ( .B1(n14006), .B2(n8597), .A(n8612), .ZN(n7799) );
  OAI21_X1 U8362 ( .B1(n7598), .B2(n7600), .A(n8820), .ZN(n13991) );
  OAI21_X1 U8363 ( .B1(n7601), .B2(n7240), .A(n14006), .ZN(n7600) );
  NAND2_X1 U8364 ( .A1(n7588), .A2(n7587), .ZN(n14021) );
  INV_X1 U8365 ( .A(n7588), .ZN(n14033) );
  AND2_X1 U8366 ( .A1(n7257), .A2(n8815), .ZN(n7630) );
  AOI21_X1 U8367 ( .B1(n7595), .B2(n7597), .A(n7247), .ZN(n7592) );
  OR2_X1 U8368 ( .A1(n8475), .A2(n11935), .ZN(n8491) );
  NAND2_X1 U8369 ( .A1(n7578), .A2(n7577), .ZN(n12059) );
  NAND2_X1 U8370 ( .A1(n8483), .A2(n8482), .ZN(n12058) );
  NAND2_X1 U8371 ( .A1(n8423), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8454) );
  INV_X1 U8372 ( .A(n8792), .ZN(n7591) );
  AOI21_X1 U8373 ( .B1(n8792), .B2(n7590), .A(n7250), .ZN(n7589) );
  NAND2_X1 U8374 ( .A1(n11002), .A2(n8311), .ZN(n11332) );
  INV_X1 U8375 ( .A(n14057), .ZN(n14071) );
  INV_X1 U8376 ( .A(n13745), .ZN(n8282) );
  NAND2_X1 U8377 ( .A1(n13745), .A2(n10984), .ZN(n11320) );
  XNOR2_X1 U8378 ( .A(n13741), .B(n8832), .ZN(n8037) );
  AND2_X1 U8379 ( .A1(n13523), .A2(n10973), .ZN(n10984) );
  AOI21_X1 U8380 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n13780) );
  INV_X1 U8381 ( .A(n13688), .ZN(n14096) );
  AND2_X1 U8382 ( .A1(n10707), .A2(n11095), .ZN(n14159) );
  AND2_X1 U8383 ( .A1(n10986), .A2(n13740), .ZN(n15861) );
  INV_X1 U8384 ( .A(n15758), .ZN(n11095) );
  AND2_X1 U8385 ( .A1(n14235), .A2(n8750), .ZN(n14904) );
  NAND2_X1 U8386 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7574) );
  INV_X1 U8387 ( .A(n8244), .ZN(n7572) );
  INV_X1 U8388 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U8389 ( .A1(n8740), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8748) );
  INV_X1 U8390 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U8391 ( .A(n8764), .B(n8763), .ZN(n12257) );
  INV_X1 U8392 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8758) );
  AND2_X1 U8393 ( .A1(n8224), .A2(n8227), .ZN(n8034) );
  OR2_X1 U8394 ( .A1(n8400), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8417) );
  INV_X1 U8395 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9521) );
  NOR2_X1 U8396 ( .A1(n14255), .A2(n8069), .ZN(n8068) );
  INV_X1 U8397 ( .A(n12600), .ZN(n8069) );
  NAND2_X1 U8398 ( .A1(n12596), .A2(n12595), .ZN(n8070) );
  OR2_X1 U8399 ( .A1(n12663), .A2(n12662), .ZN(n8133) );
  NOR2_X1 U8400 ( .A1(n9245), .A2(n9244), .ZN(n9260) );
  AND2_X1 U8401 ( .A1(n14248), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U8402 ( .A1(n14332), .A2(n7436), .ZN(n7435) );
  INV_X1 U8403 ( .A(n14331), .ZN(n7436) );
  INV_X1 U8404 ( .A(n14332), .ZN(n7437) );
  NAND2_X1 U8405 ( .A1(n11864), .A2(n8094), .ZN(n8093) );
  INV_X1 U8406 ( .A(n11866), .ZN(n8094) );
  INV_X1 U8407 ( .A(n9261), .ZN(n9272) );
  NAND2_X1 U8408 ( .A1(n14294), .A2(n14295), .ZN(n14293) );
  NAND2_X1 U8409 ( .A1(n14303), .A2(n14304), .ZN(n14302) );
  AND2_X1 U8410 ( .A1(n9295), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9306) );
  OR2_X1 U8411 ( .A1(n11205), .A2(n11206), .ZN(n7430) );
  AND2_X1 U8412 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8993) );
  AOI21_X1 U8413 ( .B1(n14375), .B2(n11435), .A(n10354), .ZN(n10355) );
  NAND2_X1 U8414 ( .A1(n10353), .A2(n10352), .ZN(n10354) );
  NAND2_X1 U8415 ( .A1(n10351), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10353) );
  AOI21_X1 U8416 ( .B1(n14375), .B2(n7192), .A(n10350), .ZN(n10913) );
  NAND2_X1 U8417 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  NAND2_X1 U8418 ( .A1(n10351), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U8419 ( .A1(n10994), .A2(n15527), .ZN(n10349) );
  OAI22_X1 U8420 ( .A1(n15529), .A2(n12706), .B1(n15565), .B2(n12640), .ZN(
        n10989) );
  NAND2_X1 U8421 ( .A1(n10634), .A2(n10624), .ZN(n11260) );
  OR2_X1 U8422 ( .A1(n9233), .A2(n9232), .ZN(n9245) );
  NAND2_X1 U8423 ( .A1(n7282), .A2(n8067), .ZN(n14341) );
  AND4_X1 U8424 ( .A1(n9314), .A2(n9313), .A3(n9312), .A4(n9311), .ZN(n12673)
         );
  AND4_X1 U8425 ( .A1(n9301), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(n12667)
         );
  AND4_X1 U8426 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n12044)
         );
  NAND2_X1 U8427 ( .A1(n8946), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U8428 ( .A1(n9406), .A2(n9405), .ZN(n14579) );
  NOR2_X1 U8429 ( .A1(n14601), .A2(n7553), .ZN(n14577) );
  INV_X1 U8430 ( .A(n14579), .ZN(n14790) );
  NAND2_X1 U8431 ( .A1(n14598), .A2(n7273), .ZN(n14573) );
  AOI21_X1 U8432 ( .B1(n7962), .B2(n7960), .A(n7254), .ZN(n7959) );
  INV_X1 U8433 ( .A(n7962), .ZN(n7961) );
  NOR2_X1 U8434 ( .A1(n14630), .A2(n7963), .ZN(n7962) );
  INV_X1 U8435 ( .A(n12462), .ZN(n7963) );
  NAND2_X1 U8436 ( .A1(n14643), .A2(n14644), .ZN(n7964) );
  NOR2_X1 U8437 ( .A1(n14645), .A2(n14817), .ZN(n14633) );
  NAND2_X1 U8438 ( .A1(n7547), .A2(n14823), .ZN(n14645) );
  INV_X1 U8439 ( .A(n7547), .ZN(n14660) );
  AND2_X1 U8440 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n9272), .ZN(n9281) );
  AND2_X1 U8441 ( .A1(n15964), .A2(n15943), .ZN(n7874) );
  NAND2_X1 U8442 ( .A1(n14741), .A2(n7875), .ZN(n14728) );
  NAND2_X1 U8443 ( .A1(n7877), .A2(n7876), .ZN(n7875) );
  XNOR2_X1 U8444 ( .A(n15964), .B(n15943), .ZN(n14729) );
  NAND2_X1 U8445 ( .A1(n7967), .A2(n7965), .ZN(n14749) );
  NAND2_X1 U8446 ( .A1(n7970), .A2(n7966), .ZN(n7965) );
  INV_X1 U8447 ( .A(n12450), .ZN(n7966) );
  NAND2_X1 U8448 ( .A1(n15918), .A2(n15920), .ZN(n15916) );
  NAND2_X1 U8449 ( .A1(n9186), .A2(n9185), .ZN(n12435) );
  OR2_X1 U8450 ( .A1(n12420), .A2(n12606), .ZN(n12421) );
  NOR2_X1 U8451 ( .A1(n12087), .A2(n12281), .ZN(n12211) );
  NAND2_X1 U8452 ( .A1(n7561), .A2(n7560), .ZN(n12087) );
  AND2_X1 U8453 ( .A1(n11221), .A2(n11634), .ZN(n11266) );
  INV_X1 U8454 ( .A(n7561), .ZN(n12102) );
  NOR2_X1 U8455 ( .A1(n15707), .A2(n15742), .ZN(n15766) );
  NOR2_X1 U8456 ( .A1(n15707), .A2(n7557), .ZN(n15764) );
  INV_X1 U8457 ( .A(n7559), .ZN(n7557) );
  NAND2_X1 U8458 ( .A1(n7958), .A2(n7957), .ZN(n15705) );
  AOI21_X1 U8459 ( .B1(n15658), .B2(n11717), .A(n7287), .ZN(n7957) );
  NOR2_X1 U8460 ( .A1(n11362), .A2(n11709), .ZN(n15656) );
  INV_X1 U8461 ( .A(n15620), .ZN(n11364) );
  INV_X1 U8462 ( .A(n15903), .ZN(n14767) );
  NAND2_X1 U8463 ( .A1(n7556), .A2(n15620), .ZN(n11362) );
  CLKBUF_X1 U8464 ( .A(n11224), .Z(n9436) );
  INV_X1 U8465 ( .A(n15901), .ZN(n14765) );
  NAND2_X1 U8466 ( .A1(n9267), .A2(n9266), .ZN(n14848) );
  INV_X1 U8467 ( .A(n12606), .ZN(n15850) );
  INV_X1 U8468 ( .A(n12408), .ZN(n15843) );
  NAND2_X1 U8469 ( .A1(n7984), .A2(n7988), .ZN(n12049) );
  INV_X1 U8470 ( .A(n7987), .ZN(n7984) );
  NOR2_X1 U8471 ( .A1(n7987), .A2(n7985), .ZN(n15807) );
  INV_X1 U8472 ( .A(n15923), .ZN(n15851) );
  OR2_X1 U8473 ( .A1(n11223), .A2(n11222), .ZN(n15744) );
  AND2_X1 U8474 ( .A1(n11264), .A2(n10621), .ZN(n15919) );
  INV_X1 U8475 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8868) );
  XNOR2_X1 U8476 ( .A(n9366), .B(n9365), .ZN(n13683) );
  OAI21_X1 U8477 ( .B1(n9359), .B2(n7946), .A(n7943), .ZN(n9366) );
  AND2_X1 U8478 ( .A1(n9377), .A2(n9376), .ZN(n13705) );
  NAND2_X1 U8479 ( .A1(n7949), .A2(n7947), .ZN(n9377) );
  NAND2_X1 U8480 ( .A1(n7949), .A2(n9361), .ZN(n9375) );
  XNOR2_X1 U8481 ( .A(n8719), .B(n8718), .ZN(n14227) );
  INV_X1 U8482 ( .A(n8896), .ZN(n8897) );
  XNOR2_X1 U8483 ( .A(n8602), .B(n15019), .ZN(n9279) );
  AND2_X1 U8485 ( .A1(n8546), .A2(n8545), .ZN(n11906) );
  NAND2_X1 U8486 ( .A1(n7953), .A2(n8222), .ZN(n8546) );
  NAND2_X1 U8487 ( .A1(n7546), .A2(n8215), .ZN(n8530) );
  NAND2_X1 U8488 ( .A1(n8205), .A2(n8204), .ZN(n8465) );
  INV_X1 U8489 ( .A(n8462), .ZN(n8204) );
  INV_X1 U8490 ( .A(n8463), .ZN(n8205) );
  OAI21_X1 U8491 ( .B1(n8433), .B2(n8432), .A(n8200), .ZN(n8447) );
  AND2_X1 U8492 ( .A1(n8197), .A2(n8196), .ZN(n8413) );
  AND2_X1 U8493 ( .A1(n8193), .A2(n8192), .ZN(n8396) );
  NAND2_X1 U8494 ( .A1(n7937), .A2(n7453), .ZN(n7452) );
  AOI21_X1 U8495 ( .B1(n7937), .B2(n7939), .A(n7936), .ZN(n7935) );
  INV_X1 U8496 ( .A(n8182), .ZN(n7453) );
  XNOR2_X1 U8497 ( .A(n8383), .B(n8382), .ZN(n10450) );
  NAND2_X1 U8498 ( .A1(n8369), .A2(n8186), .ZN(n8383) );
  NAND2_X1 U8499 ( .A1(n8367), .A2(n8366), .ZN(n8369) );
  AND2_X1 U8500 ( .A1(n8182), .A2(n8181), .ZN(n8350) );
  NAND2_X1 U8501 ( .A1(n8315), .A2(n8174), .ZN(n8330) );
  INV_X1 U8502 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8853) );
  INV_X1 U8503 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8981) );
  INV_X1 U8504 ( .A(n8312), .ZN(n8314) );
  NAND2_X1 U8505 ( .A1(n8301), .A2(n7262), .ZN(n8000) );
  AND2_X1 U8506 ( .A1(n7401), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15217) );
  INV_X1 U8507 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7401) );
  INV_X1 U8508 ( .A(n7913), .ZN(n15224) );
  OAI21_X1 U8509 ( .B1(n15220), .B2(n15221), .A(n7914), .ZN(n7913) );
  NAND2_X1 U8510 ( .A1(n14384), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7914) );
  AOI22_X1 U8511 ( .A1(n15252), .A2(n15251), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n15250), .ZN(n15255) );
  OR2_X1 U8512 ( .A1(n15250), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n15251) );
  INV_X1 U8513 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15254) );
  AND2_X1 U8514 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  INV_X1 U8515 ( .A(n7413), .ZN(n15301) );
  OAI21_X1 U8516 ( .B1(n15296), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7256), .ZN(
        n7413) );
  NOR2_X1 U8517 ( .A1(n15332), .A2(n7410), .ZN(n15333) );
  NAND2_X1 U8518 ( .A1(n12741), .A2(n12740), .ZN(n12778) );
  AND2_X1 U8519 ( .A1(n9609), .A2(n9608), .ZN(n13138) );
  INV_X1 U8520 ( .A(n12915), .ZN(n12157) );
  NAND2_X1 U8521 ( .A1(n11981), .A2(n11980), .ZN(n11983) );
  NAND2_X1 U8522 ( .A1(n11981), .A2(n7766), .ZN(n12136) );
  AND2_X1 U8523 ( .A1(n9967), .A2(n9966), .ZN(n13106) );
  NAND2_X1 U8524 ( .A1(n7756), .A2(n7764), .ZN(n12818) );
  NAND2_X1 U8525 ( .A1(n7761), .A2(n7760), .ZN(n7756) );
  OAI21_X1 U8526 ( .B1(n11041), .B2(n7750), .A(n7749), .ZN(n11477) );
  AND4_X1 U8527 ( .A1(n9902), .A2(n9901), .A3(n9900), .A4(n9899), .ZN(n13198)
         );
  NAND2_X1 U8528 ( .A1(n12352), .A2(n12351), .ZN(n12741) );
  XNOR2_X1 U8529 ( .A(n12765), .B(n12763), .ZN(n12867) );
  AOI21_X1 U8530 ( .B1(n7766), .B2(n11886), .A(n7332), .ZN(n7765) );
  NAND2_X1 U8531 ( .A1(n10919), .A2(n10918), .ZN(n10920) );
  NAND2_X1 U8532 ( .A1(n12839), .A2(n12753), .ZN(n12874) );
  INV_X1 U8533 ( .A(n15128), .ZN(n12887) );
  NAND2_X1 U8534 ( .A1(n10791), .A2(n10787), .ZN(n12897) );
  INV_X1 U8535 ( .A(n10317), .ZN(n7687) );
  AND2_X1 U8536 ( .A1(n10138), .A2(n10017), .ZN(n13064) );
  INV_X1 U8537 ( .A(n13106), .ZN(n12906) );
  INV_X1 U8538 ( .A(n12780), .ZN(n12913) );
  INV_X1 U8539 ( .A(n15574), .ZN(n12923) );
  NAND2_X1 U8540 ( .A1(n9682), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9634) );
  INV_X1 U8541 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15380) );
  OR2_X1 U8542 ( .A1(n9660), .A2(n9879), .ZN(n7494) );
  OAI22_X1 U8543 ( .A1(n10934), .A2(n10933), .B1(n10938), .B2(n10932), .ZN(
        n10936) );
  NAND2_X1 U8544 ( .A1(n7517), .A2(n15383), .ZN(n15401) );
  OR2_X1 U8545 ( .A1(n15385), .A2(n15381), .ZN(n7517) );
  NAND2_X1 U8546 ( .A1(n15385), .A2(n7515), .ZN(n7510) );
  NOR2_X1 U8547 ( .A1(n15457), .A2(n7500), .ZN(n15478) );
  AND2_X1 U8548 ( .A1(n12959), .A2(n15450), .ZN(n7500) );
  NAND2_X1 U8549 ( .A1(n15478), .A2(n15477), .ZN(n15476) );
  NOR2_X1 U8550 ( .A1(n15483), .A2(n12938), .ZN(n15519) );
  INV_X1 U8551 ( .A(n7493), .ZN(n15520) );
  AND2_X1 U8552 ( .A1(n10825), .A2(n10808), .ZN(n15517) );
  XNOR2_X1 U8553 ( .A(n12999), .B(n13014), .ZN(n12941) );
  NAND2_X1 U8554 ( .A1(n7506), .A2(n15505), .ZN(n12968) );
  NAND2_X1 U8555 ( .A1(n7507), .A2(n15504), .ZN(n7506) );
  NAND2_X1 U8556 ( .A1(n10041), .A2(n10040), .ZN(n13054) );
  NAND2_X1 U8557 ( .A1(n7678), .A2(n7683), .ZN(n10147) );
  NAND2_X1 U8558 ( .A1(n9615), .A2(n9614), .ZN(n13276) );
  NAND2_X1 U8559 ( .A1(n9931), .A2(n9930), .ZN(n13178) );
  NAND2_X1 U8560 ( .A1(n13222), .A2(n9887), .ZN(n13211) );
  NAND2_X1 U8561 ( .A1(n13230), .A2(n13229), .ZN(n13228) );
  NAND2_X1 U8562 ( .A1(n13244), .A2(n10228), .ZN(n13230) );
  NAND2_X1 U8563 ( .A1(n12328), .A2(n9857), .ZN(n13238) );
  NAND2_X1 U8564 ( .A1(n9817), .A2(n9816), .ZN(n12164) );
  INV_X1 U8565 ( .A(n10052), .ZN(n15798) );
  NAND2_X1 U8566 ( .A1(n8105), .A2(n8106), .ZN(n11993) );
  OR2_X1 U8567 ( .A1(n11855), .A2(n8108), .ZN(n8105) );
  NAND2_X1 U8568 ( .A1(n7665), .A2(n10201), .ZN(n11893) );
  AND3_X1 U8569 ( .A1(n9710), .A2(n9709), .A3(n9708), .ZN(n11686) );
  NAND2_X1 U8570 ( .A1(n10902), .A2(n15585), .ZN(n13250) );
  INV_X1 U8571 ( .A(n13250), .ZN(n15684) );
  INV_X1 U8572 ( .A(n13327), .ZN(n13265) );
  INV_X1 U8573 ( .A(n15839), .ZN(n15970) );
  INV_X1 U8574 ( .A(n10148), .ZN(n13319) );
  NAND2_X1 U8575 ( .A1(n10145), .A2(n10144), .ZN(n15975) );
  NAND2_X1 U8576 ( .A1(n9977), .A2(n9976), .ZN(n13326) );
  OR2_X1 U8577 ( .A1(n11815), .A2(n9946), .ZN(n9624) );
  NAND2_X1 U8578 ( .A1(n13148), .A2(n10260), .ZN(n13118) );
  NAND2_X1 U8579 ( .A1(n9948), .A2(n9947), .ZN(n13351) );
  NAND2_X1 U8580 ( .A1(n13181), .A2(n10248), .ZN(n13166) );
  AOI21_X1 U8581 ( .B1(n13183), .B2(n7672), .A(n13182), .ZN(n13366) );
  NAND2_X1 U8582 ( .A1(n9920), .A2(n9919), .ZN(n13362) );
  NAND2_X1 U8583 ( .A1(n9910), .A2(n9909), .ZN(n13369) );
  INV_X1 U8584 ( .A(n13391), .ZN(n15974) );
  NAND2_X1 U8585 ( .A1(n9882), .A2(n9881), .ZN(n13378) );
  NAND2_X1 U8586 ( .A1(n9849), .A2(n9848), .ZN(n13386) );
  NAND2_X1 U8587 ( .A1(n12158), .A2(n10213), .ZN(n12167) );
  INV_X1 U8588 ( .A(n10053), .ZN(n12280) );
  AND2_X2 U8589 ( .A1(n10101), .A2(n10100), .ZN(n15980) );
  OR2_X1 U8590 ( .A1(n15980), .A2(n15797), .ZN(n13391) );
  INV_X1 U8591 ( .A(n10106), .ZN(n13392) );
  INV_X1 U8592 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9590) );
  XNOR2_X1 U8593 ( .A(n9990), .B(n9988), .ZN(n12128) );
  INV_X1 U8594 ( .A(n10095), .ZN(n11930) );
  XNOR2_X1 U8595 ( .A(n9973), .B(n9971), .ZN(n11928) );
  INV_X1 U8596 ( .A(SI_25_), .ZN(n15017) );
  NAND2_X1 U8597 ( .A1(n7297), .A2(n10068), .ZN(n11816) );
  NAND2_X1 U8598 ( .A1(n9879), .A2(n9579), .ZN(n7774) );
  NAND2_X1 U8599 ( .A1(n10073), .A2(n10072), .ZN(n11756) );
  INV_X1 U8600 ( .A(n10063), .ZN(n11176) );
  AND2_X1 U8601 ( .A1(n10397), .A2(P3_U3151), .ZN(n11355) );
  NAND2_X1 U8602 ( .A1(n10030), .A2(n10029), .ZN(n11070) );
  NAND2_X1 U8603 ( .A1(n7699), .A2(n9557), .ZN(n9889) );
  OR2_X1 U8604 ( .A1(n9876), .A2(n9874), .ZN(n7699) );
  INV_X1 U8605 ( .A(SI_17_), .ZN(n15044) );
  INV_X1 U8606 ( .A(n13014), .ZN(n12993) );
  INV_X1 U8607 ( .A(SI_15_), .ZN(n15046) );
  INV_X1 U8608 ( .A(SI_14_), .ZN(n14943) );
  NAND2_X1 U8609 ( .A1(n9818), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U8610 ( .A1(n7691), .A2(n9546), .ZN(n9809) );
  NAND2_X1 U8611 ( .A1(n9795), .A2(n9794), .ZN(n7691) );
  INV_X1 U8612 ( .A(SI_11_), .ZN(n15057) );
  INV_X1 U8613 ( .A(SI_10_), .ZN(n14909) );
  INV_X1 U8614 ( .A(SI_9_), .ZN(n14910) );
  NAND2_X1 U8615 ( .A1(n7715), .A2(n9536), .ZN(n9750) );
  NAND2_X1 U8616 ( .A1(n9733), .A2(n9732), .ZN(n7715) );
  INV_X1 U8617 ( .A(n11050), .ZN(n11056) );
  INV_X1 U8618 ( .A(SI_5_), .ZN(n10406) );
  INV_X1 U8619 ( .A(SI_2_), .ZN(n15075) );
  NAND2_X1 U8620 ( .A1(n12723), .A2(n12722), .ZN(n13407) );
  NAND2_X1 U8621 ( .A1(n12723), .A2(n8060), .ZN(n13409) );
  NAND2_X1 U8622 ( .A1(n7468), .A2(n8147), .ZN(n13418) );
  INV_X1 U8623 ( .A(n13417), .ZN(n7468) );
  NOR2_X1 U8624 ( .A1(n11105), .A2(n10719), .ZN(n10723) );
  AND2_X1 U8625 ( .A1(n12512), .A2(n10718), .ZN(n10719) );
  NAND2_X1 U8626 ( .A1(n13496), .A2(n8058), .ZN(n13432) );
  NAND2_X1 U8627 ( .A1(n8240), .A2(n8239), .ZN(n14048) );
  NAND2_X1 U8628 ( .A1(n7475), .A2(n7472), .ZN(n7471) );
  NAND2_X1 U8629 ( .A1(n8061), .A2(n7473), .ZN(n7472) );
  NAND2_X1 U8630 ( .A1(n8060), .A2(n12731), .ZN(n7474) );
  AND2_X1 U8631 ( .A1(n7481), .A2(n7482), .ZN(n13449) );
  OR2_X1 U8632 ( .A1(n12526), .A2(n7216), .ZN(n8050) );
  OR2_X1 U8633 ( .A1(n13486), .A2(n13976), .ZN(n13484) );
  NAND2_X1 U8634 ( .A1(n7459), .A2(n7457), .ZN(n7456) );
  INV_X1 U8635 ( .A(n12365), .ZN(n7459) );
  NAND2_X1 U8636 ( .A1(n7460), .A2(n7463), .ZN(n12366) );
  INV_X1 U8637 ( .A(n8038), .ZN(n7460) );
  INV_X1 U8638 ( .A(n8147), .ZN(n7467) );
  NAND2_X1 U8639 ( .A1(n13418), .A2(n12547), .ZN(n13467) );
  AND2_X1 U8640 ( .A1(n13509), .A2(n11283), .ZN(n8066) );
  NAND2_X1 U8641 ( .A1(n8064), .A2(n8063), .ZN(n8062) );
  NAND2_X1 U8642 ( .A1(n7486), .A2(n13431), .ZN(n13476) );
  NAND2_X1 U8643 ( .A1(n13496), .A2(n8056), .ZN(n7486) );
  AOI21_X1 U8644 ( .B1(n8051), .B2(n7216), .A(n7292), .ZN(n8048) );
  NOR2_X1 U8645 ( .A1(n8043), .A2(n7331), .ZN(n8042) );
  INV_X1 U8646 ( .A(n8046), .ZN(n8043) );
  NAND2_X1 U8647 ( .A1(n8053), .A2(n12524), .ZN(n12530) );
  OR2_X1 U8648 ( .A1(n12526), .A2(n11840), .ZN(n8053) );
  XNOR2_X1 U8649 ( .A(n11849), .B(n11841), .ZN(n12524) );
  XNOR2_X1 U8650 ( .A(n10714), .B(n10713), .ZN(n11128) );
  NAND2_X1 U8651 ( .A1(n13510), .A2(n13509), .ZN(n13508) );
  NAND2_X1 U8652 ( .A1(n12493), .A2(n8039), .ZN(n12344) );
  NAND2_X1 U8653 ( .A1(n11124), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13479) );
  NAND2_X1 U8654 ( .A1(n10720), .A2(n8833), .ZN(n14055) );
  INV_X1 U8655 ( .A(n13690), .ZN(n13790) );
  INV_X1 U8656 ( .A(n10709), .ZN(n13816) );
  INV_X1 U8657 ( .A(n10973), .ZN(n13528) );
  XNOR2_X1 U8658 ( .A(n8295), .B(P2_IR_REG_2__SCAN_IN), .ZN(n13824) );
  XNOR2_X1 U8659 ( .A(n7360), .B(n11971), .ZN(n15161) );
  NAND2_X1 U8660 ( .A1(n12025), .A2(n7352), .ZN(n11974) );
  AOI21_X1 U8661 ( .B1(n15210), .B2(n15194), .A(n7358), .ZN(n7357) );
  INV_X1 U8662 ( .A(n15197), .ZN(n7358) );
  OR2_X1 U8663 ( .A1(n15198), .A2(n8154), .ZN(n7361) );
  AND2_X1 U8664 ( .A1(n10338), .A2(n14231), .ZN(n15201) );
  NAND2_X1 U8665 ( .A1(n13917), .A2(n8694), .ZN(n13893) );
  NAND2_X1 U8666 ( .A1(n13935), .A2(n8824), .ZN(n13912) );
  NAND2_X1 U8667 ( .A1(n7814), .A2(n7813), .ZN(n13919) );
  NAND2_X1 U8668 ( .A1(n7599), .A2(n7602), .ZN(n14003) );
  NAND2_X1 U8669 ( .A1(n8818), .A2(n7240), .ZN(n7599) );
  AOI21_X1 U8670 ( .B1(n8581), .B2(n7803), .A(n7802), .ZN(n14007) );
  NAND2_X1 U8671 ( .A1(n8818), .A2(n8817), .ZN(n7603) );
  NAND2_X1 U8672 ( .A1(n8581), .A2(n8580), .ZN(n14017) );
  NAND2_X1 U8673 ( .A1(n14081), .A2(n8562), .ZN(n14043) );
  NAND2_X1 U8674 ( .A1(n8542), .A2(n8541), .ZN(n14083) );
  NAND2_X1 U8675 ( .A1(n12184), .A2(n7817), .ZN(n12385) );
  NAND2_X1 U8676 ( .A1(n8505), .A2(n8504), .ZN(n13622) );
  NAND2_X1 U8677 ( .A1(n11805), .A2(n8806), .ZN(n12005) );
  NAND2_X1 U8678 ( .A1(n11613), .A2(n7627), .ZN(n11822) );
  AND2_X1 U8679 ( .A1(n11613), .A2(n8801), .ZN(n8138) );
  NAND2_X1 U8680 ( .A1(n7786), .A2(n8431), .ZN(n11817) );
  NAND2_X1 U8681 ( .A1(n11612), .A2(n13759), .ZN(n7786) );
  NAND2_X1 U8682 ( .A1(n7606), .A2(n7609), .ZN(n8131) );
  NAND2_X1 U8683 ( .A1(n8797), .A2(n7610), .ZN(n7606) );
  NAND2_X1 U8684 ( .A1(n11445), .A2(n8381), .ZN(n11415) );
  INV_X1 U8685 ( .A(n13984), .ZN(n15814) );
  INV_X1 U8686 ( .A(n14085), .ZN(n15824) );
  NAND2_X1 U8687 ( .A1(n11334), .A2(n8328), .ZN(n11133) );
  NAND2_X1 U8688 ( .A1(n15140), .A2(n8773), .ZN(n13959) );
  OR2_X1 U8689 ( .A1(n8844), .A2(n15194), .ZN(n13984) );
  INV_X1 U8690 ( .A(n13522), .ZN(n13534) );
  INV_X1 U8691 ( .A(n15821), .ZN(n14035) );
  INV_X1 U8692 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U8693 ( .A1(n7448), .A2(n8438), .ZN(n13600) );
  NAND2_X1 U8694 ( .A1(n10512), .A2(n13704), .ZN(n7448) );
  INV_X1 U8695 ( .A(n13883), .ZN(n14180) );
  NAND2_X1 U8696 ( .A1(n15870), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7531) );
  AND2_X1 U8697 ( .A1(n8687), .A2(n8686), .ZN(n14187) );
  AOI211_X1 U8698 ( .C1(n14107), .C2(n15859), .A(n14106), .B(n14105), .ZN(
        n14184) );
  INV_X1 U8699 ( .A(n13944), .ZN(n14191) );
  AND2_X1 U8700 ( .A1(n8658), .A2(n8657), .ZN(n14195) );
  AND3_X1 U8701 ( .A1(n14119), .A2(n14118), .A3(n14117), .ZN(n14192) );
  AND2_X1 U8702 ( .A1(n8640), .A2(n8639), .ZN(n14200) );
  INV_X1 U8703 ( .A(n14048), .ZN(n14213) );
  NAND2_X1 U8704 ( .A1(n8422), .A2(n8421), .ZN(n13591) );
  NAND2_X1 U8705 ( .A1(n14215), .A2(n15861), .ZN(n14219) );
  AND2_X1 U8706 ( .A1(n10700), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15140) );
  NAND2_X1 U8707 ( .A1(n8250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8247) );
  XNOR2_X1 U8708 ( .A(n8742), .B(P2_IR_REG_26__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U8709 ( .A1(n8746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U8710 ( .A1(n8746), .A2(n8745), .ZN(n14238) );
  OR2_X1 U8711 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  XNOR2_X1 U8712 ( .A(n8748), .B(n8747), .ZN(n14242) );
  XNOR2_X1 U8713 ( .A(n9279), .B(n8617), .ZN(n12477) );
  INV_X1 U8714 ( .A(n15194), .ZN(n13776) );
  INV_X1 U8715 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11907) );
  INV_X1 U8716 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11677) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10430) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10427) );
  INV_X1 U8719 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10422) );
  OR2_X1 U8720 ( .A1(n8318), .A2(n8756), .ZN(n8303) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10424) );
  XNOR2_X1 U8722 ( .A(n9391), .B(n9478), .ZN(n10623) );
  NAND2_X1 U8723 ( .A1(n8070), .A2(n12600), .ZN(n14254) );
  AND2_X1 U8724 ( .A1(n12067), .A2(n7223), .ZN(n8089) );
  NAND2_X1 U8725 ( .A1(n11865), .A2(n8093), .ZN(n11867) );
  NAND2_X1 U8726 ( .A1(n14312), .A2(n12654), .ZN(n14276) );
  NAND2_X1 U8727 ( .A1(n14302), .A2(n12681), .ZN(n14284) );
  NAND2_X1 U8728 ( .A1(n7423), .A2(n7421), .ZN(n7428) );
  AND2_X1 U8729 ( .A1(n7422), .A2(n11598), .ZN(n7421) );
  AND2_X1 U8730 ( .A1(n8092), .A2(n7223), .ZN(n12068) );
  INV_X1 U8731 ( .A(n15949), .ZN(n15963) );
  NOR2_X1 U8732 ( .A1(n14321), .A2(n7444), .ZN(n7443) );
  INV_X1 U8733 ( .A(n12658), .ZN(n7444) );
  NAND2_X1 U8734 ( .A1(n14274), .A2(n12658), .ZN(n14322) );
  OR2_X1 U8735 ( .A1(n10632), .A2(n11260), .ZN(n14326) );
  INV_X1 U8736 ( .A(n15965), .ZN(n14348) );
  CLKBUF_X1 U8737 ( .A(n15946), .Z(n15947) );
  INV_X1 U8738 ( .A(n14744), .ZN(n15943) );
  NAND2_X1 U8739 ( .A1(n11207), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15969) );
  AOI21_X1 U8740 ( .B1(n8083), .B2(n8085), .A(n7276), .ZN(n8081) );
  NAND2_X1 U8741 ( .A1(n9342), .A2(n9341), .ZN(n14810) );
  NAND2_X1 U8742 ( .A1(n8067), .A2(n12616), .ZN(n14343) );
  INV_X1 U8743 ( .A(n15969), .ZN(n14352) );
  NOR2_X1 U8744 ( .A1(n8023), .A2(n8024), .ZN(n8021) );
  AOI22_X1 U8745 ( .A1(n8023), .A2(n8029), .B1(n8024), .B2(n8027), .ZN(n8020)
         );
  AND2_X1 U8746 ( .A1(n9340), .A2(n9339), .ZN(n8022) );
  OR2_X1 U8747 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  INV_X1 U8748 ( .A(n12673), .ZN(n14663) );
  INV_X1 U8749 ( .A(n12237), .ZN(n14364) );
  INV_X1 U8750 ( .A(n11633), .ZN(n14370) );
  OR2_X1 U8751 ( .A1(n8919), .A2(n10367), .ZN(n8924) );
  INV_X1 U8752 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15240) );
  INV_X1 U8753 ( .A(n7548), .ZN(n14559) );
  AOI211_X1 U8754 ( .C1(n14601), .C2(n14781), .A(n7550), .B(n7549), .ZN(n7548)
         );
  AND2_X1 U8755 ( .A1(n7551), .A2(n14781), .ZN(n7549) );
  INV_X1 U8756 ( .A(n14558), .ZN(n14784) );
  NAND2_X1 U8757 ( .A1(n14598), .A2(n12465), .ZN(n12466) );
  AND2_X1 U8758 ( .A1(n9409), .A2(n8881), .ZN(n14603) );
  NAND2_X1 U8759 ( .A1(n14625), .A2(n12443), .ZN(n14610) );
  NAND2_X1 U8760 ( .A1(n9303), .A2(n9302), .ZN(n14670) );
  NAND2_X1 U8761 ( .A1(n14898), .A2(n10360), .ZN(n14692) );
  NAND2_X1 U8762 ( .A1(n14695), .A2(n12439), .ZN(n14682) );
  NAND2_X1 U8763 ( .A1(n7212), .A2(n7232), .ZN(n14700) );
  NAND2_X1 U8764 ( .A1(n7972), .A2(n7973), .ZN(n15910) );
  AND2_X1 U8765 ( .A1(n7972), .A2(n7969), .ZN(n15909) );
  NAND2_X1 U8766 ( .A1(n12449), .A2(n7975), .ZN(n7972) );
  NOR2_X1 U8767 ( .A1(n12449), .A2(n7976), .ZN(n14762) );
  NAND2_X1 U8768 ( .A1(n7898), .A2(n7899), .ZN(n12419) );
  NAND2_X1 U8769 ( .A1(n12203), .A2(n7901), .ZN(n7898) );
  AOI21_X1 U8770 ( .B1(n12203), .B2(n12202), .A(n7215), .ZN(n12411) );
  NOR2_X1 U8771 ( .A1(n7978), .A2(n7981), .ZN(n12086) );
  INV_X1 U8772 ( .A(n7980), .ZN(n7978) );
  NAND2_X1 U8773 ( .A1(n7884), .A2(n7883), .ZN(n12034) );
  AND2_X1 U8774 ( .A1(n7884), .A2(n11705), .ZN(n11707) );
  INV_X1 U8775 ( .A(n11763), .ZN(n15722) );
  OR2_X1 U8776 ( .A1(n15941), .A2(n11264), .ZN(n15723) );
  NAND2_X1 U8777 ( .A1(n14585), .A2(n14584), .ZN(n14772) );
  INV_X1 U8778 ( .A(n15930), .ZN(n14584) );
  OR2_X1 U8779 ( .A1(n15941), .A2(n15537), .ZN(n14672) );
  INV_X1 U8780 ( .A(n15723), .ZN(n15931) );
  AND2_X2 U8781 ( .A1(n10634), .A2(n10633), .ZN(n15930) );
  NAND2_X1 U8782 ( .A1(n14785), .A2(n15914), .ZN(n14795) );
  INV_X1 U8783 ( .A(n8882), .ZN(n8876) );
  NOR2_X1 U8784 ( .A1(n8887), .A2(n7904), .ZN(n7566) );
  NAND2_X1 U8785 ( .A1(n9488), .A2(n7279), .ZN(n7567) );
  NOR2_X1 U8786 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7904) );
  NOR2_X1 U8787 ( .A1(n9486), .A2(n9494), .ZN(n9495) );
  NAND2_X1 U8788 ( .A1(n9482), .A2(n9481), .ZN(n9485) );
  NAND2_X1 U8789 ( .A1(n9483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U8790 ( .A1(n8096), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U8791 ( .A1(n7442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8904) );
  INV_X1 U8792 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12112) );
  INV_X1 U8793 ( .A(n15537), .ZN(n12019) );
  NAND2_X1 U8794 ( .A1(n7545), .A2(n8215), .ZN(n8518) );
  INV_X1 U8795 ( .A(n7546), .ZN(n7545) );
  INV_X1 U8796 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11170) );
  AND2_X1 U8797 ( .A1(n9167), .A2(n9147), .ZN(n11021) );
  INV_X1 U8798 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10451) );
  NOR2_X1 U8799 ( .A1(n10397), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14880) );
  INV_X1 U8800 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10433) );
  AND3_X1 U8801 ( .A1(n8080), .A2(n8079), .A3(n8078), .ZN(n8915) );
  INV_X1 U8802 ( .A(n10418), .ZN(n8914) );
  NOR2_X1 U8803 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8954) );
  NAND2_X1 U8804 ( .A1(n8162), .A2(n8165), .ZN(n8268) );
  NAND2_X1 U8805 ( .A1(n7411), .A2(n15219), .ZN(n15227) );
  NAND2_X1 U8806 ( .A1(n15372), .A2(n15371), .ZN(n7411) );
  AOI21_X1 U8807 ( .B1(n7386), .B2(n7385), .A(n15236), .ZN(n15243) );
  INV_X1 U8808 ( .A(n15235), .ZN(n7386) );
  INV_X1 U8809 ( .A(n7387), .ZN(n15234) );
  XNOR2_X1 U8810 ( .A(n15242), .B(n7911), .ZN(n15244) );
  INV_X1 U8811 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U8812 ( .A1(n7392), .A2(n15249), .ZN(n15368) );
  NAND2_X1 U8813 ( .A1(n15248), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U8814 ( .A1(n15368), .A2(n15367), .ZN(n15366) );
  NAND2_X1 U8815 ( .A1(n7908), .A2(n15269), .ZN(n15278) );
  XNOR2_X1 U8816 ( .A(n15294), .B(n15295), .ZN(n15296) );
  INV_X1 U8817 ( .A(n7918), .ZN(n15316) );
  OAI211_X1 U8818 ( .C1(n7400), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n7393), .B(
        n7396), .ZN(n7918) );
  INV_X1 U8819 ( .A(n7394), .ZN(n7393) );
  AND2_X1 U8820 ( .A1(n15333), .A2(n15334), .ZN(n15336) );
  AND2_X1 U8821 ( .A1(n13393), .A2(n10327), .ZN(P3_U3897) );
  INV_X1 U8822 ( .A(n7363), .ZN(n7362) );
  OAI21_X1 U8823 ( .B1(n13323), .B2(n15128), .A(n12809), .ZN(n7363) );
  NAND2_X1 U8824 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  AOI211_X1 U8825 ( .C1(n15503), .C2(n13032), .A(n13021), .B(n13020), .ZN(
        n13022) );
  AOI21_X1 U8826 ( .B1(n13044), .B2(n15514), .A(n7495), .ZN(n13045) );
  NAND2_X1 U8827 ( .A1(n7359), .A2(n7355), .ZN(P2_U3233) );
  AOI21_X1 U8828 ( .B1(n15196), .B2(n15201), .A(n7356), .ZN(n7355) );
  NAND2_X1 U8829 ( .A1(n15195), .A2(n15205), .ZN(n7359) );
  NAND2_X1 U8830 ( .A1(n7361), .A2(n7357), .ZN(n7356) );
  INV_X1 U8831 ( .A(n8851), .ZN(n8852) );
  AOI21_X1 U8832 ( .B1(n14090), .B2(n14127), .A(n7580), .ZN(n7579) );
  AOI21_X1 U8833 ( .B1(n14104), .B2(n14127), .A(n7343), .ZN(n7794) );
  NAND2_X1 U8834 ( .A1(n7532), .A2(n7529), .ZN(P2_U3495) );
  INV_X1 U8835 ( .A(n7530), .ZN(n7529) );
  NAND2_X1 U8836 ( .A1(n14182), .A2(n14215), .ZN(n7532) );
  OAI21_X1 U8837 ( .B1(n14183), .B2(n14219), .A(n7531), .ZN(n7530) );
  NAND2_X1 U8838 ( .A1(n7396), .A2(n7395), .ZN(n15313) );
  XNOR2_X1 U8839 ( .A(n7916), .B(n7915), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8840 ( .A(n15365), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U8841 ( .A1(n15359), .A2(n7409), .ZN(n7916) );
  INV_X1 U8842 ( .A(n9641), .ZN(n9683) );
  AND2_X1 U8843 ( .A1(n10247), .A2(n10248), .ZN(n13185) );
  OR2_X1 U8844 ( .A1(n14609), .A2(n7213), .ZN(n7210) );
  AND2_X1 U8845 ( .A1(n14155), .A2(n14056), .ZN(n7211) );
  NAND2_X1 U8846 ( .A1(n9231), .A2(n9230), .ZN(n15953) );
  INV_X1 U8847 ( .A(n15953), .ZN(n7877) );
  AND2_X1 U8848 ( .A1(n10069), .A2(n8130), .ZN(n10067) );
  OR2_X2 U8849 ( .A1(n14713), .A2(n14714), .ZN(n7212) );
  AND2_X1 U8850 ( .A1(n14810), .A2(n12444), .ZN(n7213) );
  AND2_X1 U8851 ( .A1(n10260), .A2(n10266), .ZN(n13136) );
  AND2_X1 U8852 ( .A1(n7544), .A2(n7542), .ZN(n7214) );
  NOR2_X1 U8853 ( .A1(n12281), .A2(n12237), .ZN(n7215) );
  INV_X1 U8854 ( .A(n11876), .ZN(n11924) );
  AND3_X1 U8855 ( .A1(n9773), .A2(n9772), .A3(n9771), .ZN(n11876) );
  NAND2_X1 U8856 ( .A1(n7480), .A2(n7245), .ZN(n7216) );
  XNOR2_X1 U8857 ( .A(n14651), .B(n12673), .ZN(n14644) );
  INV_X1 U8858 ( .A(n14644), .ZN(n7960) );
  AND2_X1 U8859 ( .A1(n8106), .A2(n7326), .ZN(n7217) );
  NOR2_X1 U8860 ( .A1(n10250), .A2(n7671), .ZN(n7218) );
  AND2_X1 U8861 ( .A1(n9101), .A2(n8005), .ZN(n7219) );
  NAND2_X1 U8862 ( .A1(n14141), .A2(n14032), .ZN(n7220) );
  AND3_X1 U8863 ( .A1(n12766), .A2(n13158), .A3(n13138), .ZN(n7221) );
  OR2_X1 U8864 ( .A1(n14048), .A2(n14031), .ZN(n7222) );
  OR2_X1 U8865 ( .A1(n11945), .A2(n11944), .ZN(n7223) );
  NAND2_X1 U8866 ( .A1(n9418), .A2(n9417), .ZN(n14799) );
  INV_X1 U8867 ( .A(n14799), .ZN(n7554) );
  OR2_X1 U8868 ( .A1(n15888), .A2(n14361), .ZN(n7224) );
  AND2_X1 U8869 ( .A1(n10002), .A2(n10003), .ZN(n7225) );
  AND2_X1 U8870 ( .A1(n8234), .A2(n8235), .ZN(n7226) );
  NOR2_X1 U8871 ( .A1(n15850), .A2(n14362), .ZN(n7227) );
  INV_X1 U8872 ( .A(n9066), .ZN(n7994) );
  AND2_X1 U8873 ( .A1(n7641), .A2(n13215), .ZN(n7228) );
  INV_X1 U8874 ( .A(n12100), .ZN(n7982) );
  AND2_X1 U8875 ( .A1(n7748), .A2(n10095), .ZN(n7229) );
  XNOR2_X1 U8876 ( .A(n15310), .B(n15309), .ZN(n7230) );
  INV_X1 U8877 ( .A(n13704), .ZN(n8519) );
  OR2_X1 U8878 ( .A1(n9832), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7231) );
  AND2_X1 U8879 ( .A1(n10986), .A2(n13736), .ZN(n10708) );
  OR2_X1 U8880 ( .A1(n14721), .A2(n12454), .ZN(n7232) );
  OR2_X1 U8881 ( .A1(n11763), .A2(n11764), .ZN(n7233) );
  INV_X1 U8882 ( .A(n8323), .ZN(n8513) );
  OR2_X1 U8883 ( .A1(n11342), .A2(n13559), .ZN(n7234) );
  NOR2_X1 U8884 ( .A1(n8899), .A2(n8867), .ZN(n9486) );
  NAND2_X1 U8885 ( .A1(n9591), .A2(n9590), .ZN(n9595) );
  INV_X1 U8886 ( .A(n8861), .ZN(n8999) );
  AND2_X1 U8887 ( .A1(n7429), .A2(n11436), .ZN(n7235) );
  AND2_X1 U8888 ( .A1(n13236), .A2(n9873), .ZN(n7236) );
  NAND2_X1 U8889 ( .A1(n7964), .A2(n7962), .ZN(n14628) );
  AND4_X1 U8890 ( .A1(n8738), .A2(n8231), .A3(n8763), .A4(n8230), .ZN(n7237)
         );
  AND2_X1 U8891 ( .A1(n7935), .A2(n7452), .ZN(n7238) );
  OR2_X1 U8892 ( .A1(n12541), .A2(n12540), .ZN(n7239) );
  AND2_X1 U8893 ( .A1(n8817), .A2(n7220), .ZN(n7240) );
  AND2_X1 U8894 ( .A1(n7793), .A2(n8541), .ZN(n7241) );
  NAND2_X1 U8895 ( .A1(n9098), .A2(n9097), .ZN(n12119) );
  AND2_X1 U8896 ( .A1(n13018), .A2(n13017), .ZN(n7242) );
  NAND2_X1 U8897 ( .A1(n12726), .A2(n12722), .ZN(n8061) );
  AND2_X1 U8898 ( .A1(n8119), .A2(n9570), .ZN(n9717) );
  INV_X1 U8899 ( .A(n13971), .ZN(n7527) );
  NAND2_X1 U8900 ( .A1(n9498), .A2(n9497), .ZN(n10347) );
  NOR2_X1 U8901 ( .A1(n13580), .A2(n12488), .ZN(n7243) );
  AND3_X1 U8902 ( .A1(n8950), .A2(n8949), .A3(n8948), .ZN(n7244) );
  OR2_X1 U8903 ( .A1(n11849), .A2(n11842), .ZN(n7245) );
  NAND2_X1 U8904 ( .A1(n14293), .A2(n12622), .ZN(n15899) );
  OR2_X1 U8905 ( .A1(n14146), .A2(n14058), .ZN(n7246) );
  NAND2_X1 U8906 ( .A1(n8816), .A2(n8815), .ZN(n14068) );
  AND2_X1 U8907 ( .A1(n14168), .A2(n13800), .ZN(n7247) );
  AND2_X1 U8908 ( .A1(n13626), .A2(n13800), .ZN(n7248) );
  AND2_X1 U8909 ( .A1(n7603), .A2(n7246), .ZN(n7249) );
  NAND2_X1 U8910 ( .A1(n9822), .A2(n9821), .ZN(n12738) );
  INV_X1 U8911 ( .A(n12738), .ZN(n8116) );
  XNOR2_X1 U8912 ( .A(n8904), .B(n8903), .ZN(n8905) );
  NAND2_X1 U8913 ( .A1(n13685), .A2(n13684), .ZN(n14090) );
  INV_X1 U8914 ( .A(n14090), .ZN(n7382) );
  AND2_X1 U8915 ( .A1(n13559), .A2(n12507), .ZN(n7250) );
  INV_X1 U8916 ( .A(n11897), .ZN(n8111) );
  AND2_X1 U8917 ( .A1(n12819), .A2(n7760), .ZN(n7251) );
  INV_X1 U8918 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9584) );
  XNOR2_X1 U8919 ( .A(n8247), .B(n8246), .ZN(n8254) );
  AND2_X1 U8920 ( .A1(n12849), .A2(n12767), .ZN(n7252) );
  NAND2_X1 U8921 ( .A1(n8622), .A2(n8621), .ZN(n13994) );
  INV_X1 U8922 ( .A(n13994), .ZN(n14204) );
  NAND2_X1 U8923 ( .A1(n9316), .A2(n9315), .ZN(n14651) );
  AND2_X1 U8924 ( .A1(n14187), .A2(n14191), .ZN(n7253) );
  AND2_X1 U8925 ( .A1(n14817), .A2(n14358), .ZN(n7254) );
  OR2_X1 U8926 ( .A1(n14141), .A2(n13797), .ZN(n7255) );
  INV_X1 U8927 ( .A(n13602), .ZN(n7823) );
  OR2_X1 U8928 ( .A1(n15295), .A2(n15294), .ZN(n7256) );
  OR2_X1 U8929 ( .A1(n14155), .A2(n14056), .ZN(n7257) );
  AND4_X1 U8930 ( .A1(n7615), .A2(n8032), .A3(n8033), .A4(n7237), .ZN(n7258)
         );
  AND2_X1 U8931 ( .A1(n8237), .A2(n7226), .ZN(n7259) );
  NAND2_X1 U8932 ( .A1(n9078), .A2(n9077), .ZN(n15781) );
  NAND2_X1 U8933 ( .A1(n7964), .A2(n12462), .ZN(n14629) );
  OR2_X1 U8934 ( .A1(n15850), .A2(n12604), .ZN(n7260) );
  NAND2_X1 U8935 ( .A1(n9570), .A2(n9569), .ZN(n9688) );
  OR2_X1 U8936 ( .A1(n12606), .A2(n12604), .ZN(n7261) );
  AND2_X1 U8937 ( .A1(n8299), .A2(n8300), .ZN(n7262) );
  INV_X1 U8938 ( .A(n15260), .ZN(n7404) );
  AND2_X1 U8939 ( .A1(n7482), .A2(n13448), .ZN(n7263) );
  AND2_X1 U8940 ( .A1(n13339), .A2(n12907), .ZN(n7264) );
  AND2_X1 U8941 ( .A1(n10305), .A2(n9887), .ZN(n7265) );
  AND2_X1 U8942 ( .A1(n14048), .A2(n14031), .ZN(n7266) );
  INV_X1 U8943 ( .A(n13080), .ZN(n9985) );
  AND2_X1 U8944 ( .A1(n10158), .A2(n10156), .ZN(n13080) );
  INV_X1 U8945 ( .A(n15932), .ZN(n15920) );
  OR2_X1 U8946 ( .A1(n12045), .A2(n12044), .ZN(n7267) );
  OR2_X1 U8947 ( .A1(n13653), .A2(n13654), .ZN(n7268) );
  OR2_X1 U8948 ( .A1(n13661), .A2(n13662), .ZN(n7269) );
  NAND2_X1 U8949 ( .A1(n9251), .A2(n9250), .ZN(n15964) );
  NAND2_X1 U8950 ( .A1(n8031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U8951 ( .A1(n7942), .A2(n8685), .ZN(n8695) );
  AND2_X1 U8952 ( .A1(n7506), .A2(n7504), .ZN(n7270) );
  INV_X1 U8953 ( .A(n13579), .ZN(n7839) );
  INV_X1 U8954 ( .A(n7902), .ZN(n7901) );
  NAND2_X1 U8955 ( .A1(n12202), .A2(n7903), .ZN(n7902) );
  AND2_X1 U8956 ( .A1(n13600), .A2(n13805), .ZN(n7271) );
  NAND2_X1 U8957 ( .A1(n12769), .A2(n13128), .ZN(n7272) );
  AND2_X1 U8958 ( .A1(n9452), .A2(n12465), .ZN(n7273) );
  INV_X1 U8959 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7920) );
  XNOR2_X1 U8960 ( .A(n8784), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8772) );
  AND2_X1 U8961 ( .A1(n9872), .A2(n9857), .ZN(n7274) );
  AND2_X1 U8962 ( .A1(n12455), .A2(n7232), .ZN(n7275) );
  OR2_X1 U8963 ( .A1(n10002), .A2(n13077), .ZN(n10273) );
  INV_X1 U8964 ( .A(n15267), .ZN(n7909) );
  AND2_X1 U8965 ( .A1(n12687), .A2(n12686), .ZN(n7276) );
  NOR2_X1 U8966 ( .A1(n14638), .A2(n14358), .ZN(n12442) );
  INV_X1 U8967 ( .A(n13169), .ZN(n9940) );
  AND2_X1 U8968 ( .A1(n10249), .A2(n10056), .ZN(n13169) );
  NAND2_X1 U8969 ( .A1(n13222), .A2(n7265), .ZN(n13209) );
  INV_X1 U8970 ( .A(n8804), .ZN(n7626) );
  INV_X1 U8971 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8235) );
  NOR2_X1 U8972 ( .A1(n8867), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7277) );
  AND2_X1 U8973 ( .A1(n12534), .A2(n12533), .ZN(n7278) );
  AND2_X1 U8974 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7279) );
  NOR2_X1 U8975 ( .A1(n15742), .A2(n12044), .ZN(n7280) );
  NOR2_X1 U8976 ( .A1(n14195), .A2(n13664), .ZN(n7281) );
  OR2_X1 U8977 ( .A1(n13333), .A2(n13106), .ZN(n10152) );
  AND2_X1 U8978 ( .A1(n12616), .A2(n12615), .ZN(n7282) );
  OR2_X1 U8979 ( .A1(n15231), .A2(n7920), .ZN(n7283) );
  AND2_X1 U8980 ( .A1(n8202), .A2(n15053), .ZN(n7284) );
  INV_X1 U8981 ( .A(n9305), .ZN(n8013) );
  NAND2_X1 U8982 ( .A1(n12234), .A2(n14365), .ZN(n7285) );
  INV_X1 U8983 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U8984 ( .A1(n14104), .A2(n13790), .ZN(n7286) );
  AND2_X1 U8985 ( .A1(n11633), .A2(n15692), .ZN(n7287) );
  AND2_X1 U8986 ( .A1(n10717), .A2(n10716), .ZN(n7288) );
  AND2_X1 U8987 ( .A1(n11392), .A2(n11530), .ZN(n7289) );
  AND4_X1 U8988 ( .A1(n9576), .A2(n9575), .A3(n10022), .A4(n9574), .ZN(n7290)
         );
  NAND2_X1 U8989 ( .A1(n8222), .A2(n8221), .ZN(n7291) );
  NOR2_X1 U8990 ( .A1(n11938), .A2(n11932), .ZN(n7292) );
  AND2_X1 U8991 ( .A1(n12916), .A2(n11987), .ZN(n7293) );
  INV_X1 U8992 ( .A(n8597), .ZN(n7802) );
  NOR2_X1 U8993 ( .A1(n14804), .A2(n14356), .ZN(n7294) );
  NAND2_X1 U8994 ( .A1(n7941), .A2(n7940), .ZN(n7546) );
  INV_X1 U8995 ( .A(n12917), .ZN(n11978) );
  INV_X1 U8996 ( .A(n7977), .ZN(n7976) );
  NAND2_X1 U8997 ( .A1(n15878), .A2(n14258), .ZN(n7977) );
  OR2_X1 U8998 ( .A1(n7190), .A2(n13474), .ZN(n7295) );
  AND2_X1 U8999 ( .A1(n7554), .A2(n14586), .ZN(n7296) );
  AND2_X1 U9000 ( .A1(n7775), .A2(n7774), .ZN(n7297) );
  INV_X1 U9001 ( .A(n8061), .ZN(n8060) );
  OR2_X1 U9002 ( .A1(n10313), .A2(n8148), .ZN(n7298) );
  NAND2_X1 U9003 ( .A1(n7246), .A2(n8819), .ZN(n7299) );
  INV_X1 U9004 ( .A(n9207), .ZN(n7999) );
  INV_X1 U9005 ( .A(n7970), .ZN(n7969) );
  NAND2_X1 U9006 ( .A1(n7973), .A2(n7971), .ZN(n7970) );
  OR2_X1 U9007 ( .A1(n7554), .A2(n14586), .ZN(n7300) );
  NOR2_X1 U9008 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NAND2_X1 U9009 ( .A1(n10273), .A2(n10274), .ZN(n13068) );
  INV_X1 U9010 ( .A(n13563), .ZN(n7854) );
  OR2_X1 U9011 ( .A1(n13178), .A2(n13157), .ZN(n10249) );
  INV_X1 U9012 ( .A(n10249), .ZN(n7669) );
  AND2_X1 U9013 ( .A1(n7475), .A2(n7473), .ZN(n7301) );
  AND3_X1 U9014 ( .A1(n8263), .A2(n8261), .A3(n8262), .ZN(n7302) );
  INV_X1 U9015 ( .A(n13523), .ZN(n13529) );
  AND3_X1 U9016 ( .A1(n8279), .A2(n8277), .A3(n8278), .ZN(n7303) );
  NOR2_X1 U9017 ( .A1(n11679), .A2(n9737), .ZN(n7304) );
  AND2_X1 U9018 ( .A1(n9570), .A2(n8120), .ZN(n7305) );
  AND2_X1 U9019 ( .A1(n13920), .A2(n8824), .ZN(n7306) );
  OR2_X1 U9020 ( .A1(n14601), .A2(n7551), .ZN(n7307) );
  NAND2_X1 U9021 ( .A1(n10913), .A2(n11198), .ZN(n7308) );
  OR2_X1 U9022 ( .A1(n8010), .A2(n8008), .ZN(n7309) );
  AND2_X1 U9023 ( .A1(n7295), .A2(n8056), .ZN(n7310) );
  OR2_X1 U9024 ( .A1(n10319), .A2(n10318), .ZN(n7311) );
  AND2_X1 U9025 ( .A1(n8073), .A2(n12615), .ZN(n7312) );
  AND2_X1 U9026 ( .A1(n7951), .A2(n13726), .ZN(n7313) );
  NOR2_X1 U9027 ( .A1(n13100), .A2(n13103), .ZN(n7314) );
  AOI21_X1 U9028 ( .B1(n8073), .B2(n8075), .A(n8072), .ZN(n8071) );
  AND2_X1 U9029 ( .A1(n13117), .A2(n7647), .ZN(n7315) );
  OR2_X1 U9030 ( .A1(n13147), .A2(n13158), .ZN(n10260) );
  OR2_X1 U9031 ( .A1(n13638), .A2(n13636), .ZN(n7316) );
  OR2_X1 U9032 ( .A1(n7823), .A2(n13601), .ZN(n7317) );
  OR2_X1 U9033 ( .A1(n13590), .A2(n13588), .ZN(n7318) );
  AND2_X1 U9034 ( .A1(n7630), .A2(n7222), .ZN(n7319) );
  INV_X1 U9035 ( .A(n10002), .ZN(n13323) );
  NAND2_X1 U9036 ( .A1(n9996), .A2(n9995), .ZN(n10002) );
  AND2_X1 U9037 ( .A1(n8129), .A2(n9584), .ZN(n7320) );
  NAND2_X1 U9038 ( .A1(n10309), .A2(n7722), .ZN(n7321) );
  AND2_X1 U9039 ( .A1(n8088), .A2(n8862), .ZN(n7322) );
  NAND2_X1 U9040 ( .A1(n9067), .A2(n7994), .ZN(n7323) );
  INV_X1 U9041 ( .A(n8074), .ZN(n8073) );
  OAI21_X1 U9042 ( .B1(n14295), .B2(n8075), .A(n15897), .ZN(n8074) );
  INV_X1 U9043 ( .A(n8151), .ZN(n8125) );
  INV_X1 U9044 ( .A(n7767), .ZN(n7766) );
  NAND2_X1 U9045 ( .A1(n7768), .A2(n11980), .ZN(n7767) );
  AND2_X1 U9046 ( .A1(n7891), .A2(n7300), .ZN(n7889) );
  NAND2_X1 U9047 ( .A1(n9208), .A2(n7999), .ZN(n7324) );
  NAND2_X1 U9048 ( .A1(n9242), .A2(n7998), .ZN(n7325) );
  NAND2_X1 U9049 ( .A1(n12464), .A2(n7210), .ZN(n7893) );
  INV_X1 U9050 ( .A(n11039), .ZN(n11478) );
  NAND2_X1 U9051 ( .A1(n7533), .A2(n8603), .ZN(n14010) );
  INV_X1 U9052 ( .A(n14010), .ZN(n7586) );
  NAND2_X1 U9053 ( .A1(n8050), .A2(n8051), .ZN(n11933) );
  INV_X1 U9054 ( .A(n13431), .ZN(n8055) );
  NAND2_X1 U9055 ( .A1(n8488), .A2(n8487), .ZN(n15862) );
  INV_X1 U9056 ( .A(n15862), .ZN(n7575) );
  NAND2_X1 U9057 ( .A1(n7593), .A2(n7592), .ZN(n12371) );
  NAND2_X1 U9058 ( .A1(n7594), .A2(n8814), .ZN(n12390) );
  NAND2_X1 U9059 ( .A1(n8109), .A2(n8112), .ZN(n11896) );
  NAND2_X1 U9060 ( .A1(n12915), .A2(n10052), .ZN(n7326) );
  INV_X1 U9061 ( .A(n10201), .ZN(n7664) );
  AND2_X1 U9062 ( .A1(n8070), .A2(n8068), .ZN(n7327) );
  INV_X1 U9063 ( .A(n13615), .ZN(n7845) );
  INV_X1 U9064 ( .A(n15902), .ZN(n7876) );
  OR2_X1 U9065 ( .A1(n15405), .A2(n12931), .ZN(n7328) );
  AND2_X1 U9066 ( .A1(n12754), .A2(n13198), .ZN(n7329) );
  NAND2_X1 U9067 ( .A1(n15918), .A2(n7564), .ZN(n7565) );
  NOR2_X1 U9068 ( .A1(n8030), .A2(n9353), .ZN(n8026) );
  OR2_X1 U9069 ( .A1(n8564), .A2(SI_19_), .ZN(n7330) );
  INV_X1 U9070 ( .A(n13658), .ZN(n7850) );
  INV_X1 U9071 ( .A(n7463), .ZN(n12342) );
  NAND2_X1 U9072 ( .A1(n12493), .A2(n7461), .ZN(n7463) );
  AND2_X1 U9073 ( .A1(n8030), .A2(n9353), .ZN(n8029) );
  INV_X1 U9074 ( .A(n8029), .ZN(n8028) );
  INV_X1 U9075 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9579) );
  OR2_X1 U9076 ( .A1(n13485), .A2(n13976), .ZN(n7331) );
  NOR2_X1 U9077 ( .A1(n12143), .A2(n12135), .ZN(n7332) );
  AND2_X1 U9078 ( .A1(n12743), .A2(n12898), .ZN(n7333) );
  AND2_X1 U9079 ( .A1(n11909), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U9080 ( .A1(n12951), .A2(n15405), .ZN(n7335) );
  AND2_X1 U9081 ( .A1(n8218), .A2(n15044), .ZN(n7336) );
  AND2_X1 U9082 ( .A1(n9547), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7337) );
  INV_X1 U9083 ( .A(n9278), .ZN(n8019) );
  INV_X1 U9084 ( .A(n9241), .ZN(n7998) );
  INV_X1 U9085 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9483) );
  INV_X1 U9086 ( .A(n9171), .ZN(n7995) );
  AND2_X1 U9087 ( .A1(n7515), .A2(n7518), .ZN(n7338) );
  INV_X1 U9088 ( .A(n15427), .ZN(n7518) );
  AND2_X1 U9089 ( .A1(n7400), .A2(n7399), .ZN(n7339) );
  OR2_X1 U9090 ( .A1(n13625), .A2(n13623), .ZN(n7340) );
  AND2_X1 U9091 ( .A1(n7848), .A2(n13662), .ZN(n7341) );
  NAND2_X1 U9092 ( .A1(n9172), .A2(n7995), .ZN(n7342) );
  INV_X1 U9093 ( .A(n7193), .ZN(n8832) );
  NAND2_X1 U9094 ( .A1(n9112), .A2(n9111), .ZN(n12234) );
  INV_X1 U9095 ( .A(n12234), .ZN(n7560) );
  NAND2_X1 U9096 ( .A1(n8588), .A2(n8587), .ZN(n14141) );
  INV_X1 U9097 ( .A(n14141), .ZN(n7587) );
  NAND2_X1 U9098 ( .A1(n13508), .A2(n11280), .ZN(n11288) );
  AND2_X1 U9099 ( .A1(n7751), .A2(n11181), .ZN(n7753) );
  AND2_X1 U9100 ( .A1(n15868), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7343) );
  OR2_X1 U9101 ( .A1(n15652), .A2(n15658), .ZN(n11774) );
  OAI21_X1 U9102 ( .B1(n11337), .B2(n7591), .A(n7589), .ZN(n11100) );
  AND2_X1 U9103 ( .A1(n7428), .A2(n7426), .ZN(n11631) );
  NAND2_X1 U9104 ( .A1(n8797), .A2(n8796), .ZN(n11418) );
  NAND2_X1 U9105 ( .A1(n11337), .A2(n8791), .ZN(n11137) );
  NAND2_X1 U9106 ( .A1(n11774), .A2(n11717), .ZN(n11776) );
  INV_X1 U9107 ( .A(SI_16_), .ZN(n15047) );
  AND2_X1 U9108 ( .A1(n7510), .A2(n7512), .ZN(n7344) );
  AND2_X1 U9109 ( .A1(n11182), .A2(n7753), .ZN(n7345) );
  AND2_X1 U9110 ( .A1(n7430), .A2(n7235), .ZN(n7346) );
  AND2_X1 U9111 ( .A1(n8653), .A2(SI_24_), .ZN(n7347) );
  AND2_X1 U9112 ( .A1(n11907), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7348) );
  AND2_X1 U9113 ( .A1(n8696), .A2(n8685), .ZN(n7349) );
  AND2_X1 U9114 ( .A1(n7517), .A2(n7515), .ZN(n7350) );
  NAND2_X1 U9115 ( .A1(n8860), .A2(n8861), .ZN(n9228) );
  INV_X1 U9116 ( .A(n11705), .ZN(n7886) );
  AND2_X1 U9117 ( .A1(n7738), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U9118 ( .A1(n8037), .A2(n13776), .ZN(n10707) );
  NAND2_X1 U9119 ( .A1(n8474), .A2(n8473), .ZN(n13612) );
  INV_X1 U9120 ( .A(n13612), .ZN(n7577) );
  OR2_X1 U9121 ( .A1(n12033), .A2(n11973), .ZN(n7352) );
  NAND2_X1 U9122 ( .A1(n15596), .A2(n11513), .ZN(n11512) );
  INV_X1 U9123 ( .A(n11512), .ZN(n7556) );
  NAND2_X1 U9124 ( .A1(n11176), .A2(n10165), .ZN(n10285) );
  INV_X1 U9125 ( .A(n10412), .ZN(n7907) );
  INV_X1 U9126 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7490) );
  INV_X1 U9127 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7412) );
  INV_X1 U9128 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7385) );
  INV_X1 U9129 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15226) );
  INV_X1 U9130 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7707) );
  INV_X1 U9131 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7737) );
  INV_X1 U9132 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7398) );
  AND3_X1 U9133 ( .A1(n10347), .A2(P1_STATE_REG_SCAN_IN), .A3(n10623), .ZN(
        n10634) );
  CLKBUF_X3 U9134 ( .A(n13553), .Z(n13708) );
  NAND2_X1 U9135 ( .A1(n7859), .A2(n7857), .ZN(n7950) );
  INV_X1 U9136 ( .A(n7353), .ZN(n13585) );
  NOR2_X1 U9137 ( .A1(n13583), .A2(n13584), .ZN(n7353) );
  INV_X1 U9138 ( .A(n7354), .ZN(n13620) );
  NOR2_X1 U9139 ( .A1(n13618), .A2(n13619), .ZN(n7354) );
  AOI21_X1 U9140 ( .B1(n7855), .B2(n7856), .A(n7854), .ZN(n7852) );
  NAND2_X2 U9141 ( .A1(n10057), .A2(n10253), .ZN(n13150) );
  NAND2_X1 U9142 ( .A1(n10046), .A2(n10173), .ZN(n11540) );
  NAND2_X1 U9143 ( .A1(n12166), .A2(n10217), .ZN(n12268) );
  NAND2_X1 U9144 ( .A1(n10051), .A2(n7666), .ZN(n7665) );
  NAND2_X1 U9145 ( .A1(n7739), .A2(n7290), .ZN(n8142) );
  NOR2_X2 U9146 ( .A1(n9582), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U9147 ( .A1(n10069), .A2(n7320), .ZN(n9582) );
  NAND2_X1 U9148 ( .A1(n11974), .A2(n11975), .ZN(n15167) );
  NAND2_X1 U9149 ( .A1(n15161), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n15160) );
  AOI21_X1 U9150 ( .B1(n13865), .B2(n11081), .A(n11082), .ZN(n11374) );
  NOR2_X1 U9151 ( .A1(n11378), .A2(n11377), .ZN(n11967) );
  INV_X1 U9152 ( .A(n11970), .ZN(n7360) );
  NAND2_X1 U9153 ( .A1(n15208), .A2(n15207), .ZN(n15206) );
  AOI21_X1 U9154 ( .B1(n10646), .B2(P2_REG2_REG_4__SCAN_IN), .A(n10638), .ZN(
        n10663) );
  NOR2_X1 U9155 ( .A1(n15191), .A2(n15190), .ZN(n15193) );
  AOI21_X1 U9156 ( .B1(n10752), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10746), .ZN(
        n13853) );
  AOI21_X1 U9157 ( .B1(n10683), .B2(P2_REG2_REG_7__SCAN_IN), .A(n10677), .ZN(
        n10680) );
  AOI21_X1 U9158 ( .B1(n11078), .B2(P2_REG2_REG_10__SCAN_IN), .A(n11077), .ZN(
        n13867) );
  AOI21_X1 U9159 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10648), .A(n15148), .ZN(
        n10644) );
  NOR2_X2 U9160 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8294) );
  NAND2_X1 U9161 ( .A1(n13394), .A2(n10762), .ZN(n10763) );
  NAND2_X1 U9162 ( .A1(n7364), .A2(n7362), .ZN(P3_U3160) );
  NAND2_X1 U9163 ( .A1(n12805), .A2(n15131), .ZN(n7364) );
  NAND2_X1 U9164 ( .A1(n7743), .A2(n7742), .ZN(n12792) );
  NAND2_X1 U9165 ( .A1(n12757), .A2(n12756), .ZN(n12861) );
  INV_X1 U9166 ( .A(n11885), .ZN(n11883) );
  AOI22_X2 U9167 ( .A1(n14655), .A2(n12441), .B1(n12667), .B2(n14670), .ZN(
        n14642) );
  NAND2_X2 U9168 ( .A1(n14626), .A2(n14630), .ZN(n14625) );
  NOR2_X2 U9169 ( .A1(n12414), .A2(n12413), .ZN(n15875) );
  NAND2_X1 U9170 ( .A1(n14743), .A2(n14742), .ZN(n14741) );
  NAND2_X1 U9171 ( .A1(n7880), .A2(n7881), .ZN(n15769) );
  NAND2_X1 U9172 ( .A1(n7366), .A2(n7321), .ZN(n10283) );
  NAND3_X1 U9173 ( .A1(n7720), .A2(n7721), .A3(n7719), .ZN(n7366) );
  NAND2_X1 U9174 ( .A1(n7370), .A2(n7367), .ZN(n10271) );
  NOR2_X1 U9175 ( .A1(n10264), .A2(n10261), .ZN(n7369) );
  NAND3_X1 U9176 ( .A1(n10306), .A2(n10267), .A3(n10260), .ZN(n7370) );
  NAND2_X1 U9177 ( .A1(n9555), .A2(n9554), .ZN(n9876) );
  NAND2_X1 U9178 ( .A1(n9618), .A2(n9617), .ZN(n9621) );
  NAND2_X1 U9179 ( .A1(n9918), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U9180 ( .A1(n7733), .A2(n7351), .ZN(n7732) );
  OAI21_X1 U9181 ( .B1(n9550), .B2(n7706), .A(n9551), .ZN(n7702) );
  OAI21_X1 U9182 ( .B1(n9929), .B2(n9927), .A(n9564), .ZN(n9943) );
  NAND3_X1 U9183 ( .A1(n7687), .A2(n7311), .A3(n7638), .ZN(n7637) );
  NOR3_X2 U9184 ( .A1(n10291), .A2(n10290), .A3(n10313), .ZN(n10316) );
  OR2_X2 U9185 ( .A1(n13154), .A2(n10257), .ZN(n10057) );
  NAND2_X4 U9186 ( .A1(n10032), .A2(n12134), .ZN(n10805) );
  NAND2_X2 U9187 ( .A1(n13074), .A2(n13080), .ZN(n13076) );
  NAND2_X1 U9188 ( .A1(n12750), .A2(n7744), .ZN(n7743) );
  NAND2_X1 U9189 ( .A1(n9958), .A2(n9957), .ZN(n9973) );
  NAND2_X1 U9190 ( .A1(n9562), .A2(n9561), .ZN(n9929) );
  NAND2_X1 U9191 ( .A1(n9943), .A2(n9942), .ZN(n9945) );
  NAND2_X1 U9192 ( .A1(n9818), .A2(n7704), .ZN(n7703) );
  NAND2_X1 U9193 ( .A1(n10271), .A2(n10286), .ZN(n7720) );
  NAND2_X1 U9194 ( .A1(n7712), .A2(n7716), .ZN(n9538) );
  NOR2_X2 U9195 ( .A1(n10264), .A2(n13124), .ZN(n10306) );
  NAND3_X1 U9196 ( .A1(n13089), .A2(n13080), .A3(n13103), .ZN(n10264) );
  NOR3_X2 U9197 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_15__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U9198 ( .A1(n11518), .A2(n11508), .ZN(n11507) );
  INV_X2 U9199 ( .A(n9370), .ZN(n9408) );
  NAND2_X1 U9200 ( .A1(n14807), .A2(n14808), .ZN(n14864) );
  AOI21_X2 U9201 ( .B1(n14597), .B2(n15914), .A(n14596), .ZN(n14807) );
  NAND2_X1 U9202 ( .A1(n14711), .A2(n12437), .ZN(n14696) );
  NAND2_X1 U9203 ( .A1(n8332), .A2(n8178), .ZN(n8351) );
  NAND2_X1 U9204 ( .A1(n15454), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15453) );
  XNOR2_X1 U9205 ( .A(n12983), .B(n15450), .ZN(n15454) );
  NOR2_X1 U9206 ( .A1(n13018), .A2(n13017), .ZN(n13028) );
  NAND3_X1 U9207 ( .A1(n9194), .A2(n9193), .A3(n7324), .ZN(n7374) );
  NAND3_X1 U9208 ( .A1(n9227), .A2(n9226), .A3(n7325), .ZN(n7376) );
  NAND3_X1 U9209 ( .A1(n9157), .A2(n9156), .A3(n7342), .ZN(n7378) );
  NAND3_X1 U9210 ( .A1(n9050), .A2(n9049), .A3(n7323), .ZN(n7380) );
  OAI21_X1 U9211 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8987) );
  AOI21_X1 U9212 ( .B1(n8968), .B2(n8967), .A(n11366), .ZN(n8969) );
  NAND2_X1 U9213 ( .A1(n8265), .A2(n8165), .ZN(n8290) );
  OR2_X2 U9214 ( .A1(n11467), .A2(n13587), .ZN(n11619) );
  AND2_X2 U9215 ( .A1(n13978), .A2(n14195), .ZN(n13962) );
  NAND2_X1 U9216 ( .A1(n8299), .A2(n7383), .ZN(n8292) );
  OR2_X1 U9217 ( .A1(n8290), .A2(SI_2_), .ZN(n7383) );
  NAND2_X1 U9218 ( .A1(n8290), .A2(SI_2_), .ZN(n8299) );
  NAND2_X1 U9219 ( .A1(n7890), .A2(n7210), .ZN(n14594) );
  NAND2_X1 U9220 ( .A1(n11241), .A2(n11240), .ZN(n11700) );
  OAI21_X2 U9221 ( .B1(n12203), .B2(n7897), .A(n7895), .ZN(n12414) );
  AOI211_X2 U9222 ( .C1(n13094), .C2(n15577), .A(n13093), .B(n13092), .ZN(
        n13331) );
  NAND2_X1 U9223 ( .A1(n10069), .A2(n8129), .ZN(n7502) );
  XNOR2_X1 U9224 ( .A(n11189), .B(n12922), .ZN(n7634) );
  OAI21_X1 U9225 ( .B1(n15368), .B2(n15367), .A(P2_ADDR_REG_6__SCAN_IN), .ZN(
        n7391) );
  OAI21_X1 U9226 ( .B1(n7399), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7395), .ZN(
        n7394) );
  NAND2_X1 U9227 ( .A1(n15268), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U9228 ( .A1(n7403), .A2(n7406), .ZN(n7402) );
  NAND2_X1 U9229 ( .A1(n7406), .A2(n15260), .ZN(n15266) );
  NAND2_X1 U9230 ( .A1(n7404), .A2(n7909), .ZN(n7405) );
  NAND2_X1 U9231 ( .A1(n15347), .A2(n15348), .ZN(n15354) );
  NAND2_X1 U9232 ( .A1(n15358), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U9233 ( .A1(n15336), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n15337) );
  AOI21_X1 U9234 ( .B1(n15331), .B2(n15330), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n7410) );
  NOR2_X1 U9235 ( .A1(n15331), .A2(n15330), .ZN(n15332) );
  AND2_X1 U9236 ( .A1(n7415), .A2(n7414), .ZN(n10627) );
  NAND2_X1 U9237 ( .A1(n10355), .A2(n10913), .ZN(n7414) );
  NAND2_X4 U9238 ( .A1(n10994), .A2(n14763), .ZN(n12706) );
  INV_X1 U9239 ( .A(n12614), .ZN(n12612) );
  INV_X1 U9240 ( .A(n11597), .ZN(n7426) );
  INV_X1 U9241 ( .A(n7430), .ZN(n11434) );
  INV_X1 U9242 ( .A(n11436), .ZN(n7427) );
  INV_X1 U9243 ( .A(n11433), .ZN(n7429) );
  NAND2_X1 U9244 ( .A1(n14330), .A2(n7434), .ZN(n7432) );
  NAND2_X1 U9245 ( .A1(n14330), .A2(n14331), .ZN(n7433) );
  NAND2_X1 U9246 ( .A1(n8894), .A2(n8893), .ZN(n7442) );
  NAND2_X1 U9247 ( .A1(n8894), .A2(n7439), .ZN(n7438) );
  NAND2_X1 U9248 ( .A1(n8067), .A2(n7312), .ZN(n7447) );
  NAND2_X1 U9249 ( .A1(n7445), .A2(n8073), .ZN(n7446) );
  INV_X1 U9250 ( .A(n12616), .ZN(n7445) );
  NAND3_X1 U9251 ( .A1(n7447), .A2(n7446), .A3(n8071), .ZN(n15946) );
  NAND4_X1 U9252 ( .A1(n8861), .A2(n9182), .A3(n7322), .A4(n8859), .ZN(n8901)
         );
  NAND4_X1 U9253 ( .A1(n9181), .A2(n8859), .A3(n8861), .A4(n8088), .ZN(n8899)
         );
  NAND2_X1 U9254 ( .A1(n8353), .A2(n8182), .ZN(n8367) );
  NAND2_X1 U9255 ( .A1(n8353), .A2(n7238), .ZN(n7451) );
  OAI21_X1 U9256 ( .B1(n8353), .B2(n7938), .A(n7238), .ZN(n8397) );
  NAND2_X1 U9257 ( .A1(n12493), .A2(n7454), .ZN(n7457) );
  AOI21_X2 U9258 ( .B1(n8038), .B2(n12359), .A(n7456), .ZN(n12535) );
  NAND2_X1 U9259 ( .A1(n13417), .A2(n12547), .ZN(n7465) );
  OAI211_X1 U9260 ( .C1(n12559), .C2(n7474), .A(n7470), .B(n7469), .ZN(n12737)
         );
  NAND2_X1 U9261 ( .A1(n12559), .A2(n7301), .ZN(n7469) );
  OAI21_X1 U9262 ( .B1(n7475), .B2(n12731), .A(n7471), .ZN(n7470) );
  INV_X1 U9263 ( .A(n12731), .ZN(n7473) );
  NAND2_X1 U9264 ( .A1(n12524), .A2(n11840), .ZN(n7480) );
  NAND2_X1 U9265 ( .A1(n13496), .A2(n7310), .ZN(n7481) );
  NAND2_X1 U9266 ( .A1(n7488), .A2(n10817), .ZN(n10864) );
  INV_X1 U9267 ( .A(n10863), .ZN(n7489) );
  MUX2_X1 U9268 ( .A(n10809), .B(P3_REG2_REG_2__SCAN_IN), .S(n10892), .Z(
        n10882) );
  XNOR2_X2 U9269 ( .A(n7494), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10892) );
  INV_X1 U9270 ( .A(n9570), .ZN(n9676) );
  NAND3_X2 U9271 ( .A1(n9570), .A2(n8119), .A3(n9573), .ZN(n9811) );
  OAI22_X1 U9272 ( .A1(n15507), .A2(n7503), .B1(n7504), .B2(n13005), .ZN(
        n13031) );
  INV_X1 U9273 ( .A(n15507), .ZN(n7507) );
  NAND2_X1 U9274 ( .A1(n15385), .A2(n7338), .ZN(n7509) );
  NAND2_X1 U9275 ( .A1(n7509), .A2(n7511), .ZN(n15426) );
  NAND2_X1 U9276 ( .A1(n13970), .A2(n7525), .ZN(n7522) );
  NAND2_X1 U9277 ( .A1(n7522), .A2(n7523), .ZN(n13931) );
  NAND3_X1 U9278 ( .A1(n14103), .A2(n14101), .A3(n14102), .ZN(n14182) );
  NAND2_X1 U9279 ( .A1(n8414), .A2(n8413), .ZN(n8416) );
  NAND2_X1 U9280 ( .A1(n8214), .A2(n15047), .ZN(n7941) );
  OR2_X1 U9281 ( .A1(n8214), .A2(n15047), .ZN(n8215) );
  AND4_X2 U9282 ( .A1(n8079), .A2(n8080), .A3(n8078), .A4(n8853), .ZN(n8980)
         );
  NOR2_X2 U9283 ( .A1(n14686), .A2(n14670), .ZN(n7547) );
  NOR2_X1 U9284 ( .A1(n14601), .A2(n14799), .ZN(n14576) );
  AND2_X2 U9285 ( .A1(n7555), .A2(n8143), .ZN(n15620) );
  AND2_X1 U9286 ( .A1(n8918), .A2(n8917), .ZN(n7555) );
  NAND3_X1 U9287 ( .A1(n7562), .A2(n14737), .A3(n15918), .ZN(n14715) );
  NAND3_X1 U9288 ( .A1(n14737), .A2(n15918), .A3(n7564), .ZN(n14732) );
  INV_X1 U9289 ( .A(n7565), .ZN(n14752) );
  AND2_X2 U9290 ( .A1(n7569), .A2(n7568), .ZN(n8033) );
  NAND2_X2 U9291 ( .A1(n7573), .A2(n7570), .ZN(n14231) );
  NOR2_X2 U9292 ( .A1(n12191), .A2(n13622), .ZN(n12386) );
  NAND2_X1 U9293 ( .A1(n7582), .A2(n7579), .ZN(P2_U3530) );
  NOR2_X1 U9294 ( .A1(n15869), .A2(n7581), .ZN(n7580) );
  NAND2_X1 U9295 ( .A1(n14173), .A2(n15869), .ZN(n7582) );
  AND2_X2 U9296 ( .A1(n13962), .A2(n7583), .ZN(n13889) );
  NAND2_X1 U9297 ( .A1(n12185), .A2(n7595), .ZN(n7593) );
  XNOR2_X2 U9298 ( .A(n10709), .B(n13522), .ZN(n13745) );
  NAND2_X1 U9299 ( .A1(n7258), .A2(n7613), .ZN(n8244) );
  NOR2_X2 U9300 ( .A1(n7614), .A2(n7617), .ZN(n8237) );
  NAND3_X1 U9301 ( .A1(n7616), .A2(n7237), .A3(n8032), .ZN(n7614) );
  NAND3_X1 U9302 ( .A1(n7616), .A2(n8032), .A3(n8036), .ZN(n8238) );
  NAND2_X1 U9303 ( .A1(n13935), .A2(n7306), .ZN(n13910) );
  NAND2_X1 U9304 ( .A1(n13972), .A2(n8822), .ZN(n7618) );
  NAND2_X1 U9305 ( .A1(n7618), .A2(n7619), .ZN(n8823) );
  NAND2_X1 U9306 ( .A1(n11615), .A2(n7625), .ZN(n7622) );
  NAND2_X1 U9307 ( .A1(n8816), .A2(n7319), .ZN(n7628) );
  NAND2_X1 U9308 ( .A1(n7628), .A2(n7629), .ZN(n14029) );
  NAND2_X1 U9309 ( .A1(n11805), .A2(n7631), .ZN(n12003) );
  NAND2_X1 U9310 ( .A1(n7632), .A2(n10177), .ZN(n11678) );
  NAND2_X1 U9311 ( .A1(n11540), .A2(n10175), .ZN(n7632) );
  OAI211_X1 U9312 ( .C1(n11540), .C2(n7635), .A(n11679), .B(n7633), .ZN(n10047) );
  NAND2_X1 U9313 ( .A1(n7634), .A2(n10177), .ZN(n7633) );
  INV_X1 U9314 ( .A(n10177), .ZN(n7635) );
  NAND2_X1 U9315 ( .A1(n7636), .A2(n10323), .ZN(P3_U3296) );
  NAND2_X1 U9316 ( .A1(n7637), .A2(n10320), .ZN(n7636) );
  NAND2_X1 U9317 ( .A1(n7688), .A2(n10151), .ZN(n7638) );
  XNOR2_X2 U9318 ( .A(n15546), .B(n15580), .ZN(n15572) );
  AND2_X2 U9319 ( .A1(n10805), .A2(n10398), .ZN(n9664) );
  OAI21_X1 U9320 ( .B1(n13244), .B2(n13223), .A(n7643), .ZN(n13216) );
  NAND2_X1 U9321 ( .A1(n7642), .A2(n7228), .ZN(n13214) );
  NAND2_X1 U9322 ( .A1(n13244), .A2(n7643), .ZN(n7642) );
  NAND2_X1 U9323 ( .A1(n13150), .A2(n10260), .ZN(n7646) );
  NAND2_X1 U9324 ( .A1(n7649), .A2(n7650), .ZN(n13074) );
  NAND2_X1 U9325 ( .A1(n13110), .A2(n7652), .ZN(n7649) );
  NAND2_X1 U9326 ( .A1(n13110), .A2(n10155), .ZN(n7651) );
  NAND2_X1 U9327 ( .A1(n11996), .A2(n7657), .ZN(n7656) );
  NAND2_X1 U9328 ( .A1(n7665), .A2(n7663), .ZN(n11895) );
  NAND2_X1 U9329 ( .A1(n10051), .A2(n10195), .ZN(n11857) );
  NOR2_X1 U9330 ( .A1(n10199), .A2(n7667), .ZN(n7666) );
  INV_X1 U9331 ( .A(n10195), .ZN(n7667) );
  NAND2_X1 U9332 ( .A1(n13183), .A2(n7218), .ZN(n7670) );
  INV_X1 U9333 ( .A(n13185), .ZN(n7672) );
  NAND2_X1 U9334 ( .A1(n13076), .A2(n7684), .ZN(n7678) );
  NAND2_X1 U9335 ( .A1(n13076), .A2(n10158), .ZN(n13069) );
  XNOR2_X1 U9336 ( .A(n10149), .B(n7209), .ZN(n7688) );
  NAND2_X1 U9337 ( .A1(n7695), .A2(n7696), .ZN(n9905) );
  NAND2_X1 U9338 ( .A1(n7703), .A2(n7701), .ZN(n9846) );
  NAND2_X1 U9339 ( .A1(n7705), .A2(n9550), .ZN(n9831) );
  INV_X1 U9340 ( .A(n9830), .ZN(n7706) );
  NAND2_X1 U9341 ( .A1(n9662), .A2(n9524), .ZN(n7709) );
  NAND2_X1 U9342 ( .A1(n9523), .A2(n7708), .ZN(n7710) );
  NAND3_X1 U9343 ( .A1(n7710), .A2(n9672), .A3(n7709), .ZN(n9527) );
  NAND2_X1 U9344 ( .A1(n7711), .A2(n9524), .ZN(n9674) );
  NAND2_X1 U9345 ( .A1(n9663), .A2(n9661), .ZN(n7711) );
  NAND2_X1 U9346 ( .A1(n9534), .A2(n7713), .ZN(n7712) );
  INV_X1 U9347 ( .A(n10283), .ZN(n10289) );
  NAND2_X1 U9348 ( .A1(n9621), .A2(n7726), .ZN(n7725) );
  NAND2_X1 U9349 ( .A1(n9621), .A2(n9620), .ZN(n9958) );
  INV_X1 U9350 ( .A(n9613), .ZN(n7733) );
  NAND3_X1 U9351 ( .A1(n7732), .A2(n7734), .A3(n7729), .ZN(n9616) );
  NAND3_X1 U9352 ( .A1(n7732), .A2(n7730), .A3(n7729), .ZN(n9618) );
  NAND4_X1 U9353 ( .A1(n7741), .A2(n7740), .A3(n9577), .A4(n9833), .ZN(n10020)
         );
  NAND2_X1 U9354 ( .A1(n7748), .A2(n7747), .ZN(n10078) );
  AOI21_X1 U9355 ( .B1(n7753), .B2(n7752), .A(n7289), .ZN(n7749) );
  INV_X1 U9356 ( .A(n7753), .ZN(n7750) );
  INV_X1 U9357 ( .A(n11184), .ZN(n7751) );
  NAND2_X1 U9358 ( .A1(n12765), .A2(n7755), .ZN(n7754) );
  OAI21_X1 U9359 ( .B1(n11883), .B2(n7767), .A(n7765), .ZN(n12141) );
  OAI21_X2 U9360 ( .B1(n12352), .B2(n7771), .A(n7769), .ZN(n12826) );
  AND2_X1 U9361 ( .A1(n10069), .A2(n9578), .ZN(n10066) );
  NAND2_X1 U9362 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  NAND2_X1 U9363 ( .A1(n9531), .A2(n9530), .ZN(n9720) );
  XNOR2_X1 U9364 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9649) );
  NAND2_X1 U9365 ( .A1(n9553), .A2(n9552), .ZN(n9860) );
  AND2_X1 U9366 ( .A1(n11038), .A2(n11037), .ZN(n11041) );
  AND3_X4 U9367 ( .A1(n8274), .A2(n8273), .A3(n8272), .ZN(n13522) );
  OR2_X2 U9368 ( .A1(n11325), .A2(n13540), .ZN(n11327) );
  AND2_X2 U9369 ( .A1(n11453), .A2(n12487), .ZN(n11454) );
  OR2_X2 U9370 ( .A1(n12389), .A2(n13635), .ZN(n14077) );
  NAND2_X1 U9371 ( .A1(n9860), .A2(n9858), .ZN(n9555) );
  NAND2_X1 U9372 ( .A1(n9846), .A2(n9845), .ZN(n9553) );
  OAI21_X1 U9373 ( .B1(n13750), .B2(n7782), .A(n13751), .ZN(n7778) );
  NAND2_X1 U9374 ( .A1(n7779), .A2(n7777), .ZN(n11135) );
  INV_X1 U9375 ( .A(n7778), .ZN(n7777) );
  NAND2_X1 U9376 ( .A1(n11002), .A2(n7780), .ZN(n7779) );
  NAND2_X1 U9377 ( .A1(n11612), .A2(n7787), .ZN(n7784) );
  NAND2_X1 U9378 ( .A1(n7784), .A2(n7785), .ZN(n11804) );
  NAND2_X1 U9379 ( .A1(n7795), .A2(n7794), .ZN(P2_U3527) );
  NAND2_X1 U9380 ( .A1(n14182), .A2(n15869), .ZN(n7795) );
  NAND2_X1 U9381 ( .A1(n8237), .A2(n7796), .ZN(n8250) );
  NAND2_X1 U9382 ( .A1(n8581), .A2(n7800), .ZN(n7797) );
  NAND2_X1 U9383 ( .A1(n7797), .A2(n7798), .ZN(n13988) );
  OR2_X1 U9384 ( .A1(n13931), .A2(n13930), .ZN(n7814) );
  NAND2_X1 U9385 ( .A1(n7804), .A2(n7805), .ZN(n8728) );
  NAND2_X1 U9386 ( .A1(n12182), .A2(n7817), .ZN(n7816) );
  NAND3_X1 U9387 ( .A1(n13541), .A2(n13539), .A3(n13538), .ZN(n7820) );
  NAND3_X1 U9388 ( .A1(n7820), .A2(n7819), .A3(n7818), .ZN(n13547) );
  NAND3_X1 U9389 ( .A1(n13539), .A2(n13538), .A3(n13543), .ZN(n7818) );
  NAND2_X1 U9390 ( .A1(n7821), .A2(n7822), .ZN(n13606) );
  NAND3_X1 U9391 ( .A1(n13599), .A2(n7317), .A3(n13598), .ZN(n7821) );
  NAND2_X1 U9392 ( .A1(n7824), .A2(n7825), .ZN(n13641) );
  NAND3_X1 U9393 ( .A1(n13634), .A2(n7316), .A3(n13633), .ZN(n7824) );
  NAND2_X1 U9394 ( .A1(n7826), .A2(n7827), .ZN(n13594) );
  NAND3_X1 U9395 ( .A1(n13586), .A2(n7318), .A3(n13585), .ZN(n7826) );
  NAND2_X1 U9396 ( .A1(n7828), .A2(n7829), .ZN(n13629) );
  NAND3_X1 U9397 ( .A1(n13621), .A2(n7340), .A3(n13620), .ZN(n7828) );
  OAI21_X1 U9398 ( .B1(n13648), .B2(n7834), .A(n7833), .ZN(n13653) );
  NAND2_X1 U9399 ( .A1(n7830), .A2(n7831), .ZN(n13652) );
  NAND2_X1 U9400 ( .A1(n13648), .A2(n7833), .ZN(n7830) );
  OAI21_X1 U9401 ( .B1(n13578), .B2(n7840), .A(n7838), .ZN(n13583) );
  NAND2_X1 U9402 ( .A1(n7835), .A2(n7836), .ZN(n13582) );
  NAND2_X1 U9403 ( .A1(n13578), .A2(n7838), .ZN(n7835) );
  OAI21_X1 U9404 ( .B1(n13614), .B2(n7846), .A(n7844), .ZN(n13618) );
  NAND2_X1 U9405 ( .A1(n7841), .A2(n7842), .ZN(n13617) );
  NAND2_X1 U9406 ( .A1(n13614), .A2(n7844), .ZN(n7841) );
  OAI21_X1 U9407 ( .B1(n13657), .B2(n7851), .A(n7849), .ZN(n13661) );
  NAND2_X1 U9408 ( .A1(n7847), .A2(n7341), .ZN(n13660) );
  NAND2_X1 U9409 ( .A1(n13657), .A2(n7849), .ZN(n7847) );
  NAND2_X1 U9410 ( .A1(n13556), .A2(n7855), .ZN(n7853) );
  NAND2_X1 U9411 ( .A1(n7853), .A2(n7852), .ZN(n13561) );
  OAI21_X1 U9412 ( .B1(n13556), .B2(n7856), .A(n7855), .ZN(n13562) );
  AND2_X1 U9413 ( .A1(n13702), .A2(n13697), .ZN(n7870) );
  NAND2_X2 U9414 ( .A1(n14696), .A2(n14701), .ZN(n14695) );
  NAND2_X1 U9415 ( .A1(n15709), .A2(n7883), .ZN(n7880) );
  AOI21_X1 U9416 ( .B1(n7883), .B2(n7882), .A(n7280), .ZN(n7881) );
  NAND2_X1 U9417 ( .A1(n14625), .A2(n7889), .ZN(n7887) );
  OAI21_X1 U9418 ( .B1(n14625), .B2(n7893), .A(n7891), .ZN(n14569) );
  NAND2_X1 U9419 ( .A1(n7887), .A2(n7888), .ZN(n14571) );
  NAND2_X1 U9420 ( .A1(n14625), .A2(n7894), .ZN(n7890) );
  INV_X1 U9421 ( .A(n7897), .ZN(n7896) );
  NAND2_X2 U9422 ( .A1(n14886), .A2(n9500), .ZN(n8938) );
  INV_X2 U9423 ( .A(n7203), .ZN(n9416) );
  INV_X1 U9424 ( .A(n7906), .ZN(n7905) );
  NAND2_X1 U9425 ( .A1(n8619), .A2(n7925), .ZN(n7923) );
  NAND2_X1 U9426 ( .A1(n7942), .A2(n7349), .ZN(n8700) );
  NAND2_X1 U9427 ( .A1(n9359), .A2(n9358), .ZN(n7949) );
  NAND2_X1 U9428 ( .A1(n8160), .A2(SI_1_), .ZN(n8165) );
  NAND3_X1 U9429 ( .A1(n8266), .A2(n8162), .A3(n8165), .ZN(n8265) );
  INV_X1 U9430 ( .A(n7954), .ZN(n7953) );
  NAND3_X1 U9431 ( .A1(n8222), .A2(n7954), .A3(n7952), .ZN(n7955) );
  NAND3_X1 U9432 ( .A1(n14794), .A2(n8135), .A3(n14795), .ZN(n7956) );
  MUX2_X1 U9433 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n7956), .S(n15717), .Z(
        P1_U3557) );
  MUX2_X1 U9434 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n7956), .S(n15719), .Z(
        P1_U3525) );
  NAND2_X1 U9435 ( .A1(n15652), .A2(n11717), .ZN(n7958) );
  OAI21_X1 U9436 ( .B1(n14643), .B2(n7961), .A(n7959), .ZN(n14621) );
  NAND2_X1 U9437 ( .A1(n12449), .A2(n7968), .ZN(n7967) );
  NAND2_X1 U9438 ( .A1(n12095), .A2(n7983), .ZN(n7980) );
  INV_X1 U9439 ( .A(n14366), .ZN(n7989) );
  XNOR2_X2 U9440 ( .A(n8875), .B(n7990), .ZN(n8882) );
  AND3_X2 U9441 ( .A1(n8860), .A2(n7991), .A3(n8866), .ZN(n8887) );
  NAND2_X1 U9442 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  NAND2_X1 U9443 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
  NAND2_X1 U9444 ( .A1(n9152), .A2(n9153), .ZN(n9151) );
  NAND2_X1 U9445 ( .A1(n9254), .A2(n9255), .ZN(n9253) );
  NAND2_X1 U9446 ( .A1(n9222), .A2(n9223), .ZN(n9221) );
  AND2_X1 U9447 ( .A1(n8000), .A2(n8302), .ZN(n10418) );
  OAI21_X1 U9448 ( .B1(n9100), .B2(n7219), .A(n8004), .ZN(n9115) );
  INV_X1 U9449 ( .A(n8001), .ZN(n9114) );
  NAND2_X1 U9450 ( .A1(n8006), .A2(n8007), .ZN(n9319) );
  NAND2_X1 U9451 ( .A1(n9294), .A2(n7309), .ZN(n8006) );
  INV_X1 U9452 ( .A(n9293), .ZN(n8009) );
  NAND2_X1 U9453 ( .A1(n8014), .A2(n8016), .ZN(n9291) );
  NAND3_X1 U9454 ( .A1(n9259), .A2(n8015), .A3(n9258), .ZN(n8014) );
  INV_X1 U9455 ( .A(n9354), .ZN(n8030) );
  AOI21_X1 U9456 ( .B1(n8752), .B2(n8776), .A(n8756), .ZN(n8755) );
  NAND2_X1 U9457 ( .A1(n8547), .A2(n8738), .ZN(n8031) );
  NAND4_X1 U9458 ( .A1(n8036), .A2(n8035), .A3(n8033), .A4(n8034), .ZN(n8520)
         );
  AND2_X1 U9459 ( .A1(n8294), .A2(n8223), .ZN(n8318) );
  AND2_X2 U9460 ( .A1(n8294), .A2(n8226), .ZN(n8036) );
  NAND2_X1 U9461 ( .A1(n13441), .A2(n13442), .ZN(n11127) );
  NOR2_X2 U9462 ( .A1(n11123), .A2(n7288), .ZN(n10724) );
  XNOR2_X1 U9463 ( .A(n11104), .B(n13522), .ZN(n10710) );
  INV_X1 U9464 ( .A(n13447), .ZN(n8040) );
  NAND2_X1 U9465 ( .A1(n13447), .A2(n8045), .ZN(n8041) );
  NAND3_X1 U9466 ( .A1(n8044), .A2(n8046), .A3(n8041), .ZN(n13487) );
  NAND2_X1 U9467 ( .A1(n12526), .A2(n8051), .ZN(n8049) );
  NAND2_X1 U9468 ( .A1(n8049), .A2(n8048), .ZN(n11934) );
  INV_X1 U9469 ( .A(n12530), .ZN(n11852) );
  INV_X1 U9470 ( .A(n11291), .ZN(n8063) );
  AOI21_X2 U9471 ( .B1(n13510), .B2(n8066), .A(n8062), .ZN(n12592) );
  OAI21_X2 U9472 ( .B1(n12592), .B2(n11833), .A(n12590), .ZN(n12575) );
  NAND2_X1 U9473 ( .A1(n12614), .A2(n12613), .ZN(n12616) );
  NAND2_X1 U9474 ( .A1(n12612), .A2(n12611), .ZN(n8067) );
  NAND2_X1 U9475 ( .A1(n14303), .A2(n8083), .ZN(n8082) );
  NAND2_X1 U9476 ( .A1(n8092), .A2(n8089), .ZN(n12072) );
  NAND2_X1 U9477 ( .A1(n11865), .A2(n8090), .ZN(n8092) );
  INV_X1 U9478 ( .A(n8092), .ZN(n11946) );
  INV_X1 U9479 ( .A(n8097), .ZN(n9484) );
  NAND2_X1 U9480 ( .A1(n8097), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8096) );
  INV_X1 U9481 ( .A(n8099), .ZN(n11528) );
  NAND2_X1 U9482 ( .A1(n11533), .A2(n9681), .ZN(n11542) );
  NAND2_X1 U9483 ( .A1(n11855), .A2(n7217), .ZN(n8104) );
  INV_X1 U9484 ( .A(n8113), .ZN(n12263) );
  NAND2_X1 U9485 ( .A1(n11668), .A2(n9739), .ZN(n11792) );
  NAND2_X1 U9486 ( .A1(n9738), .A2(n11663), .ZN(n11668) );
  NAND2_X1 U9487 ( .A1(n9956), .A2(n8124), .ZN(n8123) );
  NAND2_X1 U9488 ( .A1(n9986), .A2(n9985), .ZN(n13078) );
  OAI21_X1 U9489 ( .B1(n13537), .B2(n13536), .A(n13535), .ZN(n13539) );
  XNOR2_X1 U9490 ( .A(n9359), .B(n9358), .ZN(n14224) );
  OR3_X1 U9491 ( .A1(n7209), .A2(n10063), .A3(n11070), .ZN(n10105) );
  NAND2_X1 U9492 ( .A1(n7209), .A2(n11070), .ZN(n11526) );
  NAND2_X1 U9493 ( .A1(n8939), .A2(n11503), .ZN(n11234) );
  INV_X1 U9494 ( .A(n11232), .ZN(n8962) );
  INV_X1 U9495 ( .A(n9597), .ZN(n13405) );
  OAI21_X1 U9496 ( .B1(n7259), .B2(n8756), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n8249) );
  NAND2_X1 U9497 ( .A1(n13989), .A2(n8821), .ZN(n13972) );
  AOI21_X2 U9498 ( .B1(n12448), .B2(n15914), .A(n12447), .ZN(n14801) );
  XNOR2_X1 U9499 ( .A(n8830), .B(n8829), .ZN(n8842) );
  OAI21_X1 U9500 ( .B1(n8216), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n8163), .ZN(
        n8164) );
  NAND2_X1 U9501 ( .A1(n8216), .A2(n9636), .ZN(n8163) );
  OAI21_X1 U9502 ( .B1(n8216), .B2(n10399), .A(n8159), .ZN(n8160) );
  NAND2_X1 U9503 ( .A1(n7204), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8159) );
  OAI21_X2 U9504 ( .B1(n11700), .B2(n11699), .A(n11698), .ZN(n15657) );
  NAND2_X2 U9505 ( .A1(n12082), .A2(n12081), .ZN(n12203) );
  OR2_X1 U9506 ( .A1(n8285), .A2(n8275), .ZN(n8280) );
  OR2_X1 U9507 ( .A1(n8285), .A2(n12506), .ZN(n8326) );
  NOR2_X2 U9508 ( .A1(n15762), .A2(n12048), .ZN(n12095) );
  NOR2_X1 U9509 ( .A1(n15763), .A2(n15768), .ZN(n15762) );
  NAND2_X1 U9510 ( .A1(n8870), .A2(n8889), .ZN(n9500) );
  OAI21_X1 U9511 ( .B1(n14098), .B2(n13980), .A(n8850), .ZN(n8851) );
  NAND2_X1 U9512 ( .A1(n8302), .A2(n8171), .ZN(n8312) );
  XNOR2_X1 U9513 ( .A(n14569), .B(n12467), .ZN(n12448) );
  NAND2_X1 U9514 ( .A1(n9421), .A2(n9420), .ZN(n9520) );
  INV_X1 U9515 ( .A(n14029), .ZN(n8818) );
  XNOR2_X1 U9516 ( .A(n14373), .B(n15620), .ZN(n11366) );
  NAND2_X1 U9517 ( .A1(n9484), .A2(n9483), .ZN(n9490) );
  INV_X1 U9518 ( .A(n11682), .ZN(n11680) );
  OR2_X1 U9519 ( .A1(n11201), .A2(n11200), .ZN(n11202) );
  INV_X1 U9520 ( .A(n13758), .ZN(n11419) );
  INV_X1 U9521 ( .A(n13760), .ZN(n8802) );
  AND3_X1 U9522 ( .A1(n13528), .A2(n13553), .A3(n13529), .ZN(n8134) );
  AND2_X1 U9523 ( .A1(n10722), .A2(n10721), .ZN(n13507) );
  AND2_X2 U9524 ( .A1(n11193), .A2(n15139), .ZN(n14215) );
  AND2_X1 U9525 ( .A1(n8844), .A2(n13959), .ZN(n15818) );
  INV_X1 U9526 ( .A(n13223), .ZN(n13229) );
  AND2_X1 U9527 ( .A1(n14793), .A2(n14792), .ZN(n8135) );
  OR2_X1 U9528 ( .A1(n13057), .A2(n13391), .ZN(n8136) );
  OR2_X1 U9529 ( .A1(n13057), .A2(n13316), .ZN(n8137) );
  AND2_X1 U9530 ( .A1(n14374), .A2(n11516), .ZN(n8139) );
  OR2_X1 U9531 ( .A1(n14374), .A2(n11516), .ZN(n8140) );
  INV_X1 U9532 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8937) );
  OR2_X1 U9533 ( .A1(n8938), .A2(n8926), .ZN(n8144) );
  XNOR2_X1 U9534 ( .A(n10990), .B(n10912), .ZN(n10992) );
  AND2_X1 U9535 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8145) );
  INV_X1 U9536 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8756) );
  INV_X1 U9537 ( .A(n11357), .ZN(n10320) );
  INV_X1 U9538 ( .A(n14360), .ZN(n14717) );
  OR2_X1 U9539 ( .A1(n14099), .A2(n14085), .ZN(n8146) );
  INV_X1 U9540 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9696) );
  INV_X1 U9541 ( .A(n9486), .ZN(n9493) );
  AND2_X1 U9542 ( .A1(n13795), .A2(n14076), .ZN(n8147) );
  INV_X1 U9543 ( .A(n8306), .ZN(n8341) );
  INV_X4 U9544 ( .A(n14772), .ZN(n15941) );
  AND2_X1 U9545 ( .A1(n10061), .A2(n10150), .ZN(n13240) );
  INV_X1 U9546 ( .A(n13240), .ZN(n15577) );
  AND2_X1 U9547 ( .A1(n10276), .A2(n10148), .ZN(n8148) );
  OR2_X1 U9548 ( .A1(n11249), .A2(n11261), .ZN(n15924) );
  OR2_X1 U9549 ( .A1(n11249), .A2(n11218), .ZN(n15926) );
  AND2_X1 U9550 ( .A1(n9457), .A2(n9464), .ZN(n8149) );
  INV_X1 U9551 ( .A(n12464), .ZN(n14599) );
  NOR2_X1 U9552 ( .A1(n12908), .A2(n13276), .ZN(n8150) );
  INV_X1 U9553 ( .A(n14841), .ZN(n12438) );
  INV_X1 U9554 ( .A(n10305), .ZN(n13215) );
  NOR2_X1 U9555 ( .A1(n13103), .A2(n13101), .ZN(n8151) );
  OAI22_X1 U9556 ( .A1(n13197), .A2(n9917), .B1(n13213), .B2(n13206), .ZN(
        n13184) );
  OR2_X1 U9557 ( .A1(n13553), .A2(n13529), .ZN(n13526) );
  NOR2_X1 U9558 ( .A1(n13530), .A2(n13529), .ZN(n13531) );
  NAND2_X1 U9559 ( .A1(n13533), .A2(n13532), .ZN(n13536) );
  NAND2_X1 U9560 ( .A1(n9268), .A2(n11516), .ZN(n8958) );
  NAND2_X1 U9561 ( .A1(n13552), .A2(n13551), .ZN(n13556) );
  INV_X1 U9562 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9574) );
  AND2_X1 U9563 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  AND2_X1 U9564 ( .A1(n14658), .A2(n14656), .ZN(n12459) );
  NAND2_X1 U9565 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  INV_X1 U9566 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U9567 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  INV_X1 U9568 ( .A(n8866), .ZN(n8867) );
  NOR2_X1 U9569 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  INV_X1 U9570 ( .A(n10272), .ZN(n10018) );
  INV_X1 U9571 ( .A(n12267), .ZN(n9843) );
  INV_X1 U9572 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9577) );
  AND2_X1 U9573 ( .A1(n8688), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8706) );
  NOR2_X1 U9574 ( .A1(n8589), .A2(n13451), .ZN(n8604) );
  NOR2_X1 U9575 ( .A1(n8491), .A2(n8490), .ZN(n8489) );
  INV_X1 U9576 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8229) );
  INV_X1 U9577 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8738) );
  AND2_X1 U9578 ( .A1(n11432), .A2(n11431), .ZN(n11433) );
  NAND2_X1 U9579 ( .A1(n7192), .A2(n15527), .ZN(n10352) );
  INV_X1 U9580 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9087) );
  INV_X1 U9581 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8871) );
  INV_X1 U9582 ( .A(n8582), .ZN(n8583) );
  INV_X1 U9583 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9756) );
  INV_X1 U9584 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9823) );
  INV_X1 U9585 ( .A(n12897), .ZN(n12876) );
  INV_X1 U9586 ( .A(n10785), .ZN(n10791) );
  INV_X1 U9587 ( .A(n12971), .ZN(n15405) );
  OAI22_X1 U9588 ( .A1(n13077), .A2(n15575), .B1(n13047), .B2(n11032), .ZN(
        n10039) );
  AND2_X1 U9589 ( .A1(n10105), .A2(n10285), .ZN(n10895) );
  AND2_X1 U9590 ( .A1(n10195), .A2(n10196), .ZN(n11796) );
  AND3_X1 U9591 ( .A1(n10108), .A2(n10106), .A3(n10109), .ZN(n10789) );
  INV_X1 U9592 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10121) );
  INV_X1 U9593 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U9594 ( .A1(n8405), .A2(n12584), .ZN(n8404) );
  AND2_X1 U9595 ( .A1(n10694), .A2(n10967), .ZN(n10696) );
  OR2_X1 U9596 ( .A1(n8623), .A2(n13422), .ZN(n8641) );
  OR2_X1 U9597 ( .A1(n8570), .A2(n13477), .ZN(n8589) );
  NAND2_X1 U9598 ( .A1(n8241), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8570) );
  OR2_X1 U9599 ( .A1(n8389), .A2(n8388), .ZN(n8405) );
  INV_X2 U9600 ( .A(n10329), .ZN(n8548) );
  INV_X1 U9601 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8245) );
  INV_X1 U9602 ( .A(n11759), .ZN(n11760) );
  INV_X1 U9603 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9200) );
  OR2_X1 U9604 ( .A1(n12657), .A2(n12656), .ZN(n12658) );
  AND2_X1 U9605 ( .A1(n14899), .A2(n9387), .ZN(n10359) );
  NAND2_X1 U9606 ( .A1(n9503), .A2(n8149), .ZN(n9511) );
  NOR2_X1 U9607 ( .A1(n9088), .A2(n9087), .ZN(n9119) );
  OR2_X1 U9608 ( .A1(n14848), .A2(n12454), .ZN(n12437) );
  OR2_X1 U9609 ( .A1(n12281), .A2(n14364), .ZN(n12204) );
  INV_X1 U9610 ( .A(n8961), .ZN(n8939) );
  NOR2_X1 U9611 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9494) );
  INV_X1 U9612 ( .A(SI_22_), .ZN(n15019) );
  NAND2_X1 U9613 ( .A1(n8203), .A2(SI_13_), .ZN(n8206) );
  INV_X1 U9614 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15273) );
  OR2_X1 U9615 ( .A1(n9837), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9850) );
  AND2_X1 U9616 ( .A1(n9740), .A2(n15090), .ZN(n9757) );
  NOR2_X1 U9617 ( .A1(n9802), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9824) );
  AND2_X1 U9618 ( .A1(n9866), .A2(n12829), .ZN(n9896) );
  NAND2_X1 U9619 ( .A1(n9824), .A2(n9823), .ZN(n9837) );
  NAND2_X1 U9620 ( .A1(n10791), .A2(n10790), .ZN(n15126) );
  OR2_X1 U9621 ( .A1(n9641), .A2(n9631), .ZN(n9632) );
  AND2_X1 U9622 ( .A1(n10824), .A2(n10822), .ZN(n10825) );
  INV_X1 U9623 ( .A(n13136), .ZN(n13149) );
  NOR2_X1 U9624 ( .A1(n9723), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9740) );
  INV_X1 U9625 ( .A(n10803), .ZN(n10782) );
  AND2_X1 U9626 ( .A1(n13393), .A2(n10773), .ZN(n10803) );
  AND2_X1 U9627 ( .A1(n10208), .A2(n12172), .ZN(n12138) );
  OR2_X1 U9628 ( .A1(n10788), .A2(n10285), .ZN(n15575) );
  NAND2_X1 U9629 ( .A1(n10788), .A2(n10286), .ZN(n13243) );
  INV_X1 U9630 ( .A(n13408), .ZN(n12726) );
  XNOR2_X1 U9631 ( .A(n10710), .B(n10711), .ZN(n13441) );
  INV_X1 U9632 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11843) );
  INV_X1 U9633 ( .A(n13813), .ZN(n11118) );
  NAND2_X1 U9634 ( .A1(n12363), .A2(n12358), .ZN(n12359) );
  INV_X1 U9635 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n12584) );
  INV_X1 U9636 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U9637 ( .A1(n11274), .A2(n11273), .ZN(n11275) );
  AND2_X1 U9638 ( .A1(n10696), .A2(n15140), .ZN(n10722) );
  AND2_X1 U9639 ( .A1(n8707), .A2(n8690), .ZN(n13924) );
  OR2_X1 U9640 ( .A1(n8525), .A2(n8524), .ZN(n8536) );
  NAND2_X1 U9641 ( .A1(n10720), .A2(n10341), .ZN(n14057) );
  XNOR2_X1 U9642 ( .A(n13544), .B(n12511), .ZN(n13749) );
  OR2_X1 U9643 ( .A1(n15818), .A2(n8845), .ZN(n15821) );
  INV_X1 U9644 ( .A(n13753), .ZN(n11448) );
  INV_X1 U9645 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8246) );
  INV_X1 U9646 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8336) );
  INV_X1 U9647 ( .A(n11767), .ZN(n11768) );
  OR2_X1 U9648 ( .A1(n9159), .A2(n9158), .ZN(n9175) );
  AND2_X1 U9649 ( .A1(n9119), .A2(n8879), .ZN(n9135) );
  NOR2_X1 U9650 ( .A1(n9201), .A2(n9200), .ZN(n9210) );
  AND2_X1 U9651 ( .A1(n9281), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9295) );
  NOR2_X1 U9652 ( .A1(n10990), .A2(n10989), .ZN(n10991) );
  OR2_X1 U9653 ( .A1(n9175), .A2(n9174), .ZN(n9201) );
  NAND2_X1 U9654 ( .A1(n9466), .A2(n12259), .ZN(n9467) );
  OR2_X1 U9655 ( .A1(n10364), .A2(n10363), .ZN(n10383) );
  NAND2_X1 U9656 ( .A1(n14356), .A2(n14767), .ZN(n12445) );
  INV_X1 U9657 ( .A(n15964), .ZN(n14737) );
  INV_X1 U9658 ( .A(n14361), .ZN(n15904) );
  OR2_X1 U9659 ( .A1(n9070), .A2(n9069), .ZN(n9088) );
  INV_X1 U9660 ( .A(n11214), .ZN(n10633) );
  INV_X1 U9661 ( .A(n15919), .ZN(n15887) );
  OR2_X1 U9662 ( .A1(n10628), .A2(n9500), .ZN(n15903) );
  OR2_X1 U9663 ( .A1(n10629), .A2(n10628), .ZN(n15901) );
  AND2_X1 U9664 ( .A1(n8685), .A2(n8672), .ZN(n8683) );
  INV_X1 U9665 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8903) );
  AND2_X1 U9666 ( .A1(n8186), .A2(n8185), .ZN(n8366) );
  INV_X1 U9667 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8979) );
  AOI21_X1 U9668 ( .B1(n15399), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n15277), .ZN(
        n15290) );
  OR2_X1 U9669 ( .A1(n10320), .A2(n10803), .ZN(n10824) );
  AND3_X1 U9670 ( .A1(n9939), .A2(n9938), .A3(n9937), .ZN(n13157) );
  INV_X1 U9671 ( .A(n15491), .ZN(n15503) );
  AND2_X1 U9672 ( .A1(n10825), .A2(n12955), .ZN(n15514) );
  INV_X1 U9673 ( .A(n15575), .ZN(n15547) );
  AND3_X1 U9674 ( .A1(n10110), .A2(n10803), .A3(n10109), .ZN(n10897) );
  INV_X1 U9675 ( .A(n13316), .ZN(n15971) );
  INV_X1 U9676 ( .A(n15797), .ZN(n15737) );
  INV_X1 U9677 ( .A(n15733), .ZN(n15632) );
  NAND2_X1 U9678 ( .A1(n10081), .A2(n10080), .ZN(n10106) );
  INV_X1 U9679 ( .A(n9591), .ZN(n9592) );
  XNOR2_X1 U9680 ( .A(n10094), .B(n10093), .ZN(n10804) );
  NAND2_X1 U9681 ( .A1(n10026), .A2(n10021), .ZN(n10030) );
  INV_X1 U9682 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9861) );
  INV_X1 U9683 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9706) );
  NOR2_X1 U9684 ( .A1(n12576), .A2(n11835), .ZN(n11836) );
  INV_X1 U9685 ( .A(n13499), .ZN(n13438) );
  INV_X1 U9686 ( .A(n13500), .ZN(n13439) );
  INV_X1 U9687 ( .A(n13484), .ZN(n13428) );
  NOR2_X1 U9688 ( .A1(n12535), .A2(n7278), .ZN(n13498) );
  NOR2_X1 U9689 ( .A1(n10695), .A2(n13740), .ZN(n13513) );
  AND2_X1 U9690 ( .A1(n8665), .A2(n8664), .ZN(n13664) );
  OR2_X1 U9691 ( .A1(n10326), .A2(n10325), .ZN(n10332) );
  OR2_X1 U9692 ( .A1(n8285), .A2(n8284), .ZN(n8288) );
  AND2_X1 U9693 ( .A1(n15141), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15210) );
  NAND2_X1 U9694 ( .A1(n14042), .A2(n8563), .ZN(n14027) );
  INV_X1 U9695 ( .A(n14055), .ZN(n14069) );
  AND2_X1 U9696 ( .A1(n15869), .A2(n15861), .ZN(n14127) );
  AND2_X1 U9697 ( .A1(n10966), .A2(n14902), .ZN(n11193) );
  INV_X1 U9698 ( .A(n14159), .ZN(n15859) );
  OR2_X1 U9699 ( .A1(n14235), .A2(n8768), .ZN(n8769) );
  NAND2_X1 U9700 ( .A1(n8744), .A2(n8743), .ZN(n8746) );
  AND2_X1 U9701 ( .A1(n8472), .A2(n8502), .ZN(n15209) );
  AND2_X1 U9702 ( .A1(n10397), .A2(P2_U3088), .ZN(n14234) );
  INV_X1 U9703 ( .A(n14326), .ZN(n15960) );
  AOI21_X1 U9704 ( .B1(n10993), .B2(n10992), .A(n10991), .ZN(n11204) );
  NAND2_X1 U9705 ( .A1(n10635), .A2(n14584), .ZN(n15965) );
  AND4_X1 U9706 ( .A1(n9352), .A2(n9351), .A3(n9350), .A4(n9349), .ZN(n12444)
         );
  AND4_X1 U9707 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n15902)
         );
  AND4_X1 U9708 ( .A1(n9166), .A2(n9165), .A3(n9164), .A4(n9163), .ZN(n12604)
         );
  OR2_X1 U9709 ( .A1(n10737), .A2(n10736), .ZN(n11019) );
  INV_X1 U9710 ( .A(n14548), .ZN(n14546) );
  INV_X1 U9711 ( .A(n14672), .ZN(n15935) );
  INV_X1 U9712 ( .A(n14740), .ZN(n15936) );
  NAND2_X1 U9713 ( .A1(n10619), .A2(n14874), .ZN(n11261) );
  INV_X1 U9714 ( .A(n15914), .ZN(n15890) );
  INV_X1 U9715 ( .A(n11261), .ZN(n11218) );
  AND2_X1 U9716 ( .A1(n10824), .A2(n10823), .ZN(n15502) );
  INV_X1 U9717 ( .A(n12900), .ZN(n11990) );
  AND2_X1 U9718 ( .A1(n10138), .A2(n10038), .ZN(n11032) );
  INV_X1 U9719 ( .A(n13158), .ZN(n12909) );
  INV_X1 U9720 ( .A(n12838), .ZN(n13225) );
  INV_X1 U9721 ( .A(P3_U3897), .ZN(n12925) );
  INV_X1 U9722 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15399) );
  INV_X1 U9723 ( .A(n15502), .ZN(n15417) );
  INV_X1 U9724 ( .A(n15517), .ZN(n15500) );
  AND2_X1 U9725 ( .A1(n13109), .A2(n13108), .ZN(n13271) );
  NAND2_X2 U9726 ( .A1(n10901), .A2(n13143), .ZN(n15688) );
  NAND2_X1 U9727 ( .A1(n15839), .A2(n15737), .ZN(n13316) );
  AND3_X2 U9728 ( .A1(n10114), .A2(n10897), .A3(n10113), .ZN(n15839) );
  INV_X2 U9729 ( .A(n15980), .ZN(n15978) );
  CLKBUF_X1 U9730 ( .A(n10483), .Z(n10505) );
  OR2_X1 U9731 ( .A1(n10804), .A2(P3_U3151), .ZN(n11357) );
  INV_X1 U9732 ( .A(SI_18_), .ZN(n15041) );
  INV_X1 U9733 ( .A(SI_12_), .ZN(n15053) );
  INV_X1 U9734 ( .A(n11153), .ZN(n12972) );
  INV_X1 U9735 ( .A(n15198), .ZN(n15200) );
  INV_X1 U9736 ( .A(n11111), .ZN(n11276) );
  AND2_X1 U9737 ( .A1(n10704), .A2(n13959), .ZN(n13506) );
  INV_X1 U9738 ( .A(n13665), .ZN(n13794) );
  INV_X1 U9739 ( .A(n15205), .ZN(n15180) );
  INV_X1 U9740 ( .A(n15210), .ZN(n15158) );
  INV_X1 U9741 ( .A(n7197), .ZN(n13980) );
  OR2_X1 U9742 ( .A1(n13980), .A2(n8785), .ZN(n14085) );
  OR2_X1 U9743 ( .A1(n15818), .A2(n11253), .ZN(n14066) );
  INV_X1 U9744 ( .A(n15869), .ZN(n15868) );
  AND2_X2 U9745 ( .A1(n11193), .A2(n10967), .ZN(n15869) );
  AND3_X1 U9746 ( .A1(n15867), .A2(n15866), .A3(n15865), .ZN(n15872) );
  INV_X1 U9747 ( .A(n14215), .ZN(n15870) );
  OR2_X1 U9748 ( .A1(n15137), .A2(n14904), .ZN(n14905) );
  NAND2_X1 U9749 ( .A1(n8770), .A2(n8769), .ZN(n15139) );
  INV_X1 U9750 ( .A(n11400), .ZN(n12033) );
  INV_X1 U9751 ( .A(n14604), .ZN(n14804) );
  INV_X1 U9752 ( .A(n14651), .ZN(n14823) );
  OR2_X1 U9753 ( .A1(n10632), .A2(n10622), .ZN(n15949) );
  INV_X1 U9754 ( .A(n12444), .ZN(n14357) );
  INV_X1 U9755 ( .A(n12604), .ZN(n14362) );
  INV_X1 U9756 ( .A(n14551), .ZN(n14518) );
  OR2_X1 U9757 ( .A1(n10364), .A2(n10362), .ZN(n14557) );
  OR2_X1 U9758 ( .A1(n15941), .A2(n12115), .ZN(n14740) );
  INV_X1 U9759 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14894) );
  INV_X1 U9760 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11909) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10983) );
  INV_X1 U9762 ( .A(n14880), .ZN(n14897) );
  INV_X1 U9763 ( .A(n13812), .ZN(P2_U3947) );
  NAND2_X1 U9764 ( .A1(n8146), .A2(n8852), .ZN(P2_U3236) );
  NAND4_X1 U9765 ( .A1(n8154), .A2(n8153), .A3(n8152), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n8158) );
  NAND4_X1 U9766 ( .A1(n8156), .A2(n8155), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n8157) );
  INV_X1 U9767 ( .A(n8160), .ZN(n8161) );
  INV_X1 U9768 ( .A(SI_1_), .ZN(n14953) );
  NAND2_X1 U9769 ( .A1(n8161), .A2(n14953), .ZN(n8162) );
  INV_X1 U9770 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9636) );
  NOR2_X1 U9771 ( .A1(n8164), .A2(n15067), .ZN(n8266) );
  INV_X1 U9772 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10417) );
  MUX2_X1 U9773 ( .A(n10424), .B(n10417), .S(n8216), .Z(n8291) );
  NOR2_X1 U9774 ( .A1(n8291), .A2(n15075), .ZN(n8170) );
  MUX2_X1 U9775 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8216), .Z(n8166) );
  NAND2_X1 U9776 ( .A1(n8166), .A2(SI_3_), .ZN(n8171) );
  OAI21_X1 U9777 ( .B1(n8166), .B2(SI_3_), .A(n8171), .ZN(n8300) );
  INV_X1 U9778 ( .A(n8291), .ZN(n8167) );
  NOR2_X1 U9779 ( .A1(n8167), .A2(SI_2_), .ZN(n8168) );
  NOR2_X1 U9780 ( .A1(n8300), .A2(n8168), .ZN(n8169) );
  MUX2_X1 U9781 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8216), .Z(n8172) );
  NAND2_X1 U9782 ( .A1(n8172), .A2(SI_4_), .ZN(n8174) );
  OAI21_X1 U9783 ( .B1(n8172), .B2(SI_4_), .A(n8174), .ZN(n8313) );
  INV_X1 U9784 ( .A(n8313), .ZN(n8173) );
  MUX2_X1 U9785 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8216), .Z(n8175) );
  NAND2_X1 U9786 ( .A1(n8175), .A2(SI_5_), .ZN(n8178) );
  INV_X1 U9787 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9788 ( .A1(n8176), .A2(n10406), .ZN(n8177) );
  AND2_X1 U9789 ( .A1(n8178), .A2(n8177), .ZN(n8329) );
  MUX2_X1 U9790 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7204), .Z(n8179) );
  NAND2_X1 U9791 ( .A1(n8179), .A2(SI_6_), .ZN(n8182) );
  INV_X1 U9792 ( .A(n8179), .ZN(n8180) );
  INV_X1 U9793 ( .A(SI_6_), .ZN(n10401) );
  NAND2_X1 U9794 ( .A1(n8180), .A2(n10401), .ZN(n8181) );
  NAND2_X1 U9795 ( .A1(n8351), .A2(n8350), .ZN(n8353) );
  MUX2_X1 U9796 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8216), .Z(n8183) );
  NAND2_X1 U9797 ( .A1(n8183), .A2(SI_7_), .ZN(n8186) );
  INV_X1 U9798 ( .A(n8183), .ZN(n8184) );
  INV_X1 U9799 ( .A(SI_7_), .ZN(n15062) );
  NAND2_X1 U9800 ( .A1(n8184), .A2(n15062), .ZN(n8185) );
  MUX2_X1 U9801 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7204), .Z(n8187) );
  NAND2_X1 U9802 ( .A1(n8187), .A2(SI_8_), .ZN(n8189) );
  OAI21_X1 U9803 ( .B1(SI_8_), .B2(n8187), .A(n8189), .ZN(n8382) );
  INV_X1 U9804 ( .A(n8382), .ZN(n8188) );
  MUX2_X1 U9805 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n10397), .Z(n8190) );
  NAND2_X1 U9806 ( .A1(n8190), .A2(SI_9_), .ZN(n8193) );
  INV_X1 U9807 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U9808 ( .A1(n8191), .A2(n14910), .ZN(n8192) );
  NAND2_X1 U9809 ( .A1(n8399), .A2(n8193), .ZN(n8414) );
  MUX2_X1 U9810 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10397), .Z(n8194) );
  NAND2_X1 U9811 ( .A1(n8194), .A2(SI_10_), .ZN(n8197) );
  INV_X1 U9812 ( .A(n8194), .ZN(n8195) );
  NAND2_X1 U9813 ( .A1(n8195), .A2(n14909), .ZN(n8196) );
  MUX2_X1 U9814 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n8216), .Z(n8198) );
  XNOR2_X1 U9815 ( .A(n8198), .B(SI_11_), .ZN(n8432) );
  INV_X1 U9816 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U9817 ( .A1(n8199), .A2(n15057), .ZN(n8200) );
  MUX2_X1 U9818 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8216), .Z(n8201) );
  XNOR2_X1 U9819 ( .A(n8201), .B(n15053), .ZN(n8446) );
  INV_X1 U9820 ( .A(n8201), .ZN(n8202) );
  MUX2_X1 U9821 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n10397), .Z(n8203) );
  OAI21_X1 U9822 ( .B1(n8203), .B2(SI_13_), .A(n8206), .ZN(n8462) );
  MUX2_X1 U9823 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n10397), .Z(n8207) );
  INV_X1 U9824 ( .A(n8207), .ZN(n8208) );
  NAND2_X1 U9825 ( .A1(n8208), .A2(n14943), .ZN(n8209) );
  MUX2_X1 U9826 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n10397), .Z(n8210) );
  XNOR2_X1 U9827 ( .A(n8210), .B(n15046), .ZN(n8500) );
  NAND2_X1 U9828 ( .A1(n8501), .A2(n8500), .ZN(n8213) );
  INV_X1 U9829 ( .A(n8210), .ZN(n8211) );
  NAND2_X1 U9830 ( .A1(n8211), .A2(n15046), .ZN(n8212) );
  NAND2_X1 U9831 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  INV_X1 U9832 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11402) );
  MUX2_X1 U9833 ( .A(n11402), .B(n11399), .S(n10397), .Z(n8515) );
  MUX2_X1 U9834 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n10397), .Z(n8217) );
  XNOR2_X1 U9835 ( .A(n8217), .B(SI_17_), .ZN(n8529) );
  INV_X1 U9836 ( .A(n8217), .ZN(n8218) );
  NAND2_X1 U9837 ( .A1(n8220), .A2(n15041), .ZN(n8221) );
  MUX2_X1 U9838 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n10397), .Z(n8543) );
  MUX2_X1 U9839 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n10397), .Z(n8564) );
  XNOR2_X1 U9840 ( .A(n8566), .B(n8565), .ZN(n12017) );
  NOR2_X2 U9841 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8227) );
  INV_X1 U9842 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8231) );
  INV_X1 U9843 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8230) );
  NOR2_X1 U9844 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n8233) );
  NOR2_X1 U9845 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n8232) );
  XNOR2_X2 U9846 ( .A(n8236), .B(n8235), .ZN(n10341) );
  NAND2_X2 U9847 ( .A1(n10341), .A2(n14231), .ZN(n10329) );
  NAND2_X1 U9848 ( .A1(n12017), .A2(n13704), .ZN(n8240) );
  NOR2_X2 U9849 ( .A1(n8238), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8778) );
  XNOR2_X2 U9850 ( .A(n8752), .B(P2_IR_REG_19__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U9851 ( .A1(n8420), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8548), .B2(
        n15194), .ZN(n8239) );
  AND2_X1 U9852 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8322) );
  NAND2_X1 U9853 ( .A1(n8322), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8359) );
  INV_X1 U9854 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8358) );
  NOR2_X1 U9855 ( .A1(n8359), .A2(n8358), .ZN(n8357) );
  NAND2_X1 U9856 ( .A1(n8357), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8389) );
  INV_X1 U9857 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8388) );
  INV_X1 U9858 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U9859 ( .A1(n8489), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8525) );
  INV_X1 U9860 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8524) );
  INV_X1 U9861 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8535) );
  INV_X1 U9862 ( .A(n8241), .ZN(n8554) );
  INV_X1 U9863 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9864 ( .A1(n8554), .A2(n8242), .ZN(n8243) );
  NAND2_X1 U9865 ( .A1(n8570), .A2(n8243), .ZN(n14049) );
  NAND2_X1 U9866 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8245), .ZN(n8248) );
  OR2_X1 U9867 ( .A1(n14049), .A2(n8285), .ZN(n8259) );
  AND2_X2 U9868 ( .A1(n8252), .A2(n8254), .ZN(n8306) );
  INV_X1 U9869 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14152) );
  NAND2_X1 U9870 ( .A1(n8709), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8256) );
  NAND2_X2 U9871 ( .A1(n8254), .A2(n14226), .ZN(n8572) );
  INV_X4 U9872 ( .A(n8572), .ZN(n8555) );
  NAND2_X1 U9873 ( .A1(n8555), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8255) );
  OAI211_X1 U9874 ( .C1(n8341), .C2(n14152), .A(n8256), .B(n8255), .ZN(n8257)
         );
  INV_X1 U9875 ( .A(n8257), .ZN(n8258) );
  NAND2_X1 U9876 ( .A1(n8259), .A2(n8258), .ZN(n14072) );
  XNOR2_X1 U9877 ( .A(n14048), .B(n14072), .ZN(n14054) );
  INV_X1 U9878 ( .A(n14054), .ZN(n14044) );
  NAND2_X1 U9879 ( .A1(n8477), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U9880 ( .A1(n8306), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8263) );
  INV_X1 U9881 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U9882 ( .A1(n8323), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8261) );
  INV_X1 U9883 ( .A(n8266), .ZN(n8267) );
  NAND2_X1 U9884 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  NAND2_X1 U9885 ( .A1(n8265), .A2(n8269), .ZN(n10415) );
  INV_X1 U9886 ( .A(n10415), .ZN(n8270) );
  NAND2_X1 U9887 ( .A1(n13704), .A2(n8270), .ZN(n8274) );
  NAND2_X1 U9888 ( .A1(n7198), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U9889 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8271) );
  XNOR2_X1 U9890 ( .A(n8271), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10594) );
  INV_X1 U9891 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U9892 ( .A1(n8306), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8279) );
  INV_X1 U9893 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U9894 ( .A1(n8323), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8277) );
  NOR2_X1 U9895 ( .A1(n7204), .A2(n15067), .ZN(n8281) );
  XNOR2_X1 U9896 ( .A(n8281), .B(n9521), .ZN(n14245) );
  MUX2_X1 U9897 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14245), .S(n10329), .Z(n13523)
         );
  NAND2_X1 U9898 ( .A1(n8282), .A2(n10968), .ZN(n10969) );
  NAND2_X1 U9899 ( .A1(n13521), .A2(n13522), .ZN(n8283) );
  NAND2_X1 U9900 ( .A1(n10969), .A2(n8283), .ZN(n11318) );
  NAND2_X1 U9901 ( .A1(n8306), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8289) );
  INV_X1 U9902 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U9903 ( .A1(n8555), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9904 ( .A1(n8323), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8286) );
  OR2_X1 U9905 ( .A1(n8292), .A2(n8291), .ZN(n8301) );
  NAND2_X1 U9906 ( .A1(n8292), .A2(n8291), .ZN(n8293) );
  OR2_X1 U9907 ( .A1(n8294), .A2(n8756), .ZN(n8295) );
  AOI22_X1 U9908 ( .A1(n8420), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8548), .B2(
        n13824), .ZN(n8296) );
  OAI21_X2 U9909 ( .B1(n10423), .B2(n8519), .A(n8296), .ZN(n13540) );
  NAND2_X1 U9910 ( .A1(n11004), .A2(n13540), .ZN(n11007) );
  INV_X1 U9911 ( .A(n13540), .ZN(n15604) );
  NAND2_X1 U9912 ( .A1(n15604), .A2(n13815), .ZN(n8297) );
  INV_X1 U9913 ( .A(n13747), .ZN(n11321) );
  NAND2_X1 U9914 ( .A1(n11318), .A2(n11321), .ZN(n11317) );
  NAND2_X1 U9915 ( .A1(n15604), .A2(n11004), .ZN(n8298) );
  NAND2_X1 U9916 ( .A1(n11317), .A2(n8298), .ZN(n11003) );
  NAND2_X1 U9917 ( .A1(n10418), .A2(n13704), .ZN(n8305) );
  XNOR2_X1 U9918 ( .A(n8303), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13836) );
  AOI22_X1 U9919 ( .A1(n8420), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8548), .B2(
        n13836), .ZN(n8304) );
  NAND2_X1 U9920 ( .A1(n8306), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8310) );
  INV_X1 U9921 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13833) );
  NAND2_X1 U9922 ( .A1(n8477), .A2(n13833), .ZN(n8309) );
  NAND2_X1 U9923 ( .A1(n8555), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U9924 ( .A1(n8323), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8307) );
  NAND4_X1 U9925 ( .A1(n8310), .A2(n8309), .A3(n8308), .A4(n8307), .ZN(n13814)
         );
  NAND2_X1 U9926 ( .A1(n11003), .A2(n13749), .ZN(n11002) );
  INV_X1 U9927 ( .A(n13544), .ZN(n11576) );
  NAND2_X1 U9928 ( .A1(n11576), .A2(n12511), .ZN(n8311) );
  NAND2_X1 U9929 ( .A1(n8314), .A2(n8313), .ZN(n8316) );
  AND2_X1 U9930 ( .A1(n8316), .A2(n8315), .ZN(n10412) );
  NAND2_X1 U9931 ( .A1(n10412), .A2(n13704), .ZN(n8321) );
  INV_X1 U9932 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U9933 ( .A1(n8318), .A2(n8317), .ZN(n8333) );
  NAND2_X1 U9934 ( .A1(n8333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U9935 ( .A(n8319), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U9936 ( .A1(n7198), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8548), .B2(
        n10646), .ZN(n8320) );
  NAND2_X1 U9937 ( .A1(n8321), .A2(n8320), .ZN(n13554) );
  NAND2_X1 U9938 ( .A1(n8834), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8327) );
  INV_X1 U9939 ( .A(n8322), .ZN(n8343) );
  OAI21_X1 U9940 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8343), .ZN(n12506) );
  NAND2_X1 U9941 ( .A1(n8555), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U9942 ( .A1(n8323), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8324) );
  XNOR2_X1 U9943 ( .A(n13554), .B(n11118), .ZN(n13750) );
  OR2_X1 U9944 ( .A1(n13813), .A2(n13554), .ZN(n8328) );
  OR2_X1 U9945 ( .A1(n8330), .A2(n8329), .ZN(n8331) );
  AND2_X1 U9946 ( .A1(n8332), .A2(n8331), .ZN(n10426) );
  NAND2_X1 U9947 ( .A1(n10426), .A2(n13704), .ZN(n8340) );
  NOR2_X1 U9948 ( .A1(n8333), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8337) );
  INV_X1 U9949 ( .A(n8337), .ZN(n8334) );
  NAND2_X1 U9950 ( .A1(n8334), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8335) );
  MUX2_X1 U9951 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8335), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8338) );
  NAND2_X1 U9952 ( .A1(n8337), .A2(n8336), .ZN(n8370) );
  NAND2_X1 U9953 ( .A1(n8338), .A2(n8370), .ZN(n10676) );
  INV_X1 U9954 ( .A(n10676), .ZN(n10640) );
  AOI22_X1 U9955 ( .A1(n8420), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8548), .B2(
        n10640), .ZN(n8339) );
  NAND2_X1 U9956 ( .A1(n8340), .A2(n8339), .ZN(n13559) );
  INV_X2 U9957 ( .A(n8341), .ZN(n8834) );
  NAND2_X1 U9958 ( .A1(n8834), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8348) );
  INV_X1 U9959 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U9960 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  AND2_X1 U9961 ( .A1(n8359), .A2(n8344), .ZN(n11403) );
  NAND2_X1 U9962 ( .A1(n8477), .A2(n11403), .ZN(n8347) );
  NAND2_X1 U9963 ( .A1(n8709), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U9964 ( .A1(n8555), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8345) );
  NAND4_X1 U9965 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8345), .ZN(n13811)
         );
  INV_X1 U9966 ( .A(n13811), .ZN(n12507) );
  XNOR2_X1 U9967 ( .A(n13559), .B(n12507), .ZN(n13751) );
  OR2_X1 U9968 ( .A1(n13559), .A2(n13811), .ZN(n8349) );
  NAND2_X1 U9969 ( .A1(n11135), .A2(n8349), .ZN(n11097) );
  OR2_X1 U9970 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U9971 ( .A1(n8353), .A2(n8352), .ZN(n10432) );
  OR2_X1 U9972 ( .A1(n10432), .A2(n8519), .ZN(n8356) );
  NAND2_X1 U9973 ( .A1(n8370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8354) );
  XNOR2_X1 U9974 ( .A(n8354), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U9975 ( .A1(n7198), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8548), .B2(
        n10648), .ZN(n8355) );
  NAND2_X1 U9976 ( .A1(n8356), .A2(n8355), .ZN(n13567) );
  NAND2_X1 U9977 ( .A1(n8834), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8364) );
  INV_X1 U9978 ( .A(n8357), .ZN(n8375) );
  NAND2_X1 U9979 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  AND2_X1 U9980 ( .A1(n8375), .A2(n8360), .ZN(n13514) );
  NAND2_X1 U9981 ( .A1(n8477), .A2(n13514), .ZN(n8363) );
  NAND2_X1 U9982 ( .A1(n8709), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U9983 ( .A1(n8555), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8361) );
  NAND4_X1 U9984 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(n13810)
         );
  XNOR2_X1 U9985 ( .A(n13567), .B(n13810), .ZN(n13754) );
  INV_X1 U9986 ( .A(n13754), .ZN(n11101) );
  NAND2_X1 U9987 ( .A1(n11097), .A2(n11101), .ZN(n11096) );
  INV_X1 U9988 ( .A(n13567), .ZN(n11558) );
  INV_X1 U9989 ( .A(n13810), .ZN(n11114) );
  NAND2_X1 U9990 ( .A1(n11558), .A2(n11114), .ZN(n8365) );
  NAND2_X1 U9991 ( .A1(n11096), .A2(n8365), .ZN(n11446) );
  OR2_X1 U9992 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U9993 ( .A1(n8369), .A2(n8368), .ZN(n10435) );
  OR2_X1 U9994 ( .A1(n10435), .A2(n8519), .ZN(n8373) );
  NAND2_X1 U9995 ( .A1(n8384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8371) );
  XNOR2_X1 U9996 ( .A(n8371), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U9997 ( .A1(n8420), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8548), .B2(
        n10683), .ZN(n8372) );
  NAND2_X1 U9998 ( .A1(n8373), .A2(n8372), .ZN(n13576) );
  NAND2_X1 U9999 ( .A1(n8834), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8380) );
  INV_X1 U10000 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10001 ( .A1(n8375), .A2(n8374), .ZN(n8376) );
  AND2_X1 U10002 ( .A1(n8389), .A2(n8376), .ZN(n11456) );
  NAND2_X1 U10003 ( .A1(n8477), .A2(n11456), .ZN(n8379) );
  NAND2_X1 U10004 ( .A1(n8555), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10005 ( .A1(n8709), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8377) );
  NAND4_X1 U10006 ( .A1(n8380), .A2(n8379), .A3(n8378), .A4(n8377), .ZN(n13809) );
  XNOR2_X1 U10007 ( .A(n13576), .B(n13809), .ZN(n13753) );
  OR2_X1 U10008 ( .A1(n13576), .A2(n13809), .ZN(n8381) );
  NAND2_X1 U10009 ( .A1(n10450), .A2(n13704), .ZN(n8387) );
  NAND2_X1 U10010 ( .A1(n8400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8385) );
  XNOR2_X1 U10011 ( .A(n8385), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U10012 ( .A1(n8420), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8548), .B2(
        n10752), .ZN(n8386) );
  NAND2_X1 U10013 ( .A1(n8387), .A2(n8386), .ZN(n13580) );
  NAND2_X1 U10014 ( .A1(n8834), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10015 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  AND2_X1 U10016 ( .A1(n8405), .A2(n8390), .ZN(n11425) );
  NAND2_X1 U10017 ( .A1(n8477), .A2(n11425), .ZN(n8393) );
  NAND2_X1 U10018 ( .A1(n8709), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10019 ( .A1(n8555), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8391) );
  NAND4_X1 U10020 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n13808) );
  XNOR2_X1 U10021 ( .A(n13580), .B(n12488), .ZN(n13758) );
  NAND2_X1 U10022 ( .A1(n13580), .A2(n13808), .ZN(n8395) );
  NAND2_X1 U10023 ( .A1(n11417), .A2(n8395), .ZN(n11461) );
  OR2_X1 U10024 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U10025 ( .A1(n8399), .A2(n8398), .ZN(n10455) );
  OR2_X1 U10026 ( .A1(n10455), .A2(n8519), .ZN(n8403) );
  NAND2_X1 U10027 ( .A1(n8417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8401) );
  XNOR2_X1 U10028 ( .A(n8401), .B(P2_IR_REG_9__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U10029 ( .A1(n7198), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n13860), 
        .B2(n8548), .ZN(n8402) );
  NAND2_X1 U10030 ( .A1(n8403), .A2(n8402), .ZN(n13587) );
  NAND2_X1 U10031 ( .A1(n8834), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8410) );
  INV_X1 U10032 ( .A(n8404), .ZN(n8425) );
  NAND2_X1 U10033 ( .A1(n8405), .A2(n12584), .ZN(n8406) );
  AND2_X1 U10034 ( .A1(n8425), .A2(n8406), .ZN(n12588) );
  NAND2_X1 U10035 ( .A1(n8477), .A2(n12588), .ZN(n8409) );
  NAND2_X1 U10036 ( .A1(n8555), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10037 ( .A1(n8709), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8407) );
  NAND4_X1 U10038 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n13807) );
  XNOR2_X1 U10039 ( .A(n13587), .B(n13807), .ZN(n13756) );
  INV_X1 U10040 ( .A(n13756), .ZN(n8799) );
  NAND2_X1 U10041 ( .A1(n11461), .A2(n8799), .ZN(n8412) );
  NAND2_X1 U10042 ( .A1(n13587), .A2(n13807), .ZN(n8411) );
  OR2_X1 U10043 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  NAND2_X1 U10044 ( .A1(n8416), .A2(n8415), .ZN(n10460) );
  OR2_X1 U10045 ( .A1(n10460), .A2(n8519), .ZN(n8422) );
  INV_X1 U10046 ( .A(n8435), .ZN(n8418) );
  NAND2_X1 U10047 ( .A1(n8418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8419) );
  XNOR2_X1 U10048 ( .A(n8419), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U10049 ( .A1(n11078), .A2(n8548), .B1(n7198), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U10050 ( .A1(n8306), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8430) );
  INV_X1 U10051 ( .A(n8423), .ZN(n8440) );
  INV_X1 U10052 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10053 ( .A1(n8425), .A2(n8424), .ZN(n8426) );
  AND2_X1 U10054 ( .A1(n8440), .A2(n8426), .ZN(n12571) );
  NAND2_X1 U10055 ( .A1(n8477), .A2(n12571), .ZN(n8429) );
  NAND2_X1 U10056 ( .A1(n8555), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10057 ( .A1(n8709), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8427) );
  NAND4_X1 U10058 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n13806) );
  INV_X1 U10059 ( .A(n13806), .ZN(n11823) );
  XNOR2_X1 U10060 ( .A(n13591), .B(n11823), .ZN(n13759) );
  NAND2_X1 U10061 ( .A1(n13591), .A2(n13806), .ZN(n8431) );
  INV_X1 U10062 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8434) );
  INV_X1 U10063 ( .A(n8449), .ZN(n8436) );
  NAND2_X1 U10064 ( .A1(n8436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8437) );
  XNOR2_X1 U10065 ( .A(n8437), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U10066 ( .A1(n13873), .A2(n8548), .B1(n8420), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10067 ( .A1(n8834), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8445) );
  INV_X1 U10068 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10069 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  AND2_X1 U10070 ( .A1(n8454), .A2(n8441), .ZN(n15817) );
  NAND2_X1 U10071 ( .A1(n8477), .A2(n15817), .ZN(n8444) );
  NAND2_X1 U10072 ( .A1(n8555), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10073 ( .A1(n8709), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8442) );
  NAND4_X1 U10074 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), .ZN(n13805) );
  INV_X1 U10075 ( .A(n13805), .ZN(n8803) );
  XNOR2_X1 U10076 ( .A(n13600), .B(n8803), .ZN(n13760) );
  XNOR2_X1 U10077 ( .A(n8447), .B(n8446), .ZN(n10582) );
  NAND2_X1 U10078 ( .A1(n10582), .A2(n13704), .ZN(n8453) );
  INV_X1 U10079 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8448) );
  INV_X1 U10080 ( .A(n8467), .ZN(n8450) );
  NAND2_X1 U10081 ( .A1(n8450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8451) );
  XNOR2_X1 U10082 ( .A(n8451), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U10083 ( .A1(n11086), .A2(n8548), .B1(n7198), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10084 ( .A1(n8834), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10085 ( .A1(n8454), .A2(n11843), .ZN(n8455) );
  AND2_X1 U10086 ( .A1(n8475), .A2(n8455), .ZN(n11848) );
  NAND2_X1 U10087 ( .A1(n8477), .A2(n11848), .ZN(n8458) );
  NAND2_X1 U10088 ( .A1(n8555), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10089 ( .A1(n8709), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8456) );
  NAND4_X1 U10090 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n13804) );
  XNOR2_X1 U10091 ( .A(n13603), .B(n13804), .ZN(n13761) );
  INV_X1 U10092 ( .A(n13761), .ZN(n8805) );
  NAND2_X1 U10093 ( .A1(n11804), .A2(n8805), .ZN(n8461) );
  NAND2_X1 U10094 ( .A1(n13603), .A2(n13804), .ZN(n8460) );
  NAND2_X1 U10095 ( .A1(n8461), .A2(n8460), .ZN(n12002) );
  NAND2_X1 U10096 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NAND2_X1 U10097 ( .A1(n8465), .A2(n8464), .ZN(n10692) );
  OR2_X1 U10098 ( .A1(n10692), .A2(n8519), .ZN(n8474) );
  INV_X1 U10099 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10100 ( .A1(n8467), .A2(n8466), .ZN(n8469) );
  NAND2_X1 U10101 ( .A1(n8469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8468) );
  MUX2_X1 U10102 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8468), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8472) );
  INV_X1 U10103 ( .A(n8469), .ZN(n8471) );
  INV_X1 U10104 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10105 ( .A1(n8471), .A2(n8470), .ZN(n8502) );
  AOI22_X1 U10106 ( .A1(n15209), .A2(n8548), .B1(n8420), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10107 ( .A1(n8306), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10108 ( .A1(n8475), .A2(n11935), .ZN(n8476) );
  AND2_X1 U10109 ( .A1(n8491), .A2(n8476), .ZN(n12011) );
  NAND2_X1 U10110 ( .A1(n8477), .A2(n12011), .ZN(n8480) );
  NAND2_X1 U10111 ( .A1(n8555), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10112 ( .A1(n8709), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8478) );
  NAND4_X1 U10113 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n13803) );
  XNOR2_X1 U10114 ( .A(n13612), .B(n13803), .ZN(n13762) );
  INV_X1 U10115 ( .A(n13762), .ZN(n12006) );
  NAND2_X1 U10116 ( .A1(n12002), .A2(n12006), .ZN(n8483) );
  NAND2_X1 U10117 ( .A1(n13612), .A2(n13803), .ZN(n8482) );
  XNOR2_X1 U10118 ( .A(n8485), .B(n8484), .ZN(n10980) );
  NAND2_X1 U10119 ( .A1(n10980), .A2(n13704), .ZN(n8488) );
  NAND2_X1 U10120 ( .A1(n8502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8486) );
  XNOR2_X1 U10121 ( .A(n8486), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U10122 ( .A1(n11388), .A2(n8548), .B1(n8420), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8487) );
  INV_X1 U10123 ( .A(n8489), .ZN(n8509) );
  NAND2_X1 U10124 ( .A1(n8491), .A2(n8490), .ZN(n8492) );
  AND2_X1 U10125 ( .A1(n8509), .A2(n8492), .ZN(n12494) );
  NAND2_X1 U10126 ( .A1(n12494), .A2(n8477), .ZN(n8496) );
  NAND2_X1 U10127 ( .A1(n8306), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10128 ( .A1(n8555), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10129 ( .A1(n8709), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8493) );
  NAND4_X1 U10130 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n13802) );
  XNOR2_X1 U10131 ( .A(n15862), .B(n13802), .ZN(n13764) );
  INV_X1 U10132 ( .A(n13764), .ZN(n8497) );
  NAND2_X1 U10133 ( .A1(n12058), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U10134 ( .A1(n15862), .A2(n13802), .ZN(n8498) );
  NAND2_X1 U10135 ( .A1(n8499), .A2(n8498), .ZN(n12182) );
  XNOR2_X1 U10136 ( .A(n8501), .B(n8500), .ZN(n11167) );
  NAND2_X1 U10137 ( .A1(n11167), .A2(n13704), .ZN(n8505) );
  OAI21_X1 U10138 ( .B1(n8502), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U10139 ( .A(n8503), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U10140 ( .A1(n11971), .A2(n8548), .B1(n7198), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8504) );
  INV_X1 U10141 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U10142 ( .A1(n8834), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10143 ( .A1(n8555), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8506) );
  AND2_X1 U10144 ( .A1(n8507), .A2(n8506), .ZN(n8512) );
  INV_X1 U10145 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10146 ( .A1(n8509), .A2(n8508), .ZN(n8510) );
  NAND2_X1 U10147 ( .A1(n8525), .A2(n8510), .ZN(n12341) );
  OR2_X1 U10148 ( .A1(n8285), .A2(n12341), .ZN(n8511) );
  OAI211_X1 U10149 ( .C1(n8513), .C2(n12190), .A(n8512), .B(n8511), .ZN(n13801) );
  INV_X1 U10150 ( .A(n13801), .ZN(n8813) );
  XNOR2_X1 U10151 ( .A(n13622), .B(n8813), .ZN(n13766) );
  OR2_X1 U10152 ( .A1(n13622), .A2(n13801), .ZN(n8514) );
  NAND2_X1 U10153 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  NAND2_X1 U10154 ( .A1(n8518), .A2(n8517), .ZN(n11401) );
  OR2_X1 U10155 ( .A1(n11401), .A2(n8519), .ZN(n8523) );
  NAND2_X1 U10156 ( .A1(n8520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8521) );
  XNOR2_X1 U10157 ( .A(n8521), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U10158 ( .A1(n8420), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8548), 
        .B2(n11400), .ZN(n8522) );
  NAND2_X1 U10159 ( .A1(n8525), .A2(n8524), .ZN(n8526) );
  NAND2_X1 U10160 ( .A1(n8536), .A2(n8526), .ZN(n12396) );
  AOI22_X1 U10161 ( .A1(n8306), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8555), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10162 ( .A1(n8709), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8527) );
  OAI211_X1 U10163 ( .C1(n12396), .C2(n8285), .A(n8528), .B(n8527), .ZN(n13800) );
  INV_X1 U10164 ( .A(n13800), .ZN(n12373) );
  XNOR2_X1 U10165 ( .A(n13626), .B(n12373), .ZN(n13767) );
  INV_X1 U10166 ( .A(n13767), .ZN(n12382) );
  XNOR2_X1 U10167 ( .A(n8530), .B(n8529), .ZN(n11674) );
  NAND2_X1 U10168 ( .A1(n11674), .A2(n13704), .ZN(n8533) );
  NAND2_X1 U10169 ( .A1(n8238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U10170 ( .A(n8531), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U10171 ( .A1(n7198), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8548), 
        .B2(n15174), .ZN(n8532) );
  INV_X1 U10172 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12376) );
  INV_X1 U10173 ( .A(n8534), .ZN(n8552) );
  NAND2_X1 U10174 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U10175 ( .A1(n8552), .A2(n8537), .ZN(n12375) );
  OR2_X1 U10176 ( .A1(n12375), .A2(n8285), .ZN(n8539) );
  AOI22_X1 U10177 ( .A1(n8834), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8555), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8538) );
  OAI211_X1 U10178 ( .C1(n8513), .C2(n12376), .A(n8539), .B(n8538), .ZN(n14070) );
  XNOR2_X1 U10179 ( .A(n13635), .B(n14070), .ZN(n13768) );
  INV_X1 U10180 ( .A(n13768), .ZN(n8540) );
  NAND2_X1 U10181 ( .A1(n12370), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U10182 ( .A1(n13635), .A2(n14070), .ZN(n8541) );
  INV_X1 U10183 ( .A(n8543), .ZN(n8544) );
  NAND2_X1 U10184 ( .A1(n7291), .A2(n8544), .ZN(n8545) );
  NAND2_X1 U10185 ( .A1(n11906), .A2(n13704), .ZN(n8550) );
  XNOR2_X1 U10186 ( .A(n8547), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U10187 ( .A1(n8420), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8548), 
        .B2(n15175), .ZN(n8549) );
  INV_X1 U10188 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10189 ( .A1(n8552), .A2(n8551), .ZN(n8553) );
  AND2_X1 U10190 ( .A1(n8554), .A2(n8553), .ZN(n14078) );
  NAND2_X1 U10191 ( .A1(n14078), .A2(n8477), .ZN(n8561) );
  INV_X1 U10192 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10193 ( .A1(n8555), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10194 ( .A1(n8709), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U10195 ( .C1(n8341), .C2(n8558), .A(n8557), .B(n8556), .ZN(n8559)
         );
  INV_X1 U10196 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U10197 ( .A1(n8561), .A2(n8560), .ZN(n13799) );
  XNOR2_X1 U10198 ( .A(n14155), .B(n13799), .ZN(n14084) );
  OR2_X1 U10199 ( .A1(n14155), .A2(n13799), .ZN(n8562) );
  OR2_X1 U10200 ( .A1(n14048), .A2(n14072), .ZN(n8563) );
  INV_X1 U10201 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12131) );
  MUX2_X1 U10202 ( .A(n12131), .B(n12112), .S(n10397), .Z(n8582) );
  XNOR2_X1 U10203 ( .A(n8582), .B(SI_20_), .ZN(n8567) );
  XNOR2_X1 U10204 ( .A(n8586), .B(n8567), .ZN(n12111) );
  NAND2_X1 U10205 ( .A1(n12111), .A2(n13704), .ZN(n8569) );
  NAND2_X1 U10206 ( .A1(n7198), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8568) );
  INV_X1 U10207 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U10208 ( .A1(n8570), .A2(n13477), .ZN(n8571) );
  AND2_X1 U10209 ( .A1(n8589), .A2(n8571), .ZN(n14036) );
  NAND2_X1 U10210 ( .A1(n14036), .A2(n8477), .ZN(n8578) );
  INV_X1 U10211 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10212 ( .A1(n8306), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10213 ( .A1(n8709), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8573) );
  OAI211_X1 U10214 ( .C1(n8572), .C2(n8575), .A(n8574), .B(n8573), .ZN(n8576)
         );
  INV_X1 U10215 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U10216 ( .A1(n8578), .A2(n8577), .ZN(n13798) );
  NAND2_X1 U10217 ( .A1(n14146), .A2(n13798), .ZN(n8579) );
  NAND2_X1 U10218 ( .A1(n14027), .A2(n8579), .ZN(n8581) );
  OR2_X1 U10219 ( .A1(n14146), .A2(n13798), .ZN(n8580) );
  NOR2_X1 U10220 ( .A1(n8583), .A2(SI_20_), .ZN(n8585) );
  NAND2_X1 U10221 ( .A1(n8583), .A2(SI_20_), .ZN(n8584) );
  MUX2_X1 U10222 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n10397), .Z(n8601) );
  XNOR2_X1 U10223 ( .A(n8601), .B(SI_21_), .ZN(n8598) );
  XNOR2_X1 U10224 ( .A(n8600), .B(n8598), .ZN(n12216) );
  NAND2_X1 U10225 ( .A1(n12216), .A2(n13704), .ZN(n8588) );
  NAND2_X1 U10226 ( .A1(n7198), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8587) );
  INV_X1 U10227 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13451) );
  INV_X1 U10228 ( .A(n8604), .ZN(n8605) );
  NAND2_X1 U10229 ( .A1(n8589), .A2(n13451), .ZN(n8590) );
  NAND2_X1 U10230 ( .A1(n8605), .A2(n8590), .ZN(n13450) );
  OR2_X1 U10231 ( .A1(n13450), .A2(n8285), .ZN(n8596) );
  INV_X1 U10232 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U10233 ( .A1(n8306), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U10234 ( .A1(n8709), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8591) );
  OAI211_X1 U10235 ( .C1(n8572), .C2(n8593), .A(n8592), .B(n8591), .ZN(n8594)
         );
  INV_X1 U10236 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U10237 ( .A1(n8596), .A2(n8595), .ZN(n13797) );
  NAND2_X1 U10238 ( .A1(n14141), .A2(n13797), .ZN(n8597) );
  NAND2_X1 U10239 ( .A1(n8600), .A2(n8599), .ZN(n8616) );
  NAND2_X1 U10240 ( .A1(n8601), .A2(SI_21_), .ZN(n8613) );
  NAND2_X1 U10241 ( .A1(n8616), .A2(n8613), .ZN(n8602) );
  INV_X1 U10242 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12479) );
  INV_X1 U10243 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9565) );
  MUX2_X1 U10244 ( .A(n12479), .B(n9565), .S(n10397), .Z(n8617) );
  NAND2_X1 U10245 ( .A1(n7198), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U10246 ( .A1(n8604), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8623) );
  INV_X1 U10247 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U10248 ( .A1(n8605), .A2(n13491), .ZN(n8606) );
  NAND2_X1 U10249 ( .A1(n8623), .A2(n8606), .ZN(n13490) );
  OR2_X1 U10250 ( .A1(n13490), .A2(n8285), .ZN(n8611) );
  INV_X1 U10251 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14206) );
  NAND2_X1 U10252 ( .A1(n8834), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10253 ( .A1(n8709), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8607) );
  OAI211_X1 U10254 ( .C1(n8572), .C2(n14206), .A(n8608), .B(n8607), .ZN(n8609)
         );
  INV_X1 U10255 ( .A(n8609), .ZN(n8610) );
  NAND2_X1 U10256 ( .A1(n8611), .A2(n8610), .ZN(n13796) );
  NAND2_X1 U10257 ( .A1(n14010), .A2(n13796), .ZN(n8612) );
  OAI21_X1 U10258 ( .B1(n8617), .B2(n15019), .A(n8613), .ZN(n8614) );
  INV_X1 U10259 ( .A(n8614), .ZN(n8615) );
  NAND2_X1 U10260 ( .A1(n8616), .A2(n8615), .ZN(n8619) );
  NAND2_X1 U10261 ( .A1(n8617), .A2(n15019), .ZN(n8618) );
  INV_X1 U10262 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8620) );
  MUX2_X1 U10263 ( .A(n9610), .B(n8620), .S(n10397), .Z(n8634) );
  XNOR2_X1 U10264 ( .A(n8634), .B(SI_23_), .ZN(n8633) );
  XNOR2_X1 U10265 ( .A(n8638), .B(n8633), .ZN(n12256) );
  NAND2_X1 U10266 ( .A1(n12256), .A2(n13704), .ZN(n8622) );
  NAND2_X1 U10267 ( .A1(n8420), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8621) );
  INV_X1 U10268 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U10269 ( .A1(n8623), .A2(n13422), .ZN(n8624) );
  NAND2_X1 U10270 ( .A1(n8641), .A2(n8624), .ZN(n13420) );
  OR2_X1 U10271 ( .A1(n13420), .A2(n8285), .ZN(n8629) );
  INV_X1 U10272 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U10273 ( .A1(n8306), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10274 ( .A1(n8709), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8625) );
  OAI211_X1 U10275 ( .C1(n14202), .C2(n8572), .A(n8626), .B(n8625), .ZN(n8627)
         );
  INV_X1 U10276 ( .A(n8627), .ZN(n8628) );
  NAND2_X1 U10277 ( .A1(n8629), .A2(n8628), .ZN(n13795) );
  XNOR2_X1 U10278 ( .A(n13994), .B(n13795), .ZN(n13990) );
  INV_X1 U10279 ( .A(n13990), .ZN(n8630) );
  NAND2_X1 U10280 ( .A1(n13988), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U10281 ( .A1(n13994), .A2(n13795), .ZN(n8631) );
  NAND2_X1 U10282 ( .A1(n8632), .A2(n8631), .ZN(n13970) );
  INV_X1 U10283 ( .A(n8633), .ZN(n8637) );
  INV_X1 U10284 ( .A(n8634), .ZN(n8635) );
  NAND2_X1 U10285 ( .A1(n8635), .A2(SI_23_), .ZN(n8636) );
  MUX2_X1 U10286 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n10397), .Z(n8653) );
  XNOR2_X1 U10287 ( .A(n8653), .B(SI_24_), .ZN(n8650) );
  XNOR2_X1 U10288 ( .A(n8652), .B(n8650), .ZN(n14241) );
  NAND2_X1 U10289 ( .A1(n14241), .A2(n13704), .ZN(n8640) );
  NAND2_X1 U10290 ( .A1(n7198), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8639) );
  INV_X1 U10291 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U10292 ( .A1(n8641), .A2(n13469), .ZN(n8642) );
  AND2_X1 U10293 ( .A1(n8659), .A2(n8642), .ZN(n13981) );
  NAND2_X1 U10294 ( .A1(n13981), .A2(n8477), .ZN(n8647) );
  INV_X1 U10295 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14198) );
  NAND2_X1 U10296 ( .A1(n8834), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10297 ( .A1(n8709), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8643) );
  OAI211_X1 U10298 ( .C1(n8572), .C2(n14198), .A(n8644), .B(n8643), .ZN(n8645)
         );
  INV_X1 U10299 ( .A(n8645), .ZN(n8646) );
  NAND2_X1 U10300 ( .A1(n14126), .A2(n13665), .ZN(n13950) );
  OR2_X1 U10301 ( .A1(n14126), .A2(n13665), .ZN(n8648) );
  NAND2_X1 U10302 ( .A1(n13950), .A2(n8648), .ZN(n13971) );
  OR2_X1 U10303 ( .A1(n14200), .A2(n13665), .ZN(n8649) );
  INV_X1 U10304 ( .A(n8650), .ZN(n8651) );
  INV_X1 U10305 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14240) );
  MUX2_X1 U10306 ( .A(n14240), .B(n14894), .S(n10397), .Z(n8654) );
  NAND2_X1 U10307 ( .A1(n8654), .A2(n15017), .ZN(n8667) );
  INV_X1 U10308 ( .A(n8654), .ZN(n8655) );
  NAND2_X1 U10309 ( .A1(n8655), .A2(SI_25_), .ZN(n8656) );
  NAND2_X1 U10310 ( .A1(n8667), .A2(n8656), .ZN(n8668) );
  XNOR2_X1 U10311 ( .A(n8669), .B(n8668), .ZN(n14237) );
  NAND2_X1 U10312 ( .A1(n14237), .A2(n13704), .ZN(n8658) );
  NAND2_X1 U10313 ( .A1(n8420), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8657) );
  INV_X1 U10314 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13463) );
  INV_X1 U10315 ( .A(n8675), .ZN(n8676) );
  NAND2_X1 U10316 ( .A1(n8659), .A2(n13463), .ZN(n8660) );
  NAND2_X1 U10317 ( .A1(n8676), .A2(n8660), .ZN(n13960) );
  OR2_X1 U10318 ( .A1(n13960), .A2(n8285), .ZN(n8665) );
  INV_X1 U10319 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14193) );
  NAND2_X1 U10320 ( .A1(n8306), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U10321 ( .A1(n8709), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8661) );
  OAI211_X1 U10322 ( .C1(n8572), .C2(n14193), .A(n8662), .B(n8661), .ZN(n8663)
         );
  INV_X1 U10323 ( .A(n8663), .ZN(n8664) );
  NAND2_X1 U10324 ( .A1(n13965), .A2(n13664), .ZN(n8666) );
  INV_X1 U10325 ( .A(n13966), .ZN(n13951) );
  OAI21_X2 U10326 ( .B1(n8669), .B2(n8668), .A(n8667), .ZN(n8684) );
  INV_X1 U10327 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9959) );
  INV_X1 U10328 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14891) );
  MUX2_X1 U10329 ( .A(n9959), .B(n14891), .S(n10397), .Z(n8670) );
  INV_X1 U10330 ( .A(SI_26_), .ZN(n14927) );
  NAND2_X1 U10331 ( .A1(n8670), .A2(n14927), .ZN(n8685) );
  INV_X1 U10332 ( .A(n8670), .ZN(n8671) );
  NAND2_X1 U10333 ( .A1(n8671), .A2(SI_26_), .ZN(n8672) );
  NAND2_X1 U10334 ( .A1(n14233), .A2(n13704), .ZN(n8674) );
  NAND2_X1 U10335 ( .A1(n8420), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8673) );
  INV_X1 U10336 ( .A(n8688), .ZN(n8689) );
  INV_X1 U10337 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U10338 ( .A1(n8676), .A2(n12566), .ZN(n8677) );
  NAND2_X1 U10339 ( .A1(n8689), .A2(n8677), .ZN(n13942) );
  OR2_X1 U10340 ( .A1(n13942), .A2(n8285), .ZN(n8682) );
  INV_X1 U10341 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U10342 ( .A1(n8834), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U10343 ( .A1(n8709), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8678) );
  OAI211_X1 U10344 ( .C1(n8572), .C2(n14189), .A(n8679), .B(n8678), .ZN(n8680)
         );
  INV_X1 U10345 ( .A(n8680), .ZN(n8681) );
  NAND2_X1 U10346 ( .A1(n8682), .A2(n8681), .ZN(n13792) );
  INV_X1 U10347 ( .A(n13792), .ZN(n13411) );
  XNOR2_X1 U10348 ( .A(n13944), .B(n13411), .ZN(n13933) );
  INV_X1 U10349 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14232) );
  INV_X1 U10350 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14888) );
  MUX2_X1 U10351 ( .A(n14232), .B(n14888), .S(n10397), .Z(n8697) );
  XNOR2_X1 U10352 ( .A(n8697), .B(SI_27_), .ZN(n8696) );
  NAND2_X1 U10353 ( .A1(n14230), .A2(n13704), .ZN(n8687) );
  NAND2_X1 U10354 ( .A1(n8420), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8686) );
  INV_X1 U10355 ( .A(n8706), .ZN(n8707) );
  INV_X1 U10356 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U10357 ( .A1(n8689), .A2(n13412), .ZN(n8690) );
  INV_X1 U10358 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14185) );
  NAND2_X1 U10359 ( .A1(n8306), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U10360 ( .A1(n8709), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8691) );
  OAI211_X1 U10361 ( .C1(n14185), .C2(n8572), .A(n8692), .B(n8691), .ZN(n8693)
         );
  XNOR2_X1 U10362 ( .A(n13923), .B(n13693), .ZN(n13913) );
  INV_X1 U10363 ( .A(n13913), .ZN(n13920) );
  OR2_X1 U10364 ( .A1(n14187), .A2(n13693), .ZN(n8694) );
  INV_X1 U10365 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U10366 ( .A1(n8698), .A2(SI_27_), .ZN(n8699) );
  NAND2_X1 U10367 ( .A1(n8700), .A2(n8699), .ZN(n8719) );
  INV_X1 U10368 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9993) );
  INV_X1 U10369 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14885) );
  MUX2_X1 U10370 ( .A(n9993), .B(n14885), .S(n10397), .Z(n8701) );
  NAND2_X1 U10371 ( .A1(n8701), .A2(n14919), .ZN(n8717) );
  INV_X1 U10372 ( .A(n8701), .ZN(n8702) );
  NAND2_X1 U10373 ( .A1(n8702), .A2(SI_28_), .ZN(n8703) );
  NAND2_X1 U10374 ( .A1(n8717), .A2(n8703), .ZN(n8718) );
  NAND2_X1 U10375 ( .A1(n14227), .A2(n13704), .ZN(n8705) );
  NAND2_X1 U10376 ( .A1(n8420), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10377 ( .A1(n8706), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8846) );
  INV_X1 U10378 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U10379 ( .A1(n8707), .A2(n12733), .ZN(n8708) );
  NAND2_X1 U10380 ( .A1(n8846), .A2(n8708), .ZN(n13897) );
  OR2_X1 U10381 ( .A1(n13897), .A2(n8285), .ZN(n8715) );
  INV_X1 U10382 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U10383 ( .A1(n8834), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U10384 ( .A1(n8709), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8710) );
  OAI211_X1 U10385 ( .C1(n8572), .C2(n8712), .A(n8711), .B(n8710), .ZN(n8713)
         );
  INV_X1 U10386 ( .A(n8713), .ZN(n8714) );
  NAND2_X1 U10387 ( .A1(n14104), .A2(n13690), .ZN(n8716) );
  NAND2_X1 U10388 ( .A1(n8828), .A2(n8716), .ZN(n13900) );
  INV_X1 U10389 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14225) );
  MUX2_X1 U10390 ( .A(n14225), .B(n10121), .S(n10397), .Z(n9360) );
  XNOR2_X1 U10391 ( .A(n9360), .B(SI_29_), .ZN(n9358) );
  NAND2_X1 U10392 ( .A1(n14224), .A2(n13704), .ZN(n8721) );
  NAND2_X1 U10393 ( .A1(n7198), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8720) );
  OR2_X1 U10394 ( .A1(n8846), .A2(n8285), .ZN(n8727) );
  INV_X1 U10395 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U10396 ( .A1(n8306), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10397 ( .A1(n8709), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U10398 ( .C1(n8572), .C2(n8724), .A(n8723), .B(n8722), .ZN(n8725)
         );
  INV_X1 U10399 ( .A(n8725), .ZN(n8726) );
  AND2_X1 U10400 ( .A1(n8727), .A2(n8726), .ZN(n13689) );
  INV_X1 U10401 ( .A(n13689), .ZN(n13789) );
  XNOR2_X1 U10402 ( .A(n14096), .B(n13789), .ZN(n13774) );
  XNOR2_X1 U10403 ( .A(n8728), .B(n13774), .ZN(n14099) );
  NOR4_X1 U10404 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n8737) );
  OR4_X1 U10405 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8734) );
  NOR4_X1 U10406 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8732) );
  NOR4_X1 U10407 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8731) );
  NOR4_X1 U10408 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8730) );
  NOR4_X1 U10409 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8729) );
  NAND4_X1 U10410 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n8733)
         );
  NOR4_X1 U10411 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n8734), .A4(n8733), .ZN(n8736) );
  NOR4_X1 U10412 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8735) );
  NAND3_X1 U10413 ( .A1(n8737), .A2(n8736), .A3(n8735), .ZN(n8751) );
  NAND2_X1 U10414 ( .A1(n8778), .A2(n8738), .ZN(n8781) );
  INV_X1 U10415 ( .A(n8781), .ZN(n8739) );
  NAND2_X1 U10416 ( .A1(n8739), .A2(n8141), .ZN(n8753) );
  NAND2_X1 U10417 ( .A1(n8761), .A2(n8763), .ZN(n8740) );
  NAND2_X1 U10418 ( .A1(n8748), .A2(n8747), .ZN(n8741) );
  INV_X1 U10419 ( .A(P2_B_REG_SCAN_IN), .ZN(n8837) );
  XOR2_X1 U10420 ( .A(n14242), .B(n8837), .Z(n8749) );
  NAND2_X1 U10421 ( .A1(n14238), .A2(n8749), .ZN(n8750) );
  AND2_X1 U10422 ( .A1(n8751), .A2(n14904), .ZN(n10693) );
  INV_X1 U10423 ( .A(n8784), .ZN(n8754) );
  NAND2_X1 U10424 ( .A1(n13736), .A2(n13776), .ZN(n13740) );
  NAND2_X1 U10425 ( .A1(n13740), .A2(n13779), .ZN(n13709) );
  NOR2_X1 U10426 ( .A1(n13709), .A2(n7193), .ZN(n10698) );
  NOR2_X1 U10427 ( .A1(n10693), .A2(n10698), .ZN(n10964) );
  NOR2_X1 U10428 ( .A1(n14238), .A2(n14242), .ZN(n8760) );
  NAND2_X1 U10429 ( .A1(n14235), .A2(n8760), .ZN(n10326) );
  INV_X1 U10430 ( .A(n8761), .ZN(n8762) );
  NAND2_X1 U10431 ( .A1(n8762), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8764) );
  INV_X1 U10432 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14903) );
  NAND2_X1 U10433 ( .A1(n14904), .A2(n14903), .ZN(n8767) );
  INV_X1 U10434 ( .A(n14238), .ZN(n8765) );
  OR2_X1 U10435 ( .A1(n14235), .A2(n8765), .ZN(n8766) );
  NAND2_X1 U10436 ( .A1(n8767), .A2(n8766), .ZN(n10965) );
  INV_X1 U10437 ( .A(n10965), .ZN(n8771) );
  INV_X1 U10438 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U10439 ( .A1(n14904), .A2(n15138), .ZN(n8770) );
  INV_X1 U10440 ( .A(n14242), .ZN(n8768) );
  NAND4_X1 U10441 ( .A1(n10964), .A2(n15140), .A3(n8771), .A4(n15139), .ZN(
        n8844) );
  INV_X1 U10442 ( .A(n10963), .ZN(n8773) );
  NAND2_X1 U10443 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8774) );
  NAND2_X1 U10444 ( .A1(n8774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8775) );
  OAI21_X1 U10445 ( .B1(n8776), .B2(P2_IR_REG_20__SCAN_IN), .A(n8775), .ZN(
        n8780) );
  NAND2_X1 U10446 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8777) );
  OR2_X1 U10447 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  OAI211_X1 U10448 ( .C1(n8781), .C2(P2_IR_REG_19__SCAN_IN), .A(n8780), .B(
        n8779), .ZN(n8782) );
  NAND2_X1 U10449 ( .A1(n13780), .A2(n13779), .ZN(n11253) );
  AND2_X1 U10450 ( .A1(n10707), .A2(n11253), .ZN(n8785) );
  NAND2_X1 U10451 ( .A1(n13521), .A2(n13534), .ZN(n11319) );
  NAND2_X1 U10452 ( .A1(n11320), .A2(n11319), .ZN(n8786) );
  NAND2_X1 U10453 ( .A1(n8786), .A2(n13747), .ZN(n11006) );
  NAND2_X1 U10454 ( .A1(n11006), .A2(n11007), .ZN(n8788) );
  INV_X1 U10455 ( .A(n13749), .ZN(n8787) );
  NAND2_X1 U10456 ( .A1(n8788), .A2(n8787), .ZN(n11005) );
  NAND2_X1 U10457 ( .A1(n12511), .A2(n13544), .ZN(n11335) );
  NAND2_X1 U10458 ( .A1(n11005), .A2(n11335), .ZN(n8790) );
  INV_X1 U10459 ( .A(n13750), .ZN(n8789) );
  NAND2_X1 U10460 ( .A1(n13554), .A2(n11118), .ZN(n8791) );
  OR2_X1 U10461 ( .A1(n13559), .A2(n12507), .ZN(n8792) );
  NAND2_X1 U10462 ( .A1(n11100), .A2(n13754), .ZN(n8794) );
  NAND2_X1 U10463 ( .A1(n13567), .A2(n11114), .ZN(n8793) );
  NAND2_X1 U10464 ( .A1(n8794), .A2(n8793), .ZN(n11447) );
  INV_X1 U10465 ( .A(n13809), .ZN(n11420) );
  OR2_X1 U10466 ( .A1(n13576), .A2(n11420), .ZN(n8795) );
  NAND2_X1 U10467 ( .A1(n11447), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U10468 ( .A1(n13576), .A2(n11420), .ZN(n8796) );
  NAND2_X1 U10469 ( .A1(n13580), .A2(n12488), .ZN(n8798) );
  INV_X1 U10470 ( .A(n13807), .ZN(n11421) );
  OR2_X1 U10471 ( .A1(n13587), .A2(n11421), .ZN(n8800) );
  NAND2_X1 U10472 ( .A1(n11462), .A2(n8800), .ZN(n11615) );
  INV_X1 U10473 ( .A(n13759), .ZN(n11614) );
  OR2_X1 U10474 ( .A1(n13591), .A2(n11823), .ZN(n8801) );
  NAND2_X1 U10475 ( .A1(n13600), .A2(n8803), .ZN(n8804) );
  INV_X1 U10476 ( .A(n13804), .ZN(n11824) );
  OR2_X1 U10477 ( .A1(n13603), .A2(n11824), .ZN(n8806) );
  INV_X1 U10478 ( .A(n13803), .ZN(n8807) );
  NAND2_X1 U10479 ( .A1(n13612), .A2(n8807), .ZN(n8808) );
  NAND2_X1 U10480 ( .A1(n12054), .A2(n15862), .ZN(n8809) );
  NAND2_X1 U10481 ( .A1(n8809), .A2(n13802), .ZN(n8812) );
  INV_X1 U10482 ( .A(n12054), .ZN(n8810) );
  NAND2_X1 U10483 ( .A1(n8810), .A2(n7575), .ZN(n8811) );
  NAND2_X1 U10484 ( .A1(n8812), .A2(n8811), .ZN(n12185) );
  OR2_X1 U10485 ( .A1(n13622), .A2(n8813), .ZN(n8814) );
  INV_X1 U10486 ( .A(n13626), .ZN(n14168) );
  NAND2_X1 U10487 ( .A1(n12371), .A2(n13768), .ZN(n8816) );
  INV_X1 U10488 ( .A(n14070), .ZN(n13501) );
  OR2_X1 U10489 ( .A1(n13635), .A2(n13501), .ZN(n8815) );
  INV_X1 U10490 ( .A(n13799), .ZN(n14056) );
  INV_X1 U10491 ( .A(n14072), .ZN(n14031) );
  INV_X1 U10492 ( .A(n13798), .ZN(n14058) );
  XNOR2_X1 U10493 ( .A(n14146), .B(n14058), .ZN(n14028) );
  INV_X1 U10494 ( .A(n13797), .ZN(n14032) );
  OR2_X1 U10495 ( .A1(n14141), .A2(n14032), .ZN(n8819) );
  INV_X1 U10496 ( .A(n13796), .ZN(n13485) );
  OR2_X1 U10497 ( .A1(n14010), .A2(n13485), .ZN(n8820) );
  NAND2_X1 U10498 ( .A1(n13991), .A2(n13990), .ZN(n13989) );
  INV_X1 U10499 ( .A(n13795), .ZN(n13667) );
  OR2_X1 U10500 ( .A1(n13994), .A2(n13667), .ZN(n8821) );
  AND2_X1 U10501 ( .A1(n13966), .A2(n13950), .ZN(n8822) );
  NAND2_X1 U10502 ( .A1(n8823), .A2(n13930), .ZN(n13935) );
  OR2_X1 U10503 ( .A1(n13944), .A2(n13411), .ZN(n8824) );
  INV_X1 U10504 ( .A(n13693), .ZN(n13791) );
  OR2_X1 U10505 ( .A1(n14187), .A2(n13791), .ZN(n8825) );
  INV_X1 U10506 ( .A(n13901), .ZN(n8827) );
  INV_X1 U10507 ( .A(n13900), .ZN(n8826) );
  NAND2_X1 U10508 ( .A1(n8827), .A2(n8826), .ZN(n13903) );
  NAND2_X1 U10509 ( .A1(n13903), .A2(n8828), .ZN(n8830) );
  INV_X1 U10510 ( .A(n13774), .ZN(n8829) );
  INV_X1 U10511 ( .A(n13736), .ZN(n13746) );
  NAND2_X1 U10512 ( .A1(n13746), .A2(n13779), .ZN(n8831) );
  OAI21_X2 U10513 ( .B1(n7193), .B2(n13776), .A(n8831), .ZN(n14074) );
  INV_X1 U10514 ( .A(n10341), .ZN(n8833) );
  NAND2_X1 U10515 ( .A1(n13790), .A2(n14069), .ZN(n8840) );
  INV_X1 U10516 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U10517 ( .A1(n8834), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U10518 ( .A1(n8709), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8835) );
  OAI211_X1 U10519 ( .C1(n8572), .C2(n14178), .A(n8836), .B(n8835), .ZN(n13788) );
  NOR2_X1 U10520 ( .A1(n14231), .A2(n8837), .ZN(n8838) );
  NOR2_X1 U10521 ( .A1(n14057), .A2(n8838), .ZN(n13885) );
  NAND2_X1 U10522 ( .A1(n13788), .A2(n13885), .ZN(n8839) );
  INV_X1 U10523 ( .A(n13600), .ZN(n15822) );
  INV_X1 U10524 ( .A(n13580), .ZN(n15754) );
  NAND2_X1 U10525 ( .A1(n13522), .A2(n13529), .ZN(n11325) );
  NOR2_X2 U10526 ( .A1(n11327), .A2(n13544), .ZN(n11343) );
  INV_X1 U10527 ( .A(n13554), .ZN(n15637) );
  NAND2_X1 U10528 ( .A1(n11343), .A2(n15637), .ZN(n11342) );
  NOR2_X2 U10529 ( .A1(n7234), .A2(n13567), .ZN(n11453) );
  INV_X1 U10530 ( .A(n13576), .ZN(n12487) );
  NAND2_X1 U10531 ( .A1(n15754), .A2(n11454), .ZN(n11467) );
  NOR2_X2 U10532 ( .A1(n13591), .A2(n11619), .ZN(n11818) );
  NAND2_X1 U10533 ( .A1(n15822), .A2(n11818), .ZN(n11819) );
  NAND2_X1 U10534 ( .A1(n14168), .A2(n12386), .ZN(n12389) );
  NOR2_X2 U10535 ( .A1(n14155), .A2(n14077), .ZN(n14075) );
  NAND2_X1 U10536 ( .A1(n14213), .A2(n14075), .ZN(n14045) );
  NOR2_X2 U10537 ( .A1(n13996), .A2(n14126), .ZN(n13978) );
  INV_X1 U10538 ( .A(n13895), .ZN(n8843) );
  AOI211_X1 U10539 ( .C1(n14096), .C2(n8843), .A(n14076), .B(n13889), .ZN(
        n14095) );
  AND2_X1 U10540 ( .A1(n10986), .A2(n13746), .ZN(n10703) );
  INV_X1 U10541 ( .A(n10703), .ZN(n8845) );
  INV_X1 U10542 ( .A(n8846), .ZN(n8847) );
  INV_X1 U10543 ( .A(n13959), .ZN(n15816) );
  AOI22_X1 U10544 ( .A1(n8847), .A2(n15816), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13980), .ZN(n8848) );
  OAI21_X1 U10545 ( .B1(n13688), .B2(n15821), .A(n8848), .ZN(n8849) );
  AOI21_X1 U10546 ( .B1(n14095), .B2(n15814), .A(n8849), .ZN(n8850) );
  INV_X2 U10547 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U10548 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8855) );
  NOR2_X2 U10549 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n8854) );
  NAND4_X1 U10550 ( .A1(n8855), .A2(n8854), .A3(n9108), .A4(n9030), .ZN(n8858)
         );
  NAND4_X1 U10551 ( .A1(n9094), .A2(n9127), .A3(n9059), .A4(n8856), .ZN(n8857)
         );
  NOR2_X2 U10552 ( .A1(n8858), .A2(n8857), .ZN(n9181) );
  NAND3_X1 U10553 ( .A1(n8862), .A2(n8893), .A3(n9478), .ZN(n8865) );
  NAND2_X1 U10554 ( .A1(n9479), .A2(n8863), .ZN(n8864) );
  NAND2_X1 U10555 ( .A1(n8870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8869) );
  INV_X1 U10556 ( .A(n8870), .ZN(n8872) );
  NAND2_X2 U10557 ( .A1(n8882), .A2(n8877), .ZN(n9015) );
  NAND2_X1 U10558 ( .A1(n9407), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10559 ( .A1(n9408), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8885) );
  AND2_X2 U10560 ( .A1(n8876), .A2(n14881), .ZN(n8929) );
  NAND2_X1 U10561 ( .A1(n8993), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U10562 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n8878) );
  NOR2_X1 U10563 ( .A1(n9035), .A2(n8878), .ZN(n9051) );
  NAND2_X1 U10564 ( .A1(n9051), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9070) );
  INV_X1 U10565 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9069) );
  AND2_X1 U10566 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8879) );
  NAND2_X1 U10567 ( .A1(n9135), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9159) );
  INV_X1 U10568 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9158) );
  INV_X1 U10569 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U10570 ( .A1(n9210), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9233) );
  INV_X1 U10571 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9232) );
  INV_X1 U10572 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U10573 ( .A1(n9260), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U10574 ( .A1(n9306), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9326) );
  INV_X1 U10575 ( .A(n9326), .ZN(n9307) );
  NAND2_X1 U10576 ( .A1(n9307), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9343) );
  INV_X1 U10577 ( .A(n9343), .ZN(n9325) );
  NAND2_X1 U10578 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9325), .ZN(n9345) );
  INV_X1 U10579 ( .A(n9345), .ZN(n8880) );
  NAND2_X1 U10580 ( .A1(n8880), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9409) );
  INV_X1 U10581 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U10582 ( .A1(n9345), .A2(n14250), .ZN(n8881) );
  NAND2_X1 U10583 ( .A1(n9410), .A2(n14603), .ZN(n8884) );
  NAND2_X1 U10584 ( .A1(n9411), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8883) );
  NAND4_X1 U10585 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n14356) );
  INV_X1 U10586 ( .A(n14356), .ZN(n14334) );
  INV_X1 U10587 ( .A(n8887), .ZN(n8890) );
  NAND2_X1 U10588 ( .A1(n8890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8888) );
  MUX2_X2 U10589 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8888), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8889) );
  NAND2_X1 U10590 ( .A1(n14230), .A2(n9416), .ZN(n8892) );
  NAND2_X1 U10591 ( .A1(n7206), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8891) );
  INV_X1 U10592 ( .A(n8901), .ZN(n8894) );
  INV_X1 U10593 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U10594 ( .A1(n8896), .A2(n8895), .ZN(n9390) );
  NAND2_X1 U10595 ( .A1(n8897), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U10596 ( .A1(n8899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U10597 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8900), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8902) );
  INV_X1 U10598 ( .A(n11220), .ZN(n10910) );
  NAND2_X1 U10599 ( .A1(n11229), .A2(n15537), .ZN(n11223) );
  NAND2_X1 U10600 ( .A1(n8908), .A2(n8905), .ZN(n9392) );
  NAND2_X1 U10601 ( .A1(n8906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8907) );
  INV_X1 U10602 ( .A(n15536), .ZN(n11222) );
  NAND2_X1 U10603 ( .A1(n9387), .A2(n11222), .ZN(n11230) );
  NAND2_X1 U10604 ( .A1(n8908), .A2(n11222), .ZN(n8909) );
  AND2_X4 U10605 ( .A1(n9380), .A2(n8909), .ZN(n8984) );
  MUX2_X1 U10606 ( .A(n14334), .B(n14804), .S(n9419), .Z(n9356) );
  INV_X1 U10607 ( .A(n9356), .ZN(n9357) );
  NAND2_X1 U10608 ( .A1(n8947), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8913) );
  INV_X1 U10609 ( .A(n8919), .ZN(n8946) );
  NAND2_X1 U10610 ( .A1(n8946), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U10611 ( .A1(n9103), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8911) );
  INV_X1 U10612 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U10613 ( .A1(n8929), .A2(n11363), .ZN(n8910) );
  INV_X1 U10614 ( .A(n14373), .ZN(n11239) );
  NAND2_X1 U10615 ( .A1(n7207), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8918) );
  OR2_X1 U10616 ( .A1(n8915), .A2(n8979), .ZN(n8916) );
  XNOR2_X1 U10617 ( .A(n8916), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U10618 ( .A1(n7200), .A2(n14413), .ZN(n8917) );
  AOI21_X1 U10619 ( .B1(n11239), .B2(n8984), .A(n15620), .ZN(n8973) );
  AOI21_X1 U10620 ( .B1(n14373), .B2(n9268), .A(n11364), .ZN(n8972) );
  INV_X1 U10621 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U10622 ( .A1(n8929), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8923) );
  INV_X1 U10623 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U10624 ( .A1(n9103), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U10625 ( .A1(n8953), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U10626 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8925) );
  XNOR2_X1 U10627 ( .A(n8925), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14386) );
  INV_X1 U10628 ( .A(n14386), .ZN(n8926) );
  INV_X2 U10629 ( .A(n11503), .ZN(n15565) );
  NAND2_X1 U10630 ( .A1(n15529), .A2(n15565), .ZN(n11225) );
  INV_X1 U10631 ( .A(n11225), .ZN(n8945) );
  AOI21_X1 U10632 ( .B1(n15529), .B2(n9268), .A(n15565), .ZN(n8944) );
  NAND2_X1 U10633 ( .A1(n8929), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U10634 ( .A1(n9103), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8930) );
  AND2_X2 U10635 ( .A1(n8931), .A2(n8930), .ZN(n8934) );
  NAND2_X1 U10636 ( .A1(n8946), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U10637 ( .A1(n8947), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U10638 ( .A1(n10397), .A2(SI_0_), .ZN(n8935) );
  XNOR2_X1 U10639 ( .A(n8935), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14900) );
  OAI21_X2 U10640 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n15527) );
  NOR2_X2 U10641 ( .A1(n14375), .A2(n8941), .ZN(n11233) );
  INV_X1 U10642 ( .A(n11233), .ZN(n8940) );
  NAND3_X1 U10643 ( .A1(n8940), .A2(n8984), .A3(n11234), .ZN(n8943) );
  NAND2_X1 U10644 ( .A1(n14375), .A2(n8941), .ZN(n9434) );
  OAI211_X1 U10645 ( .C1(n11233), .C2(n11219), .A(n9434), .B(n9268), .ZN(n8942) );
  OAI211_X1 U10646 ( .C1(n8945), .C2(n8944), .A(n8943), .B(n8942), .ZN(n8965)
         );
  NAND2_X1 U10647 ( .A1(n8947), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U10648 ( .A1(n9103), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U10649 ( .A1(n8929), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U10650 ( .A1(n7206), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8957) );
  OR2_X1 U10651 ( .A1(n8954), .A2(n8979), .ZN(n8955) );
  XNOR2_X1 U10652 ( .A(n8955), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U10653 ( .A1(n7199), .A2(n14397), .ZN(n8956) );
  MUX2_X1 U10654 ( .A(n14374), .B(n11516), .S(n8984), .Z(n8966) );
  NAND2_X1 U10655 ( .A1(n8960), .A2(n8966), .ZN(n8964) );
  NAND3_X1 U10656 ( .A1(n8965), .A2(n8964), .A3(n8963), .ZN(n8970) );
  INV_X1 U10657 ( .A(n8966), .ZN(n8968) );
  NAND2_X1 U10658 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  NAND2_X1 U10659 ( .A1(n9407), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10660 ( .A1(n9408), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8977) );
  NOR2_X1 U10661 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8974) );
  NOR2_X1 U10662 ( .A1(n8993), .A2(n8974), .ZN(n11442) );
  NAND2_X1 U10663 ( .A1(n9410), .A2(n11442), .ZN(n8976) );
  NAND2_X1 U10664 ( .A1(n9103), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8975) );
  NAND4_X1 U10665 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n14372) );
  OR2_X1 U10666 ( .A1(n8980), .A2(n8979), .ZN(n8982) );
  XNOR2_X1 U10667 ( .A(n8982), .B(n8981), .ZN(n10461) );
  NAND2_X1 U10668 ( .A1(n7206), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U10669 ( .A(n14372), .B(n11709), .S(n8984), .Z(n8988) );
  NAND2_X1 U10670 ( .A1(n8987), .A2(n8988), .ZN(n8986) );
  MUX2_X1 U10671 ( .A(n14372), .B(n11709), .S(n9268), .Z(n8985) );
  NAND2_X1 U10672 ( .A1(n8986), .A2(n8985), .ZN(n8992) );
  INV_X1 U10673 ( .A(n8987), .ZN(n8990) );
  INV_X1 U10674 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U10675 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NAND2_X1 U10676 ( .A1(n8992), .A2(n8991), .ZN(n9006) );
  NAND2_X1 U10677 ( .A1(n9408), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U10678 ( .A1(n9407), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8996) );
  OAI21_X1 U10679 ( .B1(n8993), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9035), .ZN(
        n11608) );
  INV_X1 U10680 ( .A(n11608), .ZN(n15666) );
  NAND2_X1 U10681 ( .A1(n9410), .A2(n15666), .ZN(n8995) );
  NAND2_X1 U10682 ( .A1(n9103), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U10683 ( .A1(n10426), .A2(n9416), .ZN(n9003) );
  NAND2_X1 U10684 ( .A1(n8999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9000) );
  MUX2_X1 U10685 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9000), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9001) );
  OR2_X1 U10686 ( .A1(n8999), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9029) );
  AND2_X1 U10687 ( .A1(n9001), .A2(n9029), .ZN(n10523) );
  AOI22_X1 U10688 ( .A1(n9249), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7200), .B2(
        n10523), .ZN(n9002) );
  NAND2_X1 U10689 ( .A1(n9003), .A2(n9002), .ZN(n11716) );
  MUX2_X1 U10690 ( .A(n14371), .B(n11716), .S(n9419), .Z(n9007) );
  NAND2_X1 U10691 ( .A1(n9006), .A2(n9007), .ZN(n9005) );
  MUX2_X1 U10692 ( .A(n14371), .B(n11716), .S(n8984), .Z(n9004) );
  NAND2_X1 U10693 ( .A1(n9005), .A2(n9004), .ZN(n9011) );
  INV_X1 U10694 ( .A(n9006), .ZN(n9009) );
  INV_X1 U10695 ( .A(n9007), .ZN(n9008) );
  NAND2_X1 U10696 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U10697 ( .A1(n9011), .A2(n9010), .ZN(n9023) );
  OR2_X1 U10698 ( .A1(n10432), .A2(n7203), .ZN(n9014) );
  NAND2_X1 U10699 ( .A1(n9029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9012) );
  XNOR2_X1 U10700 ( .A(n9012), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14430) );
  AOI22_X1 U10701 ( .A1(n9249), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7200), .B2(
        n14430), .ZN(n9013) );
  NAND2_X1 U10702 ( .A1(n9014), .A2(n9013), .ZN(n11780) );
  XNOR2_X1 U10703 ( .A(n9035), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U10704 ( .A1(n9410), .A2(n11779), .ZN(n9020) );
  NAND2_X1 U10705 ( .A1(n9411), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9019) );
  INV_X1 U10706 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9016) );
  OR2_X1 U10707 ( .A1(n9015), .A2(n9016), .ZN(n9018) );
  INV_X1 U10708 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10524) );
  OR2_X1 U10709 ( .A1(n7195), .A2(n10524), .ZN(n9017) );
  MUX2_X1 U10710 ( .A(n11780), .B(n14370), .S(n9419), .Z(n9024) );
  NAND2_X1 U10711 ( .A1(n9023), .A2(n9024), .ZN(n9022) );
  MUX2_X1 U10712 ( .A(n11780), .B(n14370), .S(n8984), .Z(n9021) );
  NAND2_X1 U10713 ( .A1(n9022), .A2(n9021), .ZN(n9028) );
  INV_X1 U10714 ( .A(n9023), .ZN(n9026) );
  INV_X1 U10715 ( .A(n9024), .ZN(n9025) );
  NAND2_X1 U10716 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  NAND2_X1 U10717 ( .A1(n9028), .A2(n9027), .ZN(n9045) );
  OR2_X1 U10718 ( .A1(n10435), .A2(n7203), .ZN(n9034) );
  INV_X1 U10719 ( .A(n9029), .ZN(n9031) );
  NAND2_X1 U10720 ( .A1(n9031), .A2(n9030), .ZN(n9058) );
  NAND2_X1 U10721 ( .A1(n9058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9032) );
  XNOR2_X1 U10722 ( .A(n9032), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U10723 ( .A1(n9249), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7200), .B2(
        n14449), .ZN(n9033) );
  INV_X1 U10724 ( .A(n9035), .ZN(n9036) );
  AOI21_X1 U10725 ( .B1(n9036), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n9037) );
  NOR2_X1 U10726 ( .A1(n9037), .A2(n9051), .ZN(n15720) );
  NAND2_X1 U10727 ( .A1(n9410), .A2(n15720), .ZN(n9042) );
  NAND2_X1 U10728 ( .A1(n9411), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9041) );
  INV_X1 U10729 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9038) );
  OR2_X1 U10730 ( .A1(n9015), .A2(n9038), .ZN(n9040) );
  INV_X1 U10731 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10527) );
  OR2_X1 U10732 ( .A1(n7195), .A2(n10527), .ZN(n9039) );
  INV_X1 U10733 ( .A(n11764), .ZN(n14369) );
  MUX2_X1 U10734 ( .A(n11763), .B(n14369), .S(n8984), .Z(n9046) );
  NAND2_X1 U10735 ( .A1(n9045), .A2(n9046), .ZN(n9044) );
  MUX2_X1 U10736 ( .A(n11763), .B(n14369), .S(n9419), .Z(n9043) );
  NAND2_X1 U10737 ( .A1(n9044), .A2(n9043), .ZN(n9050) );
  INV_X1 U10738 ( .A(n9045), .ZN(n9048) );
  INV_X1 U10739 ( .A(n9046), .ZN(n9047) );
  NAND2_X1 U10740 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NAND2_X1 U10741 ( .A1(n9103), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9057) );
  OR2_X1 U10742 ( .A1(n9051), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9052) );
  AND2_X1 U10743 ( .A1(n9070), .A2(n9052), .ZN(n11869) );
  NAND2_X1 U10744 ( .A1(n9410), .A2(n11869), .ZN(n9056) );
  INV_X1 U10745 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10530) );
  OR2_X1 U10746 ( .A1(n7195), .A2(n10530), .ZN(n9055) );
  INV_X1 U10747 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9053) );
  OR2_X1 U10748 ( .A1(n9015), .A2(n9053), .ZN(n9054) );
  INV_X1 U10749 ( .A(n12044), .ZN(n14368) );
  NAND2_X1 U10750 ( .A1(n10450), .A2(n9416), .ZN(n9065) );
  INV_X1 U10751 ( .A(n9058), .ZN(n9060) );
  NAND2_X1 U10752 ( .A1(n9060), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U10753 ( .A1(n9062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9061) );
  MUX2_X1 U10754 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9061), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9063) );
  AND2_X1 U10755 ( .A1(n9063), .A2(n9076), .ZN(n10554) );
  AOI22_X1 U10756 ( .A1(n9249), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7200), .B2(
        n10554), .ZN(n9064) );
  NAND2_X2 U10757 ( .A1(n9065), .A2(n9064), .ZN(n15742) );
  MUX2_X1 U10758 ( .A(n14368), .B(n15742), .S(n8984), .Z(n9067) );
  MUX2_X1 U10759 ( .A(n14368), .B(n15742), .S(n9419), .Z(n9066) );
  INV_X1 U10760 ( .A(n9067), .ZN(n9068) );
  NAND2_X1 U10761 ( .A1(n9407), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U10762 ( .A1(n9408), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U10763 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  AND2_X1 U10764 ( .A1(n9088), .A2(n9071), .ZN(n15780) );
  NAND2_X1 U10765 ( .A1(n9410), .A2(n15780), .ZN(n9073) );
  NAND2_X1 U10766 ( .A1(n9103), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9072) );
  NAND4_X1 U10767 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n14367) );
  OR2_X1 U10768 ( .A1(n10455), .A2(n7203), .ZN(n9078) );
  NAND2_X1 U10769 ( .A1(n9076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9095) );
  XNOR2_X1 U10770 ( .A(n9095), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U10771 ( .A1(n9249), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7200), .B2(
        n14464), .ZN(n9077) );
  MUX2_X1 U10772 ( .A(n14367), .B(n15781), .S(n9419), .Z(n9082) );
  MUX2_X1 U10773 ( .A(n14367), .B(n15781), .S(n8984), .Z(n9079) );
  NAND2_X1 U10774 ( .A1(n9080), .A2(n9079), .ZN(n9086) );
  INV_X1 U10775 ( .A(n9081), .ZN(n9084) );
  INV_X1 U10776 ( .A(n9082), .ZN(n9083) );
  NAND2_X1 U10777 ( .A1(n9084), .A2(n9083), .ZN(n9085) );
  NAND2_X1 U10778 ( .A1(n9086), .A2(n9085), .ZN(n9100) );
  NAND2_X1 U10779 ( .A1(n9408), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10780 ( .A1(n9103), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9092) );
  AND2_X1 U10781 ( .A1(n9088), .A2(n9087), .ZN(n9089) );
  NOR2_X1 U10782 ( .A1(n9119), .A2(n9089), .ZN(n12118) );
  NAND2_X1 U10783 ( .A1(n9410), .A2(n12118), .ZN(n9091) );
  NAND2_X1 U10784 ( .A1(n9407), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9090) );
  NAND4_X1 U10785 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n14366) );
  OR2_X1 U10786 ( .A1(n10460), .A2(n7203), .ZN(n9098) );
  NAND2_X1 U10787 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  NAND2_X1 U10788 ( .A1(n9096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9109) );
  XNOR2_X1 U10789 ( .A(n9109), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U10790 ( .A1(n9249), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7200), 
        .B2(n14479), .ZN(n9097) );
  MUX2_X1 U10791 ( .A(n14366), .B(n12119), .S(n8984), .Z(n9101) );
  MUX2_X1 U10792 ( .A(n14366), .B(n12119), .S(n9419), .Z(n9099) );
  NAND2_X1 U10793 ( .A1(n9407), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U10794 ( .A1(n9408), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9106) );
  INV_X1 U10795 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U10796 ( .A(n9119), .B(n9102), .ZN(n12230) );
  NAND2_X1 U10797 ( .A1(n9410), .A2(n12230), .ZN(n9105) );
  NAND2_X1 U10798 ( .A1(n9103), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9104) );
  NAND4_X1 U10799 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n14365) );
  NAND2_X1 U10800 ( .A1(n10512), .A2(n9416), .ZN(n9112) );
  NAND2_X1 U10801 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U10802 ( .A1(n9110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9128) );
  XNOR2_X1 U10803 ( .A(n9128), .B(P1_IR_REG_11__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U10804 ( .A1(n9249), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n14496), 
        .B2(n7200), .ZN(n9111) );
  MUX2_X1 U10805 ( .A(n14365), .B(n12234), .S(n9419), .Z(n9116) );
  MUX2_X1 U10806 ( .A(n14365), .B(n12234), .S(n8984), .Z(n9113) );
  NAND2_X1 U10807 ( .A1(n9114), .A2(n9113), .ZN(n9118) );
  NAND2_X1 U10808 ( .A1(n9118), .A2(n9117), .ZN(n9133) );
  AOI21_X1 U10809 ( .B1(n9119), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n9120) );
  NOR2_X1 U10810 ( .A1(n9135), .A2(n9120), .ZN(n12290) );
  NAND2_X1 U10811 ( .A1(n9410), .A2(n12290), .ZN(n9126) );
  NAND2_X1 U10812 ( .A1(n9411), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9125) );
  INV_X1 U10813 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9121) );
  OR2_X1 U10814 ( .A1(n7195), .A2(n9121), .ZN(n9124) );
  INV_X1 U10815 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9122) );
  OR2_X1 U10816 ( .A1(n9015), .A2(n9122), .ZN(n9123) );
  NAND2_X1 U10817 ( .A1(n10582), .A2(n9416), .ZN(n9131) );
  NAND2_X1 U10818 ( .A1(n9128), .A2(n9127), .ZN(n9129) );
  NAND2_X1 U10819 ( .A1(n9129), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9143) );
  XNOR2_X1 U10820 ( .A(n9143), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U10821 ( .A1(n10734), .A2(n7200), .B1(n7206), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9130) );
  MUX2_X1 U10822 ( .A(n14364), .B(n12281), .S(n8984), .Z(n9134) );
  MUX2_X1 U10823 ( .A(n14364), .B(n12281), .S(n9419), .Z(n9132) );
  OR2_X1 U10824 ( .A1(n9135), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9136) );
  AND2_X1 U10825 ( .A1(n9159), .A2(n9136), .ZN(n12253) );
  NAND2_X1 U10826 ( .A1(n9410), .A2(n12253), .ZN(n9141) );
  NAND2_X1 U10827 ( .A1(n9411), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9140) );
  INV_X1 U10828 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9137) );
  OR2_X1 U10829 ( .A1(n9015), .A2(n9137), .ZN(n9139) );
  INV_X1 U10830 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12210) );
  OR2_X1 U10831 ( .A1(n7195), .A2(n12210), .ZN(n9138) );
  INV_X1 U10832 ( .A(n12409), .ZN(n14363) );
  OR2_X1 U10833 ( .A1(n10692), .A2(n7203), .ZN(n9149) );
  INV_X1 U10834 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U10835 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  NAND2_X1 U10836 ( .A1(n9144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9146) );
  INV_X1 U10837 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U10838 ( .A1(n9146), .A2(n9145), .ZN(n9167) );
  OR2_X1 U10839 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  AOI22_X1 U10840 ( .A1(n11021), .A2(n7200), .B1(n7207), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9148) );
  MUX2_X1 U10841 ( .A(n14363), .B(n12408), .S(n9419), .Z(n9153) );
  MUX2_X1 U10842 ( .A(n14363), .B(n12408), .S(n8984), .Z(n9150) );
  NAND2_X1 U10843 ( .A1(n9151), .A2(n9150), .ZN(n9157) );
  INV_X1 U10844 ( .A(n9152), .ZN(n9155) );
  INV_X1 U10845 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U10846 ( .A1(n9155), .A2(n9154), .ZN(n9156) );
  NAND2_X1 U10847 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  AND2_X1 U10848 ( .A1(n9175), .A2(n9160), .ZN(n14261) );
  NAND2_X1 U10849 ( .A1(n9410), .A2(n14261), .ZN(n9166) );
  NAND2_X1 U10850 ( .A1(n9411), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9165) );
  INV_X1 U10851 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9161) );
  OR2_X1 U10852 ( .A1(n9015), .A2(n9161), .ZN(n9164) );
  INV_X1 U10853 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9162) );
  OR2_X1 U10854 ( .A1(n7195), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U10855 ( .A1(n10980), .A2(n9416), .ZN(n9170) );
  NAND2_X1 U10856 ( .A1(n9167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9168) );
  XNOR2_X1 U10857 ( .A(n9168), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U10858 ( .A1(n11300), .A2(n7200), .B1(n7207), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9169) );
  MUX2_X1 U10859 ( .A(n14362), .B(n12606), .S(n8984), .Z(n9172) );
  MUX2_X1 U10860 ( .A(n14362), .B(n12606), .S(n9419), .Z(n9171) );
  INV_X1 U10861 ( .A(n9172), .ZN(n9173) );
  NAND2_X1 U10862 ( .A1(n9407), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U10863 ( .A1(n9408), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U10864 ( .A1(n9175), .A2(n9174), .ZN(n9176) );
  AND2_X1 U10865 ( .A1(n9201), .A2(n9176), .ZN(n14351) );
  NAND2_X1 U10866 ( .A1(n9410), .A2(n14351), .ZN(n9178) );
  NAND2_X1 U10867 ( .A1(n9411), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9177) );
  NAND4_X1 U10868 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(n14768) );
  NAND2_X1 U10869 ( .A1(n11167), .A2(n9416), .ZN(n9186) );
  BUF_X1 U10870 ( .A(n9181), .Z(n9182) );
  INV_X1 U10871 ( .A(n9182), .ZN(n9183) );
  NOR2_X1 U10872 ( .A1(n8999), .A2(n9183), .ZN(n9196) );
  OR2_X1 U10873 ( .A1(n9196), .A2(n8979), .ZN(n9184) );
  XNOR2_X1 U10874 ( .A(n9184), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U10875 ( .A1(n9249), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7200), 
        .B2(n11305), .ZN(n9185) );
  MUX2_X1 U10876 ( .A(n14768), .B(n12435), .S(n9419), .Z(n9190) );
  MUX2_X1 U10877 ( .A(n14768), .B(n12435), .S(n8984), .Z(n9187) );
  NAND2_X1 U10878 ( .A1(n9188), .A2(n9187), .ZN(n9194) );
  INV_X1 U10879 ( .A(n9189), .ZN(n9192) );
  INV_X1 U10880 ( .A(n9190), .ZN(n9191) );
  NAND2_X1 U10881 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  OR2_X1 U10882 ( .A1(n11401), .A2(n7203), .ZN(n9199) );
  INV_X1 U10883 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U10884 ( .A1(n9196), .A2(n9195), .ZN(n9216) );
  NAND2_X1 U10885 ( .A1(n9216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U10886 ( .A(n9197), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U10887 ( .A1(n9249), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7200), 
        .B2(n14505), .ZN(n9198) );
  INV_X2 U10888 ( .A(n14775), .ZN(n15888) );
  NAND2_X1 U10889 ( .A1(n9407), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U10890 ( .A1(n9408), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9205) );
  AND2_X1 U10891 ( .A1(n9201), .A2(n9200), .ZN(n9202) );
  NOR2_X1 U10892 ( .A1(n9210), .A2(n9202), .ZN(n14771) );
  NAND2_X1 U10893 ( .A1(n9410), .A2(n14771), .ZN(n9204) );
  NAND2_X1 U10894 ( .A1(n9411), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9203) );
  NAND4_X1 U10895 ( .A1(n9206), .A2(n9205), .A3(n9204), .A4(n9203), .ZN(n14361) );
  MUX2_X1 U10896 ( .A(n15888), .B(n14361), .S(n9419), .Z(n9208) );
  MUX2_X1 U10897 ( .A(n14361), .B(n15888), .S(n9419), .Z(n9207) );
  INV_X1 U10898 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U10899 ( .A1(n9407), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U10900 ( .A1(n9408), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U10901 ( .A1(n9411), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9213) );
  OR2_X1 U10902 ( .A1(n9210), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U10903 ( .A1(n9233), .A2(n9211), .ZN(n15908) );
  INV_X1 U10904 ( .A(n15908), .ZN(n15929) );
  NAND2_X1 U10905 ( .A1(n9410), .A2(n15929), .ZN(n9212) );
  NAND4_X1 U10906 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n14766) );
  NAND2_X1 U10907 ( .A1(n11674), .A2(n9416), .ZN(n9219) );
  OAI21_X1 U10908 ( .B1(n9216), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9217) );
  XNOR2_X1 U10909 ( .A(n9217), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14523) );
  AOI22_X1 U10910 ( .A1(n9249), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7200), 
        .B2(n14523), .ZN(n9218) );
  MUX2_X1 U10911 ( .A(n14766), .B(n15932), .S(n9419), .Z(n9223) );
  MUX2_X1 U10912 ( .A(n14766), .B(n15932), .S(n8984), .Z(n9220) );
  NAND2_X1 U10913 ( .A1(n9221), .A2(n9220), .ZN(n9227) );
  INV_X1 U10914 ( .A(n9222), .ZN(n9225) );
  INV_X1 U10915 ( .A(n9223), .ZN(n9224) );
  NAND2_X1 U10916 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND2_X1 U10917 ( .A1(n11906), .A2(n9416), .ZN(n9231) );
  NAND2_X1 U10918 ( .A1(n9228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9229) );
  XNOR2_X1 U10919 ( .A(n9229), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14542) );
  AOI22_X1 U10920 ( .A1(n9249), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7200), 
        .B2(n14542), .ZN(n9230) );
  NAND2_X1 U10921 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  NAND2_X1 U10922 ( .A1(n9245), .A2(n9234), .ZN(n15956) );
  INV_X1 U10923 ( .A(n15956), .ZN(n14753) );
  NAND2_X1 U10924 ( .A1(n14753), .A2(n9410), .ZN(n9240) );
  NAND2_X1 U10925 ( .A1(n9411), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9239) );
  INV_X1 U10926 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9235) );
  OR2_X1 U10927 ( .A1(n9015), .A2(n9235), .ZN(n9238) );
  INV_X1 U10928 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9236) );
  OR2_X1 U10929 ( .A1(n7195), .A2(n9236), .ZN(n9237) );
  MUX2_X1 U10930 ( .A(n15953), .B(n7876), .S(n9419), .Z(n9242) );
  MUX2_X1 U10931 ( .A(n15953), .B(n7876), .S(n8984), .Z(n9241) );
  INV_X1 U10932 ( .A(n9242), .ZN(n9243) );
  AND2_X1 U10933 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  OR2_X1 U10934 ( .A1(n9246), .A2(n9260), .ZN(n15968) );
  INV_X1 U10935 ( .A(n9410), .ZN(n9265) );
  AOI22_X1 U10936 ( .A1(n9407), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n9408), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U10937 ( .A1(n9411), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U10938 ( .C1(n15968), .C2(n9265), .A(n9248), .B(n9247), .ZN(n14744) );
  NAND2_X1 U10939 ( .A1(n12017), .A2(n9416), .ZN(n9251) );
  AOI22_X1 U10940 ( .A1(n9249), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15537), 
        .B2(n7200), .ZN(n9250) );
  MUX2_X1 U10941 ( .A(n14744), .B(n15964), .S(n9419), .Z(n9255) );
  MUX2_X1 U10942 ( .A(n14744), .B(n15964), .S(n8984), .Z(n9252) );
  NAND2_X1 U10943 ( .A1(n9253), .A2(n9252), .ZN(n9259) );
  INV_X1 U10944 ( .A(n9254), .ZN(n9257) );
  INV_X1 U10945 ( .A(n9255), .ZN(n9256) );
  NAND2_X1 U10946 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  OR2_X1 U10947 ( .A1(n9260), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U10948 ( .A1(n9262), .A2(n9261), .ZN(n14315) );
  AOI22_X1 U10949 ( .A1(n9407), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n9408), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U10950 ( .A1(n9411), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9263) );
  OAI211_X1 U10951 ( .C1(n14315), .C2(n9265), .A(n9264), .B(n9263), .ZN(n14730) );
  NAND2_X1 U10952 ( .A1(n12111), .A2(n9416), .ZN(n9267) );
  NAND2_X1 U10953 ( .A1(n7206), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9266) );
  MUX2_X1 U10954 ( .A(n14730), .B(n14848), .S(n8984), .Z(n9278) );
  MUX2_X1 U10955 ( .A(n14730), .B(n14848), .S(n9419), .Z(n9269) );
  NAND2_X1 U10956 ( .A1(n12216), .A2(n9416), .ZN(n9271) );
  NAND2_X1 U10957 ( .A1(n7207), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U10958 ( .A1(n9407), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U10959 ( .A1(n9408), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9276) );
  NOR2_X1 U10960 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n9272), .ZN(n9273) );
  NOR2_X1 U10961 ( .A1(n9281), .A2(n9273), .ZN(n14705) );
  NAND2_X1 U10962 ( .A1(n9410), .A2(n14705), .ZN(n9275) );
  NAND2_X1 U10963 ( .A1(n9411), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9274) );
  NAND4_X1 U10964 ( .A1(n9277), .A2(n9276), .A3(n9275), .A4(n9274), .ZN(n14360) );
  XNOR2_X1 U10965 ( .A(n14841), .B(n14360), .ZN(n14701) );
  NAND2_X1 U10966 ( .A1(n9279), .A2(n10397), .ZN(n9280) );
  XNOR2_X1 U10967 ( .A(n9280), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U10968 ( .A1(n9407), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U10969 ( .A1(n9408), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9285) );
  NOR2_X1 U10970 ( .A1(n9281), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9282) );
  NOR2_X1 U10971 ( .A1(n9295), .A2(n9282), .ZN(n14689) );
  NAND2_X1 U10972 ( .A1(n9410), .A2(n14689), .ZN(n9284) );
  NAND2_X1 U10973 ( .A1(n9411), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9283) );
  NAND4_X1 U10974 ( .A1(n9286), .A2(n9285), .A3(n9284), .A4(n9283), .ZN(n14662) );
  NAND2_X1 U10975 ( .A1(n14692), .A2(n14662), .ZN(n9292) );
  NAND2_X1 U10976 ( .A1(n12440), .A2(n9292), .ZN(n14683) );
  INV_X1 U10977 ( .A(n14683), .ZN(n14678) );
  AND2_X1 U10978 ( .A1(n14360), .A2(n9419), .ZN(n9289) );
  NAND2_X1 U10979 ( .A1(n14717), .A2(n8984), .ZN(n9287) );
  NAND2_X1 U10980 ( .A1(n14841), .A2(n9287), .ZN(n9288) );
  OAI21_X1 U10981 ( .B1(n14841), .B2(n9289), .A(n9288), .ZN(n9290) );
  NAND3_X1 U10982 ( .A1(n9291), .A2(n14678), .A3(n9290), .ZN(n9294) );
  MUX2_X1 U10983 ( .A(n9292), .B(n12440), .S(n9419), .Z(n9293) );
  NAND2_X1 U10984 ( .A1(n9411), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9301) );
  NOR2_X1 U10985 ( .A1(n9295), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9296) );
  NOR2_X1 U10986 ( .A1(n9306), .A2(n9296), .ZN(n14664) );
  NAND2_X1 U10987 ( .A1(n9410), .A2(n14664), .ZN(n9300) );
  INV_X1 U10988 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14668) );
  OR2_X1 U10989 ( .A1(n7195), .A2(n14668), .ZN(n9299) );
  INV_X1 U10990 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9297) );
  OR2_X1 U10991 ( .A1(n9015), .A2(n9297), .ZN(n9298) );
  NAND2_X1 U10992 ( .A1(n12256), .A2(n9416), .ZN(n9303) );
  NAND2_X1 U10993 ( .A1(n7206), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9302) );
  MUX2_X1 U10994 ( .A(n14359), .B(n14670), .S(n9419), .Z(n9305) );
  MUX2_X1 U10995 ( .A(n14359), .B(n14670), .S(n8984), .Z(n9304) );
  INV_X1 U10996 ( .A(n9306), .ZN(n9308) );
  INV_X1 U10997 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14308) );
  AOI21_X1 U10998 ( .B1(n9308), .B2(n14308), .A(n9307), .ZN(n14647) );
  NAND2_X1 U10999 ( .A1(n9410), .A2(n14647), .ZN(n9314) );
  NAND2_X1 U11000 ( .A1(n9411), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9313) );
  INV_X1 U11001 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9309) );
  OR2_X1 U11002 ( .A1(n7195), .A2(n9309), .ZN(n9312) );
  INV_X1 U11003 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9310) );
  OR2_X1 U11004 ( .A1(n9015), .A2(n9310), .ZN(n9311) );
  NAND2_X1 U11005 ( .A1(n14241), .A2(n9416), .ZN(n9316) );
  NAND2_X1 U11006 ( .A1(n7206), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9315) );
  MUX2_X1 U11007 ( .A(n14663), .B(n14651), .S(n8984), .Z(n9320) );
  NAND2_X1 U11008 ( .A1(n9319), .A2(n9320), .ZN(n9318) );
  MUX2_X1 U11009 ( .A(n14663), .B(n14651), .S(n9419), .Z(n9317) );
  NAND2_X1 U11010 ( .A1(n9318), .A2(n9317), .ZN(n9324) );
  INV_X1 U11011 ( .A(n9319), .ZN(n9322) );
  INV_X1 U11012 ( .A(n9320), .ZN(n9321) );
  NAND2_X1 U11013 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  NAND2_X1 U11014 ( .A1(n9324), .A2(n9323), .ZN(n9335) );
  NAND2_X1 U11015 ( .A1(n9408), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11016 ( .A1(n9407), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9329) );
  INV_X1 U11017 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14288) );
  AOI21_X1 U11018 ( .B1(n14288), .B2(n9326), .A(n9325), .ZN(n14635) );
  NAND2_X1 U11019 ( .A1(n9410), .A2(n14635), .ZN(n9328) );
  NAND2_X1 U11020 ( .A1(n9411), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9327) );
  NAND4_X1 U11021 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(n14358) );
  NAND2_X1 U11022 ( .A1(n14237), .A2(n9416), .ZN(n9332) );
  NAND2_X1 U11023 ( .A1(n7207), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9331) );
  MUX2_X1 U11024 ( .A(n14358), .B(n14817), .S(n9419), .Z(n9336) );
  NAND2_X1 U11025 ( .A1(n9335), .A2(n9336), .ZN(n9334) );
  MUX2_X1 U11026 ( .A(n14358), .B(n14817), .S(n8984), .Z(n9333) );
  NAND2_X1 U11027 ( .A1(n9334), .A2(n9333), .ZN(n9340) );
  INV_X1 U11028 ( .A(n9335), .ZN(n9338) );
  INV_X1 U11029 ( .A(n9336), .ZN(n9337) );
  NAND2_X1 U11030 ( .A1(n9338), .A2(n9337), .ZN(n9339) );
  NAND2_X1 U11031 ( .A1(n14233), .A2(n9416), .ZN(n9342) );
  NAND2_X1 U11032 ( .A1(n7207), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9341) );
  INV_X1 U11033 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U11034 ( .A1(n9344), .A2(n9343), .ZN(n9346) );
  AND2_X1 U11035 ( .A1(n9346), .A2(n9345), .ZN(n14616) );
  NAND2_X1 U11036 ( .A1(n9410), .A2(n14616), .ZN(n9352) );
  NAND2_X1 U11037 ( .A1(n9411), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9351) );
  INV_X1 U11038 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9347) );
  OR2_X1 U11039 ( .A1(n9015), .A2(n9347), .ZN(n9350) );
  INV_X1 U11040 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9348) );
  OR2_X1 U11041 ( .A1(n7195), .A2(n9348), .ZN(n9349) );
  MUX2_X1 U11042 ( .A(n14810), .B(n14357), .S(n9419), .Z(n9353) );
  MUX2_X1 U11043 ( .A(n14357), .B(n14810), .S(n9419), .Z(n9354) );
  MUX2_X1 U11044 ( .A(n14604), .B(n14356), .S(n9419), .Z(n9355) );
  INV_X1 U11045 ( .A(n9431), .ZN(n9421) );
  INV_X1 U11046 ( .A(SI_29_), .ZN(n15026) );
  NAND2_X1 U11047 ( .A1(n9360), .A2(n15026), .ZN(n9361) );
  MUX2_X1 U11048 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n10397), .Z(n9362) );
  NAND2_X1 U11049 ( .A1(n9362), .A2(SI_30_), .ZN(n9363) );
  OAI21_X1 U11050 ( .B1(SI_30_), .B2(n9362), .A(n9363), .ZN(n9374) );
  MUX2_X1 U11051 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10397), .Z(n9364) );
  XNOR2_X1 U11052 ( .A(n9364), .B(SI_31_), .ZN(n9365) );
  NAND2_X1 U11053 ( .A1(n13683), .A2(n9416), .ZN(n9368) );
  NAND2_X1 U11054 ( .A1(n7206), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9367) );
  INV_X1 U11055 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11056 ( .A1(n9411), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9372) );
  INV_X1 U11057 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9369) );
  OR2_X1 U11058 ( .A1(n7195), .A2(n9369), .ZN(n9371) );
  OAI211_X1 U11059 ( .C1(n9015), .C2(n9373), .A(n9372), .B(n9371), .ZN(n14562)
         );
  NAND2_X1 U11060 ( .A1(n9375), .A2(n9374), .ZN(n9376) );
  NAND2_X1 U11061 ( .A1(n13705), .A2(n9416), .ZN(n9379) );
  NAND2_X1 U11062 ( .A1(n7207), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9378) );
  INV_X1 U11063 ( .A(n9380), .ZN(n9384) );
  INV_X1 U11064 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11065 ( .A1(n9408), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11066 ( .A1(n9411), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9381) );
  OAI211_X1 U11067 ( .C1(n9015), .C2(n9383), .A(n9382), .B(n9381), .ZN(n14581)
         );
  OAI21_X1 U11068 ( .B1(n14562), .B2(n9384), .A(n14581), .ZN(n9385) );
  INV_X1 U11069 ( .A(n9385), .ZN(n9386) );
  MUX2_X1 U11070 ( .A(n14558), .B(n9386), .S(n9419), .Z(n9476) );
  INV_X1 U11071 ( .A(n9476), .ZN(n9510) );
  INV_X1 U11072 ( .A(n11229), .ZN(n14899) );
  AND2_X1 U11073 ( .A1(n11229), .A2(n15536), .ZN(n9388) );
  OR2_X1 U11074 ( .A1(n10359), .A2(n9388), .ZN(n9389) );
  NAND2_X1 U11075 ( .A1(n11219), .A2(n15537), .ZN(n15534) );
  NAND2_X1 U11076 ( .A1(n9389), .A2(n15534), .ZN(n9457) );
  NAND2_X1 U11077 ( .A1(n9390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9391) );
  OR2_X1 U11078 ( .A1(n10623), .A2(P1_U3086), .ZN(n9508) );
  NOR2_X1 U11079 ( .A1(n9457), .A2(n9508), .ZN(n9397) );
  NAND3_X1 U11080 ( .A1(n9503), .A2(n9510), .A3(n9397), .ZN(n9399) );
  NAND2_X1 U11081 ( .A1(n14558), .A2(n9419), .ZN(n9396) );
  NAND2_X1 U11082 ( .A1(n8984), .A2(n14562), .ZN(n9393) );
  NAND2_X1 U11083 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11084 ( .A1(n9394), .A2(n14581), .ZN(n9395) );
  NAND2_X1 U11085 ( .A1(n9396), .A2(n9395), .ZN(n9509) );
  AND2_X1 U11086 ( .A1(n9509), .A2(n9397), .ZN(n9475) );
  NAND2_X1 U11087 ( .A1(n9503), .A2(n9475), .ZN(n9398) );
  NAND2_X1 U11088 ( .A1(n9399), .A2(n9398), .ZN(n9474) );
  NAND2_X1 U11089 ( .A1(n9407), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11090 ( .A1(n9408), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9403) );
  INV_X1 U11091 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9400) );
  NOR2_X1 U11092 ( .A1(n9409), .A2(n9400), .ZN(n14582) );
  NAND2_X1 U11093 ( .A1(n9410), .A2(n14582), .ZN(n9402) );
  NAND2_X1 U11094 ( .A1(n9411), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9401) );
  NAND4_X1 U11095 ( .A1(n9404), .A2(n9403), .A3(n9402), .A4(n9401), .ZN(n14355) );
  INV_X1 U11096 ( .A(n14355), .ZN(n12716) );
  NAND2_X1 U11097 ( .A1(n14224), .A2(n9416), .ZN(n9406) );
  NAND2_X1 U11098 ( .A1(n7206), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9405) );
  MUX2_X1 U11099 ( .A(n12716), .B(n14790), .S(n9419), .Z(n9425) );
  MUX2_X1 U11100 ( .A(n14355), .B(n14579), .S(n8984), .Z(n9424) );
  NAND2_X1 U11101 ( .A1(n9425), .A2(n9424), .ZN(n9468) );
  NAND2_X1 U11102 ( .A1(n9474), .A2(n9468), .ZN(n9470) );
  NAND2_X1 U11103 ( .A1(n9407), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11104 ( .A1(n9408), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9414) );
  XNOR2_X1 U11105 ( .A(n9409), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U11106 ( .A1(n9410), .A2(n12713), .ZN(n9413) );
  NAND2_X1 U11107 ( .A1(n9411), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9412) );
  NAND4_X1 U11108 ( .A1(n9415), .A2(n9414), .A3(n9413), .A4(n9412), .ZN(n14586) );
  INV_X1 U11109 ( .A(n14586), .ZN(n14568) );
  NAND2_X1 U11110 ( .A1(n14227), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U11111 ( .A1(n7207), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9417) );
  MUX2_X1 U11112 ( .A(n14568), .B(n7554), .S(n8984), .Z(n9429) );
  MUX2_X1 U11113 ( .A(n14586), .B(n14799), .S(n9419), .Z(n9428) );
  NOR2_X1 U11114 ( .A1(n9429), .A2(n9428), .ZN(n9469) );
  NOR2_X1 U11115 ( .A1(n9470), .A2(n9469), .ZN(n9420) );
  AND2_X1 U11116 ( .A1(n8905), .A2(n11222), .ZN(n9456) );
  INV_X1 U11117 ( .A(n9456), .ZN(n9464) );
  INV_X1 U11118 ( .A(n9511), .ZN(n9423) );
  AOI21_X1 U11119 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9422) );
  AND2_X1 U11120 ( .A1(n9423), .A2(n9422), .ZN(n9517) );
  INV_X1 U11121 ( .A(n9424), .ZN(n9427) );
  INV_X1 U11122 ( .A(n9425), .ZN(n9426) );
  NAND2_X1 U11123 ( .A1(n9427), .A2(n9426), .ZN(n9506) );
  NAND2_X1 U11124 ( .A1(n9517), .A2(n9506), .ZN(n9473) );
  INV_X1 U11125 ( .A(n9473), .ZN(n9430) );
  NAND2_X1 U11126 ( .A1(n9429), .A2(n9428), .ZN(n9471) );
  NAND3_X1 U11127 ( .A1(n9431), .A2(n9430), .A3(n9471), .ZN(n9519) );
  OR2_X1 U11128 ( .A1(n14799), .A2(n14586), .ZN(n9432) );
  NAND2_X1 U11129 ( .A1(n14572), .A2(n9432), .ZN(n12467) );
  INV_X1 U11130 ( .A(n12467), .ZN(n9452) );
  XNOR2_X1 U11131 ( .A(n14604), .B(n14356), .ZN(n12464) );
  XNOR2_X1 U11132 ( .A(n14810), .B(n12444), .ZN(n14620) );
  XNOR2_X1 U11133 ( .A(n14670), .B(n12667), .ZN(n14658) );
  XNOR2_X1 U11134 ( .A(n15953), .B(n15902), .ZN(n14748) );
  XNOR2_X1 U11135 ( .A(n15932), .B(n14766), .ZN(n15911) );
  NAND2_X1 U11136 ( .A1(n14775), .A2(n14361), .ZN(n9433) );
  NAND2_X1 U11137 ( .A1(n15888), .A2(n15904), .ZN(n12436) );
  XNOR2_X1 U11138 ( .A(n12606), .B(n12604), .ZN(n12427) );
  XNOR2_X1 U11139 ( .A(n12281), .B(n12237), .ZN(n12085) );
  XNOR2_X1 U11140 ( .A(n12234), .B(n14365), .ZN(n12079) );
  INV_X1 U11141 ( .A(n12079), .ZN(n9444) );
  XNOR2_X1 U11142 ( .A(n12119), .B(n14366), .ZN(n12100) );
  INV_X1 U11143 ( .A(n9434), .ZN(n9435) );
  OR2_X1 U11144 ( .A1(n9435), .A2(n11233), .ZN(n15540) );
  NAND2_X1 U11145 ( .A1(n11232), .A2(n11234), .ZN(n11224) );
  XNOR2_X1 U11146 ( .A(n14372), .B(n11712), .ZN(n11242) );
  NOR3_X1 U11147 ( .A1(n15540), .A2(n9436), .A3(n11242), .ZN(n9439) );
  INV_X1 U11148 ( .A(n11366), .ZN(n9437) );
  XNOR2_X2 U11149 ( .A(n14374), .B(n11516), .ZN(n11518) );
  AND2_X1 U11150 ( .A1(n9437), .A2(n11518), .ZN(n9438) );
  XNOR2_X1 U11151 ( .A(n11780), .B(n11633), .ZN(n11777) );
  INV_X1 U11152 ( .A(n11777), .ZN(n11784) );
  NAND4_X1 U11153 ( .A1(n9439), .A2(n9438), .A3(n11784), .A4(n15658), .ZN(
        n9440) );
  XNOR2_X1 U11154 ( .A(n11763), .B(n11764), .ZN(n15710) );
  NOR2_X1 U11155 ( .A1(n9440), .A2(n15710), .ZN(n9442) );
  OR2_X1 U11156 ( .A1(n15781), .A2(n14367), .ZN(n12047) );
  NAND2_X1 U11157 ( .A1(n15781), .A2(n14367), .ZN(n9441) );
  NAND2_X1 U11158 ( .A1(n12047), .A2(n9441), .ZN(n15768) );
  XNOR2_X1 U11159 ( .A(n15742), .B(n12044), .ZN(n11718) );
  INV_X1 U11160 ( .A(n11718), .ZN(n11706) );
  NAND4_X1 U11161 ( .A1(n12100), .A2(n9442), .A3(n15768), .A4(n11706), .ZN(
        n9443) );
  OR4_X1 U11162 ( .A1(n12410), .A2(n12085), .A3(n9444), .A4(n9443), .ZN(n9445)
         );
  NOR2_X1 U11163 ( .A1(n12427), .A2(n9445), .ZN(n9446) );
  XNOR2_X1 U11164 ( .A(n12435), .B(n14768), .ZN(n12412) );
  NAND4_X1 U11165 ( .A1(n15911), .A2(n14761), .A3(n9446), .A4(n12412), .ZN(
        n9447) );
  NOR2_X1 U11166 ( .A1(n14748), .A2(n9447), .ZN(n9448) );
  XNOR2_X1 U11167 ( .A(n14848), .B(n14730), .ZN(n14714) );
  INV_X1 U11168 ( .A(n14729), .ZN(n14725) );
  NAND4_X1 U11169 ( .A1(n14701), .A2(n9448), .A3(n14714), .A4(n14725), .ZN(
        n9449) );
  NOR2_X1 U11170 ( .A1(n14658), .A2(n9449), .ZN(n9450) );
  NAND4_X1 U11171 ( .A1(n14630), .A2(n14678), .A3(n9450), .A4(n7960), .ZN(
        n9451) );
  NOR4_X1 U11172 ( .A1(n9452), .A2(n14599), .A3(n14620), .A4(n9451), .ZN(n9454) );
  XNOR2_X1 U11173 ( .A(n14558), .B(n14581), .ZN(n9453) );
  NAND4_X1 U11174 ( .A1(n9503), .A2(n9454), .A3(n14574), .A4(n9453), .ZN(n9455) );
  XNOR2_X1 U11175 ( .A(n9455), .B(n12019), .ZN(n9465) );
  NOR2_X1 U11176 ( .A1(n14562), .A2(n9456), .ZN(n9458) );
  XNOR2_X1 U11177 ( .A(n9419), .B(n9457), .ZN(n9459) );
  AOI21_X1 U11178 ( .B1(n9458), .B2(n9459), .A(n14781), .ZN(n9463) );
  INV_X1 U11179 ( .A(n9459), .ZN(n9461) );
  AOI21_X1 U11180 ( .B1(n9461), .B2(n14562), .A(n9460), .ZN(n9462) );
  OAI22_X1 U11181 ( .A1(n9465), .A2(n9464), .B1(n9463), .B2(n9462), .ZN(n9466)
         );
  INV_X1 U11182 ( .A(n9508), .ZN(n12259) );
  INV_X1 U11183 ( .A(n9468), .ZN(n9516) );
  INV_X1 U11184 ( .A(n9469), .ZN(n9472) );
  OAI22_X1 U11185 ( .A1(n9473), .A2(n9472), .B1(n9471), .B2(n9470), .ZN(n9515)
         );
  INV_X1 U11186 ( .A(n9474), .ZN(n9507) );
  INV_X1 U11187 ( .A(n9475), .ZN(n9477) );
  NOR2_X1 U11188 ( .A1(n9477), .A2(n9476), .ZN(n9504) );
  INV_X1 U11189 ( .A(P1_B_REG_SCAN_IN), .ZN(n10441) );
  NAND2_X1 U11190 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  NAND2_X1 U11191 ( .A1(n9493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9487) );
  MUX2_X1 U11192 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9487), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9489) );
  NAND2_X1 U11193 ( .A1(n9489), .A2(n9488), .ZN(n14889) );
  NAND2_X1 U11194 ( .A1(n9490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9492) );
  INV_X1 U11195 ( .A(n10439), .ZN(n9497) );
  NAND2_X1 U11196 ( .A1(n15536), .A2(n12019), .ZN(n9499) );
  NAND2_X1 U11197 ( .A1(n10359), .A2(n9499), .ZN(n10624) );
  INV_X1 U11198 ( .A(n10359), .ZN(n10628) );
  NOR3_X1 U11199 ( .A1(n11260), .A2(n14886), .A3(n15903), .ZN(n9501) );
  AOI211_X1 U11200 ( .C1(n12259), .C2(n11229), .A(n10441), .B(n9501), .ZN(
        n9502) );
  AOI21_X1 U11201 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(n9505) );
  OAI21_X1 U11202 ( .B1(n9507), .B2(n9506), .A(n9505), .ZN(n9513) );
  NOR4_X1 U11203 ( .A1(n9511), .A2(n9510), .A3(n9509), .A4(n9508), .ZN(n9512)
         );
  AOI211_X1 U11204 ( .C1(n9517), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9518)
         );
  NAND4_X1 U11205 ( .A1(n9520), .A2(n9519), .A3(n9467), .A4(n9518), .ZN(
        P1_U3242) );
  INV_X1 U11206 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10102) );
  INV_X1 U11207 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U11208 ( .A1(n10399), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9522) );
  XNOR2_X1 U11209 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9661) );
  NAND2_X1 U11210 ( .A1(n10424), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9524) );
  INV_X1 U11211 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U11212 ( .A1(n9525), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U11213 ( .A1(n9527), .A2(n9526), .ZN(n9692) );
  NAND2_X1 U11214 ( .A1(n9692), .A2(n9690), .ZN(n9529) );
  NAND2_X1 U11215 ( .A1(n10422), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U11216 ( .A1(n9529), .A2(n9528), .ZN(n9705) );
  NAND2_X1 U11217 ( .A1(n9705), .A2(n9703), .ZN(n9531) );
  NAND2_X1 U11218 ( .A1(n10427), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11219 ( .A1(n10433), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U11220 ( .A1(n9535), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U11221 ( .A1(n10451), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11222 ( .A1(n9538), .A2(n9537), .ZN(n9765) );
  XNOR2_X1 U11223 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9764) );
  NAND2_X1 U11224 ( .A1(n9765), .A2(n9764), .ZN(n9541) );
  NAND2_X1 U11225 ( .A1(n9539), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11226 ( .A1(n9541), .A2(n9540), .ZN(n9782) );
  XNOR2_X1 U11227 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9781) );
  NAND2_X1 U11228 ( .A1(n9782), .A2(n9781), .ZN(n9544) );
  NAND2_X1 U11229 ( .A1(n9542), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9543) );
  XNOR2_X1 U11230 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9794) );
  NAND2_X1 U11231 ( .A1(n9545), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9546) );
  XNOR2_X1 U11232 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9808) );
  INV_X1 U11233 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U11234 ( .A1(n9549), .A2(n9548), .ZN(n9550) );
  XNOR2_X1 U11235 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9830) );
  NAND2_X1 U11236 ( .A1(n10983), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9551) );
  XNOR2_X1 U11237 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9845) );
  NAND2_X1 U11238 ( .A1(n11170), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9552) );
  XNOR2_X1 U11239 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9858) );
  NAND2_X1 U11240 ( .A1(n11399), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U11241 ( .A1(n11677), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9557) );
  INV_X1 U11242 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U11243 ( .A1(n11675), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U11244 ( .A1(n9557), .A2(n9556), .ZN(n9874) );
  XNOR2_X1 U11245 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9904) );
  NAND2_X1 U11246 ( .A1(n9905), .A2(n9904), .ZN(n9559) );
  INV_X1 U11247 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12018) );
  NAND2_X1 U11248 ( .A1(n12018), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U11249 ( .A1(n9560), .A2(n12131), .ZN(n9561) );
  INV_X1 U11250 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12217) );
  NAND2_X1 U11251 ( .A1(n12217), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9564) );
  INV_X1 U11252 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U11253 ( .A1(n12476), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U11254 ( .A1(n9564), .A2(n9563), .ZN(n9927) );
  NAND2_X1 U11255 ( .A1(n9565), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U11256 ( .A1(n12479), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9566) );
  NAND2_X2 U11257 ( .A1(n9945), .A2(n9567), .ZN(n9613) );
  XNOR2_X1 U11258 ( .A(n9610), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9612) );
  XNOR2_X1 U11259 ( .A(n9613), .B(n9612), .ZN(n11356) );
  NOR2_X1 U11260 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n9576) );
  NOR2_X1 U11261 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), 
        .ZN(n9575) );
  NAND2_X1 U11262 ( .A1(n9582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U11263 ( .A1(n11356), .A2(n10130), .ZN(n9586) );
  NAND2_X1 U11264 ( .A1(n10143), .A2(SI_23_), .ZN(n9585) );
  NOR2_X1 U11265 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9697) );
  NAND2_X1 U11266 ( .A1(n9697), .A2(n9696), .ZN(n9711) );
  NOR2_X1 U11267 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_REG3_REG_18__SCAN_IN), 
        .ZN(n9587) );
  INV_X1 U11268 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15108) );
  INV_X1 U11269 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15096) );
  NAND2_X1 U11270 ( .A1(n15108), .A2(n15096), .ZN(n9588) );
  INV_X1 U11271 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12868) );
  OR2_X1 U11272 ( .A1(n9951), .A2(n15015), .ZN(n9589) );
  NAND2_X1 U11273 ( .A1(n9603), .A2(n9589), .ZN(n13142) );
  NAND2_X1 U11274 ( .A1(n9592), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9593) );
  AND2_X2 U11275 ( .A1(n9599), .A2(n9598), .ZN(n9655) );
  NAND2_X1 U11276 ( .A1(n13142), .A2(n10011), .ZN(n9602) );
  AOI22_X1 U11277 ( .A1(n10133), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n10013), 
        .B2(P3_REG2_REG_23__SCAN_IN), .ZN(n9601) );
  AND2_X2 U11278 ( .A1(n9599), .A2(n13405), .ZN(n9682) );
  NAND2_X1 U11279 ( .A1(n10012), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U11280 ( .A1(n13147), .A2(n13158), .ZN(n10266) );
  OR2_X2 U11281 ( .A1(n9603), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U11282 ( .A1(n9603), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U11283 ( .A1(n9625), .A2(n9604), .ZN(n13129) );
  NAND2_X1 U11284 ( .A1(n13129), .A2(n10011), .ZN(n9609) );
  INV_X1 U11285 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13342) );
  NAND2_X1 U11286 ( .A1(n10012), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11287 ( .A1(n9667), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9605) );
  OAI211_X1 U11288 ( .C1(n9641), .C2(n13342), .A(n9606), .B(n9605), .ZN(n9607)
         );
  INV_X1 U11289 ( .A(n9607), .ZN(n9608) );
  INV_X1 U11290 ( .A(n13138), .ZN(n12908) );
  NAND2_X1 U11291 ( .A1(n9610), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9611) );
  XNOR2_X1 U11292 ( .A(n9616), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U11293 ( .A1(n11753), .A2(n10130), .ZN(n9615) );
  NAND2_X1 U11294 ( .A1(n10143), .A2(SI_24_), .ZN(n9614) );
  OR2_X1 U11295 ( .A1(n13136), .A2(n8150), .ZN(n13100) );
  INV_X1 U11296 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U11297 ( .A1(n14894), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U11298 ( .A1(n14240), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9619) );
  AND2_X1 U11299 ( .A1(n9957), .A2(n9619), .ZN(n9620) );
  OR2_X1 U11300 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  NAND2_X1 U11301 ( .A1(n9958), .A2(n9622), .ZN(n11815) );
  NAND2_X1 U11302 ( .A1(n10143), .A2(SI_25_), .ZN(n9623) );
  OR2_X2 U11303 ( .A1(n9625), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U11304 ( .A1(n9625), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U11305 ( .A1(n9980), .A2(n9626), .ZN(n13112) );
  INV_X1 U11306 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U11307 ( .A1(n9682), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U11308 ( .A1(n9667), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9627) );
  OAI211_X1 U11309 ( .C1(n9641), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9630)
         );
  NAND2_X1 U11310 ( .A1(n13339), .A2(n13128), .ZN(n10155) );
  AND2_X1 U11311 ( .A1(n10058), .A2(n10155), .ZN(n13103) );
  NAND2_X1 U11312 ( .A1(n9655), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U11313 ( .A1(n9667), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9633) );
  INV_X1 U11314 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9631) );
  INV_X1 U11315 ( .A(n9648), .ZN(n9638) );
  NAND2_X1 U11316 ( .A1(n9636), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U11317 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  MUX2_X1 U11318 ( .A(SI_0_), .B(n9639), .S(n10397), .Z(n13406) );
  MUX2_X1 U11319 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13406), .S(n10805), .Z(n10906) );
  NAND2_X1 U11320 ( .A1(n10042), .A2(n10906), .ZN(n15548) );
  NAND2_X1 U11321 ( .A1(n9655), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U11322 ( .A1(n9682), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9644) );
  NAND2_X1 U11323 ( .A1(n9667), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9643) );
  INV_X1 U11324 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9640) );
  INV_X1 U11325 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U11326 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9646) );
  XNOR2_X1 U11327 ( .A(n9647), .B(n9646), .ZN(n10954) );
  XNOR2_X1 U11328 ( .A(n9649), .B(n9648), .ZN(n10390) );
  NAND2_X1 U11329 ( .A1(n9675), .A2(n10390), .ZN(n9651) );
  NAND2_X1 U11330 ( .A1(n9664), .A2(SI_1_), .ZN(n9650) );
  OAI211_X1 U11331 ( .C1(n10805), .C2(n10954), .A(n9651), .B(n9650), .ZN(
        n15557) );
  NAND2_X1 U11332 ( .A1(n9652), .A2(n15557), .ZN(n10161) );
  INV_X1 U11333 ( .A(n9652), .ZN(n12924) );
  NAND2_X1 U11334 ( .A1(n15548), .A2(n15549), .ZN(n9654) );
  NAND2_X1 U11335 ( .A1(n9652), .A2(n15553), .ZN(n9653) );
  NAND2_X1 U11336 ( .A1(n9654), .A2(n9653), .ZN(n15573) );
  NAND2_X1 U11337 ( .A1(n9655), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U11338 ( .A1(n9683), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U11339 ( .A1(n9667), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U11340 ( .A1(n9682), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9656) );
  NAND4_X2 U11341 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n15546) );
  INV_X1 U11342 ( .A(n9661), .ZN(n9662) );
  XNOR2_X1 U11343 ( .A(n9663), .B(n9662), .ZN(n10405) );
  NAND2_X1 U11344 ( .A1(n15573), .A2(n15572), .ZN(n9666) );
  INV_X1 U11345 ( .A(n15546), .ZN(n11531) );
  NAND2_X1 U11346 ( .A1(n11531), .A2(n15580), .ZN(n9665) );
  INV_X1 U11347 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15013) );
  NAND2_X1 U11348 ( .A1(n9655), .A2(n15013), .ZN(n9671) );
  NAND2_X1 U11349 ( .A1(n9682), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9670) );
  BUF_X4 U11350 ( .A(n9667), .Z(n10013) );
  NAND2_X1 U11351 ( .A1(n9667), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U11352 ( .A1(n9683), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9668) );
  AND4_X2 U11353 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n15574)
         );
  INV_X1 U11354 ( .A(SI_3_), .ZN(n10408) );
  NAND2_X1 U11355 ( .A1(n9664), .A2(n10408), .ZN(n9680) );
  INV_X1 U11356 ( .A(n9672), .ZN(n9673) );
  XNOR2_X1 U11357 ( .A(n9674), .B(n9673), .ZN(n10409) );
  NAND2_X1 U11358 ( .A1(n9675), .A2(n10409), .ZN(n9679) );
  NAND2_X1 U11359 ( .A1(n9676), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9677) );
  XNOR2_X1 U11360 ( .A(n9677), .B(n9569), .ZN(n10835) );
  NAND2_X1 U11361 ( .A1(n9908), .A2(n10835), .ZN(n9678) );
  NAND2_X1 U11362 ( .A1(n15574), .A2(n11045), .ZN(n10173) );
  INV_X1 U11363 ( .A(n11045), .ZN(n15613) );
  NAND2_X1 U11364 ( .A1(n12923), .A2(n11045), .ZN(n9681) );
  OR2_X1 U11365 ( .A1(n8145), .A2(n9697), .ZN(n11546) );
  NAND2_X1 U11366 ( .A1(n9655), .A2(n11546), .ZN(n9687) );
  NAND2_X1 U11367 ( .A1(n9682), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U11368 ( .A1(n9683), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U11369 ( .A1(n10013), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9684) );
  NAND4_X1 U11370 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n12922) );
  NAND2_X1 U11371 ( .A1(n9688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9689) );
  XNOR2_X1 U11372 ( .A(n9689), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10875) );
  INV_X1 U11373 ( .A(n9690), .ZN(n9691) );
  XNOR2_X1 U11374 ( .A(n9692), .B(n9691), .ZN(n10404) );
  NAND2_X1 U11375 ( .A1(n9675), .A2(n10404), .ZN(n9694) );
  INV_X1 U11376 ( .A(SI_4_), .ZN(n10403) );
  NAND2_X1 U11377 ( .A1(n9664), .A2(n10403), .ZN(n9693) );
  OAI211_X1 U11378 ( .C1(n10875), .C2(n10805), .A(n9694), .B(n9693), .ZN(
        n11189) );
  NAND2_X1 U11379 ( .A1(n11542), .A2(n7634), .ZN(n11541) );
  INV_X1 U11380 ( .A(n11189), .ZN(n15628) );
  NAND2_X1 U11381 ( .A1(n12922), .A2(n15628), .ZN(n9695) );
  OR2_X1 U11382 ( .A1(n9697), .A2(n9696), .ZN(n9698) );
  NAND2_X1 U11383 ( .A1(n9711), .A2(n9698), .ZN(n11685) );
  NAND2_X1 U11384 ( .A1(n9655), .A2(n11685), .ZN(n9702) );
  NAND2_X1 U11385 ( .A1(n9682), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9701) );
  INV_X2 U11386 ( .A(n9641), .ZN(n10133) );
  NAND2_X1 U11387 ( .A1(n10133), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U11388 ( .A1(n10013), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U11389 ( .A1(n9664), .A2(n10406), .ZN(n9710) );
  INV_X1 U11390 ( .A(n9703), .ZN(n9704) );
  XNOR2_X1 U11391 ( .A(n9705), .B(n9704), .ZN(n10407) );
  NAND2_X1 U11392 ( .A1(n10130), .A2(n10407), .ZN(n9709) );
  OR2_X1 U11393 ( .A1(n7305), .A2(n9879), .ZN(n9707) );
  XNOR2_X1 U11394 ( .A(n9707), .B(n9706), .ZN(n10927) );
  NAND2_X1 U11395 ( .A1(n9908), .A2(n10927), .ZN(n9708) );
  NAND2_X1 U11396 ( .A1(n11545), .A2(n11686), .ZN(n10182) );
  INV_X1 U11397 ( .A(n11545), .ZN(n12921) );
  NAND2_X1 U11398 ( .A1(n12921), .A2(n15647), .ZN(n10183) );
  NAND2_X1 U11399 ( .A1(n9711), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U11400 ( .A1(n9723), .A2(n9712), .ZN(n15681) );
  NAND2_X1 U11401 ( .A1(n9655), .A2(n15681), .ZN(n9716) );
  NAND2_X1 U11402 ( .A1(n9682), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U11403 ( .A1(n10133), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U11404 ( .A1(n9667), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9713) );
  OR2_X1 U11405 ( .A1(n9717), .A2(n9879), .ZN(n9718) );
  XNOR2_X1 U11406 ( .A(n9718), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U11407 ( .A1(n9664), .A2(SI_6_), .ZN(n9722) );
  XNOR2_X1 U11408 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9719) );
  XNOR2_X1 U11409 ( .A(n9720), .B(n9719), .ZN(n10400) );
  NAND2_X1 U11410 ( .A1(n9675), .A2(n10400), .ZN(n9721) );
  OAI211_X1 U11411 ( .C1(n10805), .C2(n11056), .A(n9722), .B(n9721), .ZN(
        n15685) );
  AND2_X1 U11412 ( .A1(n12920), .A2(n15685), .ZN(n9737) );
  AND2_X1 U11413 ( .A1(n9723), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9724) );
  OR2_X1 U11414 ( .A1(n9724), .A2(n9740), .ZN(n11671) );
  NAND2_X1 U11415 ( .A1(n10011), .A2(n11671), .ZN(n9728) );
  NAND2_X1 U11416 ( .A1(n10012), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U11417 ( .A1(n10133), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U11418 ( .A1(n10013), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9725) );
  NAND4_X1 U11419 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n12919) );
  NAND2_X1 U11420 ( .A1(n9717), .A2(n9729), .ZN(n9746) );
  NAND2_X1 U11421 ( .A1(n9746), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9731) );
  INV_X1 U11422 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9730) );
  XNOR2_X1 U11423 ( .A(n9731), .B(n9730), .ZN(n11155) );
  INV_X1 U11424 ( .A(n11155), .ZN(n9736) );
  XNOR2_X1 U11425 ( .A(n9733), .B(n9732), .ZN(n10395) );
  NAND2_X1 U11426 ( .A1(n10130), .A2(n10395), .ZN(n9735) );
  NAND2_X1 U11427 ( .A1(n9664), .A2(n15062), .ZN(n9734) );
  OAI211_X1 U11428 ( .C1(n9736), .C2(n10805), .A(n9735), .B(n9734), .ZN(n11649) );
  XNOR2_X1 U11429 ( .A(n12919), .B(n11649), .ZN(n11661) );
  NAND2_X1 U11430 ( .A1(n11666), .A2(n15685), .ZN(n10187) );
  INV_X1 U11431 ( .A(n15685), .ZN(n11737) );
  NAND2_X1 U11432 ( .A1(n12920), .A2(n11737), .ZN(n10188) );
  NAND2_X1 U11433 ( .A1(n10187), .A2(n10188), .ZN(n11732) );
  NAND2_X1 U11434 ( .A1(n11545), .A2(n15647), .ZN(n11728) );
  AND2_X1 U11435 ( .A1(n11732), .A2(n11728), .ZN(n11729) );
  OR2_X1 U11436 ( .A1(n9737), .A2(n11729), .ZN(n11662) );
  AND2_X1 U11437 ( .A1(n11661), .A2(n11662), .ZN(n9738) );
  INV_X1 U11438 ( .A(n11649), .ZN(n15701) );
  NAND2_X1 U11439 ( .A1(n12919), .A2(n15701), .ZN(n9739) );
  NOR2_X1 U11440 ( .A1(n9740), .A2(n15090), .ZN(n9741) );
  OR2_X1 U11441 ( .A1(n9757), .A2(n9741), .ZN(n11797) );
  NAND2_X1 U11442 ( .A1(n10011), .A2(n11797), .ZN(n9745) );
  NAND2_X1 U11443 ( .A1(n10012), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U11444 ( .A1(n10133), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U11445 ( .A1(n10013), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U11446 ( .A1(n9766), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9747) );
  XNOR2_X1 U11447 ( .A(n9747), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11153) );
  INV_X1 U11448 ( .A(n9748), .ZN(n9749) );
  XNOR2_X1 U11449 ( .A(n9750), .B(n9749), .ZN(n10392) );
  NAND2_X1 U11450 ( .A1(n10130), .A2(n10392), .ZN(n9752) );
  NAND2_X1 U11451 ( .A1(n9664), .A2(SI_8_), .ZN(n9751) );
  OAI211_X1 U11452 ( .C1(n10805), .C2(n12972), .A(n9752), .B(n9751), .ZN(
        n15736) );
  NAND2_X1 U11453 ( .A1(n11879), .A2(n15736), .ZN(n10195) );
  INV_X1 U11454 ( .A(n11879), .ZN(n12918) );
  INV_X1 U11455 ( .A(n15736), .ZN(n9754) );
  NAND2_X1 U11456 ( .A1(n12918), .A2(n9754), .ZN(n10196) );
  NOR2_X1 U11457 ( .A1(n11792), .A2(n11796), .ZN(n9753) );
  INV_X1 U11458 ( .A(n9753), .ZN(n11791) );
  NAND2_X1 U11459 ( .A1(n11879), .A2(n9754), .ZN(n9755) );
  NAND2_X1 U11460 ( .A1(n11791), .A2(n9755), .ZN(n11855) );
  OR2_X1 U11461 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  NAND2_X1 U11462 ( .A1(n9775), .A2(n9758), .ZN(n11890) );
  NAND2_X1 U11463 ( .A1(n10011), .A2(n11890), .ZN(n9763) );
  NAND2_X1 U11464 ( .A1(n10012), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U11465 ( .A1(n10013), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11466 ( .A1(n10133), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9760) );
  NAND4_X1 U11467 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n12917) );
  XNOR2_X1 U11468 ( .A(n9765), .B(n9764), .ZN(n10396) );
  NAND2_X1 U11469 ( .A1(n10130), .A2(n10396), .ZN(n9773) );
  NAND2_X1 U11470 ( .A1(n10143), .A2(n14910), .ZN(n9772) );
  NOR2_X1 U11471 ( .A1(n9766), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9769) );
  OR2_X1 U11472 ( .A1(n9769), .A2(n9879), .ZN(n9767) );
  INV_X1 U11473 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U11474 ( .A(n9767), .B(P3_IR_REG_31__SCAN_IN), .S(n9768), .Z(n9770)
         );
  NAND2_X1 U11475 ( .A1(n9769), .A2(n9768), .ZN(n9796) );
  NAND2_X1 U11476 ( .A1(n9770), .A2(n9796), .ZN(n12975) );
  NAND2_X1 U11477 ( .A1(n9908), .A2(n12975), .ZN(n9771) );
  NOR2_X1 U11478 ( .A1(n12917), .A2(n11876), .ZN(n9774) );
  NAND2_X1 U11479 ( .A1(n9775), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U11480 ( .A1(n9788), .A2(n9776), .ZN(n11901) );
  NAND2_X1 U11481 ( .A1(n10011), .A2(n11901), .ZN(n9780) );
  NAND2_X1 U11482 ( .A1(n10012), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9779) );
  NAND2_X1 U11483 ( .A1(n10133), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U11484 ( .A1(n10013), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9777) );
  XNOR2_X1 U11485 ( .A(n9782), .B(n9781), .ZN(n10410) );
  NAND2_X1 U11486 ( .A1(n10130), .A2(n10410), .ZN(n9787) );
  NAND2_X1 U11487 ( .A1(n10143), .A2(n14909), .ZN(n9786) );
  NAND2_X1 U11488 ( .A1(n9796), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9784) );
  XNOR2_X1 U11489 ( .A(n9784), .B(n9783), .ZN(n12971) );
  NAND2_X1 U11490 ( .A1(n9908), .A2(n12971), .ZN(n9785) );
  NAND2_X1 U11491 ( .A1(n12143), .A2(n11987), .ZN(n10204) );
  INV_X1 U11492 ( .A(n12143), .ZN(n12916) );
  INV_X1 U11493 ( .A(n11987), .ZN(n15789) );
  NAND2_X1 U11494 ( .A1(n12916), .A2(n15789), .ZN(n10205) );
  NAND2_X1 U11495 ( .A1(n10204), .A2(n10205), .ZN(n11897) );
  NAND2_X1 U11496 ( .A1(n9788), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U11497 ( .A1(n9802), .A2(n9789), .ZN(n12145) );
  NAND2_X1 U11498 ( .A1(n10011), .A2(n12145), .ZN(n9793) );
  NAND2_X1 U11499 ( .A1(n10012), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U11500 ( .A1(n9667), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U11501 ( .A1(n10133), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9790) );
  NAND4_X1 U11502 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(n12915) );
  XNOR2_X1 U11503 ( .A(n9795), .B(n9794), .ZN(n10411) );
  NAND2_X1 U11504 ( .A1(n10130), .A2(n10411), .ZN(n9801) );
  NAND2_X1 U11505 ( .A1(n10143), .A2(n15057), .ZN(n9800) );
  OAI21_X1 U11506 ( .B1(n9796), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9798) );
  INV_X1 U11507 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9797) );
  XNOR2_X1 U11508 ( .A(n9798), .B(n9797), .ZN(n12978) );
  NAND2_X1 U11509 ( .A1(n9908), .A2(n12978), .ZN(n9799) );
  NAND2_X1 U11510 ( .A1(n12157), .A2(n15798), .ZN(n12137) );
  AND2_X1 U11511 ( .A1(n9802), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9803) );
  OR2_X1 U11512 ( .A1(n9803), .A2(n9824), .ZN(n12179) );
  NAND2_X1 U11513 ( .A1(n10011), .A2(n12179), .ZN(n9807) );
  NAND2_X1 U11514 ( .A1(n10012), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U11515 ( .A1(n10013), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U11516 ( .A1(n10133), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9804) );
  NAND4_X1 U11517 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n12914) );
  XNOR2_X1 U11518 ( .A(n9809), .B(n9808), .ZN(n10425) );
  NAND2_X1 U11519 ( .A1(n10425), .A2(n10130), .ZN(n9814) );
  NAND2_X1 U11520 ( .A1(n9811), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9810) );
  MUX2_X1 U11521 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9810), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9812) );
  OR2_X2 U11522 ( .A1(n9811), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U11523 ( .A1(n9812), .A2(n9832), .ZN(n15433) );
  AOI22_X1 U11524 ( .A1(n10143), .A2(n15053), .B1(n9908), .B2(n15433), .ZN(
        n9813) );
  NAND2_X1 U11525 ( .A1(n12914), .A2(n10053), .ZN(n9815) );
  NAND2_X1 U11526 ( .A1(n12155), .A2(n9815), .ZN(n9817) );
  INV_X1 U11527 ( .A(n12914), .ZN(n11995) );
  NAND2_X1 U11528 ( .A1(n11995), .A2(n12280), .ZN(n9816) );
  XNOR2_X1 U11529 ( .A(n9818), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U11530 ( .A1(n10437), .A2(n10130), .ZN(n9822) );
  INV_X1 U11531 ( .A(SI_13_), .ZN(n10438) );
  NAND2_X1 U11532 ( .A1(n9832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9820) );
  INV_X1 U11533 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9819) );
  XNOR2_X1 U11534 ( .A(n9820), .B(n9819), .ZN(n12982) );
  AOI22_X1 U11535 ( .A1(n10143), .A2(n10438), .B1(n9908), .B2(n12982), .ZN(
        n9821) );
  OR2_X1 U11536 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  NAND2_X1 U11537 ( .A1(n9837), .A2(n9825), .ZN(n12355) );
  NAND2_X1 U11538 ( .A1(n10011), .A2(n12355), .ZN(n9829) );
  NAND2_X1 U11539 ( .A1(n10012), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U11540 ( .A1(n10133), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U11541 ( .A1(n10013), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9826) );
  XNOR2_X1 U11542 ( .A(n9831), .B(n9830), .ZN(n10448) );
  NAND2_X1 U11543 ( .A1(n10448), .A2(n10130), .ZN(n9836) );
  NAND2_X1 U11544 ( .A1(n7231), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9834) );
  XNOR2_X1 U11545 ( .A(n9834), .B(n9833), .ZN(n12970) );
  AOI22_X1 U11546 ( .A1(n10143), .A2(n14943), .B1(n9908), .B2(n12970), .ZN(
        n9835) );
  NAND2_X1 U11547 ( .A1(n9837), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U11548 ( .A1(n9850), .A2(n9838), .ZN(n12783) );
  NAND2_X1 U11549 ( .A1(n10011), .A2(n12783), .ZN(n9842) );
  NAND2_X1 U11550 ( .A1(n10012), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U11551 ( .A1(n10133), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U11552 ( .A1(n10013), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9839) );
  NAND4_X1 U11553 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n12912) );
  OR2_X1 U11554 ( .A1(n13390), .A2(n12912), .ZN(n10055) );
  NAND2_X1 U11555 ( .A1(n13390), .A2(n12912), .ZN(n10218) );
  INV_X1 U11556 ( .A(n12912), .ZN(n12898) );
  OR2_X1 U11557 ( .A1(n13390), .A2(n12898), .ZN(n9844) );
  NAND2_X1 U11558 ( .A1(n12262), .A2(n9844), .ZN(n12330) );
  XNOR2_X1 U11559 ( .A(n9846), .B(n9845), .ZN(n10457) );
  NAND2_X1 U11560 ( .A1(n10457), .A2(n10130), .ZN(n9849) );
  OR2_X1 U11561 ( .A1(n9862), .A2(n9879), .ZN(n9847) );
  XNOR2_X1 U11562 ( .A(n9847), .B(n9861), .ZN(n15490) );
  AOI22_X1 U11563 ( .A1(n10143), .A2(n15046), .B1(n9908), .B2(n15490), .ZN(
        n9848) );
  INV_X1 U11564 ( .A(n9866), .ZN(n9852) );
  NAND2_X1 U11565 ( .A1(n9850), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11566 ( .A1(n9852), .A2(n9851), .ZN(n12901) );
  NAND2_X1 U11567 ( .A1(n9655), .A2(n12901), .ZN(n9856) );
  NAND2_X1 U11568 ( .A1(n10012), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U11569 ( .A1(n10133), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11570 ( .A1(n10013), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9853) );
  NAND4_X1 U11571 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(n12911) );
  OR2_X1 U11572 ( .A1(n13386), .A2(n12911), .ZN(n10224) );
  NAND2_X1 U11573 ( .A1(n13386), .A2(n12911), .ZN(n10225) );
  NAND2_X1 U11574 ( .A1(n10224), .A2(n10225), .ZN(n12329) );
  INV_X1 U11575 ( .A(n12911), .ZN(n13241) );
  OR2_X1 U11576 ( .A1(n13386), .A2(n13241), .ZN(n9857) );
  INV_X1 U11577 ( .A(n9858), .ZN(n9859) );
  XNOR2_X1 U11578 ( .A(n9860), .B(n9859), .ZN(n10572) );
  NAND2_X1 U11579 ( .A1(n10572), .A2(n10130), .ZN(n9865) );
  OR2_X1 U11580 ( .A1(n9878), .A2(n9879), .ZN(n9863) );
  XNOR2_X1 U11581 ( .A(n9863), .B(P3_IR_REG_16__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U11582 ( .A1(n10143), .A2(SI_16_), .B1(n9908), .B2(n15510), .ZN(
        n9864) );
  NAND2_X1 U11583 ( .A1(n9865), .A2(n9864), .ZN(n13247) );
  NOR2_X1 U11584 ( .A1(n9866), .A2(n12829), .ZN(n9867) );
  OR2_X1 U11585 ( .A1(n9896), .A2(n9867), .ZN(n13248) );
  NAND2_X1 U11586 ( .A1(n10011), .A2(n13248), .ZN(n9871) );
  NAND2_X1 U11587 ( .A1(n10012), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U11588 ( .A1(n10133), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U11589 ( .A1(n9667), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9868) );
  OR2_X1 U11590 ( .A1(n13247), .A2(n12838), .ZN(n10230) );
  NAND2_X1 U11591 ( .A1(n13247), .A2(n12838), .ZN(n10228) );
  OR2_X1 U11592 ( .A1(n13247), .A2(n13225), .ZN(n9873) );
  INV_X1 U11593 ( .A(n9874), .ZN(n9875) );
  XNOR2_X1 U11594 ( .A(n9876), .B(n9875), .ZN(n10574) );
  NAND2_X1 U11595 ( .A1(n10574), .A2(n10130), .ZN(n9882) );
  INV_X1 U11596 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9877) );
  OR2_X1 U11597 ( .A1(n9891), .A2(n9879), .ZN(n9880) );
  XNOR2_X1 U11598 ( .A(n9880), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U11599 ( .A1(n10143), .A2(n15044), .B1(n9908), .B2(n12993), .ZN(
        n9881) );
  INV_X1 U11600 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9895) );
  XNOR2_X1 U11601 ( .A(n9896), .B(n9895), .ZN(n13231) );
  NAND2_X1 U11602 ( .A1(n10011), .A2(n13231), .ZN(n9886) );
  NAND2_X1 U11603 ( .A1(n10012), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U11604 ( .A1(n10133), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U11605 ( .A1(n10013), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9883) );
  NAND4_X1 U11606 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n12910) );
  NAND2_X1 U11607 ( .A1(n13378), .A2(n12910), .ZN(n10233) );
  NAND2_X1 U11608 ( .A1(n10238), .A2(n10233), .ZN(n13223) );
  OR2_X1 U11609 ( .A1(n13378), .A2(n13242), .ZN(n9887) );
  AOI22_X1 U11610 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11907), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11909), .ZN(n9888) );
  XNOR2_X1 U11611 ( .A(n9889), .B(n9888), .ZN(n10659) );
  NAND2_X1 U11612 ( .A1(n10659), .A2(n10130), .ZN(n9894) );
  NAND2_X1 U11613 ( .A1(n9906), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9892) );
  XNOR2_X1 U11614 ( .A(n9892), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U11615 ( .A1(n10143), .A2(SI_18_), .B1(n9908), .B2(n13032), .ZN(
        n9893) );
  NAND2_X1 U11616 ( .A1(n9894), .A2(n9893), .ZN(n12878) );
  NAND2_X1 U11617 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  NAND2_X1 U11618 ( .A1(n9897), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U11619 ( .A1(n9898), .A2(n9911), .ZN(n13217) );
  NAND2_X1 U11620 ( .A1(n9655), .A2(n13217), .ZN(n9902) );
  NAND2_X1 U11621 ( .A1(n10012), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U11622 ( .A1(n10133), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U11623 ( .A1(n10013), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9899) );
  OR2_X1 U11624 ( .A1(n12878), .A2(n13198), .ZN(n10235) );
  NAND2_X1 U11625 ( .A1(n12878), .A2(n13198), .ZN(n10236) );
  NAND2_X1 U11626 ( .A1(n10235), .A2(n10236), .ZN(n10305) );
  INV_X1 U11627 ( .A(n13198), .ZN(n13224) );
  OR2_X1 U11628 ( .A1(n12878), .A2(n13224), .ZN(n9903) );
  NAND2_X1 U11629 ( .A1(n13209), .A2(n9903), .ZN(n13197) );
  XNOR2_X1 U11630 ( .A(n9905), .B(n9904), .ZN(n10744) );
  NAND2_X1 U11631 ( .A1(n10744), .A2(n10130), .ZN(n9910) );
  AOI22_X1 U11632 ( .A1(n10143), .A2(SI_19_), .B1(n7209), .B2(n9908), .ZN(
        n9909) );
  NAND2_X1 U11633 ( .A1(n9911), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U11634 ( .A1(n9932), .A2(n9912), .ZN(n13204) );
  NAND2_X1 U11635 ( .A1(n9655), .A2(n13204), .ZN(n9916) );
  NAND2_X1 U11636 ( .A1(n10012), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U11637 ( .A1(n10013), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U11638 ( .A1(n10133), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9913) );
  NAND4_X1 U11639 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n13186) );
  NOR2_X1 U11640 ( .A1(n13369), .A2(n13186), .ZN(n9917) );
  INV_X1 U11641 ( .A(n13369), .ZN(n13206) );
  XNOR2_X1 U11642 ( .A(n9918), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U11643 ( .A1(n11067), .A2(n10130), .ZN(n9920) );
  NAND2_X1 U11644 ( .A1(n10143), .A2(SI_20_), .ZN(n9919) );
  XNOR2_X1 U11645 ( .A(n9932), .B(P3_REG3_REG_20__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U11646 ( .A1(n13192), .A2(n10011), .ZN(n9924) );
  NAND2_X1 U11647 ( .A1(n10133), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U11648 ( .A1(n10013), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U11649 ( .A1(n10012), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9921) );
  OR2_X1 U11650 ( .A1(n13362), .A2(n13199), .ZN(n10247) );
  NAND2_X1 U11651 ( .A1(n13362), .A2(n13199), .ZN(n10248) );
  NAND2_X1 U11652 ( .A1(n13184), .A2(n7672), .ZN(n9926) );
  INV_X1 U11653 ( .A(n13199), .ZN(n13172) );
  NAND2_X1 U11654 ( .A1(n13362), .A2(n13172), .ZN(n9925) );
  INV_X1 U11655 ( .A(n9927), .ZN(n9928) );
  XNOR2_X1 U11656 ( .A(n9929), .B(n9928), .ZN(n11092) );
  NAND2_X1 U11657 ( .A1(n11092), .A2(n10130), .ZN(n9931) );
  NAND2_X1 U11658 ( .A1(n10143), .A2(SI_21_), .ZN(n9930) );
  OAI21_X1 U11659 ( .B1(n9932), .B2(P3_REG3_REG_20__SCAN_IN), .A(
        P3_REG3_REG_21__SCAN_IN), .ZN(n9933) );
  INV_X1 U11660 ( .A(n9933), .ZN(n9934) );
  OR2_X1 U11661 ( .A1(n9934), .A2(n9949), .ZN(n13177) );
  NAND2_X1 U11662 ( .A1(n13177), .A2(n10011), .ZN(n9939) );
  NAND2_X1 U11663 ( .A1(n10133), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U11664 ( .A1(n10013), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9935) );
  AND2_X1 U11665 ( .A1(n9936), .A2(n9935), .ZN(n9938) );
  NAND2_X1 U11666 ( .A1(n10012), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U11667 ( .A1(n13178), .A2(n13157), .ZN(n10056) );
  INV_X1 U11668 ( .A(n13157), .ZN(n13187) );
  OR2_X1 U11669 ( .A1(n13178), .A2(n13187), .ZN(n9941) );
  OR2_X1 U11670 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  NAND2_X1 U11671 ( .A1(n9945), .A2(n9944), .ZN(n11178) );
  OR2_X1 U11672 ( .A1(n11178), .A2(n9946), .ZN(n9948) );
  NAND2_X1 U11673 ( .A1(n10143), .A2(SI_22_), .ZN(n9947) );
  INV_X1 U11674 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13284) );
  NOR2_X1 U11675 ( .A1(n9949), .A2(n12868), .ZN(n9950) );
  OR2_X1 U11676 ( .A1(n9951), .A2(n9950), .ZN(n13163) );
  NAND2_X1 U11677 ( .A1(n13163), .A2(n10011), .ZN(n9953) );
  AOI22_X1 U11678 ( .A1(n10133), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n10013), 
        .B2(P3_REG2_REG_22__SCAN_IN), .ZN(n9952) );
  OAI211_X1 U11679 ( .C1(n9759), .C2(n13284), .A(n9953), .B(n9952), .ZN(n13173) );
  NAND2_X1 U11680 ( .A1(n13351), .A2(n13173), .ZN(n9954) );
  NAND2_X1 U11681 ( .A1(n13156), .A2(n9954), .ZN(n9956) );
  OR2_X1 U11682 ( .A1(n13351), .A2(n13173), .ZN(n9955) );
  NAND2_X1 U11683 ( .A1(n13276), .A2(n13138), .ZN(n10261) );
  NAND2_X1 U11684 ( .A1(n10262), .A2(n10261), .ZN(n13124) );
  NAND2_X1 U11685 ( .A1(n13147), .A2(n12909), .ZN(n13121) );
  AND2_X1 U11686 ( .A1(n13124), .A2(n13121), .ZN(n13122) );
  OR2_X1 U11687 ( .A1(n8150), .A2(n13122), .ZN(n13101) );
  INV_X1 U11688 ( .A(n13128), .ZN(n12907) );
  NAND2_X1 U11689 ( .A1(n14891), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U11690 ( .A1(n9959), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9960) );
  NAND2_X1 U11691 ( .A1(n9974), .A2(n9960), .ZN(n9971) );
  NAND2_X1 U11692 ( .A1(n11928), .A2(n10130), .ZN(n9962) );
  NAND2_X1 U11693 ( .A1(n10143), .A2(SI_26_), .ZN(n9961) );
  XNOR2_X1 U11694 ( .A(n9980), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U11695 ( .A1(n13096), .A2(n10011), .ZN(n9967) );
  INV_X1 U11696 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U11697 ( .A1(n10012), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11698 ( .A1(n10013), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U11699 ( .C1(n9641), .C2(n13332), .A(n9964), .B(n9963), .ZN(n9965)
         );
  INV_X1 U11700 ( .A(n9965), .ZN(n9966) );
  OR2_X1 U11701 ( .A1(n13333), .A2(n12906), .ZN(n9968) );
  NAND2_X1 U11702 ( .A1(n13090), .A2(n9968), .ZN(n9970) );
  NAND2_X1 U11703 ( .A1(n13333), .A2(n12906), .ZN(n9969) );
  NAND2_X1 U11704 ( .A1(n9970), .A2(n9969), .ZN(n13079) );
  INV_X1 U11705 ( .A(n13079), .ZN(n9986) );
  INV_X1 U11706 ( .A(n9971), .ZN(n9972) );
  NAND2_X1 U11707 ( .A1(n14888), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U11708 ( .A1(n14232), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U11709 ( .A1(n9991), .A2(n9975), .ZN(n9988) );
  NAND2_X1 U11710 ( .A1(n12128), .A2(n10130), .ZN(n9977) );
  NAND2_X1 U11711 ( .A1(n10143), .A2(SI_27_), .ZN(n9976) );
  OAI21_X1 U11712 ( .B1(n9980), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n9978) );
  INV_X1 U11713 ( .A(n9978), .ZN(n9981) );
  INV_X1 U11714 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15083) );
  INV_X1 U11715 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15121) );
  NAND2_X1 U11716 ( .A1(n15083), .A2(n15121), .ZN(n9979) );
  INV_X1 U11717 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U11718 ( .A1(n9682), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U11719 ( .A1(n10013), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9982) );
  OAI211_X1 U11720 ( .C1(n9641), .C2(n13325), .A(n9983), .B(n9982), .ZN(n9984)
         );
  OR2_X2 U11721 ( .A1(n13326), .A2(n13091), .ZN(n10158) );
  NAND2_X1 U11722 ( .A1(n13326), .A2(n13091), .ZN(n10156) );
  INV_X1 U11723 ( .A(n13091), .ZN(n12905) );
  OR2_X1 U11724 ( .A1(n13326), .A2(n12905), .ZN(n9987) );
  INV_X1 U11725 ( .A(n9988), .ZN(n9989) );
  NAND2_X1 U11726 ( .A1(n9990), .A2(n9989), .ZN(n9992) );
  NAND2_X1 U11727 ( .A1(n14885), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U11728 ( .A1(n9993), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U11729 ( .A1(n10007), .A2(n9994), .ZN(n10004) );
  XNOR2_X1 U11730 ( .A(n10006), .B(n10004), .ZN(n12132) );
  NAND2_X1 U11731 ( .A1(n12132), .A2(n10130), .ZN(n9996) );
  NAND2_X1 U11732 ( .A1(n10143), .A2(SI_28_), .ZN(n9995) );
  INV_X1 U11733 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12806) );
  NOR2_X1 U11734 ( .A1(n9997), .A2(n12806), .ZN(n9998) );
  INV_X1 U11735 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U11736 ( .A1(n10012), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10000) );
  NAND2_X1 U11737 ( .A1(n10013), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9999) );
  OAI211_X1 U11738 ( .C1(n9641), .C2(n13320), .A(n10000), .B(n9999), .ZN(
        n10001) );
  NAND2_X1 U11739 ( .A1(n10002), .A2(n13077), .ZN(n10274) );
  INV_X1 U11740 ( .A(n13077), .ZN(n10003) );
  INV_X1 U11741 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U11742 ( .A1(n10006), .A2(n10005), .ZN(n10008) );
  XNOR2_X1 U11743 ( .A(n10121), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n10118) );
  XNOR2_X1 U11744 ( .A(n10120), .B(n10118), .ZN(n12199) );
  NAND2_X1 U11745 ( .A1(n12199), .A2(n10130), .ZN(n10010) );
  NAND2_X1 U11746 ( .A1(n10143), .A2(SI_29_), .ZN(n10009) );
  NAND2_X1 U11747 ( .A1(n10010), .A2(n10009), .ZN(n10103) );
  NAND2_X1 U11748 ( .A1(n13055), .A2(n10011), .ZN(n10138) );
  INV_X1 U11749 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U11750 ( .A1(n10013), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U11751 ( .A1(n10133), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10014) );
  OAI211_X1 U11752 ( .C1(n10116), .C2(n9759), .A(n10015), .B(n10014), .ZN(
        n10016) );
  INV_X1 U11753 ( .A(n10016), .ZN(n10017) );
  OR2_X1 U11754 ( .A1(n10103), .A2(n13064), .ZN(n10282) );
  NAND2_X1 U11755 ( .A1(n10103), .A2(n13064), .ZN(n10139) );
  NAND2_X1 U11756 ( .A1(n10282), .A2(n10139), .ZN(n10272) );
  XNOR2_X1 U11757 ( .A(n10019), .B(n10018), .ZN(n10031) );
  NOR2_X2 U11758 ( .A1(n7231), .A2(n10020), .ZN(n10026) );
  NAND2_X1 U11759 ( .A1(n10092), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10023) );
  XNOR2_X1 U11760 ( .A(n10023), .B(n10022), .ZN(n10063) );
  NAND2_X1 U11761 ( .A1(n7209), .A2(n11176), .ZN(n10061) );
  NAND2_X1 U11762 ( .A1(n10030), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10024) );
  MUX2_X1 U11763 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10024), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n10025) );
  INV_X1 U11764 ( .A(n10026), .ZN(n10027) );
  NAND2_X1 U11765 ( .A1(n10027), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10028) );
  MUX2_X1 U11766 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10028), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n10029) );
  INV_X1 U11767 ( .A(n11070), .ZN(n10060) );
  NAND2_X1 U11768 ( .A1(n10165), .A2(n10060), .ZN(n10150) );
  NAND2_X1 U11769 ( .A1(n10031), .A2(n15577), .ZN(n10041) );
  INV_X1 U11770 ( .A(n12134), .ZN(n10820) );
  NAND2_X1 U11771 ( .A1(n10820), .A2(n7384), .ZN(n10807) );
  NAND2_X1 U11772 ( .A1(n10807), .A2(n10805), .ZN(n10788) );
  INV_X1 U11773 ( .A(P3_B_REG_SCAN_IN), .ZN(n10033) );
  NOR2_X1 U11774 ( .A1(n12134), .A2(n10033), .ZN(n10034) );
  OR2_X1 U11775 ( .A1(n13243), .A2(n10034), .ZN(n13047) );
  NAND2_X1 U11776 ( .A1(n10012), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U11777 ( .A1(n10133), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10036) );
  NAND2_X1 U11778 ( .A1(n10013), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10035) );
  AND3_X1 U11779 ( .A1(n10037), .A2(n10036), .A3(n10035), .ZN(n10038) );
  INV_X1 U11780 ( .A(n10039), .ZN(n10040) );
  INV_X1 U11781 ( .A(n15572), .ZN(n10044) );
  INV_X1 U11782 ( .A(n10906), .ZN(n15127) );
  NOR2_X2 U11783 ( .A1(n10042), .A2(n15127), .ZN(n15544) );
  NAND2_X1 U11784 ( .A1(n15544), .A2(n10160), .ZN(n10043) );
  NAND2_X1 U11785 ( .A1(n10044), .A2(n10163), .ZN(n10045) );
  INV_X1 U11786 ( .A(n15580), .ZN(n15586) );
  NAND2_X1 U11787 ( .A1(n11531), .A2(n15586), .ZN(n10171) );
  NAND2_X1 U11788 ( .A1(n10045), .A2(n10171), .ZN(n11527) );
  NAND2_X1 U11789 ( .A1(n11527), .A2(n11528), .ZN(n10046) );
  INV_X1 U11790 ( .A(n12922), .ZN(n11530) );
  NAND2_X1 U11791 ( .A1(n11530), .A2(n15628), .ZN(n10177) );
  NAND2_X1 U11792 ( .A1(n10047), .A2(n10182), .ZN(n11727) );
  INV_X1 U11793 ( .A(n11732), .ZN(n10185) );
  NAND2_X1 U11794 ( .A1(n11727), .A2(n10185), .ZN(n10048) );
  NAND2_X1 U11795 ( .A1(n10048), .A2(n10187), .ZN(n11660) );
  INV_X1 U11796 ( .A(n11661), .ZN(n11664) );
  NAND2_X1 U11797 ( .A1(n11660), .A2(n11664), .ZN(n10050) );
  INV_X1 U11798 ( .A(n12919), .ZN(n11794) );
  NAND2_X1 U11799 ( .A1(n11794), .A2(n15701), .ZN(n10049) );
  NAND2_X1 U11800 ( .A1(n10050), .A2(n10049), .ZN(n11795) );
  NAND2_X1 U11801 ( .A1(n11795), .A2(n11796), .ZN(n10051) );
  NOR2_X1 U11802 ( .A1(n12917), .A2(n11924), .ZN(n10199) );
  NAND2_X1 U11803 ( .A1(n12917), .A2(n11924), .ZN(n10201) );
  NAND2_X1 U11804 ( .A1(n11895), .A2(n10204), .ZN(n11997) );
  NAND2_X1 U11805 ( .A1(n12157), .A2(n10052), .ZN(n10208) );
  NAND2_X1 U11806 ( .A1(n12915), .A2(n15798), .ZN(n12172) );
  NAND2_X1 U11807 ( .A1(n11995), .A2(n10053), .ZN(n10213) );
  NAND2_X1 U11808 ( .A1(n12914), .A2(n12280), .ZN(n10212) );
  NAND2_X1 U11809 ( .A1(n12738), .A2(n12913), .ZN(n10054) );
  NAND2_X1 U11810 ( .A1(n12268), .A2(n12267), .ZN(n12266) );
  NAND2_X1 U11811 ( .A1(n12266), .A2(n10055), .ZN(n12335) );
  INV_X1 U11812 ( .A(n12329), .ZN(n12334) );
  NAND2_X1 U11813 ( .A1(n12335), .A2(n12334), .ZN(n12333) );
  NAND2_X1 U11814 ( .A1(n13214), .A2(n10236), .ZN(n13202) );
  INV_X1 U11815 ( .A(n10056), .ZN(n10250) );
  INV_X1 U11816 ( .A(n13173), .ZN(n13137) );
  NOR2_X1 U11817 ( .A1(n13351), .A2(n13137), .ZN(n10257) );
  NAND2_X1 U11818 ( .A1(n13351), .A2(n13137), .ZN(n10253) );
  INV_X1 U11819 ( .A(n13124), .ZN(n13117) );
  NAND2_X1 U11820 ( .A1(n13333), .A2(n13106), .ZN(n10154) );
  INV_X1 U11821 ( .A(n13068), .ZN(n10307) );
  INV_X1 U11822 ( .A(n10273), .ZN(n10059) );
  XOR2_X1 U11823 ( .A(n10272), .B(n10147), .Z(n13059) );
  NAND2_X1 U11824 ( .A1(n11525), .A2(n10060), .ZN(n10761) );
  OR2_X1 U11825 ( .A1(n10061), .A2(n10761), .ZN(n10774) );
  NAND3_X1 U11826 ( .A1(n10783), .A2(n10774), .A3(n10285), .ZN(n10778) );
  INV_X1 U11827 ( .A(n7209), .ZN(n13042) );
  NAND2_X1 U11828 ( .A1(n13042), .A2(n11070), .ZN(n10318) );
  OR2_X1 U11829 ( .A1(n10318), .A2(n15737), .ZN(n10062) );
  OR2_X1 U11830 ( .A1(n10778), .A2(n10062), .ZN(n10064) );
  OR2_X1 U11831 ( .A1(n11526), .A2(n11176), .ZN(n15732) );
  AND2_X1 U11832 ( .A1(n13059), .A2(n15802), .ZN(n10065) );
  NOR2_X1 U11833 ( .A1(n13054), .A2(n10065), .ZN(n10115) );
  INV_X1 U11834 ( .A(n10067), .ZN(n10068) );
  INV_X1 U11835 ( .A(n10069), .ZN(n10070) );
  NAND2_X1 U11836 ( .A1(n10070), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U11837 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10071), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n10073) );
  INV_X1 U11838 ( .A(n10066), .ZN(n10072) );
  XNOR2_X1 U11839 ( .A(n11756), .B(P3_B_REG_SCAN_IN), .ZN(n10074) );
  INV_X1 U11840 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U11841 ( .A1(n11930), .A2(n11756), .ZN(n10077) );
  INV_X1 U11842 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11843 ( .A1(n7229), .A2(n10079), .ZN(n10081) );
  NAND2_X1 U11844 ( .A1(n11930), .A2(n11816), .ZN(n10080) );
  NOR2_X1 U11845 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n10085) );
  NOR4_X1 U11846 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10084) );
  NOR4_X1 U11847 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10083) );
  NOR4_X1 U11848 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10082) );
  NAND4_X1 U11849 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10091) );
  NOR4_X1 U11850 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10089) );
  NOR4_X1 U11851 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10088) );
  NOR4_X1 U11852 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n10087) );
  NOR4_X1 U11853 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n10086) );
  NAND4_X1 U11854 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10090) );
  OAI21_X1 U11855 ( .B1(n10091), .B2(n10090), .A(n7229), .ZN(n10109) );
  INV_X1 U11856 ( .A(n11816), .ZN(n10097) );
  INV_X1 U11857 ( .A(n11756), .ZN(n10096) );
  NAND3_X1 U11858 ( .A1(n10097), .A2(n10096), .A3(n10095), .ZN(n10773) );
  NAND2_X1 U11859 ( .A1(n10789), .A2(n10803), .ZN(n10098) );
  OR2_X1 U11860 ( .A1(n10778), .A2(n10098), .ZN(n10101) );
  INV_X1 U11861 ( .A(n10108), .ZN(n13394) );
  AND3_X1 U11862 ( .A1(n13392), .A2(n13394), .A3(n10109), .ZN(n10777) );
  AND2_X1 U11863 ( .A1(n10777), .A2(n10803), .ZN(n10781) );
  OR2_X1 U11864 ( .A1(n10318), .A2(n10285), .ZN(n10899) );
  NAND2_X1 U11865 ( .A1(n10899), .A2(n10774), .ZN(n10099) );
  NAND2_X1 U11866 ( .A1(n10781), .A2(n10099), .ZN(n10100) );
  MUX2_X1 U11867 ( .A(n10102), .B(n10115), .S(n15978), .Z(n10104) );
  INV_X1 U11868 ( .A(n10103), .ZN(n13057) );
  NAND2_X1 U11869 ( .A1(n10104), .A2(n8136), .ZN(P3_U3456) );
  NAND2_X1 U11870 ( .A1(n10895), .A2(n10783), .ZN(n10107) );
  NAND2_X1 U11871 ( .A1(n10107), .A2(n10106), .ZN(n10114) );
  XNOR2_X1 U11872 ( .A(n13392), .B(n10108), .ZN(n10110) );
  NAND2_X1 U11873 ( .A1(n10318), .A2(n10286), .ZN(n10896) );
  INV_X1 U11874 ( .A(n10895), .ZN(n10111) );
  NAND2_X1 U11875 ( .A1(n10896), .A2(n10111), .ZN(n10112) );
  NAND2_X1 U11876 ( .A1(n10112), .A2(n13392), .ZN(n10113) );
  MUX2_X1 U11877 ( .A(n10116), .B(n10115), .S(n15839), .Z(n10117) );
  NAND2_X1 U11878 ( .A1(n10117), .A2(n8137), .ZN(P3_U3488) );
  INV_X1 U11879 ( .A(n10118), .ZN(n10119) );
  NAND2_X1 U11880 ( .A1(n10120), .A2(n10119), .ZN(n10123) );
  NAND2_X1 U11881 ( .A1(n10121), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U11882 ( .A1(n10123), .A2(n10122), .ZN(n10142) );
  XNOR2_X1 U11883 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n10140) );
  NAND2_X1 U11884 ( .A1(n10142), .A2(n10140), .ZN(n10126) );
  INV_X1 U11885 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U11886 ( .A1(n10124), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U11887 ( .A1(n10126), .A2(n10125), .ZN(n10129) );
  INV_X1 U11888 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10127) );
  XNOR2_X1 U11889 ( .A(n10127), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n10128) );
  XNOR2_X1 U11890 ( .A(n10129), .B(n10128), .ZN(n13395) );
  NAND2_X1 U11891 ( .A1(n13395), .A2(n10130), .ZN(n10132) );
  NAND2_X1 U11892 ( .A1(n10143), .A2(SI_31_), .ZN(n10131) );
  NAND2_X1 U11893 ( .A1(n10132), .A2(n10131), .ZN(n10148) );
  NAND2_X1 U11894 ( .A1(n10012), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U11895 ( .A1(n10133), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U11896 ( .A1(n9667), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10134) );
  AND3_X1 U11897 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(n10137) );
  AND2_X1 U11898 ( .A1(n10138), .A2(n10137), .ZN(n13048) );
  OR2_X1 U11899 ( .A1(n10148), .A2(n13048), .ZN(n10277) );
  NAND2_X1 U11900 ( .A1(n10277), .A2(n10139), .ZN(n10284) );
  INV_X1 U11901 ( .A(n10140), .ZN(n10141) );
  XNOR2_X1 U11902 ( .A(n10142), .B(n10141), .ZN(n13400) );
  NAND2_X1 U11903 ( .A1(n13400), .A2(n10130), .ZN(n10145) );
  NAND2_X1 U11904 ( .A1(n10143), .A2(SI_30_), .ZN(n10144) );
  INV_X1 U11905 ( .A(n15975), .ZN(n13053) );
  INV_X1 U11906 ( .A(n13048), .ZN(n12904) );
  NAND2_X1 U11907 ( .A1(n15975), .A2(n11032), .ZN(n10279) );
  OAI21_X1 U11908 ( .B1(n13053), .B2(n12904), .A(n10279), .ZN(n10146) );
  NOR2_X1 U11909 ( .A1(n13319), .A2(n12904), .ZN(n10313) );
  NOR2_X1 U11910 ( .A1(n15975), .A2(n11032), .ZN(n10276) );
  INV_X1 U11911 ( .A(n10150), .ZN(n10151) );
  INV_X1 U11912 ( .A(n10152), .ZN(n10153) );
  AOI21_X1 U11913 ( .B1(n10155), .B2(n10154), .A(n10153), .ZN(n10159) );
  INV_X1 U11914 ( .A(n10156), .ZN(n10157) );
  AOI21_X1 U11915 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(n10263) );
  NAND2_X1 U11916 ( .A1(n10042), .A2(n15127), .ZN(n10294) );
  AND2_X1 U11917 ( .A1(n10160), .A2(n10294), .ZN(n10164) );
  INV_X1 U11918 ( .A(n10164), .ZN(n10162) );
  NAND2_X1 U11919 ( .A1(n10162), .A2(n10161), .ZN(n10167) );
  AOI21_X1 U11920 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(n10166) );
  MUX2_X1 U11921 ( .A(n10167), .B(n10166), .S(n10285), .Z(n10170) );
  INV_X1 U11922 ( .A(n10176), .ZN(n10168) );
  AOI21_X1 U11923 ( .B1(n15546), .B2(n15580), .A(n10168), .ZN(n10169) );
  OAI22_X1 U11924 ( .A1(n10170), .A2(n15572), .B1(n10169), .B2(n10285), .ZN(
        n10174) );
  AOI21_X1 U11925 ( .B1(n10173), .B2(n10171), .A(n10286), .ZN(n10172) );
  AOI21_X1 U11926 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10181) );
  OAI21_X1 U11927 ( .B1(n10286), .B2(n10176), .A(n10175), .ZN(n10180) );
  NAND2_X1 U11928 ( .A1(n12922), .A2(n11189), .ZN(n10178) );
  MUX2_X1 U11929 ( .A(n10178), .B(n10177), .S(n10285), .Z(n10179) );
  OAI211_X1 U11930 ( .C1(n10181), .C2(n10180), .A(n11679), .B(n10179), .ZN(
        n10186) );
  MUX2_X1 U11931 ( .A(n10183), .B(n10182), .S(n10286), .Z(n10184) );
  NAND3_X1 U11932 ( .A1(n10186), .A2(n10185), .A3(n10184), .ZN(n10190) );
  MUX2_X1 U11933 ( .A(n10188), .B(n10187), .S(n10285), .Z(n10189) );
  NAND3_X1 U11934 ( .A1(n10190), .A2(n11664), .A3(n10189), .ZN(n10194) );
  NAND2_X1 U11935 ( .A1(n15701), .A2(n10286), .ZN(n10192) );
  NAND2_X1 U11936 ( .A1(n11649), .A2(n10285), .ZN(n10191) );
  MUX2_X1 U11937 ( .A(n10192), .B(n10191), .S(n12919), .Z(n10193) );
  NAND3_X1 U11938 ( .A1(n10194), .A2(n11796), .A3(n10193), .ZN(n10198) );
  OR2_X1 U11939 ( .A1(n7664), .A2(n10199), .ZN(n10296) );
  INV_X1 U11940 ( .A(n10296), .ZN(n11858) );
  MUX2_X1 U11941 ( .A(n10196), .B(n10195), .S(n10285), .Z(n10197) );
  NAND3_X1 U11942 ( .A1(n10198), .A2(n11858), .A3(n10197), .ZN(n10203) );
  INV_X1 U11943 ( .A(n10199), .ZN(n10200) );
  MUX2_X1 U11944 ( .A(n10201), .B(n10200), .S(n10286), .Z(n10202) );
  NAND3_X1 U11945 ( .A1(n10203), .A2(n8111), .A3(n10202), .ZN(n10207) );
  MUX2_X1 U11946 ( .A(n10205), .B(n10204), .S(n10285), .Z(n10206) );
  INV_X1 U11947 ( .A(n12138), .ZN(n11992) );
  AOI21_X1 U11948 ( .B1(n10207), .B2(n10206), .A(n11992), .ZN(n10215) );
  NAND2_X1 U11949 ( .A1(n10213), .A2(n10208), .ZN(n10209) );
  OAI211_X1 U11950 ( .C1(n10215), .C2(n10209), .A(n10285), .B(n10212), .ZN(
        n10211) );
  NOR2_X1 U11951 ( .A1(n12780), .A2(n10286), .ZN(n10210) );
  AOI22_X1 U11952 ( .A1(n10211), .A2(n12350), .B1(n10210), .B2(n12738), .ZN(
        n10223) );
  NAND2_X1 U11953 ( .A1(n12172), .A2(n10212), .ZN(n10214) );
  OAI211_X1 U11954 ( .C1(n10215), .C2(n10214), .A(n10286), .B(n10213), .ZN(
        n10216) );
  NAND2_X1 U11955 ( .A1(n10216), .A2(n12267), .ZN(n10222) );
  INV_X1 U11956 ( .A(n10217), .ZN(n10220) );
  XNOR2_X1 U11957 ( .A(n10218), .B(n10286), .ZN(n10219) );
  OAI21_X1 U11958 ( .B1(n9843), .B2(n10220), .A(n10219), .ZN(n10221) );
  OAI211_X1 U11959 ( .C1(n10223), .C2(n10222), .A(n12334), .B(n10221), .ZN(
        n10227) );
  MUX2_X1 U11960 ( .A(n10225), .B(n10224), .S(n10285), .Z(n10226) );
  NAND3_X1 U11961 ( .A1(n10227), .A2(n13245), .A3(n10226), .ZN(n10232) );
  AND2_X1 U11962 ( .A1(n10236), .A2(n10228), .ZN(n10229) );
  MUX2_X1 U11963 ( .A(n10230), .B(n10229), .S(n10286), .Z(n10231) );
  NAND4_X1 U11964 ( .A1(n10232), .A2(n13229), .A3(n10235), .A4(n10231), .ZN(
        n10246) );
  INV_X1 U11965 ( .A(n10236), .ZN(n10234) );
  OAI211_X1 U11966 ( .C1(n10234), .C2(n10233), .A(n10243), .B(n10235), .ZN(
        n10241) );
  INV_X1 U11967 ( .A(n10235), .ZN(n10239) );
  INV_X1 U11968 ( .A(n10292), .ZN(n10237) );
  OAI211_X1 U11969 ( .C1(n10239), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10240) );
  MUX2_X1 U11970 ( .A(n10241), .B(n10240), .S(n10285), .Z(n10242) );
  INV_X1 U11971 ( .A(n10242), .ZN(n10245) );
  INV_X1 U11972 ( .A(n10243), .ZN(n10293) );
  MUX2_X1 U11973 ( .A(n10292), .B(n10293), .S(n10285), .Z(n10244) );
  AOI211_X1 U11974 ( .C1(n10246), .C2(n10245), .A(n10244), .B(n7672), .ZN(
        n10255) );
  MUX2_X1 U11975 ( .A(n10248), .B(n10247), .S(n10286), .Z(n10252) );
  MUX2_X1 U11976 ( .A(n10250), .B(n7669), .S(n10285), .Z(n10251) );
  AOI21_X1 U11977 ( .B1(n13169), .B2(n10252), .A(n10251), .ZN(n10254) );
  INV_X1 U11978 ( .A(n10253), .ZN(n10256) );
  AOI211_X1 U11979 ( .C1(n10255), .C2(n13169), .A(n10254), .B(n13155), .ZN(
        n10259) );
  MUX2_X1 U11980 ( .A(n10257), .B(n10256), .S(n10286), .Z(n10258) );
  OR3_X1 U11981 ( .A1(n10259), .A2(n10258), .A3(n13149), .ZN(n10267) );
  INV_X1 U11982 ( .A(n10262), .ZN(n10265) );
  OAI21_X1 U11983 ( .B1(n10265), .B2(n10264), .A(n10263), .ZN(n10269) );
  NAND3_X1 U11984 ( .A1(n10267), .A2(n10306), .A3(n10266), .ZN(n10268) );
  NAND2_X1 U11985 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  MUX2_X1 U11986 ( .A(n10274), .B(n10273), .S(n10286), .Z(n10275) );
  INV_X1 U11987 ( .A(n10276), .ZN(n10278) );
  AND2_X1 U11988 ( .A1(n10278), .A2(n10279), .ZN(n10309) );
  INV_X1 U11989 ( .A(n10277), .ZN(n10311) );
  NAND2_X1 U11990 ( .A1(n10278), .A2(n10286), .ZN(n10280) );
  NAND2_X1 U11991 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  AOI211_X1 U11992 ( .C1(n10283), .C2(n10282), .A(n10311), .B(n10281), .ZN(
        n10291) );
  INV_X1 U11993 ( .A(n10284), .ZN(n10287) );
  INV_X1 U11994 ( .A(n10316), .ZN(n10319) );
  OR2_X1 U11995 ( .A1(n10293), .A2(n10292), .ZN(n13196) );
  INV_X1 U11996 ( .A(n13196), .ZN(n13203) );
  INV_X1 U11997 ( .A(n11679), .ZN(n11681) );
  INV_X1 U11998 ( .A(n10294), .ZN(n10295) );
  OR2_X1 U11999 ( .A1(n10295), .A2(n15544), .ZN(n15130) );
  NOR4_X1 U12000 ( .A1(n11681), .A2(n11732), .A3(n15130), .A4(n15549), .ZN(
        n10298) );
  NOR2_X1 U12001 ( .A1(n10296), .A2(n11661), .ZN(n10297) );
  NAND4_X1 U12002 ( .A1(n10298), .A2(n11528), .A3(n11796), .A4(n10297), .ZN(
        n10299) );
  NOR4_X1 U12003 ( .A1(n10299), .A2(n7634), .A3(n15572), .A4(n11897), .ZN(
        n10300) );
  NAND4_X1 U12004 ( .A1(n10300), .A2(n12138), .A3(n12175), .A4(n12350), .ZN(
        n10301) );
  NOR3_X1 U12005 ( .A1(n10301), .A2(n9843), .A3(n12329), .ZN(n10302) );
  NAND3_X1 U12006 ( .A1(n13203), .A2(n13245), .A3(n10302), .ZN(n10304) );
  NAND4_X1 U12007 ( .A1(n13136), .A2(n13169), .A3(n13185), .A4(n13153), .ZN(
        n10303) );
  NOR4_X1 U12008 ( .A1(n10305), .A2(n13223), .A3(n10304), .A4(n10303), .ZN(
        n10308) );
  NAND4_X1 U12009 ( .A1(n10308), .A2(n10018), .A3(n10307), .A4(n10306), .ZN(
        n10312) );
  INV_X1 U12010 ( .A(n10309), .ZN(n10310) );
  NOR4_X1 U12011 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10314) );
  XNOR2_X1 U12012 ( .A(n10314), .B(n7209), .ZN(n10315) );
  OAI22_X1 U12013 ( .A1(n10316), .A2(n11526), .B1(n10761), .B2(n10315), .ZN(
        n10317) );
  INV_X2 U12014 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR2_X1 U12015 ( .A1(n10899), .A2(n10782), .ZN(n10785) );
  NOR3_X1 U12016 ( .A1(n10785), .A2(n7384), .A3(n12134), .ZN(n10322) );
  OAI21_X1 U12017 ( .B1(n11357), .B2(n11176), .A(P3_B_REG_SCAN_IN), .ZN(n10321) );
  OR2_X1 U12018 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  NOR2_X1 U12019 ( .A1(n10347), .A2(P1_U3086), .ZN(n10324) );
  AND2_X2 U12020 ( .A1(n10324), .A2(n10623), .ZN(P1_U4016) );
  INV_X1 U12021 ( .A(n12257), .ZN(n10325) );
  INV_X1 U12022 ( .A(n10773), .ZN(n10327) );
  NAND2_X1 U12023 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10336) );
  INV_X1 U12024 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10328) );
  MUX2_X1 U12025 ( .A(n10328), .B(P2_REG2_REG_1__SCAN_IN), .S(n10594), .Z(
        n10335) );
  OR2_X1 U12026 ( .A1(n10335), .A2(n10336), .ZN(n13822) );
  INV_X1 U12027 ( .A(n13822), .ZN(n10334) );
  NAND2_X1 U12028 ( .A1(n10720), .A2(n12257), .ZN(n10330) );
  NAND2_X1 U12029 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  NAND2_X1 U12030 ( .A1(n10332), .A2(n10331), .ZN(n10342) );
  NOR2_X1 U12031 ( .A1(n10341), .A2(P2_U3088), .ZN(n14228) );
  AND2_X1 U12032 ( .A1(n10342), .A2(n14228), .ZN(n10338) );
  INV_X1 U12033 ( .A(n14231), .ZN(n10333) );
  AND2_X1 U12034 ( .A1(n10338), .A2(n10333), .ZN(n15205) );
  AOI211_X1 U12035 ( .C1(n10336), .C2(n10335), .A(n10334), .B(n15180), .ZN(
        n10346) );
  INV_X1 U12036 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10977) );
  MUX2_X1 U12037 ( .A(n10977), .B(P2_REG1_REG_1__SCAN_IN), .S(n10594), .Z(
        n10340) );
  INV_X1 U12038 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10337) );
  INV_X1 U12039 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10988) );
  OR2_X1 U12040 ( .A1(n10337), .A2(n10988), .ZN(n10339) );
  NOR3_X1 U12041 ( .A1(n10340), .A2(n10988), .A3(n10337), .ZN(n13829) );
  INV_X1 U12042 ( .A(n15201), .ZN(n11089) );
  AOI211_X1 U12043 ( .C1(n10340), .C2(n10339), .A(n13829), .B(n11089), .ZN(
        n10345) );
  AND2_X1 U12044 ( .A1(n10342), .A2(n10341), .ZN(n15141) );
  INV_X1 U12045 ( .A(n10594), .ZN(n10587) );
  NOR2_X1 U12046 ( .A1(n15158), .A2(n10587), .ZN(n10344) );
  OR2_X1 U12047 ( .A1(n10342), .A2(P2_U3088), .ZN(n15198) );
  INV_X1 U12048 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11311) );
  OAI22_X1 U12049 ( .A1(n15198), .A2(n7412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11311), .ZN(n10343) );
  OR4_X1 U12050 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        P2_U3215) );
  NAND2_X1 U12051 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14390) );
  AND2_X4 U12052 ( .A1(n10347), .A2(n10909), .ZN(n10994) );
  INV_X1 U12053 ( .A(n10347), .ZN(n10351) );
  MUX2_X1 U12054 ( .A(n14390), .B(n10627), .S(n14886), .Z(n10357) );
  INV_X1 U12055 ( .A(n9500), .ZN(n10629) );
  OAI21_X1 U12056 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14886), .A(n10629), .ZN(
        n14377) );
  NAND2_X1 U12057 ( .A1(n14377), .A2(n8937), .ZN(n10356) );
  OAI211_X1 U12058 ( .C1(n10357), .C2(n9500), .A(P1_U4016), .B(n10356), .ZN(
        n14408) );
  INV_X1 U12059 ( .A(n14408), .ZN(n10389) );
  INV_X1 U12060 ( .A(n10623), .ZN(n10358) );
  OAI21_X1 U12061 ( .B1(n10347), .B2(n10358), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n10364) );
  NAND2_X1 U12062 ( .A1(n10359), .A2(n10623), .ZN(n10361) );
  NAND2_X1 U12063 ( .A1(n10361), .A2(n10360), .ZN(n10363) );
  INV_X1 U12064 ( .A(n10363), .ZN(n10362) );
  INV_X1 U12065 ( .A(n14886), .ZN(n14560) );
  NAND2_X1 U12066 ( .A1(n10629), .A2(n14560), .ZN(n10365) );
  NOR2_X2 U12067 ( .A1(n10383), .A2(n10365), .ZN(n14553) );
  INV_X1 U12068 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10366) );
  MUX2_X1 U12069 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10366), .S(n14397), .Z(
        n10370) );
  MUX2_X1 U12070 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10367), .S(n14386), .Z(
        n14391) );
  AND2_X1 U12071 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10368) );
  NAND2_X1 U12072 ( .A1(n14391), .A2(n10368), .ZN(n14399) );
  NAND2_X1 U12073 ( .A1(n14386), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U12074 ( .A1(n14399), .A2(n14398), .ZN(n10369) );
  NAND2_X1 U12075 ( .A1(n10370), .A2(n10369), .ZN(n14416) );
  NAND2_X1 U12076 ( .A1(n14397), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14415) );
  NAND2_X1 U12077 ( .A1(n14416), .A2(n14415), .ZN(n10372) );
  INV_X1 U12078 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14414) );
  MUX2_X1 U12079 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14414), .S(n14413), .Z(
        n10371) );
  NAND2_X1 U12080 ( .A1(n10372), .A2(n10371), .ZN(n14419) );
  NAND2_X1 U12081 ( .A1(n14413), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U12082 ( .A1(n14419), .A2(n10376), .ZN(n10375) );
  INV_X1 U12083 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U12084 ( .A(n10373), .B(P1_REG2_REG_4__SCAN_IN), .S(n10461), .Z(
        n10374) );
  NAND2_X1 U12085 ( .A1(n10375), .A2(n10374), .ZN(n10471) );
  MUX2_X1 U12086 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10373), .S(n10461), .Z(
        n10377) );
  NAND3_X1 U12087 ( .A1(n10377), .A2(n14419), .A3(n10376), .ZN(n10378) );
  NAND3_X1 U12088 ( .A1(n14553), .A2(n10471), .A3(n10378), .ZN(n10379) );
  NAND2_X1 U12089 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n11439) );
  OAI211_X1 U12090 ( .C1(n15240), .C2(n14557), .A(n10379), .B(n11439), .ZN(
        n10388) );
  NOR2_X1 U12091 ( .A1(n10383), .A2(n10629), .ZN(n14551) );
  INV_X1 U12092 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11252) );
  MUX2_X1 U12093 ( .A(n11252), .B(P1_REG1_REG_4__SCAN_IN), .S(n10461), .Z(
        n10385) );
  INV_X1 U12094 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15600) );
  MUX2_X1 U12095 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n15600), .S(n14397), .Z(
        n14404) );
  INV_X1 U12096 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15570) );
  MUX2_X1 U12097 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15570), .S(n14386), .Z(
        n14389) );
  AND2_X1 U12098 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14388) );
  NAND2_X1 U12099 ( .A1(n14389), .A2(n14388), .ZN(n14387) );
  NAND2_X1 U12100 ( .A1(n14386), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U12101 ( .A1(n14387), .A2(n10380), .ZN(n14403) );
  NAND2_X1 U12102 ( .A1(n14404), .A2(n14403), .ZN(n14402) );
  NAND2_X1 U12103 ( .A1(n14397), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10381) );
  NAND2_X1 U12104 ( .A1(n14402), .A2(n10381), .ZN(n14410) );
  INV_X1 U12105 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15624) );
  MUX2_X1 U12106 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n15624), .S(n14413), .Z(
        n14411) );
  NAND2_X1 U12107 ( .A1(n14410), .A2(n14411), .ZN(n14409) );
  NAND2_X1 U12108 ( .A1(n14413), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U12109 ( .A1(n14409), .A2(n10382), .ZN(n10384) );
  INV_X1 U12110 ( .A(n10383), .ZN(n14379) );
  NAND2_X1 U12111 ( .A1(n14379), .A2(n14886), .ZN(n14548) );
  NAND2_X1 U12112 ( .A1(n10384), .A2(n10385), .ZN(n10463) );
  OAI211_X1 U12113 ( .C1(n10385), .C2(n10384), .A(n14546), .B(n10463), .ZN(
        n10386) );
  OAI21_X1 U12114 ( .B1(n14518), .B2(n10461), .A(n10386), .ZN(n10387) );
  OR3_X1 U12115 ( .A1(n10389), .A2(n10388), .A3(n10387), .ZN(P1_U3247) );
  NOR2_X1 U12116 ( .A1(n10397), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13397) );
  INV_X2 U12117 ( .A(n13397), .ZN(n13403) );
  INV_X2 U12118 ( .A(n11355), .ZN(n13402) );
  INV_X1 U12119 ( .A(n10390), .ZN(n10391) );
  OAI222_X1 U12120 ( .A1(P3_U3151), .A2(n10954), .B1(n13403), .B2(n14953), 
        .C1(n13402), .C2(n10391), .ZN(P3_U3294) );
  INV_X1 U12121 ( .A(SI_8_), .ZN(n10394) );
  INV_X1 U12122 ( .A(n10392), .ZN(n10393) );
  OAI222_X1 U12123 ( .A1(P3_U3151), .A2(n12972), .B1(n13403), .B2(n10394), 
        .C1(n13402), .C2(n10393), .ZN(P3_U3287) );
  OAI222_X1 U12124 ( .A1(P3_U3151), .A2(n11155), .B1(n13403), .B2(n15062), 
        .C1(n13402), .C2(n10395), .ZN(P3_U3288) );
  OAI222_X1 U12125 ( .A1(P3_U3151), .A2(n12975), .B1(n13403), .B2(n14910), 
        .C1(n13402), .C2(n10396), .ZN(P3_U3286) );
  INV_X1 U12126 ( .A(n14234), .ZN(n14244) );
  OAI222_X1 U12127 ( .A1(n14244), .A2(n10399), .B1(n14239), .B2(n10415), .C1(
        n10587), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U12128 ( .A(n10400), .ZN(n10402) );
  OAI222_X1 U12129 ( .A1(P3_U3151), .A2(n11056), .B1(n13402), .B2(n10402), 
        .C1(n10401), .C2(n13403), .ZN(P3_U3289) );
  INV_X1 U12130 ( .A(n10875), .ZN(n10819) );
  OAI222_X1 U12131 ( .A1(n10819), .A2(P3_U3151), .B1(n13402), .B2(n10404), 
        .C1(n10403), .C2(n13403), .ZN(P3_U3291) );
  INV_X1 U12132 ( .A(n10892), .ZN(n10833) );
  OAI222_X1 U12133 ( .A1(n10833), .A2(P3_U3151), .B1(n13402), .B2(n10405), 
        .C1(n15075), .C2(n13403), .ZN(P3_U3293) );
  OAI222_X1 U12134 ( .A1(n10927), .A2(P3_U3151), .B1(n13402), .B2(n10407), 
        .C1(n10406), .C2(n13403), .ZN(P3_U3290) );
  OAI222_X1 U12135 ( .A1(n10835), .A2(P3_U3151), .B1(n13402), .B2(n10409), 
        .C1(n10408), .C2(n13403), .ZN(P3_U3292) );
  OAI222_X1 U12136 ( .A1(P3_U3151), .A2(n12971), .B1(n13403), .B2(n14909), 
        .C1(n13402), .C2(n10410), .ZN(P3_U3285) );
  OAI222_X1 U12137 ( .A1(n12978), .A2(P3_U3151), .B1(n13402), .B2(n10411), 
        .C1(n13403), .C2(n15057), .ZN(P3_U3284) );
  INV_X1 U12138 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10413) );
  OAI222_X1 U12139 ( .A1(n14897), .A2(n10413), .B1(n14893), .B2(n7907), .C1(
        n10461), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12140 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10414) );
  OAI222_X1 U12141 ( .A1(P1_U3086), .A2(n8926), .B1(n14893), .B2(n10415), .C1(
        n10414), .C2(n14897), .ZN(P1_U3354) );
  INV_X1 U12142 ( .A(n14397), .ZN(n10416) );
  OAI222_X1 U12143 ( .A1(n14897), .A2(n10417), .B1(n14893), .B2(n10423), .C1(
        n10416), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U12144 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10420) );
  INV_X1 U12145 ( .A(n14413), .ZN(n10419) );
  OAI222_X1 U12146 ( .A1(n14897), .A2(n10420), .B1(n14893), .B2(n8914), .C1(
        n10419), .C2(P1_U3086), .ZN(P1_U3352) );
  AOI22_X1 U12147 ( .A1(n13836), .A2(P2_STATE_REG_SCAN_IN), .B1(n14234), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n10421) );
  OAI21_X1 U12148 ( .B1(n8914), .B2(n14239), .A(n10421), .ZN(P2_U3324) );
  INV_X1 U12149 ( .A(n10646), .ZN(n10605) );
  OAI222_X1 U12150 ( .A1(n14244), .A2(n10422), .B1(n14239), .B2(n7907), .C1(
        n10605), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U12151 ( .A(n13824), .ZN(n10596) );
  OAI222_X1 U12152 ( .A1(n14244), .A2(n10424), .B1(n14239), .B2(n10423), .C1(
        n10596), .C2(P2_U3088), .ZN(P2_U3325) );
  OAI222_X1 U12153 ( .A1(n15433), .A2(P3_U3151), .B1(n13402), .B2(n10425), 
        .C1(n13403), .C2(n15053), .ZN(P3_U3283) );
  INV_X1 U12154 ( .A(n10426), .ZN(n10428) );
  OAI222_X1 U12155 ( .A1(n14244), .A2(n10427), .B1(n14239), .B2(n10428), .C1(
        n10676), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U12156 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10429) );
  INV_X1 U12157 ( .A(n10523), .ZN(n10515) );
  OAI222_X1 U12158 ( .A1(n14897), .A2(n10429), .B1(n14893), .B2(n10428), .C1(
        n10515), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U12159 ( .A(n10648), .ZN(n15142) );
  OAI222_X1 U12160 ( .A1(n14244), .A2(n10430), .B1(n14239), .B2(n10432), .C1(
        n15142), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12161 ( .A(n14430), .ZN(n10431) );
  OAI222_X1 U12162 ( .A1(n14897), .A2(n10433), .B1(n14893), .B2(n10432), .C1(
        n10431), .C2(P1_U3086), .ZN(P1_U3349) );
  AOI22_X1 U12163 ( .A1(n14449), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14880), .ZN(n10434) );
  OAI21_X1 U12164 ( .B1(n10435), .B2(n14893), .A(n10434), .ZN(P1_U3348) );
  INV_X1 U12165 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10436) );
  INV_X1 U12166 ( .A(n10683), .ZN(n10658) );
  OAI222_X1 U12167 ( .A1(n14244), .A2(n10436), .B1(n14239), .B2(n10435), .C1(
        n10658), .C2(P2_U3088), .ZN(P2_U3320) );
  OAI222_X1 U12168 ( .A1(P3_U3151), .A2(n12982), .B1(n13403), .B2(n10438), 
        .C1(n13402), .C2(n10437), .ZN(P3_U3282) );
  NAND3_X1 U12169 ( .A1(n10439), .A2(P1_B_REG_SCAN_IN), .A3(n10440), .ZN(
        n10444) );
  INV_X1 U12170 ( .A(n10440), .ZN(n10442) );
  AOI21_X1 U12171 ( .B1(n10442), .B2(n10441), .A(n14889), .ZN(n10443) );
  INV_X1 U12172 ( .A(n10618), .ZN(n10445) );
  NAND2_X1 U12173 ( .A1(n10634), .A2(n10445), .ZN(n14901) );
  INV_X1 U12174 ( .A(n14901), .ZN(n10447) );
  INV_X1 U12175 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U12176 ( .A1(n10439), .A2(n14889), .ZN(n11212) );
  NAND2_X1 U12177 ( .A1(n10447), .A2(n11212), .ZN(n10446) );
  OAI21_X1 U12178 ( .B1(n10447), .B2(n10616), .A(n10446), .ZN(P1_U3446) );
  OAI222_X1 U12179 ( .A1(n12970), .A2(P3_U3151), .B1(n13402), .B2(n10448), 
        .C1(n13403), .C2(n14943), .ZN(P3_U3281) );
  AOI22_X1 U12180 ( .A1(n14464), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14880), .ZN(n10449) );
  OAI21_X1 U12181 ( .B1(n10455), .B2(n14893), .A(n10449), .ZN(P1_U3346) );
  INV_X1 U12182 ( .A(n10450), .ZN(n10452) );
  INV_X1 U12183 ( .A(n10554), .ZN(n10543) );
  OAI222_X1 U12184 ( .A1(n14897), .A2(n10451), .B1(n14893), .B2(n10452), .C1(
        P1_U3086), .C2(n10543), .ZN(P1_U3347) );
  INV_X1 U12185 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10453) );
  INV_X1 U12186 ( .A(n10752), .ZN(n10691) );
  OAI222_X1 U12187 ( .A1(n14244), .A2(n10453), .B1(n14239), .B2(n10452), .C1(
        P2_U3088), .C2(n10691), .ZN(P2_U3319) );
  INV_X1 U12188 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10456) );
  INV_X1 U12189 ( .A(n13860), .ZN(n10454) );
  OAI222_X1 U12190 ( .A1(n14244), .A2(n10456), .B1(n14239), .B2(n10455), .C1(
        n10454), .C2(P2_U3088), .ZN(P2_U3318) );
  OAI222_X1 U12191 ( .A1(n15490), .A2(P3_U3151), .B1(n13402), .B2(n10457), 
        .C1(n13403), .C2(n15046), .ZN(P3_U3280) );
  AOI22_X1 U12192 ( .A1(n14479), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14880), .ZN(n10458) );
  OAI21_X1 U12193 ( .B1(n10460), .B2(n14893), .A(n10458), .ZN(P1_U3345) );
  INV_X1 U12194 ( .A(n11078), .ZN(n11072) );
  INV_X1 U12195 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10459) );
  OAI222_X1 U12196 ( .A1(P2_U3088), .A2(n11072), .B1(n14239), .B2(n10460), 
        .C1(n10459), .C2(n14244), .ZN(P2_U3317) );
  INV_X1 U12197 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10514) );
  XNOR2_X1 U12198 ( .A(n10523), .B(n10514), .ZN(n10465) );
  INV_X1 U12199 ( .A(n10461), .ZN(n10466) );
  NAND2_X1 U12200 ( .A1(n10466), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10462) );
  AND2_X1 U12201 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  NAND2_X1 U12202 ( .A1(n10464), .A2(n10465), .ZN(n10517) );
  OAI21_X1 U12203 ( .B1(n10465), .B2(n10464), .A(n10517), .ZN(n10475) );
  NAND2_X1 U12204 ( .A1(n10466), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U12205 ( .A1(n10471), .A2(n10470), .ZN(n10469) );
  INV_X1 U12206 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10467) );
  MUX2_X1 U12207 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10467), .S(n10523), .Z(
        n10468) );
  NAND2_X1 U12208 ( .A1(n10469), .A2(n10468), .ZN(n14433) );
  MUX2_X1 U12209 ( .A(n10467), .B(P1_REG2_REG_5__SCAN_IN), .S(n10523), .Z(
        n10472) );
  NAND3_X1 U12210 ( .A1(n10472), .A2(n10471), .A3(n10470), .ZN(n10473) );
  AND3_X1 U12211 ( .A1(n14553), .A2(n14433), .A3(n10473), .ZN(n10474) );
  AOI21_X1 U12212 ( .B1(n14546), .B2(n10475), .A(n10474), .ZN(n10478) );
  INV_X1 U12213 ( .A(n14557), .ZN(n14521) );
  AND2_X1 U12214 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10476) );
  AOI21_X1 U12215 ( .B1(n14521), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10476), .ZN(
        n10477) );
  OAI211_X1 U12216 ( .C1(n10515), .C2(n14518), .A(n10478), .B(n10477), .ZN(
        P1_U3248) );
  INV_X1 U12217 ( .A(n13393), .ZN(n10479) );
  NOR2_X1 U12218 ( .A1(n10479), .A2(n7229), .ZN(n10483) );
  INV_X1 U12219 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10480) );
  NOR2_X1 U12220 ( .A1(n10505), .A2(n10480), .ZN(P3_U3240) );
  INV_X1 U12221 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10481) );
  NOR2_X1 U12222 ( .A1(n10483), .A2(n10481), .ZN(P3_U3260) );
  INV_X1 U12223 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10482) );
  NOR2_X1 U12224 ( .A1(n10483), .A2(n10482), .ZN(P3_U3262) );
  INV_X1 U12225 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10484) );
  NOR2_X1 U12226 ( .A1(n10505), .A2(n10484), .ZN(P3_U3254) );
  INV_X1 U12227 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10485) );
  NOR2_X1 U12228 ( .A1(n10483), .A2(n10485), .ZN(P3_U3258) );
  INV_X1 U12229 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10486) );
  NOR2_X1 U12230 ( .A1(n10505), .A2(n10486), .ZN(P3_U3256) );
  INV_X1 U12231 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10487) );
  NOR2_X1 U12232 ( .A1(n10483), .A2(n10487), .ZN(P3_U3244) );
  INV_X1 U12233 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10488) );
  NOR2_X1 U12234 ( .A1(n10505), .A2(n10488), .ZN(P3_U3253) );
  INV_X1 U12235 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10489) );
  NOR2_X1 U12236 ( .A1(n10505), .A2(n10489), .ZN(P3_U3252) );
  INV_X1 U12237 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10490) );
  NOR2_X1 U12238 ( .A1(n10505), .A2(n10490), .ZN(P3_U3257) );
  INV_X1 U12239 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10491) );
  NOR2_X1 U12240 ( .A1(n10505), .A2(n10491), .ZN(P3_U3246) );
  INV_X1 U12241 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10492) );
  NOR2_X1 U12242 ( .A1(n10505), .A2(n10492), .ZN(P3_U3255) );
  INV_X1 U12243 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10493) );
  NOR2_X1 U12244 ( .A1(n10505), .A2(n10493), .ZN(P3_U3251) );
  INV_X1 U12245 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10494) );
  NOR2_X1 U12246 ( .A1(n10505), .A2(n10494), .ZN(P3_U3259) );
  INV_X1 U12247 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10495) );
  NOR2_X1 U12248 ( .A1(n10483), .A2(n10495), .ZN(P3_U3239) );
  INV_X1 U12249 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10496) );
  NOR2_X1 U12250 ( .A1(n10483), .A2(n10496), .ZN(P3_U3237) );
  INV_X1 U12251 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10497) );
  NOR2_X1 U12252 ( .A1(n10483), .A2(n10497), .ZN(P3_U3241) );
  INV_X1 U12253 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10498) );
  NOR2_X1 U12254 ( .A1(n10483), .A2(n10498), .ZN(P3_U3242) );
  INV_X1 U12255 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10499) );
  NOR2_X1 U12256 ( .A1(n10505), .A2(n10499), .ZN(P3_U3250) );
  INV_X1 U12257 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10500) );
  NOR2_X1 U12258 ( .A1(n10505), .A2(n10500), .ZN(P3_U3261) );
  INV_X1 U12259 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10501) );
  NOR2_X1 U12260 ( .A1(n10505), .A2(n10501), .ZN(P3_U3263) );
  INV_X1 U12261 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10502) );
  NOR2_X1 U12262 ( .A1(n10505), .A2(n10502), .ZN(P3_U3249) );
  INV_X1 U12263 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10503) );
  NOR2_X1 U12264 ( .A1(n10505), .A2(n10503), .ZN(P3_U3248) );
  INV_X1 U12265 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10504) );
  NOR2_X1 U12266 ( .A1(n10505), .A2(n10504), .ZN(P3_U3247) );
  INV_X1 U12267 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10506) );
  NOR2_X1 U12268 ( .A1(n10483), .A2(n10506), .ZN(P3_U3238) );
  INV_X1 U12269 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10507) );
  NOR2_X1 U12270 ( .A1(n10483), .A2(n10507), .ZN(P3_U3245) );
  INV_X1 U12271 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10508) );
  NOR2_X1 U12272 ( .A1(n10483), .A2(n10508), .ZN(P3_U3234) );
  INV_X1 U12273 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10509) );
  NOR2_X1 U12274 ( .A1(n10505), .A2(n10509), .ZN(P3_U3235) );
  INV_X1 U12275 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10510) );
  NOR2_X1 U12276 ( .A1(n10505), .A2(n10510), .ZN(P3_U3236) );
  INV_X1 U12277 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10511) );
  NOR2_X1 U12278 ( .A1(n10505), .A2(n10511), .ZN(P3_U3243) );
  INV_X1 U12279 ( .A(n10512), .ZN(n10570) );
  AOI22_X1 U12280 ( .A1(n14496), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n14880), .ZN(n10513) );
  OAI21_X1 U12281 ( .B1(n10570), .B2(n14893), .A(n10513), .ZN(P1_U3344) );
  INV_X1 U12282 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10542) );
  XNOR2_X1 U12283 ( .A(n10554), .B(n10542), .ZN(n10522) );
  NAND2_X1 U12284 ( .A1(n10515), .A2(n10514), .ZN(n10516) );
  NAND2_X1 U12285 ( .A1(n10517), .A2(n10516), .ZN(n14425) );
  INV_X1 U12286 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10518) );
  MUX2_X1 U12287 ( .A(n10518), .B(P1_REG1_REG_6__SCAN_IN), .S(n14430), .Z(
        n14424) );
  OR2_X1 U12288 ( .A1(n14425), .A2(n14424), .ZN(n14427) );
  NAND2_X1 U12289 ( .A1(n14430), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10519) );
  NAND2_X1 U12290 ( .A1(n14427), .A2(n10519), .ZN(n14440) );
  INV_X1 U12291 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15716) );
  MUX2_X1 U12292 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15716), .S(n14449), .Z(
        n14441) );
  NAND2_X1 U12293 ( .A1(n14440), .A2(n14441), .ZN(n14439) );
  NAND2_X1 U12294 ( .A1(n14449), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10520) );
  AND2_X1 U12295 ( .A1(n14439), .A2(n10520), .ZN(n10521) );
  NAND2_X1 U12296 ( .A1(n10521), .A2(n10522), .ZN(n10545) );
  OAI21_X1 U12297 ( .B1(n10522), .B2(n10521), .A(n10545), .ZN(n10539) );
  NAND2_X1 U12298 ( .A1(n10523), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U12299 ( .A1(n14433), .A2(n14432), .ZN(n10526) );
  MUX2_X1 U12300 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10524), .S(n14430), .Z(
        n10525) );
  NAND2_X1 U12301 ( .A1(n10526), .A2(n10525), .ZN(n14446) );
  NAND2_X1 U12302 ( .A1(n14430), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14445) );
  NAND2_X1 U12303 ( .A1(n14446), .A2(n14445), .ZN(n10529) );
  MUX2_X1 U12304 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10527), .S(n14449), .Z(
        n10528) );
  NAND2_X1 U12305 ( .A1(n10529), .A2(n10528), .ZN(n14448) );
  NAND2_X1 U12306 ( .A1(n14449), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U12307 ( .A1(n14448), .A2(n10534), .ZN(n10532) );
  MUX2_X1 U12308 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10530), .S(n10554), .Z(
        n10531) );
  NAND2_X1 U12309 ( .A1(n10532), .A2(n10531), .ZN(n14462) );
  MUX2_X1 U12310 ( .A(n10530), .B(P1_REG2_REG_8__SCAN_IN), .S(n10554), .Z(
        n10533) );
  NAND3_X1 U12311 ( .A1(n14448), .A2(n10534), .A3(n10533), .ZN(n10535) );
  AND3_X1 U12312 ( .A1(n14553), .A2(n14462), .A3(n10535), .ZN(n10538) );
  NAND2_X1 U12313 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U12314 ( .A1(n14521), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10536) );
  OAI211_X1 U12315 ( .C1(n14518), .C2(n10543), .A(n11870), .B(n10536), .ZN(
        n10537) );
  AOI211_X1 U12316 ( .C1(n14546), .C2(n10539), .A(n10538), .B(n10537), .ZN(
        n10540) );
  INV_X1 U12317 ( .A(n10540), .ZN(P1_U3251) );
  INV_X1 U12318 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10541) );
  MUX2_X1 U12319 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10541), .S(n10734), .Z(
        n10552) );
  NAND2_X1 U12320 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  NAND2_X1 U12321 ( .A1(n10545), .A2(n10544), .ZN(n14455) );
  INV_X1 U12322 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10546) );
  MUX2_X1 U12323 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10546), .S(n14464), .Z(
        n14456) );
  NAND2_X1 U12324 ( .A1(n14455), .A2(n14456), .ZN(n14454) );
  OR2_X1 U12325 ( .A1(n14464), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U12326 ( .A1(n14454), .A2(n10547), .ZN(n14470) );
  MUX2_X1 U12327 ( .A(n12110), .B(P1_REG1_REG_10__SCAN_IN), .S(n14479), .Z(
        n14469) );
  OR2_X1 U12328 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  NAND2_X1 U12329 ( .A1(n14479), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10548) );
  AND2_X1 U12330 ( .A1(n14471), .A2(n10548), .ZN(n14486) );
  INV_X1 U12331 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10549) );
  MUX2_X1 U12332 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10549), .S(n14496), .Z(
        n14485) );
  NAND2_X1 U12333 ( .A1(n14486), .A2(n14485), .ZN(n14484) );
  OR2_X1 U12334 ( .A1(n14496), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U12335 ( .A1(n14484), .A2(n10550), .ZN(n10551) );
  NAND2_X1 U12336 ( .A1(n10551), .A2(n10552), .ZN(n10729) );
  OAI21_X1 U12337 ( .B1(n10552), .B2(n10551), .A(n10729), .ZN(n10553) );
  NAND2_X1 U12338 ( .A1(n10553), .A2(n14546), .ZN(n10569) );
  MUX2_X1 U12339 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9121), .S(n10734), .Z(
        n10563) );
  NAND2_X1 U12340 ( .A1(n10554), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U12341 ( .A1(n14462), .A2(n14461), .ZN(n10557) );
  INV_X1 U12342 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10555) );
  MUX2_X1 U12343 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10555), .S(n14464), .Z(
        n10556) );
  NAND2_X1 U12344 ( .A1(n10557), .A2(n10556), .ZN(n14477) );
  NAND2_X1 U12345 ( .A1(n14464), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U12346 ( .A1(n14477), .A2(n14476), .ZN(n10560) );
  INV_X1 U12347 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U12348 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10558), .S(n14479), .Z(
        n10559) );
  NAND2_X1 U12349 ( .A1(n10560), .A2(n10559), .ZN(n14493) );
  NAND2_X1 U12350 ( .A1(n14479), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n14492) );
  INV_X1 U12351 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10561) );
  MUX2_X1 U12352 ( .A(n10561), .B(P1_REG2_REG_11__SCAN_IN), .S(n14496), .Z(
        n14491) );
  AOI21_X1 U12353 ( .B1(n14493), .B2(n14492), .A(n14491), .ZN(n14490) );
  AOI21_X1 U12354 ( .B1(n14496), .B2(P1_REG2_REG_11__SCAN_IN), .A(n14490), 
        .ZN(n10562) );
  NAND2_X1 U12355 ( .A1(n10562), .A2(n10563), .ZN(n10733) );
  OAI21_X1 U12356 ( .B1(n10563), .B2(n10562), .A(n10733), .ZN(n10567) );
  INV_X1 U12357 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U12358 ( .A1(n14551), .A2(n10734), .ZN(n10564) );
  NAND2_X1 U12359 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12287)
         );
  OAI211_X1 U12360 ( .C1(n10565), .C2(n14557), .A(n10564), .B(n12287), .ZN(
        n10566) );
  AOI21_X1 U12361 ( .B1(n10567), .B2(n14553), .A(n10566), .ZN(n10568) );
  NAND2_X1 U12362 ( .A1(n10569), .A2(n10568), .ZN(P1_U3255) );
  INV_X1 U12363 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10571) );
  INV_X1 U12364 ( .A(n13873), .ZN(n11080) );
  OAI222_X1 U12365 ( .A1(n14244), .A2(n10571), .B1(n14239), .B2(n10570), .C1(
        P2_U3088), .C2(n11080), .ZN(P2_U3316) );
  INV_X1 U12366 ( .A(n15510), .ZN(n12988) );
  INV_X1 U12367 ( .A(n10572), .ZN(n10573) );
  OAI222_X1 U12368 ( .A1(P3_U3151), .A2(n12988), .B1(n13403), .B2(n15047), 
        .C1(n13402), .C2(n10573), .ZN(P3_U3279) );
  OAI222_X1 U12369 ( .A1(P3_U3151), .A2(n12993), .B1(n13402), .B2(n10574), 
        .C1(n13403), .C2(n15044), .ZN(P3_U3278) );
  AOI22_X1 U12370 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15201), .B1(n15205), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10579) );
  INV_X1 U12371 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U12372 ( .A1(n15205), .A2(n10575), .ZN(n10577) );
  NAND2_X1 U12373 ( .A1(n15201), .A2(n10988), .ZN(n10576) );
  AND3_X1 U12374 ( .A1(n15158), .A2(n10577), .A3(n10576), .ZN(n10578) );
  MUX2_X1 U12375 ( .A(n10579), .B(n10578), .S(P2_IR_REG_0__SCAN_IN), .Z(n10581) );
  AOI22_X1 U12376 ( .A1(n15200), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10580) );
  NAND2_X1 U12377 ( .A1(n10581), .A2(n10580), .ZN(P2_U3214) );
  NOR2_X1 U12378 ( .A1(n14521), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12379 ( .A(n10582), .ZN(n10586) );
  AOI22_X1 U12380 ( .A1(n10734), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14880), .ZN(n10583) );
  OAI21_X1 U12381 ( .B1(n10586), .B2(n14893), .A(n10583), .ZN(P1_U3343) );
  AOI22_X1 U12382 ( .A1(n11021), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n14880), .ZN(n10584) );
  OAI21_X1 U12383 ( .B1(n10692), .B2(n14893), .A(n10584), .ZN(P1_U3342) );
  INV_X1 U12384 ( .A(n11086), .ZN(n11380) );
  INV_X1 U12385 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10585) );
  OAI222_X1 U12386 ( .A1(P2_U3088), .A2(n11380), .B1(n14239), .B2(n10586), 
        .C1(n10585), .C2(n14244), .ZN(P2_U3315) );
  NAND2_X1 U12387 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n12505) );
  NOR2_X1 U12388 ( .A1(n10587), .A2(n10977), .ZN(n13825) );
  INV_X1 U12389 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10588) );
  MUX2_X1 U12390 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10588), .S(n13824), .Z(
        n10589) );
  OAI21_X1 U12391 ( .B1(n13829), .B2(n13825), .A(n10589), .ZN(n13845) );
  NAND2_X1 U12392 ( .A1(n13824), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13844) );
  INV_X1 U12393 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11014) );
  MUX2_X1 U12394 ( .A(n11014), .B(P2_REG1_REG_3__SCAN_IN), .S(n13836), .Z(
        n13843) );
  AOI21_X1 U12395 ( .B1(n13845), .B2(n13844), .A(n13843), .ZN(n13842) );
  AOI21_X1 U12396 ( .B1(n13836), .B2(P2_REG1_REG_3__SCAN_IN), .A(n13842), .ZN(
        n10591) );
  INV_X1 U12397 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15642) );
  MUX2_X1 U12398 ( .A(n15642), .B(P2_REG1_REG_4__SCAN_IN), .S(n10646), .Z(
        n10590) );
  NOR2_X1 U12399 ( .A1(n10591), .A2(n10590), .ZN(n10673) );
  AOI211_X1 U12400 ( .C1(n10591), .C2(n10590), .A(n10673), .B(n11089), .ZN(
        n10592) );
  INV_X1 U12401 ( .A(n10592), .ZN(n10593) );
  NAND2_X1 U12402 ( .A1(n12505), .A2(n10593), .ZN(n10603) );
  NAND2_X1 U12403 ( .A1(n10594), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n13820) );
  INV_X1 U12404 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10595) );
  MUX2_X1 U12405 ( .A(n10595), .B(P2_REG2_REG_2__SCAN_IN), .S(n13824), .Z(
        n13821) );
  NOR2_X1 U12406 ( .A1(n10596), .A2(n10595), .ZN(n13835) );
  INV_X1 U12407 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U12408 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11349), .S(n13836), .Z(
        n10597) );
  OAI21_X1 U12409 ( .B1(n13819), .B2(n13835), .A(n10597), .ZN(n13841) );
  NAND2_X1 U12410 ( .A1(n13836), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10600) );
  INV_X1 U12411 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10598) );
  MUX2_X1 U12412 ( .A(n10598), .B(P2_REG2_REG_4__SCAN_IN), .S(n10646), .Z(
        n10599) );
  AOI21_X1 U12413 ( .B1(n13841), .B2(n10600), .A(n10599), .ZN(n10638) );
  AND3_X1 U12414 ( .A1(n13841), .A2(n10600), .A3(n10599), .ZN(n10601) );
  NOR3_X1 U12415 ( .A1(n15180), .A2(n10638), .A3(n10601), .ZN(n10602) );
  AOI211_X1 U12416 ( .C1(n15200), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10603), .B(
        n10602), .ZN(n10604) );
  OAI21_X1 U12417 ( .B1(n10605), .B2(n15158), .A(n10604), .ZN(P2_U3218) );
  NOR2_X1 U12418 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10609) );
  NOR4_X1 U12419 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10608) );
  NOR4_X1 U12420 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10607) );
  NOR4_X1 U12421 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U12422 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10615) );
  NOR4_X1 U12423 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10613) );
  NOR4_X1 U12424 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10612) );
  NOR4_X1 U12425 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10611) );
  NOR4_X1 U12426 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U12427 ( .A1(n10613), .A2(n10612), .A3(n10611), .A4(n10610), .ZN(
        n10614) );
  OAI21_X1 U12428 ( .B1(n10615), .B2(n10614), .A(n10618), .ZN(n11215) );
  NAND2_X1 U12429 ( .A1(n10618), .A2(n10616), .ZN(n11213) );
  AND3_X1 U12430 ( .A1(n11215), .A2(n11213), .A3(n11212), .ZN(n11262) );
  INV_X1 U12431 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U12432 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  NAND2_X1 U12433 ( .A1(n10440), .A2(n14889), .ZN(n14874) );
  NAND2_X1 U12434 ( .A1(n11262), .A2(n11218), .ZN(n10632) );
  INV_X1 U12435 ( .A(n15526), .ZN(n10620) );
  OR2_X1 U12436 ( .A1(n10620), .A2(n15536), .ZN(n11264) );
  OR2_X1 U12437 ( .A1(n10620), .A2(n12019), .ZN(n10621) );
  NAND3_X1 U12438 ( .A1(n10634), .A2(n15919), .A3(n10628), .ZN(n10622) );
  NAND2_X1 U12439 ( .A1(n10632), .A2(n11214), .ZN(n10626) );
  AND3_X1 U12440 ( .A1(n10624), .A2(n10347), .A3(n10623), .ZN(n10625) );
  NAND2_X1 U12441 ( .A1(n10626), .A2(n10625), .ZN(n11207) );
  OR2_X1 U12442 ( .A1(n11207), .A2(P1_U3086), .ZN(n10999) );
  AOI22_X1 U12443 ( .A1(n10627), .A2(n15963), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10999), .ZN(n10637) );
  NAND2_X1 U12444 ( .A1(n15960), .A2(n14765), .ZN(n15942) );
  INV_X1 U12445 ( .A(n15942), .ZN(n14316) );
  INV_X1 U12446 ( .A(n11264), .ZN(n10630) );
  NAND2_X1 U12447 ( .A1(n10634), .A2(n10630), .ZN(n10631) );
  OR2_X1 U12448 ( .A1(n10632), .A2(n10631), .ZN(n10635) );
  AOI22_X1 U12449 ( .A1(n14316), .A2(n8961), .B1(n15527), .B2(n15965), .ZN(
        n10636) );
  NAND2_X1 U12450 ( .A1(n10637), .A2(n10636), .ZN(P1_U3232) );
  INV_X1 U12451 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10639) );
  MUX2_X1 U12452 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10639), .S(n10676), .Z(
        n10662) );
  NOR2_X1 U12453 ( .A1(n10663), .A2(n10662), .ZN(n10661) );
  AOI21_X1 U12454 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10640), .A(n10661), .ZN(
        n15150) );
  INV_X1 U12455 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10641) );
  MUX2_X1 U12456 ( .A(n10641), .B(P2_REG2_REG_6__SCAN_IN), .S(n10648), .Z(
        n15149) );
  NOR2_X1 U12457 ( .A1(n15150), .A2(n15149), .ZN(n15148) );
  INV_X1 U12458 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10642) );
  MUX2_X1 U12459 ( .A(n10642), .B(P2_REG2_REG_7__SCAN_IN), .S(n10683), .Z(
        n10643) );
  NOR2_X1 U12460 ( .A1(n10644), .A2(n10643), .ZN(n10677) );
  AOI211_X1 U12461 ( .C1(n10644), .C2(n10643), .A(n10677), .B(n15180), .ZN(
        n10645) );
  INV_X1 U12462 ( .A(n10645), .ZN(n10654) );
  INV_X1 U12463 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10649) );
  INV_X1 U12464 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10667) );
  AND2_X1 U12465 ( .A1(n10646), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10668) );
  MUX2_X1 U12466 ( .A(n10667), .B(P2_REG1_REG_5__SCAN_IN), .S(n10676), .Z(
        n10647) );
  OAI21_X1 U12467 ( .B1(n10673), .B2(n10668), .A(n10647), .ZN(n10671) );
  OAI21_X1 U12468 ( .B1(n10667), .B2(n10676), .A(n10671), .ZN(n15147) );
  MUX2_X1 U12469 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10649), .S(n10648), .Z(
        n15146) );
  NAND2_X1 U12470 ( .A1(n15147), .A2(n15146), .ZN(n15145) );
  OAI21_X1 U12471 ( .B1(n10649), .B2(n15142), .A(n15145), .ZN(n10652) );
  INV_X1 U12472 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10650) );
  MUX2_X1 U12473 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10650), .S(n10683), .Z(
        n10651) );
  NAND2_X1 U12474 ( .A1(n10652), .A2(n10651), .ZN(n10686) );
  OAI211_X1 U12475 ( .C1(n10652), .C2(n10651), .A(n15201), .B(n10686), .ZN(
        n10653) );
  NAND2_X1 U12476 ( .A1(n10654), .A2(n10653), .ZN(n10656) );
  NAND2_X1 U12477 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n12485) );
  INV_X1 U12478 ( .A(n12485), .ZN(n10655) );
  AOI211_X1 U12479 ( .C1(n15200), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10656), .B(
        n10655), .ZN(n10657) );
  OAI21_X1 U12480 ( .B1(n15158), .B2(n10658), .A(n10657), .ZN(P2_U3221) );
  INV_X1 U12481 ( .A(n10659), .ZN(n10660) );
  OAI222_X1 U12482 ( .A1(P3_U3151), .A2(n13029), .B1(n13403), .B2(n15041), 
        .C1(n13402), .C2(n10660), .ZN(P3_U3277) );
  NAND2_X1 U12483 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11112) );
  AOI211_X1 U12484 ( .C1(n10663), .C2(n10662), .A(n10661), .B(n15180), .ZN(
        n10664) );
  INV_X1 U12485 ( .A(n10664), .ZN(n10665) );
  NAND2_X1 U12486 ( .A1(n11112), .A2(n10665), .ZN(n10666) );
  AOI21_X1 U12487 ( .B1(n15200), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10666), .ZN(
        n10675) );
  MUX2_X1 U12488 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10667), .S(n10676), .Z(
        n10670) );
  INV_X1 U12489 ( .A(n10668), .ZN(n10669) );
  NAND2_X1 U12490 ( .A1(n10670), .A2(n10669), .ZN(n10672) );
  OAI211_X1 U12491 ( .C1(n10673), .C2(n10672), .A(n15201), .B(n10671), .ZN(
        n10674) );
  OAI211_X1 U12492 ( .C1(n15158), .C2(n10676), .A(n10675), .B(n10674), .ZN(
        P2_U3219) );
  NAND2_X1 U12493 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11284) );
  INV_X1 U12494 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10678) );
  MUX2_X1 U12495 ( .A(n10678), .B(P2_REG2_REG_8__SCAN_IN), .S(n10752), .Z(
        n10679) );
  NOR2_X1 U12496 ( .A1(n10680), .A2(n10679), .ZN(n10746) );
  AOI211_X1 U12497 ( .C1(n10680), .C2(n10679), .A(n10746), .B(n15180), .ZN(
        n10681) );
  INV_X1 U12498 ( .A(n10681), .ZN(n10682) );
  NAND2_X1 U12499 ( .A1(n11284), .A2(n10682), .ZN(n10689) );
  NAND2_X1 U12500 ( .A1(n10683), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10685) );
  INV_X1 U12501 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15759) );
  MUX2_X1 U12502 ( .A(n15759), .B(P2_REG1_REG_8__SCAN_IN), .S(n10752), .Z(
        n10684) );
  AOI21_X1 U12503 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(n10751) );
  AND3_X1 U12504 ( .A1(n10686), .A2(n10685), .A3(n10684), .ZN(n10687) );
  NOR3_X1 U12505 ( .A1(n11089), .A2(n10751), .A3(n10687), .ZN(n10688) );
  AOI211_X1 U12506 ( .C1(n15200), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10689), .B(
        n10688), .ZN(n10690) );
  OAI21_X1 U12507 ( .B1(n10691), .B2(n15158), .A(n10690), .ZN(P2_U3222) );
  INV_X1 U12508 ( .A(n15209), .ZN(n11382) );
  OAI222_X1 U12509 ( .A1(n14244), .A2(n7707), .B1(n14239), .B2(n10692), .C1(
        n11382), .C2(P2_U3088), .ZN(P2_U3314) );
  NOR2_X1 U12510 ( .A1(n10965), .A2(n10693), .ZN(n10694) );
  INV_X1 U12511 ( .A(n15139), .ZN(n10967) );
  INV_X1 U12512 ( .A(n10722), .ZN(n10695) );
  NAND2_X1 U12513 ( .A1(n13513), .A2(n14071), .ZN(n13499) );
  INV_X1 U12514 ( .A(n10696), .ZN(n10697) );
  NAND2_X1 U12515 ( .A1(n10697), .A2(n10963), .ZN(n10702) );
  INV_X1 U12516 ( .A(n10698), .ZN(n10699) );
  AND2_X1 U12517 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U12518 ( .A1(n10702), .A2(n10701), .ZN(n11124) );
  OAI22_X1 U12519 ( .A1(n13479), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n13833), .ZN(n10706) );
  NAND2_X1 U12520 ( .A1(n13513), .A2(n14069), .ZN(n13500) );
  NAND2_X1 U12521 ( .A1(n10722), .A2(n10703), .ZN(n10704) );
  OAI22_X1 U12522 ( .A1(n11004), .A2(n13500), .B1(n13506), .B2(n11576), .ZN(
        n10705) );
  AOI211_X1 U12523 ( .C1(n13438), .C2(n13813), .A(n10706), .B(n10705), .ZN(
        n10726) );
  XNOR2_X1 U12524 ( .A(n11104), .B(n13540), .ZN(n10714) );
  INV_X1 U12525 ( .A(n10714), .ZN(n10717) );
  AND2_X1 U12526 ( .A1(n14076), .A2(n13815), .ZN(n10713) );
  INV_X1 U12527 ( .A(n10713), .ZN(n10716) );
  AOI21_X1 U12528 ( .B1(n11109), .B2(n13529), .A(n11174), .ZN(n13442) );
  NOR2_X1 U12529 ( .A1(n10709), .A2(n10708), .ZN(n10711) );
  INV_X1 U12530 ( .A(n10711), .ZN(n10712) );
  NAND2_X1 U12531 ( .A1(n10710), .A2(n10712), .ZN(n10715) );
  NAND2_X1 U12532 ( .A1(n14076), .A2(n13814), .ZN(n10718) );
  NOR2_X1 U12533 ( .A1(n12512), .A2(n10718), .ZN(n11105) );
  NOR2_X1 U12534 ( .A1(n15861), .A2(n10720), .ZN(n10721) );
  OAI211_X1 U12535 ( .C1(n10724), .C2(n10723), .A(n12510), .B(n13507), .ZN(
        n10725) );
  NAND2_X1 U12536 ( .A1(n10726), .A2(n10725), .ZN(P2_U3190) );
  INV_X1 U12537 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U12538 ( .A(n10727), .B(P1_REG1_REG_13__SCAN_IN), .S(n11021), .Z(
        n10732) );
  OR2_X1 U12539 ( .A1(n10734), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U12540 ( .A1(n10729), .A2(n10728), .ZN(n10731) );
  INV_X1 U12541 ( .A(n11023), .ZN(n10730) );
  AOI211_X1 U12542 ( .C1(n10732), .C2(n10731), .A(n14548), .B(n10730), .ZN(
        n10743) );
  OAI21_X1 U12543 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10734), .A(n10733), 
        .ZN(n10737) );
  MUX2_X1 U12544 ( .A(n12210), .B(P1_REG2_REG_13__SCAN_IN), .S(n11021), .Z(
        n10736) );
  INV_X1 U12545 ( .A(n14553), .ZN(n11308) );
  INV_X1 U12546 ( .A(n11019), .ZN(n10735) );
  AOI211_X1 U12547 ( .C1(n10737), .C2(n10736), .A(n11308), .B(n10735), .ZN(
        n10742) );
  INV_X1 U12548 ( .A(n11021), .ZN(n10740) );
  INV_X1 U12549 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12250) );
  NOR2_X1 U12550 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12250), .ZN(n10738) );
  AOI21_X1 U12551 ( .B1(n14521), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10738), 
        .ZN(n10739) );
  OAI21_X1 U12552 ( .B1(n14518), .B2(n10740), .A(n10739), .ZN(n10741) );
  OR3_X1 U12553 ( .A1(n10743), .A2(n10742), .A3(n10741), .ZN(P1_U3256) );
  INV_X1 U12554 ( .A(SI_19_), .ZN(n15020) );
  INV_X1 U12555 ( .A(n10744), .ZN(n10745) );
  OAI222_X1 U12556 ( .A1(n13403), .A2(n15020), .B1(n13402), .B2(n10745), .C1(
        n13042), .C2(P3_U3151), .ZN(P3_U3276) );
  INV_X1 U12557 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10747) );
  MUX2_X1 U12558 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10747), .S(n13860), .Z(
        n13852) );
  NAND2_X1 U12559 ( .A1(n13853), .A2(n13852), .ZN(n13851) );
  OAI21_X1 U12560 ( .B1(n13860), .B2(P2_REG2_REG_9__SCAN_IN), .A(n13851), .ZN(
        n10750) );
  INV_X1 U12561 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10748) );
  MUX2_X1 U12562 ( .A(n10748), .B(P2_REG2_REG_10__SCAN_IN), .S(n11078), .Z(
        n10749) );
  NOR2_X1 U12563 ( .A1(n10750), .A2(n10749), .ZN(n11077) );
  AOI211_X1 U12564 ( .C1(n10750), .C2(n10749), .A(n15180), .B(n11077), .ZN(
        n10759) );
  AOI21_X1 U12565 ( .B1(n10752), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10751), .ZN(
        n13858) );
  INV_X1 U12566 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10753) );
  MUX2_X1 U12567 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10753), .S(n13860), .Z(
        n13857) );
  NAND2_X1 U12568 ( .A1(n13858), .A2(n13857), .ZN(n13856) );
  OAI21_X1 U12569 ( .B1(n13860), .B2(P2_REG1_REG_9__SCAN_IN), .A(n13856), .ZN(
        n10755) );
  INV_X1 U12570 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11071) );
  MUX2_X1 U12571 ( .A(n11071), .B(P2_REG1_REG_10__SCAN_IN), .S(n11078), .Z(
        n10754) );
  NOR2_X1 U12572 ( .A1(n10755), .A2(n10754), .ZN(n13879) );
  AOI211_X1 U12573 ( .C1(n10755), .C2(n10754), .A(n11089), .B(n13879), .ZN(
        n10758) );
  NAND2_X1 U12574 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12572)
         );
  NAND2_X1 U12575 ( .A1(n15200), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10756) );
  OAI211_X1 U12576 ( .C1(n15158), .C2(n11072), .A(n12572), .B(n10756), .ZN(
        n10757) );
  OR3_X1 U12577 ( .A1(n10759), .A2(n10758), .A3(n10757), .ZN(P2_U3224) );
  NAND2_X1 U12578 ( .A1(n13025), .A2(n11525), .ZN(n10760) );
  NAND2_X1 U12579 ( .A1(n10760), .A2(n11070), .ZN(n10764) );
  INV_X1 U12580 ( .A(n10761), .ZN(n10762) );
  XNOR2_X1 U12581 ( .A(n15557), .B(n7191), .ZN(n10917) );
  XNOR2_X1 U12582 ( .A(n9652), .B(n10917), .ZN(n10768) );
  NAND2_X1 U12583 ( .A1(n15127), .A2(n11039), .ZN(n10765) );
  NAND2_X1 U12584 ( .A1(n15548), .A2(n10765), .ZN(n10767) );
  INV_X1 U12585 ( .A(n10919), .ZN(n10766) );
  AOI21_X1 U12586 ( .B1(n10768), .B2(n10767), .A(n10766), .ZN(n10796) );
  INV_X1 U12587 ( .A(n10778), .ZN(n10769) );
  NAND3_X1 U12588 ( .A1(n10769), .A2(n10781), .A3(n15797), .ZN(n10772) );
  INV_X1 U12589 ( .A(n10774), .ZN(n10770) );
  NAND3_X1 U12590 ( .A1(n10770), .A2(n10803), .A3(n10789), .ZN(n10771) );
  INV_X1 U12591 ( .A(n15131), .ZN(n12890) );
  OAI211_X1 U12592 ( .C1(n10774), .C2(n10789), .A(n10896), .B(n10773), .ZN(
        n10775) );
  INV_X1 U12593 ( .A(n10775), .ZN(n10776) );
  OAI21_X1 U12594 ( .B1(n10778), .B2(n10777), .A(n10776), .ZN(n10780) );
  NOR2_X1 U12595 ( .A1(n10785), .A2(n10789), .ZN(n10779) );
  AOI21_X1 U12596 ( .B1(n10780), .B2(P3_STATE_REG_SCAN_IN), .A(n10779), .ZN(
        n11034) );
  AND2_X1 U12597 ( .A1(n11034), .A2(n13393), .ZN(n15132) );
  INV_X1 U12598 ( .A(n15132), .ZN(n10794) );
  NAND2_X1 U12599 ( .A1(n10781), .A2(n15737), .ZN(n10784) );
  INV_X1 U12600 ( .A(n10788), .ZN(n10786) );
  AND2_X1 U12601 ( .A1(n10786), .A2(n10789), .ZN(n10787) );
  AND2_X1 U12602 ( .A1(n10789), .A2(n10788), .ZN(n10790) );
  INV_X1 U12603 ( .A(n15126), .ZN(n12895) );
  AOI22_X1 U12604 ( .A1(n12876), .A2(n10042), .B1(n12895), .B2(n15546), .ZN(
        n10792) );
  OAI21_X1 U12605 ( .B1(n15553), .B2(n15128), .A(n10792), .ZN(n10793) );
  AOI21_X1 U12606 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10794), .A(n10793), .ZN(
        n10795) );
  OAI21_X1 U12607 ( .B1(n10796), .B2(n12890), .A(n10795), .ZN(P3_U3162) );
  INV_X2 U12608 ( .A(n7384), .ZN(n12955) );
  MUX2_X1 U12609 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12955), .Z(n10928) );
  XNOR2_X1 U12610 ( .A(n10928), .B(n10927), .ZN(n10929) );
  MUX2_X1 U12611 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12955), .Z(n10797) );
  XNOR2_X1 U12612 ( .A(n10797), .B(n10954), .ZN(n10949) );
  INV_X1 U12613 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10905) );
  INV_X1 U12614 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10826) );
  MUX2_X1 U12615 ( .A(n10905), .B(n10826), .S(n12955), .Z(n15375) );
  NAND2_X1 U12616 ( .A1(n15375), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15374) );
  OAI22_X1 U12617 ( .A1(n10949), .A2(n15374), .B1(n10797), .B2(n10954), .ZN(
        n10878) );
  MUX2_X1 U12618 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12955), .Z(n10798) );
  XNOR2_X1 U12619 ( .A(n10798), .B(n10892), .ZN(n10879) );
  INV_X1 U12620 ( .A(n10798), .ZN(n10799) );
  AOI22_X1 U12621 ( .A1(n10878), .A2(n10879), .B1(n10892), .B2(n10799), .ZN(
        n10848) );
  MUX2_X1 U12622 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12955), .Z(n10800) );
  XNOR2_X1 U12623 ( .A(n10800), .B(n10835), .ZN(n10849) );
  OAI22_X1 U12624 ( .A1(n10848), .A2(n10849), .B1(n10800), .B2(n10835), .ZN(
        n10861) );
  MUX2_X1 U12625 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12955), .Z(n10801) );
  XNOR2_X1 U12626 ( .A(n10801), .B(n10875), .ZN(n10862) );
  INV_X1 U12627 ( .A(n10801), .ZN(n10802) );
  AOI22_X1 U12628 ( .A1(n10861), .A2(n10862), .B1(n10875), .B2(n10802), .ZN(
        n10930) );
  XOR2_X1 U12629 ( .A(n10929), .B(n10930), .Z(n10847) );
  NAND2_X1 U12630 ( .A1(P3_U3897), .A2(n12134), .ZN(n15460) );
  NAND2_X1 U12631 ( .A1(n10286), .A2(n10804), .ZN(n10806) );
  AND2_X1 U12632 ( .A1(n10806), .A2(n10805), .ZN(n10822) );
  INV_X1 U12633 ( .A(n10807), .ZN(n10808) );
  INV_X1 U12634 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10809) );
  NAND2_X1 U12635 ( .A1(n9660), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U12636 ( .A1(n10954), .A2(n10813), .ZN(n10812) );
  INV_X1 U12637 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U12638 ( .A1(n10827), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10810) );
  OR2_X1 U12639 ( .A1(n10810), .A2(n9660), .ZN(n10811) );
  NAND2_X1 U12640 ( .A1(n10812), .A2(n10811), .ZN(n10950) );
  NAND2_X1 U12641 ( .A1(n10950), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U12642 ( .A1(n10814), .A2(n10813), .ZN(n10881) );
  NAND2_X1 U12643 ( .A1(n10833), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U12644 ( .A1(n10880), .A2(n10815), .ZN(n10816) );
  INV_X1 U12645 ( .A(n10835), .ZN(n10858) );
  NAND2_X1 U12646 ( .A1(n10816), .A2(n10835), .ZN(n10817) );
  INV_X1 U12647 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10818) );
  MUX2_X1 U12648 ( .A(n10818), .B(P3_REG2_REG_4__SCAN_IN), .S(n10875), .Z(
        n10863) );
  AOI21_X1 U12649 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10819), .A(n10866), .ZN(
        n10937) );
  INV_X1 U12650 ( .A(n10927), .ZN(n10938) );
  XNOR2_X1 U12651 ( .A(n10937), .B(n10938), .ZN(n10939) );
  INV_X1 U12652 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11684) );
  XNOR2_X1 U12653 ( .A(n10939), .B(n11684), .ZN(n10845) );
  INV_X1 U12654 ( .A(n10825), .ZN(n10821) );
  MUX2_X1 U12655 ( .A(n10821), .B(n12925), .S(n10820), .Z(n15491) );
  INV_X1 U12656 ( .A(n10822), .ZN(n10823) );
  NOR2_X1 U12657 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9696), .ZN(n11394) );
  AOI21_X1 U12658 ( .B1(n15502), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11394), .ZN(
        n10843) );
  MUX2_X1 U12659 ( .A(n15582), .B(P3_REG1_REG_2__SCAN_IN), .S(n10892), .Z(
        n10886) );
  NAND2_X1 U12660 ( .A1(n9660), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U12661 ( .A1(n10954), .A2(n10831), .ZN(n10830) );
  NAND2_X1 U12662 ( .A1(n10827), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10828) );
  OR2_X1 U12663 ( .A1(n10828), .A2(n9660), .ZN(n10829) );
  NAND2_X1 U12664 ( .A1(n10830), .A2(n10829), .ZN(n10951) );
  NAND2_X1 U12665 ( .A1(n10951), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U12666 ( .A1(n10832), .A2(n10831), .ZN(n10885) );
  NAND2_X1 U12667 ( .A1(n10886), .A2(n10885), .ZN(n10884) );
  NAND2_X1 U12668 ( .A1(n10833), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U12669 ( .A1(n10884), .A2(n10834), .ZN(n10836) );
  XNOR2_X1 U12670 ( .A(n10836), .B(n10858), .ZN(n10852) );
  NAND2_X1 U12671 ( .A1(n10852), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U12672 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  NAND2_X1 U12673 ( .A1(n10838), .A2(n10837), .ZN(n10868) );
  INV_X1 U12674 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10839) );
  MUX2_X1 U12675 ( .A(n10839), .B(P3_REG1_REG_4__SCAN_IN), .S(n10875), .Z(
        n10869) );
  NAND2_X1 U12676 ( .A1(n10868), .A2(n10869), .ZN(n10867) );
  OR2_X1 U12677 ( .A1(n10875), .A2(n10839), .ZN(n10840) );
  NAND2_X1 U12678 ( .A1(n10867), .A2(n10840), .ZN(n10931) );
  XNOR2_X1 U12679 ( .A(n10931), .B(n10927), .ZN(n10934) );
  INV_X1 U12680 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10933) );
  XNOR2_X1 U12681 ( .A(n10934), .B(n10933), .ZN(n10841) );
  NAND2_X1 U12682 ( .A1(n15514), .A2(n10841), .ZN(n10842) );
  OAI211_X1 U12683 ( .C1(n15491), .C2(n10927), .A(n10843), .B(n10842), .ZN(
        n10844) );
  AOI21_X1 U12684 ( .B1(n15517), .B2(n10845), .A(n10844), .ZN(n10846) );
  OAI21_X1 U12685 ( .B1(n10847), .B2(n15460), .A(n10846), .ZN(P3_U3187) );
  XOR2_X1 U12686 ( .A(n10849), .B(n10848), .Z(n10860) );
  XNOR2_X1 U12687 ( .A(n10850), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U12688 ( .A1(n15517), .A2(n10851), .ZN(n10856) );
  XNOR2_X1 U12689 ( .A(n10852), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U12690 ( .A1(n15514), .A2(n10853), .ZN(n10855) );
  NOR2_X1 U12691 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15013), .ZN(n11042) );
  AOI21_X1 U12692 ( .B1(n15502), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11042), .ZN(
        n10854) );
  NAND3_X1 U12693 ( .A1(n10856), .A2(n10855), .A3(n10854), .ZN(n10857) );
  AOI21_X1 U12694 ( .B1(n15503), .B2(n10858), .A(n10857), .ZN(n10859) );
  OAI21_X1 U12695 ( .B1(n10860), .B2(n15460), .A(n10859), .ZN(P3_U3185) );
  XOR2_X1 U12696 ( .A(n10862), .B(n10861), .Z(n10877) );
  NOR2_X1 U12697 ( .A1(n10864), .A2(n10863), .ZN(n10865) );
  OAI21_X1 U12698 ( .B1(n10866), .B2(n10865), .A(n15517), .ZN(n10873) );
  INV_X1 U12699 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15098) );
  NOR2_X1 U12700 ( .A1(n15098), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11185) );
  AOI21_X1 U12701 ( .B1(n15502), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11185), .ZN(
        n10872) );
  OAI21_X1 U12702 ( .B1(n10869), .B2(n10868), .A(n10867), .ZN(n10870) );
  NAND2_X1 U12703 ( .A1(n15514), .A2(n10870), .ZN(n10871) );
  NAND3_X1 U12704 ( .A1(n10873), .A2(n10872), .A3(n10871), .ZN(n10874) );
  AOI21_X1 U12705 ( .B1(n15503), .B2(n10875), .A(n10874), .ZN(n10876) );
  OAI21_X1 U12706 ( .B1(n10877), .B2(n15460), .A(n10876), .ZN(P3_U3186) );
  XOR2_X1 U12707 ( .A(n10879), .B(n10878), .Z(n10894) );
  OAI21_X1 U12708 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(n10883) );
  NAND2_X1 U12709 ( .A1(n15517), .A2(n10883), .ZN(n10890) );
  OAI21_X1 U12710 ( .B1(n10886), .B2(n10885), .A(n10884), .ZN(n10887) );
  NAND2_X1 U12711 ( .A1(n15514), .A2(n10887), .ZN(n10889) );
  AOI22_X1 U12712 ( .A1(n15502), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10888) );
  NAND3_X1 U12713 ( .A1(n10890), .A2(n10889), .A3(n10888), .ZN(n10891) );
  AOI21_X1 U12714 ( .B1(n15503), .B2(n10892), .A(n10891), .ZN(n10893) );
  OAI21_X1 U12715 ( .B1(n10894), .B2(n15460), .A(n10893), .ZN(P3_U3184) );
  XNOR2_X1 U12716 ( .A(n10895), .B(n13392), .ZN(n10898) );
  NAND3_X1 U12717 ( .A1(n10898), .A2(n10897), .A3(n10896), .ZN(n10901) );
  NAND3_X1 U12718 ( .A1(n15130), .A2(n15797), .A3(n10899), .ZN(n10900) );
  OAI21_X1 U12719 ( .B1(n9652), .B2(n13243), .A(n10900), .ZN(n10961) );
  NAND2_X1 U12720 ( .A1(n10961), .A2(n15688), .ZN(n10904) );
  INV_X1 U12721 ( .A(n10901), .ZN(n10902) );
  AND2_X1 U12722 ( .A1(n11526), .A2(n15737), .ZN(n15585) );
  INV_X2 U12723 ( .A(n13143), .ZN(n15680) );
  AOI22_X1 U12724 ( .A1(n15684), .A2(n10906), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15680), .ZN(n10903) );
  OAI211_X1 U12725 ( .C1(n10905), .C2(n15688), .A(n10904), .B(n10903), .ZN(
        P3_U3233) );
  INV_X1 U12726 ( .A(n10961), .ZN(n10908) );
  AOI22_X1 U12727 ( .A1(n15971), .A2(n10906), .B1(n15970), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10907) );
  OAI21_X1 U12728 ( .B1(n10908), .B2(n15970), .A(n10907), .ZN(P3_U3459) );
  NAND2_X2 U12729 ( .A1(n10910), .A2(n10909), .ZN(n11634) );
  INV_X1 U12730 ( .A(n10989), .ZN(n10912) );
  XOR2_X1 U12731 ( .A(n10992), .B(n10993), .Z(n10916) );
  NOR2_X1 U12732 ( .A1(n14326), .A2(n15903), .ZN(n14345) );
  AOI22_X1 U12733 ( .A1(n14345), .A2(n14375), .B1(n11503), .B2(n15965), .ZN(
        n10915) );
  AOI22_X1 U12734 ( .A1(n14316), .A2(n14374), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10999), .ZN(n10914) );
  OAI211_X1 U12735 ( .C1(n10916), .C2(n15949), .A(n10915), .B(n10914), .ZN(
        P1_U3222) );
  INV_X1 U12736 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10926) );
  XNOR2_X1 U12737 ( .A(n15580), .B(n11039), .ZN(n11035) );
  XNOR2_X1 U12738 ( .A(n11035), .B(n11531), .ZN(n10921) );
  NAND2_X1 U12739 ( .A1(n9652), .A2(n10917), .ZN(n10918) );
  NAND2_X1 U12740 ( .A1(n10920), .A2(n10921), .ZN(n11038) );
  OAI21_X1 U12741 ( .B1(n10921), .B2(n10920), .A(n11038), .ZN(n10922) );
  NAND2_X1 U12742 ( .A1(n10922), .A2(n15131), .ZN(n10925) );
  OAI22_X1 U12743 ( .A1(n9652), .A2(n12897), .B1(n15574), .B2(n15126), .ZN(
        n10923) );
  AOI21_X1 U12744 ( .B1(n15586), .B2(n12887), .A(n10923), .ZN(n10924) );
  OAI211_X1 U12745 ( .C1(n15132), .C2(n10926), .A(n10925), .B(n10924), .ZN(
        P3_U3177) );
  MUX2_X1 U12746 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12955), .Z(n11048) );
  XNOR2_X1 U12747 ( .A(n11048), .B(n11050), .ZN(n11051) );
  OAI22_X1 U12748 ( .A1(n10930), .A2(n10929), .B1(n10928), .B2(n10927), .ZN(
        n11052) );
  XOR2_X1 U12749 ( .A(n11051), .B(n11052), .Z(n10948) );
  INV_X1 U12750 ( .A(n10931), .ZN(n10932) );
  INV_X1 U12751 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U12752 ( .A1(n11050), .A2(n15679), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n11056), .ZN(n10935) );
  NAND2_X1 U12753 ( .A1(n10935), .A2(n10936), .ZN(n11053) );
  OAI21_X1 U12754 ( .B1(n10936), .B2(n10935), .A(n11053), .ZN(n10946) );
  INV_X1 U12755 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U12756 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15120), .ZN(n11481) );
  AOI21_X1 U12757 ( .B1(n15502), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11481), .ZN(
        n10944) );
  OAI22_X1 U12758 ( .A1(n10939), .A2(n11684), .B1(n10938), .B2(n10937), .ZN(
        n10941) );
  INV_X1 U12759 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15687) );
  AOI22_X1 U12760 ( .A1(n11050), .A2(n15687), .B1(P3_REG2_REG_6__SCAN_IN), 
        .B2(n11056), .ZN(n10940) );
  NAND2_X1 U12761 ( .A1(n10940), .A2(n10941), .ZN(n11057) );
  OAI21_X1 U12762 ( .B1(n10941), .B2(n10940), .A(n11057), .ZN(n10942) );
  NAND2_X1 U12763 ( .A1(n15517), .A2(n10942), .ZN(n10943) );
  OAI211_X1 U12764 ( .C1(n15491), .C2(n11056), .A(n10944), .B(n10943), .ZN(
        n10945) );
  AOI21_X1 U12765 ( .B1(n15514), .B2(n10946), .A(n10945), .ZN(n10947) );
  OAI21_X1 U12766 ( .B1(n10948), .B2(n15460), .A(n10947), .ZN(P3_U3188) );
  XOR2_X1 U12767 ( .A(n15374), .B(n10949), .Z(n10959) );
  XNOR2_X1 U12768 ( .A(n10950), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n10957) );
  INV_X1 U12769 ( .A(n15514), .ZN(n15373) );
  XOR2_X1 U12770 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n10951), .Z(n10953) );
  AOI22_X1 U12771 ( .A1(n15502), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10952) );
  OAI21_X1 U12772 ( .B1(n15373), .B2(n10953), .A(n10952), .ZN(n10956) );
  NOR2_X1 U12773 ( .A1(n15491), .A2(n10954), .ZN(n10955) );
  AOI211_X1 U12774 ( .C1(n15517), .C2(n10957), .A(n10956), .B(n10955), .ZN(
        n10958) );
  OAI21_X1 U12775 ( .B1(n15460), .B2(n10959), .A(n10958), .ZN(P3_U3183) );
  OAI22_X1 U12776 ( .A1(n15127), .A2(n13391), .B1(n15978), .B2(n9631), .ZN(
        n10960) );
  AOI21_X1 U12777 ( .B1(n15978), .B2(n10961), .A(n10960), .ZN(n10962) );
  INV_X1 U12778 ( .A(n10962), .ZN(P3_U3390) );
  AND2_X1 U12779 ( .A1(n10964), .A2(n10963), .ZN(n10966) );
  AND2_X1 U12780 ( .A1(n15140), .A2(n10965), .ZN(n14902) );
  INV_X1 U12781 ( .A(n14127), .ZN(n14165) );
  INV_X1 U12782 ( .A(n10968), .ZN(n10971) );
  INV_X1 U12783 ( .A(n10969), .ZN(n10970) );
  AOI21_X1 U12784 ( .B1(n10971), .B2(n13745), .A(n10970), .ZN(n11316) );
  OAI21_X1 U12785 ( .B1(n10984), .B2(n13745), .A(n11320), .ZN(n10976) );
  OAI22_X1 U12786 ( .A1(n11004), .A2(n14057), .B1(n10973), .B2(n14055), .ZN(
        n10975) );
  NOR2_X1 U12787 ( .A1(n11316), .A2(n10707), .ZN(n10974) );
  AOI211_X1 U12788 ( .C1(n14074), .C2(n10976), .A(n10975), .B(n10974), .ZN(
        n11310) );
  OAI211_X1 U12789 ( .C1(n13522), .C2(n13529), .A(n13976), .B(n11325), .ZN(
        n11312) );
  OAI211_X1 U12790 ( .C1(n11316), .C2(n11095), .A(n11310), .B(n11312), .ZN(
        n11413) );
  NOR2_X1 U12791 ( .A1(n15869), .A2(n10977), .ZN(n10978) );
  AOI21_X1 U12792 ( .B1(n11413), .B2(n15869), .A(n10978), .ZN(n10979) );
  OAI21_X1 U12793 ( .B1(n13522), .B2(n14165), .A(n10979), .ZN(P2_U3500) );
  INV_X1 U12794 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10981) );
  INV_X1 U12795 ( .A(n10980), .ZN(n10982) );
  INV_X1 U12796 ( .A(n11388), .ZN(n11969) );
  OAI222_X1 U12797 ( .A1(n14244), .A2(n10981), .B1(n14239), .B2(n10982), .C1(
        P2_U3088), .C2(n11969), .ZN(P2_U3313) );
  INV_X1 U12798 ( .A(n11300), .ZN(n11025) );
  OAI222_X1 U12799 ( .A1(n14897), .A2(n10983), .B1(n14893), .B2(n10982), .C1(
        P1_U3086), .C2(n11025), .ZN(P1_U3341) );
  AOI21_X1 U12800 ( .B1(n13529), .B2(n13528), .A(n10984), .ZN(n13748) );
  AOI21_X1 U12801 ( .B1(n14063), .B2(n10707), .A(n13748), .ZN(n10985) );
  NOR2_X1 U12802 ( .A1(n13521), .A2(n14057), .ZN(n11171) );
  NOR2_X1 U12803 ( .A1(n10985), .A2(n11171), .ZN(n11254) );
  NAND2_X1 U12804 ( .A1(n10986), .A2(n13523), .ZN(n11255) );
  OAI211_X1 U12805 ( .C1(n13748), .C2(n11095), .A(n11254), .B(n11255), .ZN(
        n11194) );
  NAND2_X1 U12806 ( .A1(n15869), .A2(n11194), .ZN(n10987) );
  OAI21_X1 U12807 ( .B1(n15869), .B2(n10988), .A(n10987), .ZN(P2_U3499) );
  NAND2_X1 U12808 ( .A1(n14374), .A2(n7192), .ZN(n10996) );
  NAND2_X1 U12809 ( .A1(n11516), .A2(n10994), .ZN(n10995) );
  NAND2_X1 U12810 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  XNOR2_X1 U12811 ( .A(n10997), .B(n11634), .ZN(n11201) );
  INV_X1 U12812 ( .A(n14374), .ZN(n11236) );
  OAI22_X1 U12813 ( .A1(n11236), .A2(n12706), .B1(n15596), .B2(n12640), .ZN(
        n11200) );
  XNOR2_X1 U12814 ( .A(n11201), .B(n11200), .ZN(n11203) );
  XOR2_X1 U12815 ( .A(n11204), .B(n11203), .Z(n11001) );
  AOI22_X1 U12816 ( .A1(n8961), .A2(n14767), .B1(n14765), .B2(n14373), .ZN(
        n11509) );
  OAI22_X1 U12817 ( .A1(n11509), .A2(n14326), .B1(n14348), .B2(n15596), .ZN(
        n10998) );
  AOI21_X1 U12818 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10999), .A(n10998), .ZN(
        n11000) );
  OAI21_X1 U12819 ( .B1(n11001), .B2(n15949), .A(n11000), .ZN(P1_U3237) );
  OAI21_X1 U12820 ( .B1(n11003), .B2(n13749), .A(n11002), .ZN(n11011) );
  INV_X1 U12821 ( .A(n11011), .ZN(n11354) );
  INV_X1 U12822 ( .A(n10707), .ZN(n14060) );
  OAI22_X1 U12823 ( .A1(n11118), .A2(n14057), .B1(n11004), .B2(n14055), .ZN(
        n11010) );
  NAND3_X1 U12824 ( .A1(n11006), .A2(n13749), .A3(n11007), .ZN(n11008) );
  AOI21_X1 U12825 ( .B1(n11005), .B2(n11008), .A(n14063), .ZN(n11009) );
  AOI211_X1 U12826 ( .C1(n14060), .C2(n11011), .A(n11010), .B(n11009), .ZN(
        n11348) );
  NAND2_X1 U12827 ( .A1(n11327), .A2(n13544), .ZN(n11012) );
  NAND2_X1 U12828 ( .A1(n11012), .A2(n13976), .ZN(n11013) );
  OR2_X1 U12829 ( .A1(n11013), .A2(n11343), .ZN(n11350) );
  OAI211_X1 U12830 ( .C1(n11354), .C2(n11095), .A(n11348), .B(n11350), .ZN(
        n11578) );
  OAI22_X1 U12831 ( .A1(n14165), .A2(n11576), .B1(n15869), .B2(n11014), .ZN(
        n11015) );
  AOI21_X1 U12832 ( .B1(n15869), .B2(n11578), .A(n11015), .ZN(n11016) );
  INV_X1 U12833 ( .A(n11016), .ZN(P2_U3502) );
  NAND2_X1 U12834 ( .A1(n11021), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11018) );
  MUX2_X1 U12835 ( .A(n9162), .B(P1_REG2_REG_14__SCAN_IN), .S(n11300), .Z(
        n11017) );
  AOI21_X1 U12836 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11295) );
  NAND3_X1 U12837 ( .A1(n11019), .A2(n11018), .A3(n11017), .ZN(n11020) );
  NAND2_X1 U12838 ( .A1(n11020), .A2(n14553), .ZN(n11030) );
  NAND2_X1 U12839 ( .A1(n11021), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11022) );
  NAND2_X1 U12840 ( .A1(n11023), .A2(n11022), .ZN(n11299) );
  XNOR2_X1 U12841 ( .A(n11299), .B(n11025), .ZN(n11024) );
  NAND2_X1 U12842 ( .A1(n11024), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11297) );
  OAI211_X1 U12843 ( .C1(n11024), .C2(P1_REG1_REG_14__SCAN_IN), .A(n11297), 
        .B(n14546), .ZN(n11029) );
  NAND2_X1 U12844 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14256)
         );
  INV_X1 U12845 ( .A(n14256), .ZN(n11027) );
  NOR2_X1 U12846 ( .A1(n14518), .A2(n11025), .ZN(n11026) );
  AOI211_X1 U12847 ( .C1(n14521), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11027), 
        .B(n11026), .ZN(n11028) );
  OAI211_X1 U12848 ( .C1(n11295), .C2(n11030), .A(n11029), .B(n11028), .ZN(
        P1_U3257) );
  NAND2_X1 U12849 ( .A1(n12925), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11031) );
  OAI21_X1 U12850 ( .B1(n11032), .B2(n12925), .A(n11031), .ZN(P3_U3521) );
  NAND2_X1 U12851 ( .A1(n12925), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11033) );
  OAI21_X1 U12852 ( .B1(n13064), .B2(n12925), .A(n11033), .ZN(P3_U3520) );
  INV_X1 U12853 ( .A(n11035), .ZN(n11036) );
  NAND2_X1 U12854 ( .A1(n11036), .A2(n11531), .ZN(n11037) );
  XNOR2_X1 U12855 ( .A(n11045), .B(n11478), .ZN(n11179) );
  XNOR2_X1 U12856 ( .A(n11179), .B(n15574), .ZN(n11040) );
  OAI211_X1 U12857 ( .C1(n11041), .C2(n11040), .A(n11182), .B(n15131), .ZN(
        n11047) );
  AOI21_X1 U12858 ( .B1(n12876), .B2(n15546), .A(n11042), .ZN(n11043) );
  OAI21_X1 U12859 ( .B1(n11530), .B2(n15126), .A(n11043), .ZN(n11044) );
  AOI21_X1 U12860 ( .B1(n11045), .B2(n12887), .A(n11044), .ZN(n11046) );
  OAI211_X1 U12861 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11990), .A(n11047), .B(
        n11046), .ZN(P3_U3158) );
  MUX2_X1 U12862 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12955), .Z(n11142) );
  XNOR2_X1 U12863 ( .A(n11142), .B(n11155), .ZN(n11143) );
  INV_X1 U12864 ( .A(n11048), .ZN(n11049) );
  AOI22_X1 U12865 ( .A1(n11052), .A2(n11051), .B1(n11050), .B2(n11049), .ZN(
        n11144) );
  XOR2_X1 U12866 ( .A(n11143), .B(n11144), .Z(n11066) );
  NAND2_X1 U12867 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n11056), .ZN(n11054) );
  NAND2_X1 U12868 ( .A1(n11054), .A2(n11053), .ZN(n11148) );
  XOR2_X1 U12869 ( .A(n11148), .B(n11155), .Z(n11055) );
  NAND2_X1 U12870 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n11055), .ZN(n11149) );
  OAI21_X1 U12871 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11055), .A(n11149), .ZN(
        n11064) );
  NAND2_X1 U12872 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n11056), .ZN(n11058) );
  OAI21_X1 U12873 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11059), .A(n11156), .ZN(
        n11060) );
  NAND2_X1 U12874 ( .A1(n11060), .A2(n15517), .ZN(n11062) );
  INV_X1 U12875 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15080) );
  NOR2_X1 U12876 ( .A1(n15080), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11652) );
  AOI21_X1 U12877 ( .B1(n15502), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11652), .ZN(
        n11061) );
  OAI211_X1 U12878 ( .C1(n15491), .C2(n11155), .A(n11062), .B(n11061), .ZN(
        n11063) );
  AOI21_X1 U12879 ( .B1(n15514), .B2(n11064), .A(n11063), .ZN(n11065) );
  OAI21_X1 U12880 ( .B1(n11066), .B2(n15460), .A(n11065), .ZN(P3_U3189) );
  INV_X1 U12881 ( .A(n11067), .ZN(n11069) );
  INV_X1 U12882 ( .A(SI_20_), .ZN(n11068) );
  OAI222_X1 U12883 ( .A1(P3_U3151), .A2(n11070), .B1(n13402), .B2(n11069), 
        .C1(n11068), .C2(n13403), .ZN(P3_U3275) );
  INV_X1 U12884 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n13874) );
  NOR2_X1 U12885 ( .A1(n11072), .A2(n11071), .ZN(n13872) );
  MUX2_X1 U12886 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13874), .S(n13873), .Z(
        n11073) );
  OAI21_X1 U12887 ( .B1(n13879), .B2(n13872), .A(n11073), .ZN(n13877) );
  OAI21_X1 U12888 ( .B1(n13874), .B2(n11080), .A(n13877), .ZN(n11076) );
  INV_X1 U12889 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11074) );
  MUX2_X1 U12890 ( .A(n11074), .B(P2_REG1_REG_12__SCAN_IN), .S(n11086), .Z(
        n11075) );
  NOR2_X1 U12891 ( .A1(n11076), .A2(n11075), .ZN(n11379) );
  AOI21_X1 U12892 ( .B1(n11076), .B2(n11075), .A(n11379), .ZN(n11090) );
  INV_X1 U12893 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11079) );
  MUX2_X1 U12894 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11079), .S(n13873), .Z(
        n13866) );
  NAND2_X1 U12895 ( .A1(n13867), .A2(n13866), .ZN(n13865) );
  NAND2_X1 U12896 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  MUX2_X1 U12897 ( .A(n11375), .B(P2_REG2_REG_12__SCAN_IN), .S(n11086), .Z(
        n11082) );
  AND3_X1 U12898 ( .A1(n13865), .A2(n11082), .A3(n11081), .ZN(n11083) );
  OAI21_X1 U12899 ( .B1(n11374), .B2(n11083), .A(n15205), .ZN(n11088) );
  NAND2_X1 U12900 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11084)
         );
  OAI21_X1 U12901 ( .B1(n15198), .B2(n7398), .A(n11084), .ZN(n11085) );
  AOI21_X1 U12902 ( .B1(n11086), .B2(n15210), .A(n11085), .ZN(n11087) );
  OAI211_X1 U12903 ( .C1(n11090), .C2(n11089), .A(n11088), .B(n11087), .ZN(
        P2_U3226) );
  NAND2_X1 U12904 ( .A1(n12925), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11091) );
  OAI21_X1 U12905 ( .B1(n13077), .B2(n12925), .A(n11091), .ZN(P3_U3519) );
  INV_X1 U12906 ( .A(n11092), .ZN(n11094) );
  INV_X1 U12907 ( .A(SI_21_), .ZN(n11093) );
  OAI222_X1 U12908 ( .A1(n13402), .A2(n11094), .B1(n13403), .B2(n11093), .C1(
        P3_U3151), .C2(n11525), .ZN(P3_U3274) );
  OAI21_X1 U12909 ( .B1(n11097), .B2(n11101), .A(n11096), .ZN(n11555) );
  NAND2_X1 U12910 ( .A1(n7234), .A2(n13567), .ZN(n11098) );
  NAND2_X1 U12911 ( .A1(n11098), .A2(n13976), .ZN(n11099) );
  NOR2_X1 U12912 ( .A1(n11453), .A2(n11099), .ZN(n11550) );
  XNOR2_X1 U12913 ( .A(n11100), .B(n11101), .ZN(n11102) );
  AOI22_X1 U12914 ( .A1(n14071), .A2(n13809), .B1(n13811), .B2(n14069), .ZN(
        n13511) );
  OAI21_X1 U12915 ( .B1(n11102), .B2(n14063), .A(n13511), .ZN(n11552) );
  AOI211_X1 U12916 ( .C1(n15859), .C2(n11555), .A(n11550), .B(n11552), .ZN(
        n11561) );
  AOI22_X1 U12917 ( .A1(n14127), .A2(n13567), .B1(n15868), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11103) );
  OAI21_X1 U12918 ( .B1(n11561), .B2(n15868), .A(n11103), .ZN(P2_U3505) );
  XNOR2_X1 U12919 ( .A(n13554), .B(n11104), .ZN(n11107) );
  NAND2_X1 U12920 ( .A1(n14076), .A2(n13813), .ZN(n11108) );
  XNOR2_X1 U12921 ( .A(n11107), .B(n11108), .ZN(n12513) );
  INV_X1 U12922 ( .A(n11105), .ZN(n11106) );
  INV_X1 U12923 ( .A(n11107), .ZN(n11117) );
  NAND2_X1 U12924 ( .A1(n11117), .A2(n11108), .ZN(n11110) );
  XNOR2_X1 U12925 ( .A(n13559), .B(n11109), .ZN(n11274) );
  NAND2_X1 U12926 ( .A1(n14076), .A2(n13811), .ZN(n11273) );
  XNOR2_X1 U12927 ( .A(n11274), .B(n11273), .ZN(n11120) );
  AOI21_X1 U12928 ( .B1(n12519), .B2(n11110), .A(n11120), .ZN(n11111) );
  INV_X1 U12929 ( .A(n11403), .ZN(n11113) );
  OAI21_X1 U12930 ( .B1(n13479), .B2(n11113), .A(n11112), .ZN(n11116) );
  INV_X1 U12931 ( .A(n13559), .ZN(n11567) );
  OAI22_X1 U12932 ( .A1(n11114), .A2(n13499), .B1(n13506), .B2(n11567), .ZN(
        n11115) );
  AOI211_X1 U12933 ( .C1(n13439), .C2(n13813), .A(n11116), .B(n11115), .ZN(
        n11122) );
  INV_X2 U12934 ( .A(n13507), .ZN(n13486) );
  OAI22_X1 U12935 ( .A1(n13484), .A2(n11118), .B1(n11117), .B2(n13486), .ZN(
        n11119) );
  NAND3_X1 U12936 ( .A1(n12519), .A2(n11120), .A3(n11119), .ZN(n11121) );
  OAI211_X1 U12937 ( .C1(n11276), .C2(n13486), .A(n11122), .B(n11121), .ZN(
        P2_U3199) );
  INV_X1 U12938 ( .A(n11123), .ZN(n11132) );
  OR2_X1 U12939 ( .A1(n11124), .A2(P2_U3088), .ZN(n13440) );
  NOR2_X1 U12940 ( .A1(n13506), .A2(n15604), .ZN(n11126) );
  OAI22_X1 U12941 ( .A1(n13521), .A2(n13500), .B1(n13499), .B2(n12511), .ZN(
        n11125) );
  AOI211_X1 U12942 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n13440), .A(n11126), .B(
        n11125), .ZN(n11131) );
  OAI22_X1 U12943 ( .A1(n13484), .A2(n13521), .B1(n10710), .B2(n13486), .ZN(
        n11129) );
  NAND3_X1 U12944 ( .A1(n11129), .A2(n11128), .A3(n11127), .ZN(n11130) );
  OAI211_X1 U12945 ( .C1(n13486), .C2(n11132), .A(n11131), .B(n11130), .ZN(
        P2_U3209) );
  OR2_X1 U12946 ( .A1(n11133), .A2(n13751), .ZN(n11134) );
  NAND2_X1 U12947 ( .A1(n11135), .A2(n11134), .ZN(n11409) );
  AOI21_X1 U12948 ( .B1(n11342), .B2(n13559), .A(n14076), .ZN(n11136) );
  AND2_X1 U12949 ( .A1(n11136), .A2(n7234), .ZN(n11404) );
  XNOR2_X1 U12950 ( .A(n11137), .B(n13751), .ZN(n11140) );
  NAND2_X1 U12951 ( .A1(n11409), .A2(n14060), .ZN(n11139) );
  AOI22_X1 U12952 ( .A1(n14071), .A2(n13810), .B1(n13813), .B2(n14069), .ZN(
        n11138) );
  OAI211_X1 U12953 ( .C1(n14063), .C2(n11140), .A(n11139), .B(n11138), .ZN(
        n11406) );
  AOI211_X1 U12954 ( .C1(n15758), .C2(n11409), .A(n11404), .B(n11406), .ZN(
        n11570) );
  AOI22_X1 U12955 ( .A1(n14127), .A2(n13559), .B1(n15868), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n11141) );
  OAI21_X1 U12956 ( .B1(n11570), .B2(n15868), .A(n11141), .ZN(P2_U3504) );
  OAI22_X1 U12957 ( .A1(n11144), .A2(n11143), .B1(n11142), .B2(n11155), .ZN(
        n11146) );
  MUX2_X1 U12958 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12955), .Z(n12946) );
  XNOR2_X1 U12959 ( .A(n12946), .B(n11153), .ZN(n11145) );
  NAND2_X1 U12960 ( .A1(n11146), .A2(n11145), .ZN(n12947) );
  OAI21_X1 U12961 ( .B1(n11146), .B2(n11145), .A(n12947), .ZN(n11147) );
  INV_X1 U12962 ( .A(n15460), .ZN(n15515) );
  NAND2_X1 U12963 ( .A1(n11147), .A2(n15515), .ZN(n11166) );
  INV_X1 U12964 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15738) );
  AOI22_X1 U12965 ( .A1(n11153), .A2(n15738), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n12972), .ZN(n11152) );
  NAND2_X1 U12966 ( .A1(n11155), .A2(n11148), .ZN(n11150) );
  NAND2_X1 U12967 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  NAND2_X1 U12968 ( .A1(n11152), .A2(n11151), .ZN(n12973) );
  OAI21_X1 U12969 ( .B1(n11152), .B2(n11151), .A(n12973), .ZN(n11164) );
  INV_X1 U12970 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U12971 ( .A1(n11153), .A2(n11799), .B1(P3_REG2_REG_8__SCAN_IN), 
        .B2(n12972), .ZN(n11159) );
  NAND2_X1 U12972 ( .A1(n11155), .A2(n11154), .ZN(n11157) );
  NAND2_X1 U12973 ( .A1(n11159), .A2(n11158), .ZN(n12927) );
  OAI21_X1 U12974 ( .B1(n11159), .B2(n11158), .A(n12927), .ZN(n11160) );
  NAND2_X1 U12975 ( .A1(n11160), .A2(n15517), .ZN(n11162) );
  NOR2_X1 U12976 ( .A1(n15090), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11746) );
  AOI21_X1 U12977 ( .B1(n15502), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11746), .ZN(
        n11161) );
  OAI211_X1 U12978 ( .C1(n15491), .C2(n12972), .A(n11162), .B(n11161), .ZN(
        n11163) );
  AOI21_X1 U12979 ( .B1(n15514), .B2(n11164), .A(n11163), .ZN(n11165) );
  NAND2_X1 U12980 ( .A1(n11166), .A2(n11165), .ZN(P3_U3190) );
  INV_X1 U12981 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11168) );
  INV_X1 U12982 ( .A(n11167), .ZN(n11169) );
  INV_X1 U12983 ( .A(n11971), .ZN(n15157) );
  OAI222_X1 U12984 ( .A1(n14244), .A2(n11168), .B1(n14239), .B2(n11169), .C1(
        n15157), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U12985 ( .A(n11305), .ZN(n11587) );
  OAI222_X1 U12986 ( .A1(n14897), .A2(n11170), .B1(n14893), .B2(n11169), .C1(
        n11587), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI22_X1 U12987 ( .A1(n13428), .A2(n13528), .B1(n13523), .B2(n13507), .ZN(
        n11175) );
  AOI22_X1 U12988 ( .A1(n13513), .A2(n11171), .B1(n13440), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n11173) );
  INV_X1 U12989 ( .A(n13506), .ZN(n13516) );
  NAND2_X1 U12990 ( .A1(n13516), .A2(n13523), .ZN(n11172) );
  OAI211_X1 U12991 ( .C1(n11175), .C2(n11174), .A(n11173), .B(n11172), .ZN(
        P2_U3204) );
  OAI22_X1 U12992 ( .A1(n11176), .A2(P3_U3151), .B1(SI_22_), .B2(n13403), .ZN(
        n11177) );
  AOI21_X1 U12993 ( .B1(n11178), .B2(n11355), .A(n11177), .ZN(P3_U3273) );
  XNOR2_X1 U12994 ( .A(n11189), .B(n11039), .ZN(n11391) );
  XNOR2_X1 U12995 ( .A(n11391), .B(n12922), .ZN(n11184) );
  INV_X1 U12996 ( .A(n11179), .ZN(n11180) );
  OR2_X1 U12997 ( .A1(n15574), .A2(n11180), .ZN(n11181) );
  AOI21_X1 U12998 ( .B1(n11184), .B2(n11183), .A(n7345), .ZN(n11192) );
  INV_X1 U12999 ( .A(n11185), .ZN(n11186) );
  OAI21_X1 U13000 ( .B1(n15574), .B2(n12897), .A(n11186), .ZN(n11187) );
  AOI21_X1 U13001 ( .B1(n12895), .B2(n12921), .A(n11187), .ZN(n11188) );
  OAI21_X1 U13002 ( .B1(n15128), .B2(n11189), .A(n11188), .ZN(n11190) );
  AOI21_X1 U13003 ( .B1(n11546), .B2(n12900), .A(n11190), .ZN(n11191) );
  OAI21_X1 U13004 ( .B1(n11192), .B2(n12890), .A(n11191), .ZN(P3_U3170) );
  NAND2_X1 U13005 ( .A1(n14215), .A2(n11194), .ZN(n11195) );
  OAI21_X1 U13006 ( .B1(n14215), .B2(n8276), .A(n11195), .ZN(P2_U3430) );
  NAND2_X1 U13007 ( .A1(n14373), .A2(n7192), .ZN(n11197) );
  NAND2_X1 U13008 ( .A1(n11364), .A2(n10994), .ZN(n11196) );
  NAND2_X1 U13009 ( .A1(n11197), .A2(n11196), .ZN(n11199) );
  XNOR2_X1 U13010 ( .A(n11199), .B(n11634), .ZN(n11432) );
  OAI22_X1 U13011 ( .A1(n11239), .A2(n12706), .B1(n15620), .B2(n12640), .ZN(
        n11431) );
  XNOR2_X1 U13012 ( .A(n11432), .B(n11431), .ZN(n11206) );
  OAI21_X1 U13013 ( .B1(n11204), .B2(n11203), .A(n11202), .ZN(n11205) );
  AOI211_X1 U13014 ( .C1(n11206), .C2(n11205), .A(n15949), .B(n11434), .ZN(
        n11211) );
  AOI22_X1 U13015 ( .A1(n15969), .A2(n11363), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n11210) );
  INV_X1 U13016 ( .A(n14345), .ZN(n15945) );
  AOI22_X1 U13017 ( .A1(n14316), .A2(n14372), .B1(n11364), .B2(n15965), .ZN(
        n11208) );
  OAI21_X1 U13018 ( .B1(n11236), .B2(n15945), .A(n11208), .ZN(n11209) );
  OR3_X1 U13019 ( .A1(n11211), .A2(n11210), .A3(n11209), .ZN(P1_U3218) );
  NAND2_X1 U13020 ( .A1(n11213), .A2(n11212), .ZN(n11216) );
  NAND3_X1 U13021 ( .A1(n11216), .A2(n11215), .A3(n11214), .ZN(n11217) );
  OR2_X1 U13022 ( .A1(n11217), .A2(n11260), .ZN(n11249) );
  INV_X2 U13023 ( .A(n15926), .ZN(n15719) );
  INV_X1 U13024 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U13025 ( .A1(n11220), .A2(n11219), .ZN(n11221) );
  NAND2_X1 U13026 ( .A1(n11266), .A2(n12019), .ZN(n15771) );
  NAND2_X1 U13027 ( .A1(n14375), .A2(n15527), .ZN(n11499) );
  NAND2_X1 U13028 ( .A1(n11224), .A2(n11499), .ZN(n11226) );
  NAND2_X1 U13029 ( .A1(n11226), .A2(n11225), .ZN(n11517) );
  INV_X1 U13030 ( .A(n11517), .ZN(n11227) );
  AOI21_X1 U13031 ( .B1(n11227), .B2(n8140), .A(n8139), .ZN(n11361) );
  NAND2_X1 U13032 ( .A1(n11361), .A2(n11366), .ZN(n11360) );
  NAND2_X1 U13033 ( .A1(n11239), .A2(n15620), .ZN(n11228) );
  NAND2_X1 U13034 ( .A1(n11360), .A2(n11228), .ZN(n11711) );
  XOR2_X1 U13035 ( .A(n11711), .B(n11242), .Z(n11267) );
  OR2_X1 U13036 ( .A1(n11229), .A2(n12019), .ZN(n11231) );
  NAND2_X1 U13037 ( .A1(n11233), .A2(n11232), .ZN(n11235) );
  NAND2_X1 U13038 ( .A1(n11235), .A2(n11234), .ZN(n11508) );
  NAND2_X1 U13039 ( .A1(n11236), .A2(n11516), .ZN(n11237) );
  NAND2_X1 U13040 ( .A1(n11507), .A2(n11237), .ZN(n11367) );
  NAND2_X1 U13041 ( .A1(n14373), .A2(n15620), .ZN(n11238) );
  NAND2_X1 U13042 ( .A1(n11367), .A2(n11238), .ZN(n11241) );
  NAND2_X1 U13043 ( .A1(n11239), .A2(n11364), .ZN(n11240) );
  XOR2_X1 U13044 ( .A(n11700), .B(n11242), .Z(n11243) );
  AOI222_X1 U13045 ( .A1(n15914), .A2(n11243), .B1(n14373), .B2(n14767), .C1(
        n14371), .C2(n14765), .ZN(n11272) );
  NAND2_X1 U13046 ( .A1(n11362), .A2(n11709), .ZN(n11244) );
  NAND2_X1 U13047 ( .A1(n11244), .A2(n15917), .ZN(n11245) );
  NOR2_X1 U13048 ( .A1(n15656), .A2(n11245), .ZN(n11270) );
  AOI21_X1 U13049 ( .B1(n11709), .B2(n15887), .A(n11270), .ZN(n11246) );
  OAI211_X1 U13050 ( .C1(n15851), .C2(n11267), .A(n11272), .B(n11246), .ZN(
        n11250) );
  NAND2_X1 U13051 ( .A1(n11250), .A2(n15719), .ZN(n11247) );
  OAI21_X1 U13052 ( .B1(n15719), .B2(n11248), .A(n11247), .ZN(P1_U3471) );
  INV_X2 U13053 ( .A(n15924), .ZN(n15717) );
  NAND2_X1 U13054 ( .A1(n11250), .A2(n15717), .ZN(n11251) );
  OAI21_X1 U13055 ( .B1(n15717), .B2(n11252), .A(n11251), .ZN(P1_U3532) );
  OAI21_X1 U13056 ( .B1(n13780), .B2(n11255), .A(n11254), .ZN(n11256) );
  AOI21_X1 U13057 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n15816), .A(n11256), .ZN(
        n11257) );
  NOR2_X1 U13058 ( .A1(n11257), .A2(n13980), .ZN(n11258) );
  AOI21_X1 U13059 ( .B1(n15818), .B2(P2_REG2_REG_0__SCAN_IN), .A(n11258), .ZN(
        n11259) );
  OAI21_X1 U13060 ( .B1(n13748), .B2(n14066), .A(n11259), .ZN(P2_U3265) );
  INV_X1 U13061 ( .A(n11260), .ZN(n11263) );
  NAND3_X1 U13062 ( .A1(n11263), .A2(n11262), .A3(n11261), .ZN(n14585) );
  AOI22_X1 U13063 ( .A1(n15941), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n11442), 
        .B2(n15930), .ZN(n11265) );
  OAI21_X1 U13064 ( .B1(n15723), .B2(n11712), .A(n11265), .ZN(n11269) );
  INV_X1 U13065 ( .A(n11266), .ZN(n12115) );
  NOR2_X1 U13066 ( .A1(n11267), .A2(n14740), .ZN(n11268) );
  AOI211_X1 U13067 ( .C1(n11270), .C2(n15935), .A(n11269), .B(n11268), .ZN(
        n11271) );
  OAI21_X1 U13068 ( .B1(n15941), .B2(n11272), .A(n11271), .ZN(P1_U3289) );
  AND2_X2 U13069 ( .A1(n11276), .A2(n11275), .ZN(n13510) );
  XNOR2_X1 U13070 ( .A(n13567), .B(n11109), .ZN(n12481) );
  NAND2_X1 U13071 ( .A1(n14076), .A2(n13810), .ZN(n11277) );
  NOR2_X1 U13072 ( .A1(n12481), .A2(n11277), .ZN(n11278) );
  AOI21_X1 U13073 ( .B1(n12481), .B2(n11277), .A(n11278), .ZN(n13509) );
  XNOR2_X1 U13074 ( .A(n13576), .B(n12728), .ZN(n11281) );
  NAND2_X1 U13075 ( .A1(n14076), .A2(n13809), .ZN(n11282) );
  XNOR2_X1 U13076 ( .A(n11281), .B(n11282), .ZN(n12482) );
  INV_X1 U13077 ( .A(n11278), .ZN(n11279) );
  INV_X1 U13078 ( .A(n11281), .ZN(n11289) );
  NAND2_X1 U13079 ( .A1(n11289), .A2(n11282), .ZN(n11283) );
  XNOR2_X1 U13080 ( .A(n13580), .B(n12728), .ZN(n12589) );
  NOR2_X1 U13081 ( .A1(n12488), .A2(n13976), .ZN(n11832) );
  XNOR2_X1 U13082 ( .A(n12589), .B(n11832), .ZN(n11291) );
  INV_X1 U13083 ( .A(n12592), .ZN(n11294) );
  INV_X1 U13084 ( .A(n11425), .ZN(n11286) );
  AOI22_X1 U13085 ( .A1(n13438), .A2(n13807), .B1(n13439), .B2(n13809), .ZN(
        n11285) );
  OAI211_X1 U13086 ( .C1(n11286), .C2(n13479), .A(n11285), .B(n11284), .ZN(
        n11287) );
  AOI21_X1 U13087 ( .B1(n13580), .B2(n13516), .A(n11287), .ZN(n11293) );
  OAI22_X1 U13088 ( .A1(n13484), .A2(n11420), .B1(n11289), .B2(n13486), .ZN(
        n11290) );
  NAND3_X1 U13089 ( .A1(n11288), .A2(n11291), .A3(n11290), .ZN(n11292) );
  OAI211_X1 U13090 ( .C1(n11294), .C2(n13486), .A(n11293), .B(n11292), .ZN(
        P2_U3193) );
  AOI21_X1 U13091 ( .B1(n11300), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11295), 
        .ZN(n11588) );
  XNOR2_X1 U13092 ( .A(n11588), .B(n11587), .ZN(n11296) );
  NOR2_X1 U13093 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11296), .ZN(n11586) );
  AOI21_X1 U13094 ( .B1(n11296), .B2(P1_REG2_REG_15__SCAN_IN), .A(n11586), 
        .ZN(n11309) );
  INV_X1 U13095 ( .A(n11297), .ZN(n11298) );
  AOI21_X1 U13096 ( .B1(n11300), .B2(n11299), .A(n11298), .ZN(n11580) );
  XNOR2_X1 U13097 ( .A(n11580), .B(n11305), .ZN(n11301) );
  INV_X1 U13098 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15882) );
  NAND2_X1 U13099 ( .A1(n11301), .A2(n15882), .ZN(n11581) );
  OAI21_X1 U13100 ( .B1(n11301), .B2(n15882), .A(n11581), .ZN(n11302) );
  NAND2_X1 U13101 ( .A1(n11302), .A2(n14546), .ZN(n11307) );
  INV_X1 U13102 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U13103 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14346)
         );
  OAI21_X1 U13104 ( .B1(n14557), .B2(n11303), .A(n14346), .ZN(n11304) );
  AOI21_X1 U13105 ( .B1(n14551), .B2(n11305), .A(n11304), .ZN(n11306) );
  OAI211_X1 U13106 ( .C1(n11309), .C2(n11308), .A(n11307), .B(n11306), .ZN(
        P1_U3258) );
  MUX2_X1 U13107 ( .A(n10328), .B(n11310), .S(n7197), .Z(n11315) );
  OAI22_X1 U13108 ( .A1(n13984), .A2(n11312), .B1(n11311), .B2(n13959), .ZN(
        n11313) );
  AOI21_X1 U13109 ( .B1(n14035), .B2(n13534), .A(n11313), .ZN(n11314) );
  OAI211_X1 U13110 ( .C1(n11316), .C2(n14066), .A(n11315), .B(n11314), .ZN(
        P2_U3264) );
  OAI21_X1 U13111 ( .B1(n11318), .B2(n11321), .A(n11317), .ZN(n15608) );
  INV_X1 U13112 ( .A(n15608), .ZN(n11331) );
  OAI22_X1 U13113 ( .A1(n12511), .A2(n14057), .B1(n13521), .B2(n14055), .ZN(
        n11324) );
  NAND3_X1 U13114 ( .A1(n11321), .A2(n11320), .A3(n11319), .ZN(n11322) );
  AOI21_X1 U13115 ( .B1(n11322), .B2(n11006), .A(n14063), .ZN(n11323) );
  AOI211_X1 U13116 ( .C1(n14060), .C2(n15608), .A(n11324), .B(n11323), .ZN(
        n15605) );
  MUX2_X1 U13117 ( .A(n15605), .B(n10595), .S(n15818), .Z(n11330) );
  NAND2_X1 U13118 ( .A1(n13540), .A2(n11325), .ZN(n11326) );
  NAND3_X1 U13119 ( .A1(n11327), .A2(n13976), .A3(n11326), .ZN(n15603) );
  OAI22_X1 U13120 ( .A1(n13984), .A2(n15603), .B1(n8284), .B2(n13959), .ZN(
        n11328) );
  AOI21_X1 U13121 ( .B1(n14035), .B2(n13540), .A(n11328), .ZN(n11329) );
  OAI211_X1 U13122 ( .C1(n11331), .C2(n14066), .A(n11330), .B(n11329), .ZN(
        P2_U3263) );
  OR2_X1 U13123 ( .A1(n11332), .A2(n13750), .ZN(n11333) );
  NAND2_X1 U13124 ( .A1(n11334), .A2(n11333), .ZN(n15639) );
  INV_X1 U13125 ( .A(n15639), .ZN(n11347) );
  NAND3_X1 U13126 ( .A1(n11005), .A2(n13750), .A3(n11335), .ZN(n11336) );
  NAND2_X1 U13127 ( .A1(n11337), .A2(n11336), .ZN(n11338) );
  NAND2_X1 U13128 ( .A1(n11338), .A2(n14074), .ZN(n11340) );
  AOI22_X1 U13129 ( .A1(n14069), .A2(n13814), .B1(n13811), .B2(n14071), .ZN(
        n11339) );
  NAND2_X1 U13130 ( .A1(n11340), .A2(n11339), .ZN(n11341) );
  AOI21_X1 U13131 ( .B1(n15639), .B2(n14060), .A(n11341), .ZN(n15641) );
  MUX2_X1 U13132 ( .A(n10598), .B(n15641), .S(n7197), .Z(n11346) );
  OAI211_X1 U13133 ( .C1(n11343), .C2(n15637), .A(n13976), .B(n11342), .ZN(
        n15636) );
  OAI22_X1 U13134 ( .A1(n13984), .A2(n15636), .B1(n12506), .B2(n13959), .ZN(
        n11344) );
  AOI21_X1 U13135 ( .B1(n14035), .B2(n13554), .A(n11344), .ZN(n11345) );
  OAI211_X1 U13136 ( .C1(n11347), .C2(n14066), .A(n11346), .B(n11345), .ZN(
        P2_U3261) );
  MUX2_X1 U13137 ( .A(n11349), .B(n11348), .S(n7197), .Z(n11353) );
  OAI22_X1 U13138 ( .A1(n13984), .A2(n11350), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13959), .ZN(n11351) );
  AOI21_X1 U13139 ( .B1(n14035), .B2(n13544), .A(n11351), .ZN(n11352) );
  OAI211_X1 U13140 ( .C1(n11354), .C2(n14066), .A(n11353), .B(n11352), .ZN(
        P2_U3262) );
  INV_X1 U13141 ( .A(SI_23_), .ZN(n11359) );
  NAND2_X1 U13142 ( .A1(n11356), .A2(n11355), .ZN(n11358) );
  OAI211_X1 U13143 ( .C1(n11359), .C2(n13403), .A(n11358), .B(n11357), .ZN(
        P3_U3272) );
  OR2_X1 U13144 ( .A1(n15941), .A2(n15534), .ZN(n12122) );
  INV_X1 U13145 ( .A(n12122), .ZN(n15784) );
  OAI21_X1 U13146 ( .B1(n11361), .B2(n11366), .A(n11360), .ZN(n15623) );
  OAI211_X1 U13147 ( .C1(n7556), .C2(n15620), .A(n15917), .B(n11362), .ZN(
        n15619) );
  AOI22_X1 U13148 ( .A1(n15931), .A2(n11364), .B1(n15930), .B2(n11363), .ZN(
        n11365) );
  OAI21_X1 U13149 ( .B1(n14672), .B2(n15619), .A(n11365), .ZN(n11372) );
  XNOR2_X1 U13150 ( .A(n11367), .B(n11366), .ZN(n11370) );
  INV_X1 U13151 ( .A(n15771), .ZN(n15749) );
  NAND2_X1 U13152 ( .A1(n15623), .A2(n15749), .ZN(n11369) );
  AOI22_X1 U13153 ( .A1(n14767), .A2(n14374), .B1(n14372), .B2(n14765), .ZN(
        n11368) );
  OAI211_X1 U13154 ( .C1(n15890), .C2(n11370), .A(n11369), .B(n11368), .ZN(
        n15621) );
  MUX2_X1 U13155 ( .A(n15621), .B(P1_REG2_REG_3__SCAN_IN), .S(n15941), .Z(
        n11371) );
  AOI211_X1 U13156 ( .C1(n15784), .C2(n15623), .A(n11372), .B(n11371), .ZN(
        n11373) );
  INV_X1 U13157 ( .A(n11373), .ZN(P1_U3290) );
  INV_X1 U13158 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13159 ( .A1(n11388), .A2(n11968), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n11969), .ZN(n11378) );
  NAND2_X1 U13160 ( .A1(n15209), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11376) );
  INV_X1 U13161 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11375) );
  AOI21_X1 U13162 ( .B1(n11375), .B2(n11380), .A(n11374), .ZN(n15208) );
  XNOR2_X1 U13163 ( .A(n11382), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n15207) );
  NAND2_X1 U13164 ( .A1(n11376), .A2(n15206), .ZN(n11377) );
  AOI21_X1 U13165 ( .B1(n11378), .B2(n11377), .A(n11967), .ZN(n11390) );
  INV_X1 U13166 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U13167 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12495)
         );
  INV_X1 U13168 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11381) );
  AOI21_X1 U13169 ( .B1(n11074), .B2(n11380), .A(n11379), .ZN(n15204) );
  XNOR2_X1 U13170 ( .A(n11382), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15203) );
  NAND2_X1 U13171 ( .A1(n15204), .A2(n15203), .ZN(n15202) );
  OAI21_X1 U13172 ( .B1(n11382), .B2(n11381), .A(n15202), .ZN(n11385) );
  INV_X1 U13173 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11383) );
  MUX2_X1 U13174 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n11383), .S(n11388), .Z(
        n11384) );
  NAND2_X1 U13175 ( .A1(n11384), .A2(n11385), .ZN(n11957) );
  OAI211_X1 U13176 ( .C1(n11385), .C2(n11384), .A(n15201), .B(n11957), .ZN(
        n11386) );
  OAI211_X1 U13177 ( .C1(n15319), .C2(n15198), .A(n12495), .B(n11386), .ZN(
        n11387) );
  AOI21_X1 U13178 ( .B1(n15210), .B2(n11388), .A(n11387), .ZN(n11389) );
  OAI21_X1 U13179 ( .B1(n11390), .B2(n15180), .A(n11389), .ZN(P2_U3228) );
  XNOR2_X1 U13180 ( .A(n11686), .B(n7205), .ZN(n11473) );
  XNOR2_X1 U13181 ( .A(n11473), .B(n11545), .ZN(n11476) );
  INV_X1 U13182 ( .A(n11391), .ZN(n11392) );
  XOR2_X1 U13183 ( .A(n11476), .B(n11477), .Z(n11398) );
  NOR2_X1 U13184 ( .A1(n11530), .A2(n12897), .ZN(n11393) );
  AOI211_X1 U13185 ( .C1(n12895), .C2(n12920), .A(n11394), .B(n11393), .ZN(
        n11395) );
  OAI21_X1 U13186 ( .B1(n15128), .B2(n15647), .A(n11395), .ZN(n11396) );
  AOI21_X1 U13187 ( .B1(n11685), .B2(n12900), .A(n11396), .ZN(n11397) );
  OAI21_X1 U13188 ( .B1(n11398), .B2(n12890), .A(n11397), .ZN(P3_U3167) );
  INV_X1 U13189 ( .A(n14505), .ZN(n14512) );
  OAI222_X1 U13190 ( .A1(n14897), .A2(n11399), .B1(n14893), .B2(n11401), .C1(
        n14512), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U13191 ( .A1(n14244), .A2(n11402), .B1(n14239), .B2(n11401), .C1(
        n12033), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13192 ( .A(n14066), .ZN(n11410) );
  AOI22_X1 U13193 ( .A1(n15814), .A2(n11404), .B1(n11403), .B2(n15816), .ZN(
        n11405) );
  OAI21_X1 U13194 ( .B1(n11567), .B2(n15821), .A(n11405), .ZN(n11408) );
  MUX2_X1 U13195 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11406), .S(n7197), .Z(
        n11407) );
  AOI211_X1 U13196 ( .C1(n11410), .C2(n11409), .A(n11408), .B(n11407), .ZN(
        n11411) );
  INV_X1 U13197 ( .A(n11411), .ZN(P2_U3260) );
  NOR2_X1 U13198 ( .A1(n14215), .A2(n8260), .ZN(n11412) );
  AOI21_X1 U13199 ( .B1(n11413), .B2(n14215), .A(n11412), .ZN(n11414) );
  OAI21_X1 U13200 ( .B1(n13522), .B2(n14219), .A(n11414), .ZN(P2_U3433) );
  NAND2_X1 U13201 ( .A1(n11415), .A2(n11419), .ZN(n11416) );
  NAND2_X1 U13202 ( .A1(n11417), .A2(n11416), .ZN(n15751) );
  XNOR2_X1 U13203 ( .A(n11418), .B(n11419), .ZN(n11423) );
  OAI22_X1 U13204 ( .A1(n11421), .A2(n14057), .B1(n11420), .B2(n14055), .ZN(
        n11422) );
  AOI21_X1 U13205 ( .B1(n11423), .B2(n14074), .A(n11422), .ZN(n11424) );
  OAI21_X1 U13206 ( .B1(n15751), .B2(n10707), .A(n11424), .ZN(n15755) );
  NAND2_X1 U13207 ( .A1(n15755), .A2(n7197), .ZN(n11430) );
  OAI211_X1 U13208 ( .C1(n15754), .C2(n11454), .A(n13976), .B(n11467), .ZN(
        n15752) );
  INV_X1 U13209 ( .A(n15752), .ZN(n11428) );
  AOI22_X1 U13210 ( .A1(n15818), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11425), 
        .B2(n15816), .ZN(n11426) );
  OAI21_X1 U13211 ( .B1(n15821), .B2(n15754), .A(n11426), .ZN(n11427) );
  AOI21_X1 U13212 ( .B1(n15814), .B2(n11428), .A(n11427), .ZN(n11429) );
  OAI211_X1 U13213 ( .C1(n15751), .C2(n14066), .A(n11430), .B(n11429), .ZN(
        P2_U3257) );
  AOI22_X1 U13214 ( .A1(n14372), .A2(n11435), .B1(n7192), .B2(n11709), .ZN(
        n11436) );
  NOR2_X1 U13215 ( .A1(n11597), .A2(n7346), .ZN(n11438) );
  INV_X1 U13216 ( .A(n14372), .ZN(n11713) );
  OAI22_X1 U13217 ( .A1(n11713), .A2(n12640), .B1(n11712), .B2(n12708), .ZN(
        n11437) );
  XNOR2_X1 U13218 ( .A(n11437), .B(n11634), .ZN(n11598) );
  XNOR2_X1 U13219 ( .A(n11438), .B(n11598), .ZN(n11444) );
  AOI22_X1 U13220 ( .A1(n14316), .A2(n14371), .B1(n14345), .B2(n14373), .ZN(
        n11440) );
  OAI211_X1 U13221 ( .C1(n11712), .C2(n14348), .A(n11440), .B(n11439), .ZN(
        n11441) );
  AOI21_X1 U13222 ( .B1(n11442), .B2(n14352), .A(n11441), .ZN(n11443) );
  OAI21_X1 U13223 ( .B1(n11444), .B2(n15949), .A(n11443), .ZN(P1_U3230) );
  OAI21_X1 U13224 ( .B1(n11446), .B2(n11448), .A(n11445), .ZN(n11489) );
  INV_X1 U13225 ( .A(n11489), .ZN(n11460) );
  XNOR2_X1 U13226 ( .A(n11447), .B(n11448), .ZN(n11451) );
  NAND2_X1 U13227 ( .A1(n11489), .A2(n14060), .ZN(n11450) );
  AOI22_X1 U13228 ( .A1(n14071), .A2(n13808), .B1(n13810), .B2(n14069), .ZN(
        n11449) );
  OAI211_X1 U13229 ( .C1(n14063), .C2(n11451), .A(n11450), .B(n11449), .ZN(
        n11487) );
  INV_X1 U13230 ( .A(n11487), .ZN(n11452) );
  MUX2_X1 U13231 ( .A(n10642), .B(n11452), .S(n7197), .Z(n11459) );
  OAI21_X1 U13232 ( .B1(n11453), .B2(n12487), .A(n13976), .ZN(n11455) );
  NOR2_X1 U13233 ( .A1(n11455), .A2(n11454), .ZN(n11488) );
  INV_X1 U13234 ( .A(n11456), .ZN(n12486) );
  OAI22_X1 U13235 ( .A1(n15821), .A2(n12487), .B1(n12486), .B2(n13959), .ZN(
        n11457) );
  AOI21_X1 U13236 ( .B1(n15814), .B2(n11488), .A(n11457), .ZN(n11458) );
  OAI211_X1 U13237 ( .C1(n11460), .C2(n14066), .A(n11459), .B(n11458), .ZN(
        P2_U3258) );
  XNOR2_X1 U13238 ( .A(n11461), .B(n13756), .ZN(n11523) );
  INV_X1 U13239 ( .A(n11523), .ZN(n11472) );
  OAI211_X1 U13240 ( .C1(n8131), .C2(n13756), .A(n14074), .B(n11462), .ZN(
        n11465) );
  NAND2_X1 U13241 ( .A1(n13806), .A2(n14071), .ZN(n11464) );
  NAND2_X1 U13242 ( .A1(n13808), .A2(n14069), .ZN(n11463) );
  AND2_X1 U13243 ( .A1(n11464), .A2(n11463), .ZN(n12585) );
  NAND2_X1 U13244 ( .A1(n11465), .A2(n12585), .ZN(n11521) );
  INV_X1 U13245 ( .A(n13587), .ZN(n12583) );
  INV_X1 U13246 ( .A(n11619), .ZN(n11466) );
  AOI211_X1 U13247 ( .C1(n13587), .C2(n11467), .A(n14076), .B(n11466), .ZN(
        n11522) );
  NAND2_X1 U13248 ( .A1(n11522), .A2(n15814), .ZN(n11469) );
  AOI22_X1 U13249 ( .A1(n15818), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n12588), 
        .B2(n15816), .ZN(n11468) );
  OAI211_X1 U13250 ( .C1(n12583), .C2(n15821), .A(n11469), .B(n11468), .ZN(
        n11470) );
  AOI21_X1 U13251 ( .B1(n7197), .B2(n11521), .A(n11470), .ZN(n11471) );
  OAI21_X1 U13252 ( .B1(n11472), .B2(n14085), .A(n11471), .ZN(P2_U3256) );
  INV_X1 U13253 ( .A(n15681), .ZN(n11486) );
  INV_X1 U13254 ( .A(n11473), .ZN(n11474) );
  AND2_X1 U13255 ( .A1(n11474), .A2(n11545), .ZN(n11475) );
  XNOR2_X1 U13256 ( .A(n7205), .B(n15685), .ZN(n11645) );
  XNOR2_X1 U13257 ( .A(n11645), .B(n11666), .ZN(n11479) );
  NAND2_X1 U13258 ( .A1(n11480), .A2(n11479), .ZN(n11648) );
  OAI211_X1 U13259 ( .C1(n11480), .C2(n11479), .A(n11648), .B(n15131), .ZN(
        n11485) );
  AOI21_X1 U13260 ( .B1(n12921), .B2(n12876), .A(n11481), .ZN(n11482) );
  OAI21_X1 U13261 ( .B1(n11794), .B2(n15126), .A(n11482), .ZN(n11483) );
  AOI21_X1 U13262 ( .B1(n15685), .B2(n12887), .A(n11483), .ZN(n11484) );
  OAI211_X1 U13263 ( .C1(n11486), .C2(n11990), .A(n11485), .B(n11484), .ZN(
        P3_U3179) );
  AOI211_X1 U13264 ( .C1(n15758), .C2(n11489), .A(n11488), .B(n11487), .ZN(
        n11565) );
  AOI22_X1 U13265 ( .A1(n14127), .A2(n13576), .B1(n15868), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11490) );
  OAI21_X1 U13266 ( .B1(n11565), .B2(n15868), .A(n11490), .ZN(P2_U3506) );
  INV_X1 U13267 ( .A(n11513), .ZN(n11492) );
  NAND2_X1 U13268 ( .A1(n11503), .A2(n15527), .ZN(n11491) );
  NAND2_X1 U13269 ( .A1(n11492), .A2(n11491), .ZN(n11500) );
  XNOR2_X1 U13270 ( .A(n11500), .B(n15529), .ZN(n11493) );
  INV_X1 U13271 ( .A(n14375), .ZN(n11494) );
  OAI21_X1 U13272 ( .B1(n11493), .B2(n15890), .A(n11494), .ZN(n11498) );
  OAI21_X1 U13273 ( .B1(n9436), .B2(n11494), .A(n15914), .ZN(n11495) );
  NAND2_X1 U13274 ( .A1(n11495), .A2(n15903), .ZN(n11497) );
  AND2_X1 U13275 ( .A1(n14374), .A2(n14765), .ZN(n11496) );
  AOI21_X1 U13276 ( .B1(n11498), .B2(n11497), .A(n11496), .ZN(n15569) );
  XNOR2_X1 U13277 ( .A(n11499), .B(n9436), .ZN(n15567) );
  INV_X1 U13278 ( .A(n11500), .ZN(n11501) );
  NAND2_X1 U13279 ( .A1(n11501), .A2(n15917), .ZN(n15564) );
  INV_X1 U13280 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14383) );
  OAI22_X1 U13281 ( .A1(n14772), .A2(n10367), .B1(n14383), .B2(n14584), .ZN(
        n11502) );
  AOI21_X1 U13282 ( .B1(n15931), .B2(n11503), .A(n11502), .ZN(n11504) );
  OAI21_X1 U13283 ( .B1(n14672), .B2(n15564), .A(n11504), .ZN(n11505) );
  AOI21_X1 U13284 ( .B1(n15936), .B2(n15567), .A(n11505), .ZN(n11506) );
  OAI21_X1 U13285 ( .B1(n15941), .B2(n15569), .A(n11506), .ZN(P1_U3292) );
  OAI21_X1 U13286 ( .B1(n11508), .B2(n11518), .A(n11507), .ZN(n11511) );
  INV_X1 U13287 ( .A(n11509), .ZN(n11510) );
  AOI21_X1 U13288 ( .B1(n11511), .B2(n15914), .A(n11510), .ZN(n15595) );
  OAI211_X1 U13289 ( .C1(n11513), .C2(n15596), .A(n11512), .B(n15917), .ZN(
        n15594) );
  NOR2_X1 U13290 ( .A1(n14672), .A2(n15594), .ZN(n11515) );
  INV_X1 U13291 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14395) );
  OAI22_X1 U13292 ( .A1(n14772), .A2(n10366), .B1(n14395), .B2(n14584), .ZN(
        n11514) );
  AOI211_X1 U13293 ( .C1(n15931), .C2(n11516), .A(n11515), .B(n11514), .ZN(
        n11520) );
  XOR2_X1 U13294 ( .A(n11518), .B(n11517), .Z(n15599) );
  NAND2_X1 U13295 ( .A1(n15599), .A2(n15936), .ZN(n11519) );
  OAI211_X1 U13296 ( .C1(n15941), .C2(n15595), .A(n11520), .B(n11519), .ZN(
        P1_U3291) );
  AOI211_X1 U13297 ( .C1(n11523), .C2(n15859), .A(n11522), .B(n11521), .ZN(
        n11574) );
  AOI22_X1 U13298 ( .A1(n14127), .A2(n13587), .B1(n15868), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11524) );
  OAI21_X1 U13299 ( .B1(n11574), .B2(n15868), .A(n11524), .ZN(P2_U3508) );
  OR2_X1 U13300 ( .A1(n11526), .A2(n11525), .ZN(n15588) );
  AOI21_X2 U13301 ( .B1(n15733), .B2(n15588), .A(n15690), .ZN(n13252) );
  INV_X1 U13302 ( .A(n13252), .ZN(n11689) );
  XNOR2_X1 U13303 ( .A(n11527), .B(n11528), .ZN(n15615) );
  INV_X1 U13304 ( .A(n15615), .ZN(n11539) );
  AOI21_X1 U13305 ( .B1(n11529), .B2(n11528), .A(n13240), .ZN(n11534) );
  OAI22_X1 U13306 ( .A1(n11531), .A2(n15575), .B1(n11530), .B2(n13243), .ZN(
        n11532) );
  AOI21_X1 U13307 ( .B1(n11534), .B2(n11533), .A(n11532), .ZN(n15612) );
  INV_X1 U13308 ( .A(n15612), .ZN(n11537) );
  NOR2_X1 U13309 ( .A1(n15688), .A2(n7490), .ZN(n11536) );
  OAI22_X1 U13310 ( .A1(n13250), .A2(n15613), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n13143), .ZN(n11535) );
  AOI211_X1 U13311 ( .C1(n11537), .C2(n15688), .A(n11536), .B(n11535), .ZN(
        n11538) );
  OAI21_X1 U13312 ( .B1(n11689), .B2(n11539), .A(n11538), .ZN(P3_U3230) );
  XNOR2_X1 U13313 ( .A(n7634), .B(n11540), .ZN(n15630) );
  OAI211_X1 U13314 ( .C1(n11542), .C2(n7634), .A(n11541), .B(n15577), .ZN(
        n11544) );
  OR2_X1 U13315 ( .A1(n15574), .A2(n15575), .ZN(n11543) );
  OAI211_X1 U13316 ( .C1(n11545), .C2(n13243), .A(n11544), .B(n11543), .ZN(
        n15627) );
  AOI22_X1 U13317 ( .A1(n15684), .A2(n15628), .B1(n15680), .B2(n11546), .ZN(
        n11547) );
  OAI21_X1 U13318 ( .B1(n10818), .B2(n15688), .A(n11547), .ZN(n11548) );
  AOI21_X1 U13319 ( .B1(n15627), .B2(n15688), .A(n11548), .ZN(n11549) );
  OAI21_X1 U13320 ( .B1(n11689), .B2(n15630), .A(n11549), .ZN(P3_U3229) );
  AOI22_X1 U13321 ( .A1(n15814), .A2(n11550), .B1(n13514), .B2(n15816), .ZN(
        n11551) );
  OAI21_X1 U13322 ( .B1(n11558), .B2(n15821), .A(n11551), .ZN(n11554) );
  MUX2_X1 U13323 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11552), .S(n7197), .Z(
        n11553) );
  AOI211_X1 U13324 ( .C1(n15824), .C2(n11555), .A(n11554), .B(n11553), .ZN(
        n11556) );
  INV_X1 U13325 ( .A(n11556), .ZN(P2_U3259) );
  INV_X1 U13326 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11557) );
  OAI22_X1 U13327 ( .A1(n14219), .A2(n11558), .B1(n14215), .B2(n11557), .ZN(
        n11559) );
  INV_X1 U13328 ( .A(n11559), .ZN(n11560) );
  OAI21_X1 U13329 ( .B1(n11561), .B2(n15870), .A(n11560), .ZN(P2_U3448) );
  INV_X1 U13330 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11562) );
  OAI22_X1 U13331 ( .A1(n14219), .A2(n12487), .B1(n14215), .B2(n11562), .ZN(
        n11563) );
  INV_X1 U13332 ( .A(n11563), .ZN(n11564) );
  OAI21_X1 U13333 ( .B1(n11565), .B2(n15870), .A(n11564), .ZN(P2_U3451) );
  INV_X1 U13334 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11566) );
  OAI22_X1 U13335 ( .A1(n14219), .A2(n11567), .B1(n14215), .B2(n11566), .ZN(
        n11568) );
  INV_X1 U13336 ( .A(n11568), .ZN(n11569) );
  OAI21_X1 U13337 ( .B1(n11570), .B2(n15870), .A(n11569), .ZN(P2_U3445) );
  INV_X1 U13338 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11571) );
  OAI22_X1 U13339 ( .A1(n14219), .A2(n12583), .B1(n14215), .B2(n11571), .ZN(
        n11572) );
  INV_X1 U13340 ( .A(n11572), .ZN(n11573) );
  OAI21_X1 U13341 ( .B1(n11574), .B2(n15870), .A(n11573), .ZN(P2_U3457) );
  INV_X1 U13342 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11575) );
  OAI22_X1 U13343 ( .A1(n14219), .A2(n11576), .B1(n14215), .B2(n11575), .ZN(
        n11577) );
  AOI21_X1 U13344 ( .B1(n11578), .B2(n14215), .A(n11577), .ZN(n11579) );
  INV_X1 U13345 ( .A(n11579), .ZN(P2_U3439) );
  NAND2_X1 U13346 ( .A1(n11580), .A2(n11587), .ZN(n11582) );
  NAND2_X1 U13347 ( .A1(n11582), .A2(n11581), .ZN(n11585) );
  INV_X1 U13348 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15894) );
  NOR2_X1 U13349 ( .A1(n14505), .A2(n15894), .ZN(n11583) );
  AOI21_X1 U13350 ( .B1(n14505), .B2(n15894), .A(n11583), .ZN(n11584) );
  NOR2_X1 U13351 ( .A1(n11584), .A2(n11585), .ZN(n14504) );
  AOI211_X1 U13352 ( .C1(n11585), .C2(n11584), .A(n14504), .B(n14548), .ZN(
        n11596) );
  AOI21_X1 U13353 ( .B1(n11588), .B2(n11587), .A(n11586), .ZN(n11591) );
  INV_X1 U13354 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14511) );
  NOR2_X1 U13355 ( .A1(n14512), .A2(n14511), .ZN(n11589) );
  AOI21_X1 U13356 ( .B1(n14511), .B2(n14512), .A(n11589), .ZN(n11590) );
  NAND2_X1 U13357 ( .A1(n11590), .A2(n11591), .ZN(n14510) );
  OAI211_X1 U13358 ( .C1(n11591), .C2(n11590), .A(n14553), .B(n14510), .ZN(
        n11594) );
  NAND2_X1 U13359 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14297)
         );
  INV_X1 U13360 ( .A(n14297), .ZN(n11592) );
  AOI21_X1 U13361 ( .B1(n14521), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11592), 
        .ZN(n11593) );
  OAI211_X1 U13362 ( .C1(n14518), .C2(n14512), .A(n11594), .B(n11593), .ZN(
        n11595) );
  OR2_X1 U13363 ( .A1(n11596), .A2(n11595), .ZN(P1_U3259) );
  NAND2_X1 U13364 ( .A1(n14371), .A2(n7192), .ZN(n11600) );
  NAND2_X1 U13365 ( .A1(n11716), .A2(n10994), .ZN(n11599) );
  NAND2_X1 U13366 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  XNOR2_X1 U13367 ( .A(n11601), .B(n11634), .ZN(n11627) );
  NAND2_X1 U13368 ( .A1(n14371), .A2(n11435), .ZN(n11603) );
  NAND2_X1 U13369 ( .A1(n11716), .A2(n7192), .ZN(n11602) );
  NAND2_X1 U13370 ( .A1(n11603), .A2(n11602), .ZN(n11626) );
  INV_X1 U13371 ( .A(n11626), .ZN(n11628) );
  XNOR2_X1 U13372 ( .A(n11627), .B(n11628), .ZN(n11604) );
  XNOR2_X1 U13373 ( .A(n11631), .B(n11604), .ZN(n11610) );
  NAND2_X1 U13374 ( .A1(n14372), .A2(n14767), .ZN(n11605) );
  OAI21_X1 U13375 ( .B1(n11633), .B2(n15901), .A(n11605), .ZN(n15660) );
  AOI22_X1 U13376 ( .A1(n15960), .A2(n15660), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11607) );
  NAND2_X1 U13377 ( .A1(n15965), .A2(n11716), .ZN(n11606) );
  OAI211_X1 U13378 ( .C1(n15969), .C2(n11608), .A(n11607), .B(n11606), .ZN(
        n11609) );
  AOI21_X1 U13379 ( .B1(n11610), .B2(n15963), .A(n11609), .ZN(n11611) );
  INV_X1 U13380 ( .A(n11611), .ZN(P1_U3227) );
  XNOR2_X1 U13381 ( .A(n11612), .B(n11614), .ZN(n11692) );
  INV_X1 U13382 ( .A(n11692), .ZN(n11625) );
  OAI211_X1 U13383 ( .C1(n11615), .C2(n11614), .A(n11613), .B(n14074), .ZN(
        n11618) );
  NAND2_X1 U13384 ( .A1(n13805), .A2(n14071), .ZN(n11617) );
  NAND2_X1 U13385 ( .A1(n13807), .A2(n14069), .ZN(n11616) );
  AND2_X1 U13386 ( .A1(n11617), .A2(n11616), .ZN(n12574) );
  NAND2_X1 U13387 ( .A1(n11618), .A2(n12574), .ZN(n11690) );
  INV_X1 U13388 ( .A(n13591), .ZN(n11622) );
  AOI211_X1 U13389 ( .C1(n13591), .C2(n11619), .A(n14076), .B(n11818), .ZN(
        n11691) );
  NAND2_X1 U13390 ( .A1(n11691), .A2(n15814), .ZN(n11621) );
  AOI22_X1 U13391 ( .A1(n15818), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12571), 
        .B2(n15816), .ZN(n11620) );
  OAI211_X1 U13392 ( .C1(n11622), .C2(n15821), .A(n11621), .B(n11620), .ZN(
        n11623) );
  AOI21_X1 U13393 ( .B1(n7197), .B2(n11690), .A(n11623), .ZN(n11624) );
  OAI21_X1 U13394 ( .B1(n11625), .B2(n14085), .A(n11624), .ZN(P2_U3255) );
  NOR2_X1 U13395 ( .A1(n11627), .A2(n11626), .ZN(n11630) );
  INV_X1 U13396 ( .A(n11627), .ZN(n11629) );
  OAI22_X1 U13397 ( .A1(n11631), .A2(n11630), .B1(n11629), .B2(n11628), .ZN(
        n11758) );
  NAND2_X1 U13398 ( .A1(n11780), .A2(n10994), .ZN(n11632) );
  OAI21_X1 U13399 ( .B1(n11633), .B2(n12640), .A(n11632), .ZN(n11635) );
  XNOR2_X1 U13400 ( .A(n11635), .B(n11198), .ZN(n11637) );
  AOI22_X1 U13401 ( .A1(n14370), .A2(n11435), .B1(n11780), .B2(n7192), .ZN(
        n11636) );
  NOR2_X1 U13402 ( .A1(n11637), .A2(n11636), .ZN(n11759) );
  NAND2_X1 U13403 ( .A1(n11637), .A2(n11636), .ZN(n11757) );
  INV_X1 U13404 ( .A(n11757), .ZN(n11638) );
  NOR2_X1 U13405 ( .A1(n11759), .A2(n11638), .ZN(n11639) );
  XNOR2_X1 U13406 ( .A(n11758), .B(n11639), .ZN(n11644) );
  NAND2_X1 U13407 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n14428) );
  OAI21_X1 U13408 ( .B1(n15942), .B2(n11764), .A(n14428), .ZN(n11642) );
  INV_X1 U13409 ( .A(n14371), .ZN(n11640) );
  INV_X1 U13410 ( .A(n11780), .ZN(n15692) );
  OAI22_X1 U13411 ( .A1(n15945), .A2(n11640), .B1(n15692), .B2(n14348), .ZN(
        n11641) );
  AOI211_X1 U13412 ( .C1(n11779), .C2(n14352), .A(n11642), .B(n11641), .ZN(
        n11643) );
  OAI21_X1 U13413 ( .B1(n11644), .B2(n15949), .A(n11643), .ZN(P1_U3239) );
  INV_X1 U13414 ( .A(n11671), .ZN(n11658) );
  INV_X1 U13415 ( .A(n11645), .ZN(n11646) );
  OR2_X1 U13416 ( .A1(n11666), .A2(n11646), .ZN(n11647) );
  NAND2_X1 U13417 ( .A1(n11648), .A2(n11647), .ZN(n11651) );
  XNOR2_X1 U13418 ( .A(n11649), .B(n12802), .ZN(n11741) );
  XNOR2_X1 U13419 ( .A(n11794), .B(n11741), .ZN(n11650) );
  NAND2_X1 U13420 ( .A1(n11651), .A2(n11650), .ZN(n11743) );
  OAI211_X1 U13421 ( .C1(n11651), .C2(n11650), .A(n11743), .B(n15131), .ZN(
        n11657) );
  NAND2_X1 U13422 ( .A1(n12920), .A2(n12876), .ZN(n11654) );
  INV_X1 U13423 ( .A(n11652), .ZN(n11653) );
  OAI211_X1 U13424 ( .C1(n11879), .C2(n15126), .A(n11654), .B(n11653), .ZN(
        n11655) );
  AOI21_X1 U13425 ( .B1(n15701), .B2(n12887), .A(n11655), .ZN(n11656) );
  OAI211_X1 U13426 ( .C1(n11658), .C2(n11990), .A(n11657), .B(n11656), .ZN(
        P3_U3153) );
  INV_X1 U13427 ( .A(n15588), .ZN(n11659) );
  NAND2_X1 U13428 ( .A1(n15688), .A2(n11659), .ZN(n13195) );
  INV_X1 U13429 ( .A(n13195), .ZN(n15682) );
  AOI21_X1 U13430 ( .B1(n15632), .B2(n15688), .A(n15682), .ZN(n13135) );
  XNOR2_X1 U13431 ( .A(n11660), .B(n11661), .ZN(n15697) );
  INV_X1 U13432 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11670) );
  NAND2_X1 U13433 ( .A1(n11663), .A2(n11662), .ZN(n11665) );
  AOI21_X1 U13434 ( .B1(n11665), .B2(n11664), .A(n13240), .ZN(n11669) );
  OAI22_X1 U13435 ( .A1(n11666), .A2(n15575), .B1(n11879), .B2(n13243), .ZN(
        n11667) );
  AOI21_X1 U13436 ( .B1(n11669), .B2(n11668), .A(n11667), .ZN(n15698) );
  MUX2_X1 U13437 ( .A(n11670), .B(n15698), .S(n15688), .Z(n11673) );
  AOI22_X1 U13438 ( .A1(n15684), .A2(n15701), .B1(n15680), .B2(n11671), .ZN(
        n11672) );
  OAI211_X1 U13439 ( .C1(n13135), .C2(n15697), .A(n11673), .B(n11672), .ZN(
        P3_U3226) );
  INV_X1 U13440 ( .A(n11674), .ZN(n11676) );
  INV_X1 U13441 ( .A(n14523), .ZN(n14530) );
  OAI222_X1 U13442 ( .A1(n14897), .A2(n11675), .B1(n14893), .B2(n11676), .C1(
        P1_U3086), .C2(n14530), .ZN(P1_U3338) );
  INV_X1 U13443 ( .A(n15174), .ZN(n15168) );
  OAI222_X1 U13444 ( .A1(n14244), .A2(n11677), .B1(n14239), .B2(n11676), .C1(
        P2_U3088), .C2(n15168), .ZN(P2_U3310) );
  XNOR2_X1 U13445 ( .A(n11678), .B(n11681), .ZN(n15645) );
  OR2_X1 U13446 ( .A1(n11680), .A2(n11679), .ZN(n11730) );
  OAI21_X1 U13447 ( .B1(n11682), .B2(n11681), .A(n11730), .ZN(n11683) );
  INV_X1 U13448 ( .A(n13243), .ZN(n15545) );
  AOI222_X1 U13449 ( .A1(n15577), .A2(n11683), .B1(n12920), .B2(n15545), .C1(
        n12922), .C2(n15547), .ZN(n15646) );
  MUX2_X1 U13450 ( .A(n11684), .B(n15646), .S(n15688), .Z(n11688) );
  AOI22_X1 U13451 ( .A1(n15684), .A2(n11686), .B1(n15680), .B2(n11685), .ZN(
        n11687) );
  OAI211_X1 U13452 ( .C1(n11689), .C2(n15645), .A(n11688), .B(n11687), .ZN(
        P3_U3228) );
  AOI211_X1 U13453 ( .C1(n11692), .C2(n15859), .A(n11691), .B(n11690), .ZN(
        n11697) );
  AOI22_X1 U13454 ( .A1(n14127), .A2(n13591), .B1(n15868), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11693) );
  OAI21_X1 U13455 ( .B1(n11697), .B2(n15868), .A(n11693), .ZN(P2_U3509) );
  INV_X1 U13456 ( .A(n14219), .ZN(n12151) );
  INV_X1 U13457 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11694) );
  NOR2_X1 U13458 ( .A1(n14215), .A2(n11694), .ZN(n11695) );
  AOI21_X1 U13459 ( .B1(n12151), .B2(n13591), .A(n11695), .ZN(n11696) );
  OAI21_X1 U13460 ( .B1(n11697), .B2(n15870), .A(n11696), .ZN(P2_U3460) );
  NAND2_X1 U13461 ( .A1(n14372), .A2(n11712), .ZN(n11698) );
  NAND2_X1 U13462 ( .A1(n15657), .A2(n15658), .ZN(n11702) );
  INV_X1 U13463 ( .A(n11716), .ZN(n15668) );
  NAND2_X1 U13464 ( .A1(n15668), .A2(n14371), .ZN(n11701) );
  NAND2_X1 U13465 ( .A1(n11702), .A2(n11701), .ZN(n11783) );
  NAND2_X1 U13466 ( .A1(n11783), .A2(n11784), .ZN(n11704) );
  NAND2_X1 U13467 ( .A1(n15692), .A2(n14370), .ZN(n11703) );
  NAND2_X1 U13468 ( .A1(n11763), .A2(n11764), .ZN(n11705) );
  OAI211_X1 U13469 ( .C1(n11707), .C2(n11706), .A(n15914), .B(n12034), .ZN(
        n11708) );
  AOI22_X1 U13470 ( .A1(n14369), .A2(n14767), .B1(n14765), .B2(n14367), .ZN(
        n11872) );
  NAND2_X1 U13471 ( .A1(n11708), .A2(n11872), .ZN(n15747) );
  INV_X1 U13472 ( .A(n15747), .ZN(n11726) );
  NAND2_X1 U13473 ( .A1(n14372), .A2(n11709), .ZN(n11710) );
  NAND2_X1 U13474 ( .A1(n11711), .A2(n11710), .ZN(n11715) );
  NAND2_X1 U13475 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  NAND2_X1 U13476 ( .A1(n11715), .A2(n11714), .ZN(n15652) );
  NAND2_X1 U13477 ( .A1(n14371), .A2(n11716), .ZN(n11775) );
  AND2_X1 U13478 ( .A1(n11777), .A2(n11775), .ZN(n11717) );
  AOI22_X1 U13479 ( .A1(n15705), .A2(n15710), .B1(n15722), .B2(n11764), .ZN(
        n11719) );
  NAND2_X1 U13480 ( .A1(n11719), .A2(n11718), .ZN(n12046) );
  OAI21_X1 U13481 ( .B1(n11719), .B2(n11718), .A(n12046), .ZN(n15745) );
  INV_X1 U13482 ( .A(n15745), .ZN(n15748) );
  INV_X1 U13483 ( .A(n15742), .ZN(n12045) );
  AND2_X1 U13484 ( .A1(n15656), .A2(n15668), .ZN(n15654) );
  NAND2_X1 U13485 ( .A1(n15654), .A2(n15692), .ZN(n15706) );
  NAND2_X1 U13486 ( .A1(n15707), .A2(n15742), .ZN(n11720) );
  NAND2_X1 U13487 ( .A1(n11720), .A2(n15917), .ZN(n11721) );
  NOR2_X1 U13488 ( .A1(n15766), .A2(n11721), .ZN(n15741) );
  NAND2_X1 U13489 ( .A1(n15741), .A2(n15935), .ZN(n11723) );
  AOI22_X1 U13490 ( .A1(n15941), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11869), 
        .B2(n15930), .ZN(n11722) );
  OAI211_X1 U13491 ( .C1(n12045), .C2(n15723), .A(n11723), .B(n11722), .ZN(
        n11724) );
  AOI21_X1 U13492 ( .B1(n15748), .B2(n15936), .A(n11724), .ZN(n11725) );
  OAI21_X1 U13493 ( .B1(n15941), .B2(n11726), .A(n11725), .ZN(P1_U3285) );
  XNOR2_X1 U13494 ( .A(n11727), .B(n11732), .ZN(n11738) );
  AND2_X1 U13495 ( .A1(n11730), .A2(n11728), .ZN(n11733) );
  NAND2_X1 U13496 ( .A1(n11730), .A2(n11729), .ZN(n11731) );
  OAI211_X1 U13497 ( .C1(n11733), .C2(n11732), .A(n11731), .B(n15577), .ZN(
        n11735) );
  AOI22_X1 U13498 ( .A1(n12921), .A2(n15547), .B1(n15545), .B2(n12919), .ZN(
        n11734) );
  OAI211_X1 U13499 ( .C1(n15733), .C2(n11738), .A(n11735), .B(n11734), .ZN(
        n11736) );
  INV_X1 U13500 ( .A(n11736), .ZN(n15689) );
  OAI21_X1 U13501 ( .B1(n11737), .B2(n15797), .A(n15689), .ZN(n15677) );
  INV_X1 U13502 ( .A(n15677), .ZN(n11740) );
  INV_X1 U13503 ( .A(n11738), .ZN(n15683) );
  NOR2_X1 U13504 ( .A1(n15980), .A2(n15732), .ZN(n13330) );
  AOI22_X1 U13505 ( .A1(n15683), .A2(n13330), .B1(P3_REG0_REG_6__SCAN_IN), 
        .B2(n15980), .ZN(n11739) );
  OAI21_X1 U13506 ( .B1(n11740), .B2(n15980), .A(n11739), .ZN(P3_U3408) );
  INV_X1 U13507 ( .A(n11797), .ZN(n11752) );
  NAND2_X1 U13508 ( .A1(n11741), .A2(n12919), .ZN(n11742) );
  NAND2_X1 U13509 ( .A1(n11743), .A2(n11742), .ZN(n11745) );
  XNOR2_X1 U13510 ( .A(n7205), .B(n15736), .ZN(n11877) );
  XNOR2_X1 U13511 ( .A(n11877), .B(n11879), .ZN(n11744) );
  NAND2_X1 U13512 ( .A1(n11745), .A2(n11744), .ZN(n11881) );
  OAI211_X1 U13513 ( .C1(n11745), .C2(n11744), .A(n11881), .B(n15131), .ZN(
        n11751) );
  NAND2_X1 U13514 ( .A1(n12876), .A2(n12919), .ZN(n11748) );
  INV_X1 U13515 ( .A(n11746), .ZN(n11747) );
  OAI211_X1 U13516 ( .C1(n11978), .C2(n15126), .A(n11748), .B(n11747), .ZN(
        n11749) );
  AOI21_X1 U13517 ( .B1(n15736), .B2(n12887), .A(n11749), .ZN(n11750) );
  OAI211_X1 U13518 ( .C1(n11752), .C2(n11990), .A(n11751), .B(n11750), .ZN(
        P3_U3161) );
  INV_X1 U13519 ( .A(SI_24_), .ZN(n11755) );
  INV_X1 U13520 ( .A(n11753), .ZN(n11754) );
  OAI222_X1 U13521 ( .A1(P3_U3151), .A2(n11756), .B1(n13403), .B2(n11755), 
        .C1(n13402), .C2(n11754), .ZN(P3_U3271) );
  NAND2_X1 U13522 ( .A1(n11758), .A2(n11757), .ZN(n11761) );
  NAND2_X1 U13523 ( .A1(n11761), .A2(n11760), .ZN(n11769) );
  INV_X1 U13524 ( .A(n11769), .ZN(n11766) );
  NOR2_X1 U13525 ( .A1(n11764), .A2(n12706), .ZN(n11762) );
  AOI21_X1 U13526 ( .B1(n11763), .B2(n7192), .A(n11762), .ZN(n11866) );
  OAI22_X1 U13527 ( .A1(n15722), .A2(n12708), .B1(n11764), .B2(n12640), .ZN(
        n11765) );
  XNOR2_X1 U13528 ( .A(n11765), .B(n11634), .ZN(n11864) );
  XOR2_X1 U13529 ( .A(n11866), .B(n11864), .Z(n11767) );
  AOI21_X1 U13530 ( .B1(n11766), .B2(n11767), .A(n15949), .ZN(n11770) );
  NAND2_X1 U13531 ( .A1(n11769), .A2(n11768), .ZN(n11865) );
  NAND2_X1 U13532 ( .A1(n11770), .A2(n11865), .ZN(n11773) );
  AOI22_X1 U13533 ( .A1(n14767), .A2(n14370), .B1(n14368), .B2(n14765), .ZN(
        n15711) );
  INV_X1 U13534 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n14442) );
  OAI22_X1 U13535 ( .A1(n15711), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14442), .ZN(n11771) );
  AOI21_X1 U13536 ( .B1(n15720), .B2(n14352), .A(n11771), .ZN(n11772) );
  OAI211_X1 U13537 ( .C1(n15722), .C2(n14348), .A(n11773), .B(n11772), .ZN(
        P1_U3213) );
  AND2_X1 U13538 ( .A1(n11774), .A2(n11775), .ZN(n11778) );
  OAI21_X1 U13539 ( .B1(n11778), .B2(n11777), .A(n11776), .ZN(n15695) );
  OAI211_X1 U13540 ( .C1(n15654), .C2(n15692), .A(n15917), .B(n15706), .ZN(
        n15691) );
  NAND2_X1 U13541 ( .A1(n15930), .A2(n11779), .ZN(n11782) );
  NAND2_X1 U13542 ( .A1(n15931), .A2(n11780), .ZN(n11781) );
  OAI211_X1 U13543 ( .C1(n15691), .C2(n14672), .A(n11782), .B(n11781), .ZN(
        n11789) );
  XNOR2_X1 U13544 ( .A(n11783), .B(n11784), .ZN(n11787) );
  NAND2_X1 U13545 ( .A1(n15695), .A2(n15749), .ZN(n11786) );
  AOI22_X1 U13546 ( .A1(n14369), .A2(n14765), .B1(n14767), .B2(n14371), .ZN(
        n11785) );
  OAI211_X1 U13547 ( .C1(n15890), .C2(n11787), .A(n11786), .B(n11785), .ZN(
        n15693) );
  MUX2_X1 U13548 ( .A(n15693), .B(P1_REG2_REG_6__SCAN_IN), .S(n15941), .Z(
        n11788) );
  AOI211_X1 U13549 ( .C1(n15784), .C2(n15695), .A(n11789), .B(n11788), .ZN(
        n11790) );
  INV_X1 U13550 ( .A(n11790), .ZN(P1_U3287) );
  AOI21_X1 U13551 ( .B1(n11796), .B2(n11792), .A(n9753), .ZN(n11793) );
  OAI222_X1 U13552 ( .A1(n13243), .A2(n11978), .B1(n15575), .B2(n11794), .C1(
        n13240), .C2(n11793), .ZN(n15734) );
  INV_X1 U13553 ( .A(n15734), .ZN(n11803) );
  XOR2_X1 U13554 ( .A(n11795), .B(n11796), .Z(n15731) );
  INV_X1 U13555 ( .A(n15731), .ZN(n11801) );
  AOI22_X1 U13556 ( .A1(n15684), .A2(n15736), .B1(n15680), .B2(n11797), .ZN(
        n11798) );
  OAI21_X1 U13557 ( .B1(n11799), .B2(n15688), .A(n11798), .ZN(n11800) );
  AOI21_X1 U13558 ( .B1(n11801), .B2(n13252), .A(n11800), .ZN(n11802) );
  OAI21_X1 U13559 ( .B1(n11803), .B2(n15690), .A(n11802), .ZN(P3_U3225) );
  XNOR2_X1 U13560 ( .A(n11804), .B(n13761), .ZN(n11912) );
  INV_X1 U13561 ( .A(n11912), .ZN(n11814) );
  OAI211_X1 U13562 ( .C1(n8132), .C2(n13761), .A(n14074), .B(n11805), .ZN(
        n11808) );
  NAND2_X1 U13563 ( .A1(n13803), .A2(n14071), .ZN(n11807) );
  NAND2_X1 U13564 ( .A1(n13805), .A2(n14069), .ZN(n11806) );
  AND2_X1 U13565 ( .A1(n11807), .A2(n11806), .ZN(n11844) );
  NAND2_X1 U13566 ( .A1(n11808), .A2(n11844), .ZN(n11910) );
  INV_X1 U13567 ( .A(n13603), .ZN(n11845) );
  AOI21_X1 U13568 ( .B1(n11819), .B2(n13603), .A(n14076), .ZN(n11809) );
  AND2_X1 U13569 ( .A1(n11809), .A2(n12009), .ZN(n11911) );
  NAND2_X1 U13570 ( .A1(n11911), .A2(n15814), .ZN(n11811) );
  AOI22_X1 U13571 ( .A1(n15818), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11848), 
        .B2(n15816), .ZN(n11810) );
  OAI211_X1 U13572 ( .C1(n11845), .C2(n15821), .A(n11811), .B(n11810), .ZN(
        n11812) );
  AOI21_X1 U13573 ( .B1(n11910), .B2(n7197), .A(n11812), .ZN(n11813) );
  OAI21_X1 U13574 ( .B1(n11814), .B2(n14085), .A(n11813), .ZN(P2_U3253) );
  OAI222_X1 U13575 ( .A1(P3_U3151), .A2(n11816), .B1(n13403), .B2(n15017), 
        .C1(n13402), .C2(n11815), .ZN(P3_U3270) );
  XOR2_X1 U13576 ( .A(n13760), .B(n11817), .Z(n15825) );
  INV_X1 U13577 ( .A(n11818), .ZN(n11821) );
  INV_X1 U13578 ( .A(n11819), .ZN(n11820) );
  AOI211_X1 U13579 ( .C1(n13600), .C2(n11821), .A(n14076), .B(n11820), .ZN(
        n15815) );
  OAI21_X1 U13580 ( .B1(n8138), .B2(n8802), .A(n11822), .ZN(n11825) );
  OAI22_X1 U13581 ( .A1(n11824), .A2(n14057), .B1(n11823), .B2(n14055), .ZN(
        n12520) );
  AOI21_X1 U13582 ( .B1(n11825), .B2(n14074), .A(n12520), .ZN(n15827) );
  INV_X1 U13583 ( .A(n15827), .ZN(n11826) );
  AOI211_X1 U13584 ( .C1(n15859), .C2(n15825), .A(n15815), .B(n11826), .ZN(
        n11831) );
  AOI22_X1 U13585 ( .A1(n13600), .A2(n14127), .B1(n15868), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11827) );
  OAI21_X1 U13586 ( .B1(n11831), .B2(n15868), .A(n11827), .ZN(P2_U3510) );
  INV_X1 U13587 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11828) );
  OAI22_X1 U13588 ( .A1(n15822), .A2(n14219), .B1(n14215), .B2(n11828), .ZN(
        n11829) );
  INV_X1 U13589 ( .A(n11829), .ZN(n11830) );
  OAI21_X1 U13590 ( .B1(n11831), .B2(n15870), .A(n11830), .ZN(P2_U3463) );
  NOR2_X1 U13591 ( .A1(n12589), .A2(n11832), .ZN(n11833) );
  XNOR2_X1 U13592 ( .A(n13587), .B(n12728), .ZN(n12576) );
  NAND2_X1 U13593 ( .A1(n14076), .A2(n13807), .ZN(n11834) );
  XNOR2_X1 U13594 ( .A(n12576), .B(n11834), .ZN(n12590) );
  INV_X1 U13595 ( .A(n12575), .ZN(n11837) );
  INV_X1 U13596 ( .A(n11834), .ZN(n11835) );
  XNOR2_X1 U13597 ( .A(n13591), .B(n12728), .ZN(n12523) );
  NAND2_X1 U13598 ( .A1(n14076), .A2(n13806), .ZN(n11838) );
  XNOR2_X1 U13599 ( .A(n12523), .B(n11838), .ZN(n12577) );
  INV_X1 U13600 ( .A(n11838), .ZN(n11839) );
  NOR2_X1 U13601 ( .A1(n12523), .A2(n11839), .ZN(n11840) );
  XNOR2_X1 U13602 ( .A(n13600), .B(n12728), .ZN(n11849) );
  NAND2_X1 U13603 ( .A1(n14076), .A2(n13805), .ZN(n11841) );
  INV_X1 U13604 ( .A(n11841), .ZN(n11842) );
  XNOR2_X1 U13605 ( .A(n13603), .B(n12728), .ZN(n11938) );
  NAND2_X1 U13606 ( .A1(n14076), .A2(n13804), .ZN(n11931) );
  XNOR2_X1 U13607 ( .A(n11938), .B(n11931), .ZN(n11850) );
  INV_X1 U13608 ( .A(n13479), .ZN(n13515) );
  INV_X1 U13609 ( .A(n13513), .ZN(n13492) );
  OAI22_X1 U13610 ( .A1(n13492), .A2(n11844), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11843), .ZN(n11847) );
  NOR2_X1 U13611 ( .A1(n11845), .A2(n13506), .ZN(n11846) );
  AOI211_X1 U13612 ( .C1(n13515), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n11854) );
  AOI22_X1 U13613 ( .A1(n11849), .A2(n13507), .B1(n13428), .B2(n13805), .ZN(
        n11851) );
  OR3_X1 U13614 ( .A1(n11852), .A2(n11851), .A3(n11850), .ZN(n11853) );
  OAI211_X1 U13615 ( .C1(n11933), .C2(n13486), .A(n11854), .B(n11853), .ZN(
        P2_U3196) );
  XNOR2_X1 U13616 ( .A(n11855), .B(n11858), .ZN(n11856) );
  OAI222_X1 U13617 ( .A1(n13243), .A2(n12143), .B1(n15575), .B2(n11879), .C1(
        n13240), .C2(n11856), .ZN(n11918) );
  INV_X1 U13618 ( .A(n11918), .ZN(n11862) );
  XNOR2_X1 U13619 ( .A(n11857), .B(n11858), .ZN(n11919) );
  INV_X1 U13620 ( .A(n13135), .ZN(n12170) );
  INV_X1 U13621 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U13622 ( .A1(n15684), .A2(n11876), .B1(n15680), .B2(n11890), .ZN(
        n11859) );
  OAI21_X1 U13623 ( .B1(n12944), .B2(n15688), .A(n11859), .ZN(n11860) );
  AOI21_X1 U13624 ( .B1(n11919), .B2(n12170), .A(n11860), .ZN(n11861) );
  OAI21_X1 U13625 ( .B1(n11862), .B2(n15690), .A(n11861), .ZN(P3_U3224) );
  OAI22_X1 U13626 ( .A1(n12045), .A2(n12708), .B1(n12044), .B2(n12640), .ZN(
        n11863) );
  XNOR2_X1 U13627 ( .A(n11863), .B(n11634), .ZN(n11945) );
  OAI22_X1 U13628 ( .A1(n12045), .A2(n12640), .B1(n12044), .B2(n12706), .ZN(
        n11944) );
  XNOR2_X1 U13629 ( .A(n11945), .B(n11944), .ZN(n11868) );
  AOI21_X1 U13630 ( .B1(n11868), .B2(n11867), .A(n11946), .ZN(n11875) );
  NAND2_X1 U13631 ( .A1(n14352), .A2(n11869), .ZN(n11871) );
  OAI211_X1 U13632 ( .C1(n11872), .C2(n14326), .A(n11871), .B(n11870), .ZN(
        n11873) );
  AOI21_X1 U13633 ( .B1(n15742), .B2(n15965), .A(n11873), .ZN(n11874) );
  OAI21_X1 U13634 ( .B1(n11875), .B2(n15949), .A(n11874), .ZN(P1_U3221) );
  XNOR2_X1 U13635 ( .A(n11876), .B(n12802), .ZN(n11979) );
  XNOR2_X1 U13636 ( .A(n11979), .B(n11978), .ZN(n11886) );
  INV_X1 U13637 ( .A(n11877), .ZN(n11878) );
  OR2_X1 U13638 ( .A1(n11879), .A2(n11878), .ZN(n11880) );
  NAND2_X1 U13639 ( .A1(n11881), .A2(n11880), .ZN(n11885) );
  INV_X1 U13640 ( .A(n11886), .ZN(n11882) );
  INV_X1 U13641 ( .A(n11981), .ZN(n11884) );
  AOI21_X1 U13642 ( .B1(n11886), .B2(n11885), .A(n11884), .ZN(n11892) );
  NAND2_X1 U13643 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15397) );
  OAI21_X1 U13644 ( .B1(n12143), .B2(n15126), .A(n15397), .ZN(n11887) );
  AOI21_X1 U13645 ( .B1(n12876), .B2(n12918), .A(n11887), .ZN(n11888) );
  OAI21_X1 U13646 ( .B1(n15128), .B2(n11924), .A(n11888), .ZN(n11889) );
  AOI21_X1 U13647 ( .B1(n11890), .B2(n12900), .A(n11889), .ZN(n11891) );
  OAI21_X1 U13648 ( .B1(n11892), .B2(n12890), .A(n11891), .ZN(P3_U3171) );
  NAND2_X1 U13649 ( .A1(n11893), .A2(n11897), .ZN(n11894) );
  NAND2_X1 U13650 ( .A1(n11895), .A2(n11894), .ZN(n15792) );
  INV_X1 U13651 ( .A(n15792), .ZN(n11905) );
  XNOR2_X1 U13652 ( .A(n11896), .B(n11897), .ZN(n11900) );
  OAI22_X1 U13653 ( .A1(n11978), .A2(n15575), .B1(n12157), .B2(n13243), .ZN(
        n11898) );
  AOI21_X1 U13654 ( .B1(n15792), .B2(n15632), .A(n11898), .ZN(n11899) );
  OAI21_X1 U13655 ( .B1(n11900), .B2(n13240), .A(n11899), .ZN(n15790) );
  NAND2_X1 U13656 ( .A1(n15790), .A2(n15688), .ZN(n11904) );
  INV_X1 U13657 ( .A(n11901), .ZN(n11991) );
  OAI22_X1 U13658 ( .A1(n13250), .A2(n15789), .B1(n11991), .B2(n13143), .ZN(
        n11902) );
  AOI21_X1 U13659 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15690), .A(n11902), 
        .ZN(n11903) );
  OAI211_X1 U13660 ( .C1(n11905), .C2(n13195), .A(n11904), .B(n11903), .ZN(
        P3_U3223) );
  INV_X1 U13661 ( .A(n11906), .ZN(n11908) );
  INV_X1 U13662 ( .A(n15175), .ZN(n15186) );
  OAI222_X1 U13663 ( .A1(n14244), .A2(n11907), .B1(n14239), .B2(n11908), .C1(
        n15186), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13664 ( .A(n14542), .ZN(n14535) );
  OAI222_X1 U13665 ( .A1(n14897), .A2(n11909), .B1(n14893), .B2(n11908), .C1(
        n14535), .C2(P1_U3086), .ZN(P1_U3337) );
  AOI211_X1 U13666 ( .C1(n15859), .C2(n11912), .A(n11911), .B(n11910), .ZN(
        n11917) );
  AOI22_X1 U13667 ( .A1(n13603), .A2(n14127), .B1(n15868), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11913) );
  OAI21_X1 U13668 ( .B1(n11917), .B2(n15868), .A(n11913), .ZN(P2_U3511) );
  INV_X1 U13669 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11914) );
  NOR2_X1 U13670 ( .A1(n14215), .A2(n11914), .ZN(n11915) );
  AOI21_X1 U13671 ( .B1(n13603), .B2(n12151), .A(n11915), .ZN(n11916) );
  OAI21_X1 U13672 ( .B1(n11917), .B2(n15870), .A(n11916), .ZN(P2_U3466) );
  AOI21_X1 U13673 ( .B1(n11919), .B2(n15802), .A(n11918), .ZN(n11927) );
  INV_X1 U13674 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11920) );
  OAI22_X1 U13675 ( .A1(n11924), .A2(n13391), .B1(n15978), .B2(n11920), .ZN(
        n11921) );
  INV_X1 U13676 ( .A(n11921), .ZN(n11922) );
  OAI21_X1 U13677 ( .B1(n11927), .B2(n15980), .A(n11922), .ZN(P3_U3417) );
  INV_X1 U13678 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11923) );
  OAI22_X1 U13679 ( .A1(n13316), .A2(n11924), .B1(n15839), .B2(n11923), .ZN(
        n11925) );
  INV_X1 U13680 ( .A(n11925), .ZN(n11926) );
  OAI21_X1 U13681 ( .B1(n11927), .B2(n15970), .A(n11926), .ZN(P3_U3468) );
  INV_X1 U13682 ( .A(n11928), .ZN(n11929) );
  OAI222_X1 U13683 ( .A1(n11930), .A2(P3_U3151), .B1(n13402), .B2(n11929), 
        .C1(n14927), .C2(n13403), .ZN(P3_U3269) );
  INV_X1 U13684 ( .A(n11931), .ZN(n11932) );
  XNOR2_X1 U13685 ( .A(n13612), .B(n12728), .ZN(n12498) );
  NAND2_X1 U13686 ( .A1(n14076), .A2(n13803), .ZN(n12293) );
  XNOR2_X1 U13687 ( .A(n12498), .B(n12293), .ZN(n11939) );
  NAND2_X1 U13688 ( .A1(n11934), .A2(n11939), .ZN(n12296) );
  AOI22_X1 U13689 ( .A1(n14071), .A2(n13802), .B1(n13804), .B2(n14069), .ZN(
        n12007) );
  OAI22_X1 U13690 ( .A1(n13492), .A2(n12007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11935), .ZN(n11937) );
  NOR2_X1 U13691 ( .A1(n7577), .A2(n13506), .ZN(n11936) );
  AOI211_X1 U13692 ( .C1(n13515), .C2(n12011), .A(n11937), .B(n11936), .ZN(
        n11943) );
  INV_X1 U13693 ( .A(n11933), .ZN(n11941) );
  AOI22_X1 U13694 ( .A1(n11938), .A2(n13507), .B1(n13428), .B2(n13804), .ZN(
        n11940) );
  OR3_X1 U13695 ( .A1(n11941), .A2(n11940), .A3(n11939), .ZN(n11942) );
  OAI211_X1 U13696 ( .C1(n12296), .C2(n13486), .A(n11943), .B(n11942), .ZN(
        P2_U3206) );
  NAND2_X1 U13697 ( .A1(n15781), .A2(n7192), .ZN(n11948) );
  NAND2_X1 U13698 ( .A1(n14367), .A2(n11435), .ZN(n11947) );
  NAND2_X1 U13699 ( .A1(n11948), .A2(n11947), .ZN(n12069) );
  NAND2_X1 U13700 ( .A1(n15781), .A2(n10994), .ZN(n11950) );
  NAND2_X1 U13701 ( .A1(n14367), .A2(n7192), .ZN(n11949) );
  NAND2_X1 U13702 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  XNOR2_X1 U13703 ( .A(n11951), .B(n11634), .ZN(n12070) );
  XOR2_X1 U13704 ( .A(n12069), .B(n12070), .Z(n11952) );
  XNOR2_X1 U13705 ( .A(n12068), .B(n11952), .ZN(n11956) );
  AOI22_X1 U13706 ( .A1(n14368), .A2(n14767), .B1(n14765), .B2(n14366), .ZN(
        n15770) );
  NAND2_X1 U13707 ( .A1(n14352), .A2(n15780), .ZN(n11953) );
  NAND2_X1 U13708 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14458) );
  OAI211_X1 U13709 ( .C1(n15770), .C2(n14326), .A(n11953), .B(n14458), .ZN(
        n11954) );
  AOI21_X1 U13710 ( .B1(n15781), .B2(n15965), .A(n11954), .ZN(n11955) );
  OAI21_X1 U13711 ( .B1(n11956), .B2(n15949), .A(n11955), .ZN(P1_U3231) );
  NAND2_X1 U13712 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n12360)
         );
  INV_X1 U13713 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14163) );
  XNOR2_X1 U13714 ( .A(n15174), .B(n14163), .ZN(n11962) );
  INV_X1 U13715 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11960) );
  XNOR2_X1 U13716 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n12033), .ZN(n12023) );
  OAI21_X1 U13717 ( .B1(n11383), .B2(n11969), .A(n11957), .ZN(n11958) );
  NAND2_X1 U13718 ( .A1(n11971), .A2(n11958), .ZN(n11959) );
  XNOR2_X1 U13719 ( .A(n15157), .B(n11958), .ZN(n15163) );
  NAND2_X1 U13720 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15163), .ZN(n15162) );
  NAND2_X1 U13721 ( .A1(n11959), .A2(n15162), .ZN(n12024) );
  NAND2_X1 U13722 ( .A1(n12023), .A2(n12024), .ZN(n12022) );
  OAI21_X1 U13723 ( .B1(n11960), .B2(n12033), .A(n12022), .ZN(n11961) );
  NAND2_X1 U13724 ( .A1(n11962), .A2(n11961), .ZN(n15172) );
  OAI211_X1 U13725 ( .C1(n11962), .C2(n11961), .A(n15172), .B(n15201), .ZN(
        n11963) );
  NAND2_X1 U13726 ( .A1(n12360), .A2(n11963), .ZN(n11964) );
  AOI21_X1 U13727 ( .B1(n15200), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11964), 
        .ZN(n11977) );
  NOR2_X1 U13728 ( .A1(n15168), .A2(n12376), .ZN(n11965) );
  AOI21_X1 U13729 ( .B1(n12376), .B2(n15168), .A(n11965), .ZN(n11975) );
  INV_X1 U13730 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11973) );
  NOR2_X1 U13731 ( .A1(n11973), .A2(n12033), .ZN(n11966) );
  AOI21_X1 U13732 ( .B1(n11973), .B2(n12033), .A(n11966), .ZN(n12026) );
  AOI21_X1 U13733 ( .B1(n11969), .B2(n11968), .A(n11967), .ZN(n11970) );
  NAND2_X1 U13734 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  NAND2_X1 U13735 ( .A1(n11972), .A2(n15160), .ZN(n12027) );
  NAND2_X1 U13736 ( .A1(n12026), .A2(n12027), .ZN(n12025) );
  OAI211_X1 U13737 ( .C1(n11975), .C2(n11974), .A(n15205), .B(n15167), .ZN(
        n11976) );
  OAI211_X1 U13738 ( .C1(n15158), .C2(n15168), .A(n11977), .B(n11976), .ZN(
        P2_U3231) );
  NAND2_X1 U13739 ( .A1(n11979), .A2(n11978), .ZN(n11980) );
  XNOR2_X1 U13740 ( .A(n11987), .B(n12802), .ZN(n12135) );
  XNOR2_X1 U13741 ( .A(n12135), .B(n12143), .ZN(n11982) );
  AOI21_X1 U13742 ( .B1(n11983), .B2(n11982), .A(n12890), .ZN(n11984) );
  NAND2_X1 U13743 ( .A1(n11984), .A2(n12136), .ZN(n11989) );
  NAND2_X1 U13744 ( .A1(n12876), .A2(n12917), .ZN(n11985) );
  NAND2_X1 U13745 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15415)
         );
  OAI211_X1 U13746 ( .C1(n12157), .C2(n15126), .A(n11985), .B(n15415), .ZN(
        n11986) );
  AOI21_X1 U13747 ( .B1(n11987), .B2(n12887), .A(n11986), .ZN(n11988) );
  OAI211_X1 U13748 ( .C1(n11991), .C2(n11990), .A(n11989), .B(n11988), .ZN(
        P3_U3157) );
  XNOR2_X1 U13749 ( .A(n11993), .B(n11992), .ZN(n11994) );
  OAI222_X1 U13750 ( .A1(n13243), .A2(n11995), .B1(n15575), .B2(n12143), .C1(
        n11994), .C2(n13240), .ZN(n15799) );
  INV_X1 U13751 ( .A(n15799), .ZN(n12001) );
  OAI21_X1 U13752 ( .B1(n11997), .B2(n12138), .A(n11996), .ZN(n15801) );
  AOI22_X1 U13753 ( .A1(n15690), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15680), 
        .B2(n12145), .ZN(n11998) );
  OAI21_X1 U13754 ( .B1(n15798), .B2(n13250), .A(n11998), .ZN(n11999) );
  AOI21_X1 U13755 ( .B1(n15801), .B2(n13252), .A(n11999), .ZN(n12000) );
  OAI21_X1 U13756 ( .B1(n12001), .B2(n15690), .A(n12000), .ZN(P3_U3222) );
  XNOR2_X1 U13757 ( .A(n12002), .B(n13762), .ZN(n12150) );
  INV_X1 U13758 ( .A(n12150), .ZN(n12016) );
  INV_X1 U13759 ( .A(n12003), .ZN(n12004) );
  AOI21_X1 U13760 ( .B1(n12006), .B2(n12005), .A(n12004), .ZN(n12008) );
  OAI21_X1 U13761 ( .B1(n12008), .B2(n14063), .A(n12007), .ZN(n12148) );
  AOI21_X1 U13762 ( .B1(n13612), .B2(n12009), .A(n14076), .ZN(n12010) );
  AND2_X1 U13763 ( .A1(n12010), .A2(n12059), .ZN(n12149) );
  NAND2_X1 U13764 ( .A1(n12149), .A2(n15814), .ZN(n12013) );
  AOI22_X1 U13765 ( .A1(n15818), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12011), 
        .B2(n15816), .ZN(n12012) );
  OAI211_X1 U13766 ( .C1(n7577), .C2(n15821), .A(n12013), .B(n12012), .ZN(
        n12014) );
  AOI21_X1 U13767 ( .B1(n12148), .B2(n7197), .A(n12014), .ZN(n12015) );
  OAI21_X1 U13768 ( .B1(n12016), .B2(n14085), .A(n12015), .ZN(P2_U3252) );
  INV_X1 U13769 ( .A(n12017), .ZN(n12020) );
  OAI222_X1 U13770 ( .A1(n14244), .A2(n12018), .B1(n14239), .B2(n12020), .C1(
        n13776), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U13771 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12021) );
  OAI222_X1 U13772 ( .A1(n14897), .A2(n12021), .B1(n14893), .B2(n12020), .C1(
        P1_U3086), .C2(n12019), .ZN(P1_U3336) );
  OAI211_X1 U13773 ( .C1(n12024), .C2(n12023), .A(n15201), .B(n12022), .ZN(
        n12029) );
  OAI211_X1 U13774 ( .C1(n12027), .C2(n12026), .A(n15205), .B(n12025), .ZN(
        n12028) );
  NAND2_X1 U13775 ( .A1(n12029), .A2(n12028), .ZN(n12031) );
  NAND2_X1 U13776 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n12304)
         );
  INV_X1 U13777 ( .A(n12304), .ZN(n12030) );
  AOI211_X1 U13778 ( .C1(n15200), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n12031), 
        .B(n12030), .ZN(n12032) );
  OAI21_X1 U13779 ( .B1(n15158), .B2(n12033), .A(n12032), .ZN(P2_U3230) );
  INV_X1 U13780 ( .A(n14367), .ZN(n12036) );
  NAND2_X1 U13781 ( .A1(n15781), .A2(n12036), .ZN(n12035) );
  NAND2_X1 U13782 ( .A1(n15769), .A2(n12035), .ZN(n12038) );
  OR2_X1 U13783 ( .A1(n15781), .A2(n12036), .ZN(n12037) );
  NAND2_X1 U13784 ( .A1(n12038), .A2(n12037), .ZN(n12099) );
  NAND2_X1 U13785 ( .A1(n12099), .A2(n12100), .ZN(n12040) );
  OR2_X1 U13786 ( .A1(n12119), .A2(n7989), .ZN(n12039) );
  NAND2_X1 U13787 ( .A1(n12040), .A2(n12039), .ZN(n12080) );
  XNOR2_X1 U13788 ( .A(n12080), .B(n12079), .ZN(n12041) );
  AOI22_X1 U13789 ( .A1(n14364), .A2(n14765), .B1(n14767), .B2(n14366), .ZN(
        n12232) );
  OAI21_X1 U13790 ( .B1(n12041), .B2(n15890), .A(n12232), .ZN(n15808) );
  INV_X1 U13791 ( .A(n15808), .ZN(n12053) );
  INV_X1 U13792 ( .A(n15781), .ZN(n15767) );
  INV_X1 U13793 ( .A(n12119), .ZN(n12103) );
  INV_X1 U13794 ( .A(n12087), .ZN(n12042) );
  AOI211_X1 U13795 ( .C1(n12234), .C2(n12102), .A(n14763), .B(n12042), .ZN(
        n15810) );
  AOI22_X1 U13796 ( .A1(n15941), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12230), 
        .B2(n15930), .ZN(n12043) );
  OAI21_X1 U13797 ( .B1(n7560), .B2(n15723), .A(n12043), .ZN(n12051) );
  NAND2_X1 U13798 ( .A1(n12046), .A2(n7267), .ZN(n15763) );
  INV_X1 U13799 ( .A(n12047), .ZN(n12048) );
  AND2_X1 U13800 ( .A1(n12049), .A2(n12079), .ZN(n15806) );
  NOR3_X1 U13801 ( .A1(n15807), .A2(n15806), .A3(n14740), .ZN(n12050) );
  AOI211_X1 U13802 ( .C1(n15935), .C2(n15810), .A(n12051), .B(n12050), .ZN(
        n12052) );
  OAI21_X1 U13803 ( .B1(n15941), .B2(n12053), .A(n12052), .ZN(P1_U3282) );
  XNOR2_X1 U13804 ( .A(n12054), .B(n13764), .ZN(n12055) );
  NAND2_X1 U13805 ( .A1(n12055), .A2(n14074), .ZN(n12057) );
  AOI22_X1 U13806 ( .A1(n13801), .A2(n14071), .B1(n13803), .B2(n14069), .ZN(
        n12056) );
  AND2_X1 U13807 ( .A1(n12057), .A2(n12056), .ZN(n15867) );
  XNOR2_X1 U13808 ( .A(n12058), .B(n13764), .ZN(n15860) );
  AOI21_X1 U13809 ( .B1(n15862), .B2(n12059), .A(n14076), .ZN(n12060) );
  NAND2_X1 U13810 ( .A1(n12060), .A2(n12191), .ZN(n15864) );
  AOI22_X1 U13811 ( .A1(n15818), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12494), 
        .B2(n15816), .ZN(n12062) );
  NAND2_X1 U13812 ( .A1(n15862), .A2(n14035), .ZN(n12061) );
  OAI211_X1 U13813 ( .C1(n15864), .C2(n13984), .A(n12062), .B(n12061), .ZN(
        n12063) );
  AOI21_X1 U13814 ( .B1(n15860), .B2(n15824), .A(n12063), .ZN(n12064) );
  OAI21_X1 U13815 ( .B1(n15867), .B2(n13980), .A(n12064), .ZN(P2_U3251) );
  INV_X1 U13816 ( .A(n12070), .ZN(n12066) );
  INV_X1 U13817 ( .A(n12069), .ZN(n12065) );
  NAND2_X1 U13818 ( .A1(n12070), .A2(n12069), .ZN(n12071) );
  NAND2_X1 U13819 ( .A1(n12072), .A2(n12071), .ZN(n12220) );
  OAI22_X1 U13820 ( .A1(n12103), .A2(n12708), .B1(n7989), .B2(n12640), .ZN(
        n12073) );
  XNOR2_X1 U13821 ( .A(n12073), .B(n11634), .ZN(n12223) );
  AND2_X1 U13822 ( .A1(n14366), .A2(n11435), .ZN(n12074) );
  AOI21_X1 U13823 ( .B1(n12119), .B2(n7192), .A(n12074), .ZN(n12221) );
  XNOR2_X1 U13824 ( .A(n12223), .B(n12221), .ZN(n12219) );
  XNOR2_X1 U13825 ( .A(n12220), .B(n12219), .ZN(n12078) );
  NAND2_X1 U13826 ( .A1(n14367), .A2(n14767), .ZN(n12116) );
  NAND2_X1 U13827 ( .A1(n14365), .A2(n14765), .ZN(n12114) );
  AND2_X1 U13828 ( .A1(n12116), .A2(n12114), .ZN(n12097) );
  NAND2_X1 U13829 ( .A1(n14352), .A2(n12118), .ZN(n12075) );
  NAND2_X1 U13830 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n14473)
         );
  OAI211_X1 U13831 ( .C1(n12097), .C2(n14326), .A(n12075), .B(n14473), .ZN(
        n12076) );
  AOI21_X1 U13832 ( .B1(n12119), .B2(n15965), .A(n12076), .ZN(n12077) );
  OAI21_X1 U13833 ( .B1(n12078), .B2(n15949), .A(n12077), .ZN(P1_U3217) );
  INV_X1 U13834 ( .A(n14365), .ZN(n12084) );
  NAND2_X1 U13835 ( .A1(n12080), .A2(n12079), .ZN(n12082) );
  OR2_X1 U13836 ( .A1(n12234), .A2(n12084), .ZN(n12081) );
  INV_X1 U13837 ( .A(n12085), .ZN(n12202) );
  XNOR2_X1 U13838 ( .A(n12203), .B(n12202), .ZN(n12083) );
  OAI222_X1 U13839 ( .A1(n15903), .A2(n12084), .B1(n15901), .B2(n12409), .C1(
        n12083), .C2(n15890), .ZN(n15831) );
  INV_X1 U13840 ( .A(n15831), .ZN(n12094) );
  OAI21_X1 U13841 ( .B1(n12086), .B2(n12085), .A(n12205), .ZN(n15832) );
  NAND2_X1 U13842 ( .A1(n12087), .A2(n12281), .ZN(n12088) );
  NAND2_X1 U13843 ( .A1(n12088), .A2(n15917), .ZN(n12089) );
  OR2_X1 U13844 ( .A1(n12211), .A2(n12089), .ZN(n15828) );
  AOI22_X1 U13845 ( .A1(n15941), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12290), 
        .B2(n15930), .ZN(n12091) );
  NAND2_X1 U13846 ( .A1(n12281), .A2(n15931), .ZN(n12090) );
  OAI211_X1 U13847 ( .C1(n15828), .C2(n14672), .A(n12091), .B(n12090), .ZN(
        n12092) );
  AOI21_X1 U13848 ( .B1(n15832), .B2(n15936), .A(n12092), .ZN(n12093) );
  OAI21_X1 U13849 ( .B1(n15941), .B2(n12094), .A(n12093), .ZN(P1_U3281) );
  INV_X1 U13850 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n12107) );
  XOR2_X1 U13851 ( .A(n12100), .B(n12095), .Z(n12123) );
  INV_X1 U13852 ( .A(n12123), .ZN(n12096) );
  NAND2_X1 U13853 ( .A1(n12096), .A2(n15923), .ZN(n12105) );
  INV_X1 U13854 ( .A(n12097), .ZN(n12098) );
  AOI21_X1 U13855 ( .B1(n12119), .B2(n15887), .A(n12098), .ZN(n12104) );
  XNOR2_X1 U13856 ( .A(n12099), .B(n7982), .ZN(n12101) );
  NAND2_X1 U13857 ( .A1(n12101), .A2(n15914), .ZN(n12117) );
  OAI211_X1 U13858 ( .C1(n15764), .C2(n12103), .A(n15917), .B(n12102), .ZN(
        n12113) );
  NAND4_X1 U13859 ( .A1(n12105), .A2(n12104), .A3(n12117), .A4(n12113), .ZN(
        n12108) );
  NAND2_X1 U13860 ( .A1(n12108), .A2(n15719), .ZN(n12106) );
  OAI21_X1 U13861 ( .B1(n15719), .B2(n12107), .A(n12106), .ZN(P1_U3489) );
  INV_X1 U13862 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n12110) );
  NAND2_X1 U13863 ( .A1(n12108), .A2(n15717), .ZN(n12109) );
  OAI21_X1 U13864 ( .B1(n15717), .B2(n12110), .A(n12109), .ZN(P1_U3538) );
  INV_X1 U13865 ( .A(n12111), .ZN(n12130) );
  OAI222_X1 U13866 ( .A1(n14897), .A2(n12112), .B1(n14893), .B2(n12130), .C1(
        n15536), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI211_X1 U13867 ( .C1(n12123), .C2(n12115), .A(n12114), .B(n12113), .ZN(
        n12126) );
  AOI21_X1 U13868 ( .B1(n12117), .B2(n12116), .A(n15941), .ZN(n12125) );
  AOI22_X1 U13869 ( .A1(n15941), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12118), 
        .B2(n15930), .ZN(n12121) );
  NAND2_X1 U13870 ( .A1(n12119), .A2(n15931), .ZN(n12120) );
  OAI211_X1 U13871 ( .C1(n12123), .C2(n12122), .A(n12121), .B(n12120), .ZN(
        n12124) );
  AOI211_X1 U13872 ( .C1(n15935), .C2(n12126), .A(n12125), .B(n12124), .ZN(
        n12127) );
  INV_X1 U13873 ( .A(n12127), .ZN(P1_U3283) );
  INV_X1 U13874 ( .A(n12128), .ZN(n12129) );
  INV_X1 U13875 ( .A(SI_27_), .ZN(n15029) );
  OAI222_X1 U13876 ( .A1(P3_U3151), .A2(n12955), .B1(n13402), .B2(n12129), 
        .C1(n15029), .C2(n13403), .ZN(P3_U3268) );
  OAI222_X1 U13877 ( .A1(n14244), .A2(n12131), .B1(P2_U3088), .B2(n13736), 
        .C1(n14239), .C2(n12130), .ZN(P2_U3307) );
  INV_X1 U13878 ( .A(n12132), .ZN(n12133) );
  OAI222_X1 U13879 ( .A1(P3_U3151), .A2(n12134), .B1(n13402), .B2(n12133), 
        .C1(n14919), .C2(n13403), .ZN(P3_U3267) );
  AND2_X1 U13880 ( .A1(n7326), .A2(n12137), .ZN(n12139) );
  MUX2_X1 U13881 ( .A(n12139), .B(n12138), .S(n12802), .Z(n12140) );
  NAND2_X1 U13882 ( .A1(n12141), .A2(n12140), .ZN(n12174) );
  OAI211_X1 U13883 ( .C1(n12141), .C2(n12140), .A(n12174), .B(n15131), .ZN(
        n12147) );
  NAND2_X1 U13884 ( .A1(n12895), .A2(n12914), .ZN(n12142) );
  NAND2_X1 U13885 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n15430)
         );
  OAI211_X1 U13886 ( .C1(n12143), .C2(n12897), .A(n12142), .B(n15430), .ZN(
        n12144) );
  AOI21_X1 U13887 ( .B1(n12900), .B2(n12145), .A(n12144), .ZN(n12146) );
  OAI211_X1 U13888 ( .C1(n15128), .C2(n15798), .A(n12147), .B(n12146), .ZN(
        P3_U3176) );
  AOI211_X1 U13889 ( .C1(n15859), .C2(n12150), .A(n12149), .B(n12148), .ZN(
        n12154) );
  AOI22_X1 U13890 ( .A1(n13612), .A2(n12151), .B1(P2_REG0_REG_13__SCAN_IN), 
        .B2(n15870), .ZN(n12152) );
  OAI21_X1 U13891 ( .B1(n12154), .B2(n15870), .A(n12152), .ZN(P2_U3469) );
  AOI22_X1 U13892 ( .A1(n13612), .A2(n14127), .B1(P2_REG1_REG_13__SCAN_IN), 
        .B2(n15868), .ZN(n12153) );
  OAI21_X1 U13893 ( .B1(n12154), .B2(n15868), .A(n12153), .ZN(P2_U3512) );
  XNOR2_X1 U13894 ( .A(n12155), .B(n12175), .ZN(n12156) );
  OAI222_X1 U13895 ( .A1(n13243), .A2(n12780), .B1(n15575), .B2(n12157), .C1(
        n13240), .C2(n12156), .ZN(n12273) );
  INV_X1 U13896 ( .A(n12273), .ZN(n12163) );
  OAI21_X1 U13897 ( .B1(n12159), .B2(n12175), .A(n12158), .ZN(n12274) );
  AOI22_X1 U13898 ( .A1(n15690), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15680), 
        .B2(n12179), .ZN(n12160) );
  OAI21_X1 U13899 ( .B1(n12280), .B2(n13250), .A(n12160), .ZN(n12161) );
  AOI21_X1 U13900 ( .B1(n12274), .B2(n13252), .A(n12161), .ZN(n12162) );
  OAI21_X1 U13901 ( .B1(n12163), .B2(n15690), .A(n12162), .ZN(P3_U3221) );
  XOR2_X1 U13902 ( .A(n12350), .B(n12164), .Z(n12165) );
  AOI222_X1 U13903 ( .A1(n15577), .A2(n12165), .B1(n12912), .B2(n15545), .C1(
        n12914), .C2(n15547), .ZN(n12325) );
  OAI21_X1 U13904 ( .B1(n12167), .B2(n12350), .A(n12166), .ZN(n15834) );
  AOI22_X1 U13905 ( .A1(n15690), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15680), 
        .B2(n12355), .ZN(n12168) );
  OAI21_X1 U13906 ( .B1(n12738), .B2(n13250), .A(n12168), .ZN(n12169) );
  AOI21_X1 U13907 ( .B1(n15834), .B2(n12170), .A(n12169), .ZN(n12171) );
  OAI21_X1 U13908 ( .B1(n12325), .B2(n15690), .A(n12171), .ZN(P3_U3220) );
  MUX2_X1 U13909 ( .A(n7326), .B(n12172), .S(n11039), .Z(n12173) );
  XNOR2_X1 U13910 ( .A(n12175), .B(n11039), .ZN(n12348) );
  XNOR2_X1 U13911 ( .A(n12349), .B(n12348), .ZN(n12181) );
  NOR2_X1 U13912 ( .A1(n15128), .A2(n12280), .ZN(n12178) );
  NAND2_X1 U13913 ( .A1(n12876), .A2(n12915), .ZN(n12176) );
  NAND2_X1 U13914 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15447)
         );
  OAI211_X1 U13915 ( .C1(n12780), .C2(n15126), .A(n12176), .B(n15447), .ZN(
        n12177) );
  AOI211_X1 U13916 ( .C1(n12179), .C2(n12900), .A(n12178), .B(n12177), .ZN(
        n12180) );
  OAI21_X1 U13917 ( .B1(n12181), .B2(n12890), .A(n12180), .ZN(P3_U3164) );
  NAND2_X1 U13918 ( .A1(n12182), .A2(n12186), .ZN(n12183) );
  NAND2_X1 U13919 ( .A1(n12184), .A2(n12183), .ZN(n12313) );
  INV_X1 U13920 ( .A(n12313), .ZN(n12198) );
  XNOR2_X1 U13921 ( .A(n12185), .B(n12186), .ZN(n12189) );
  NAND2_X1 U13922 ( .A1(n12313), .A2(n14060), .ZN(n12188) );
  AOI22_X1 U13923 ( .A1(n13800), .A2(n14071), .B1(n14069), .B2(n13802), .ZN(
        n12187) );
  OAI211_X1 U13924 ( .C1(n12189), .C2(n14063), .A(n12188), .B(n12187), .ZN(
        n12317) );
  NAND2_X1 U13925 ( .A1(n12317), .A2(n7197), .ZN(n12197) );
  OAI22_X1 U13926 ( .A1(n7197), .A2(n12190), .B1(n12341), .B2(n13959), .ZN(
        n12195) );
  NAND2_X1 U13927 ( .A1(n13622), .A2(n12191), .ZN(n12192) );
  NAND2_X1 U13928 ( .A1(n12192), .A2(n13976), .ZN(n12193) );
  OR2_X1 U13929 ( .A1(n12386), .A2(n12193), .ZN(n12314) );
  NOR2_X1 U13930 ( .A1(n12314), .A2(n13984), .ZN(n12194) );
  AOI211_X1 U13931 ( .C1(n14035), .C2(n13622), .A(n12195), .B(n12194), .ZN(
        n12196) );
  OAI211_X1 U13932 ( .C1(n12198), .C2(n14066), .A(n12197), .B(n12196), .ZN(
        P2_U3250) );
  INV_X1 U13933 ( .A(n12199), .ZN(n12200) );
  OAI222_X1 U13934 ( .A1(P3_U3151), .A2(n12201), .B1(n13402), .B2(n12200), 
        .C1(n15026), .C2(n13403), .ZN(P3_U3266) );
  XNOR2_X1 U13935 ( .A(n12411), .B(n12410), .ZN(n15840) );
  OR2_X1 U13936 ( .A1(n15941), .A2(n15890), .ZN(n14779) );
  NAND2_X1 U13937 ( .A1(n12205), .A2(n12204), .ZN(n12400) );
  XNOR2_X1 U13938 ( .A(n12400), .B(n12410), .ZN(n15846) );
  NAND2_X1 U13939 ( .A1(n15846), .A2(n15936), .ZN(n12215) );
  NAND2_X1 U13940 ( .A1(n14362), .A2(n14765), .ZN(n12207) );
  NAND2_X1 U13941 ( .A1(n14364), .A2(n14767), .ZN(n12206) );
  AND2_X1 U13942 ( .A1(n12207), .A2(n12206), .ZN(n15841) );
  INV_X1 U13943 ( .A(n15841), .ZN(n12208) );
  AOI22_X1 U13944 ( .A1(n12208), .A2(n14772), .B1(n12253), .B2(n15930), .ZN(
        n12209) );
  OAI21_X1 U13945 ( .B1(n12210), .B2(n14772), .A(n12209), .ZN(n12213) );
  NAND2_X1 U13946 ( .A1(n12211), .A2(n15843), .ZN(n12420) );
  OAI211_X1 U13947 ( .C1(n12211), .C2(n15843), .A(n12420), .B(n15917), .ZN(
        n15842) );
  NOR2_X1 U13948 ( .A1(n15842), .A2(n14672), .ZN(n12212) );
  AOI211_X1 U13949 ( .C1(n15931), .C2(n12408), .A(n12213), .B(n12212), .ZN(
        n12214) );
  OAI211_X1 U13950 ( .C1(n15840), .C2(n14779), .A(n12215), .B(n12214), .ZN(
        P1_U3280) );
  INV_X1 U13951 ( .A(n12216), .ZN(n12475) );
  OAI222_X1 U13952 ( .A1(n14897), .A2(n12217), .B1(n14893), .B2(n12475), .C1(
        P1_U3086), .C2(n8905), .ZN(P1_U3334) );
  AOI22_X1 U13953 ( .A1(n12234), .A2(n10994), .B1(n7192), .B2(n14365), .ZN(
        n12218) );
  XNOR2_X1 U13954 ( .A(n12218), .B(n11634), .ZN(n12240) );
  AOI22_X1 U13955 ( .A1(n12234), .A2(n7192), .B1(n11435), .B2(n14365), .ZN(
        n12241) );
  XNOR2_X1 U13956 ( .A(n12240), .B(n12241), .ZN(n12229) );
  NAND2_X1 U13957 ( .A1(n12220), .A2(n12219), .ZN(n12227) );
  INV_X1 U13958 ( .A(n12221), .ZN(n12222) );
  NAND2_X1 U13959 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U13960 ( .A1(n12227), .A2(n12224), .ZN(n12228) );
  INV_X1 U13961 ( .A(n12229), .ZN(n12225) );
  AND2_X1 U13962 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  NAND2_X1 U13963 ( .A1(n12227), .A2(n12226), .ZN(n12245) );
  INV_X1 U13964 ( .A(n12245), .ZN(n12284) );
  AOI21_X1 U13965 ( .B1(n12229), .B2(n12228), .A(n12284), .ZN(n12236) );
  NAND2_X1 U13966 ( .A1(n14352), .A2(n12230), .ZN(n12231) );
  NAND2_X1 U13967 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14488)
         );
  OAI211_X1 U13968 ( .C1(n12232), .C2(n14326), .A(n12231), .B(n14488), .ZN(
        n12233) );
  AOI21_X1 U13969 ( .B1(n12234), .B2(n15965), .A(n12233), .ZN(n12235) );
  OAI21_X1 U13970 ( .B1(n12236), .B2(n15949), .A(n12235), .ZN(P1_U3236) );
  NOR2_X1 U13971 ( .A1(n12237), .A2(n12706), .ZN(n12238) );
  AOI21_X1 U13972 ( .B1(n12281), .B2(n7192), .A(n12238), .ZN(n12247) );
  AOI22_X1 U13973 ( .A1(n12281), .A2(n10994), .B1(n7192), .B2(n14364), .ZN(
        n12239) );
  XNOR2_X1 U13974 ( .A(n12239), .B(n11634), .ZN(n12246) );
  XNOR2_X1 U13975 ( .A(n12246), .B(n12247), .ZN(n12282) );
  INV_X1 U13976 ( .A(n12240), .ZN(n12243) );
  INV_X1 U13977 ( .A(n12241), .ZN(n12242) );
  NOR2_X1 U13978 ( .A1(n12243), .A2(n12242), .ZN(n12283) );
  NOR2_X1 U13979 ( .A1(n12282), .A2(n12283), .ZN(n12244) );
  NAND2_X1 U13980 ( .A1(n12245), .A2(n12244), .ZN(n12285) );
  OAI21_X1 U13981 ( .B1(n12247), .B2(n12246), .A(n12285), .ZN(n12596) );
  OAI22_X1 U13982 ( .A1(n15843), .A2(n12708), .B1(n12409), .B2(n12640), .ZN(
        n12248) );
  XNOR2_X1 U13983 ( .A(n12248), .B(n11634), .ZN(n12597) );
  NOR2_X1 U13984 ( .A1(n12409), .A2(n12706), .ZN(n12249) );
  AOI21_X1 U13985 ( .B1(n12408), .B2(n7192), .A(n12249), .ZN(n12598) );
  XNOR2_X1 U13986 ( .A(n12597), .B(n12598), .ZN(n12595) );
  XNOR2_X1 U13987 ( .A(n12596), .B(n12595), .ZN(n12255) );
  OAI22_X1 U13988 ( .A1(n15841), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12250), .ZN(n12252) );
  NOR2_X1 U13989 ( .A1(n15843), .A2(n14348), .ZN(n12251) );
  AOI211_X1 U13990 ( .C1(n14352), .C2(n12253), .A(n12252), .B(n12251), .ZN(
        n12254) );
  OAI21_X1 U13991 ( .B1(n12255), .B2(n15949), .A(n12254), .ZN(P1_U3234) );
  INV_X1 U13992 ( .A(n12256), .ZN(n12261) );
  NOR2_X1 U13993 ( .A1(n12257), .A2(P2_U3088), .ZN(n13782) );
  AOI21_X1 U13994 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14234), .A(n13782), 
        .ZN(n12258) );
  OAI21_X1 U13995 ( .B1(n12261), .B2(n14239), .A(n12258), .ZN(P2_U3304) );
  AOI21_X1 U13996 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n14880), .A(n12259), 
        .ZN(n12260) );
  OAI21_X1 U13997 ( .B1(n12261), .B2(n14893), .A(n12260), .ZN(P1_U3332) );
  OAI211_X1 U13998 ( .C1(n12263), .C2(n9843), .A(n15577), .B(n12262), .ZN(
        n12265) );
  AOI22_X1 U13999 ( .A1(n12913), .A2(n15547), .B1(n15545), .B2(n12911), .ZN(
        n12264) );
  NAND2_X1 U14000 ( .A1(n12265), .A2(n12264), .ZN(n13312) );
  INV_X1 U14001 ( .A(n13312), .ZN(n12272) );
  OAI21_X1 U14002 ( .B1(n12268), .B2(n12267), .A(n12266), .ZN(n13313) );
  AOI22_X1 U14003 ( .A1(n15690), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15680), 
        .B2(n12783), .ZN(n12269) );
  OAI21_X1 U14004 ( .B1(n13390), .B2(n13250), .A(n12269), .ZN(n12270) );
  AOI21_X1 U14005 ( .B1(n13313), .B2(n13252), .A(n12270), .ZN(n12271) );
  OAI21_X1 U14006 ( .B1(n12272), .B2(n15690), .A(n12271), .ZN(P3_U3219) );
  INV_X1 U14007 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12275) );
  AOI21_X1 U14008 ( .B1(n15802), .B2(n12274), .A(n12273), .ZN(n12277) );
  MUX2_X1 U14009 ( .A(n12275), .B(n12277), .S(n15839), .Z(n12276) );
  OAI21_X1 U14010 ( .B1(n13316), .B2(n12280), .A(n12276), .ZN(P3_U3471) );
  INV_X1 U14011 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12278) );
  MUX2_X1 U14012 ( .A(n12278), .B(n12277), .S(n15978), .Z(n12279) );
  OAI21_X1 U14013 ( .B1(n13391), .B2(n12280), .A(n12279), .ZN(P3_U3426) );
  INV_X1 U14014 ( .A(n12281), .ZN(n15829) );
  OAI21_X1 U14015 ( .B1(n12284), .B2(n12283), .A(n12282), .ZN(n12286) );
  NAND3_X1 U14016 ( .A1(n12286), .A2(n15963), .A3(n12285), .ZN(n12292) );
  NAND2_X1 U14017 ( .A1(n14345), .A2(n14365), .ZN(n12288) );
  OAI211_X1 U14018 ( .C1(n15942), .C2(n12409), .A(n12288), .B(n12287), .ZN(
        n12289) );
  AOI21_X1 U14019 ( .B1(n12290), .B2(n14352), .A(n12289), .ZN(n12291) );
  OAI211_X1 U14020 ( .C1(n15829), .C2(n14348), .A(n12292), .B(n12291), .ZN(
        P1_U3224) );
  NAND2_X1 U14021 ( .A1(n14076), .A2(n13802), .ZN(n12297) );
  INV_X1 U14022 ( .A(n12297), .ZN(n12300) );
  XNOR2_X1 U14023 ( .A(n15862), .B(n12728), .ZN(n12299) );
  INV_X1 U14024 ( .A(n12293), .ZN(n12294) );
  NAND2_X1 U14025 ( .A1(n12296), .A2(n12295), .ZN(n12298) );
  XNOR2_X1 U14026 ( .A(n12299), .B(n12297), .ZN(n12499) );
  NAND2_X1 U14027 ( .A1(n12298), .A2(n12499), .ZN(n12493) );
  XNOR2_X1 U14028 ( .A(n13622), .B(n12728), .ZN(n12307) );
  AND2_X1 U14029 ( .A1(n13801), .A2(n14076), .ZN(n12301) );
  NAND2_X1 U14030 ( .A1(n12307), .A2(n12301), .ZN(n12302) );
  OAI21_X1 U14031 ( .B1(n12307), .B2(n12301), .A(n12302), .ZN(n12343) );
  INV_X1 U14032 ( .A(n12302), .ZN(n12303) );
  XNOR2_X1 U14033 ( .A(n13626), .B(n11109), .ZN(n12363) );
  NAND2_X1 U14034 ( .A1(n13800), .A2(n14076), .ZN(n12358) );
  XNOR2_X1 U14035 ( .A(n12363), .B(n12358), .ZN(n12309) );
  AOI22_X1 U14036 ( .A1(n13439), .A2(n13801), .B1(n13438), .B2(n14070), .ZN(
        n12305) );
  OAI211_X1 U14037 ( .C1(n12396), .C2(n13479), .A(n12305), .B(n12304), .ZN(
        n12306) );
  AOI21_X1 U14038 ( .B1(n13626), .B2(n13516), .A(n12306), .ZN(n12312) );
  NAND3_X1 U14039 ( .A1(n12307), .A2(n13428), .A3(n13801), .ZN(n12308) );
  OAI21_X1 U14040 ( .B1(n7463), .B2(n13486), .A(n12308), .ZN(n12310) );
  NAND2_X1 U14041 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  OAI211_X1 U14042 ( .C1(n12366), .C2(n13486), .A(n12312), .B(n12311), .ZN(
        P2_U3198) );
  INV_X1 U14043 ( .A(n13622), .ZN(n12323) );
  INV_X1 U14044 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U14045 ( .A1(n12313), .A2(n15758), .ZN(n12315) );
  NAND2_X1 U14046 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  NOR2_X1 U14047 ( .A1(n12317), .A2(n12316), .ZN(n12320) );
  MUX2_X1 U14048 ( .A(n12318), .B(n12320), .S(n14215), .Z(n12319) );
  OAI21_X1 U14049 ( .B1(n12323), .B2(n14219), .A(n12319), .ZN(P2_U3475) );
  INV_X1 U14050 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n12321) );
  MUX2_X1 U14051 ( .A(n12321), .B(n12320), .S(n15869), .Z(n12322) );
  OAI21_X1 U14052 ( .B1(n12323), .B2(n14165), .A(n12322), .ZN(P2_U3514) );
  NAND2_X1 U14053 ( .A1(n15834), .A2(n15632), .ZN(n12324) );
  OAI211_X1 U14054 ( .C1(n12738), .C2(n15797), .A(n12325), .B(n12324), .ZN(
        n15836) );
  INV_X1 U14055 ( .A(n15836), .ZN(n12327) );
  AOI22_X1 U14056 ( .A1(n15834), .A2(n13330), .B1(P3_REG0_REG_13__SCAN_IN), 
        .B2(n15980), .ZN(n12326) );
  OAI21_X1 U14057 ( .B1(n12327), .B2(n15980), .A(n12326), .ZN(P3_U3429) );
  OAI211_X1 U14058 ( .C1(n12330), .C2(n12329), .A(n12328), .B(n15577), .ZN(
        n12332) );
  AOI22_X1 U14059 ( .A1(n13225), .A2(n15545), .B1(n15547), .B2(n12912), .ZN(
        n12331) );
  NAND2_X1 U14060 ( .A1(n12332), .A2(n12331), .ZN(n13308) );
  INV_X1 U14061 ( .A(n13308), .ZN(n12339) );
  OAI21_X1 U14062 ( .B1(n12335), .B2(n12334), .A(n12333), .ZN(n13309) );
  AOI22_X1 U14063 ( .A1(n15690), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15680), 
        .B2(n12901), .ZN(n12336) );
  OAI21_X1 U14064 ( .B1(n13386), .B2(n13250), .A(n12336), .ZN(n12337) );
  AOI21_X1 U14065 ( .B1(n13309), .B2(n13252), .A(n12337), .ZN(n12338) );
  OAI21_X1 U14066 ( .B1(n12339), .B2(n15690), .A(n12338), .ZN(P3_U3218) );
  AOI22_X1 U14067 ( .A1(n13438), .A2(n13800), .B1(n13439), .B2(n13802), .ZN(
        n12340) );
  NAND2_X1 U14068 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15156)
         );
  OAI211_X1 U14069 ( .C1(n13479), .C2(n12341), .A(n12340), .B(n15156), .ZN(
        n12346) );
  AOI211_X1 U14070 ( .C1(n12344), .C2(n12343), .A(n13486), .B(n12342), .ZN(
        n12345) );
  AOI211_X1 U14071 ( .C1(n13622), .C2(n13516), .A(n12346), .B(n12345), .ZN(
        n12347) );
  INV_X1 U14072 ( .A(n12347), .ZN(P2_U3213) );
  MUX2_X2 U14073 ( .A(n12914), .B(n12349), .S(n12348), .Z(n12352) );
  XNOR2_X1 U14074 ( .A(n12350), .B(n12802), .ZN(n12351) );
  OAI211_X1 U14075 ( .C1(n12352), .C2(n12351), .A(n12741), .B(n15131), .ZN(
        n12357) );
  NAND2_X1 U14076 ( .A1(n12876), .A2(n12914), .ZN(n12353) );
  NAND2_X1 U14077 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_U3151), .ZN(n15463)
         );
  OAI211_X1 U14078 ( .C1(n12898), .C2(n15126), .A(n12353), .B(n15463), .ZN(
        n12354) );
  AOI21_X1 U14079 ( .B1(n12900), .B2(n12355), .A(n12354), .ZN(n12356) );
  OAI211_X1 U14080 ( .C1(n15128), .C2(n12738), .A(n12357), .B(n12356), .ZN(
        P3_U3174) );
  XNOR2_X1 U14081 ( .A(n13635), .B(n12728), .ZN(n12531) );
  NOR2_X1 U14082 ( .A1(n13501), .A2(n13976), .ZN(n12532) );
  XNOR2_X1 U14083 ( .A(n12531), .B(n12532), .ZN(n12365) );
  INV_X1 U14084 ( .A(n12535), .ZN(n12369) );
  AOI22_X1 U14085 ( .A1(n13439), .A2(n13800), .B1(n13438), .B2(n13799), .ZN(
        n12361) );
  OAI211_X1 U14086 ( .C1(n12375), .C2(n13479), .A(n12361), .B(n12360), .ZN(
        n12362) );
  AOI21_X1 U14087 ( .B1(n13635), .B2(n13516), .A(n12362), .ZN(n12368) );
  OAI22_X1 U14088 ( .A1(n12363), .A2(n13486), .B1(n12373), .B2(n13484), .ZN(
        n12364) );
  NAND3_X1 U14089 ( .A1(n12366), .A2(n12365), .A3(n12364), .ZN(n12367) );
  OAI211_X1 U14090 ( .C1(n12369), .C2(n13486), .A(n12368), .B(n12367), .ZN(
        P2_U3200) );
  XNOR2_X1 U14091 ( .A(n12370), .B(n13768), .ZN(n14162) );
  INV_X1 U14092 ( .A(n14162), .ZN(n12381) );
  XNOR2_X1 U14093 ( .A(n12371), .B(n13768), .ZN(n12372) );
  OAI222_X1 U14094 ( .A1(n14057), .A2(n14056), .B1(n14055), .B2(n12373), .C1(
        n12372), .C2(n14063), .ZN(n14160) );
  NAND2_X1 U14095 ( .A1(n14160), .A2(n7197), .ZN(n12380) );
  INV_X1 U14096 ( .A(n14077), .ZN(n12374) );
  AOI211_X1 U14097 ( .C1(n13635), .C2(n12389), .A(n14076), .B(n12374), .ZN(
        n14161) );
  INV_X1 U14098 ( .A(n13635), .ZN(n14220) );
  NOR2_X1 U14099 ( .A1(n14220), .A2(n15821), .ZN(n12378) );
  OAI22_X1 U14100 ( .A1(n7197), .A2(n12376), .B1(n12375), .B2(n13959), .ZN(
        n12377) );
  AOI211_X1 U14101 ( .C1(n14161), .C2(n15814), .A(n12378), .B(n12377), .ZN(
        n12379) );
  OAI211_X1 U14102 ( .C1(n12381), .C2(n14085), .A(n12380), .B(n12379), .ZN(
        P2_U3248) );
  NAND2_X1 U14103 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  NAND2_X1 U14104 ( .A1(n12385), .A2(n12384), .ZN(n14166) );
  INV_X1 U14105 ( .A(n12386), .ZN(n12387) );
  AOI21_X1 U14106 ( .B1(n13626), .B2(n12387), .A(n14076), .ZN(n12388) );
  NAND2_X1 U14107 ( .A1(n12389), .A2(n12388), .ZN(n14167) );
  OR2_X1 U14108 ( .A1(n14166), .A2(n10707), .ZN(n12394) );
  AOI22_X1 U14109 ( .A1(n14070), .A2(n14071), .B1(n14069), .B2(n13801), .ZN(
        n12393) );
  XNOR2_X1 U14110 ( .A(n12390), .B(n13767), .ZN(n12391) );
  NAND2_X1 U14111 ( .A1(n12391), .A2(n14074), .ZN(n12392) );
  OAI21_X1 U14112 ( .B1(n15194), .B2(n14167), .A(n14172), .ZN(n12395) );
  NAND2_X1 U14113 ( .A1(n12395), .A2(n7197), .ZN(n12399) );
  OAI22_X1 U14114 ( .A1(n7197), .A2(n11973), .B1(n12396), .B2(n13959), .ZN(
        n12397) );
  AOI21_X1 U14115 ( .B1(n13626), .B2(n14035), .A(n12397), .ZN(n12398) );
  OAI211_X1 U14116 ( .C1(n14166), .C2(n14066), .A(n12399), .B(n12398), .ZN(
        P2_U3249) );
  AOI22_X1 U14117 ( .A1(n12400), .A2(n12410), .B1(n15843), .B2(n12409), .ZN(
        n12428) );
  NAND2_X1 U14118 ( .A1(n12429), .A2(n7260), .ZN(n12401) );
  NOR2_X2 U14119 ( .A1(n12401), .A2(n12412), .ZN(n12449) );
  AOI21_X1 U14120 ( .B1(n12412), .B2(n12401), .A(n12449), .ZN(n15873) );
  NAND2_X1 U14121 ( .A1(n12435), .A2(n12421), .ZN(n12402) );
  NAND3_X1 U14122 ( .A1(n14764), .A2(n15917), .A3(n12402), .ZN(n15877) );
  INV_X1 U14123 ( .A(n15877), .ZN(n12417) );
  INV_X1 U14124 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U14125 ( .A1(n12435), .A2(n15931), .ZN(n12406) );
  AOI22_X1 U14126 ( .A1(n14362), .A2(n14767), .B1(n14765), .B2(n14361), .ZN(
        n15876) );
  NAND2_X1 U14127 ( .A1(n15930), .A2(n14351), .ZN(n12403) );
  NAND2_X1 U14128 ( .A1(n15876), .A2(n12403), .ZN(n12404) );
  NAND2_X1 U14129 ( .A1(n12404), .A2(n14772), .ZN(n12405) );
  OAI211_X1 U14130 ( .C1(n12407), .C2(n14772), .A(n12406), .B(n12405), .ZN(
        n12416) );
  INV_X1 U14131 ( .A(n12412), .ZN(n12413) );
  AND2_X1 U14132 ( .A1(n12414), .A2(n12413), .ZN(n15874) );
  NOR3_X1 U14133 ( .A1(n15875), .A2(n15874), .A3(n14779), .ZN(n12415) );
  AOI211_X1 U14134 ( .C1(n12417), .C2(n15935), .A(n12416), .B(n12415), .ZN(
        n12418) );
  OAI21_X1 U14135 ( .B1(n15873), .B2(n14740), .A(n12418), .ZN(P1_U3278) );
  XNOR2_X1 U14136 ( .A(n12419), .B(n12427), .ZN(n15856) );
  INV_X1 U14137 ( .A(n14779), .ZN(n12432) );
  AOI21_X1 U14138 ( .B1(n12420), .B2(n12606), .A(n14763), .ZN(n12422) );
  NAND2_X1 U14139 ( .A1(n12422), .A2(n12421), .ZN(n15849) );
  AOI22_X1 U14140 ( .A1(n14363), .A2(n14767), .B1(n14765), .B2(n14768), .ZN(
        n15848) );
  NAND2_X1 U14141 ( .A1(n15930), .A2(n14261), .ZN(n12424) );
  NAND2_X1 U14142 ( .A1(n15941), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12423) );
  OAI211_X1 U14143 ( .C1(n15848), .C2(n15941), .A(n12424), .B(n12423), .ZN(
        n12425) );
  AOI21_X1 U14144 ( .B1(n12606), .B2(n15931), .A(n12425), .ZN(n12426) );
  OAI21_X1 U14145 ( .B1(n15849), .B2(n14672), .A(n12426), .ZN(n12431) );
  NOR2_X1 U14146 ( .A1(n12428), .A2(n12427), .ZN(n15853) );
  INV_X1 U14147 ( .A(n12429), .ZN(n15852) );
  NOR3_X1 U14148 ( .A1(n15853), .A2(n15852), .A3(n14740), .ZN(n12430) );
  AOI211_X1 U14149 ( .C1(n15856), .C2(n12432), .A(n12431), .B(n12430), .ZN(
        n12433) );
  INV_X1 U14150 ( .A(n12433), .ZN(P1_U3279) );
  INV_X1 U14151 ( .A(n13705), .ZN(n14879) );
  INV_X1 U14152 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12434) );
  OAI222_X1 U14153 ( .A1(n14239), .A2(n14879), .B1(P2_U3088), .B2(n8254), .C1(
        n12434), .C2(n14244), .ZN(P2_U3297) );
  AOI21_X1 U14154 ( .B1(n15878), .B2(n14768), .A(n15875), .ZN(n14759) );
  NAND2_X1 U14155 ( .A1(n14759), .A2(n14761), .ZN(n14758) );
  INV_X1 U14156 ( .A(n14766), .ZN(n15944) );
  INV_X1 U14157 ( .A(n14748), .ZN(n14742) );
  NAND2_X1 U14158 ( .A1(n14712), .A2(n14714), .ZN(n14711) );
  INV_X1 U14159 ( .A(n14730), .ZN(n12454) );
  NAND2_X1 U14160 ( .A1(n12438), .A2(n14360), .ZN(n12439) );
  INV_X1 U14161 ( .A(n14658), .ZN(n12441) );
  AOI22_X1 U14162 ( .A1(n14642), .A2(n7960), .B1(n14823), .B2(n14663), .ZN(
        n14626) );
  INV_X1 U14163 ( .A(n14817), .ZN(n14638) );
  INV_X1 U14164 ( .A(n12442), .ZN(n12443) );
  INV_X1 U14165 ( .A(n14620), .ZN(n14609) );
  NAND2_X1 U14166 ( .A1(n14355), .A2(n14765), .ZN(n12446) );
  NAND2_X1 U14167 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  INV_X1 U14168 ( .A(n14768), .ZN(n14258) );
  NOR2_X1 U14169 ( .A1(n15920), .A2(n15944), .ZN(n12450) );
  NAND2_X1 U14170 ( .A1(n14749), .A2(n14748), .ZN(n14747) );
  NAND2_X1 U14171 ( .A1(n7877), .A2(n15902), .ZN(n12451) );
  NAND2_X1 U14172 ( .A1(n14747), .A2(n12451), .ZN(n14726) );
  NAND2_X1 U14173 ( .A1(n14726), .A2(n14729), .ZN(n12453) );
  NAND2_X1 U14174 ( .A1(n14737), .A2(n15943), .ZN(n12452) );
  NAND2_X1 U14175 ( .A1(n12453), .A2(n12452), .ZN(n14713) );
  INV_X1 U14176 ( .A(n14848), .ZN(n14721) );
  INV_X1 U14177 ( .A(n14701), .ZN(n12455) );
  NAND2_X1 U14178 ( .A1(n12438), .A2(n14717), .ZN(n14677) );
  INV_X1 U14179 ( .A(n14662), .ZN(n14270) );
  NAND2_X1 U14180 ( .A1(n14692), .A2(n14270), .ZN(n12457) );
  AND2_X1 U14181 ( .A1(n14677), .A2(n12457), .ZN(n12456) );
  NAND2_X1 U14182 ( .A1(n14675), .A2(n12456), .ZN(n14657) );
  INV_X1 U14183 ( .A(n12457), .ZN(n12458) );
  OR2_X1 U14184 ( .A1(n12458), .A2(n14683), .ZN(n14656) );
  NAND2_X1 U14185 ( .A1(n14657), .A2(n12459), .ZN(n12461) );
  INV_X1 U14186 ( .A(n14670), .ZN(n14830) );
  NAND2_X1 U14187 ( .A1(n14830), .A2(n12667), .ZN(n12460) );
  NAND2_X1 U14188 ( .A1(n12461), .A2(n12460), .ZN(n14643) );
  NAND2_X1 U14189 ( .A1(n14823), .A2(n12673), .ZN(n12462) );
  NAND2_X1 U14190 ( .A1(n14621), .A2(n14620), .ZN(n14619) );
  NAND2_X1 U14191 ( .A1(n14810), .A2(n14357), .ZN(n12463) );
  NAND2_X1 U14192 ( .A1(n14804), .A2(n14334), .ZN(n12465) );
  NAND2_X1 U14193 ( .A1(n12466), .A2(n12467), .ZN(n14796) );
  NAND3_X1 U14194 ( .A1(n14797), .A2(n14796), .A3(n15936), .ZN(n12474) );
  NAND2_X1 U14195 ( .A1(n14692), .A2(n14704), .ZN(n14686) );
  INV_X1 U14196 ( .A(n14810), .ZN(n14618) );
  OR2_X2 U14197 ( .A1(n14612), .A2(n14604), .ZN(n14601) );
  NAND2_X1 U14198 ( .A1(n14799), .A2(n14601), .ZN(n12468) );
  NAND2_X1 U14199 ( .A1(n12468), .A2(n15917), .ZN(n12469) );
  NOR2_X1 U14200 ( .A1(n14576), .A2(n12469), .ZN(n14798) );
  NAND2_X1 U14201 ( .A1(n14799), .A2(n15931), .ZN(n12471) );
  AOI22_X1 U14202 ( .A1(n15941), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n12713), 
        .B2(n15930), .ZN(n12470) );
  NAND2_X1 U14203 ( .A1(n12471), .A2(n12470), .ZN(n12472) );
  AOI21_X1 U14204 ( .B1(n14798), .B2(n15935), .A(n12472), .ZN(n12473) );
  OAI211_X1 U14205 ( .C1(n14801), .C2(n15941), .A(n12474), .B(n12473), .ZN(
        P1_U3265) );
  OAI222_X1 U14206 ( .A1(n14244), .A2(n12476), .B1(n14239), .B2(n12475), .C1(
        n8772), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U14207 ( .A(n12477), .ZN(n12478) );
  OAI222_X1 U14208 ( .A1(n14244), .A2(n12479), .B1(n14239), .B2(n12478), .C1(
        n7193), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14209 ( .A1(n13428), .A2(n13810), .ZN(n12480) );
  OAI22_X1 U14210 ( .A1(n13508), .A2(n13486), .B1(n12481), .B2(n12480), .ZN(
        n12484) );
  INV_X1 U14211 ( .A(n12482), .ZN(n12483) );
  NAND2_X1 U14212 ( .A1(n12484), .A2(n12483), .ZN(n12492) );
  OAI21_X1 U14213 ( .B1(n13479), .B2(n12486), .A(n12485), .ZN(n12490) );
  OAI22_X1 U14214 ( .A1(n12488), .A2(n13499), .B1(n13506), .B2(n12487), .ZN(
        n12489) );
  AOI211_X1 U14215 ( .C1(n13439), .C2(n13810), .A(n12490), .B(n12489), .ZN(
        n12491) );
  OAI211_X1 U14216 ( .C1(n11288), .C2(n13486), .A(n12492), .B(n12491), .ZN(
        P2_U3185) );
  INV_X1 U14217 ( .A(n12494), .ZN(n12497) );
  AOI22_X1 U14218 ( .A1(n13438), .A2(n13801), .B1(n13439), .B2(n13803), .ZN(
        n12496) );
  OAI211_X1 U14219 ( .C1(n12497), .C2(n13479), .A(n12496), .B(n12495), .ZN(
        n12503) );
  INV_X1 U14220 ( .A(n12296), .ZN(n12501) );
  AOI22_X1 U14221 ( .A1(n12498), .A2(n13507), .B1(n13428), .B2(n13803), .ZN(
        n12500) );
  NOR3_X1 U14222 ( .A1(n12501), .A2(n12500), .A3(n12499), .ZN(n12502) );
  AOI211_X1 U14223 ( .C1(n15862), .C2(n13516), .A(n12503), .B(n12502), .ZN(
        n12504) );
  OAI21_X1 U14224 ( .B1(n12493), .B2(n13486), .A(n12504), .ZN(P2_U3187) );
  OAI21_X1 U14225 ( .B1(n13479), .B2(n12506), .A(n12505), .ZN(n12509) );
  OAI22_X1 U14226 ( .A1(n12507), .A2(n13499), .B1(n13506), .B2(n15637), .ZN(
        n12508) );
  AOI211_X1 U14227 ( .C1(n13439), .C2(n13814), .A(n12509), .B(n12508), .ZN(
        n12518) );
  NOR2_X1 U14228 ( .A1(n12510), .A2(n13486), .ZN(n12516) );
  NOR3_X1 U14229 ( .A1(n13484), .A2(n12512), .A3(n12511), .ZN(n12515) );
  INV_X1 U14230 ( .A(n12513), .ZN(n12514) );
  OAI21_X1 U14231 ( .B1(n12516), .B2(n12515), .A(n12514), .ZN(n12517) );
  OAI211_X1 U14232 ( .C1(n13486), .C2(n12519), .A(n12518), .B(n12517), .ZN(
        P2_U3202) );
  INV_X1 U14233 ( .A(n15817), .ZN(n12522) );
  NAND2_X1 U14234 ( .A1(n13513), .A2(n12520), .ZN(n12521) );
  NAND2_X1 U14235 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n13869)
         );
  OAI211_X1 U14236 ( .C1(n13479), .C2(n12522), .A(n12521), .B(n13869), .ZN(
        n12528) );
  AOI22_X1 U14237 ( .A1(n12523), .A2(n13507), .B1(n13428), .B2(n13806), .ZN(
        n12525) );
  NOR3_X1 U14238 ( .A1(n12526), .A2(n12525), .A3(n12524), .ZN(n12527) );
  AOI211_X1 U14239 ( .C1(n13600), .C2(n13516), .A(n12528), .B(n12527), .ZN(
        n12529) );
  OAI21_X1 U14240 ( .B1(n12530), .B2(n13486), .A(n12529), .ZN(P2_U3208) );
  XNOR2_X1 U14241 ( .A(n14141), .B(n12728), .ZN(n12539) );
  INV_X1 U14242 ( .A(n12539), .ZN(n12541) );
  NAND2_X1 U14243 ( .A1(n13797), .A2(n14076), .ZN(n12540) );
  XNOR2_X1 U14244 ( .A(n14155), .B(n12728), .ZN(n12536) );
  NAND2_X1 U14245 ( .A1(n13799), .A2(n14076), .ZN(n12537) );
  INV_X1 U14246 ( .A(n12531), .ZN(n12534) );
  INV_X1 U14247 ( .A(n12532), .ZN(n12533) );
  XNOR2_X1 U14248 ( .A(n12536), .B(n12537), .ZN(n13497) );
  NAND2_X1 U14249 ( .A1(n13498), .A2(n13497), .ZN(n13496) );
  XNOR2_X1 U14250 ( .A(n14048), .B(n11109), .ZN(n13430) );
  NAND2_X1 U14251 ( .A1(n14072), .A2(n14076), .ZN(n12538) );
  NOR2_X1 U14252 ( .A1(n13430), .A2(n12538), .ZN(n13427) );
  NAND2_X1 U14253 ( .A1(n13430), .A2(n12538), .ZN(n13431) );
  NAND2_X1 U14254 ( .A1(n13798), .A2(n14076), .ZN(n13474) );
  XNOR2_X1 U14255 ( .A(n12539), .B(n12540), .ZN(n13448) );
  XNOR2_X1 U14256 ( .A(n14010), .B(n12728), .ZN(n12542) );
  NAND2_X1 U14257 ( .A1(n12543), .A2(n12542), .ZN(n12544) );
  XNOR2_X1 U14258 ( .A(n13994), .B(n12728), .ZN(n12545) );
  NAND2_X1 U14259 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  XNOR2_X1 U14260 ( .A(n14200), .B(n11104), .ZN(n13458) );
  NAND2_X1 U14261 ( .A1(n13794), .A2(n14076), .ZN(n12548) );
  NOR2_X1 U14262 ( .A1(n13458), .A2(n12548), .ZN(n12549) );
  AOI21_X1 U14263 ( .B1(n13458), .B2(n12548), .A(n12549), .ZN(n13468) );
  INV_X1 U14264 ( .A(n12549), .ZN(n12550) );
  NAND2_X1 U14265 ( .A1(n13455), .A2(n12550), .ZN(n12555) );
  XNOR2_X1 U14266 ( .A(n14195), .B(n11109), .ZN(n12551) );
  NOR2_X1 U14267 ( .A1(n13664), .A2(n13976), .ZN(n12552) );
  NAND2_X1 U14268 ( .A1(n12551), .A2(n12552), .ZN(n12556) );
  INV_X1 U14269 ( .A(n12551), .ZN(n12560) );
  INV_X1 U14270 ( .A(n12552), .ZN(n12553) );
  NAND2_X1 U14271 ( .A1(n12560), .A2(n12553), .ZN(n12554) );
  NAND2_X1 U14272 ( .A1(n12555), .A2(n13456), .ZN(n12559) );
  XNOR2_X1 U14273 ( .A(n13944), .B(n11109), .ZN(n12721) );
  NAND2_X1 U14274 ( .A1(n13792), .A2(n14076), .ZN(n12720) );
  XNOR2_X1 U14275 ( .A(n12721), .B(n12720), .ZN(n12561) );
  INV_X1 U14276 ( .A(n12556), .ZN(n12557) );
  NOR2_X1 U14277 ( .A1(n12561), .A2(n12557), .ZN(n12558) );
  NOR2_X1 U14278 ( .A1(n12559), .A2(n13486), .ZN(n12563) );
  NOR3_X1 U14279 ( .A1(n12560), .A2(n13664), .A3(n13484), .ZN(n12562) );
  OAI21_X1 U14280 ( .B1(n12563), .B2(n12562), .A(n12561), .ZN(n12570) );
  OR2_X1 U14281 ( .A1(n13693), .A2(n14057), .ZN(n12565) );
  INV_X1 U14282 ( .A(n13664), .ZN(n13793) );
  NAND2_X1 U14283 ( .A1(n13793), .A2(n14069), .ZN(n12564) );
  NAND2_X1 U14284 ( .A1(n12565), .A2(n12564), .ZN(n13936) );
  OAI22_X1 U14285 ( .A1(n13942), .A2(n13479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12566), .ZN(n12568) );
  NOR2_X1 U14286 ( .A1(n14191), .A2(n13506), .ZN(n12567) );
  AOI211_X1 U14287 ( .C1(n13513), .C2(n13936), .A(n12568), .B(n12567), .ZN(
        n12569) );
  OAI211_X1 U14288 ( .C1(n13486), .C2(n12723), .A(n12570), .B(n12569), .ZN(
        P2_U3212) );
  NAND2_X1 U14289 ( .A1(n13515), .A2(n12571), .ZN(n12573) );
  OAI211_X1 U14290 ( .C1(n13492), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12580) );
  AOI22_X1 U14291 ( .A1(n13428), .A2(n13807), .B1(n12576), .B2(n13507), .ZN(
        n12578) );
  NOR3_X1 U14292 ( .A1(n11837), .A2(n12578), .A3(n12577), .ZN(n12579) );
  AOI211_X1 U14293 ( .C1(n13591), .C2(n13516), .A(n12580), .B(n12579), .ZN(
        n12581) );
  OAI21_X1 U14294 ( .B1(n12582), .B2(n13486), .A(n12581), .ZN(P2_U3189) );
  NOR2_X1 U14295 ( .A1(n13506), .A2(n12583), .ZN(n12587) );
  OAI22_X1 U14296 ( .A1(n13492), .A2(n12585), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12584), .ZN(n12586) );
  AOI211_X1 U14297 ( .C1(n13515), .C2(n12588), .A(n12587), .B(n12586), .ZN(
        n12594) );
  AOI22_X1 U14298 ( .A1(n13428), .A2(n13808), .B1(n13507), .B2(n12589), .ZN(
        n12591) );
  OR3_X1 U14299 ( .A1(n12592), .A2(n12591), .A3(n12590), .ZN(n12593) );
  OAI211_X1 U14300 ( .C1(n12575), .C2(n13486), .A(n12594), .B(n12593), .ZN(
        P2_U3203) );
  INV_X1 U14301 ( .A(n12597), .ZN(n12599) );
  OR2_X1 U14302 ( .A1(n12599), .A2(n12598), .ZN(n12600) );
  NAND2_X1 U14303 ( .A1(n12606), .A2(n10994), .ZN(n12602) );
  NAND2_X1 U14304 ( .A1(n14362), .A2(n7192), .ZN(n12601) );
  NAND2_X1 U14305 ( .A1(n12602), .A2(n12601), .ZN(n12603) );
  XNOR2_X1 U14306 ( .A(n12603), .B(n11198), .ZN(n12608) );
  NOR2_X1 U14307 ( .A1(n12604), .A2(n12706), .ZN(n12605) );
  AOI21_X1 U14308 ( .B1(n12606), .B2(n7192), .A(n12605), .ZN(n12607) );
  NAND2_X1 U14309 ( .A1(n12608), .A2(n12607), .ZN(n12609) );
  OAI21_X1 U14310 ( .B1(n12608), .B2(n12607), .A(n12609), .ZN(n14255) );
  OAI22_X1 U14311 ( .A1(n15878), .A2(n12708), .B1(n14258), .B2(n12640), .ZN(
        n12610) );
  XOR2_X1 U14312 ( .A(n11634), .B(n12610), .Z(n12613) );
  INV_X1 U14313 ( .A(n12613), .ZN(n12611) );
  OAI22_X1 U14314 ( .A1(n15878), .A2(n12640), .B1(n14258), .B2(n12706), .ZN(
        n14344) );
  INV_X1 U14315 ( .A(n14344), .ZN(n12615) );
  OAI22_X1 U14316 ( .A1(n14775), .A2(n12640), .B1(n15904), .B2(n12706), .ZN(
        n12619) );
  OAI22_X1 U14317 ( .A1(n14775), .A2(n12708), .B1(n15904), .B2(n12640), .ZN(
        n12617) );
  XNOR2_X1 U14318 ( .A(n12617), .B(n11634), .ZN(n12618) );
  XOR2_X1 U14319 ( .A(n12619), .B(n12618), .Z(n14295) );
  INV_X1 U14320 ( .A(n12618), .ZN(n12621) );
  INV_X1 U14321 ( .A(n12619), .ZN(n12620) );
  NAND2_X1 U14322 ( .A1(n12621), .A2(n12620), .ZN(n12622) );
  NAND2_X1 U14323 ( .A1(n15932), .A2(n10994), .ZN(n12624) );
  NAND2_X1 U14324 ( .A1(n14766), .A2(n7192), .ZN(n12623) );
  NAND2_X1 U14325 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  XNOR2_X1 U14326 ( .A(n12625), .B(n11634), .ZN(n12628) );
  NAND2_X1 U14327 ( .A1(n15932), .A2(n7192), .ZN(n12627) );
  NAND2_X1 U14328 ( .A1(n14766), .A2(n11435), .ZN(n12626) );
  NAND2_X1 U14329 ( .A1(n12627), .A2(n12626), .ZN(n12629) );
  NAND2_X1 U14330 ( .A1(n12628), .A2(n12629), .ZN(n15897) );
  INV_X1 U14331 ( .A(n12628), .ZN(n12631) );
  INV_X1 U14332 ( .A(n12629), .ZN(n12630) );
  NAND2_X1 U14333 ( .A1(n12631), .A2(n12630), .ZN(n15898) );
  NAND2_X1 U14334 ( .A1(n15953), .A2(n10994), .ZN(n12633) );
  NAND2_X1 U14335 ( .A1(n7876), .A2(n7192), .ZN(n12632) );
  NAND2_X1 U14336 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  XNOR2_X1 U14337 ( .A(n12634), .B(n11634), .ZN(n12635) );
  AOI22_X1 U14338 ( .A1(n15953), .A2(n7192), .B1(n11435), .B2(n7876), .ZN(
        n12636) );
  XNOR2_X1 U14339 ( .A(n12635), .B(n12636), .ZN(n15948) );
  NAND2_X1 U14340 ( .A1(n15946), .A2(n15948), .ZN(n12639) );
  INV_X1 U14341 ( .A(n12635), .ZN(n12637) );
  NAND2_X1 U14342 ( .A1(n12637), .A2(n12636), .ZN(n12638) );
  NAND2_X1 U14343 ( .A1(n12639), .A2(n12638), .ZN(n15957) );
  OAI22_X1 U14344 ( .A1(n14737), .A2(n12640), .B1(n15943), .B2(n12706), .ZN(
        n12644) );
  NAND2_X1 U14345 ( .A1(n15964), .A2(n10994), .ZN(n12642) );
  NAND2_X1 U14346 ( .A1(n14744), .A2(n7192), .ZN(n12641) );
  NAND2_X1 U14347 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  XNOR2_X1 U14348 ( .A(n12643), .B(n11634), .ZN(n12645) );
  XOR2_X1 U14349 ( .A(n12644), .B(n12645), .Z(n15958) );
  NOR2_X1 U14350 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  AOI21_X2 U14351 ( .B1(n15957), .B2(n15958), .A(n12646), .ZN(n14314) );
  NAND2_X1 U14352 ( .A1(n14848), .A2(n10994), .ZN(n12648) );
  NAND2_X1 U14353 ( .A1(n14730), .A2(n7192), .ZN(n12647) );
  NAND2_X1 U14354 ( .A1(n12648), .A2(n12647), .ZN(n12649) );
  XNOR2_X1 U14355 ( .A(n12649), .B(n11634), .ZN(n12653) );
  AND2_X1 U14356 ( .A1(n14730), .A2(n11435), .ZN(n12650) );
  AOI21_X1 U14357 ( .B1(n14848), .B2(n7192), .A(n12650), .ZN(n12651) );
  XNOR2_X1 U14358 ( .A(n12653), .B(n12651), .ZN(n14313) );
  INV_X1 U14359 ( .A(n12651), .ZN(n12652) );
  NAND2_X1 U14360 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  OAI22_X1 U14361 ( .A1(n12438), .A2(n12708), .B1(n14717), .B2(n12640), .ZN(
        n12655) );
  XNOR2_X1 U14362 ( .A(n12655), .B(n11634), .ZN(n12657) );
  OAI22_X1 U14363 ( .A1(n12438), .A2(n12640), .B1(n14717), .B2(n12706), .ZN(
        n12656) );
  XNOR2_X1 U14364 ( .A(n12657), .B(n12656), .ZN(n14277) );
  OAI22_X1 U14365 ( .A1(n14692), .A2(n12708), .B1(n14270), .B2(n12640), .ZN(
        n12659) );
  XNOR2_X1 U14366 ( .A(n12659), .B(n11634), .ZN(n12660) );
  OAI22_X1 U14367 ( .A1(n14692), .A2(n12640), .B1(n14270), .B2(n12706), .ZN(
        n12661) );
  XNOR2_X1 U14368 ( .A(n12660), .B(n12661), .ZN(n14321) );
  INV_X1 U14369 ( .A(n12660), .ZN(n12663) );
  INV_X1 U14370 ( .A(n12661), .ZN(n12662) );
  NAND2_X1 U14371 ( .A1(n14670), .A2(n10994), .ZN(n12665) );
  NAND2_X1 U14372 ( .A1(n14359), .A2(n7192), .ZN(n12664) );
  NAND2_X1 U14373 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  XNOR2_X1 U14374 ( .A(n12666), .B(n11634), .ZN(n12668) );
  OAI22_X1 U14375 ( .A1(n14830), .A2(n12640), .B1(n12667), .B2(n12706), .ZN(
        n12669) );
  XNOR2_X1 U14376 ( .A(n12668), .B(n12669), .ZN(n14267) );
  INV_X1 U14377 ( .A(n12668), .ZN(n12671) );
  INV_X1 U14378 ( .A(n12669), .ZN(n12670) );
  NAND2_X1 U14379 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U14380 ( .A1(n14264), .A2(n12672), .ZN(n14303) );
  OAI22_X1 U14381 ( .A1(n14823), .A2(n12640), .B1(n12673), .B2(n12706), .ZN(
        n12678) );
  NAND2_X1 U14382 ( .A1(n14651), .A2(n10994), .ZN(n12675) );
  NAND2_X1 U14383 ( .A1(n14663), .A2(n7192), .ZN(n12674) );
  NAND2_X1 U14384 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  XNOR2_X1 U14385 ( .A(n12676), .B(n11634), .ZN(n12677) );
  XOR2_X1 U14386 ( .A(n12678), .B(n12677), .Z(n14304) );
  INV_X1 U14387 ( .A(n12677), .ZN(n12680) );
  INV_X1 U14388 ( .A(n12678), .ZN(n12679) );
  NAND2_X1 U14389 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  NAND2_X1 U14390 ( .A1(n14817), .A2(n10994), .ZN(n12683) );
  NAND2_X1 U14391 ( .A1(n14358), .A2(n7192), .ZN(n12682) );
  NAND2_X1 U14392 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  XNOR2_X1 U14393 ( .A(n12684), .B(n11634), .ZN(n12685) );
  AOI22_X1 U14394 ( .A1(n14817), .A2(n7192), .B1(n11435), .B2(n14358), .ZN(
        n12686) );
  XNOR2_X1 U14395 ( .A(n12685), .B(n12686), .ZN(n14285) );
  INV_X1 U14396 ( .A(n12685), .ZN(n12687) );
  NAND2_X1 U14397 ( .A1(n14810), .A2(n10994), .ZN(n12689) );
  NAND2_X1 U14398 ( .A1(n14357), .A2(n7192), .ZN(n12688) );
  NAND2_X1 U14399 ( .A1(n12689), .A2(n12688), .ZN(n12690) );
  XNOR2_X1 U14400 ( .A(n12690), .B(n11634), .ZN(n12694) );
  NAND2_X1 U14401 ( .A1(n14810), .A2(n7192), .ZN(n12693) );
  NAND2_X1 U14402 ( .A1(n14357), .A2(n11435), .ZN(n12692) );
  NAND2_X1 U14403 ( .A1(n12693), .A2(n12692), .ZN(n12695) );
  NAND2_X1 U14404 ( .A1(n12694), .A2(n12695), .ZN(n14331) );
  INV_X1 U14405 ( .A(n12694), .ZN(n12697) );
  INV_X1 U14406 ( .A(n12695), .ZN(n12696) );
  NAND2_X1 U14407 ( .A1(n12697), .A2(n12696), .ZN(n14332) );
  NAND2_X1 U14408 ( .A1(n14604), .A2(n10994), .ZN(n12699) );
  NAND2_X1 U14409 ( .A1(n14356), .A2(n7192), .ZN(n12698) );
  NAND2_X1 U14410 ( .A1(n12699), .A2(n12698), .ZN(n12700) );
  XNOR2_X1 U14411 ( .A(n12700), .B(n11634), .ZN(n12704) );
  NAND2_X1 U14412 ( .A1(n14604), .A2(n7192), .ZN(n12702) );
  NAND2_X1 U14413 ( .A1(n14356), .A2(n11435), .ZN(n12701) );
  NAND2_X1 U14414 ( .A1(n12702), .A2(n12701), .ZN(n12703) );
  NOR2_X1 U14415 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  AOI21_X1 U14416 ( .B1(n12704), .B2(n12703), .A(n12705), .ZN(n14248) );
  OAI22_X1 U14417 ( .A1(n7554), .A2(n12640), .B1(n14568), .B2(n12706), .ZN(
        n12707) );
  XNOR2_X1 U14418 ( .A(n12707), .B(n11634), .ZN(n12710) );
  OAI22_X1 U14419 ( .A1(n7554), .A2(n12708), .B1(n14568), .B2(n12640), .ZN(
        n12709) );
  XNOR2_X1 U14420 ( .A(n12710), .B(n12709), .ZN(n12711) );
  XNOR2_X1 U14421 ( .A(n12712), .B(n12711), .ZN(n12719) );
  AOI22_X1 U14422 ( .A1(n14345), .A2(n14356), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12715) );
  NAND2_X1 U14423 ( .A1(n14352), .A2(n12713), .ZN(n12714) );
  OAI211_X1 U14424 ( .C1(n12716), .C2(n15942), .A(n12715), .B(n12714), .ZN(
        n12717) );
  AOI21_X1 U14425 ( .B1(n14799), .B2(n15965), .A(n12717), .ZN(n12718) );
  OAI21_X1 U14426 ( .B1(n12719), .B2(n15949), .A(n12718), .ZN(P1_U3220) );
  NAND2_X1 U14427 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  XNOR2_X1 U14428 ( .A(n14187), .B(n11109), .ZN(n12725) );
  NOR2_X1 U14429 ( .A1(n13693), .A2(n13976), .ZN(n12724) );
  NAND2_X1 U14430 ( .A1(n12725), .A2(n12724), .ZN(n12727) );
  OAI21_X1 U14431 ( .B1(n12725), .B2(n12724), .A(n12727), .ZN(n13408) );
  NOR2_X1 U14432 ( .A1(n13690), .A2(n13976), .ZN(n12729) );
  XNOR2_X1 U14433 ( .A(n12729), .B(n12728), .ZN(n12730) );
  OR2_X1 U14434 ( .A1(n13693), .A2(n14055), .ZN(n12732) );
  OAI21_X1 U14435 ( .B1(n13689), .B2(n14057), .A(n12732), .ZN(n13904) );
  OAI22_X1 U14436 ( .A1(n13897), .A2(n13479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12733), .ZN(n12735) );
  NOR2_X1 U14437 ( .A1(n14183), .A2(n13506), .ZN(n12734) );
  AOI211_X1 U14438 ( .C1(n13513), .C2(n13904), .A(n12735), .B(n12734), .ZN(
        n12736) );
  OAI21_X1 U14439 ( .B1(n12737), .B2(n13486), .A(n12736), .ZN(P2_U3192) );
  XNOR2_X1 U14440 ( .A(n13326), .B(n12802), .ZN(n12799) );
  XNOR2_X1 U14441 ( .A(n12799), .B(n12905), .ZN(n12800) );
  XNOR2_X1 U14442 ( .A(n12738), .B(n12802), .ZN(n12739) );
  NAND2_X1 U14443 ( .A1(n12739), .A2(n12913), .ZN(n12740) );
  XNOR2_X1 U14444 ( .A(n13390), .B(n12802), .ZN(n12742) );
  XNOR2_X1 U14445 ( .A(n12742), .B(n12912), .ZN(n12777) );
  INV_X1 U14446 ( .A(n12742), .ZN(n12743) );
  XNOR2_X1 U14447 ( .A(n13247), .B(n7205), .ZN(n12825) );
  XNOR2_X1 U14448 ( .A(n13386), .B(n12802), .ZN(n12893) );
  AOI22_X1 U14449 ( .A1(n12825), .A2(n13225), .B1(n12911), .B2(n12893), .ZN(
        n12744) );
  NAND2_X1 U14450 ( .A1(n12826), .A2(n12744), .ZN(n12749) );
  INV_X1 U14451 ( .A(n12825), .ZN(n12837) );
  OAI21_X1 U14452 ( .B1(n12893), .B2(n12911), .A(n13225), .ZN(n12747) );
  INV_X1 U14453 ( .A(n12893), .ZN(n12746) );
  AND2_X1 U14454 ( .A1(n13241), .A2(n12838), .ZN(n12745) );
  AOI22_X1 U14455 ( .A1(n12837), .A2(n12747), .B1(n12746), .B2(n12745), .ZN(
        n12748) );
  NAND2_X1 U14456 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  XNOR2_X1 U14457 ( .A(n13378), .B(n12802), .ZN(n12751) );
  XNOR2_X1 U14458 ( .A(n12751), .B(n13242), .ZN(n12836) );
  INV_X1 U14459 ( .A(n12751), .ZN(n12752) );
  NAND2_X1 U14460 ( .A1(n12752), .A2(n13242), .ZN(n12753) );
  XNOR2_X1 U14461 ( .A(n12878), .B(n12802), .ZN(n12754) );
  XNOR2_X1 U14462 ( .A(n12754), .B(n13224), .ZN(n12875) );
  XNOR2_X1 U14463 ( .A(n13369), .B(n12802), .ZN(n12755) );
  XNOR2_X1 U14464 ( .A(n12755), .B(n13186), .ZN(n12791) );
  NAND2_X1 U14465 ( .A1(n12792), .A2(n12791), .ZN(n12757) );
  NAND2_X1 U14466 ( .A1(n12755), .A2(n13213), .ZN(n12756) );
  XNOR2_X1 U14467 ( .A(n13362), .B(n7205), .ZN(n12758) );
  NAND2_X1 U14468 ( .A1(n12758), .A2(n13172), .ZN(n12858) );
  NAND2_X1 U14469 ( .A1(n12861), .A2(n12858), .ZN(n12760) );
  INV_X1 U14470 ( .A(n12758), .ZN(n12759) );
  NAND2_X1 U14471 ( .A1(n12759), .A2(n13199), .ZN(n12859) );
  NAND2_X1 U14472 ( .A1(n12760), .A2(n12859), .ZN(n12812) );
  XNOR2_X1 U14473 ( .A(n13178), .B(n12802), .ZN(n12810) );
  OAI21_X1 U14474 ( .B1(n12812), .B2(n13157), .A(n12810), .ZN(n12762) );
  NAND2_X1 U14475 ( .A1(n12812), .A2(n13157), .ZN(n12761) );
  XNOR2_X1 U14476 ( .A(n13351), .B(n7205), .ZN(n12763) );
  INV_X1 U14477 ( .A(n12763), .ZN(n12764) );
  XNOR2_X1 U14478 ( .A(n13276), .B(n12802), .ZN(n12849) );
  XNOR2_X1 U14479 ( .A(n13147), .B(n12802), .ZN(n12766) );
  OAI22_X1 U14480 ( .A1(n12849), .A2(n13138), .B1(n13158), .B2(n12766), .ZN(
        n12768) );
  INV_X1 U14481 ( .A(n12766), .ZN(n12846) );
  OAI21_X1 U14482 ( .B1(n12846), .B2(n12909), .A(n12908), .ZN(n12767) );
  XNOR2_X1 U14483 ( .A(n13339), .B(n12802), .ZN(n12769) );
  XNOR2_X1 U14484 ( .A(n12769), .B(n12907), .ZN(n12819) );
  XNOR2_X1 U14485 ( .A(n13333), .B(n7191), .ZN(n12770) );
  XNOR2_X1 U14486 ( .A(n12770), .B(n13106), .ZN(n12884) );
  INV_X1 U14487 ( .A(n12770), .ZN(n12771) );
  XOR2_X1 U14488 ( .A(n12800), .B(n12801), .Z(n12776) );
  OAI22_X1 U14489 ( .A1(n13077), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15083), .ZN(n12772) );
  AOI21_X1 U14490 ( .B1(n13085), .B2(n12900), .A(n12772), .ZN(n12773) );
  OAI21_X1 U14491 ( .B1(n13106), .B2(n12897), .A(n12773), .ZN(n12774) );
  AOI21_X1 U14492 ( .B1(n13326), .B2(n12887), .A(n12774), .ZN(n12775) );
  OAI21_X1 U14493 ( .B1(n12776), .B2(n12890), .A(n12775), .ZN(P3_U3154) );
  XOR2_X1 U14494 ( .A(n12778), .B(n12777), .Z(n12785) );
  NAND2_X1 U14495 ( .A1(n12895), .A2(n12911), .ZN(n12779) );
  NAND2_X1 U14496 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15480)
         );
  OAI211_X1 U14497 ( .C1(n12780), .C2(n12897), .A(n12779), .B(n15480), .ZN(
        n12782) );
  NOR2_X1 U14498 ( .A1(n13390), .A2(n15128), .ZN(n12781) );
  AOI211_X1 U14499 ( .C1(n12783), .C2(n12900), .A(n12782), .B(n12781), .ZN(
        n12784) );
  OAI21_X1 U14500 ( .B1(n12785), .B2(n12890), .A(n12784), .ZN(P3_U3155) );
  INV_X1 U14501 ( .A(n13147), .ZN(n13348) );
  XNOR2_X1 U14502 ( .A(n12847), .B(n12846), .ZN(n12848) );
  XNOR2_X1 U14503 ( .A(n12848), .B(n12909), .ZN(n12786) );
  NAND2_X1 U14504 ( .A1(n12786), .A2(n15131), .ZN(n12790) );
  OAI22_X1 U14505 ( .A1(n13137), .A2(n12897), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15015), .ZN(n12788) );
  NOR2_X1 U14506 ( .A1(n13138), .A2(n15126), .ZN(n12787) );
  AOI211_X1 U14507 ( .C1(n13142), .C2(n12900), .A(n12788), .B(n12787), .ZN(
        n12789) );
  OAI211_X1 U14508 ( .C1(n13348), .C2(n15128), .A(n12790), .B(n12789), .ZN(
        P3_U3156) );
  XNOR2_X1 U14509 ( .A(n12792), .B(n12791), .ZN(n12793) );
  NAND2_X1 U14510 ( .A1(n12793), .A2(n15131), .ZN(n12798) );
  NOR2_X1 U14511 ( .A1(n13198), .A2(n12897), .ZN(n12796) );
  INV_X1 U14512 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12794) );
  OAI22_X1 U14513 ( .A1(n13199), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12794), .ZN(n12795) );
  AOI211_X1 U14514 ( .C1(n12900), .C2(n13204), .A(n12796), .B(n12795), .ZN(
        n12797) );
  OAI211_X1 U14515 ( .C1(n13206), .C2(n15128), .A(n12798), .B(n12797), .ZN(
        P3_U3159) );
  XNOR2_X1 U14516 ( .A(n13068), .B(n12802), .ZN(n12803) );
  XNOR2_X1 U14517 ( .A(n12804), .B(n12803), .ZN(n12805) );
  NOR2_X1 U14518 ( .A1(n13091), .A2(n12897), .ZN(n12808) );
  OAI22_X1 U14519 ( .A1(n13064), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12806), .ZN(n12807) );
  AOI211_X1 U14520 ( .C1(n13070), .C2(n12900), .A(n12808), .B(n12807), .ZN(
        n12809) );
  INV_X1 U14521 ( .A(n13178), .ZN(n13356) );
  XNOR2_X1 U14522 ( .A(n12810), .B(n13187), .ZN(n12811) );
  XNOR2_X1 U14523 ( .A(n12812), .B(n12811), .ZN(n12813) );
  NAND2_X1 U14524 ( .A1(n12813), .A2(n15131), .ZN(n12817) );
  NOR2_X1 U14525 ( .A1(n13199), .A2(n12897), .ZN(n12815) );
  OAI22_X1 U14526 ( .A1(n13137), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15096), .ZN(n12814) );
  AOI211_X1 U14527 ( .C1(n13177), .C2(n12900), .A(n12815), .B(n12814), .ZN(
        n12816) );
  OAI211_X1 U14528 ( .C1(n13356), .C2(n15128), .A(n12817), .B(n12816), .ZN(
        P3_U3163) );
  XOR2_X1 U14529 ( .A(n12819), .B(n12818), .Z(n12824) );
  AOI22_X1 U14530 ( .A1(n12908), .A2(n12876), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12821) );
  NAND2_X1 U14531 ( .A1(n12900), .A2(n13112), .ZN(n12820) );
  OAI211_X1 U14532 ( .C1(n13106), .C2(n15126), .A(n12821), .B(n12820), .ZN(
        n12822) );
  AOI21_X1 U14533 ( .B1(n13339), .B2(n12887), .A(n12822), .ZN(n12823) );
  OAI21_X1 U14534 ( .B1(n12824), .B2(n12890), .A(n12823), .ZN(P3_U3165) );
  XNOR2_X1 U14535 ( .A(n12825), .B(n13225), .ZN(n12828) );
  XNOR2_X1 U14536 ( .A(n12826), .B(n12911), .ZN(n12894) );
  NAND2_X1 U14537 ( .A1(n12894), .A2(n12893), .ZN(n12892) );
  OAI21_X1 U14538 ( .B1(n13241), .B2(n12826), .A(n12892), .ZN(n12827) );
  NOR2_X1 U14539 ( .A1(n12827), .A2(n12828), .ZN(n12835) );
  AOI21_X1 U14540 ( .B1(n12828), .B2(n12827), .A(n12835), .ZN(n12834) );
  NOR2_X1 U14541 ( .A1(n13241), .A2(n12897), .ZN(n12831) );
  OAI22_X1 U14542 ( .A1(n13242), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12829), .ZN(n12830) );
  AOI211_X1 U14543 ( .C1(n12900), .C2(n13248), .A(n12831), .B(n12830), .ZN(
        n12833) );
  NAND2_X1 U14544 ( .A1(n13247), .A2(n12887), .ZN(n12832) );
  OAI211_X1 U14545 ( .C1(n12834), .C2(n12890), .A(n12833), .B(n12832), .ZN(
        P3_U3166) );
  AOI211_X1 U14546 ( .C1(n12838), .C2(n12837), .A(n12836), .B(n12835), .ZN(
        n12841) );
  INV_X1 U14547 ( .A(n12839), .ZN(n12840) );
  OAI21_X1 U14548 ( .B1(n12841), .B2(n12840), .A(n15131), .ZN(n12845) );
  NAND2_X1 U14549 ( .A1(n13225), .A2(n12876), .ZN(n12842) );
  NAND2_X1 U14550 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12992)
         );
  OAI211_X1 U14551 ( .C1(n13198), .C2(n15126), .A(n12842), .B(n12992), .ZN(
        n12843) );
  AOI21_X1 U14552 ( .B1(n12900), .B2(n13231), .A(n12843), .ZN(n12844) );
  OAI211_X1 U14553 ( .C1(n15128), .C2(n13378), .A(n12845), .B(n12844), .ZN(
        P3_U3168) );
  OAI22_X1 U14554 ( .A1(n12848), .A2(n12909), .B1(n12847), .B2(n12846), .ZN(
        n12851) );
  XNOR2_X1 U14555 ( .A(n12849), .B(n13138), .ZN(n12850) );
  XNOR2_X1 U14556 ( .A(n12851), .B(n12850), .ZN(n12857) );
  INV_X1 U14557 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12852) );
  OAI22_X1 U14558 ( .A1(n13158), .A2(n12897), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12852), .ZN(n12854) );
  NOR2_X1 U14559 ( .A1(n13128), .A2(n15126), .ZN(n12853) );
  AOI211_X1 U14560 ( .C1(n13129), .C2(n12900), .A(n12854), .B(n12853), .ZN(
        n12856) );
  NAND2_X1 U14561 ( .A1(n13276), .A2(n12887), .ZN(n12855) );
  OAI211_X1 U14562 ( .C1(n12857), .C2(n12890), .A(n12856), .B(n12855), .ZN(
        P3_U3169) );
  NAND2_X1 U14563 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  XNOR2_X1 U14564 ( .A(n12861), .B(n12860), .ZN(n12866) );
  NOR2_X1 U14565 ( .A1(n13213), .A2(n12897), .ZN(n12863) );
  OAI22_X1 U14566 ( .A1(n13157), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15108), .ZN(n12862) );
  AOI211_X1 U14567 ( .C1(n13192), .C2(n12900), .A(n12863), .B(n12862), .ZN(
        n12865) );
  NAND2_X1 U14568 ( .A1(n13362), .A2(n12887), .ZN(n12864) );
  OAI211_X1 U14569 ( .C1(n12866), .C2(n12890), .A(n12865), .B(n12864), .ZN(
        P3_U3173) );
  XNOR2_X1 U14570 ( .A(n12867), .B(n13173), .ZN(n12873) );
  NOR2_X1 U14571 ( .A1(n13157), .A2(n12897), .ZN(n12870) );
  OAI22_X1 U14572 ( .A1(n13158), .A2(n15126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12868), .ZN(n12869) );
  AOI211_X1 U14573 ( .C1(n13163), .C2(n12900), .A(n12870), .B(n12869), .ZN(
        n12872) );
  NAND2_X1 U14574 ( .A1(n13351), .A2(n12887), .ZN(n12871) );
  OAI211_X1 U14575 ( .C1(n12873), .C2(n12890), .A(n12872), .B(n12871), .ZN(
        P3_U3175) );
  XOR2_X1 U14576 ( .A(n12875), .B(n12874), .Z(n12882) );
  NAND2_X1 U14577 ( .A1(n12876), .A2(n12910), .ZN(n12877) );
  NAND2_X1 U14578 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13010)
         );
  OAI211_X1 U14579 ( .C1(n13213), .C2(n15126), .A(n12877), .B(n13010), .ZN(
        n12880) );
  INV_X1 U14580 ( .A(n12878), .ZN(n13374) );
  NOR2_X1 U14581 ( .A1(n13374), .A2(n15128), .ZN(n12879) );
  AOI211_X1 U14582 ( .C1(n13217), .C2(n12900), .A(n12880), .B(n12879), .ZN(
        n12881) );
  OAI21_X1 U14583 ( .B1(n12882), .B2(n12890), .A(n12881), .ZN(P3_U3178) );
  XOR2_X1 U14584 ( .A(n12884), .B(n12883), .Z(n12891) );
  OAI22_X1 U14585 ( .A1(n13128), .A2(n12897), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15121), .ZN(n12886) );
  NOR2_X1 U14586 ( .A1(n13091), .A2(n15126), .ZN(n12885) );
  AOI211_X1 U14587 ( .C1(n13096), .C2(n12900), .A(n12886), .B(n12885), .ZN(
        n12889) );
  NAND2_X1 U14588 ( .A1(n13333), .A2(n12887), .ZN(n12888) );
  OAI211_X1 U14589 ( .C1(n12891), .C2(n12890), .A(n12889), .B(n12888), .ZN(
        P3_U3180) );
  OAI211_X1 U14590 ( .C1(n12894), .C2(n12893), .A(n12892), .B(n15131), .ZN(
        n12903) );
  INV_X1 U14591 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U14592 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15118), .ZN(n15488) );
  AOI21_X1 U14593 ( .B1(n13225), .B2(n12895), .A(n15488), .ZN(n12896) );
  OAI21_X1 U14594 ( .B1(n12898), .B2(n12897), .A(n12896), .ZN(n12899) );
  AOI21_X1 U14595 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12902) );
  OAI211_X1 U14596 ( .C1(n15128), .C2(n13386), .A(n12903), .B(n12902), .ZN(
        P3_U3181) );
  MUX2_X1 U14597 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12904), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14598 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12905), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14599 ( .A(n12906), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12925), .Z(
        P3_U3517) );
  MUX2_X1 U14600 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12907), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14601 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12908), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14602 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12909), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14603 ( .A(n13173), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12925), .Z(
        P3_U3513) );
  MUX2_X1 U14604 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13187), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14605 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13172), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14606 ( .A(n13186), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12925), .Z(
        P3_U3510) );
  MUX2_X1 U14607 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13224), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14608 ( .A(n12910), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12925), .Z(
        P3_U3508) );
  MUX2_X1 U14609 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13225), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14610 ( .A(n12911), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12925), .Z(
        P3_U3506) );
  MUX2_X1 U14611 ( .A(n12912), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12925), .Z(
        P3_U3505) );
  MUX2_X1 U14612 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12913), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14613 ( .A(n12914), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12925), .Z(
        P3_U3503) );
  MUX2_X1 U14614 ( .A(n12915), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12925), .Z(
        P3_U3502) );
  MUX2_X1 U14615 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12916), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14616 ( .A(n12917), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12925), .Z(
        P3_U3500) );
  MUX2_X1 U14617 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12918), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14618 ( .A(n12919), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12925), .Z(
        P3_U3498) );
  MUX2_X1 U14619 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12920), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14620 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12921), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14621 ( .A(n12922), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12925), .Z(
        P3_U3495) );
  MUX2_X1 U14622 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12923), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14623 ( .A(n15546), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12925), .Z(
        P3_U3493) );
  MUX2_X1 U14624 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12924), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14625 ( .A(n10042), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12925), .Z(
        P3_U3491) );
  INV_X1 U14626 ( .A(n15490), .ZN(n12936) );
  INV_X1 U14627 ( .A(n12970), .ZN(n15468) );
  INV_X1 U14628 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n15467) );
  NAND2_X1 U14629 ( .A1(n15468), .A2(n15467), .ZN(n15466) );
  NAND2_X1 U14630 ( .A1(n15433), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12956) );
  OR2_X1 U14631 ( .A1(n15433), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12926) );
  AND2_X1 U14632 ( .A1(n12956), .A2(n12926), .ZN(n15437) );
  INV_X1 U14633 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U14634 ( .A1(n15405), .A2(n12931), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n12971), .ZN(n15403) );
  NAND2_X1 U14635 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n12972), .ZN(n12928) );
  NAND2_X1 U14636 ( .A1(n12928), .A2(n12927), .ZN(n12929) );
  NAND2_X1 U14637 ( .A1(n12975), .A2(n12929), .ZN(n12930) );
  INV_X1 U14638 ( .A(n12975), .ZN(n15388) );
  XNOR2_X1 U14639 ( .A(n15388), .B(n12929), .ZN(n15391) );
  NAND2_X1 U14640 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n15391), .ZN(n15390) );
  NAND2_X1 U14641 ( .A1(n12978), .A2(n12932), .ZN(n12933) );
  INV_X1 U14642 ( .A(n12978), .ZN(n15419) );
  NAND2_X1 U14643 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n15421), .ZN(n15420) );
  NAND2_X1 U14644 ( .A1(n12933), .A2(n15420), .ZN(n15436) );
  NAND2_X1 U14645 ( .A1(n15437), .A2(n15436), .ZN(n15435) );
  NAND2_X1 U14646 ( .A1(n12956), .A2(n15435), .ZN(n12934) );
  NAND2_X1 U14647 ( .A1(n12982), .A2(n12934), .ZN(n12935) );
  INV_X1 U14648 ( .A(n12982), .ZN(n15450) );
  NOR2_X1 U14649 ( .A1(n12936), .A2(n12937), .ZN(n12938) );
  INV_X1 U14650 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15485) );
  XNOR2_X1 U14651 ( .A(n12937), .B(n12936), .ZN(n15484) );
  NOR2_X1 U14652 ( .A1(n15485), .A2(n15484), .ZN(n15483) );
  NAND2_X1 U14653 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12988), .ZN(n12939) );
  OAI21_X1 U14654 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12988), .A(n12939), 
        .ZN(n15518) );
  INV_X1 U14655 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12940) );
  NOR2_X1 U14656 ( .A1(n12940), .A2(n12941), .ZN(n13000) );
  AOI21_X1 U14657 ( .B1(n12941), .B2(n12940), .A(n13000), .ZN(n12998) );
  MUX2_X1 U14658 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12955), .Z(n12942) );
  AND2_X1 U14659 ( .A1(n12993), .A2(n12942), .ZN(n13005) );
  NOR2_X1 U14660 ( .A1(n12993), .A2(n12942), .ZN(n12943) );
  OR2_X1 U14661 ( .A1(n13005), .A2(n12943), .ZN(n12969) );
  MUX2_X1 U14662 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12955), .Z(n12960) );
  NAND2_X1 U14663 ( .A1(n12960), .A2(n12970), .ZN(n12961) );
  MUX2_X1 U14664 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12955), .Z(n12958) );
  INV_X1 U14665 ( .A(n12958), .ZN(n12959) );
  MUX2_X1 U14666 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12955), .Z(n12952) );
  INV_X1 U14667 ( .A(n12952), .ZN(n12953) );
  MUX2_X1 U14668 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12955), .Z(n12950) );
  INV_X1 U14669 ( .A(n12950), .ZN(n12951) );
  MUX2_X1 U14670 ( .A(n12944), .B(n11923), .S(n12955), .Z(n12945) );
  AND2_X1 U14671 ( .A1(n12945), .A2(n15388), .ZN(n15381) );
  OR2_X1 U14672 ( .A1(n12946), .A2(n12972), .ZN(n12948) );
  NAND2_X1 U14673 ( .A1(n12948), .A2(n12947), .ZN(n15385) );
  MUX2_X1 U14674 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12955), .Z(n12949) );
  NAND2_X1 U14675 ( .A1(n12949), .A2(n12975), .ZN(n15383) );
  XNOR2_X1 U14676 ( .A(n12950), .B(n12971), .ZN(n15400) );
  XNOR2_X1 U14677 ( .A(n12952), .B(n12978), .ZN(n15427) );
  AOI21_X1 U14678 ( .B1(n15419), .B2(n12953), .A(n15426), .ZN(n15445) );
  NAND2_X1 U14679 ( .A1(n15433), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12981) );
  OR2_X1 U14680 ( .A1(n15433), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12954) );
  AND2_X1 U14681 ( .A1(n12981), .A2(n12954), .ZN(n15440) );
  MUX2_X1 U14682 ( .A(n15437), .B(n15440), .S(n12955), .Z(n15444) );
  NAND2_X1 U14683 ( .A1(n15445), .A2(n15444), .ZN(n15443) );
  MUX2_X1 U14684 ( .A(n12956), .B(n12981), .S(n12955), .Z(n12957) );
  NAND2_X1 U14685 ( .A1(n15443), .A2(n12957), .ZN(n15458) );
  XNOR2_X1 U14686 ( .A(n12958), .B(n12982), .ZN(n15459) );
  NOR2_X1 U14687 ( .A1(n15458), .A2(n15459), .ZN(n15457) );
  XNOR2_X1 U14688 ( .A(n12960), .B(n15468), .ZN(n15477) );
  NOR2_X1 U14689 ( .A1(n15490), .A2(n12962), .ZN(n12964) );
  INV_X1 U14690 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13310) );
  MUX2_X1 U14691 ( .A(n15485), .B(n13310), .S(n12955), .Z(n15495) );
  XNOR2_X1 U14692 ( .A(n15490), .B(n12963), .ZN(n15494) );
  AND2_X1 U14693 ( .A1(n15495), .A2(n15494), .ZN(n15497) );
  NOR2_X1 U14694 ( .A1(n12964), .A2(n15497), .ZN(n15507) );
  MUX2_X1 U14695 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12955), .Z(n12965) );
  NAND2_X1 U14696 ( .A1(n12965), .A2(n12988), .ZN(n15504) );
  INV_X1 U14697 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12966) );
  INV_X1 U14698 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n15509) );
  MUX2_X1 U14699 ( .A(n12966), .B(n15509), .S(n12955), .Z(n12967) );
  NAND2_X1 U14700 ( .A1(n12967), .A2(n15510), .ZN(n15505) );
  AOI211_X1 U14701 ( .C1(n12969), .C2(n12968), .A(n15460), .B(n7270), .ZN(
        n12996) );
  INV_X1 U14702 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13303) );
  NAND2_X1 U14703 ( .A1(n15510), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U14704 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n12970), .ZN(n12985) );
  INV_X1 U14705 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14706 ( .A1(n15468), .A2(n13314), .B1(P3_REG1_REG_14__SCAN_IN), 
        .B2(n12970), .ZN(n15473) );
  INV_X1 U14707 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15794) );
  AOI22_X1 U14708 ( .A1(n15405), .A2(n15794), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n12971), .ZN(n15409) );
  NAND2_X1 U14709 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n12972), .ZN(n12974) );
  NAND2_X1 U14710 ( .A1(n12974), .A2(n12973), .ZN(n12976) );
  NAND2_X1 U14711 ( .A1(n12975), .A2(n12976), .ZN(n12977) );
  XNOR2_X1 U14712 ( .A(n15388), .B(n12976), .ZN(n15387) );
  NAND2_X1 U14713 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15387), .ZN(n15386) );
  NAND2_X1 U14714 ( .A1(n12977), .A2(n15386), .ZN(n15408) );
  NAND2_X1 U14715 ( .A1(n15409), .A2(n15408), .ZN(n15407) );
  NAND2_X1 U14716 ( .A1(n12978), .A2(n12979), .ZN(n12980) );
  XNOR2_X1 U14717 ( .A(n15419), .B(n12979), .ZN(n15423) );
  NAND2_X1 U14718 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15423), .ZN(n15422) );
  NAND2_X1 U14719 ( .A1(n12980), .A2(n15422), .ZN(n15439) );
  NAND2_X1 U14720 ( .A1(n15440), .A2(n15439), .ZN(n15438) );
  NAND2_X1 U14721 ( .A1(n12981), .A2(n15438), .ZN(n12983) );
  NAND2_X1 U14722 ( .A1(n12982), .A2(n12983), .ZN(n12984) );
  NAND2_X1 U14723 ( .A1(n12984), .A2(n15453), .ZN(n15472) );
  NAND2_X1 U14724 ( .A1(n15473), .A2(n15472), .ZN(n15471) );
  NAND2_X1 U14725 ( .A1(n15490), .A2(n12986), .ZN(n12987) );
  NAND2_X1 U14726 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n15487), .ZN(n15486) );
  NAND2_X1 U14727 ( .A1(n12987), .A2(n15486), .ZN(n15512) );
  XNOR2_X1 U14728 ( .A(n13013), .B(n13014), .ZN(n12989) );
  NOR2_X1 U14729 ( .A1(n13303), .A2(n12989), .ZN(n13015) );
  AOI21_X1 U14730 ( .B1(n13303), .B2(n12989), .A(n13015), .ZN(n12990) );
  NOR2_X1 U14731 ( .A1(n12990), .A2(n15373), .ZN(n12995) );
  NAND2_X1 U14732 ( .A1(n15502), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12991) );
  OAI211_X1 U14733 ( .C1(n15491), .C2(n12993), .A(n12992), .B(n12991), .ZN(
        n12994) );
  NOR3_X1 U14734 ( .A1(n12996), .A2(n12995), .A3(n12994), .ZN(n12997) );
  OAI21_X1 U14735 ( .B1(n12998), .B2(n15500), .A(n12997), .ZN(P3_U3199) );
  NOR2_X1 U14736 ( .A1(n13014), .A2(n12999), .ZN(n13001) );
  NOR2_X1 U14737 ( .A1(n13001), .A2(n13000), .ZN(n13004) );
  NAND2_X1 U14738 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n13029), .ZN(n13002) );
  OAI21_X1 U14739 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13029), .A(n13002), 
        .ZN(n13003) );
  NOR2_X1 U14740 ( .A1(n13004), .A2(n13003), .ZN(n13024) );
  AOI21_X1 U14741 ( .B1(n13004), .B2(n13003), .A(n13024), .ZN(n13023) );
  INV_X1 U14742 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13012) );
  XNOR2_X1 U14743 ( .A(n13029), .B(n13031), .ZN(n13008) );
  INV_X1 U14744 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13006) );
  INV_X1 U14745 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13299) );
  MUX2_X1 U14746 ( .A(n13006), .B(n13299), .S(n12955), .Z(n13007) );
  NAND2_X1 U14747 ( .A1(n13008), .A2(n13007), .ZN(n13034) );
  OAI21_X1 U14748 ( .B1(n13008), .B2(n13007), .A(n13034), .ZN(n13009) );
  NAND2_X1 U14749 ( .A1(n13009), .A2(n15515), .ZN(n13011) );
  OAI211_X1 U14750 ( .C1(n15417), .C2(n13012), .A(n13011), .B(n13010), .ZN(
        n13021) );
  NOR2_X1 U14751 ( .A1(n13014), .A2(n13013), .ZN(n13016) );
  NOR2_X1 U14752 ( .A1(n13016), .A2(n13015), .ZN(n13018) );
  AOI22_X1 U14753 ( .A1(n13032), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n13299), 
        .B2(n13029), .ZN(n13017) );
  NOR2_X1 U14754 ( .A1(n13019), .A2(n15373), .ZN(n13020) );
  OAI21_X1 U14755 ( .B1(n13023), .B2(n15500), .A(n13022), .ZN(P3_U3200) );
  AOI21_X1 U14756 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13029), .A(n13024), 
        .ZN(n13027) );
  INV_X1 U14757 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13026) );
  MUX2_X1 U14758 ( .A(n13026), .B(P3_REG2_REG_19__SCAN_IN), .S(n7209), .Z(
        n13037) );
  XNOR2_X1 U14759 ( .A(n13027), .B(n13037), .ZN(n13046) );
  AOI21_X1 U14760 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n13029), .A(n13028), 
        .ZN(n13030) );
  XNOR2_X1 U14761 ( .A(n13042), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13035) );
  XNOR2_X1 U14762 ( .A(n13030), .B(n13035), .ZN(n13044) );
  NAND2_X1 U14763 ( .A1(n13032), .A2(n13031), .ZN(n13033) );
  INV_X1 U14764 ( .A(n13035), .ZN(n13038) );
  MUX2_X1 U14765 ( .A(n13038), .B(n13037), .S(n7384), .Z(n13039) );
  NAND2_X1 U14766 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n13041)
         );
  NAND2_X1 U14767 ( .A1(n15502), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13040) );
  OAI211_X1 U14768 ( .C1(n15491), .C2(n13042), .A(n13041), .B(n13040), .ZN(
        n13043) );
  OAI21_X1 U14769 ( .B1(n13046), .B2(n15500), .A(n13045), .ZN(P3_U3201) );
  NAND2_X1 U14770 ( .A1(n13055), .A2(n15680), .ZN(n13049) );
  OR2_X1 U14771 ( .A1(n13048), .A2(n13047), .ZN(n15979) );
  NAND3_X1 U14772 ( .A1(n15688), .A2(n13049), .A3(n15979), .ZN(n13051) );
  OAI21_X1 U14773 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15688), .A(n13051), 
        .ZN(n13050) );
  OAI21_X1 U14774 ( .B1(n13319), .B2(n13250), .A(n13050), .ZN(P3_U3202) );
  OAI21_X1 U14775 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15688), .A(n13051), 
        .ZN(n13052) );
  OAI21_X1 U14776 ( .B1(n13053), .B2(n13250), .A(n13052), .ZN(P3_U3203) );
  INV_X1 U14777 ( .A(n13054), .ZN(n13061) );
  AOI22_X1 U14778 ( .A1(n13055), .A2(n15680), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15690), .ZN(n13056) );
  OAI21_X1 U14779 ( .B1(n13057), .B2(n13250), .A(n13056), .ZN(n13058) );
  AOI21_X1 U14780 ( .B1(n13059), .B2(n13252), .A(n13058), .ZN(n13060) );
  OAI21_X1 U14781 ( .B1(n13061), .B2(n15690), .A(n13060), .ZN(P3_U3204) );
  OAI211_X1 U14782 ( .C1(n13063), .C2(n13068), .A(n13062), .B(n15577), .ZN(
        n13067) );
  OAI22_X1 U14783 ( .A1(n13064), .A2(n13243), .B1(n13091), .B2(n15575), .ZN(
        n13065) );
  INV_X1 U14784 ( .A(n13065), .ZN(n13066) );
  XNOR2_X1 U14785 ( .A(n13069), .B(n13068), .ZN(n13257) );
  AOI22_X1 U14786 ( .A1(n13070), .A2(n15680), .B1(n15690), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13071) );
  OAI21_X1 U14787 ( .B1(n13323), .B2(n13250), .A(n13071), .ZN(n13072) );
  AOI21_X1 U14788 ( .B1(n13257), .B2(n13252), .A(n13072), .ZN(n13073) );
  OAI21_X1 U14789 ( .B1(n13259), .B2(n15690), .A(n13073), .ZN(P3_U3205) );
  OR2_X1 U14790 ( .A1(n13074), .A2(n13080), .ZN(n13075) );
  INV_X1 U14791 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13084) );
  OAI22_X1 U14792 ( .A1(n13077), .A2(n13243), .B1(n13106), .B2(n15575), .ZN(
        n13083) );
  NAND2_X1 U14793 ( .A1(n13079), .A2(n13080), .ZN(n13081) );
  AOI21_X1 U14794 ( .B1(n13078), .B2(n13081), .A(n13240), .ZN(n13082) );
  AOI211_X1 U14795 ( .C1(n13327), .C2(n15632), .A(n13083), .B(n13082), .ZN(
        n13324) );
  MUX2_X1 U14796 ( .A(n13084), .B(n13324), .S(n15688), .Z(n13087) );
  AOI22_X1 U14797 ( .A1(n13326), .A2(n15684), .B1(n15680), .B2(n13085), .ZN(
        n13086) );
  OAI211_X1 U14798 ( .C1(n13265), .C2(n13195), .A(n13087), .B(n13086), .ZN(
        P3_U3206) );
  INV_X1 U14799 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13095) );
  XNOR2_X1 U14800 ( .A(n13090), .B(n13089), .ZN(n13094) );
  NOR2_X1 U14801 ( .A1(n13336), .A2(n15733), .ZN(n13093) );
  OAI22_X1 U14802 ( .A1(n13091), .A2(n13243), .B1(n13128), .B2(n15575), .ZN(
        n13092) );
  MUX2_X1 U14803 ( .A(n13095), .B(n13331), .S(n15688), .Z(n13098) );
  AOI22_X1 U14804 ( .A1(n13333), .A2(n15684), .B1(n13096), .B2(n15680), .ZN(
        n13097) );
  OAI211_X1 U14805 ( .C1(n13336), .C2(n13195), .A(n13098), .B(n13097), .ZN(
        P3_U3207) );
  OR2_X1 U14806 ( .A1(n13099), .A2(n13100), .ZN(n13102) );
  NAND2_X1 U14807 ( .A1(n13102), .A2(n13101), .ZN(n13105) );
  INV_X1 U14808 ( .A(n13103), .ZN(n13111) );
  OAI211_X1 U14809 ( .C1(n13105), .C2(n13111), .A(n13104), .B(n15577), .ZN(
        n13109) );
  OAI22_X1 U14810 ( .A1(n13106), .A2(n13243), .B1(n13138), .B2(n15575), .ZN(
        n13107) );
  INV_X1 U14811 ( .A(n13107), .ZN(n13108) );
  XNOR2_X1 U14812 ( .A(n13110), .B(n13111), .ZN(n13269) );
  INV_X1 U14813 ( .A(n13339), .ZN(n13114) );
  AOI22_X1 U14814 ( .A1(n15690), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13112), 
        .B2(n15680), .ZN(n13113) );
  OAI21_X1 U14815 ( .B1(n13114), .B2(n13250), .A(n13113), .ZN(n13115) );
  AOI21_X1 U14816 ( .B1(n13269), .B2(n13252), .A(n13115), .ZN(n13116) );
  OAI21_X1 U14817 ( .B1(n13271), .B2(n15690), .A(n13116), .ZN(P3_U3208) );
  OR2_X1 U14818 ( .A1(n13118), .A2(n13117), .ZN(n13119) );
  NAND2_X1 U14819 ( .A1(n13120), .A2(n13119), .ZN(n13344) );
  AND2_X1 U14820 ( .A1(n13140), .A2(n13121), .ZN(n13125) );
  NAND2_X1 U14821 ( .A1(n13140), .A2(n13122), .ZN(n13123) );
  OAI21_X1 U14822 ( .B1(n13125), .B2(n13124), .A(n13123), .ZN(n13126) );
  INV_X1 U14823 ( .A(n13126), .ZN(n13127) );
  OAI222_X1 U14824 ( .A1(n13243), .A2(n13128), .B1(n15575), .B2(n13158), .C1(
        n13240), .C2(n13127), .ZN(n13274) );
  NAND2_X1 U14825 ( .A1(n13274), .A2(n15688), .ZN(n13134) );
  INV_X1 U14826 ( .A(n13129), .ZN(n13131) );
  INV_X1 U14827 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13130) );
  OAI22_X1 U14828 ( .A1(n13131), .A2(n13143), .B1(n15688), .B2(n13130), .ZN(
        n13132) );
  AOI21_X1 U14829 ( .B1(n13276), .B2(n15684), .A(n13132), .ZN(n13133) );
  OAI211_X1 U14830 ( .C1(n13135), .C2(n13344), .A(n13134), .B(n13133), .ZN(
        P3_U3209) );
  AOI21_X1 U14831 ( .B1(n13099), .B2(n13136), .A(n13240), .ZN(n13141) );
  OAI22_X1 U14832 ( .A1(n13138), .A2(n13243), .B1(n13137), .B2(n15575), .ZN(
        n13139) );
  AOI21_X1 U14833 ( .B1(n13141), .B2(n13140), .A(n13139), .ZN(n13281) );
  INV_X1 U14834 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13145) );
  INV_X1 U14835 ( .A(n13142), .ZN(n13144) );
  OAI22_X1 U14836 ( .A1(n15688), .A2(n13145), .B1(n13144), .B2(n13143), .ZN(
        n13146) );
  AOI21_X1 U14837 ( .B1(n13147), .B2(n15684), .A(n13146), .ZN(n13152) );
  NAND2_X1 U14838 ( .A1(n13150), .A2(n13149), .ZN(n13279) );
  NAND3_X1 U14839 ( .A1(n13148), .A2(n13279), .A3(n13252), .ZN(n13151) );
  OAI211_X1 U14840 ( .C1(n13281), .C2(n15690), .A(n13152), .B(n13151), .ZN(
        P3_U3210) );
  XNOR2_X1 U14841 ( .A(n13154), .B(n13153), .ZN(n13354) );
  INV_X1 U14842 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13162) );
  XNOR2_X1 U14843 ( .A(n13156), .B(n13155), .ZN(n13161) );
  NOR2_X1 U14844 ( .A1(n13354), .A2(n15733), .ZN(n13160) );
  OAI22_X1 U14845 ( .A1(n13158), .A2(n13243), .B1(n13157), .B2(n15575), .ZN(
        n13159) );
  AOI211_X1 U14846 ( .C1(n13161), .C2(n15577), .A(n13160), .B(n13159), .ZN(
        n13349) );
  MUX2_X1 U14847 ( .A(n13162), .B(n13349), .S(n15688), .Z(n13165) );
  AOI22_X1 U14848 ( .A1(n13351), .A2(n15684), .B1(n15680), .B2(n13163), .ZN(
        n13164) );
  OAI211_X1 U14849 ( .C1(n13354), .C2(n13195), .A(n13165), .B(n13164), .ZN(
        P3_U3211) );
  XNOR2_X1 U14850 ( .A(n13166), .B(n9940), .ZN(n13357) );
  NAND2_X1 U14851 ( .A1(n13168), .A2(n13169), .ZN(n13170) );
  NAND2_X1 U14852 ( .A1(n13167), .A2(n13170), .ZN(n13171) );
  NAND2_X1 U14853 ( .A1(n13171), .A2(n15577), .ZN(n13175) );
  AOI22_X1 U14854 ( .A1(n15545), .A2(n13173), .B1(n13172), .B2(n15547), .ZN(
        n13174) );
  OAI211_X1 U14855 ( .C1(n15733), .C2(n13357), .A(n13175), .B(n13174), .ZN(
        n13355) );
  MUX2_X1 U14856 ( .A(n13355), .B(P3_REG2_REG_21__SCAN_IN), .S(n15690), .Z(
        n13176) );
  INV_X1 U14857 ( .A(n13176), .ZN(n13180) );
  AOI22_X1 U14858 ( .A1(n13178), .A2(n15684), .B1(n15680), .B2(n13177), .ZN(
        n13179) );
  OAI211_X1 U14859 ( .C1(n13357), .C2(n13195), .A(n13180), .B(n13179), .ZN(
        P3_U3212) );
  INV_X1 U14860 ( .A(n13181), .ZN(n13182) );
  INV_X1 U14861 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13191) );
  XNOR2_X1 U14862 ( .A(n13184), .B(n13185), .ZN(n13190) );
  AOI22_X1 U14863 ( .A1(n13187), .A2(n15545), .B1(n15547), .B2(n13186), .ZN(
        n13188) );
  OAI21_X1 U14864 ( .B1(n13366), .B2(n15733), .A(n13188), .ZN(n13189) );
  AOI21_X1 U14865 ( .B1(n13190), .B2(n15577), .A(n13189), .ZN(n13360) );
  MUX2_X1 U14866 ( .A(n13191), .B(n13360), .S(n15688), .Z(n13194) );
  AOI22_X1 U14867 ( .A1(n13362), .A2(n15684), .B1(n15680), .B2(n13192), .ZN(
        n13193) );
  OAI211_X1 U14868 ( .C1(n13366), .C2(n13195), .A(n13194), .B(n13193), .ZN(
        P3_U3213) );
  XNOR2_X1 U14869 ( .A(n13197), .B(n13196), .ZN(n13201) );
  OAI22_X1 U14870 ( .A1(n13199), .A2(n13243), .B1(n13198), .B2(n15575), .ZN(
        n13200) );
  AOI21_X1 U14871 ( .B1(n13201), .B2(n15577), .A(n13200), .ZN(n13294) );
  XNOR2_X1 U14872 ( .A(n13202), .B(n13203), .ZN(n13292) );
  AOI22_X1 U14873 ( .A1(n15690), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15680), 
        .B2(n13204), .ZN(n13205) );
  OAI21_X1 U14874 ( .B1(n13206), .B2(n13250), .A(n13205), .ZN(n13207) );
  AOI21_X1 U14875 ( .B1(n13292), .B2(n13252), .A(n13207), .ZN(n13208) );
  OAI21_X1 U14876 ( .B1(n13294), .B2(n15690), .A(n13208), .ZN(P3_U3214) );
  INV_X1 U14877 ( .A(n13209), .ZN(n13210) );
  AOI21_X1 U14878 ( .B1(n13215), .B2(n13211), .A(n13210), .ZN(n13212) );
  OAI222_X1 U14879 ( .A1(n13243), .A2(n13213), .B1(n15575), .B2(n13242), .C1(
        n13240), .C2(n13212), .ZN(n13297) );
  INV_X1 U14880 ( .A(n13297), .ZN(n13221) );
  OAI21_X1 U14881 ( .B1(n13216), .B2(n13215), .A(n13214), .ZN(n13298) );
  AOI22_X1 U14882 ( .A1(n15690), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15680), 
        .B2(n13217), .ZN(n13218) );
  OAI21_X1 U14883 ( .B1(n13374), .B2(n13250), .A(n13218), .ZN(n13219) );
  AOI21_X1 U14884 ( .B1(n13298), .B2(n13252), .A(n13219), .ZN(n13220) );
  OAI21_X1 U14885 ( .B1(n13221), .B2(n15690), .A(n13220), .ZN(P3_U3215) );
  OAI211_X1 U14886 ( .C1(n7236), .C2(n13223), .A(n15577), .B(n13222), .ZN(
        n13227) );
  AOI22_X1 U14887 ( .A1(n15547), .A2(n13225), .B1(n13224), .B2(n15545), .ZN(
        n13226) );
  NAND2_X1 U14888 ( .A1(n13227), .A2(n13226), .ZN(n13301) );
  INV_X1 U14889 ( .A(n13301), .ZN(n13235) );
  OAI21_X1 U14890 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(n13302) );
  AOI22_X1 U14891 ( .A1(n15690), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13231), 
        .B2(n15680), .ZN(n13232) );
  OAI21_X1 U14892 ( .B1(n13378), .B2(n13250), .A(n13232), .ZN(n13233) );
  AOI21_X1 U14893 ( .B1(n13302), .B2(n13252), .A(n13233), .ZN(n13234) );
  OAI21_X1 U14894 ( .B1(n13235), .B2(n15690), .A(n13234), .ZN(P3_U3216) );
  INV_X1 U14895 ( .A(n13236), .ZN(n13237) );
  AOI21_X1 U14896 ( .B1(n13245), .B2(n13238), .A(n13237), .ZN(n13239) );
  OAI222_X1 U14897 ( .A1(n13243), .A2(n13242), .B1(n15575), .B2(n13241), .C1(
        n13240), .C2(n13239), .ZN(n13305) );
  INV_X1 U14898 ( .A(n13305), .ZN(n13254) );
  OAI21_X1 U14899 ( .B1(n13246), .B2(n13245), .A(n13244), .ZN(n13306) );
  INV_X1 U14900 ( .A(n13247), .ZN(n13382) );
  AOI22_X1 U14901 ( .A1(n15690), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15680), 
        .B2(n13248), .ZN(n13249) );
  OAI21_X1 U14902 ( .B1(n13382), .B2(n13250), .A(n13249), .ZN(n13251) );
  AOI21_X1 U14903 ( .B1(n13306), .B2(n13252), .A(n13251), .ZN(n13253) );
  OAI21_X1 U14904 ( .B1(n13254), .B2(n15690), .A(n13253), .ZN(P3_U3217) );
  NAND2_X1 U14905 ( .A1(n15970), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13256) );
  INV_X1 U14906 ( .A(n15979), .ZN(n13255) );
  NAND2_X1 U14907 ( .A1(n13255), .A2(n15839), .ZN(n15972) );
  OAI211_X1 U14908 ( .C1(n13319), .C2(n13316), .A(n13256), .B(n15972), .ZN(
        P3_U3490) );
  NAND2_X1 U14909 ( .A1(n13257), .A2(n15802), .ZN(n13258) );
  INV_X1 U14910 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13260) );
  OAI21_X1 U14911 ( .B1(n13323), .B2(n13316), .A(n13261), .ZN(P3_U3487) );
  INV_X1 U14912 ( .A(n15732), .ZN(n15793) );
  NAND2_X1 U14913 ( .A1(n15839), .A2(n15793), .ZN(n15676) );
  INV_X1 U14914 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13262) );
  MUX2_X1 U14915 ( .A(n13262), .B(n13324), .S(n15839), .Z(n13264) );
  NAND2_X1 U14916 ( .A1(n13326), .A2(n15971), .ZN(n13263) );
  OAI211_X1 U14917 ( .C1(n13265), .C2(n15676), .A(n13264), .B(n13263), .ZN(
        P3_U3486) );
  INV_X1 U14918 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13266) );
  MUX2_X1 U14919 ( .A(n13266), .B(n13331), .S(n15839), .Z(n13268) );
  NAND2_X1 U14920 ( .A1(n13333), .A2(n15971), .ZN(n13267) );
  OAI211_X1 U14921 ( .C1(n13336), .C2(n15676), .A(n13268), .B(n13267), .ZN(
        P3_U3485) );
  NAND2_X1 U14922 ( .A1(n13269), .A2(n15802), .ZN(n13270) );
  NAND2_X1 U14923 ( .A1(n13271), .A2(n13270), .ZN(n13337) );
  MUX2_X1 U14924 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13337), .S(n15839), .Z(
        n13272) );
  AOI21_X1 U14925 ( .B1(n15971), .B2(n13339), .A(n13272), .ZN(n13273) );
  INV_X1 U14926 ( .A(n13273), .ZN(P3_U3484) );
  INV_X1 U14927 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13277) );
  NOR2_X1 U14928 ( .A1(n13344), .A2(n15733), .ZN(n13275) );
  AOI211_X1 U14929 ( .C1(n15737), .C2(n13276), .A(n13275), .B(n13274), .ZN(
        n13341) );
  MUX2_X1 U14930 ( .A(n13277), .B(n13341), .S(n15839), .Z(n13278) );
  OAI21_X1 U14931 ( .B1(n13344), .B2(n15676), .A(n13278), .ZN(P3_U3483) );
  NAND3_X1 U14932 ( .A1(n13148), .A2(n13279), .A3(n15802), .ZN(n13280) );
  AND2_X1 U14933 ( .A1(n13281), .A2(n13280), .ZN(n13346) );
  INV_X1 U14934 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13282) );
  MUX2_X1 U14935 ( .A(n13346), .B(n13282), .S(n15970), .Z(n13283) );
  OAI21_X1 U14936 ( .B1(n13348), .B2(n13316), .A(n13283), .ZN(P3_U3482) );
  MUX2_X1 U14937 ( .A(n13284), .B(n13349), .S(n15839), .Z(n13286) );
  NAND2_X1 U14938 ( .A1(n13351), .A2(n15971), .ZN(n13285) );
  OAI211_X1 U14939 ( .C1(n13354), .C2(n15676), .A(n13286), .B(n13285), .ZN(
        P3_U3481) );
  MUX2_X1 U14940 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13355), .S(n15839), .Z(
        n13288) );
  OAI22_X1 U14941 ( .A1(n13357), .A2(n15676), .B1(n13356), .B2(n13316), .ZN(
        n13287) );
  OR2_X1 U14942 ( .A1(n13288), .A2(n13287), .ZN(P3_U3480) );
  INV_X1 U14943 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13289) );
  MUX2_X1 U14944 ( .A(n13289), .B(n13360), .S(n15839), .Z(n13291) );
  NAND2_X1 U14945 ( .A1(n13362), .A2(n15971), .ZN(n13290) );
  OAI211_X1 U14946 ( .C1(n13366), .C2(n15676), .A(n13291), .B(n13290), .ZN(
        P3_U3479) );
  NAND2_X1 U14947 ( .A1(n13292), .A2(n15802), .ZN(n13293) );
  NAND2_X1 U14948 ( .A1(n13294), .A2(n13293), .ZN(n13367) );
  MUX2_X1 U14949 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13367), .S(n15839), .Z(
        n13295) );
  AOI21_X1 U14950 ( .B1(n15971), .B2(n13369), .A(n13295), .ZN(n13296) );
  INV_X1 U14951 ( .A(n13296), .ZN(P3_U3478) );
  AOI21_X1 U14952 ( .B1(n15802), .B2(n13298), .A(n13297), .ZN(n13371) );
  MUX2_X1 U14953 ( .A(n13299), .B(n13371), .S(n15839), .Z(n13300) );
  OAI21_X1 U14954 ( .B1(n13374), .B2(n13316), .A(n13300), .ZN(P3_U3477) );
  AOI21_X1 U14955 ( .B1(n15802), .B2(n13302), .A(n13301), .ZN(n13375) );
  MUX2_X1 U14956 ( .A(n13303), .B(n13375), .S(n15839), .Z(n13304) );
  OAI21_X1 U14957 ( .B1(n13316), .B2(n13378), .A(n13304), .ZN(P3_U3476) );
  AOI21_X1 U14958 ( .B1(n15802), .B2(n13306), .A(n13305), .ZN(n13379) );
  MUX2_X1 U14959 ( .A(n15509), .B(n13379), .S(n15839), .Z(n13307) );
  OAI21_X1 U14960 ( .B1(n13382), .B2(n13316), .A(n13307), .ZN(P3_U3475) );
  AOI21_X1 U14961 ( .B1(n15802), .B2(n13309), .A(n13308), .ZN(n13383) );
  MUX2_X1 U14962 ( .A(n13310), .B(n13383), .S(n15839), .Z(n13311) );
  OAI21_X1 U14963 ( .B1(n13316), .B2(n13386), .A(n13311), .ZN(P3_U3474) );
  AOI21_X1 U14964 ( .B1(n15802), .B2(n13313), .A(n13312), .ZN(n13387) );
  MUX2_X1 U14965 ( .A(n13314), .B(n13387), .S(n15839), .Z(n13315) );
  OAI21_X1 U14966 ( .B1(n13316), .B2(n13390), .A(n13315), .ZN(P3_U3473) );
  NOR2_X1 U14967 ( .A1(n15979), .A2(n15980), .ZN(n13317) );
  AOI21_X1 U14968 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15980), .A(n13317), 
        .ZN(n13318) );
  OAI21_X1 U14969 ( .B1(n13319), .B2(n13391), .A(n13318), .ZN(P3_U3458) );
  OAI21_X1 U14970 ( .B1(n13323), .B2(n13391), .A(n13322), .ZN(P3_U3455) );
  MUX2_X1 U14971 ( .A(n13325), .B(n13324), .S(n15978), .Z(n13329) );
  AOI22_X1 U14972 ( .A1(n13327), .A2(n13330), .B1(n15974), .B2(n13326), .ZN(
        n13328) );
  NAND2_X1 U14973 ( .A1(n13329), .A2(n13328), .ZN(P3_U3454) );
  INV_X1 U14974 ( .A(n13330), .ZN(n13365) );
  MUX2_X1 U14975 ( .A(n13332), .B(n13331), .S(n15978), .Z(n13335) );
  NAND2_X1 U14976 ( .A1(n13333), .A2(n15974), .ZN(n13334) );
  OAI211_X1 U14977 ( .C1(n13336), .C2(n13365), .A(n13335), .B(n13334), .ZN(
        P3_U3453) );
  MUX2_X1 U14978 ( .A(n13337), .B(P3_REG0_REG_25__SCAN_IN), .S(n15980), .Z(
        n13338) );
  AOI21_X1 U14979 ( .B1(n15974), .B2(n13339), .A(n13338), .ZN(n13340) );
  INV_X1 U14980 ( .A(n13340), .ZN(P3_U3452) );
  MUX2_X1 U14981 ( .A(n13342), .B(n13341), .S(n15978), .Z(n13343) );
  OAI21_X1 U14982 ( .B1(n13344), .B2(n13365), .A(n13343), .ZN(P3_U3451) );
  INV_X1 U14983 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13345) );
  MUX2_X1 U14984 ( .A(n13346), .B(n13345), .S(n15980), .Z(n13347) );
  OAI21_X1 U14985 ( .B1(n13348), .B2(n13391), .A(n13347), .ZN(P3_U3450) );
  INV_X1 U14986 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13350) );
  MUX2_X1 U14987 ( .A(n13350), .B(n13349), .S(n15978), .Z(n13353) );
  NAND2_X1 U14988 ( .A1(n13351), .A2(n15974), .ZN(n13352) );
  OAI211_X1 U14989 ( .C1(n13354), .C2(n13365), .A(n13353), .B(n13352), .ZN(
        P3_U3449) );
  MUX2_X1 U14990 ( .A(n13355), .B(P3_REG0_REG_21__SCAN_IN), .S(n15980), .Z(
        n13359) );
  OAI22_X1 U14991 ( .A1(n13357), .A2(n13365), .B1(n13356), .B2(n13391), .ZN(
        n13358) );
  OR2_X1 U14992 ( .A1(n13359), .A2(n13358), .ZN(P3_U3448) );
  INV_X1 U14993 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13361) );
  MUX2_X1 U14994 ( .A(n13361), .B(n13360), .S(n15978), .Z(n13364) );
  NAND2_X1 U14995 ( .A1(n13362), .A2(n15974), .ZN(n13363) );
  OAI211_X1 U14996 ( .C1(n13366), .C2(n13365), .A(n13364), .B(n13363), .ZN(
        P3_U3447) );
  MUX2_X1 U14997 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13367), .S(n15978), .Z(
        n13368) );
  AOI21_X1 U14998 ( .B1(n15974), .B2(n13369), .A(n13368), .ZN(n13370) );
  INV_X1 U14999 ( .A(n13370), .ZN(P3_U3446) );
  INV_X1 U15000 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13372) );
  MUX2_X1 U15001 ( .A(n13372), .B(n13371), .S(n15978), .Z(n13373) );
  OAI21_X1 U15002 ( .B1(n13374), .B2(n13391), .A(n13373), .ZN(P3_U3444) );
  INV_X1 U15003 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13376) );
  MUX2_X1 U15004 ( .A(n13376), .B(n13375), .S(n15978), .Z(n13377) );
  OAI21_X1 U15005 ( .B1(n13391), .B2(n13378), .A(n13377), .ZN(P3_U3441) );
  INV_X1 U15006 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13380) );
  MUX2_X1 U15007 ( .A(n13380), .B(n13379), .S(n15978), .Z(n13381) );
  OAI21_X1 U15008 ( .B1(n13382), .B2(n13391), .A(n13381), .ZN(P3_U3438) );
  INV_X1 U15009 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13384) );
  MUX2_X1 U15010 ( .A(n13384), .B(n13383), .S(n15978), .Z(n13385) );
  OAI21_X1 U15011 ( .B1(n13391), .B2(n13386), .A(n13385), .ZN(P3_U3435) );
  INV_X1 U15012 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13388) );
  MUX2_X1 U15013 ( .A(n13388), .B(n13387), .S(n15978), .Z(n13389) );
  OAI21_X1 U15014 ( .B1(n13391), .B2(n13390), .A(n13389), .ZN(P3_U3432) );
  MUX2_X1 U15015 ( .A(P3_D_REG_1__SCAN_IN), .B(n13392), .S(n13393), .Z(
        P3_U3377) );
  MUX2_X1 U15016 ( .A(P3_D_REG_0__SCAN_IN), .B(n13394), .S(n13393), .Z(
        P3_U3376) );
  INV_X1 U15017 ( .A(n13395), .ZN(n13399) );
  NOR4_X1 U15018 ( .A1(n9595), .A2(P3_IR_REG_30__SCAN_IN), .A3(n9879), .A4(
        P3_U3151), .ZN(n13396) );
  AOI21_X1 U15019 ( .B1(SI_31_), .B2(n13397), .A(n13396), .ZN(n13398) );
  OAI21_X1 U15020 ( .B1(n13399), .B2(n13402), .A(n13398), .ZN(P3_U3264) );
  INV_X1 U15021 ( .A(SI_30_), .ZN(n15023) );
  INV_X1 U15022 ( .A(n13400), .ZN(n13401) );
  OAI222_X1 U15023 ( .A1(n13405), .A2(P3_U3151), .B1(n13403), .B2(n15023), 
        .C1(n13402), .C2(n13401), .ZN(P3_U3265) );
  MUX2_X1 U15024 ( .A(n13406), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15025 ( .B1(n13407), .B2(n13408), .A(n13486), .ZN(n13410) );
  NAND2_X1 U15026 ( .A1(n13410), .A2(n13409), .ZN(n13416) );
  OAI22_X1 U15027 ( .A1(n13690), .A2(n14057), .B1(n13411), .B2(n14055), .ZN(
        n13914) );
  INV_X1 U15028 ( .A(n13924), .ZN(n13413) );
  OAI22_X1 U15029 ( .A1(n13413), .A2(n13479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13412), .ZN(n13414) );
  AOI21_X1 U15030 ( .B1(n13914), .B2(n13513), .A(n13414), .ZN(n13415) );
  OAI211_X1 U15031 ( .C1(n14187), .C2(n13506), .A(n13416), .B(n13415), .ZN(
        P2_U3186) );
  OAI22_X1 U15032 ( .A1(n13417), .A2(n13486), .B1(n13667), .B2(n13484), .ZN(
        n13419) );
  NAND2_X1 U15033 ( .A1(n13419), .A2(n13418), .ZN(n13425) );
  INV_X1 U15034 ( .A(n13420), .ZN(n13997) );
  OAI22_X1 U15035 ( .A1(n13665), .A2(n14057), .B1(n13485), .B2(n14055), .ZN(
        n13421) );
  INV_X1 U15036 ( .A(n13421), .ZN(n13992) );
  OAI22_X1 U15037 ( .A1(n13992), .A2(n13492), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13422), .ZN(n13423) );
  AOI21_X1 U15038 ( .B1(n13997), .B2(n13515), .A(n13423), .ZN(n13424) );
  OAI211_X1 U15039 ( .C1(n14204), .C2(n13506), .A(n13425), .B(n13424), .ZN(
        P2_U3188) );
  AOI22_X1 U15040 ( .A1(n13439), .A2(n13799), .B1(n13438), .B2(n13798), .ZN(
        n13426) );
  NAND2_X1 U15041 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n15197)
         );
  OAI211_X1 U15042 ( .C1(n13479), .C2(n14049), .A(n13426), .B(n15197), .ZN(
        n13436) );
  NOR3_X1 U15043 ( .A1(n13427), .A2(n8055), .A3(n13486), .ZN(n13434) );
  NAND2_X1 U15044 ( .A1(n13428), .A2(n14072), .ZN(n13429) );
  OAI22_X1 U15045 ( .A1(n13431), .A2(n13486), .B1(n13430), .B2(n13429), .ZN(
        n13433) );
  MUX2_X1 U15046 ( .A(n13434), .B(n13433), .S(n13432), .Z(n13435) );
  AOI211_X1 U15047 ( .C1(n14048), .C2(n13516), .A(n13436), .B(n13435), .ZN(
        n13437) );
  INV_X1 U15048 ( .A(n13437), .ZN(P2_U3191) );
  AOI22_X1 U15049 ( .A1(n13439), .A2(n13528), .B1(n13438), .B2(n13815), .ZN(
        n13446) );
  AOI22_X1 U15050 ( .A1(n13516), .A2(n13534), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13440), .ZN(n13445) );
  OAI21_X1 U15051 ( .B1(n13442), .B2(n13441), .A(n11127), .ZN(n13443) );
  NAND2_X1 U15052 ( .A1(n13507), .A2(n13443), .ZN(n13444) );
  NAND3_X1 U15053 ( .A1(n13446), .A2(n13445), .A3(n13444), .ZN(P2_U3194) );
  OAI211_X1 U15054 ( .C1(n13449), .C2(n13448), .A(n13447), .B(n13507), .ZN(
        n13454) );
  INV_X1 U15055 ( .A(n13450), .ZN(n14022) );
  AOI22_X1 U15056 ( .A1(n13796), .A2(n14071), .B1(n14069), .B2(n13798), .ZN(
        n14019) );
  OAI22_X1 U15057 ( .A1(n14019), .A2(n13492), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13451), .ZN(n13452) );
  AOI21_X1 U15058 ( .B1(n14022), .B2(n13515), .A(n13452), .ZN(n13453) );
  OAI211_X1 U15059 ( .C1(n7587), .C2(n13506), .A(n13454), .B(n13453), .ZN(
        P2_U3195) );
  INV_X1 U15060 ( .A(n13456), .ZN(n13457) );
  AOI21_X1 U15061 ( .B1(n13455), .B2(n13457), .A(n13486), .ZN(n13460) );
  NOR3_X1 U15062 ( .A1(n13458), .A2(n13665), .A3(n13484), .ZN(n13459) );
  OAI21_X1 U15063 ( .B1(n13460), .B2(n13459), .A(n12559), .ZN(n13466) );
  NAND2_X1 U15064 ( .A1(n13792), .A2(n14071), .ZN(n13462) );
  NAND2_X1 U15065 ( .A1(n13794), .A2(n14069), .ZN(n13461) );
  NAND2_X1 U15066 ( .A1(n13462), .A2(n13461), .ZN(n13955) );
  OAI22_X1 U15067 ( .A1(n13960), .A2(n13479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13463), .ZN(n13464) );
  AOI21_X1 U15068 ( .B1(n13955), .B2(n13513), .A(n13464), .ZN(n13465) );
  OAI211_X1 U15069 ( .C1(n14195), .C2(n13506), .A(n13466), .B(n13465), .ZN(
        P2_U3197) );
  OAI211_X1 U15070 ( .C1(n13468), .C2(n13467), .A(n13455), .B(n13507), .ZN(
        n13473) );
  OAI22_X1 U15071 ( .A1(n13664), .A2(n14057), .B1(n13667), .B2(n14055), .ZN(
        n13974) );
  INV_X1 U15072 ( .A(n13981), .ZN(n13470) );
  OAI22_X1 U15073 ( .A1(n13470), .A2(n13479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13469), .ZN(n13471) );
  AOI21_X1 U15074 ( .B1(n13974), .B2(n13513), .A(n13471), .ZN(n13472) );
  OAI211_X1 U15075 ( .C1(n14200), .C2(n13506), .A(n13473), .B(n13472), .ZN(
        P2_U3201) );
  XNOR2_X1 U15076 ( .A(n7190), .B(n13474), .ZN(n13475) );
  XNOR2_X1 U15077 ( .A(n13476), .B(n13475), .ZN(n13483) );
  INV_X1 U15078 ( .A(n14036), .ZN(n13478) );
  OAI22_X1 U15079 ( .A1(n13479), .A2(n13478), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13477), .ZN(n13481) );
  OAI22_X1 U15080 ( .A1(n14031), .A2(n13500), .B1(n13499), .B2(n14032), .ZN(
        n13480) );
  AOI211_X1 U15081 ( .C1(n14146), .C2(n13516), .A(n13481), .B(n13480), .ZN(
        n13482) );
  OAI21_X1 U15082 ( .B1(n13483), .B2(n13486), .A(n13482), .ZN(P2_U3205) );
  OAI22_X1 U15083 ( .A1(n13487), .A2(n13486), .B1(n13485), .B2(n13484), .ZN(
        n13489) );
  NAND2_X1 U15084 ( .A1(n13489), .A2(n13488), .ZN(n13495) );
  INV_X1 U15085 ( .A(n13490), .ZN(n14011) );
  AOI22_X1 U15086 ( .A1(n13795), .A2(n14071), .B1(n14069), .B2(n13797), .ZN(
        n14004) );
  OAI22_X1 U15087 ( .A1(n14004), .A2(n13492), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13491), .ZN(n13493) );
  AOI21_X1 U15088 ( .B1(n14011), .B2(n13515), .A(n13493), .ZN(n13494) );
  OAI211_X1 U15089 ( .C1(n7586), .C2(n13506), .A(n13495), .B(n13494), .ZN(
        P2_U3207) );
  INV_X1 U15090 ( .A(n14155), .ZN(n14080) );
  OAI211_X1 U15091 ( .C1(n13498), .C2(n13497), .A(n13496), .B(n13507), .ZN(
        n13505) );
  NAND2_X1 U15092 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n15182)
         );
  INV_X1 U15093 ( .A(n15182), .ZN(n13503) );
  OAI22_X1 U15094 ( .A1(n13501), .A2(n13500), .B1(n13499), .B2(n14031), .ZN(
        n13502) );
  AOI211_X1 U15095 ( .C1(n14078), .C2(n13515), .A(n13503), .B(n13502), .ZN(
        n13504) );
  OAI211_X1 U15096 ( .C1(n14080), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        P2_U3210) );
  OAI211_X1 U15097 ( .C1(n13510), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        n13519) );
  INV_X1 U15098 ( .A(n13511), .ZN(n13512) );
  AOI22_X1 U15099 ( .A1(n13513), .A2(n13512), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13518) );
  AOI22_X1 U15100 ( .A1(n13516), .A2(n13567), .B1(n13515), .B2(n13514), .ZN(
        n13517) );
  NAND3_X1 U15101 ( .A1(n13519), .A2(n13518), .A3(n13517), .ZN(P2_U3211) );
  INV_X1 U15102 ( .A(n15140), .ZN(n15137) );
  NOR4_X1 U15103 ( .A1(n15137), .A2(n14231), .A3(n13740), .A4(n14055), .ZN(
        n13787) );
  INV_X1 U15104 ( .A(n13782), .ZN(n13520) );
  OAI21_X1 U15105 ( .B1(n13520), .B2(n8832), .A(P2_B_REG_SCAN_IN), .ZN(n13786)
         );
  AND2_X4 U15106 ( .A1(n15758), .A2(n13779), .ZN(n13553) );
  INV_X4 U15107 ( .A(n13553), .ZN(n13703) );
  MUX2_X1 U15108 ( .A(n13522), .B(n13521), .S(n13703), .Z(n13537) );
  INV_X1 U15109 ( .A(n13741), .ZN(n13525) );
  NAND2_X1 U15110 ( .A1(n7193), .A2(n15194), .ZN(n13524) );
  NAND2_X1 U15111 ( .A1(n13525), .A2(n13524), .ZN(n13530) );
  NAND2_X1 U15112 ( .A1(n13526), .A2(n13530), .ZN(n13527) );
  NAND2_X1 U15113 ( .A1(n10973), .A2(n13527), .ZN(n13533) );
  NOR2_X1 U15114 ( .A1(n8134), .A2(n13531), .ZN(n13532) );
  MUX2_X1 U15115 ( .A(n13816), .B(n13534), .S(n13703), .Z(n13535) );
  NAND2_X1 U15116 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  MUX2_X1 U15117 ( .A(n13815), .B(n13540), .S(n13703), .Z(n13542) );
  MUX2_X1 U15118 ( .A(n13815), .B(n13540), .S(n13708), .Z(n13541) );
  INV_X1 U15119 ( .A(n13542), .ZN(n13543) );
  MUX2_X1 U15120 ( .A(n13544), .B(n13814), .S(n13703), .Z(n13548) );
  NAND2_X1 U15121 ( .A1(n13547), .A2(n13548), .ZN(n13546) );
  MUX2_X1 U15122 ( .A(n13544), .B(n13814), .S(n13708), .Z(n13545) );
  NAND2_X1 U15123 ( .A1(n13546), .A2(n13545), .ZN(n13552) );
  INV_X1 U15124 ( .A(n13547), .ZN(n13550) );
  INV_X1 U15125 ( .A(n13548), .ZN(n13549) );
  NAND2_X1 U15126 ( .A1(n13550), .A2(n13549), .ZN(n13551) );
  MUX2_X1 U15127 ( .A(n13813), .B(n13554), .S(n13703), .Z(n13557) );
  MUX2_X1 U15128 ( .A(n13813), .B(n13554), .S(n13708), .Z(n13555) );
  INV_X1 U15129 ( .A(n13557), .ZN(n13558) );
  MUX2_X1 U15130 ( .A(n13559), .B(n13811), .S(n13703), .Z(n13563) );
  MUX2_X1 U15131 ( .A(n13811), .B(n13559), .S(n13703), .Z(n13560) );
  NAND2_X1 U15132 ( .A1(n13561), .A2(n13560), .ZN(n13566) );
  INV_X1 U15133 ( .A(n13562), .ZN(n13564) );
  NAND2_X1 U15134 ( .A1(n13564), .A2(n7854), .ZN(n13565) );
  MUX2_X1 U15135 ( .A(n13567), .B(n13810), .S(n13708), .Z(n13571) );
  NAND2_X1 U15136 ( .A1(n13570), .A2(n13571), .ZN(n13569) );
  MUX2_X1 U15137 ( .A(n13567), .B(n13810), .S(n13703), .Z(n13568) );
  NAND2_X1 U15138 ( .A1(n13569), .A2(n13568), .ZN(n13575) );
  INV_X1 U15139 ( .A(n13570), .ZN(n13573) );
  INV_X1 U15140 ( .A(n13571), .ZN(n13572) );
  NAND2_X1 U15141 ( .A1(n13573), .A2(n13572), .ZN(n13574) );
  NAND2_X1 U15142 ( .A1(n13575), .A2(n13574), .ZN(n13578) );
  MUX2_X1 U15143 ( .A(n13576), .B(n13809), .S(n13703), .Z(n13579) );
  MUX2_X1 U15144 ( .A(n13576), .B(n13809), .S(n13708), .Z(n13577) );
  MUX2_X1 U15145 ( .A(n13808), .B(n13580), .S(n13703), .Z(n13584) );
  MUX2_X1 U15146 ( .A(n13808), .B(n13580), .S(n13708), .Z(n13581) );
  NAND2_X1 U15147 ( .A1(n13582), .A2(n13581), .ZN(n13586) );
  MUX2_X1 U15148 ( .A(n13807), .B(n13587), .S(n13708), .Z(n13589) );
  MUX2_X1 U15149 ( .A(n13807), .B(n13587), .S(n13703), .Z(n13588) );
  INV_X1 U15150 ( .A(n13589), .ZN(n13590) );
  MUX2_X1 U15151 ( .A(n13806), .B(n13591), .S(n13703), .Z(n13595) );
  NAND2_X1 U15152 ( .A1(n13594), .A2(n13595), .ZN(n13593) );
  MUX2_X1 U15153 ( .A(n13806), .B(n13591), .S(n13708), .Z(n13592) );
  NAND2_X1 U15154 ( .A1(n13593), .A2(n13592), .ZN(n13599) );
  INV_X1 U15155 ( .A(n13594), .ZN(n13597) );
  INV_X1 U15156 ( .A(n13595), .ZN(n13596) );
  NAND2_X1 U15157 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  MUX2_X1 U15158 ( .A(n13805), .B(n13600), .S(n13708), .Z(n13602) );
  MUX2_X1 U15159 ( .A(n13805), .B(n13600), .S(n13703), .Z(n13601) );
  MUX2_X1 U15160 ( .A(n13804), .B(n13603), .S(n13703), .Z(n13607) );
  NAND2_X1 U15161 ( .A1(n13606), .A2(n13607), .ZN(n13605) );
  MUX2_X1 U15162 ( .A(n13804), .B(n13603), .S(n13708), .Z(n13604) );
  NAND2_X1 U15163 ( .A1(n13605), .A2(n13604), .ZN(n13611) );
  INV_X1 U15164 ( .A(n13606), .ZN(n13609) );
  INV_X1 U15165 ( .A(n13607), .ZN(n13608) );
  NAND2_X1 U15166 ( .A1(n13609), .A2(n13608), .ZN(n13610) );
  NAND2_X1 U15167 ( .A1(n13611), .A2(n13610), .ZN(n13614) );
  MUX2_X1 U15168 ( .A(n13803), .B(n13612), .S(n13708), .Z(n13615) );
  MUX2_X1 U15169 ( .A(n13803), .B(n13612), .S(n13703), .Z(n13613) );
  MUX2_X1 U15170 ( .A(n13802), .B(n15862), .S(n13703), .Z(n13619) );
  MUX2_X1 U15171 ( .A(n13802), .B(n15862), .S(n13708), .Z(n13616) );
  NAND2_X1 U15172 ( .A1(n13617), .A2(n13616), .ZN(n13621) );
  MUX2_X1 U15173 ( .A(n13801), .B(n13622), .S(n13708), .Z(n13624) );
  MUX2_X1 U15174 ( .A(n13801), .B(n13622), .S(n13703), .Z(n13623) );
  INV_X1 U15175 ( .A(n13624), .ZN(n13625) );
  MUX2_X1 U15176 ( .A(n13800), .B(n13626), .S(n13703), .Z(n13630) );
  NAND2_X1 U15177 ( .A1(n13629), .A2(n13630), .ZN(n13628) );
  MUX2_X1 U15178 ( .A(n13626), .B(n13800), .S(n13703), .Z(n13627) );
  NAND2_X1 U15179 ( .A1(n13628), .A2(n13627), .ZN(n13634) );
  INV_X1 U15180 ( .A(n13629), .ZN(n13632) );
  INV_X1 U15181 ( .A(n13630), .ZN(n13631) );
  NAND2_X1 U15182 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  MUX2_X1 U15183 ( .A(n14070), .B(n13635), .S(n13708), .Z(n13637) );
  MUX2_X1 U15184 ( .A(n14070), .B(n13635), .S(n13703), .Z(n13636) );
  INV_X1 U15185 ( .A(n13637), .ZN(n13638) );
  MUX2_X1 U15186 ( .A(n14155), .B(n13799), .S(n13708), .Z(n13642) );
  NAND2_X1 U15187 ( .A1(n13641), .A2(n13642), .ZN(n13640) );
  MUX2_X1 U15188 ( .A(n14155), .B(n13799), .S(n13703), .Z(n13639) );
  NAND2_X1 U15189 ( .A1(n13640), .A2(n13639), .ZN(n13646) );
  INV_X1 U15190 ( .A(n13641), .ZN(n13644) );
  INV_X1 U15191 ( .A(n13642), .ZN(n13643) );
  NAND2_X1 U15192 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U15193 ( .A1(n13646), .A2(n13645), .ZN(n13648) );
  MUX2_X1 U15194 ( .A(n14072), .B(n14048), .S(n13553), .Z(n13649) );
  MUX2_X1 U15195 ( .A(n14072), .B(n14048), .S(n13703), .Z(n13647) );
  INV_X1 U15196 ( .A(n13649), .ZN(n13650) );
  MUX2_X1 U15197 ( .A(n13798), .B(n14146), .S(n13703), .Z(n13654) );
  MUX2_X1 U15198 ( .A(n13798), .B(n14146), .S(n13553), .Z(n13651) );
  NAND2_X1 U15199 ( .A1(n13652), .A2(n13651), .ZN(n13655) );
  NAND2_X1 U15200 ( .A1(n13655), .A2(n7268), .ZN(n13657) );
  MUX2_X1 U15201 ( .A(n13797), .B(n14141), .S(n13708), .Z(n13658) );
  MUX2_X1 U15202 ( .A(n13797), .B(n14141), .S(n13703), .Z(n13656) );
  MUX2_X1 U15203 ( .A(n13796), .B(n14010), .S(n13703), .Z(n13662) );
  MUX2_X1 U15204 ( .A(n13796), .B(n14010), .S(n13708), .Z(n13659) );
  NAND2_X1 U15205 ( .A1(n13660), .A2(n13659), .ZN(n13663) );
  NAND2_X1 U15206 ( .A1(n13663), .A2(n7269), .ZN(n13670) );
  MUX2_X1 U15207 ( .A(n13795), .B(n13994), .S(n13553), .Z(n13669) );
  MUX2_X1 U15208 ( .A(n13664), .B(n14195), .S(n13708), .Z(n13674) );
  MUX2_X1 U15209 ( .A(n13793), .B(n13965), .S(n13703), .Z(n13673) );
  NAND2_X1 U15210 ( .A1(n13674), .A2(n13673), .ZN(n13678) );
  MUX2_X1 U15211 ( .A(n13665), .B(n14200), .S(n13708), .Z(n13672) );
  MUX2_X1 U15212 ( .A(n13794), .B(n14126), .S(n13703), .Z(n13671) );
  NAND2_X1 U15213 ( .A1(n13672), .A2(n13671), .ZN(n13666) );
  MUX2_X1 U15214 ( .A(n13667), .B(n14204), .S(n13703), .Z(n13668) );
  NOR2_X1 U15215 ( .A1(n13672), .A2(n13671), .ZN(n13677) );
  INV_X1 U15216 ( .A(n13673), .ZN(n13676) );
  INV_X1 U15217 ( .A(n13674), .ZN(n13675) );
  AOI22_X1 U15218 ( .A1(n13678), .A2(n13677), .B1(n13676), .B2(n13675), .ZN(
        n13681) );
  MUX2_X1 U15219 ( .A(n13944), .B(n13792), .S(n13708), .Z(n13695) );
  INV_X1 U15220 ( .A(n13695), .ZN(n13679) );
  MUX2_X1 U15221 ( .A(n13944), .B(n13792), .S(n13703), .Z(n13694) );
  NAND2_X1 U15222 ( .A1(n13679), .A2(n13694), .ZN(n13680) );
  NAND2_X1 U15223 ( .A1(n13683), .A2(n13704), .ZN(n13685) );
  NAND2_X1 U15224 ( .A1(n8420), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13684) );
  INV_X1 U15225 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U15226 ( .A1(n8306), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n13687) );
  NAND2_X1 U15227 ( .A1(n8709), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13686) );
  OAI211_X1 U15228 ( .C1(n8572), .C2(n14175), .A(n13687), .B(n13686), .ZN(
        n13884) );
  XNOR2_X1 U15229 ( .A(n14090), .B(n13884), .ZN(n13718) );
  MUX2_X1 U15230 ( .A(n13689), .B(n13688), .S(n13708), .Z(n13715) );
  MUX2_X1 U15231 ( .A(n13789), .B(n14096), .S(n13703), .Z(n13714) );
  NAND2_X1 U15232 ( .A1(n13715), .A2(n13714), .ZN(n13722) );
  MUX2_X1 U15233 ( .A(n13690), .B(n14183), .S(n13708), .Z(n13720) );
  MUX2_X1 U15234 ( .A(n13790), .B(n14104), .S(n13703), .Z(n13719) );
  NAND2_X1 U15235 ( .A1(n13720), .A2(n13719), .ZN(n13691) );
  AND2_X1 U15236 ( .A1(n13722), .A2(n13691), .ZN(n13692) );
  AND2_X1 U15237 ( .A1(n13718), .A2(n13692), .ZN(n13702) );
  MUX2_X1 U15238 ( .A(n14187), .B(n13693), .S(n13703), .Z(n13699) );
  MUX2_X1 U15239 ( .A(n13791), .B(n13923), .S(n13703), .Z(n13698) );
  INV_X1 U15240 ( .A(n13694), .ZN(n13696) );
  AOI22_X1 U15241 ( .A1(n13699), .A2(n13698), .B1(n13696), .B2(n13695), .ZN(
        n13697) );
  INV_X1 U15242 ( .A(n13698), .ZN(n13701) );
  INV_X1 U15243 ( .A(n13699), .ZN(n13700) );
  NAND3_X1 U15244 ( .A1(n13702), .A2(n13701), .A3(n13700), .ZN(n13726) );
  NAND2_X1 U15245 ( .A1(n13884), .A2(n13703), .ZN(n13711) );
  MUX2_X1 U15246 ( .A(n13711), .B(n13884), .S(n14090), .Z(n13717) );
  NAND2_X1 U15247 ( .A1(n13705), .A2(n13704), .ZN(n13707) );
  NAND2_X1 U15248 ( .A1(n8420), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13706) );
  MUX2_X1 U15249 ( .A(n13883), .B(n13788), .S(n13708), .Z(n13728) );
  AND2_X1 U15250 ( .A1(n8832), .A2(n13780), .ZN(n13734) );
  NOR2_X1 U15251 ( .A1(n13734), .A2(n13709), .ZN(n13712) );
  INV_X1 U15252 ( .A(n13788), .ZN(n13710) );
  AOI21_X1 U15253 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(n13713) );
  AOI21_X1 U15254 ( .B1(n13883), .B2(n13708), .A(n13713), .ZN(n13727) );
  OAI22_X1 U15255 ( .A1(n13728), .A2(n13727), .B1(n13715), .B2(n13714), .ZN(
        n13716) );
  NAND2_X1 U15256 ( .A1(n13717), .A2(n13716), .ZN(n13725) );
  INV_X1 U15257 ( .A(n13719), .ZN(n13723) );
  INV_X1 U15258 ( .A(n13720), .ZN(n13721) );
  NAND4_X1 U15259 ( .A1(n13718), .A2(n13723), .A3(n13722), .A4(n13721), .ZN(
        n13724) );
  NAND2_X1 U15260 ( .A1(n13728), .A2(n13727), .ZN(n13733) );
  INV_X1 U15261 ( .A(n13884), .ZN(n13729) );
  NOR2_X1 U15262 ( .A1(n14090), .A2(n13729), .ZN(n13731) );
  AND2_X1 U15263 ( .A1(n14090), .A2(n13729), .ZN(n13730) );
  MUX2_X1 U15264 ( .A(n13731), .B(n13730), .S(n13703), .Z(n13732) );
  NAND2_X1 U15265 ( .A1(n13779), .A2(n15194), .ZN(n13737) );
  INV_X1 U15266 ( .A(n13734), .ZN(n13735) );
  OAI21_X1 U15267 ( .B1(n13737), .B2(n13736), .A(n13735), .ZN(n13738) );
  INV_X1 U15268 ( .A(n13738), .ZN(n13744) );
  NAND2_X1 U15269 ( .A1(n13779), .A2(n13776), .ZN(n13739) );
  OAI211_X1 U15270 ( .C1(n13741), .C2(n8832), .A(n13740), .B(n13739), .ZN(
        n13742) );
  NAND2_X1 U15271 ( .A1(n13781), .A2(n13742), .ZN(n13743) );
  OAI21_X1 U15272 ( .B1(n13781), .B2(n13744), .A(n13743), .ZN(n13784) );
  XOR2_X1 U15273 ( .A(n13797), .B(n14141), .Z(n14018) );
  NAND4_X1 U15274 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13752) );
  NOR4_X1 U15275 ( .A1(n13752), .A2(n13751), .A3(n13750), .A4(n13749), .ZN(
        n13755) );
  NAND4_X1 U15276 ( .A1(n13756), .A2(n13755), .A3(n13754), .A4(n13753), .ZN(
        n13757) );
  NOR4_X1 U15277 ( .A1(n13760), .A2(n13759), .A3(n13758), .A4(n13757), .ZN(
        n13763) );
  NAND4_X1 U15278 ( .A1(n13764), .A2(n13763), .A3(n13762), .A4(n13761), .ZN(
        n13765) );
  NOR3_X1 U15279 ( .A1(n13767), .A2(n13766), .A3(n13765), .ZN(n13769) );
  NAND4_X1 U15280 ( .A1(n14054), .A2(n13769), .A3(n13768), .A4(n14084), .ZN(
        n13770) );
  NOR4_X1 U15281 ( .A1(n13971), .A2(n14018), .A3(n14028), .A4(n13770), .ZN(
        n13771) );
  NAND4_X1 U15282 ( .A1(n13771), .A2(n13966), .A3(n13990), .A4(n14006), .ZN(
        n13772) );
  NOR4_X1 U15283 ( .A1(n13900), .A2(n13913), .A3(n13933), .A4(n13772), .ZN(
        n13775) );
  XNOR2_X1 U15284 ( .A(n13883), .B(n13788), .ZN(n13773) );
  NAND4_X1 U15285 ( .A1(n13718), .A2(n13775), .A3(n13774), .A4(n13773), .ZN(
        n13777) );
  XNOR2_X1 U15286 ( .A(n13777), .B(n13776), .ZN(n13778) );
  AOI211_X1 U15287 ( .C1(n13781), .C2(n13780), .A(n13779), .B(n13778), .ZN(
        n13783) );
  OAI21_X1 U15288 ( .B1(n13784), .B2(n13783), .A(n13782), .ZN(n13785) );
  OAI21_X1 U15289 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(P2_U3328) );
  MUX2_X1 U15290 ( .A(n13884), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13812), .Z(
        P2_U3562) );
  MUX2_X1 U15291 ( .A(n13788), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13812), .Z(
        P2_U3561) );
  MUX2_X1 U15292 ( .A(n13789), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13812), .Z(
        P2_U3560) );
  MUX2_X1 U15293 ( .A(n13790), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13812), .Z(
        P2_U3559) );
  MUX2_X1 U15294 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13791), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15295 ( .A(n13792), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13812), .Z(
        P2_U3557) );
  MUX2_X1 U15296 ( .A(n13793), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13812), .Z(
        P2_U3556) );
  MUX2_X1 U15297 ( .A(n13794), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13812), .Z(
        P2_U3555) );
  MUX2_X1 U15298 ( .A(n13795), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13812), .Z(
        P2_U3554) );
  MUX2_X1 U15299 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13796), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15300 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13797), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15301 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13798), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15302 ( .A(n14072), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13812), .Z(
        P2_U3550) );
  MUX2_X1 U15303 ( .A(n13799), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13812), .Z(
        P2_U3549) );
  MUX2_X1 U15304 ( .A(n14070), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13812), .Z(
        P2_U3548) );
  MUX2_X1 U15305 ( .A(n13800), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13812), .Z(
        P2_U3547) );
  MUX2_X1 U15306 ( .A(n13801), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13812), .Z(
        P2_U3546) );
  MUX2_X1 U15307 ( .A(n13802), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13812), .Z(
        P2_U3545) );
  MUX2_X1 U15308 ( .A(n13803), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13812), .Z(
        P2_U3544) );
  MUX2_X1 U15309 ( .A(n13804), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13812), .Z(
        P2_U3543) );
  MUX2_X1 U15310 ( .A(n13805), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13812), .Z(
        P2_U3542) );
  MUX2_X1 U15311 ( .A(n13806), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13812), .Z(
        P2_U3541) );
  MUX2_X1 U15312 ( .A(n13807), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13812), .Z(
        P2_U3540) );
  MUX2_X1 U15313 ( .A(n13808), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13812), .Z(
        P2_U3539) );
  MUX2_X1 U15314 ( .A(n13809), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13812), .Z(
        P2_U3538) );
  MUX2_X1 U15315 ( .A(n13810), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13812), .Z(
        P2_U3537) );
  MUX2_X1 U15316 ( .A(n13811), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13812), .Z(
        P2_U3536) );
  MUX2_X1 U15317 ( .A(n13813), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13812), .Z(
        P2_U3535) );
  MUX2_X1 U15318 ( .A(n13814), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13812), .Z(
        P2_U3534) );
  MUX2_X1 U15319 ( .A(n13815), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13812), .Z(
        P2_U3533) );
  MUX2_X1 U15320 ( .A(n13816), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13812), .Z(
        P2_U3532) );
  MUX2_X1 U15321 ( .A(n13528), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13812), .Z(
        P2_U3531) );
  INV_X1 U15322 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n13817) );
  OAI22_X1 U15323 ( .A1(n15198), .A2(n13817), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8284), .ZN(n13818) );
  AOI21_X1 U15324 ( .B1(n13824), .B2(n15210), .A(n13818), .ZN(n13832) );
  INV_X1 U15325 ( .A(n13819), .ZN(n13839) );
  NAND3_X1 U15326 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n13823) );
  NAND3_X1 U15327 ( .A1(n15205), .A2(n13839), .A3(n13823), .ZN(n13831) );
  MUX2_X1 U15328 ( .A(n10588), .B(P2_REG1_REG_2__SCAN_IN), .S(n13824), .Z(
        n13827) );
  INV_X1 U15329 ( .A(n13825), .ZN(n13826) );
  NAND2_X1 U15330 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  OAI211_X1 U15331 ( .C1(n13829), .C2(n13828), .A(n15201), .B(n13845), .ZN(
        n13830) );
  NAND3_X1 U15332 ( .A1(n13832), .A2(n13831), .A3(n13830), .ZN(P2_U3216) );
  OAI22_X1 U15333 ( .A1(n15198), .A2(n7385), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13833), .ZN(n13834) );
  AOI21_X1 U15334 ( .B1(n13836), .B2(n15210), .A(n13834), .ZN(n13850) );
  INV_X1 U15335 ( .A(n13835), .ZN(n13838) );
  MUX2_X1 U15336 ( .A(n11349), .B(P2_REG2_REG_3__SCAN_IN), .S(n13836), .Z(
        n13837) );
  NAND3_X1 U15337 ( .A1(n13839), .A2(n13838), .A3(n13837), .ZN(n13840) );
  NAND3_X1 U15338 ( .A1(n15205), .A2(n13841), .A3(n13840), .ZN(n13849) );
  INV_X1 U15339 ( .A(n13842), .ZN(n13847) );
  NAND3_X1 U15340 ( .A1(n13845), .A2(n13844), .A3(n13843), .ZN(n13846) );
  NAND3_X1 U15341 ( .A1(n15201), .A2(n13847), .A3(n13846), .ZN(n13848) );
  NAND3_X1 U15342 ( .A1(n13850), .A2(n13849), .A3(n13848), .ZN(P2_U3217) );
  OAI21_X1 U15343 ( .B1(n13853), .B2(n13852), .A(n13851), .ZN(n13854) );
  NAND2_X1 U15344 ( .A1(n13854), .A2(n15205), .ZN(n13864) );
  AND2_X1 U15345 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n13855) );
  AOI21_X1 U15346 ( .B1(n15200), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n13855), .ZN(
        n13863) );
  OAI21_X1 U15347 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13859) );
  NAND2_X1 U15348 ( .A1(n13859), .A2(n15201), .ZN(n13862) );
  NAND2_X1 U15349 ( .A1(n15210), .A2(n13860), .ZN(n13861) );
  NAND4_X1 U15350 ( .A1(n13864), .A2(n13863), .A3(n13862), .A4(n13861), .ZN(
        P2_U3223) );
  OAI21_X1 U15351 ( .B1(n13867), .B2(n13866), .A(n13865), .ZN(n13868) );
  NAND2_X1 U15352 ( .A1(n13868), .A2(n15205), .ZN(n13882) );
  INV_X1 U15353 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n13870) );
  OAI21_X1 U15354 ( .B1(n15198), .B2(n13870), .A(n13869), .ZN(n13871) );
  AOI21_X1 U15355 ( .B1(n13873), .B2(n15210), .A(n13871), .ZN(n13881) );
  INV_X1 U15356 ( .A(n13872), .ZN(n13876) );
  MUX2_X1 U15357 ( .A(n13874), .B(P2_REG1_REG_11__SCAN_IN), .S(n13873), .Z(
        n13875) );
  NAND2_X1 U15358 ( .A1(n13876), .A2(n13875), .ZN(n13878) );
  OAI211_X1 U15359 ( .C1(n13879), .C2(n13878), .A(n13877), .B(n15201), .ZN(
        n13880) );
  NAND3_X1 U15360 ( .A1(n13882), .A2(n13881), .A3(n13880), .ZN(P2_U3225) );
  NAND2_X1 U15361 ( .A1(n14180), .A2(n13889), .ZN(n13888) );
  NAND2_X1 U15362 ( .A1(n13885), .A2(n13884), .ZN(n14091) );
  NOR2_X1 U15363 ( .A1(n13980), .A2(n14091), .ZN(n13891) );
  NOR2_X1 U15364 ( .A1(n7382), .A2(n15821), .ZN(n13886) );
  AOI211_X1 U15365 ( .C1(n15818), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13891), 
        .B(n13886), .ZN(n13887) );
  OAI21_X1 U15366 ( .B1(n13984), .B2(n14089), .A(n13887), .ZN(P2_U3234) );
  OAI211_X1 U15367 ( .C1(n14180), .C2(n13889), .A(n13976), .B(n13888), .ZN(
        n14092) );
  NOR2_X1 U15368 ( .A1(n14180), .A2(n15821), .ZN(n13890) );
  AOI211_X1 U15369 ( .C1(n15818), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13891), 
        .B(n13890), .ZN(n13892) );
  OAI21_X1 U15370 ( .B1(n13984), .B2(n14092), .A(n13892), .ZN(P2_U3235) );
  XNOR2_X1 U15371 ( .A(n13893), .B(n8826), .ZN(n14100) );
  OAI21_X1 U15372 ( .B1(n13921), .B2(n14183), .A(n13976), .ZN(n13894) );
  INV_X1 U15373 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13896) );
  OAI22_X1 U15374 ( .A1(n13897), .A2(n13959), .B1(n13896), .B2(n7197), .ZN(
        n13898) );
  AOI21_X1 U15375 ( .B1(n14104), .B2(n14035), .A(n13898), .ZN(n13899) );
  OAI21_X1 U15376 ( .B1(n14101), .B2(n13984), .A(n13899), .ZN(n13908) );
  NAND2_X1 U15377 ( .A1(n13901), .A2(n13900), .ZN(n13902) );
  NAND3_X1 U15378 ( .A1(n13903), .A2(n13902), .A3(n14074), .ZN(n13906) );
  INV_X1 U15379 ( .A(n13904), .ZN(n13905) );
  NOR2_X1 U15380 ( .A1(n14102), .A2(n13980), .ZN(n13907) );
  AOI211_X1 U15381 ( .C1(n14100), .C2(n15824), .A(n13908), .B(n13907), .ZN(
        n13909) );
  INV_X1 U15382 ( .A(n13909), .ZN(P2_U3237) );
  INV_X1 U15383 ( .A(n13910), .ZN(n13911) );
  AOI21_X1 U15384 ( .B1(n13913), .B2(n13912), .A(n13911), .ZN(n13916) );
  INV_X1 U15385 ( .A(n13914), .ZN(n13915) );
  OAI21_X1 U15386 ( .B1(n13916), .B2(n14063), .A(n13915), .ZN(n14105) );
  INV_X1 U15387 ( .A(n14105), .ZN(n13929) );
  INV_X1 U15388 ( .A(n13917), .ZN(n13918) );
  AOI21_X1 U15389 ( .B1(n13920), .B2(n13919), .A(n13918), .ZN(n14107) );
  INV_X1 U15390 ( .A(n13940), .ZN(n13922) );
  AOI211_X1 U15391 ( .C1(n13923), .C2(n13922), .A(n14076), .B(n13921), .ZN(
        n14106) );
  NAND2_X1 U15392 ( .A1(n14106), .A2(n15814), .ZN(n13926) );
  AOI22_X1 U15393 ( .A1(n13924), .A2(n15816), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13980), .ZN(n13925) );
  OAI211_X1 U15394 ( .C1(n14187), .C2(n15821), .A(n13926), .B(n13925), .ZN(
        n13927) );
  AOI21_X1 U15395 ( .B1(n14107), .B2(n15824), .A(n13927), .ZN(n13928) );
  OAI21_X1 U15396 ( .B1(n13929), .B2(n13980), .A(n13928), .ZN(P2_U3238) );
  XNOR2_X1 U15397 ( .A(n13931), .B(n13930), .ZN(n14113) );
  INV_X1 U15398 ( .A(n14113), .ZN(n13948) );
  NAND3_X1 U15399 ( .A1(n13953), .A2(n13933), .A3(n13932), .ZN(n13934) );
  NAND3_X1 U15400 ( .A1(n13935), .A2(n14074), .A3(n13934), .ZN(n13938) );
  INV_X1 U15401 ( .A(n13936), .ZN(n13937) );
  NAND2_X1 U15402 ( .A1(n13938), .A2(n13937), .ZN(n14111) );
  OAI21_X1 U15403 ( .B1(n13962), .B2(n14191), .A(n13976), .ZN(n13939) );
  OR2_X1 U15404 ( .A1(n13940), .A2(n13939), .ZN(n14110) );
  INV_X1 U15405 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13941) );
  OAI22_X1 U15406 ( .A1(n13942), .A2(n13959), .B1(n13941), .B2(n7197), .ZN(
        n13943) );
  AOI21_X1 U15407 ( .B1(n13944), .B2(n14035), .A(n13943), .ZN(n13945) );
  OAI21_X1 U15408 ( .B1(n14110), .B2(n13984), .A(n13945), .ZN(n13946) );
  AOI21_X1 U15409 ( .B1(n14111), .B2(n7197), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15410 ( .B1(n13948), .B2(n14085), .A(n13947), .ZN(P2_U3239) );
  NAND2_X1 U15411 ( .A1(n13949), .A2(n13950), .ZN(n13952) );
  NAND2_X1 U15412 ( .A1(n13952), .A2(n13951), .ZN(n13954) );
  NAND3_X1 U15413 ( .A1(n13954), .A2(n14074), .A3(n13953), .ZN(n13957) );
  INV_X1 U15414 ( .A(n13955), .ZN(n13956) );
  AND2_X1 U15415 ( .A1(n13957), .A2(n13956), .ZN(n14119) );
  INV_X1 U15416 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13958) );
  OAI22_X1 U15417 ( .A1(n13960), .A2(n13959), .B1(n13958), .B2(n7197), .ZN(
        n13964) );
  OAI21_X1 U15418 ( .B1(n13978), .B2(n14195), .A(n13976), .ZN(n13961) );
  OR2_X1 U15419 ( .A1(n13962), .A2(n13961), .ZN(n14117) );
  NOR2_X1 U15420 ( .A1(n14117), .A2(n13984), .ZN(n13963) );
  AOI211_X1 U15421 ( .C1(n14035), .C2(n13965), .A(n13964), .B(n13963), .ZN(
        n13969) );
  XNOR2_X1 U15422 ( .A(n13967), .B(n13966), .ZN(n14116) );
  NAND2_X1 U15423 ( .A1(n14116), .A2(n15824), .ZN(n13968) );
  OAI211_X1 U15424 ( .C1(n15818), .C2(n14119), .A(n13969), .B(n13968), .ZN(
        P2_U3240) );
  XNOR2_X1 U15425 ( .A(n13970), .B(n13971), .ZN(n14124) );
  NAND2_X1 U15426 ( .A1(n13972), .A2(n13971), .ZN(n13973) );
  NAND2_X1 U15427 ( .A1(n13949), .A2(n13973), .ZN(n13975) );
  AOI21_X1 U15428 ( .B1(n13975), .B2(n14074), .A(n13974), .ZN(n14123) );
  INV_X1 U15429 ( .A(n14123), .ZN(n13986) );
  NAND2_X1 U15430 ( .A1(n13996), .A2(n14126), .ZN(n13977) );
  NAND2_X1 U15431 ( .A1(n13977), .A2(n13976), .ZN(n13979) );
  OR2_X1 U15432 ( .A1(n13979), .A2(n13978), .ZN(n14122) );
  AOI22_X1 U15433 ( .A1(n13981), .A2(n15816), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13980), .ZN(n13983) );
  NAND2_X1 U15434 ( .A1(n14126), .A2(n14035), .ZN(n13982) );
  OAI211_X1 U15435 ( .C1(n14122), .C2(n13984), .A(n13983), .B(n13982), .ZN(
        n13985) );
  AOI21_X1 U15436 ( .B1(n13986), .B2(n7197), .A(n13985), .ZN(n13987) );
  OAI21_X1 U15437 ( .B1(n14085), .B2(n14124), .A(n13987), .ZN(P2_U3241) );
  XNOR2_X1 U15438 ( .A(n13988), .B(n13990), .ZN(n14131) );
  INV_X1 U15439 ( .A(n14131), .ZN(n14002) );
  OAI211_X1 U15440 ( .C1(n13991), .C2(n13990), .A(n13989), .B(n14074), .ZN(
        n13993) );
  NAND2_X1 U15441 ( .A1(n13993), .A2(n13992), .ZN(n14129) );
  AOI21_X1 U15442 ( .B1(n14008), .B2(n13994), .A(n14076), .ZN(n13995) );
  AND2_X1 U15443 ( .A1(n13996), .A2(n13995), .ZN(n14130) );
  NAND2_X1 U15444 ( .A1(n14130), .A2(n15814), .ZN(n13999) );
  AOI22_X1 U15445 ( .A1(n13997), .A2(n15816), .B1(n15818), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13998) );
  OAI211_X1 U15446 ( .C1(n14204), .C2(n15821), .A(n13999), .B(n13998), .ZN(
        n14000) );
  AOI21_X1 U15447 ( .B1(n14129), .B2(n7197), .A(n14000), .ZN(n14001) );
  OAI21_X1 U15448 ( .B1(n14085), .B2(n14002), .A(n14001), .ZN(P2_U3242) );
  XNOR2_X1 U15449 ( .A(n14003), .B(n14006), .ZN(n14005) );
  OAI21_X1 U15450 ( .B1(n14005), .B2(n14063), .A(n14004), .ZN(n14135) );
  INV_X1 U15451 ( .A(n14135), .ZN(n14016) );
  XOR2_X1 U15452 ( .A(n14007), .B(n14006), .Z(n14136) );
  INV_X1 U15453 ( .A(n14008), .ZN(n14009) );
  AOI211_X1 U15454 ( .C1(n14010), .C2(n14021), .A(n14076), .B(n14009), .ZN(
        n14134) );
  NAND2_X1 U15455 ( .A1(n14134), .A2(n15814), .ZN(n14013) );
  AOI22_X1 U15456 ( .A1(n15818), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14011), 
        .B2(n15816), .ZN(n14012) );
  OAI211_X1 U15457 ( .C1(n7586), .C2(n15821), .A(n14013), .B(n14012), .ZN(
        n14014) );
  AOI21_X1 U15458 ( .B1(n15824), .B2(n14136), .A(n14014), .ZN(n14015) );
  OAI21_X1 U15459 ( .B1(n15818), .B2(n14016), .A(n14015), .ZN(P2_U3243) );
  XOR2_X1 U15460 ( .A(n14018), .B(n14017), .Z(n14143) );
  XNOR2_X1 U15461 ( .A(n7249), .B(n14018), .ZN(n14020) );
  OAI21_X1 U15462 ( .B1(n14020), .B2(n14063), .A(n14019), .ZN(n14139) );
  NAND2_X1 U15463 ( .A1(n14139), .A2(n7197), .ZN(n14026) );
  AOI211_X1 U15464 ( .C1(n14141), .C2(n14033), .A(n14076), .B(n7196), .ZN(
        n14140) );
  AOI22_X1 U15465 ( .A1(n15818), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14022), 
        .B2(n15816), .ZN(n14023) );
  OAI21_X1 U15466 ( .B1(n7587), .B2(n15821), .A(n14023), .ZN(n14024) );
  AOI21_X1 U15467 ( .B1(n14140), .B2(n15814), .A(n14024), .ZN(n14025) );
  OAI211_X1 U15468 ( .C1(n14143), .C2(n14085), .A(n14026), .B(n14025), .ZN(
        P2_U3244) );
  XOR2_X1 U15469 ( .A(n14027), .B(n14028), .Z(n14148) );
  XNOR2_X1 U15470 ( .A(n14029), .B(n14028), .ZN(n14030) );
  OAI222_X1 U15471 ( .A1(n14057), .A2(n14032), .B1(n14055), .B2(n14031), .C1(
        n14030), .C2(n14063), .ZN(n14144) );
  NAND2_X1 U15472 ( .A1(n14144), .A2(n7197), .ZN(n14041) );
  AOI21_X1 U15473 ( .B1(n14146), .B2(n14045), .A(n14076), .ZN(n14034) );
  AND2_X1 U15474 ( .A1(n14034), .A2(n14033), .ZN(n14145) );
  NAND2_X1 U15475 ( .A1(n14146), .A2(n14035), .ZN(n14038) );
  AOI22_X1 U15476 ( .A1(n15818), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14036), 
        .B2(n15816), .ZN(n14037) );
  NAND2_X1 U15477 ( .A1(n14038), .A2(n14037), .ZN(n14039) );
  AOI21_X1 U15478 ( .B1(n14145), .B2(n15814), .A(n14039), .ZN(n14040) );
  OAI211_X1 U15479 ( .C1(n14148), .C2(n14085), .A(n14041), .B(n14040), .ZN(
        P2_U3245) );
  OAI21_X1 U15480 ( .B1(n14044), .B2(n14043), .A(n14042), .ZN(n14151) );
  INV_X1 U15481 ( .A(n14151), .ZN(n14067) );
  INV_X1 U15482 ( .A(n14075), .ZN(n14047) );
  INV_X1 U15483 ( .A(n14045), .ZN(n14046) );
  AOI211_X1 U15484 ( .C1(n14048), .C2(n14047), .A(n14076), .B(n14046), .ZN(
        n14150) );
  INV_X1 U15485 ( .A(n14049), .ZN(n14050) );
  AOI22_X1 U15486 ( .A1(n15818), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14050), 
        .B2(n15816), .ZN(n14051) );
  OAI21_X1 U15487 ( .B1(n14213), .B2(n15821), .A(n14051), .ZN(n14052) );
  AOI21_X1 U15488 ( .B1(n14150), .B2(n15814), .A(n14052), .ZN(n14065) );
  XNOR2_X1 U15489 ( .A(n14054), .B(n14053), .ZN(n14062) );
  OAI22_X1 U15490 ( .A1(n14058), .A2(n14057), .B1(n14056), .B2(n14055), .ZN(
        n14059) );
  AOI21_X1 U15491 ( .B1(n14151), .B2(n14060), .A(n14059), .ZN(n14061) );
  OAI21_X1 U15492 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(n14149) );
  NAND2_X1 U15493 ( .A1(n14149), .A2(n7197), .ZN(n14064) );
  OAI211_X1 U15494 ( .C1(n14067), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        P2_U3246) );
  XOR2_X1 U15495 ( .A(n14068), .B(n14084), .Z(n14073) );
  AOI222_X1 U15496 ( .A1(n14074), .A2(n14073), .B1(n14072), .B2(n14071), .C1(
        n14070), .C2(n14069), .ZN(n14157) );
  AOI211_X1 U15497 ( .C1(n14155), .C2(n14077), .A(n14076), .B(n14075), .ZN(
        n14154) );
  AOI22_X1 U15498 ( .A1(n15818), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14078), 
        .B2(n15816), .ZN(n14079) );
  OAI21_X1 U15499 ( .B1(n14080), .B2(n15821), .A(n14079), .ZN(n14087) );
  INV_X1 U15500 ( .A(n14081), .ZN(n14082) );
  AOI21_X1 U15501 ( .B1(n14084), .B2(n14083), .A(n14082), .ZN(n14158) );
  NOR2_X1 U15502 ( .A1(n14158), .A2(n14085), .ZN(n14086) );
  AOI211_X1 U15503 ( .C1(n14154), .C2(n15814), .A(n14087), .B(n14086), .ZN(
        n14088) );
  OAI21_X1 U15504 ( .B1(n15818), .B2(n14157), .A(n14088), .ZN(P2_U3247) );
  INV_X1 U15505 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14093) );
  AND2_X1 U15506 ( .A1(n14092), .A2(n14091), .ZN(n14177) );
  MUX2_X1 U15507 ( .A(n14093), .B(n14177), .S(n15869), .Z(n14094) );
  OAI21_X1 U15508 ( .B1(n14180), .B2(n14165), .A(n14094), .ZN(P2_U3529) );
  AOI21_X1 U15509 ( .B1(n15861), .B2(n14096), .A(n14095), .ZN(n14097) );
  OAI211_X1 U15510 ( .C1(n14159), .C2(n14099), .A(n14098), .B(n14097), .ZN(
        n14181) );
  MUX2_X1 U15511 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14181), .S(n15869), .Z(
        P2_U3528) );
  NAND2_X1 U15512 ( .A1(n14100), .A2(n15859), .ZN(n14103) );
  INV_X1 U15513 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14108) );
  MUX2_X1 U15514 ( .A(n14108), .B(n14184), .S(n15869), .Z(n14109) );
  OAI21_X1 U15515 ( .B1(n14187), .B2(n14165), .A(n14109), .ZN(P2_U3526) );
  INV_X1 U15516 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14114) );
  INV_X1 U15517 ( .A(n14110), .ZN(n14112) );
  AOI211_X1 U15518 ( .C1(n15859), .C2(n14113), .A(n14112), .B(n14111), .ZN(
        n14188) );
  MUX2_X1 U15519 ( .A(n14114), .B(n14188), .S(n15869), .Z(n14115) );
  OAI21_X1 U15520 ( .B1(n14191), .B2(n14165), .A(n14115), .ZN(P2_U3525) );
  INV_X1 U15521 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U15522 ( .A1(n14116), .A2(n15859), .ZN(n14118) );
  MUX2_X1 U15523 ( .A(n14120), .B(n14192), .S(n15869), .Z(n14121) );
  OAI21_X1 U15524 ( .B1(n14195), .B2(n14165), .A(n14121), .ZN(P2_U3524) );
  OAI211_X1 U15525 ( .C1(n14159), .C2(n14124), .A(n14123), .B(n14122), .ZN(
        n14196) );
  MUX2_X1 U15526 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14196), .S(n15869), .Z(
        n14125) );
  AOI21_X1 U15527 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n14128) );
  INV_X1 U15528 ( .A(n14128), .ZN(P2_U3523) );
  INV_X1 U15529 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14132) );
  AOI211_X1 U15530 ( .C1(n15859), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        n14201) );
  MUX2_X1 U15531 ( .A(n14132), .B(n14201), .S(n15869), .Z(n14133) );
  OAI21_X1 U15532 ( .B1(n14204), .B2(n14165), .A(n14133), .ZN(P2_U3522) );
  INV_X1 U15533 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14137) );
  AOI211_X1 U15534 ( .C1(n15859), .C2(n14136), .A(n14135), .B(n14134), .ZN(
        n14205) );
  MUX2_X1 U15535 ( .A(n14137), .B(n14205), .S(n15869), .Z(n14138) );
  OAI21_X1 U15536 ( .B1(n7586), .B2(n14165), .A(n14138), .ZN(P2_U3521) );
  AOI211_X1 U15537 ( .C1(n15861), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14142) );
  OAI21_X1 U15538 ( .B1(n14159), .B2(n14143), .A(n14142), .ZN(n14208) );
  MUX2_X1 U15539 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14208), .S(n15869), .Z(
        P2_U3520) );
  AOI211_X1 U15540 ( .C1(n15861), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14147) );
  OAI21_X1 U15541 ( .B1(n14159), .B2(n14148), .A(n14147), .ZN(n14209) );
  MUX2_X1 U15542 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14209), .S(n15869), .Z(
        P2_U3519) );
  MUX2_X1 U15543 ( .A(n14152), .B(n14210), .S(n15869), .Z(n14153) );
  OAI21_X1 U15544 ( .B1(n14213), .B2(n14165), .A(n14153), .ZN(P2_U3518) );
  AOI21_X1 U15545 ( .B1(n15861), .B2(n14155), .A(n14154), .ZN(n14156) );
  OAI211_X1 U15546 ( .C1(n14159), .C2(n14158), .A(n14157), .B(n14156), .ZN(
        n14214) );
  MUX2_X1 U15547 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14214), .S(n15869), .Z(
        P2_U3517) );
  AOI211_X1 U15548 ( .C1(n15859), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        n14216) );
  MUX2_X1 U15549 ( .A(n14163), .B(n14216), .S(n15869), .Z(n14164) );
  OAI21_X1 U15550 ( .B1(n14220), .B2(n14165), .A(n14164), .ZN(P2_U3516) );
  INV_X1 U15551 ( .A(n14166), .ZN(n14170) );
  INV_X1 U15552 ( .A(n15861), .ZN(n15753) );
  OAI21_X1 U15553 ( .B1(n14168), .B2(n15753), .A(n14167), .ZN(n14169) );
  AOI21_X1 U15554 ( .B1(n14170), .B2(n15758), .A(n14169), .ZN(n14171) );
  NAND2_X1 U15555 ( .A1(n14172), .A2(n14171), .ZN(n14221) );
  MUX2_X1 U15556 ( .A(n14221), .B(P2_REG1_REG_16__SCAN_IN), .S(n15868), .Z(
        P2_U3515) );
  INV_X1 U15557 ( .A(n14173), .ZN(n14174) );
  MUX2_X1 U15558 ( .A(n14175), .B(n14174), .S(n14215), .Z(n14176) );
  OAI21_X1 U15559 ( .B1(n7382), .B2(n14219), .A(n14176), .ZN(P2_U3498) );
  MUX2_X1 U15560 ( .A(n14178), .B(n14177), .S(n14215), .Z(n14179) );
  OAI21_X1 U15561 ( .B1(n14180), .B2(n14219), .A(n14179), .ZN(P2_U3497) );
  MUX2_X1 U15562 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14181), .S(n14215), .Z(
        P2_U3496) );
  MUX2_X1 U15563 ( .A(n14185), .B(n14184), .S(n14215), .Z(n14186) );
  OAI21_X1 U15564 ( .B1(n14187), .B2(n14219), .A(n14186), .ZN(P2_U3494) );
  MUX2_X1 U15565 ( .A(n14189), .B(n14188), .S(n14215), .Z(n14190) );
  OAI21_X1 U15566 ( .B1(n14191), .B2(n14219), .A(n14190), .ZN(P2_U3493) );
  MUX2_X1 U15567 ( .A(n14193), .B(n14192), .S(n14215), .Z(n14194) );
  OAI21_X1 U15568 ( .B1(n14195), .B2(n14219), .A(n14194), .ZN(P2_U3492) );
  INV_X1 U15569 ( .A(n14196), .ZN(n14197) );
  MUX2_X1 U15570 ( .A(n14198), .B(n14197), .S(n14215), .Z(n14199) );
  OAI21_X1 U15571 ( .B1(n14200), .B2(n14219), .A(n14199), .ZN(P2_U3491) );
  MUX2_X1 U15572 ( .A(n14202), .B(n14201), .S(n14215), .Z(n14203) );
  OAI21_X1 U15573 ( .B1(n14204), .B2(n14219), .A(n14203), .ZN(P2_U3490) );
  MUX2_X1 U15574 ( .A(n14206), .B(n14205), .S(n14215), .Z(n14207) );
  OAI21_X1 U15575 ( .B1(n7586), .B2(n14219), .A(n14207), .ZN(P2_U3489) );
  MUX2_X1 U15576 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14208), .S(n14215), .Z(
        P2_U3488) );
  MUX2_X1 U15577 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14209), .S(n14215), .Z(
        P2_U3487) );
  INV_X1 U15578 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14211) );
  MUX2_X1 U15579 ( .A(n14211), .B(n14210), .S(n14215), .Z(n14212) );
  OAI21_X1 U15580 ( .B1(n14213), .B2(n14219), .A(n14212), .ZN(P2_U3486) );
  MUX2_X1 U15581 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14214), .S(n14215), .Z(
        P2_U3484) );
  INV_X1 U15582 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14217) );
  MUX2_X1 U15583 ( .A(n14217), .B(n14216), .S(n14215), .Z(n14218) );
  OAI21_X1 U15584 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(P2_U3481) );
  MUX2_X1 U15585 ( .A(n14221), .B(P2_REG0_REG_16__SCAN_IN), .S(n15870), .Z(
        P2_U3478) );
  INV_X1 U15586 ( .A(n13683), .ZN(n14877) );
  NOR4_X1 U15587 ( .A1(n8250), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8756), .A4(
        P2_U3088), .ZN(n14222) );
  AOI21_X1 U15588 ( .B1(n14234), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14222), 
        .ZN(n14223) );
  OAI21_X1 U15589 ( .B1(n14877), .B2(n14239), .A(n14223), .ZN(P2_U3296) );
  INV_X1 U15590 ( .A(n14224), .ZN(n14883) );
  OAI222_X1 U15591 ( .A1(n14239), .A2(n14883), .B1(P2_U3088), .B2(n14226), 
        .C1(n14225), .C2(n14244), .ZN(P2_U3298) );
  INV_X1 U15592 ( .A(n14227), .ZN(n14884) );
  AOI21_X1 U15593 ( .B1(n14234), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14228), 
        .ZN(n14229) );
  OAI21_X1 U15594 ( .B1(n14884), .B2(n14239), .A(n14229), .ZN(P2_U3299) );
  INV_X1 U15595 ( .A(n14230), .ZN(n14887) );
  OAI222_X1 U15596 ( .A1(n14244), .A2(n14232), .B1(n14239), .B2(n14887), .C1(
        n14231), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15597 ( .A(n14233), .ZN(n14890) );
  AOI22_X1 U15598 ( .A1(n14235), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14234), .ZN(n14236) );
  OAI21_X1 U15599 ( .B1(n14890), .B2(n14239), .A(n14236), .ZN(P2_U3301) );
  INV_X1 U15600 ( .A(n14237), .ZN(n14892) );
  OAI222_X1 U15601 ( .A1(n14244), .A2(n14240), .B1(n14239), .B2(n14892), .C1(
        n14238), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15602 ( .A(n14241), .ZN(n14896) );
  OAI222_X1 U15603 ( .A1(n14244), .A2(n14243), .B1(n14239), .B2(n14896), .C1(
        n14242), .C2(P2_U3088), .ZN(P2_U3303) );
  MUX2_X1 U15604 ( .A(n14245), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15605 ( .B1(n14248), .B2(n14247), .A(n14246), .ZN(n14249) );
  NAND2_X1 U15606 ( .A1(n14249), .A2(n15963), .ZN(n14253) );
  AOI22_X1 U15607 ( .A1(n14357), .A2(n14767), .B1(n14765), .B2(n14586), .ZN(
        n14595) );
  OAI22_X1 U15608 ( .A1(n14595), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14250), .ZN(n14251) );
  AOI21_X1 U15609 ( .B1(n14603), .B2(n14352), .A(n14251), .ZN(n14252) );
  OAI211_X1 U15610 ( .C1(n14804), .C2(n14348), .A(n14253), .B(n14252), .ZN(
        P1_U3214) );
  AOI21_X1 U15611 ( .B1(n14255), .B2(n14254), .A(n7327), .ZN(n14263) );
  NAND2_X1 U15612 ( .A1(n14345), .A2(n14363), .ZN(n14257) );
  OAI211_X1 U15613 ( .C1(n15942), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14260) );
  NOR2_X1 U15614 ( .A1(n15850), .A2(n14348), .ZN(n14259) );
  AOI211_X1 U15615 ( .C1(n14352), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        n14262) );
  OAI21_X1 U15616 ( .B1(n14263), .B2(n15949), .A(n14262), .ZN(P1_U3215) );
  INV_X1 U15617 ( .A(n14264), .ZN(n14265) );
  AOI21_X1 U15618 ( .B1(n14267), .B2(n14266), .A(n14265), .ZN(n14273) );
  AOI22_X1 U15619 ( .A1(n14316), .A2(n14663), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14269) );
  NAND2_X1 U15620 ( .A1(n14352), .A2(n14664), .ZN(n14268) );
  OAI211_X1 U15621 ( .C1(n14270), .C2(n15945), .A(n14269), .B(n14268), .ZN(
        n14271) );
  AOI21_X1 U15622 ( .B1(n14670), .B2(n15965), .A(n14271), .ZN(n14272) );
  OAI21_X1 U15623 ( .B1(n14273), .B2(n15949), .A(n14272), .ZN(P1_U3216) );
  INV_X1 U15624 ( .A(n14274), .ZN(n14275) );
  AOI21_X1 U15625 ( .B1(n14277), .B2(n14276), .A(n14275), .ZN(n14283) );
  AND2_X1 U15626 ( .A1(n14662), .A2(n14765), .ZN(n14278) );
  AOI21_X1 U15627 ( .B1(n14730), .B2(n14767), .A(n14278), .ZN(n14697) );
  INV_X1 U15628 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14279) );
  OAI22_X1 U15629 ( .A1(n14697), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14279), .ZN(n14281) );
  NOR2_X1 U15630 ( .A1(n12438), .A2(n14348), .ZN(n14280) );
  AOI211_X1 U15631 ( .C1(n14352), .C2(n14705), .A(n14281), .B(n14280), .ZN(
        n14282) );
  OAI21_X1 U15632 ( .B1(n14283), .B2(n15949), .A(n14282), .ZN(P1_U3223) );
  XOR2_X1 U15633 ( .A(n14285), .B(n14284), .Z(n14292) );
  NAND2_X1 U15634 ( .A1(n14663), .A2(n14767), .ZN(n14287) );
  NAND2_X1 U15635 ( .A1(n14357), .A2(n14765), .ZN(n14286) );
  AND2_X1 U15636 ( .A1(n14287), .A2(n14286), .ZN(n14634) );
  OAI22_X1 U15637 ( .A1(n14634), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14288), .ZN(n14290) );
  NOR2_X1 U15638 ( .A1(n14638), .A2(n14348), .ZN(n14289) );
  AOI211_X1 U15639 ( .C1(n14352), .C2(n14635), .A(n14290), .B(n14289), .ZN(
        n14291) );
  OAI21_X1 U15640 ( .B1(n14292), .B2(n15949), .A(n14291), .ZN(P1_U3225) );
  OAI21_X1 U15641 ( .B1(n14295), .B2(n14294), .A(n14293), .ZN(n14296) );
  NAND2_X1 U15642 ( .A1(n14296), .A2(n15963), .ZN(n14301) );
  NAND2_X1 U15643 ( .A1(n14345), .A2(n14768), .ZN(n14298) );
  OAI211_X1 U15644 ( .C1(n15942), .C2(n15944), .A(n14298), .B(n14297), .ZN(
        n14299) );
  AOI21_X1 U15645 ( .B1(n14771), .B2(n14352), .A(n14299), .ZN(n14300) );
  OAI211_X1 U15646 ( .C1(n14775), .C2(n14348), .A(n14301), .B(n14300), .ZN(
        P1_U3226) );
  OAI21_X1 U15647 ( .B1(n14304), .B2(n14303), .A(n14302), .ZN(n14305) );
  NAND2_X1 U15648 ( .A1(n14305), .A2(n15963), .ZN(n14311) );
  NAND2_X1 U15649 ( .A1(n14359), .A2(n14767), .ZN(n14307) );
  NAND2_X1 U15650 ( .A1(n14358), .A2(n14765), .ZN(n14306) );
  AND2_X1 U15651 ( .A1(n14307), .A2(n14306), .ZN(n14821) );
  OAI22_X1 U15652 ( .A1(n14821), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14308), .ZN(n14309) );
  AOI21_X1 U15653 ( .B1(n14647), .B2(n14352), .A(n14309), .ZN(n14310) );
  OAI211_X1 U15654 ( .C1(n14823), .C2(n14348), .A(n14311), .B(n14310), .ZN(
        P1_U3229) );
  OAI211_X1 U15655 ( .C1(n14314), .C2(n14313), .A(n14312), .B(n15963), .ZN(
        n14320) );
  INV_X1 U15656 ( .A(n14315), .ZN(n14718) );
  AOI22_X1 U15657 ( .A1(n14316), .A2(n14360), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14317) );
  OAI21_X1 U15658 ( .B1(n15943), .B2(n15945), .A(n14317), .ZN(n14318) );
  AOI21_X1 U15659 ( .B1(n14718), .B2(n14352), .A(n14318), .ZN(n14319) );
  OAI211_X1 U15660 ( .C1(n14721), .C2(n14348), .A(n14320), .B(n14319), .ZN(
        P1_U3233) );
  AOI21_X1 U15661 ( .B1(n14322), .B2(n14321), .A(n15949), .ZN(n14324) );
  NAND2_X1 U15662 ( .A1(n14324), .A2(n14323), .ZN(n14329) );
  AOI22_X1 U15663 ( .A1(n14359), .A2(n14765), .B1(n14767), .B2(n14360), .ZN(
        n14684) );
  INV_X1 U15664 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14325) );
  OAI22_X1 U15665 ( .A1(n14684), .A2(n14326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14325), .ZN(n14327) );
  AOI21_X1 U15666 ( .B1(n14689), .B2(n14352), .A(n14327), .ZN(n14328) );
  OAI211_X1 U15667 ( .C1(n14348), .C2(n14692), .A(n14329), .B(n14328), .ZN(
        P1_U3235) );
  NAND2_X1 U15668 ( .A1(n14332), .A2(n14331), .ZN(n14333) );
  XNOR2_X1 U15669 ( .A(n14330), .B(n14333), .ZN(n14340) );
  INV_X1 U15670 ( .A(n14616), .ZN(n14337) );
  INV_X1 U15671 ( .A(n14358), .ZN(n14335) );
  OAI22_X1 U15672 ( .A1(n14335), .A2(n15903), .B1(n14334), .B2(n15901), .ZN(
        n14613) );
  AOI22_X1 U15673 ( .A1(n14613), .A2(n15960), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14336) );
  OAI21_X1 U15674 ( .B1(n14337), .B2(n15969), .A(n14336), .ZN(n14338) );
  AOI21_X1 U15675 ( .B1(n14810), .B2(n15965), .A(n14338), .ZN(n14339) );
  OAI21_X1 U15676 ( .B1(n14340), .B2(n15949), .A(n14339), .ZN(P1_U3240) );
  INV_X1 U15677 ( .A(n14341), .ZN(n14342) );
  AOI21_X1 U15678 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14354) );
  NAND2_X1 U15679 ( .A1(n14345), .A2(n14362), .ZN(n14347) );
  OAI211_X1 U15680 ( .C1(n15942), .C2(n15904), .A(n14347), .B(n14346), .ZN(
        n14350) );
  NOR2_X1 U15681 ( .A1(n15878), .A2(n14348), .ZN(n14349) );
  AOI211_X1 U15682 ( .C1(n14352), .C2(n14351), .A(n14350), .B(n14349), .ZN(
        n14353) );
  OAI21_X1 U15683 ( .B1(n14354), .B2(n15949), .A(n14353), .ZN(P1_U3241) );
  MUX2_X1 U15684 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14562), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15685 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14581), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15686 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14355), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15687 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14586), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15688 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14356), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15689 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14357), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15690 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14358), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15691 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14663), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15692 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14359), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15693 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14662), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14360), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14730), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14744), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15697 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n7876), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15698 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14766), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15699 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14361), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15700 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14768), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14362), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14363), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14364), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14365), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14366), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15706 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14367), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15707 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14368), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15708 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14369), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15709 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14370), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15710 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14371), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15711 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14372), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15712 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14373), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15713 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14374), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15714 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8961), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15715 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14375), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U15716 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15531) );
  NAND3_X1 U15717 ( .A1(n14546), .A2(P1_IR_REG_0__SCAN_IN), .A3(n15531), .ZN(
        n14382) );
  AOI22_X1 U15718 ( .A1(n14521), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14381) );
  AOI21_X1 U15719 ( .B1(n15531), .B2(n14886), .A(n14377), .ZN(n14376) );
  MUX2_X1 U15720 ( .A(n14377), .B(n14376), .S(n8937), .Z(n14378) );
  NAND2_X1 U15721 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  NAND3_X1 U15722 ( .A1(n14382), .A2(n14381), .A3(n14380), .ZN(P1_U3243) );
  INV_X1 U15723 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14384) );
  OAI22_X1 U15724 ( .A1(n14557), .A2(n14384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14383), .ZN(n14385) );
  AOI21_X1 U15725 ( .B1(n14551), .B2(n14386), .A(n14385), .ZN(n14394) );
  OAI211_X1 U15726 ( .C1(n14389), .C2(n14388), .A(n14546), .B(n14387), .ZN(
        n14393) );
  OAI211_X1 U15727 ( .C1(n10368), .C2(n14391), .A(n14553), .B(n14399), .ZN(
        n14392) );
  NAND3_X1 U15728 ( .A1(n14394), .A2(n14393), .A3(n14392), .ZN(P1_U3244) );
  OAI22_X1 U15729 ( .A1(n14557), .A2(n15226), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14395), .ZN(n14396) );
  AOI21_X1 U15730 ( .B1(n14551), .B2(n14397), .A(n14396), .ZN(n14407) );
  MUX2_X1 U15731 ( .A(n10366), .B(P1_REG2_REG_2__SCAN_IN), .S(n14397), .Z(
        n14400) );
  NAND3_X1 U15732 ( .A1(n14400), .A2(n14399), .A3(n14398), .ZN(n14401) );
  NAND3_X1 U15733 ( .A1(n14553), .A2(n14416), .A3(n14401), .ZN(n14406) );
  OAI211_X1 U15734 ( .C1(n14404), .C2(n14403), .A(n14546), .B(n14402), .ZN(
        n14405) );
  NAND4_X1 U15735 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        P1_U3245) );
  OAI211_X1 U15736 ( .C1(n14411), .C2(n14410), .A(n14546), .B(n14409), .ZN(
        n14423) );
  NOR2_X1 U15737 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11363), .ZN(n14412) );
  AOI21_X1 U15738 ( .B1(n14521), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14412), .ZN(
        n14422) );
  NAND2_X1 U15739 ( .A1(n14551), .A2(n14413), .ZN(n14421) );
  MUX2_X1 U15740 ( .A(n14414), .B(P1_REG2_REG_3__SCAN_IN), .S(n14413), .Z(
        n14417) );
  NAND3_X1 U15741 ( .A1(n14417), .A2(n14416), .A3(n14415), .ZN(n14418) );
  NAND3_X1 U15742 ( .A1(n14553), .A2(n14419), .A3(n14418), .ZN(n14420) );
  NAND4_X1 U15743 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        P1_U3246) );
  NAND2_X1 U15744 ( .A1(n14425), .A2(n14424), .ZN(n14426) );
  NAND3_X1 U15745 ( .A1(n14546), .A2(n14427), .A3(n14426), .ZN(n14438) );
  INV_X1 U15746 ( .A(n14428), .ZN(n14429) );
  AOI21_X1 U15747 ( .B1(n14521), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14429), .ZN(
        n14437) );
  NAND2_X1 U15748 ( .A1(n14551), .A2(n14430), .ZN(n14436) );
  MUX2_X1 U15749 ( .A(n10524), .B(P1_REG2_REG_6__SCAN_IN), .S(n14430), .Z(
        n14431) );
  NAND3_X1 U15750 ( .A1(n14433), .A2(n14432), .A3(n14431), .ZN(n14434) );
  NAND3_X1 U15751 ( .A1(n14553), .A2(n14446), .A3(n14434), .ZN(n14435) );
  NAND4_X1 U15752 ( .A1(n14438), .A2(n14437), .A3(n14436), .A4(n14435), .ZN(
        P1_U3249) );
  OAI211_X1 U15753 ( .C1(n14441), .C2(n14440), .A(n14546), .B(n14439), .ZN(
        n14453) );
  NOR2_X1 U15754 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14442), .ZN(n14443) );
  AOI21_X1 U15755 ( .B1(n14521), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14443), .ZN(
        n14452) );
  MUX2_X1 U15756 ( .A(n10527), .B(P1_REG2_REG_7__SCAN_IN), .S(n14449), .Z(
        n14444) );
  NAND3_X1 U15757 ( .A1(n14446), .A2(n14445), .A3(n14444), .ZN(n14447) );
  NAND3_X1 U15758 ( .A1(n14553), .A2(n14448), .A3(n14447), .ZN(n14451) );
  NAND2_X1 U15759 ( .A1(n14551), .A2(n14449), .ZN(n14450) );
  NAND4_X1 U15760 ( .A1(n14453), .A2(n14452), .A3(n14451), .A4(n14450), .ZN(
        P1_U3250) );
  OAI21_X1 U15761 ( .B1(n14456), .B2(n14455), .A(n14454), .ZN(n14457) );
  NAND2_X1 U15762 ( .A1(n14546), .A2(n14457), .ZN(n14468) );
  INV_X1 U15763 ( .A(n14458), .ZN(n14459) );
  AOI21_X1 U15764 ( .B1(n14521), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14459), .ZN(
        n14467) );
  MUX2_X1 U15765 ( .A(n10555), .B(P1_REG2_REG_9__SCAN_IN), .S(n14464), .Z(
        n14460) );
  NAND3_X1 U15766 ( .A1(n14462), .A2(n14461), .A3(n14460), .ZN(n14463) );
  NAND3_X1 U15767 ( .A1(n14553), .A2(n14477), .A3(n14463), .ZN(n14466) );
  NAND2_X1 U15768 ( .A1(n14551), .A2(n14464), .ZN(n14465) );
  NAND4_X1 U15769 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        P1_U3252) );
  AOI21_X1 U15770 ( .B1(n14470), .B2(n14469), .A(n14548), .ZN(n14472) );
  NAND2_X1 U15771 ( .A1(n14472), .A2(n14471), .ZN(n14483) );
  INV_X1 U15772 ( .A(n14473), .ZN(n14474) );
  AOI21_X1 U15773 ( .B1(n14521), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14474), 
        .ZN(n14482) );
  MUX2_X1 U15774 ( .A(n10558), .B(P1_REG2_REG_10__SCAN_IN), .S(n14479), .Z(
        n14475) );
  NAND3_X1 U15775 ( .A1(n14477), .A2(n14476), .A3(n14475), .ZN(n14478) );
  NAND3_X1 U15776 ( .A1(n14553), .A2(n14493), .A3(n14478), .ZN(n14481) );
  NAND2_X1 U15777 ( .A1(n14551), .A2(n14479), .ZN(n14480) );
  NAND4_X1 U15778 ( .A1(n14483), .A2(n14482), .A3(n14481), .A4(n14480), .ZN(
        P1_U3253) );
  OAI21_X1 U15779 ( .B1(n14486), .B2(n14485), .A(n14484), .ZN(n14487) );
  NAND2_X1 U15780 ( .A1(n14487), .A2(n14546), .ZN(n14500) );
  INV_X1 U15781 ( .A(n14488), .ZN(n14489) );
  AOI21_X1 U15782 ( .B1(n14521), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n14489), 
        .ZN(n14499) );
  INV_X1 U15783 ( .A(n14490), .ZN(n14495) );
  NAND3_X1 U15784 ( .A1(n14493), .A2(n14492), .A3(n14491), .ZN(n14494) );
  NAND3_X1 U15785 ( .A1(n14495), .A2(n14553), .A3(n14494), .ZN(n14498) );
  NAND2_X1 U15786 ( .A1(n14551), .A2(n14496), .ZN(n14497) );
  NAND4_X1 U15787 ( .A1(n14500), .A2(n14499), .A3(n14498), .A4(n14497), .ZN(
        P1_U3254) );
  NAND2_X1 U15788 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n15906)
         );
  INV_X1 U15789 ( .A(n15906), .ZN(n14502) );
  NOR2_X1 U15790 ( .A1(n14518), .A2(n14530), .ZN(n14501) );
  AOI211_X1 U15791 ( .C1(n14521), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n14502), 
        .B(n14501), .ZN(n14517) );
  INV_X1 U15792 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15925) );
  NOR2_X1 U15793 ( .A1(n14523), .A2(n15925), .ZN(n14503) );
  AOI21_X1 U15794 ( .B1(n14523), .B2(n15925), .A(n14503), .ZN(n14507) );
  AOI21_X1 U15795 ( .B1(n14505), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14504), 
        .ZN(n14506) );
  NOR2_X1 U15796 ( .A1(n14506), .A2(n14507), .ZN(n14522) );
  AOI211_X1 U15797 ( .C1(n14507), .C2(n14506), .A(n14522), .B(n14548), .ZN(
        n14508) );
  INV_X1 U15798 ( .A(n14508), .ZN(n14516) );
  INV_X1 U15799 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14529) );
  NOR2_X1 U15800 ( .A1(n14530), .A2(n14529), .ZN(n14509) );
  AOI21_X1 U15801 ( .B1(n14529), .B2(n14530), .A(n14509), .ZN(n14514) );
  OAI21_X1 U15802 ( .B1(n14512), .B2(n14511), .A(n14510), .ZN(n14513) );
  NAND2_X1 U15803 ( .A1(n14514), .A2(n14513), .ZN(n14528) );
  OAI211_X1 U15804 ( .C1(n14514), .C2(n14513), .A(n14553), .B(n14528), .ZN(
        n14515) );
  NAND3_X1 U15805 ( .A1(n14517), .A2(n14516), .A3(n14515), .ZN(P1_U3260) );
  NAND2_X1 U15806 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n15954)
         );
  INV_X1 U15807 ( .A(n15954), .ZN(n14520) );
  NOR2_X1 U15808 ( .A1(n14518), .A2(n14535), .ZN(n14519) );
  AOI211_X1 U15809 ( .C1(n14521), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14520), 
        .B(n14519), .ZN(n14534) );
  AOI21_X1 U15810 ( .B1(n14523), .B2(P1_REG1_REG_17__SCAN_IN), .A(n14522), 
        .ZN(n14536) );
  XNOR2_X1 U15811 ( .A(n14535), .B(n14536), .ZN(n14524) );
  INV_X1 U15812 ( .A(n14524), .ZN(n14527) );
  INV_X1 U15813 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U15814 ( .A1(n14525), .A2(n14524), .ZN(n14538) );
  INV_X1 U15815 ( .A(n14538), .ZN(n14526) );
  OAI211_X1 U15816 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14527), .A(n14546), 
        .B(n14526), .ZN(n14533) );
  OAI21_X1 U15817 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n14541) );
  XNOR2_X1 U15818 ( .A(n14535), .B(n14541), .ZN(n14531) );
  NAND2_X1 U15819 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14531), .ZN(n14544) );
  OAI211_X1 U15820 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14531), .A(n14553), 
        .B(n14544), .ZN(n14532) );
  NAND3_X1 U15821 ( .A1(n14534), .A2(n14533), .A3(n14532), .ZN(P1_U3261) );
  NOR2_X1 U15822 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  NOR2_X1 U15823 ( .A1(n14538), .A2(n14537), .ZN(n14540) );
  INV_X1 U15824 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14539) );
  XOR2_X1 U15825 ( .A(n14540), .B(n14539), .Z(n14549) );
  NAND2_X1 U15826 ( .A1(n14542), .A2(n14541), .ZN(n14543) );
  NAND2_X1 U15827 ( .A1(n14544), .A2(n14543), .ZN(n14545) );
  XOR2_X1 U15828 ( .A(n14545), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14547) );
  AOI22_X1 U15829 ( .A1(n14549), .A2(n14546), .B1(n14553), .B2(n14547), .ZN(
        n14555) );
  INV_X1 U15830 ( .A(n14547), .ZN(n14552) );
  NOR2_X1 U15831 ( .A1(n14549), .A2(n14548), .ZN(n14550) );
  AOI211_X1 U15832 ( .C1(n14553), .C2(n14552), .A(n14551), .B(n14550), .ZN(
        n14554) );
  MUX2_X1 U15833 ( .A(n14555), .B(n14554), .S(n15537), .Z(n14556) );
  NAND2_X1 U15834 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n15966)
         );
  OAI211_X1 U15835 ( .C1(n8152), .C2(n14557), .A(n14556), .B(n15966), .ZN(
        P1_U3262) );
  NAND2_X1 U15836 ( .A1(n14559), .A2(n15917), .ZN(n14780) );
  NAND2_X1 U15837 ( .A1(n14560), .A2(P1_B_REG_SCAN_IN), .ZN(n14561) );
  AND2_X1 U15838 ( .A1(n14765), .A2(n14561), .ZN(n14580) );
  NAND2_X1 U15839 ( .A1(n14562), .A2(n14580), .ZN(n14782) );
  NOR2_X1 U15840 ( .A1(n15941), .A2(n14782), .ZN(n14566) );
  NOR2_X1 U15841 ( .A1(n14781), .A2(n15723), .ZN(n14563) );
  AOI211_X1 U15842 ( .C1(n15941), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14566), 
        .B(n14563), .ZN(n14564) );
  OAI21_X1 U15843 ( .B1(n14672), .B2(n14780), .A(n14564), .ZN(P1_U3263) );
  OAI211_X1 U15844 ( .C1(n14784), .C2(n14577), .A(n15917), .B(n7307), .ZN(
        n14783) );
  NOR2_X1 U15845 ( .A1(n14784), .A2(n15723), .ZN(n14565) );
  AOI211_X1 U15846 ( .C1(n15941), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14566), 
        .B(n14565), .ZN(n14567) );
  OAI21_X1 U15847 ( .B1(n14672), .B2(n14783), .A(n14567), .ZN(P1_U3264) );
  XNOR2_X1 U15848 ( .A(n14571), .B(n14570), .ZN(n14785) );
  INV_X1 U15849 ( .A(n14785), .ZN(n14593) );
  NAND2_X1 U15850 ( .A1(n14573), .A2(n14572), .ZN(n14575) );
  XNOR2_X1 U15851 ( .A(n14575), .B(n14574), .ZN(n14786) );
  NAND2_X1 U15852 ( .A1(n14786), .A2(n15936), .ZN(n14592) );
  INV_X1 U15853 ( .A(n14576), .ZN(n14578) );
  NAND2_X1 U15854 ( .A1(n14581), .A2(n14580), .ZN(n14788) );
  INV_X1 U15855 ( .A(n14582), .ZN(n14583) );
  OAI22_X1 U15856 ( .A1(n14585), .A2(n14788), .B1(n14584), .B2(n14583), .ZN(
        n14588) );
  NAND2_X1 U15857 ( .A1(n14586), .A2(n14767), .ZN(n14789) );
  NOR2_X1 U15858 ( .A1(n15941), .A2(n14789), .ZN(n14587) );
  AOI211_X1 U15859 ( .C1(n15941), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14588), 
        .B(n14587), .ZN(n14589) );
  OAI21_X1 U15860 ( .B1(n14790), .B2(n15723), .A(n14589), .ZN(n14590) );
  AOI21_X1 U15861 ( .B1(n14787), .B2(n15935), .A(n14590), .ZN(n14591) );
  OAI211_X1 U15862 ( .C1(n14593), .C2(n14779), .A(n14592), .B(n14591), .ZN(
        P1_U3356) );
  XNOR2_X1 U15863 ( .A(n14594), .B(n14599), .ZN(n14597) );
  INV_X1 U15864 ( .A(n14595), .ZN(n14596) );
  OAI21_X1 U15865 ( .B1(n14600), .B2(n14599), .A(n14598), .ZN(n14806) );
  AOI21_X1 U15866 ( .B1(n14612), .B2(n14604), .A(n14763), .ZN(n14602) );
  NAND2_X1 U15867 ( .A1(n14602), .A2(n14601), .ZN(n14803) );
  AOI22_X1 U15868 ( .A1(n15941), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14603), 
        .B2(n15930), .ZN(n14606) );
  NAND2_X1 U15869 ( .A1(n14604), .A2(n15931), .ZN(n14605) );
  OAI211_X1 U15870 ( .C1(n14803), .C2(n14672), .A(n14606), .B(n14605), .ZN(
        n14607) );
  AOI21_X1 U15871 ( .B1(n14806), .B2(n15936), .A(n14607), .ZN(n14608) );
  OAI21_X1 U15872 ( .B1(n15941), .B2(n14807), .A(n14608), .ZN(P1_U3266) );
  XNOR2_X1 U15873 ( .A(n14610), .B(n14609), .ZN(n14611) );
  NAND2_X1 U15874 ( .A1(n14611), .A2(n15914), .ZN(n14811) );
  OAI211_X1 U15875 ( .C1(n14633), .C2(n14618), .A(n14612), .B(n15917), .ZN(
        n14615) );
  INV_X1 U15876 ( .A(n14613), .ZN(n14614) );
  NAND2_X1 U15877 ( .A1(n14615), .A2(n14614), .ZN(n14809) );
  AOI22_X1 U15878 ( .A1(n15941), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14616), 
        .B2(n15930), .ZN(n14617) );
  OAI21_X1 U15879 ( .B1(n14618), .B2(n15723), .A(n14617), .ZN(n14623) );
  OAI21_X1 U15880 ( .B1(n14621), .B2(n14620), .A(n14619), .ZN(n14813) );
  NOR2_X1 U15881 ( .A1(n14813), .A2(n14740), .ZN(n14622) );
  AOI211_X1 U15882 ( .C1(n15935), .C2(n14809), .A(n14623), .B(n14622), .ZN(
        n14624) );
  OAI21_X1 U15883 ( .B1(n15941), .B2(n14811), .A(n14624), .ZN(P1_U3267) );
  OAI21_X1 U15884 ( .B1(n14626), .B2(n14630), .A(n14625), .ZN(n14627) );
  INV_X1 U15885 ( .A(n14627), .ZN(n14820) );
  NAND2_X1 U15886 ( .A1(n14629), .A2(n14630), .ZN(n14814) );
  NAND3_X1 U15887 ( .A1(n14628), .A2(n14814), .A3(n15936), .ZN(n14641) );
  NAND2_X1 U15888 ( .A1(n14645), .A2(n14817), .ZN(n14631) );
  NAND2_X1 U15889 ( .A1(n14631), .A2(n15917), .ZN(n14632) );
  NOR2_X1 U15890 ( .A1(n14633), .A2(n14632), .ZN(n14815) );
  INV_X1 U15891 ( .A(n14634), .ZN(n14816) );
  AOI22_X1 U15892 ( .A1(n14816), .A2(n14772), .B1(n14635), .B2(n15930), .ZN(
        n14637) );
  NAND2_X1 U15893 ( .A1(n15941), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14636) );
  OAI211_X1 U15894 ( .C1(n14638), .C2(n15723), .A(n14637), .B(n14636), .ZN(
        n14639) );
  AOI21_X1 U15895 ( .B1(n14815), .B2(n15935), .A(n14639), .ZN(n14640) );
  OAI211_X1 U15896 ( .C1(n14820), .C2(n14779), .A(n14641), .B(n14640), .ZN(
        P1_U3268) );
  XNOR2_X1 U15897 ( .A(n14642), .B(n7960), .ZN(n14827) );
  XNOR2_X1 U15898 ( .A(n14643), .B(n14644), .ZN(n14825) );
  AOI21_X1 U15899 ( .B1(n14660), .B2(n14651), .A(n14763), .ZN(n14646) );
  NAND2_X1 U15900 ( .A1(n14646), .A2(n14645), .ZN(n14822) );
  NAND2_X1 U15901 ( .A1(n15930), .A2(n14647), .ZN(n14649) );
  NAND2_X1 U15902 ( .A1(n15941), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n14648) );
  OAI211_X1 U15903 ( .C1(n14821), .C2(n15941), .A(n14649), .B(n14648), .ZN(
        n14650) );
  AOI21_X1 U15904 ( .B1(n14651), .B2(n15931), .A(n14650), .ZN(n14652) );
  OAI21_X1 U15905 ( .B1(n14822), .B2(n14672), .A(n14652), .ZN(n14653) );
  AOI21_X1 U15906 ( .B1(n14825), .B2(n15936), .A(n14653), .ZN(n14654) );
  OAI21_X1 U15907 ( .B1(n14827), .B2(n14779), .A(n14654), .ZN(P1_U3269) );
  XNOR2_X1 U15908 ( .A(n14655), .B(n14658), .ZN(n14834) );
  AND2_X1 U15909 ( .A1(n14657), .A2(n14656), .ZN(n14659) );
  XNOR2_X1 U15910 ( .A(n14659), .B(n14658), .ZN(n14832) );
  AOI21_X1 U15911 ( .B1(n14686), .B2(n14670), .A(n14763), .ZN(n14661) );
  NAND2_X1 U15912 ( .A1(n14661), .A2(n14660), .ZN(n14829) );
  AOI22_X1 U15913 ( .A1(n14663), .A2(n14765), .B1(n14767), .B2(n14662), .ZN(
        n14828) );
  NAND2_X1 U15914 ( .A1(n15930), .A2(n14664), .ZN(n14665) );
  NAND2_X1 U15915 ( .A1(n14828), .A2(n14665), .ZN(n14666) );
  NAND2_X1 U15916 ( .A1(n14666), .A2(n14772), .ZN(n14667) );
  OAI21_X1 U15917 ( .B1(n14772), .B2(n14668), .A(n14667), .ZN(n14669) );
  AOI21_X1 U15918 ( .B1(n14670), .B2(n15931), .A(n14669), .ZN(n14671) );
  OAI21_X1 U15919 ( .B1(n14829), .B2(n14672), .A(n14671), .ZN(n14673) );
  AOI21_X1 U15920 ( .B1(n14832), .B2(n15936), .A(n14673), .ZN(n14674) );
  OAI21_X1 U15921 ( .B1(n14834), .B2(n14779), .A(n14674), .ZN(P1_U3270) );
  NAND2_X1 U15922 ( .A1(n14676), .A2(n14677), .ZN(n14679) );
  XNOR2_X1 U15923 ( .A(n14679), .B(n14678), .ZN(n14839) );
  INV_X1 U15924 ( .A(n14680), .ZN(n14681) );
  AOI21_X1 U15925 ( .B1(n14683), .B2(n14682), .A(n14681), .ZN(n14685) );
  OAI21_X1 U15926 ( .B1(n14685), .B2(n15890), .A(n14684), .ZN(n14835) );
  INV_X1 U15927 ( .A(n14692), .ZN(n14837) );
  INV_X1 U15928 ( .A(n14704), .ZN(n14688) );
  INV_X1 U15929 ( .A(n14686), .ZN(n14687) );
  AOI211_X1 U15930 ( .C1(n14837), .C2(n14688), .A(n14763), .B(n14687), .ZN(
        n14836) );
  NAND2_X1 U15931 ( .A1(n14836), .A2(n15935), .ZN(n14691) );
  AOI22_X1 U15932 ( .A1(n15941), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14689), 
        .B2(n15930), .ZN(n14690) );
  OAI211_X1 U15933 ( .C1(n15723), .C2(n14692), .A(n14691), .B(n14690), .ZN(
        n14693) );
  AOI21_X1 U15934 ( .B1(n14835), .B2(n14772), .A(n14693), .ZN(n14694) );
  OAI21_X1 U15935 ( .B1(n14839), .B2(n14740), .A(n14694), .ZN(P1_U3271) );
  OAI211_X1 U15936 ( .C1(n14696), .C2(n14701), .A(n14695), .B(n15914), .ZN(
        n14698) );
  AND2_X1 U15937 ( .A1(n14698), .A2(n14697), .ZN(n14843) );
  INV_X1 U15938 ( .A(n14676), .ZN(n14699) );
  AOI21_X1 U15939 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14844) );
  INV_X1 U15940 ( .A(n14844), .ZN(n14709) );
  NAND2_X1 U15941 ( .A1(n14841), .A2(n14715), .ZN(n14702) );
  NAND2_X1 U15942 ( .A1(n14702), .A2(n15917), .ZN(n14703) );
  NOR2_X1 U15943 ( .A1(n14704), .A2(n14703), .ZN(n14840) );
  NAND2_X1 U15944 ( .A1(n14840), .A2(n15935), .ZN(n14707) );
  AOI22_X1 U15945 ( .A1(n15941), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14705), 
        .B2(n15930), .ZN(n14706) );
  OAI211_X1 U15946 ( .C1(n12438), .C2(n15723), .A(n14707), .B(n14706), .ZN(
        n14708) );
  AOI21_X1 U15947 ( .B1(n14709), .B2(n15936), .A(n14708), .ZN(n14710) );
  OAI21_X1 U15948 ( .B1(n15941), .B2(n14843), .A(n14710), .ZN(P1_U3272) );
  OAI21_X1 U15949 ( .B1(n14712), .B2(n14714), .A(n14711), .ZN(n14851) );
  NAND2_X1 U15950 ( .A1(n14713), .A2(n14714), .ZN(n14845) );
  NAND3_X1 U15951 ( .A1(n7212), .A2(n14845), .A3(n15936), .ZN(n14724) );
  AOI21_X1 U15952 ( .B1(n14848), .B2(n14732), .A(n14763), .ZN(n14716) );
  AND2_X1 U15953 ( .A1(n14716), .A2(n14715), .ZN(n14846) );
  OAI22_X1 U15954 ( .A1(n15943), .A2(n15903), .B1(n14717), .B2(n15901), .ZN(
        n14847) );
  AOI22_X1 U15955 ( .A1(n14847), .A2(n14772), .B1(n14718), .B2(n15930), .ZN(
        n14720) );
  NAND2_X1 U15956 ( .A1(n15941), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14719) );
  OAI211_X1 U15957 ( .C1(n14721), .C2(n15723), .A(n14720), .B(n14719), .ZN(
        n14722) );
  AOI21_X1 U15958 ( .B1(n15935), .B2(n14846), .A(n14722), .ZN(n14723) );
  OAI211_X1 U15959 ( .C1(n14851), .C2(n14779), .A(n14724), .B(n14723), .ZN(
        P1_U3273) );
  XNOR2_X1 U15960 ( .A(n14726), .B(n14725), .ZN(n14855) );
  AOI21_X1 U15961 ( .B1(n14729), .B2(n14728), .A(n14727), .ZN(n14731) );
  AOI22_X1 U15962 ( .A1(n14765), .A2(n14730), .B1(n7876), .B2(n14767), .ZN(
        n15959) );
  OAI21_X1 U15963 ( .B1(n14731), .B2(n15890), .A(n15959), .ZN(n14852) );
  INV_X1 U15964 ( .A(n14732), .ZN(n14733) );
  AOI211_X1 U15965 ( .C1(n15964), .C2(n7565), .A(n14763), .B(n14733), .ZN(
        n14853) );
  NAND2_X1 U15966 ( .A1(n14853), .A2(n15935), .ZN(n14736) );
  INV_X1 U15967 ( .A(n15968), .ZN(n14734) );
  AOI22_X1 U15968 ( .A1(n15941), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14734), 
        .B2(n15930), .ZN(n14735) );
  OAI211_X1 U15969 ( .C1(n14737), .C2(n15723), .A(n14736), .B(n14735), .ZN(
        n14738) );
  AOI21_X1 U15970 ( .B1(n14852), .B2(n14772), .A(n14738), .ZN(n14739) );
  OAI21_X1 U15971 ( .B1(n14855), .B2(n14740), .A(n14739), .ZN(P1_U3274) );
  OAI211_X1 U15972 ( .C1(n14743), .C2(n14742), .A(n14741), .B(n15914), .ZN(
        n14746) );
  AOI22_X1 U15973 ( .A1(n14744), .A2(n14765), .B1(n14767), .B2(n14766), .ZN(
        n14745) );
  AND2_X1 U15974 ( .A1(n14746), .A2(n14745), .ZN(n14859) );
  OAI21_X1 U15975 ( .B1(n14749), .B2(n14748), .A(n14747), .ZN(n14856) );
  NAND2_X1 U15976 ( .A1(n15953), .A2(n15916), .ZN(n14750) );
  NAND2_X1 U15977 ( .A1(n14750), .A2(n15917), .ZN(n14751) );
  NOR2_X1 U15978 ( .A1(n14752), .A2(n14751), .ZN(n14857) );
  NAND2_X1 U15979 ( .A1(n14857), .A2(n15935), .ZN(n14755) );
  AOI22_X1 U15980 ( .A1(n15941), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14753), 
        .B2(n15930), .ZN(n14754) );
  OAI211_X1 U15981 ( .C1(n7877), .C2(n15723), .A(n14755), .B(n14754), .ZN(
        n14756) );
  AOI21_X1 U15982 ( .B1(n14856), .B2(n15936), .A(n14756), .ZN(n14757) );
  OAI21_X1 U15983 ( .B1(n15941), .B2(n14859), .A(n14757), .ZN(P1_U3275) );
  OAI21_X1 U15984 ( .B1(n14759), .B2(n14761), .A(n14758), .ZN(n14760) );
  INV_X1 U15985 ( .A(n14760), .ZN(n15891) );
  XNOR2_X1 U15986 ( .A(n14762), .B(n14761), .ZN(n15893) );
  NAND2_X1 U15987 ( .A1(n15893), .A2(n15936), .ZN(n14778) );
  AOI211_X1 U15988 ( .C1(n15888), .C2(n14764), .A(n14763), .B(n15918), .ZN(
        n15885) );
  NAND2_X1 U15989 ( .A1(n14766), .A2(n14765), .ZN(n14770) );
  NAND2_X1 U15990 ( .A1(n14768), .A2(n14767), .ZN(n14769) );
  NAND2_X1 U15991 ( .A1(n14770), .A2(n14769), .ZN(n15886) );
  AOI22_X1 U15992 ( .A1(n14772), .A2(n15886), .B1(n14771), .B2(n15930), .ZN(
        n14774) );
  NAND2_X1 U15993 ( .A1(n15941), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14773) );
  OAI211_X1 U15994 ( .C1(n14775), .C2(n15723), .A(n14774), .B(n14773), .ZN(
        n14776) );
  AOI21_X1 U15995 ( .B1(n15885), .B2(n15935), .A(n14776), .ZN(n14777) );
  OAI211_X1 U15996 ( .C1(n15891), .C2(n14779), .A(n14778), .B(n14777), .ZN(
        P1_U3277) );
  OAI211_X1 U15997 ( .C1(n15919), .C2(n14781), .A(n14780), .B(n14782), .ZN(
        n14861) );
  MUX2_X1 U15998 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14861), .S(n15717), .Z(
        P1_U3559) );
  OAI211_X1 U15999 ( .C1(n15919), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14862) );
  MUX2_X1 U16000 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14862), .S(n15717), .Z(
        P1_U3558) );
  NAND2_X1 U16001 ( .A1(n14786), .A2(n15923), .ZN(n14794) );
  OAI211_X1 U16002 ( .C1(n14790), .C2(n15919), .A(n14789), .B(n14788), .ZN(
        n14791) );
  INV_X1 U16003 ( .A(n14791), .ZN(n14792) );
  NAND3_X1 U16004 ( .A1(n14797), .A2(n14796), .A3(n15923), .ZN(n14802) );
  AOI21_X1 U16005 ( .B1(n14799), .B2(n15887), .A(n14798), .ZN(n14800) );
  NAND3_X1 U16006 ( .A1(n14802), .A2(n14801), .A3(n14800), .ZN(n14863) );
  MUX2_X1 U16007 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14863), .S(n15717), .Z(
        P1_U3556) );
  OAI21_X1 U16008 ( .B1(n14804), .B2(n15919), .A(n14803), .ZN(n14805) );
  AOI21_X1 U16009 ( .B1(n14806), .B2(n15923), .A(n14805), .ZN(n14808) );
  MUX2_X1 U16010 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14864), .S(n15717), .Z(
        P1_U3555) );
  AOI21_X1 U16011 ( .B1(n14810), .B2(n15887), .A(n14809), .ZN(n14812) );
  OAI211_X1 U16012 ( .C1(n14813), .C2(n15851), .A(n14812), .B(n14811), .ZN(
        n14865) );
  MUX2_X1 U16013 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14865), .S(n15717), .Z(
        P1_U3554) );
  NAND3_X1 U16014 ( .A1(n14628), .A2(n14814), .A3(n15923), .ZN(n14819) );
  AOI211_X1 U16015 ( .C1(n14817), .C2(n15887), .A(n14816), .B(n14815), .ZN(
        n14818) );
  OAI211_X1 U16016 ( .C1(n15890), .C2(n14820), .A(n14819), .B(n14818), .ZN(
        n14866) );
  MUX2_X1 U16017 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14866), .S(n15717), .Z(
        P1_U3553) );
  OAI211_X1 U16018 ( .C1(n14823), .C2(n15919), .A(n14822), .B(n14821), .ZN(
        n14824) );
  AOI21_X1 U16019 ( .B1(n14825), .B2(n15923), .A(n14824), .ZN(n14826) );
  OAI21_X1 U16020 ( .B1(n15890), .B2(n14827), .A(n14826), .ZN(n14867) );
  MUX2_X1 U16021 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14867), .S(n15717), .Z(
        P1_U3552) );
  OAI211_X1 U16022 ( .C1(n14830), .C2(n15919), .A(n14829), .B(n14828), .ZN(
        n14831) );
  AOI21_X1 U16023 ( .B1(n14832), .B2(n15923), .A(n14831), .ZN(n14833) );
  OAI21_X1 U16024 ( .B1(n15890), .B2(n14834), .A(n14833), .ZN(n14868) );
  MUX2_X1 U16025 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14868), .S(n15717), .Z(
        P1_U3551) );
  AOI211_X1 U16026 ( .C1(n14837), .C2(n15887), .A(n14836), .B(n14835), .ZN(
        n14838) );
  OAI21_X1 U16027 ( .B1(n14839), .B2(n15851), .A(n14838), .ZN(n14869) );
  MUX2_X1 U16028 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14869), .S(n15717), .Z(
        P1_U3550) );
  AOI21_X1 U16029 ( .B1(n14841), .B2(n15887), .A(n14840), .ZN(n14842) );
  OAI211_X1 U16030 ( .C1(n14844), .C2(n15851), .A(n14843), .B(n14842), .ZN(
        n14870) );
  MUX2_X1 U16031 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14870), .S(n15717), .Z(
        P1_U3549) );
  NAND3_X1 U16032 ( .A1(n7212), .A2(n14845), .A3(n15923), .ZN(n14850) );
  AOI211_X1 U16033 ( .C1(n14848), .C2(n15887), .A(n14847), .B(n14846), .ZN(
        n14849) );
  OAI211_X1 U16034 ( .C1(n15890), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        n14871) );
  MUX2_X1 U16035 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14871), .S(n15717), .Z(
        P1_U3548) );
  AOI211_X1 U16036 ( .C1(n15964), .C2(n15887), .A(n14853), .B(n14852), .ZN(
        n14854) );
  OAI21_X1 U16037 ( .B1(n14855), .B2(n15851), .A(n14854), .ZN(n14872) );
  MUX2_X1 U16038 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14872), .S(n15717), .Z(
        P1_U3547) );
  INV_X1 U16039 ( .A(n14856), .ZN(n14860) );
  AOI21_X1 U16040 ( .B1(n15953), .B2(n15887), .A(n14857), .ZN(n14858) );
  OAI211_X1 U16041 ( .C1(n14860), .C2(n15851), .A(n14859), .B(n14858), .ZN(
        n14873) );
  MUX2_X1 U16042 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14873), .S(n15717), .Z(
        P1_U3546) );
  MUX2_X1 U16043 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14861), .S(n15719), .Z(
        P1_U3527) );
  MUX2_X1 U16044 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14862), .S(n15719), .Z(
        P1_U3526) );
  MUX2_X1 U16045 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14863), .S(n15719), .Z(
        P1_U3524) );
  MUX2_X1 U16046 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14864), .S(n15719), .Z(
        P1_U3523) );
  MUX2_X1 U16047 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14865), .S(n15719), .Z(
        P1_U3522) );
  MUX2_X1 U16048 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14866), .S(n15719), .Z(
        P1_U3521) );
  MUX2_X1 U16049 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14867), .S(n15719), .Z(
        P1_U3520) );
  MUX2_X1 U16050 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14868), .S(n15719), .Z(
        P1_U3519) );
  MUX2_X1 U16051 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14869), .S(n15719), .Z(
        P1_U3518) );
  MUX2_X1 U16052 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14870), .S(n15719), .Z(
        P1_U3517) );
  MUX2_X1 U16053 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14871), .S(n15719), .Z(
        P1_U3516) );
  MUX2_X1 U16054 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14872), .S(n15719), .Z(
        P1_U3515) );
  MUX2_X1 U16055 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14873), .S(n15719), .Z(
        P1_U3513) );
  MUX2_X1 U16056 ( .A(n14874), .B(P1_D_REG_0__SCAN_IN), .S(n14901), .Z(
        P1_U3445) );
  NOR4_X1 U16057 ( .A1(n8874), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8979), .A4(
        P1_U3086), .ZN(n14875) );
  AOI21_X1 U16058 ( .B1(n14880), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14875), 
        .ZN(n14876) );
  OAI21_X1 U16059 ( .B1(n14877), .B2(n14893), .A(n14876), .ZN(P1_U3324) );
  AOI22_X1 U16060 ( .A1(n8876), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n14880), .ZN(n14878) );
  OAI21_X1 U16061 ( .B1(n14879), .B2(n14893), .A(n14878), .ZN(P1_U3325) );
  AOI22_X1 U16062 ( .A1(n14881), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n14880), .ZN(n14882) );
  OAI21_X1 U16063 ( .B1(n14883), .B2(n14893), .A(n14882), .ZN(P1_U3326) );
  OAI222_X1 U16064 ( .A1(n14897), .A2(n14885), .B1(n14893), .B2(n14884), .C1(
        P1_U3086), .C2(n9500), .ZN(P1_U3327) );
  OAI222_X1 U16065 ( .A1(n14897), .A2(n14888), .B1(n14893), .B2(n14887), .C1(
        n14886), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16066 ( .A1(n14897), .A2(n14891), .B1(n14893), .B2(n14890), .C1(
        n14889), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U16067 ( .A1(n14897), .A2(n14894), .B1(n14893), .B2(n14892), .C1(
        P1_U3086), .C2(n10439), .ZN(P1_U3330) );
  OAI222_X1 U16068 ( .A1(n14897), .A2(n7737), .B1(n14893), .B2(n14896), .C1(
        P1_U3086), .C2(n10440), .ZN(P1_U3331) );
  MUX2_X1 U16069 ( .A(n14899), .B(n14898), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16070 ( .A(n14900), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16071 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14901), .ZN(P1_U3323) );
  AND2_X1 U16072 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14901), .ZN(P1_U3322) );
  AND2_X1 U16073 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14901), .ZN(P1_U3321) );
  AND2_X1 U16074 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14901), .ZN(P1_U3320) );
  AND2_X1 U16075 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14901), .ZN(P1_U3319) );
  AND2_X1 U16076 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14901), .ZN(P1_U3318) );
  AND2_X1 U16077 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14901), .ZN(P1_U3317) );
  AND2_X1 U16078 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14901), .ZN(P1_U3316) );
  AND2_X1 U16079 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14901), .ZN(P1_U3315) );
  AND2_X1 U16080 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14901), .ZN(P1_U3314) );
  AND2_X1 U16081 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14901), .ZN(P1_U3313) );
  AND2_X1 U16082 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14901), .ZN(P1_U3312) );
  AND2_X1 U16083 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14901), .ZN(P1_U3311) );
  AND2_X1 U16084 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14901), .ZN(P1_U3310) );
  AND2_X1 U16085 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14901), .ZN(P1_U3309) );
  AND2_X1 U16086 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14901), .ZN(P1_U3308) );
  AND2_X1 U16087 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14901), .ZN(P1_U3307) );
  AND2_X1 U16088 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14901), .ZN(P1_U3306) );
  AND2_X1 U16089 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14901), .ZN(P1_U3305) );
  AND2_X1 U16090 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14901), .ZN(P1_U3304) );
  AND2_X1 U16091 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14901), .ZN(P1_U3303) );
  AND2_X1 U16092 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14901), .ZN(P1_U3302) );
  AND2_X1 U16093 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14901), .ZN(P1_U3301) );
  AND2_X1 U16094 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14901), .ZN(P1_U3300) );
  AND2_X1 U16095 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14901), .ZN(P1_U3299) );
  AND2_X1 U16096 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14901), .ZN(P1_U3298) );
  AND2_X1 U16097 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14901), .ZN(P1_U3297) );
  AND2_X1 U16098 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14901), .ZN(P1_U3296) );
  AND2_X1 U16099 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14901), .ZN(P1_U3295) );
  AND2_X1 U16100 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14901), .ZN(P1_U3294) );
  AOI21_X1 U16101 ( .B1(n14903), .B2(n15137), .A(n14902), .ZN(P2_U3417) );
  AND2_X1 U16102 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14905), .ZN(P2_U3295) );
  AND2_X1 U16103 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14905), .ZN(P2_U3294) );
  AND2_X1 U16104 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14905), .ZN(P2_U3293) );
  AND2_X1 U16105 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14905), .ZN(P2_U3292) );
  AND2_X1 U16106 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14905), .ZN(P2_U3291) );
  AND2_X1 U16107 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14905), .ZN(P2_U3290) );
  AND2_X1 U16108 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14905), .ZN(P2_U3289) );
  AND2_X1 U16109 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14905), .ZN(P2_U3288) );
  AND2_X1 U16110 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14905), .ZN(P2_U3287) );
  AND2_X1 U16111 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14905), .ZN(P2_U3286) );
  AND2_X1 U16112 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14905), .ZN(P2_U3285) );
  AND2_X1 U16113 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14905), .ZN(P2_U3284) );
  AND2_X1 U16114 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14905), .ZN(P2_U3283) );
  AND2_X1 U16115 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14905), .ZN(P2_U3282) );
  AND2_X1 U16116 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14905), .ZN(P2_U3281) );
  AND2_X1 U16117 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14905), .ZN(P2_U3280) );
  AND2_X1 U16118 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14905), .ZN(P2_U3279) );
  AND2_X1 U16119 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14905), .ZN(P2_U3278) );
  AND2_X1 U16120 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14905), .ZN(P2_U3277) );
  AND2_X1 U16121 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14905), .ZN(P2_U3276) );
  AND2_X1 U16122 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14905), .ZN(P2_U3275) );
  AND2_X1 U16123 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14905), .ZN(P2_U3274) );
  AND2_X1 U16124 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14905), .ZN(P2_U3273) );
  AND2_X1 U16125 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14905), .ZN(P2_U3272) );
  AND2_X1 U16126 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14905), .ZN(P2_U3271) );
  AND2_X1 U16127 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14905), .ZN(P2_U3270) );
  AND2_X1 U16128 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14905), .ZN(P2_U3269) );
  AND2_X1 U16129 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14905), .ZN(P2_U3268) );
  AND2_X1 U16130 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14905), .ZN(P2_U3267) );
  AND2_X1 U16131 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14905), .ZN(P2_U3266) );
  NOR2_X1 U16132 ( .A1(n15200), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16133 ( .A1(P3_U3897), .A2(n15502), .ZN(P3_U3150) );
  OAI22_X1 U16134 ( .A1(n15121), .A2(keyinput_126), .B1(n15118), .B2(
        keyinput_127), .ZN(n14906) );
  AOI221_X1 U16135 ( .B1(n15121), .B2(keyinput_126), .C1(keyinput_127), .C2(
        n15118), .A(n14906), .ZN(n15003) );
  INV_X1 U16136 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15117) );
  INV_X1 U16137 ( .A(keyinput_124), .ZN(n15001) );
  INV_X1 U16138 ( .A(keyinput_123), .ZN(n14999) );
  OAI22_X1 U16139 ( .A1(n9823), .A2(keyinput_120), .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .ZN(n14907) );
  AOI221_X1 U16140 ( .B1(n9823), .B2(keyinput_120), .C1(keyinput_121), .C2(
        P3_REG3_REG_22__SCAN_IN), .A(n14907), .ZN(n14996) );
  INV_X1 U16141 ( .A(keyinput_119), .ZN(n14994) );
  INV_X1 U16142 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15105) );
  INV_X1 U16143 ( .A(keyinput_118), .ZN(n14992) );
  INV_X1 U16144 ( .A(keyinput_109), .ZN(n14978) );
  INV_X1 U16145 ( .A(keyinput_108), .ZN(n14976) );
  INV_X1 U16146 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15092) );
  INV_X1 U16147 ( .A(keyinput_107), .ZN(n14974) );
  INV_X1 U16148 ( .A(keyinput_100), .ZN(n14964) );
  AOI22_X1 U16149 ( .A1(SI_4_), .A2(keyinput_92), .B1(SI_5_), .B2(keyinput_91), 
        .ZN(n14908) );
  OAI221_X1 U16150 ( .B1(SI_4_), .B2(keyinput_92), .C1(SI_5_), .C2(keyinput_91), .A(n14908), .ZN(n14917) );
  XOR2_X1 U16151 ( .A(n14909), .B(keyinput_86), .Z(n14916) );
  XNOR2_X1 U16152 ( .A(n14910), .B(keyinput_87), .ZN(n14914) );
  XNOR2_X1 U16153 ( .A(SI_8_), .B(keyinput_88), .ZN(n14913) );
  XNOR2_X1 U16154 ( .A(SI_7_), .B(keyinput_89), .ZN(n14912) );
  XNOR2_X1 U16155 ( .A(SI_6_), .B(keyinput_90), .ZN(n14911) );
  NAND4_X1 U16156 ( .A1(n14914), .A2(n14913), .A3(n14912), .A4(n14911), .ZN(
        n14915) );
  NOR3_X1 U16157 ( .A1(n14917), .A2(n14916), .A3(n14915), .ZN(n14962) );
  INV_X1 U16158 ( .A(keyinput_85), .ZN(n14950) );
  INV_X1 U16159 ( .A(keyinput_84), .ZN(n14948) );
  INV_X1 U16160 ( .A(keyinput_79), .ZN(n14940) );
  INV_X1 U16161 ( .A(keyinput_78), .ZN(n14938) );
  INV_X1 U16162 ( .A(SI_28_), .ZN(n14919) );
  OAI22_X1 U16163 ( .A1(n14919), .A2(keyinput_68), .B1(keyinput_69), .B2(
        SI_27_), .ZN(n14918) );
  AOI221_X1 U16164 ( .B1(n14919), .B2(keyinput_68), .C1(SI_27_), .C2(
        keyinput_69), .A(n14918), .ZN(n14936) );
  INV_X1 U16165 ( .A(keyinput_67), .ZN(n14924) );
  INV_X1 U16166 ( .A(keyinput_66), .ZN(n14922) );
  AOI22_X1 U16167 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n14920) );
  OAI221_X1 U16168 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n14920), .ZN(n14921) );
  OAI221_X1 U16169 ( .B1(SI_30_), .B2(n14922), .C1(n15023), .C2(keyinput_66), 
        .A(n14921), .ZN(n14923) );
  OAI221_X1 U16170 ( .B1(SI_29_), .B2(n14924), .C1(n15026), .C2(keyinput_67), 
        .A(n14923), .ZN(n14935) );
  OAI22_X1 U16171 ( .A1(n15017), .A2(keyinput_71), .B1(n11068), .B2(
        keyinput_76), .ZN(n14925) );
  AOI221_X1 U16172 ( .B1(n15017), .B2(keyinput_71), .C1(keyinput_76), .C2(
        n11068), .A(n14925), .ZN(n14933) );
  OAI22_X1 U16173 ( .A1(n14927), .A2(keyinput_70), .B1(n15020), .B2(
        keyinput_77), .ZN(n14926) );
  AOI221_X1 U16174 ( .B1(n14927), .B2(keyinput_70), .C1(keyinput_77), .C2(
        n15020), .A(n14926), .ZN(n14932) );
  OAI22_X1 U16175 ( .A1(SI_24_), .A2(keyinput_72), .B1(SI_21_), .B2(
        keyinput_75), .ZN(n14928) );
  AOI221_X1 U16176 ( .B1(SI_24_), .B2(keyinput_72), .C1(keyinput_75), .C2(
        SI_21_), .A(n14928), .ZN(n14931) );
  OAI22_X1 U16177 ( .A1(n15019), .A2(keyinput_74), .B1(keyinput_73), .B2(
        SI_23_), .ZN(n14929) );
  AOI221_X1 U16178 ( .B1(n15019), .B2(keyinput_74), .C1(SI_23_), .C2(
        keyinput_73), .A(n14929), .ZN(n14930) );
  NAND4_X1 U16179 ( .A1(n14933), .A2(n14932), .A3(n14931), .A4(n14930), .ZN(
        n14934) );
  AOI21_X1 U16180 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14937) );
  AOI221_X1 U16181 ( .B1(SI_18_), .B2(n14938), .C1(n15041), .C2(keyinput_78), 
        .A(n14937), .ZN(n14939) );
  AOI221_X1 U16182 ( .B1(SI_17_), .B2(keyinput_79), .C1(n15044), .C2(n14940), 
        .A(n14939), .ZN(n14946) );
  AOI22_X1 U16183 ( .A1(n15047), .A2(keyinput_80), .B1(keyinput_81), .B2(
        n15046), .ZN(n14941) );
  OAI221_X1 U16184 ( .B1(n15047), .B2(keyinput_80), .C1(n15046), .C2(
        keyinput_81), .A(n14941), .ZN(n14945) );
  OAI22_X1 U16185 ( .A1(n14943), .A2(keyinput_82), .B1(keyinput_83), .B2(
        SI_13_), .ZN(n14942) );
  AOI221_X1 U16186 ( .B1(n14943), .B2(keyinput_82), .C1(SI_13_), .C2(
        keyinput_83), .A(n14942), .ZN(n14944) );
  OAI21_X1 U16187 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14947) );
  OAI221_X1 U16188 ( .B1(SI_12_), .B2(n14948), .C1(n15053), .C2(keyinput_84), 
        .A(n14947), .ZN(n14949) );
  OAI221_X1 U16189 ( .B1(SI_11_), .B2(n14950), .C1(n15057), .C2(keyinput_85), 
        .A(n14949), .ZN(n14961) );
  AOI22_X1 U16190 ( .A1(SI_0_), .A2(keyinput_96), .B1(P3_REG3_REG_7__SCAN_IN), 
        .B2(keyinput_99), .ZN(n14951) );
  OAI221_X1 U16191 ( .B1(SI_0_), .B2(keyinput_96), .C1(P3_REG3_REG_7__SCAN_IN), 
        .C2(keyinput_99), .A(n14951), .ZN(n14960) );
  INV_X1 U16192 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15525) );
  XOR2_X1 U16193 ( .A(keyinput_97), .B(n15525), .Z(n14957) );
  XNOR2_X1 U16194 ( .A(n15075), .B(keyinput_94), .ZN(n14952) );
  AOI21_X1 U16195 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_98), .A(n14952), 
        .ZN(n14956) );
  XNOR2_X1 U16196 ( .A(n14953), .B(keyinput_95), .ZN(n14955) );
  XNOR2_X1 U16197 ( .A(SI_3_), .B(keyinput_93), .ZN(n14954) );
  AND4_X1 U16198 ( .A1(n14957), .A2(n14956), .A3(n14955), .A4(n14954), .ZN(
        n14958) );
  OAI21_X1 U16199 ( .B1(keyinput_98), .B2(P3_STATE_REG_SCAN_IN), .A(n14958), 
        .ZN(n14959) );
  AOI211_X1 U16200 ( .C1(n14962), .C2(n14961), .A(n14960), .B(n14959), .ZN(
        n14963) );
  AOI221_X1 U16201 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(n14964), .C1(n15083), 
        .C2(keyinput_100), .A(n14963), .ZN(n14972) );
  AOI22_X1 U16202 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_102), .B1(
        n12794), .B2(keyinput_105), .ZN(n14965) );
  OAI221_X1 U16203 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .C1(
        n12794), .C2(keyinput_105), .A(n14965), .ZN(n14971) );
  AOI22_X1 U16204 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(
        n15013), .B2(keyinput_104), .ZN(n14966) );
  OAI221_X1 U16205 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        n15013), .C2(keyinput_104), .A(n14966), .ZN(n14970) );
  INV_X1 U16206 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U16207 ( .A1(n12806), .A2(keyinput_106), .B1(keyinput_103), .B2(
        n14968), .ZN(n14967) );
  OAI221_X1 U16208 ( .B1(n12806), .B2(keyinput_106), .C1(n14968), .C2(
        keyinput_103), .A(n14967), .ZN(n14969) );
  NOR4_X1 U16209 ( .A1(n14972), .A2(n14971), .A3(n14970), .A4(n14969), .ZN(
        n14973) );
  AOI221_X1 U16210 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n15090), .C2(n14974), .A(n14973), .ZN(n14975) );
  AOI221_X1 U16211 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n14976), .C1(n15092), 
        .C2(keyinput_108), .A(n14975), .ZN(n14977) );
  AOI221_X1 U16212 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        n15096), .C2(n14978), .A(n14977), .ZN(n14990) );
  INV_X1 U16213 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n14981) );
  INV_X1 U16214 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n14980) );
  AOI22_X1 U16215 ( .A1(n14981), .A2(keyinput_111), .B1(keyinput_110), .B2(
        n14980), .ZN(n14979) );
  OAI221_X1 U16216 ( .B1(n14981), .B2(keyinput_111), .C1(n14980), .C2(
        keyinput_110), .A(n14979), .ZN(n14984) );
  AOI22_X1 U16217 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_114), .B1(n9696), .B2(keyinput_113), .ZN(n14982) );
  OAI221_X1 U16218 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        n9696), .C2(keyinput_113), .A(n14982), .ZN(n14983) );
  AOI211_X1 U16219 ( .C1(keyinput_112), .C2(P3_REG3_REG_16__SCAN_IN), .A(
        n14984), .B(n14983), .ZN(n14985) );
  OAI21_X1 U16220 ( .B1(keyinput_112), .B2(P3_REG3_REG_16__SCAN_IN), .A(n14985), .ZN(n14989) );
  OAI22_X1 U16221 ( .A1(n15098), .A2(keyinput_116), .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .ZN(n14986) );
  AOI221_X1 U16222 ( .B1(n15098), .B2(keyinput_116), .C1(keyinput_117), .C2(
        P3_REG3_REG_9__SCAN_IN), .A(n14986), .ZN(n14988) );
  XNOR2_X1 U16223 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n14987)
         );
  OAI211_X1 U16224 ( .C1(n14990), .C2(n14989), .A(n14988), .B(n14987), .ZN(
        n14991) );
  OAI221_X1 U16225 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(
        n15105), .C2(n14992), .A(n14991), .ZN(n14993) );
  OAI221_X1 U16226 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        n15108), .C2(n14994), .A(n14993), .ZN(n14995) );
  AOI22_X1 U16227 ( .A1(n14996), .A2(n14995), .B1(keyinput_122), .B2(
        P3_REG3_REG_11__SCAN_IN), .ZN(n14997) );
  OAI21_X1 U16228 ( .B1(keyinput_122), .B2(P3_REG3_REG_11__SCAN_IN), .A(n14997), .ZN(n14998) );
  OAI221_X1 U16229 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(
        n10926), .C2(n14999), .A(n14998), .ZN(n15000) );
  OAI221_X1 U16230 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        n15117), .C2(n15001), .A(n15000), .ZN(n15002) );
  OAI211_X1 U16231 ( .C1(P3_REG3_REG_6__SCAN_IN), .C2(keyinput_125), .A(n15003), .B(n15002), .ZN(n15004) );
  AOI21_X1 U16232 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .A(n15004), 
        .ZN(n15125) );
  INV_X1 U16233 ( .A(keyinput_60), .ZN(n15116) );
  INV_X1 U16234 ( .A(keyinput_59), .ZN(n15114) );
  INV_X1 U16235 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U16236 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .ZN(n15005) );
  OAI221_X1 U16237 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n15005), .ZN(n15110) );
  INV_X1 U16238 ( .A(keyinput_55), .ZN(n15107) );
  INV_X1 U16239 ( .A(keyinput_54), .ZN(n15104) );
  OAI22_X1 U16240 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_48), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .ZN(n15006) );
  AOI221_X1 U16241 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(
        keyinput_46), .C2(P3_REG3_REG_12__SCAN_IN), .A(n15006), .ZN(n15009) );
  OAI22_X1 U16242 ( .A1(n9696), .A2(keyinput_49), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(keyinput_47), .ZN(n15007) );
  AOI221_X1 U16243 ( .B1(n9696), .B2(keyinput_49), .C1(keyinput_47), .C2(
        P3_REG3_REG_25__SCAN_IN), .A(n15007), .ZN(n15008) );
  OAI211_X1 U16244 ( .C1(P3_REG3_REG_17__SCAN_IN), .C2(keyinput_50), .A(n15009), .B(n15008), .ZN(n15010) );
  AOI21_X1 U16245 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .A(n15010), 
        .ZN(n15102) );
  INV_X1 U16246 ( .A(keyinput_45), .ZN(n15095) );
  INV_X1 U16247 ( .A(keyinput_44), .ZN(n15093) );
  INV_X1 U16248 ( .A(keyinput_43), .ZN(n15089) );
  OAI22_X1 U16249 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .ZN(n15011) );
  AOI221_X1 U16250 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        keyinput_39), .C2(P3_REG3_REG_10__SCAN_IN), .A(n15011), .ZN(n15087) );
  OAI22_X1 U16251 ( .A1(n12794), .A2(keyinput_41), .B1(n15013), .B2(
        keyinput_40), .ZN(n15012) );
  AOI221_X1 U16252 ( .B1(n12794), .B2(keyinput_41), .C1(keyinput_40), .C2(
        n15013), .A(n15012), .ZN(n15086) );
  OAI22_X1 U16253 ( .A1(n12806), .A2(keyinput_42), .B1(n15015), .B2(
        keyinput_38), .ZN(n15014) );
  AOI221_X1 U16254 ( .B1(n12806), .B2(keyinput_42), .C1(keyinput_38), .C2(
        n15015), .A(n15014), .ZN(n15085) );
  INV_X1 U16255 ( .A(keyinput_36), .ZN(n15082) );
  INV_X1 U16256 ( .A(keyinput_21), .ZN(n15056) );
  INV_X1 U16257 ( .A(keyinput_20), .ZN(n15054) );
  INV_X1 U16258 ( .A(keyinput_15), .ZN(n15043) );
  INV_X1 U16259 ( .A(keyinput_14), .ZN(n15040) );
  AOI22_X1 U16260 ( .A1(SI_24_), .A2(keyinput_8), .B1(n15017), .B2(keyinput_7), 
        .ZN(n15016) );
  OAI221_X1 U16261 ( .B1(SI_24_), .B2(keyinput_8), .C1(n15017), .C2(keyinput_7), .A(n15016), .ZN(n15038) );
  AOI22_X1 U16262 ( .A1(n15020), .A2(keyinput_13), .B1(n15019), .B2(
        keyinput_10), .ZN(n15018) );
  OAI221_X1 U16263 ( .B1(n15020), .B2(keyinput_13), .C1(n15019), .C2(
        keyinput_10), .A(n15018), .ZN(n15037) );
  INV_X1 U16264 ( .A(keyinput_3), .ZN(n15027) );
  INV_X1 U16265 ( .A(keyinput_2), .ZN(n15024) );
  OAI22_X1 U16266 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15021) );
  AOI221_X1 U16267 ( .B1(SI_31_), .B2(keyinput_1), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n15021), .ZN(n15022) );
  AOI221_X1 U16268 ( .B1(SI_30_), .B2(n15024), .C1(n15023), .C2(keyinput_2), 
        .A(n15022), .ZN(n15025) );
  AOI221_X1 U16269 ( .B1(SI_29_), .B2(n15027), .C1(n15026), .C2(keyinput_3), 
        .A(n15025), .ZN(n15035) );
  AOI22_X1 U16270 ( .A1(SI_28_), .A2(keyinput_4), .B1(n15029), .B2(keyinput_5), 
        .ZN(n15028) );
  OAI221_X1 U16271 ( .B1(SI_28_), .B2(keyinput_4), .C1(n15029), .C2(keyinput_5), .A(n15028), .ZN(n15034) );
  OAI22_X1 U16272 ( .A1(SI_26_), .A2(keyinput_6), .B1(keyinput_11), .B2(SI_21_), .ZN(n15030) );
  AOI221_X1 U16273 ( .B1(SI_26_), .B2(keyinput_6), .C1(SI_21_), .C2(
        keyinput_11), .A(n15030), .ZN(n15033) );
  OAI22_X1 U16274 ( .A1(SI_23_), .A2(keyinput_9), .B1(SI_20_), .B2(keyinput_12), .ZN(n15031) );
  AOI221_X1 U16275 ( .B1(SI_23_), .B2(keyinput_9), .C1(keyinput_12), .C2(
        SI_20_), .A(n15031), .ZN(n15032) );
  OAI211_X1 U16276 ( .C1(n15035), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        n15036) );
  NOR3_X1 U16277 ( .A1(n15038), .A2(n15037), .A3(n15036), .ZN(n15039) );
  AOI221_X1 U16278 ( .B1(SI_18_), .B2(keyinput_14), .C1(n15041), .C2(n15040), 
        .A(n15039), .ZN(n15042) );
  AOI221_X1 U16279 ( .B1(SI_17_), .B2(keyinput_15), .C1(n15044), .C2(n15043), 
        .A(n15042), .ZN(n15051) );
  AOI22_X1 U16280 ( .A1(n15047), .A2(keyinput_16), .B1(keyinput_17), .B2(
        n15046), .ZN(n15045) );
  OAI221_X1 U16281 ( .B1(n15047), .B2(keyinput_16), .C1(n15046), .C2(
        keyinput_17), .A(n15045), .ZN(n15050) );
  OAI22_X1 U16282 ( .A1(SI_14_), .A2(keyinput_18), .B1(keyinput_19), .B2(
        SI_13_), .ZN(n15048) );
  AOI221_X1 U16283 ( .B1(SI_14_), .B2(keyinput_18), .C1(SI_13_), .C2(
        keyinput_19), .A(n15048), .ZN(n15049) );
  OAI21_X1 U16284 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n15052) );
  OAI221_X1 U16285 ( .B1(SI_12_), .B2(n15054), .C1(n15053), .C2(keyinput_20), 
        .A(n15052), .ZN(n15055) );
  OAI221_X1 U16286 ( .B1(SI_11_), .B2(keyinput_21), .C1(n15057), .C2(n15056), 
        .A(n15055), .ZN(n15074) );
  AOI22_X1 U16287 ( .A1(SI_5_), .A2(keyinput_27), .B1(SI_10_), .B2(keyinput_22), .ZN(n15058) );
  OAI221_X1 U16288 ( .B1(SI_5_), .B2(keyinput_27), .C1(SI_10_), .C2(
        keyinput_22), .A(n15058), .ZN(n15066) );
  XOR2_X1 U16289 ( .A(SI_8_), .B(keyinput_24), .Z(n15061) );
  XNOR2_X1 U16290 ( .A(SI_6_), .B(keyinput_26), .ZN(n15060) );
  XNOR2_X1 U16291 ( .A(SI_4_), .B(keyinput_28), .ZN(n15059) );
  NAND3_X1 U16292 ( .A1(n15061), .A2(n15060), .A3(n15059), .ZN(n15065) );
  XNOR2_X1 U16293 ( .A(n15062), .B(keyinput_25), .ZN(n15064) );
  XNOR2_X1 U16294 ( .A(SI_9_), .B(keyinput_23), .ZN(n15063) );
  NOR4_X1 U16295 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        n15073) );
  INV_X1 U16296 ( .A(SI_0_), .ZN(n15067) );
  XOR2_X1 U16297 ( .A(n15067), .B(keyinput_32), .Z(n15071) );
  XNOR2_X1 U16298 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n15070) );
  XNOR2_X1 U16299 ( .A(SI_1_), .B(keyinput_31), .ZN(n15069) );
  XNOR2_X1 U16300 ( .A(SI_3_), .B(keyinput_29), .ZN(n15068) );
  NAND4_X1 U16301 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15072) );
  AOI21_X1 U16302 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15079) );
  XNOR2_X1 U16303 ( .A(n15075), .B(keyinput_30), .ZN(n15077) );
  XNOR2_X1 U16304 ( .A(n15525), .B(keyinput_33), .ZN(n15076) );
  AOI211_X1 U16305 ( .C1(keyinput_35), .C2(n15080), .A(n15077), .B(n15076), 
        .ZN(n15078) );
  OAI211_X1 U16306 ( .C1(keyinput_35), .C2(n15080), .A(n15079), .B(n15078), 
        .ZN(n15081) );
  OAI221_X1 U16307 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n15083), .C2(n15082), .A(n15081), .ZN(n15084) );
  NAND4_X1 U16308 ( .A1(n15087), .A2(n15086), .A3(n15085), .A4(n15084), .ZN(
        n15088) );
  OAI221_X1 U16309 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(n15090), .C2(n15089), .A(n15088), .ZN(n15091) );
  OAI221_X1 U16310 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n15093), .C1(n15092), 
        .C2(keyinput_44), .A(n15091), .ZN(n15094) );
  OAI221_X1 U16311 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        n15096), .C2(n15095), .A(n15094), .ZN(n15101) );
  XOR2_X1 U16312 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .Z(n15100) );
  AOI22_X1 U16313 ( .A1(n15098), .A2(keyinput_52), .B1(n9756), .B2(keyinput_53), .ZN(n15097) );
  OAI221_X1 U16314 ( .B1(n15098), .B2(keyinput_52), .C1(n9756), .C2(
        keyinput_53), .A(n15097), .ZN(n15099) );
  AOI211_X1 U16315 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15103) );
  AOI221_X1 U16316 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n15105), .C2(n15104), .A(n15103), .ZN(n15106) );
  AOI221_X1 U16317 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        n15108), .C2(n15107), .A(n15106), .ZN(n15109) );
  OAI22_X1 U16318 ( .A1(keyinput_58), .A2(n15112), .B1(n15110), .B2(n15109), 
        .ZN(n15111) );
  AOI21_X1 U16319 ( .B1(keyinput_58), .B2(n15112), .A(n15111), .ZN(n15113) );
  AOI221_X1 U16320 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n15114), .C1(n10926), 
        .C2(keyinput_59), .A(n15113), .ZN(n15115) );
  AOI221_X1 U16321 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        n15117), .C2(n15116), .A(n15115), .ZN(n15124) );
  XOR2_X1 U16322 ( .A(n15118), .B(keyinput_63), .Z(n15123) );
  AOI22_X1 U16323 ( .A1(n15121), .A2(keyinput_62), .B1(keyinput_61), .B2(
        n15120), .ZN(n15119) );
  OAI221_X1 U16324 ( .B1(n15121), .B2(keyinput_62), .C1(n15120), .C2(
        keyinput_61), .A(n15119), .ZN(n15122) );
  NOR4_X1 U16325 ( .A1(n15125), .A2(n15124), .A3(n15123), .A4(n15122), .ZN(
        n15136) );
  OAI22_X1 U16326 ( .A1(n15128), .A2(n15127), .B1(n9652), .B2(n15126), .ZN(
        n15129) );
  AOI21_X1 U16327 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15134) );
  OR2_X1 U16328 ( .A1(n15132), .A2(n15105), .ZN(n15133) );
  AND2_X1 U16329 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  XNOR2_X1 U16330 ( .A(n15136), .B(n15135), .ZN(P3_U3172) );
  AOI22_X1 U16331 ( .A1(n15140), .A2(n15139), .B1(n15138), .B2(n15137), .ZN(
        P2_U3416) );
  INV_X1 U16332 ( .A(n15141), .ZN(n15143) );
  OAI21_X1 U16333 ( .B1(n15143), .B2(n15142), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15144) );
  OAI21_X1 U16334 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15144), .ZN(n15155) );
  OAI211_X1 U16335 ( .C1(n15147), .C2(n15146), .A(n15201), .B(n15145), .ZN(
        n15154) );
  AOI211_X1 U16336 ( .C1(n15150), .C2(n15149), .A(n15148), .B(n15180), .ZN(
        n15151) );
  INV_X1 U16337 ( .A(n15151), .ZN(n15153) );
  NAND2_X1 U16338 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n15200), .ZN(n15152) );
  NAND4_X1 U16339 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        P2_U3220) );
  OAI21_X1 U16340 ( .B1(n15158), .B2(n15157), .A(n15156), .ZN(n15159) );
  AOI21_X1 U16341 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15200), .A(n15159), 
        .ZN(n15166) );
  OAI211_X1 U16342 ( .C1(n15161), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15205), 
        .B(n15160), .ZN(n15165) );
  OAI211_X1 U16343 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15163), .A(n15201), 
        .B(n15162), .ZN(n15164) );
  NAND3_X1 U16344 ( .A1(n15166), .A2(n15165), .A3(n15164), .ZN(P2_U3229) );
  INV_X1 U16345 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15356) );
  OAI21_X1 U16346 ( .B1(n15168), .B2(n12376), .A(n15167), .ZN(n15169) );
  INV_X1 U16347 ( .A(n15169), .ZN(n15170) );
  OAI21_X1 U16348 ( .B1(n15170), .B2(n15186), .A(n15189), .ZN(n15171) );
  NOR2_X1 U16349 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15171), .ZN(n15190) );
  AOI21_X1 U16350 ( .B1(n15171), .B2(P2_REG2_REG_18__SCAN_IN), .A(n15190), 
        .ZN(n15179) );
  NAND2_X1 U16351 ( .A1(n15210), .A2(n15175), .ZN(n15178) );
  INV_X1 U16352 ( .A(n15172), .ZN(n15173) );
  AOI21_X1 U16353 ( .B1(n15174), .B2(P2_REG1_REG_17__SCAN_IN), .A(n15173), 
        .ZN(n15185) );
  XNOR2_X1 U16354 ( .A(n15175), .B(n15185), .ZN(n15176) );
  NAND2_X1 U16355 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n15176), .ZN(n15184) );
  OAI211_X1 U16356 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n15176), .A(n15201), 
        .B(n15184), .ZN(n15177) );
  OAI211_X1 U16357 ( .C1(n15180), .C2(n15179), .A(n15178), .B(n15177), .ZN(
        n15181) );
  INV_X1 U16358 ( .A(n15181), .ZN(n15183) );
  OAI211_X1 U16359 ( .C1(n15356), .C2(n15198), .A(n15183), .B(n15182), .ZN(
        P2_U3232) );
  XNOR2_X1 U16360 ( .A(n15194), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n15188) );
  OAI21_X1 U16361 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15187) );
  XNOR2_X1 U16362 ( .A(n15188), .B(n15187), .ZN(n15196) );
  INV_X1 U16363 ( .A(n15189), .ZN(n15191) );
  XNOR2_X1 U16364 ( .A(n15194), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n15192) );
  XNOR2_X1 U16365 ( .A(n15193), .B(n15192), .ZN(n15195) );
  AOI22_X1 U16366 ( .A1(n15200), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15214) );
  OAI211_X1 U16367 ( .C1(n15204), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15213) );
  OAI211_X1 U16368 ( .C1(n15208), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n15212) );
  NAND2_X1 U16369 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  NAND4_X1 U16370 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        P2_U3227) );
  AOI21_X1 U16371 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15380), .A(n15217), .ZN(
        n15216) );
  INV_X1 U16372 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15215) );
  NOR2_X1 U16373 ( .A1(n15216), .A2(n15215), .ZN(n15371) );
  AOI21_X1 U16374 ( .B1(n15216), .B2(n15215), .A(n15371), .ZN(SUB_1596_U53) );
  INV_X1 U16375 ( .A(n15217), .ZN(n15221) );
  NAND2_X1 U16376 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15218), .ZN(n15219) );
  XNOR2_X1 U16377 ( .A(n15226), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n15223) );
  XNOR2_X1 U16378 ( .A(n15224), .B(n15223), .ZN(n15228) );
  NOR2_X1 U16379 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  AOI21_X1 U16380 ( .B1(n15227), .B2(n15228), .A(n15229), .ZN(n15222) );
  XOR2_X1 U16381 ( .A(n15222), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  NOR2_X1 U16382 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  XNOR2_X1 U16383 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15232), .ZN(n15233) );
  NAND2_X1 U16384 ( .A1(n15228), .A2(n15227), .ZN(n15230) );
  XNOR2_X1 U16385 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15235), .ZN(SUB_1596_U60)
         );
  XNOR2_X1 U16386 ( .A(n15240), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n15237) );
  XNOR2_X1 U16387 ( .A(n15238), .B(n15237), .ZN(n15242) );
  NOR2_X1 U16388 ( .A1(n15234), .A2(n15233), .ZN(n15236) );
  XOR2_X1 U16389 ( .A(n15244), .B(n15243), .Z(SUB_1596_U59) );
  XOR2_X1 U16390 ( .A(n15250), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n15241) );
  NOR2_X1 U16391 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  XOR2_X1 U16392 ( .A(n15241), .B(n15252), .Z(n15247) );
  NAND2_X1 U16393 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15242), .ZN(n15245) );
  XOR2_X1 U16394 ( .A(n15248), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  NAND2_X1 U16395 ( .A1(n15247), .A2(n15246), .ZN(n15249) );
  XOR2_X1 U16396 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(n15254), .Z(n15253) );
  XNOR2_X1 U16397 ( .A(n15253), .B(n15255), .ZN(n15367) );
  INV_X1 U16398 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15369) );
  AND2_X1 U16399 ( .A1(n15254), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n15256) );
  XOR2_X1 U16400 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15261), .Z(n15263) );
  XNOR2_X1 U16401 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15263), .ZN(n15258) );
  XOR2_X1 U16402 ( .A(n15259), .B(n15258), .Z(SUB_1596_U56) );
  NAND2_X1 U16403 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15257), .ZN(n15260) );
  XOR2_X1 U16404 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n15273), .Z(n15271) );
  INV_X1 U16405 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15262) );
  NOR2_X1 U16406 ( .A1(n15262), .A2(n15261), .ZN(n15265) );
  XOR2_X1 U16407 ( .A(n15271), .B(n15270), .Z(n15267) );
  XOR2_X1 U16408 ( .A(n15268), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  NAND2_X1 U16409 ( .A1(n15267), .A2(n15266), .ZN(n15269) );
  NAND2_X1 U16410 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  XOR2_X1 U16411 ( .A(n15399), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n15276) );
  XOR2_X1 U16412 ( .A(n15275), .B(n15276), .Z(n15279) );
  NAND2_X1 U16413 ( .A1(n15279), .A2(n15278), .ZN(n15280) );
  OAI21_X1 U16414 ( .B1(n15278), .B2(n15279), .A(n15280), .ZN(n15274) );
  INV_X1 U16415 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15281) );
  XOR2_X1 U16416 ( .A(n15274), .B(n15281), .Z(SUB_1596_U54) );
  INV_X1 U16417 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15418) );
  INV_X1 U16418 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15292) );
  XNOR2_X1 U16419 ( .A(n15418), .B(n15292), .ZN(n15289) );
  XNOR2_X1 U16420 ( .A(n15290), .B(n15289), .ZN(n15285) );
  NOR2_X1 U16421 ( .A1(n15279), .A2(n15278), .ZN(n15282) );
  OAI21_X1 U16422 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15284) );
  NAND2_X1 U16423 ( .A1(n15285), .A2(n15284), .ZN(n15286) );
  OAI21_X1 U16424 ( .B1(n15285), .B2(n15284), .A(n15286), .ZN(n15283) );
  INV_X1 U16425 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15287) );
  XOR2_X1 U16426 ( .A(n15283), .B(n15287), .Z(SUB_1596_U70) );
  NOR2_X1 U16427 ( .A1(n15285), .A2(n15284), .ZN(n15288) );
  INV_X1 U16428 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15297) );
  XOR2_X1 U16429 ( .A(n15297), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n15293) );
  XOR2_X1 U16430 ( .A(n15293), .B(n15299), .Z(n15295) );
  XNOR2_X1 U16431 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15296), .ZN(SUB_1596_U69)
         );
  INV_X1 U16432 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15307) );
  XOR2_X1 U16433 ( .A(n15307), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n15305) );
  OR2_X1 U16434 ( .A1(n15297), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n15298) );
  XNOR2_X1 U16435 ( .A(n15305), .B(n15304), .ZN(n15300) );
  XNOR2_X1 U16436 ( .A(n15301), .B(n15300), .ZN(n15302) );
  XNOR2_X1 U16437 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15302), .ZN(SUB_1596_U68)
         );
  NOR2_X1 U16438 ( .A1(n15301), .A2(n15300), .ZN(n15303) );
  XOR2_X1 U16439 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n15310) );
  NAND2_X1 U16440 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  NOR2_X1 U16441 ( .A1(n15313), .A2(n7339), .ZN(n15308) );
  XOR2_X1 U16442 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n15308), .Z(SUB_1596_U67)
         );
  INV_X1 U16443 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15312) );
  NOR2_X1 U16444 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  AOI21_X1 U16445 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n15312), .A(n15311), 
        .ZN(n15322) );
  XOR2_X1 U16446 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n15321) );
  XOR2_X1 U16447 ( .A(n15322), .B(n15321), .Z(n15315) );
  NOR2_X1 U16448 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  AOI21_X1 U16449 ( .B1(n15315), .B2(n15316), .A(n15317), .ZN(n15314) );
  XOR2_X1 U16450 ( .A(n15314), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NAND2_X1 U16451 ( .A1(n15316), .A2(n15315), .ZN(n15318) );
  AOI21_X1 U16452 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(n15331) );
  INV_X1 U16453 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U16454 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15329), .ZN(n15320) );
  AOI21_X1 U16455 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15329), .A(n15320), 
        .ZN(n15327) );
  INV_X1 U16456 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15324) );
  NOR2_X1 U16457 ( .A1(n15322), .A2(n15321), .ZN(n15323) );
  AOI21_X1 U16458 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15324), .A(n15323), 
        .ZN(n15326) );
  XNOR2_X1 U16459 ( .A(n15327), .B(n15326), .ZN(n15330) );
  AOI21_X1 U16460 ( .B1(n15331), .B2(n15330), .A(n15332), .ZN(n15325) );
  XOR2_X1 U16461 ( .A(n15325), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  NAND2_X1 U16462 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  XOR2_X1 U16463 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15340), .Z(n15341) );
  XOR2_X1 U16464 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15341), .Z(n15334) );
  NOR2_X1 U16465 ( .A1(n15334), .A2(n15333), .ZN(n15338) );
  NOR2_X1 U16466 ( .A1(n15338), .A2(n15336), .ZN(n15335) );
  XOR2_X1 U16467 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15335), .Z(SUB_1596_U64)
         );
  NOR2_X1 U16468 ( .A1(n15338), .A2(n15337), .ZN(n15346) );
  INV_X1 U16469 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16470 ( .A1(n15340), .A2(n15339), .ZN(n15343) );
  NOR2_X1 U16471 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15341), .ZN(n15342) );
  NOR2_X1 U16472 ( .A1(n15343), .A2(n15342), .ZN(n15350) );
  XOR2_X1 U16473 ( .A(n15350), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n15351) );
  XOR2_X1 U16474 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15351), .Z(n15344) );
  XOR2_X1 U16475 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15344), .Z(n15345) );
  XOR2_X1 U16476 ( .A(n15346), .B(n15345), .Z(SUB_1596_U63) );
  NAND2_X1 U16477 ( .A1(n15344), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U16478 ( .A1(n15346), .A2(n15345), .ZN(n15347) );
  INV_X1 U16479 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16480 ( .A1(n15350), .A2(n15349), .ZN(n15353) );
  NOR2_X1 U16481 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15351), .ZN(n15352) );
  NOR2_X1 U16482 ( .A1(n15353), .A2(n15352), .ZN(n15361) );
  XOR2_X1 U16483 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n15360) );
  XOR2_X1 U16484 ( .A(n15361), .B(n15360), .Z(n15355) );
  NAND2_X1 U16485 ( .A1(n15355), .A2(n15354), .ZN(n15359) );
  NAND2_X1 U16486 ( .A1(n15358), .A2(n15359), .ZN(n15357) );
  XOR2_X1 U16487 ( .A(n15357), .B(n15356), .Z(SUB_1596_U62) );
  NOR2_X1 U16488 ( .A1(n15361), .A2(n15360), .ZN(n15362) );
  AOI21_X1 U16489 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13012), .A(n15362), 
        .ZN(n15364) );
  XNOR2_X1 U16490 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15363) );
  XNOR2_X1 U16491 ( .A(n15364), .B(n15363), .ZN(n15365) );
  OAI21_X1 U16492 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(n15370) );
  XOR2_X1 U16493 ( .A(n15370), .B(n15369), .Z(SUB_1596_U57) );
  XOR2_X1 U16494 ( .A(n15372), .B(n15371), .Z(SUB_1596_U5) );
  AOI22_X1 U16495 ( .A1(n15503), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15379) );
  NAND3_X1 U16496 ( .A1(n15500), .A2(n15373), .A3(n15460), .ZN(n15377) );
  OAI21_X1 U16497 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15375), .A(n15374), .ZN(
        n15376) );
  NAND2_X1 U16498 ( .A1(n15377), .A2(n15376), .ZN(n15378) );
  OAI211_X1 U16499 ( .C1(n15380), .C2(n15417), .A(n15379), .B(n15378), .ZN(
        P3_U3182) );
  INV_X1 U16500 ( .A(n15381), .ZN(n15382) );
  NAND2_X1 U16501 ( .A1(n15383), .A2(n15382), .ZN(n15384) );
  XNOR2_X1 U16502 ( .A(n15385), .B(n15384), .ZN(n15395) );
  OAI21_X1 U16503 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15387), .A(n15386), .ZN(
        n15389) );
  AOI22_X1 U16504 ( .A1(n15389), .A2(n15514), .B1(n15388), .B2(n15503), .ZN(
        n15394) );
  OAI21_X1 U16505 ( .B1(n15391), .B2(P3_REG2_REG_9__SCAN_IN), .A(n15390), .ZN(
        n15392) );
  NAND2_X1 U16506 ( .A1(n15392), .A2(n15517), .ZN(n15393) );
  OAI211_X1 U16507 ( .C1(n15395), .C2(n15460), .A(n15394), .B(n15393), .ZN(
        n15396) );
  INV_X1 U16508 ( .A(n15396), .ZN(n15398) );
  OAI211_X1 U16509 ( .C1(n15399), .C2(n15417), .A(n15398), .B(n15397), .ZN(
        P3_U3191) );
  AOI21_X1 U16510 ( .B1(n15401), .B2(n15400), .A(n7350), .ZN(n15413) );
  OAI21_X1 U16511 ( .B1(n15404), .B2(n15403), .A(n15402), .ZN(n15406) );
  AOI22_X1 U16512 ( .A1(n15406), .A2(n15517), .B1(n15405), .B2(n15503), .ZN(
        n15412) );
  OAI21_X1 U16513 ( .B1(n15409), .B2(n15408), .A(n15407), .ZN(n15410) );
  NAND2_X1 U16514 ( .A1(n15410), .A2(n15514), .ZN(n15411) );
  OAI211_X1 U16515 ( .C1(n15413), .C2(n15460), .A(n15412), .B(n15411), .ZN(
        n15414) );
  INV_X1 U16516 ( .A(n15414), .ZN(n15416) );
  OAI211_X1 U16517 ( .C1(n15418), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        P3_U3192) );
  AOI22_X1 U16518 ( .A1(n15503), .A2(n15419), .B1(n15502), .B2(
        P3_ADDR_REG_11__SCAN_IN), .ZN(n15432) );
  OAI21_X1 U16519 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n15421), .A(n15420), 
        .ZN(n15425) );
  OAI21_X1 U16520 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15423), .A(n15422), 
        .ZN(n15424) );
  AOI22_X1 U16521 ( .A1(n15517), .A2(n15425), .B1(n15424), .B2(n15514), .ZN(
        n15431) );
  AOI21_X1 U16522 ( .B1(n7344), .B2(n15427), .A(n15426), .ZN(n15428) );
  OR2_X1 U16523 ( .A1(n15428), .A2(n15460), .ZN(n15429) );
  NAND4_X1 U16524 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        P3_U3193) );
  INV_X1 U16525 ( .A(n15433), .ZN(n15434) );
  AOI22_X1 U16526 ( .A1(n15503), .A2(n15434), .B1(n15502), .B2(
        P3_ADDR_REG_12__SCAN_IN), .ZN(n15449) );
  OAI21_X1 U16527 ( .B1(n15437), .B2(n15436), .A(n15435), .ZN(n15442) );
  OAI21_X1 U16528 ( .B1(n15440), .B2(n15439), .A(n15438), .ZN(n15441) );
  AOI22_X1 U16529 ( .A1(n15517), .A2(n15442), .B1(n15441), .B2(n15514), .ZN(
        n15448) );
  OAI211_X1 U16530 ( .C1(n15445), .C2(n15444), .A(n15443), .B(n15515), .ZN(
        n15446) );
  NAND4_X1 U16531 ( .A1(n15449), .A2(n15448), .A3(n15447), .A4(n15446), .ZN(
        P3_U3194) );
  AOI22_X1 U16532 ( .A1(n15503), .A2(n15450), .B1(n15502), .B2(
        P3_ADDR_REG_13__SCAN_IN), .ZN(n15465) );
  OAI21_X1 U16533 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n15452), .A(n15451), 
        .ZN(n15456) );
  OAI21_X1 U16534 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15454), .A(n15453), 
        .ZN(n15455) );
  AOI22_X1 U16535 ( .A1(n15517), .A2(n15456), .B1(n15455), .B2(n15514), .ZN(
        n15464) );
  AOI21_X1 U16536 ( .B1(n15459), .B2(n15458), .A(n15457), .ZN(n15461) );
  OR2_X1 U16537 ( .A1(n15461), .A2(n15460), .ZN(n15462) );
  NAND4_X1 U16538 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        P3_U3195) );
  AOI22_X1 U16539 ( .A1(n15503), .A2(n15468), .B1(n15502), .B2(
        P3_ADDR_REG_14__SCAN_IN), .ZN(n15482) );
  OAI21_X1 U16540 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15469) );
  XOR2_X1 U16541 ( .A(n15470), .B(n15469), .Z(n15475) );
  OAI21_X1 U16542 ( .B1(n15473), .B2(n15472), .A(n15471), .ZN(n15474) );
  AOI22_X1 U16543 ( .A1(n15517), .A2(n15475), .B1(n15474), .B2(n15514), .ZN(
        n15481) );
  OAI211_X1 U16544 ( .C1(n15478), .C2(n15477), .A(n15476), .B(n15515), .ZN(
        n15479) );
  NAND4_X1 U16545 ( .A1(n15482), .A2(n15481), .A3(n15480), .A4(n15479), .ZN(
        P3_U3196) );
  AOI21_X1 U16546 ( .B1(n15485), .B2(n15484), .A(n15483), .ZN(n15501) );
  OAI21_X1 U16547 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n15487), .A(n15486), 
        .ZN(n15493) );
  AOI21_X1 U16548 ( .B1(n15502), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15488), 
        .ZN(n15489) );
  OAI21_X1 U16549 ( .B1(n15491), .B2(n15490), .A(n15489), .ZN(n15492) );
  AOI21_X1 U16550 ( .B1(n15493), .B2(n15514), .A(n15492), .ZN(n15499) );
  NOR2_X1 U16551 ( .A1(n15495), .A2(n15494), .ZN(n15496) );
  OAI21_X1 U16552 ( .B1(n15497), .B2(n15496), .A(n15515), .ZN(n15498) );
  OAI211_X1 U16553 ( .C1(n15501), .C2(n15500), .A(n15499), .B(n15498), .ZN(
        P3_U3197) );
  AOI22_X1 U16554 ( .A1(n15503), .A2(n15510), .B1(n15502), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U16555 ( .A1(n15505), .A2(n15504), .ZN(n15506) );
  XNOR2_X1 U16556 ( .A(n15507), .B(n15506), .ZN(n15516) );
  OAI21_X1 U16557 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n15511) );
  XOR2_X1 U16558 ( .A(n15512), .B(n15511), .Z(n15513) );
  AOI22_X1 U16559 ( .A1(n15516), .A2(n15515), .B1(n15514), .B2(n15513), .ZN(
        n15523) );
  NAND2_X1 U16560 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n15522)
         );
  OAI221_X1 U16561 ( .B1(n15520), .B2(n15519), .C1(n15520), .C2(n15518), .A(
        n15517), .ZN(n15521) );
  NAND4_X1 U16562 ( .A1(n15524), .A2(n15523), .A3(n15522), .A4(n15521), .ZN(
        P3_U3198) );
  OAI221_X1 U16563 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8155), .C2(n8153), .A(n15525), .ZN(U29) );
  INV_X1 U16564 ( .A(n15744), .ZN(n15777) );
  NAND2_X1 U16565 ( .A1(n15527), .A2(n15526), .ZN(n15535) );
  INV_X1 U16566 ( .A(n15535), .ZN(n15530) );
  OAI21_X1 U16567 ( .B1(n15749), .B2(n15914), .A(n15540), .ZN(n15528) );
  OAI21_X1 U16568 ( .B1(n15529), .B2(n15901), .A(n15528), .ZN(n15538) );
  AOI211_X1 U16569 ( .C1(n15777), .C2(n15540), .A(n15530), .B(n15538), .ZN(
        n15533) );
  AOI22_X1 U16570 ( .A1(n15717), .A2(n15533), .B1(n15531), .B2(n15924), .ZN(
        P1_U3528) );
  INV_X1 U16571 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U16572 ( .A1(n15719), .A2(n15533), .B1(n15532), .B2(n15926), .ZN(
        P1_U3459) );
  INV_X1 U16573 ( .A(n15534), .ZN(n15541) );
  AOI21_X1 U16574 ( .B1(n15537), .B2(n15536), .A(n15535), .ZN(n15539) );
  AOI211_X1 U16575 ( .C1(n15541), .C2(n15540), .A(n15539), .B(n15538), .ZN(
        n15543) );
  AOI22_X1 U16576 ( .A1(n15930), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n15941), .ZN(n15542) );
  OAI21_X1 U16577 ( .B1(n15941), .B2(n15543), .A(n15542), .ZN(P1_U3293) );
  XNOR2_X1 U16578 ( .A(n15549), .B(n15544), .ZN(n15559) );
  AOI22_X1 U16579 ( .A1(n15547), .A2(n10042), .B1(n15546), .B2(n15545), .ZN(
        n15552) );
  XNOR2_X1 U16580 ( .A(n15549), .B(n15548), .ZN(n15550) );
  NAND2_X1 U16581 ( .A1(n15550), .A2(n15577), .ZN(n15551) );
  OAI211_X1 U16582 ( .C1(n15559), .C2(n15733), .A(n15552), .B(n15551), .ZN(
        n15561) );
  OAI22_X1 U16583 ( .A1(n15559), .A2(n15732), .B1(n15553), .B2(n15797), .ZN(
        n15554) );
  NOR2_X1 U16584 ( .A1(n15561), .A2(n15554), .ZN(n15556) );
  INV_X1 U16585 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U16586 ( .A1(n15839), .A2(n15556), .B1(n15555), .B2(n15970), .ZN(
        P3_U3460) );
  AOI22_X1 U16587 ( .A1(n15980), .A2(n9640), .B1(n15556), .B2(n15978), .ZN(
        P3_U3393) );
  INV_X1 U16588 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U16589 ( .A1(n15680), .A2(P3_REG3_REG_1__SCAN_IN), .B1(n15585), 
        .B2(n15557), .ZN(n15558) );
  OAI21_X1 U16590 ( .B1(n15559), .B2(n15588), .A(n15558), .ZN(n15560) );
  NOR2_X1 U16591 ( .A1(n15561), .A2(n15560), .ZN(n15562) );
  AOI22_X1 U16592 ( .A1(n15690), .A2(n15563), .B1(n15562), .B2(n15688), .ZN(
        P3_U3232) );
  OAI21_X1 U16593 ( .B1(n15565), .B2(n15919), .A(n15564), .ZN(n15566) );
  AOI21_X1 U16594 ( .B1(n15567), .B2(n15923), .A(n15566), .ZN(n15568) );
  AND2_X1 U16595 ( .A1(n15569), .A2(n15568), .ZN(n15571) );
  AOI22_X1 U16596 ( .A1(n15717), .A2(n15571), .B1(n15570), .B2(n15924), .ZN(
        P1_U3529) );
  AOI22_X1 U16597 ( .A1(n15719), .A2(n15571), .B1(n8920), .B2(n15926), .ZN(
        P1_U3462) );
  XNOR2_X1 U16598 ( .A(n10163), .B(n15572), .ZN(n15589) );
  XNOR2_X1 U16599 ( .A(n15573), .B(n15572), .ZN(n15578) );
  OAI22_X1 U16600 ( .A1(n9652), .A2(n15575), .B1(n15574), .B2(n13243), .ZN(
        n15576) );
  AOI21_X1 U16601 ( .B1(n15578), .B2(n15577), .A(n15576), .ZN(n15579) );
  OAI21_X1 U16602 ( .B1(n15733), .B2(n15589), .A(n15579), .ZN(n15591) );
  OAI22_X1 U16603 ( .A1(n15589), .A2(n15732), .B1(n15797), .B2(n15580), .ZN(
        n15581) );
  NOR2_X1 U16604 ( .A1(n15591), .A2(n15581), .ZN(n15583) );
  INV_X1 U16605 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15582) );
  AOI22_X1 U16606 ( .A1(n15839), .A2(n15583), .B1(n15582), .B2(n15970), .ZN(
        P3_U3461) );
  INV_X1 U16607 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U16608 ( .A1(n15980), .A2(n15584), .B1(n15583), .B2(n15978), .ZN(
        P3_U3396) );
  AOI22_X1 U16609 ( .A1(n15680), .A2(P3_REG3_REG_2__SCAN_IN), .B1(n15586), 
        .B2(n15585), .ZN(n15587) );
  OAI21_X1 U16610 ( .B1(n15589), .B2(n15588), .A(n15587), .ZN(n15590) );
  NOR2_X1 U16611 ( .A1(n15591), .A2(n15590), .ZN(n15592) );
  AOI22_X1 U16612 ( .A1(n15690), .A2(n10809), .B1(n15592), .B2(n15688), .ZN(
        P3_U3231) );
  INV_X1 U16613 ( .A(n15599), .ZN(n15593) );
  NOR2_X1 U16614 ( .A1(n15593), .A2(n15744), .ZN(n15598) );
  OAI211_X1 U16615 ( .C1(n15596), .C2(n15919), .A(n15595), .B(n15594), .ZN(
        n15597) );
  AOI211_X1 U16616 ( .C1(n15599), .C2(n15749), .A(n15598), .B(n15597), .ZN(
        n15602) );
  AOI22_X1 U16617 ( .A1(n15717), .A2(n15602), .B1(n15600), .B2(n15924), .ZN(
        P1_U3530) );
  INV_X1 U16618 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U16619 ( .A1(n15719), .A2(n15602), .B1(n15601), .B2(n15926), .ZN(
        P1_U3465) );
  OAI21_X1 U16620 ( .B1(n15604), .B2(n15753), .A(n15603), .ZN(n15607) );
  INV_X1 U16621 ( .A(n15605), .ZN(n15606) );
  AOI211_X1 U16622 ( .C1(n15758), .C2(n15608), .A(n15607), .B(n15606), .ZN(
        n15610) );
  AOI22_X1 U16623 ( .A1(n15869), .A2(n15610), .B1(n10588), .B2(n15868), .ZN(
        P2_U3501) );
  INV_X1 U16624 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15609) );
  AOI22_X1 U16625 ( .A1(n14215), .A2(n15610), .B1(n15609), .B2(n15870), .ZN(
        P2_U3436) );
  NAND2_X1 U16626 ( .A1(n15615), .A2(n15793), .ZN(n15611) );
  OAI211_X1 U16627 ( .C1(n15613), .C2(n15797), .A(n15612), .B(n15611), .ZN(
        n15614) );
  AOI21_X1 U16628 ( .B1(n15615), .B2(n15632), .A(n15614), .ZN(n15617) );
  INV_X1 U16629 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U16630 ( .A1(n15839), .A2(n15617), .B1(n15616), .B2(n15970), .ZN(
        P3_U3462) );
  INV_X1 U16631 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U16632 ( .A1(n15980), .A2(n15618), .B1(n15617), .B2(n15978), .ZN(
        P3_U3399) );
  OAI21_X1 U16633 ( .B1(n15620), .B2(n15919), .A(n15619), .ZN(n15622) );
  AOI211_X1 U16634 ( .C1(n15777), .C2(n15623), .A(n15622), .B(n15621), .ZN(
        n15626) );
  AOI22_X1 U16635 ( .A1(n15717), .A2(n15626), .B1(n15624), .B2(n15924), .ZN(
        P1_U3531) );
  INV_X1 U16636 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U16637 ( .A1(n15719), .A2(n15626), .B1(n15625), .B2(n15926), .ZN(
        P1_U3468) );
  INV_X1 U16638 ( .A(n15630), .ZN(n15633) );
  AOI21_X1 U16639 ( .B1(n15737), .B2(n15628), .A(n15627), .ZN(n15629) );
  OAI21_X1 U16640 ( .B1(n15732), .B2(n15630), .A(n15629), .ZN(n15631) );
  AOI21_X1 U16641 ( .B1(n15633), .B2(n15632), .A(n15631), .ZN(n15634) );
  AOI22_X1 U16642 ( .A1(n15839), .A2(n15634), .B1(n10839), .B2(n15970), .ZN(
        P3_U3463) );
  INV_X1 U16643 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U16644 ( .A1(n15980), .A2(n15635), .B1(n15634), .B2(n15978), .ZN(
        P3_U3402) );
  OAI21_X1 U16645 ( .B1(n15637), .B2(n15753), .A(n15636), .ZN(n15638) );
  AOI21_X1 U16646 ( .B1(n15639), .B2(n15758), .A(n15638), .ZN(n15640) );
  AND2_X1 U16647 ( .A1(n15641), .A2(n15640), .ZN(n15644) );
  AOI22_X1 U16648 ( .A1(n15869), .A2(n15644), .B1(n15642), .B2(n15868), .ZN(
        P2_U3503) );
  INV_X1 U16649 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15643) );
  AOI22_X1 U16650 ( .A1(n14215), .A2(n15644), .B1(n15643), .B2(n15870), .ZN(
        P2_U3442) );
  INV_X1 U16651 ( .A(n15645), .ZN(n15649) );
  OAI21_X1 U16652 ( .B1(n15797), .B2(n15647), .A(n15646), .ZN(n15648) );
  AOI21_X1 U16653 ( .B1(n15649), .B2(n15802), .A(n15648), .ZN(n15650) );
  AOI22_X1 U16654 ( .A1(n15839), .A2(n15650), .B1(n10933), .B2(n15970), .ZN(
        P3_U3464) );
  INV_X1 U16655 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15651) );
  AOI22_X1 U16656 ( .A1(n15980), .A2(n15651), .B1(n15650), .B2(n15978), .ZN(
        P3_U3405) );
  INV_X1 U16657 ( .A(n11774), .ZN(n15653) );
  AOI21_X1 U16658 ( .B1(n15658), .B2(n15652), .A(n15653), .ZN(n15672) );
  INV_X1 U16659 ( .A(n15654), .ZN(n15655) );
  OAI211_X1 U16660 ( .C1(n15668), .C2(n15656), .A(n15655), .B(n15917), .ZN(
        n15670) );
  OAI21_X1 U16661 ( .B1(n15668), .B2(n15919), .A(n15670), .ZN(n15663) );
  XNOR2_X1 U16662 ( .A(n15657), .B(n15658), .ZN(n15659) );
  NOR2_X1 U16663 ( .A1(n15659), .A2(n15890), .ZN(n15661) );
  AOI211_X1 U16664 ( .C1(n15672), .C2(n15749), .A(n15661), .B(n15660), .ZN(
        n15675) );
  INV_X1 U16665 ( .A(n15675), .ZN(n15662) );
  AOI211_X1 U16666 ( .C1(n15777), .C2(n15672), .A(n15663), .B(n15662), .ZN(
        n15665) );
  AOI22_X1 U16667 ( .A1(n15717), .A2(n15665), .B1(n10514), .B2(n15924), .ZN(
        P1_U3533) );
  INV_X1 U16668 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U16669 ( .A1(n15719), .A2(n15665), .B1(n15664), .B2(n15926), .ZN(
        P1_U3474) );
  AOI22_X1 U16670 ( .A1(n15941), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15666), 
        .B2(n15930), .ZN(n15667) );
  OAI21_X1 U16671 ( .B1(n15723), .B2(n15668), .A(n15667), .ZN(n15669) );
  INV_X1 U16672 ( .A(n15669), .ZN(n15674) );
  INV_X1 U16673 ( .A(n15670), .ZN(n15671) );
  AOI22_X1 U16674 ( .A1(n15672), .A2(n15784), .B1(n15935), .B2(n15671), .ZN(
        n15673) );
  OAI211_X1 U16675 ( .C1(n15941), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        P1_U3288) );
  INV_X1 U16676 ( .A(n15676), .ZN(n15835) );
  AOI22_X1 U16677 ( .A1(n15677), .A2(n15839), .B1(n15835), .B2(n15683), .ZN(
        n15678) );
  OAI21_X1 U16678 ( .B1(n15839), .B2(n15679), .A(n15678), .ZN(P3_U3465) );
  AOI222_X1 U16679 ( .A1(n15685), .A2(n15684), .B1(n15683), .B2(n15682), .C1(
        n15681), .C2(n15680), .ZN(n15686) );
  OAI221_X1 U16680 ( .B1(n15690), .B2(n15689), .C1(n15688), .C2(n15687), .A(
        n15686), .ZN(P3_U3227) );
  OAI21_X1 U16681 ( .B1(n15692), .B2(n15919), .A(n15691), .ZN(n15694) );
  AOI211_X1 U16682 ( .C1(n15777), .C2(n15695), .A(n15694), .B(n15693), .ZN(
        n15696) );
  AOI22_X1 U16683 ( .A1(n15717), .A2(n15696), .B1(n10518), .B2(n15924), .ZN(
        P1_U3534) );
  AOI22_X1 U16684 ( .A1(n15719), .A2(n15696), .B1(n9016), .B2(n15926), .ZN(
        P1_U3477) );
  AOI21_X1 U16685 ( .B1(n15733), .B2(n15732), .A(n15697), .ZN(n15700) );
  INV_X1 U16686 ( .A(n15698), .ZN(n15699) );
  AOI211_X1 U16687 ( .C1(n15737), .C2(n15701), .A(n15700), .B(n15699), .ZN(
        n15703) );
  INV_X1 U16688 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15702) );
  AOI22_X1 U16689 ( .A1(n15839), .A2(n15703), .B1(n15702), .B2(n15970), .ZN(
        P3_U3466) );
  INV_X1 U16690 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15704) );
  AOI22_X1 U16691 ( .A1(n15980), .A2(n15704), .B1(n15703), .B2(n15978), .ZN(
        P3_U3411) );
  XNOR2_X1 U16692 ( .A(n15705), .B(n15710), .ZN(n15727) );
  INV_X1 U16693 ( .A(n15706), .ZN(n15708) );
  OAI211_X1 U16694 ( .C1(n15708), .C2(n15722), .A(n15917), .B(n15707), .ZN(
        n15725) );
  OAI21_X1 U16695 ( .B1(n15722), .B2(n15919), .A(n15725), .ZN(n15715) );
  XOR2_X1 U16696 ( .A(n15709), .B(n15710), .Z(n15712) );
  OAI21_X1 U16697 ( .B1(n15712), .B2(n15890), .A(n15711), .ZN(n15713) );
  AOI21_X1 U16698 ( .B1(n15727), .B2(n15749), .A(n15713), .ZN(n15730) );
  INV_X1 U16699 ( .A(n15730), .ZN(n15714) );
  AOI211_X1 U16700 ( .C1(n15777), .C2(n15727), .A(n15715), .B(n15714), .ZN(
        n15718) );
  AOI22_X1 U16701 ( .A1(n15717), .A2(n15718), .B1(n15716), .B2(n15924), .ZN(
        P1_U3535) );
  AOI22_X1 U16702 ( .A1(n15719), .A2(n15718), .B1(n9038), .B2(n15926), .ZN(
        P1_U3480) );
  AOI22_X1 U16703 ( .A1(n15941), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n15720), 
        .B2(n15930), .ZN(n15721) );
  OAI21_X1 U16704 ( .B1(n15723), .B2(n15722), .A(n15721), .ZN(n15724) );
  INV_X1 U16705 ( .A(n15724), .ZN(n15729) );
  INV_X1 U16706 ( .A(n15725), .ZN(n15726) );
  AOI22_X1 U16707 ( .A1(n15727), .A2(n15784), .B1(n15935), .B2(n15726), .ZN(
        n15728) );
  OAI211_X1 U16708 ( .C1(n15941), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        P1_U3286) );
  AOI21_X1 U16709 ( .B1(n15733), .B2(n15732), .A(n15731), .ZN(n15735) );
  AOI211_X1 U16710 ( .C1(n15737), .C2(n15736), .A(n15735), .B(n15734), .ZN(
        n15739) );
  AOI22_X1 U16711 ( .A1(n15839), .A2(n15739), .B1(n15738), .B2(n15970), .ZN(
        P3_U3467) );
  INV_X1 U16712 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15740) );
  AOI22_X1 U16713 ( .A1(n15980), .A2(n15740), .B1(n15739), .B2(n15978), .ZN(
        P3_U3414) );
  AOI21_X1 U16714 ( .B1(n15742), .B2(n15887), .A(n15741), .ZN(n15743) );
  OAI21_X1 U16715 ( .B1(n15745), .B2(n15744), .A(n15743), .ZN(n15746) );
  AOI211_X1 U16716 ( .C1(n15749), .C2(n15748), .A(n15747), .B(n15746), .ZN(
        n15750) );
  AOI22_X1 U16717 ( .A1(n15717), .A2(n15750), .B1(n10542), .B2(n15924), .ZN(
        P1_U3536) );
  AOI22_X1 U16718 ( .A1(n15719), .A2(n15750), .B1(n9053), .B2(n15926), .ZN(
        P1_U3483) );
  INV_X1 U16719 ( .A(n15751), .ZN(n15757) );
  OAI21_X1 U16720 ( .B1(n15754), .B2(n15753), .A(n15752), .ZN(n15756) );
  AOI211_X1 U16721 ( .C1(n15758), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15761) );
  AOI22_X1 U16722 ( .A1(n15869), .A2(n15761), .B1(n15759), .B2(n15868), .ZN(
        P2_U3507) );
  INV_X1 U16723 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U16724 ( .A1(n14215), .A2(n15761), .B1(n15760), .B2(n15870), .ZN(
        P2_U3454) );
  AOI21_X1 U16725 ( .B1(n15768), .B2(n15763), .A(n15762), .ZN(n15772) );
  INV_X1 U16726 ( .A(n15772), .ZN(n15785) );
  INV_X1 U16727 ( .A(n15764), .ZN(n15765) );
  OAI211_X1 U16728 ( .C1(n15767), .C2(n15766), .A(n15765), .B(n15917), .ZN(
        n15782) );
  OAI21_X1 U16729 ( .B1(n15767), .B2(n15919), .A(n15782), .ZN(n15776) );
  XOR2_X1 U16730 ( .A(n15769), .B(n15768), .Z(n15774) );
  OAI21_X1 U16731 ( .B1(n15772), .B2(n15771), .A(n15770), .ZN(n15773) );
  AOI21_X1 U16732 ( .B1(n15774), .B2(n15914), .A(n15773), .ZN(n15788) );
  INV_X1 U16733 ( .A(n15788), .ZN(n15775) );
  AOI211_X1 U16734 ( .C1(n15777), .C2(n15785), .A(n15776), .B(n15775), .ZN(
        n15779) );
  AOI22_X1 U16735 ( .A1(n15717), .A2(n15779), .B1(n10546), .B2(n15924), .ZN(
        P1_U3537) );
  INV_X1 U16736 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U16737 ( .A1(n15719), .A2(n15779), .B1(n15778), .B2(n15926), .ZN(
        P1_U3486) );
  AOI222_X1 U16738 ( .A1(n15781), .A2(n15931), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n15941), .C1(n15930), .C2(n15780), .ZN(n15787) );
  INV_X1 U16739 ( .A(n15782), .ZN(n15783) );
  AOI22_X1 U16740 ( .A1(n15785), .A2(n15784), .B1(n15935), .B2(n15783), .ZN(
        n15786) );
  OAI211_X1 U16741 ( .C1(n15941), .C2(n15788), .A(n15787), .B(n15786), .ZN(
        P1_U3284) );
  NOR2_X1 U16742 ( .A1(n15789), .A2(n15797), .ZN(n15791) );
  AOI211_X1 U16743 ( .C1(n15793), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15795) );
  AOI22_X1 U16744 ( .A1(n15839), .A2(n15795), .B1(n15794), .B2(n15970), .ZN(
        P3_U3469) );
  INV_X1 U16745 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15796) );
  AOI22_X1 U16746 ( .A1(n15980), .A2(n15796), .B1(n15795), .B2(n15978), .ZN(
        P3_U3420) );
  NOR2_X1 U16747 ( .A1(n15798), .A2(n15797), .ZN(n15800) );
  AOI211_X1 U16748 ( .C1(n15802), .C2(n15801), .A(n15800), .B(n15799), .ZN(
        n15804) );
  INV_X1 U16749 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15803) );
  AOI22_X1 U16750 ( .A1(n15839), .A2(n15804), .B1(n15803), .B2(n15970), .ZN(
        P3_U3470) );
  INV_X1 U16751 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15805) );
  AOI22_X1 U16752 ( .A1(n15980), .A2(n15805), .B1(n15804), .B2(n15978), .ZN(
        P3_U3423) );
  NOR3_X1 U16753 ( .A1(n15807), .A2(n15806), .A3(n15851), .ZN(n15811) );
  NOR2_X1 U16754 ( .A1(n7560), .A2(n15919), .ZN(n15809) );
  NOR4_X1 U16755 ( .A1(n15811), .A2(n15810), .A3(n15809), .A4(n15808), .ZN(
        n15813) );
  AOI22_X1 U16756 ( .A1(n15717), .A2(n15813), .B1(n10549), .B2(n15924), .ZN(
        P1_U3539) );
  INV_X1 U16757 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U16758 ( .A1(n15719), .A2(n15813), .B1(n15812), .B2(n15926), .ZN(
        P1_U3492) );
  NAND2_X1 U16759 ( .A1(n15815), .A2(n15814), .ZN(n15820) );
  AOI22_X1 U16760 ( .A1(n15818), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n15817), 
        .B2(n15816), .ZN(n15819) );
  OAI211_X1 U16761 ( .C1(n15822), .C2(n15821), .A(n15820), .B(n15819), .ZN(
        n15823) );
  AOI21_X1 U16762 ( .B1(n15825), .B2(n15824), .A(n15823), .ZN(n15826) );
  OAI21_X1 U16763 ( .B1(n13980), .B2(n15827), .A(n15826), .ZN(P2_U3254) );
  OAI21_X1 U16764 ( .B1(n15829), .B2(n15919), .A(n15828), .ZN(n15830) );
  AOI211_X1 U16765 ( .C1(n15832), .C2(n15923), .A(n15831), .B(n15830), .ZN(
        n15833) );
  AOI22_X1 U16766 ( .A1(n15717), .A2(n15833), .B1(n10541), .B2(n15924), .ZN(
        P1_U3540) );
  AOI22_X1 U16767 ( .A1(n15719), .A2(n15833), .B1(n9122), .B2(n15926), .ZN(
        P1_U3495) );
  INV_X1 U16768 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15838) );
  AOI22_X1 U16769 ( .A1(n15836), .A2(n15839), .B1(n15835), .B2(n15834), .ZN(
        n15837) );
  OAI21_X1 U16770 ( .B1(n15839), .B2(n15838), .A(n15837), .ZN(P3_U3472) );
  NOR2_X1 U16771 ( .A1(n15840), .A2(n15890), .ZN(n15845) );
  OAI211_X1 U16772 ( .C1(n15843), .C2(n15919), .A(n15842), .B(n15841), .ZN(
        n15844) );
  AOI211_X1 U16773 ( .C1(n15846), .C2(n15923), .A(n15845), .B(n15844), .ZN(
        n15847) );
  AOI22_X1 U16774 ( .A1(n15717), .A2(n15847), .B1(n10727), .B2(n15924), .ZN(
        P1_U3541) );
  AOI22_X1 U16775 ( .A1(n15719), .A2(n15847), .B1(n9137), .B2(n15926), .ZN(
        P1_U3498) );
  OAI211_X1 U16776 ( .C1(n15850), .C2(n15919), .A(n15849), .B(n15848), .ZN(
        n15855) );
  NOR3_X1 U16777 ( .A1(n15853), .A2(n15852), .A3(n15851), .ZN(n15854) );
  AOI211_X1 U16778 ( .C1(n15856), .C2(n15914), .A(n15855), .B(n15854), .ZN(
        n15858) );
  INV_X1 U16779 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15857) );
  AOI22_X1 U16780 ( .A1(n15717), .A2(n15858), .B1(n15857), .B2(n15924), .ZN(
        P1_U3542) );
  AOI22_X1 U16781 ( .A1(n15719), .A2(n15858), .B1(n9161), .B2(n15926), .ZN(
        P1_U3501) );
  NAND2_X1 U16782 ( .A1(n15860), .A2(n15859), .ZN(n15866) );
  NAND2_X1 U16783 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  AND2_X1 U16784 ( .A1(n15864), .A2(n15863), .ZN(n15865) );
  AOI22_X1 U16785 ( .A1(n15869), .A2(n15872), .B1(n11383), .B2(n15868), .ZN(
        P2_U3513) );
  INV_X1 U16786 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U16787 ( .A1(n14215), .A2(n15872), .B1(n15871), .B2(n15870), .ZN(
        P2_U3472) );
  INV_X1 U16788 ( .A(n15873), .ZN(n15881) );
  NOR3_X1 U16789 ( .A1(n15875), .A2(n15874), .A3(n15890), .ZN(n15880) );
  OAI211_X1 U16790 ( .C1(n15878), .C2(n15919), .A(n15877), .B(n15876), .ZN(
        n15879) );
  AOI211_X1 U16791 ( .C1(n15881), .C2(n15923), .A(n15880), .B(n15879), .ZN(
        n15884) );
  AOI22_X1 U16792 ( .A1(n15717), .A2(n15884), .B1(n15882), .B2(n15924), .ZN(
        P1_U3543) );
  INV_X1 U16793 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U16794 ( .A1(n15719), .A2(n15884), .B1(n15883), .B2(n15926), .ZN(
        P1_U3504) );
  AOI211_X1 U16795 ( .C1(n15888), .C2(n15887), .A(n15886), .B(n15885), .ZN(
        n15889) );
  OAI21_X1 U16796 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(n15892) );
  AOI21_X1 U16797 ( .B1(n15893), .B2(n15923), .A(n15892), .ZN(n15896) );
  AOI22_X1 U16798 ( .A1(n15717), .A2(n15896), .B1(n15894), .B2(n15924), .ZN(
        P1_U3544) );
  INV_X1 U16799 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15895) );
  AOI22_X1 U16800 ( .A1(n15719), .A2(n15896), .B1(n15895), .B2(n15926), .ZN(
        P1_U3507) );
  NAND2_X1 U16801 ( .A1(n15898), .A2(n15897), .ZN(n15900) );
  XOR2_X1 U16802 ( .A(n15900), .B(n15899), .Z(n15905) );
  OAI22_X1 U16803 ( .A1(n15904), .A2(n15903), .B1(n15902), .B2(n15901), .ZN(
        n15913) );
  AOI222_X1 U16804 ( .A1(n15965), .A2(n15932), .B1(n15963), .B2(n15905), .C1(
        n15913), .C2(n15960), .ZN(n15907) );
  OAI211_X1 U16805 ( .C1(n15969), .C2(n15908), .A(n15907), .B(n15906), .ZN(
        P1_U3228) );
  AOI21_X1 U16806 ( .B1(n15911), .B2(n15910), .A(n15909), .ZN(n15937) );
  XNOR2_X1 U16807 ( .A(n15912), .B(n15911), .ZN(n15915) );
  AOI21_X1 U16808 ( .B1(n15915), .B2(n15914), .A(n15913), .ZN(n15940) );
  INV_X1 U16809 ( .A(n15940), .ZN(n15922) );
  OAI211_X1 U16810 ( .C1(n15920), .C2(n15918), .A(n15917), .B(n15916), .ZN(
        n15933) );
  OAI21_X1 U16811 ( .B1(n15920), .B2(n15919), .A(n15933), .ZN(n15921) );
  AOI211_X1 U16812 ( .C1(n15937), .C2(n15923), .A(n15922), .B(n15921), .ZN(
        n15928) );
  AOI22_X1 U16813 ( .A1(n15717), .A2(n15928), .B1(n15925), .B2(n15924), .ZN(
        P1_U3545) );
  INV_X1 U16814 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15927) );
  AOI22_X1 U16815 ( .A1(n15719), .A2(n15928), .B1(n15927), .B2(n15926), .ZN(
        P1_U3510) );
  AOI222_X1 U16816 ( .A1(n15932), .A2(n15931), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n15941), .C1(n15930), .C2(n15929), .ZN(n15939) );
  INV_X1 U16817 ( .A(n15933), .ZN(n15934) );
  AOI22_X1 U16818 ( .A1(n15937), .A2(n15936), .B1(n15935), .B2(n15934), .ZN(
        n15938) );
  OAI211_X1 U16819 ( .C1(n15941), .C2(n15940), .A(n15939), .B(n15938), .ZN(
        P1_U3276) );
  OAI22_X1 U16820 ( .A1(n15945), .A2(n15944), .B1(n15943), .B2(n15942), .ZN(
        n15952) );
  XOR2_X1 U16821 ( .A(n15947), .B(n15948), .Z(n15950) );
  NOR2_X1 U16822 ( .A1(n15950), .A2(n15949), .ZN(n15951) );
  AOI211_X1 U16823 ( .C1(n15953), .C2(n15965), .A(n15952), .B(n15951), .ZN(
        n15955) );
  OAI211_X1 U16824 ( .C1(n15969), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P1_U3238) );
  XNOR2_X1 U16825 ( .A(n15957), .B(n15958), .ZN(n15962) );
  INV_X1 U16826 ( .A(n15959), .ZN(n15961) );
  AOI222_X1 U16827 ( .A1(n15965), .A2(n15964), .B1(n15963), .B2(n15962), .C1(
        n15961), .C2(n15960), .ZN(n15967) );
  OAI211_X1 U16828 ( .C1(n15969), .C2(n15968), .A(n15967), .B(n15966), .ZN(
        P1_U3219) );
  AOI22_X1 U16829 ( .A1(n15975), .A2(n15971), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15970), .ZN(n15973) );
  NAND2_X1 U16830 ( .A1(n15973), .A2(n15972), .ZN(P3_U3489) );
  INV_X1 U16831 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U16832 ( .A1(n15975), .A2(n15974), .ZN(n15976) );
  OAI221_X1 U16833 ( .B1(n15980), .B2(n15979), .C1(n15978), .C2(n15977), .A(
        n15976), .ZN(P3_U3457) );
  AOI21_X1 U16834 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15981) );
  OAI21_X1 U16835 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n15981), 
        .ZN(U28) );
  AOI21_X1 U7546 ( .B1(n7761), .B2(n7251), .A(n7757), .ZN(n12883) );
  CLKBUF_X1 U7332 ( .A(n8919), .Z(n9370) );
  OAI21_X1 U7357 ( .B1(n12765), .B2(n7763), .A(n7754), .ZN(n7761) );
  CLKBUF_X1 U7542 ( .A(n8901), .Z(n8906) );
  OR2_X1 U7560 ( .A1(n9981), .A2(n9997), .ZN(n13085) );
  CLKBUF_X1 U7681 ( .A(n13025), .Z(n7209) );
  CLKBUF_X1 U7929 ( .A(n10708), .Z(n13976) );
endmodule

