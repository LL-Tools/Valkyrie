

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312;

  CLKBUF_X2 U2551 ( .A(n2941), .Z(n4375) );
  INV_X2 U2552 ( .A(IR_REG_31__SCAN_IN), .ZN(n4908) );
  INV_X2 U2553 ( .A(n3843), .ZN(n3824) );
  NAND2_X1 U2554 ( .A1(n3191), .A2(n3094), .ZN(n3190) );
  NAND2_X1 U2555 ( .A1(n4774), .A2(n2535), .ZN(n4754) );
  INV_X1 U2556 ( .A(n3446), .ZN(n3310) );
  NAND2_X2 U2557 ( .A1(n3807), .A2(n2599), .ZN(n4708) );
  AOI22_X2 U2558 ( .A1(n4699), .A2(n3659), .B1(n4684), .B2(n4711), .ZN(n4689)
         );
  BUF_X2 U2560 ( .A(n2792), .Z(n2517) );
  XNOR2_X1 U2561 ( .A(n2747), .B(n2746), .ZN(n2792) );
  NAND2_X2 U2562 ( .A1(n2782), .A2(IR_REG_31__SCAN_IN), .ZN(n2781) );
  NOR2_X1 U2563 ( .A1(n2525), .A2(n4852), .ZN(n2560) );
  NAND2_X1 U2564 ( .A1(n4482), .A2(n4369), .ZN(n3491) );
  INV_X1 U2565 ( .A(n3505), .ZN(n3504) );
  OR2_X1 U2566 ( .A1(n3394), .A2(n3393), .ZN(n3471) );
  NAND2_X1 U2567 ( .A1(n3246), .A2(n4371), .ZN(n3259) );
  NAND2_X1 U2568 ( .A1(n3182), .A2(n4387), .ZN(n3241) );
  NAND2_X1 U2569 ( .A1(n3173), .A2(n4439), .ZN(n3245) );
  OR2_X1 U2570 ( .A1(n3172), .A2(n3171), .ZN(n3173) );
  NAND2_X1 U2571 ( .A1(n4979), .A2(n2917), .ZN(n4990) );
  XNOR2_X1 U2572 ( .A(n2843), .B(n3843), .ZN(n2654) );
  AOI21_X1 U2573 ( .B1(n3023), .B2(n3828), .A(n2844), .ZN(n2925) );
  AOI21_X1 U2574 ( .B1(n3114), .B2(n3029), .A(n3028), .ZN(n3031) );
  NAND2_X1 U2575 ( .A1(n3042), .A2(n4388), .ZN(n3105) );
  XNOR2_X1 U2576 ( .A(n2842), .B(n4915), .ZN(n2841) );
  INV_X1 U2577 ( .A(n4540), .ZN(n3159) );
  NAND2_X1 U2578 ( .A1(n2812), .A2(IR_REG_31__SCAN_IN), .ZN(n2747) );
  INV_X2 U2579 ( .A(n2966), .ZN(n3130) );
  BUF_X2 U2580 ( .A(n2937), .Z(n3612) );
  CLKBUF_X3 U2581 ( .A(n2955), .Z(n4404) );
  NAND2_X1 U2582 ( .A1(n2763), .A2(n2772), .ZN(n2955) );
  AND2_X1 U2583 ( .A1(n4561), .A2(n2628), .ZN(n2908) );
  NAND2_X1 U2584 ( .A1(n2651), .A2(n2836), .ZN(n2906) );
  INV_X1 U2585 ( .A(IR_REG_14__SCAN_IN), .ZN(n3959) );
  INV_X1 U2586 ( .A(IR_REG_10__SCAN_IN), .ZN(n3949) );
  INV_X1 U2587 ( .A(IR_REG_4__SCAN_IN), .ZN(n3944) );
  NOR2_X1 U2588 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2718)
         );
  NOR2_X1 U2589 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2717)
         );
  NOR2_X2 U2590 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2880)
         );
  INV_X1 U2591 ( .A(IR_REG_20__SCAN_IN), .ZN(n2746) );
  INV_X1 U2592 ( .A(IR_REG_18__SCAN_IN), .ZN(n4160) );
  INV_X1 U2593 ( .A(IR_REG_13__SCAN_IN), .ZN(n4156) );
  INV_X1 U2594 ( .A(IR_REG_2__SCAN_IN), .ZN(n4132) );
  INV_X1 U2595 ( .A(IR_REG_16__SCAN_IN), .ZN(n2742) );
  OAI21_X2 U2596 ( .B1(n4286), .B2(n4342), .A(n4341), .ZN(n4340) );
  AOI21_X2 U2597 ( .B1(n3730), .B2(n4288), .A(n4287), .ZN(n4286) );
  OAI22_X2 U2598 ( .A1(n3784), .A2(n3763), .B1(n3762), .B2(n3761), .ZN(n4322)
         );
  NAND2_X2 U2599 ( .A1(n2678), .A2(n2676), .ZN(n3784) );
  OR2_X2 U2600 ( .A1(n4322), .A2(n4323), .ZN(n3775) );
  OAI21_X2 U2601 ( .B1(n3326), .B2(n3325), .A(n3791), .ZN(n3352) );
  NAND2_X2 U2602 ( .A1(n3789), .A2(n3324), .ZN(n3791) );
  NAND2_X1 U2603 ( .A1(n2624), .A2(n4170), .ZN(n2623) );
  INV_X1 U2604 ( .A(n2625), .ZN(n2624) );
  NAND2_X1 U2605 ( .A1(n3442), .A2(n3443), .ZN(n2696) );
  NOR2_X2 U2606 ( .A1(n3456), .A2(n2793), .ZN(n3828) );
  INV_X1 U2607 ( .A(n5229), .ZN(n2793) );
  AND2_X1 U2608 ( .A1(n3243), .A2(n3240), .ZN(n2615) );
  AND2_X1 U2609 ( .A1(n4915), .A2(n4916), .ZN(n2853) );
  INV_X1 U2610 ( .A(n3612), .ZN(n3680) );
  NAND2_X1 U2611 ( .A1(n4990), .A2(n4989), .ZN(n4988) );
  OR2_X1 U2612 ( .A1(n4622), .A2(n2555), .ZN(n2554) );
  NOR2_X1 U2613 ( .A1(n2523), .A2(n4675), .ZN(n5297) );
  AOI21_X1 U2614 ( .B1(n4689), .B2(n3671), .A(n3670), .ZN(n4663) );
  NAND2_X1 U2615 ( .A1(n3636), .A2(REG3_REG_24__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U2616 ( .A1(n2590), .A2(n2593), .ZN(n4789) );
  INV_X1 U2617 ( .A(n2594), .ZN(n2593) );
  OAI21_X1 U2618 ( .B1(n4817), .B2(n2595), .A(n4793), .ZN(n2594) );
  NAND2_X1 U2619 ( .A1(n4818), .A2(n4817), .ZN(n4816) );
  AND2_X1 U2620 ( .A1(n3388), .A2(n3387), .ZN(n3390) );
  OR2_X1 U2621 ( .A1(n5229), .A2(n4848), .ZN(n4856) );
  NAND2_X1 U2622 ( .A1(n2723), .A2(n2565), .ZN(n2783) );
  NOR2_X1 U2623 ( .A1(n2707), .A2(IR_REG_25__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U2624 ( .A1(n2530), .A2(n2708), .ZN(n2707) );
  INV_X1 U2625 ( .A(IR_REG_28__SCAN_IN), .ZN(n3983) );
  NAND3_X1 U2626 ( .A1(n2697), .A2(n2616), .A3(n2622), .ZN(n2761) );
  AND2_X1 U2627 ( .A1(n2640), .A2(n2722), .ZN(n2616) );
  AND2_X1 U2628 ( .A1(n4174), .A2(n2708), .ZN(n2640) );
  AND2_X1 U2629 ( .A1(n2721), .A2(n2698), .ZN(n2697) );
  NOR2_X1 U2630 ( .A1(n2700), .A2(IR_REG_21__SCAN_IN), .ZN(n2698) );
  NAND3_X1 U2631 ( .A1(n4913), .A2(n4912), .A3(n4914), .ZN(n2821) );
  AOI21_X1 U2632 ( .B1(n2664), .B2(n2667), .A(n2536), .ZN(n2663) );
  INV_X1 U2633 ( .A(n3838), .ZN(n2666) );
  INV_X1 U2634 ( .A(n3520), .ZN(n2684) );
  INV_X1 U2635 ( .A(n2689), .ZN(n2685) );
  INV_X1 U2636 ( .A(n2938), .ZN(n2966) );
  NAND2_X1 U2637 ( .A1(n4624), .A2(n4625), .ZN(n4639) );
  NOR2_X1 U2638 ( .A1(n2606), .A2(n3644), .ZN(n2604) );
  OR2_X1 U2639 ( .A1(n4763), .A2(n3635), .ZN(n4395) );
  NAND2_X1 U2640 ( .A1(n3479), .A2(n5199), .ZN(n2632) );
  OAI21_X1 U2641 ( .B1(n3245), .B2(n3244), .A(n4438), .ZN(n3246) );
  NAND2_X1 U2642 ( .A1(n4778), .A2(n4493), .ZN(n3703) );
  INV_X1 U2643 ( .A(n5182), .ZN(n5199) );
  NOR2_X1 U2644 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2722)
         );
  INV_X1 U2645 ( .A(n2728), .ZN(n2725) );
  INV_X1 U2646 ( .A(IR_REG_24__SCAN_IN), .ZN(n3975) );
  OR2_X1 U2647 ( .A1(n2730), .A2(n4908), .ZN(n2733) );
  INV_X1 U2648 ( .A(IR_REG_23__SCAN_IN), .ZN(n3974) );
  NOR2_X1 U2649 ( .A1(n2588), .A2(n2587), .ZN(n2721) );
  NOR2_X1 U2650 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2589)
         );
  NAND2_X1 U2651 ( .A1(n3949), .A2(n2626), .ZN(n2625) );
  INV_X1 U2652 ( .A(IR_REG_9__SCAN_IN), .ZN(n2626) );
  NOR2_X1 U2653 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2720)
         );
  INV_X1 U2654 ( .A(IR_REG_5__SCAN_IN), .ZN(n4140) );
  NAND2_X1 U2655 ( .A1(n2691), .A2(n2690), .ZN(n2689) );
  INV_X1 U2656 ( .A(n5183), .ZN(n2690) );
  AOI21_X1 U2657 ( .B1(n2691), .B2(n2688), .A(n2529), .ZN(n2687) );
  NOR2_X1 U2658 ( .A1(n5183), .A2(n2693), .ZN(n2688) );
  NOR2_X1 U2659 ( .A1(n2657), .A2(n2716), .ZN(n2656) );
  INV_X1 U2660 ( .A(n2663), .ZN(n2657) );
  NAND2_X1 U2661 ( .A1(n2663), .A2(n2660), .ZN(n2659) );
  NAND2_X1 U2662 ( .A1(n2665), .A2(n2661), .ZN(n2660) );
  INV_X1 U2663 ( .A(n2716), .ZN(n2661) );
  NAND2_X1 U2664 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  INV_X1 U2665 ( .A(n3039), .ZN(n2854) );
  AOI21_X1 U2666 ( .B1(n2704), .B2(n2703), .A(n3819), .ZN(n2702) );
  INV_X1 U2667 ( .A(n3774), .ZN(n2703) );
  OAI22_X1 U2668 ( .A1(n3030), .A2(n3446), .B1(n3037), .B2(n3719), .ZN(n2956)
         );
  XNOR2_X1 U2669 ( .A(n2948), .B(n3843), .ZN(n2959) );
  NAND2_X1 U2670 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  NOR2_X1 U2671 ( .A1(n3228), .A2(n4313), .ZN(n3261) );
  AOI21_X1 U2672 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2795), .A(n2845), .ZN(n2847)
         );
  OR2_X1 U2673 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  AND2_X1 U2674 ( .A1(n2696), .A2(n3350), .ZN(n2693) );
  OR2_X1 U2675 ( .A1(n2694), .A2(n2692), .ZN(n2691) );
  INV_X1 U2676 ( .A(n2696), .ZN(n2692) );
  AND2_X1 U2677 ( .A1(n3444), .A2(n2695), .ZN(n2694) );
  NAND2_X1 U2678 ( .A1(n3351), .A2(n3350), .ZN(n2695) );
  NAND2_X1 U2679 ( .A1(n4925), .A2(REG2_REG_2__SCAN_IN), .ZN(n2628) );
  XNOR2_X1 U2680 ( .A(n2909), .B(n2888), .ZN(n5044) );
  NAND2_X1 U2681 ( .A1(n5044), .A2(REG2_REG_4__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U2682 ( .A1(n4583), .A2(n2896), .ZN(n2897) );
  NAND2_X1 U2683 ( .A1(n4588), .A2(n2915), .ZN(n2916) );
  NAND2_X1 U2684 ( .A1(n4985), .A2(n2899), .ZN(n2548) );
  NAND2_X1 U2685 ( .A1(n3212), .A2(n3213), .ZN(n4606) );
  NAND2_X1 U2686 ( .A1(n4998), .A2(REG2_REG_13__SCAN_IN), .ZN(n2621) );
  XNOR2_X1 U2687 ( .A(n4639), .B(n4919), .ZN(n4626) );
  NOR2_X1 U2688 ( .A1(n4626), .A2(REG2_REG_16__SCAN_IN), .ZN(n4640) );
  OR2_X1 U2689 ( .A1(n5036), .A2(n4636), .ZN(n2650) );
  INV_X1 U2690 ( .A(IR_REG_19__SCAN_IN), .ZN(n4161) );
  NAND2_X1 U2691 ( .A1(n2745), .A2(IR_REG_31__SCAN_IN), .ZN(n2813) );
  INV_X1 U2692 ( .A(n5035), .ZN(n2649) );
  AOI21_X1 U2693 ( .B1(n2647), .B2(n4636), .A(n2543), .ZN(n2646) );
  AND2_X1 U2694 ( .A1(n4475), .A2(n4463), .ZN(n4664) );
  NAND2_X1 U2695 ( .A1(n2637), .A2(n2522), .ZN(n2636) );
  OR3_X1 U2696 ( .A1(n3652), .A2(n3651), .A3(n3650), .ZN(n3662) );
  AOI21_X1 U2697 ( .B1(n4708), .B2(n3705), .A(n4465), .ZN(n4682) );
  INV_X1 U2698 ( .A(n4521), .ZN(n4683) );
  AOI21_X1 U2699 ( .B1(n2600), .B2(n2598), .A(n2597), .ZN(n4699) );
  NOR2_X1 U2700 ( .A1(n2602), .A2(n2599), .ZN(n2598) );
  OAI21_X1 U2701 ( .B1(n2601), .B2(n2599), .A(n2539), .ZN(n2597) );
  INV_X1 U2702 ( .A(n4754), .ZN(n2600) );
  OAI21_X1 U2703 ( .B1(n2609), .B2(n2607), .A(n4395), .ZN(n2606) );
  OR2_X1 U2704 ( .A1(n4810), .A2(n5262), .ZN(n3609) );
  NAND2_X1 U2705 ( .A1(n4834), .A2(n3592), .ZN(n4818) );
  AND2_X1 U2706 ( .A1(n3601), .A2(n3600), .ZN(n4817) );
  NAND2_X1 U2707 ( .A1(n2542), .A2(n2519), .ZN(n2596) );
  AND2_X1 U2708 ( .A1(n4422), .A2(n4449), .ZN(n4369) );
  OR2_X1 U2709 ( .A1(n3385), .A2(n3384), .ZN(n5191) );
  OAI21_X1 U2710 ( .B1(n3241), .B2(n2612), .A(n2610), .ZN(n3301) );
  INV_X1 U2711 ( .A(n2611), .ZN(n2610) );
  NAND2_X1 U2712 ( .A1(n3241), .A2(n2615), .ZN(n3273) );
  AND4_X1 U2713 ( .A1(n2972), .A2(n2971), .A3(n2970), .A4(n2969), .ZN(n3095)
         );
  AND2_X1 U2714 ( .A1(n3092), .A2(n3091), .ZN(n3191) );
  INV_X1 U2715 ( .A(n4368), .ZN(n3094) );
  AND4_X1 U2716 ( .A1(n2852), .A2(n2851), .A3(n2850), .A4(n2849), .ZN(n3102)
         );
  NAND2_X1 U2717 ( .A1(n4385), .A2(n3065), .ZN(n3064) );
  INV_X1 U2718 ( .A(n5283), .ZN(n5293) );
  NAND2_X1 U2719 ( .A1(n3036), .A2(n5230), .ZN(n5257) );
  NAND2_X1 U2720 ( .A1(n2782), .A2(n2785), .ZN(n2787) );
  MUX2_X1 U2721 ( .A(IR_REG_31__SCAN_IN), .B(n2784), .S(IR_REG_29__SCAN_IN), 
        .Z(n2785) );
  NAND2_X1 U2722 ( .A1(n2761), .A2(IR_REG_31__SCAN_IN), .ZN(n2762) );
  INV_X1 U2723 ( .A(n2720), .ZN(n2700) );
  INV_X1 U2724 ( .A(n2721), .ZN(n2701) );
  INV_X1 U2725 ( .A(IR_REG_15__SCAN_IN), .ZN(n3421) );
  INV_X1 U2726 ( .A(IR_REG_11__SCAN_IN), .ZN(n4151) );
  AND2_X1 U2727 ( .A1(n2879), .A2(n2865), .ZN(n2874) );
  AOI22_X1 U2728 ( .A1(IR_REG_0__SCAN_IN), .A2(n2653), .B1(n2652), .B2(n4908), 
        .ZN(n2651) );
  INV_X1 U2729 ( .A(IR_REG_1__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U2730 ( .A1(n3775), .A2(n3774), .ZN(n3820) );
  AND2_X1 U2731 ( .A1(n3637), .A2(n3628), .ZN(n4749) );
  AND2_X1 U2732 ( .A1(n3790), .A2(n3792), .ZN(n3324) );
  NAND2_X1 U2733 ( .A1(n4267), .A2(n4268), .ZN(n4266) );
  AOI21_X1 U2734 ( .B1(n2679), .B2(n2681), .A(n2677), .ZN(n2676) );
  NAND2_X1 U2735 ( .A1(n4267), .A2(n2679), .ZN(n2678) );
  INV_X1 U2736 ( .A(n5266), .ZN(n2677) );
  AND2_X1 U2737 ( .A1(n3643), .A2(n3642), .ZN(n4407) );
  OR2_X1 U2738 ( .A1(n2830), .A2(n2817), .ZN(n4363) );
  INV_X1 U2739 ( .A(n3174), .ZN(n4536) );
  NAND2_X1 U2740 ( .A1(n4957), .A2(REG2_REG_3__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U2741 ( .A1(n4585), .A2(n2552), .ZN(n4583) );
  INV_X1 U2742 ( .A(n2553), .ZN(n2552) );
  OAI21_X1 U2743 ( .B1(n4923), .B2(REG1_REG_7__SCAN_IN), .A(n2896), .ZN(n2553)
         );
  XNOR2_X1 U2744 ( .A(n2897), .B(n2617), .ZN(n4977) );
  XNOR2_X1 U2745 ( .A(n4606), .B(n4596), .ZN(n3214) );
  NAND2_X1 U2746 ( .A1(n3214), .A2(REG2_REG_12__SCAN_IN), .ZN(n4608) );
  AOI211_X1 U2747 ( .C1(REG1_REG_15__SCAN_IN), .C2(n4920), .A(n4602), .B(n4604), .ZN(n4622) );
  NOR2_X1 U2748 ( .A1(n4623), .A2(REG1_REG_16__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U2749 ( .A1(n2650), .A2(n5035), .ZN(n5034) );
  NAND2_X1 U2750 ( .A1(n5034), .A2(n4638), .ZN(n2550) );
  AOI21_X1 U2751 ( .B1(n2650), .B2(n2647), .A(n5049), .ZN(n2551) );
  NAND2_X1 U2752 ( .A1(n2564), .A2(n2562), .ZN(n4851) );
  INV_X1 U2753 ( .A(n2563), .ZN(n2562) );
  NAND2_X1 U2754 ( .A1(n4673), .A2(n5151), .ZN(n2564) );
  OAI21_X1 U2755 ( .B1(n4683), .B2(n5154), .A(n4677), .ZN(n2563) );
  NAND2_X1 U2756 ( .A1(n2832), .A2(n2831), .ZN(n5216) );
  OR2_X1 U2757 ( .A1(n2778), .A2(n4908), .ZN(n2586) );
  AND2_X1 U2758 ( .A1(n2758), .A2(n2757), .ZN(n2778) );
  INV_X1 U2759 ( .A(n2761), .ZN(n2758) );
  INV_X1 U2760 ( .A(n4589), .ZN(n2570) );
  INV_X1 U2761 ( .A(n2915), .ZN(n2574) );
  INV_X1 U2762 ( .A(IR_REG_22__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U2763 ( .A1(n3774), .A2(n4323), .ZN(n2706) );
  NAND2_X1 U2764 ( .A1(n3221), .A2(n2668), .ZN(n2673) );
  INV_X1 U2765 ( .A(n3145), .ZN(n2668) );
  OAI22_X1 U2766 ( .A1(n3102), .A2(n3446), .B1(n3165), .B2(n3456), .ZN(n2930)
         );
  OAI21_X1 U2767 ( .B1(n3842), .B2(n3102), .A(n2931), .ZN(n2933) );
  NAND2_X1 U2768 ( .A1(n3403), .A2(REG3_REG_15__SCAN_IN), .ZN(n3425) );
  NOR2_X1 U2769 ( .A1(n4978), .A2(n2570), .ZN(n2567) );
  NAND2_X1 U2770 ( .A1(n2572), .A2(n2570), .ZN(n2569) );
  NAND2_X1 U2771 ( .A1(n2617), .A2(n2574), .ZN(n2573) );
  NOR2_X1 U2772 ( .A1(n2617), .A2(n2574), .ZN(n2572) );
  INV_X1 U2773 ( .A(n4989), .ZN(n2579) );
  INV_X1 U2774 ( .A(n2918), .ZN(n2583) );
  INV_X1 U2775 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4116) );
  NOR2_X1 U2776 ( .A1(n4703), .A2(n4279), .ZN(n2637) );
  NAND2_X1 U2777 ( .A1(n2559), .A2(n4457), .ZN(n3807) );
  NAND2_X1 U2778 ( .A1(n4722), .A2(n4462), .ZN(n2559) );
  NOR2_X1 U2779 ( .A1(n3619), .A2(n4325), .ZN(n3626) );
  INV_X1 U2780 ( .A(n3601), .ZN(n2595) );
  NOR2_X1 U2781 ( .A1(n2595), .A2(n2592), .ZN(n2591) );
  INV_X1 U2782 ( .A(n3592), .ZN(n2592) );
  OR2_X1 U2783 ( .A1(n4811), .A2(n4839), .ZN(n3592) );
  NOR2_X1 U2784 ( .A1(n4839), .A2(n4292), .ZN(n2639) );
  NAND2_X1 U2785 ( .A1(n2596), .A2(n2538), .ZN(n3505) );
  INV_X1 U2786 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3905) );
  INV_X1 U2787 ( .A(n3272), .ZN(n2612) );
  OAI21_X1 U2788 ( .B1(n2615), .B2(n2612), .A(n3298), .ZN(n2611) );
  NOR2_X1 U2789 ( .A1(n3202), .A2(n3179), .ZN(n2627) );
  AND2_X1 U2790 ( .A1(n4415), .A2(n3093), .ZN(n4368) );
  AND2_X1 U2791 ( .A1(n4514), .A2(n4426), .ZN(n2815) );
  AND2_X1 U2792 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2653)
         );
  NAND2_X1 U2793 ( .A1(n3125), .A2(n3124), .ZN(n2672) );
  INV_X1 U2794 ( .A(n2680), .ZN(n2679) );
  OAI21_X1 U2795 ( .B1(n4268), .B2(n2681), .A(n5267), .ZN(n2680) );
  INV_X1 U2796 ( .A(n3748), .ZN(n2681) );
  INV_X1 U2797 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3337) );
  NOR2_X1 U2798 ( .A1(n3425), .A2(n4116), .ZN(n3495) );
  XNOR2_X1 U2799 ( .A(n2959), .B(n2960), .ZN(n2981) );
  NOR2_X1 U2800 ( .A1(n3593), .A2(n4271), .ZN(n3602) );
  NAND2_X1 U2801 ( .A1(n3287), .A2(REG3_REG_11__SCAN_IN), .ZN(n3338) );
  AOI21_X1 U2802 ( .B1(n2929), .B2(n2928), .A(n2927), .ZN(n4332) );
  NOR2_X1 U2803 ( .A1(n2935), .A2(n2934), .ZN(n4333) );
  AND2_X1 U2804 ( .A1(n2933), .A2(n2932), .ZN(n2934) );
  NAND2_X1 U2805 ( .A1(n4332), .A2(n4333), .ZN(n4331) );
  INV_X1 U2806 ( .A(n3545), .ZN(n3546) );
  NAND2_X1 U2807 ( .A1(n3546), .A2(REG3_REG_18__SCAN_IN), .ZN(n3593) );
  AND2_X1 U2808 ( .A1(n3526), .A2(n3525), .ZN(n3570) );
  AOI21_X1 U2809 ( .B1(n2682), .B2(n2518), .A(n2683), .ZN(n3574) );
  AND4_X1 U2810 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3174)
         );
  AND4_X1 U2811 ( .A1(n3000), .A2(n2999), .A3(n2998), .A4(n2997), .ZN(n3138)
         );
  NAND4_X1 U2812 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(n3022)
         );
  NAND2_X1 U2813 ( .A1(n2938), .A2(REG1_REG_1__SCAN_IN), .ZN(n2829) );
  NAND2_X1 U2814 ( .A1(n2941), .A2(REG0_REG_1__SCAN_IN), .ZN(n2828) );
  AOI21_X1 U2815 ( .B1(n4959), .B2(REG1_REG_3__SCAN_IN), .A(n2556), .ZN(n2889)
         );
  NAND2_X1 U2816 ( .A1(n4966), .A2(n2914), .ZN(n4590) );
  NAND2_X1 U2817 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  OAI211_X1 U2818 ( .C1(n4590), .C2(n2571), .A(n2568), .B(n2566), .ZN(n4980)
         );
  INV_X1 U2819 ( .A(n2572), .ZN(n2571) );
  AND2_X1 U2820 ( .A1(n2569), .A2(n2573), .ZN(n2568) );
  NAND2_X1 U2821 ( .A1(n4590), .A2(n2567), .ZN(n2566) );
  NAND2_X1 U2822 ( .A1(n4980), .A2(REG2_REG_8__SCAN_IN), .ZN(n4979) );
  INV_X1 U2823 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4313) );
  NOR2_X1 U2824 ( .A1(n4921), .A2(n2579), .ZN(n2576) );
  NAND2_X1 U2825 ( .A1(n2581), .A2(n2579), .ZN(n2578) );
  NAND2_X1 U2826 ( .A1(n2618), .A2(n2583), .ZN(n2582) );
  NOR2_X1 U2827 ( .A1(n2618), .A2(n2583), .ZN(n2581) );
  NAND2_X1 U2828 ( .A1(n4988), .A2(n2918), .ZN(n3011) );
  AOI22_X1 U2829 ( .A1(n4598), .A2(REG1_REG_12__SCAN_IN), .B1(n2544), .B2(
        n4607), .ZN(n5001) );
  NAND2_X1 U2830 ( .A1(n4999), .A2(n4601), .ZN(n2642) );
  XNOR2_X1 U2831 ( .A(n2642), .B(n2619), .ZN(n5014) );
  NAND2_X1 U2832 ( .A1(n5017), .A2(n4610), .ZN(n4614) );
  NOR2_X1 U2833 ( .A1(n4640), .A2(n2527), .ZN(n5029) );
  NAND2_X1 U2834 ( .A1(n4701), .A2(n4690), .ZN(n4692) );
  AND2_X1 U2835 ( .A1(n3658), .A2(n3657), .ZN(n4684) );
  AND2_X1 U2836 ( .A1(n3669), .A2(n3668), .ZN(n4712) );
  NOR2_X1 U2837 ( .A1(n4727), .A2(n2635), .ZN(n4701) );
  INV_X1 U2838 ( .A(n2637), .ZN(n2635) );
  INV_X1 U2839 ( .A(n3826), .ZN(n4279) );
  NOR2_X1 U2840 ( .A1(n4727), .A2(n4279), .ZN(n4700) );
  AOI21_X1 U2841 ( .B1(n2604), .B2(n2609), .A(n2528), .ZN(n2601) );
  INV_X1 U2842 ( .A(n2604), .ZN(n2602) );
  OR2_X1 U2843 ( .A1(n4747), .A2(n3711), .ZN(n4727) );
  AND2_X1 U2844 ( .A1(n4764), .A2(n4765), .ZN(n4767) );
  OR2_X1 U2845 ( .A1(n3610), .A2(n4112), .ZN(n3619) );
  OR2_X1 U2846 ( .A1(n4757), .A2(n3617), .ZN(n4777) );
  NAND2_X1 U2847 ( .A1(n3697), .A2(n4412), .ZN(n4792) );
  AND2_X1 U2848 ( .A1(n3555), .A2(n2638), .ZN(n4797) );
  AND2_X1 U2849 ( .A1(n2520), .A2(n3752), .ZN(n2638) );
  NAND2_X1 U2850 ( .A1(n3555), .A2(n2520), .ZN(n4819) );
  AOI21_X1 U2851 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n4836) );
  NAND2_X1 U2852 ( .A1(n3555), .A2(n3723), .ZN(n4838) );
  INV_X1 U2853 ( .A(n3582), .ZN(n3562) );
  AND2_X1 U2854 ( .A1(n3508), .A2(n3562), .ZN(n3555) );
  NOR2_X1 U2855 ( .A1(n3434), .A2(n3524), .ZN(n3508) );
  NAND2_X1 U2856 ( .A1(n2631), .A2(n2630), .ZN(n2629) );
  INV_X1 U2857 ( .A(n2632), .ZN(n2631) );
  NOR2_X1 U2858 ( .A1(n3413), .A2(n3453), .ZN(n2630) );
  NOR2_X1 U2859 ( .A1(n3338), .A2(n3337), .ZN(n3356) );
  NOR3_X1 U2860 ( .A1(n5145), .A2(n3413), .A3(n2633), .ZN(n5194) );
  OR2_X1 U2861 ( .A1(n3383), .A2(n5141), .ZN(n3466) );
  NOR2_X1 U2862 ( .A1(n5145), .A2(n3413), .ZN(n5146) );
  AND2_X1 U2863 ( .A1(n3381), .A2(n3380), .ZN(n5149) );
  AND2_X1 U2864 ( .A1(n4419), .A2(n3470), .ZN(n4366) );
  OR2_X1 U2865 ( .A1(n5125), .A2(n3382), .ZN(n5145) );
  AND4_X1 U2866 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n4314)
         );
  INV_X1 U2867 ( .A(n4312), .ZN(n3311) );
  AND4_X1 U2868 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n5155)
         );
  INV_X1 U2869 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U2870 ( .A1(n2627), .A2(n3176), .ZN(n3251) );
  NOR2_X1 U2871 ( .A1(n3251), .A2(n3252), .ZN(n3275) );
  AND4_X1 U2872 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3312)
         );
  INV_X1 U2873 ( .A(n2627), .ZN(n2710) );
  INV_X1 U2874 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4117) );
  NOR2_X1 U2875 ( .A1(n3108), .A2(n3090), .ZN(n3201) );
  NAND2_X1 U2876 ( .A1(n3102), .A2(n4335), .ZN(n4428) );
  INV_X1 U2877 ( .A(n5151), .ZN(n5206) );
  OR2_X1 U2878 ( .A1(n2763), .A2(n2848), .ZN(n5154) );
  OR2_X1 U2879 ( .A1(n3164), .A2(n3053), .ZN(n3108) );
  NAND2_X1 U2880 ( .A1(n3156), .A2(n3027), .ZN(n3114) );
  AND2_X1 U2881 ( .A1(n4434), .A2(n4430), .ZN(n4388) );
  INV_X1 U2882 ( .A(n4335), .ZN(n3165) );
  INV_X1 U2883 ( .A(n3041), .ZN(n4389) );
  INV_X1 U2884 ( .A(n3038), .ZN(n4385) );
  MUX2_X1 U2885 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2955), .Z(n4384) );
  AND2_X1 U2886 ( .A1(n3070), .A2(n5057), .ZN(n3166) );
  INV_X1 U2887 ( .A(n4809), .ZN(n5200) );
  INV_X1 U2888 ( .A(n5229), .ZN(n5304) );
  AND2_X1 U2889 ( .A1(n2821), .A2(n2750), .ZN(n2831) );
  OAI21_X1 U2890 ( .B1(n2709), .B2(n4174), .A(n2726), .ZN(n2809) );
  NOR2_X1 U2891 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  XNOR2_X1 U2892 ( .A(n2732), .B(n3975), .ZN(n2753) );
  INV_X1 U2893 ( .A(IR_REG_17__SCAN_IN), .ZN(n3537) );
  OAI21_X2 U2894 ( .B1(n2741), .B2(IR_REG_13__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3379) );
  OR2_X1 U2895 ( .A1(n2879), .A2(n4908), .ZN(n2885) );
  XNOR2_X1 U2896 ( .A(n2584), .B(IR_REG_2__SCAN_IN), .ZN(n4558) );
  OAI21_X1 U2897 ( .B1(n3352), .B2(n2689), .A(n2687), .ZN(n3521) );
  AND4_X1 U2898 ( .A1(n2954), .A2(n2953), .A3(n2952), .A4(n2951), .ZN(n3030)
         );
  NAND2_X1 U2899 ( .A1(n2664), .A2(n2716), .ZN(n2662) );
  NAND2_X1 U2900 ( .A1(n2659), .A2(n2524), .ZN(n2658) );
  AOI21_X1 U2901 ( .B1(n3222), .B2(n3221), .A(n2714), .ZN(n3318) );
  INV_X1 U2902 ( .A(n3070), .ZN(n2838) );
  INV_X1 U2903 ( .A(n4384), .ZN(n5057) );
  INV_X1 U2904 ( .A(n3023), .ZN(n5058) );
  NAND2_X1 U2905 ( .A1(n4266), .A2(n3748), .ZN(n5268) );
  NAND2_X1 U2906 ( .A1(n2686), .A2(n2691), .ZN(n5184) );
  NAND2_X1 U2907 ( .A1(n3352), .A2(n2693), .ZN(n2686) );
  OR3_X1 U2908 ( .A1(n3033), .A2(n2848), .A3(n4895), .ZN(n4345) );
  INV_X1 U2909 ( .A(n4833), .ZN(n4839) );
  NAND2_X1 U2910 ( .A1(n2833), .A2(n5216), .ZN(n5263) );
  INV_X1 U2911 ( .A(n5263), .ZN(n4324) );
  INV_X1 U2912 ( .A(n4358), .ZN(n5272) );
  INV_X1 U2913 ( .A(n4363), .ZN(n5274) );
  INV_X1 U2914 ( .A(n5154), .ZN(n5204) );
  INV_X1 U2915 ( .A(n4405), .ZN(n4520) );
  AND3_X1 U2916 ( .A1(n3677), .A2(n3676), .A3(n3675), .ZN(n3678) );
  OR2_X1 U2917 ( .A1(n3851), .A2(n3680), .ZN(n3679) );
  INV_X1 U2918 ( .A(n4712), .ZN(n4522) );
  INV_X1 U2919 ( .A(n4684), .ZN(n4523) );
  NAND2_X1 U2920 ( .A1(n3649), .A2(n3648), .ZN(n4726) );
  INV_X1 U2921 ( .A(n4407), .ZN(n4524) );
  NAND2_X1 U2922 ( .A1(n3634), .A2(n3633), .ZN(n4763) );
  NAND2_X1 U2923 ( .A1(n3625), .A2(n3624), .ZN(n4525) );
  NAND4_X1 U2924 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n4810)
         );
  INV_X1 U2925 ( .A(n3564), .ZN(n4528) );
  INV_X1 U2926 ( .A(n5155), .ZN(n4533) );
  INV_X1 U2927 ( .A(n3095), .ZN(n4538) );
  INV_X1 U2928 ( .A(n3030), .ZN(n4539) );
  NAND4_X1 U2929 ( .A1(n2945), .A2(n2944), .A3(n2943), .A4(n2942), .ZN(n4540)
         );
  NAND2_X1 U2930 ( .A1(n2938), .A2(REG1_REG_0__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U2931 ( .A1(n4541), .A2(n2907), .ZN(n4563) );
  XNOR2_X1 U2932 ( .A(n2908), .B(n4958), .ZN(n4957) );
  XNOR2_X1 U2933 ( .A(n2889), .B(n5045), .ZN(n5041) );
  NAND2_X1 U2934 ( .A1(n5042), .A2(n2910), .ZN(n4572) );
  NAND2_X1 U2935 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U2936 ( .A1(n4968), .A2(n2895), .ZN(n4585) );
  NAND2_X1 U2937 ( .A1(n4976), .A2(n2898), .ZN(n4987) );
  NAND2_X1 U2938 ( .A1(n4987), .A2(n4986), .ZN(n4985) );
  XNOR2_X1 U2939 ( .A(n2548), .B(n2618), .ZN(n3007) );
  OAI211_X1 U2940 ( .C1(n4990), .C2(n2580), .A(n2577), .B(n2575), .ZN(n2921)
         );
  INV_X1 U2941 ( .A(n2581), .ZN(n2580) );
  AND2_X1 U2942 ( .A1(n2578), .A2(n2582), .ZN(n2577) );
  NAND2_X1 U2943 ( .A1(n4990), .A2(n2576), .ZN(n2575) );
  NAND2_X1 U2944 ( .A1(n2921), .A2(REG2_REG_10__SCAN_IN), .ZN(n3012) );
  NOR2_X1 U2945 ( .A1(n3010), .A2(n2541), .ZN(n3208) );
  AND2_X1 U2946 ( .A1(n3328), .A2(n5161), .ZN(n2545) );
  AND2_X1 U2947 ( .A1(n2547), .A2(n2546), .ZN(n3010) );
  NAND2_X1 U2948 ( .A1(n2548), .A2(n4921), .ZN(n2546) );
  NAND2_X1 U2949 ( .A1(n3007), .A2(REG1_REG_10__SCAN_IN), .ZN(n2547) );
  XNOR2_X1 U2950 ( .A(n2544), .B(n4596), .ZN(n4598) );
  NAND2_X1 U2951 ( .A1(n4608), .A2(n4609), .ZN(n5005) );
  XNOR2_X1 U2952 ( .A(n2620), .B(n2619), .ZN(n5018) );
  NAND2_X1 U2953 ( .A1(n5018), .A2(REG2_REG_14__SCAN_IN), .ZN(n5017) );
  AOI21_X1 U2954 ( .B1(n5014), .B2(REG1_REG_14__SCAN_IN), .A(n2641), .ZN(n4604) );
  AND2_X1 U2955 ( .A1(n2642), .A2(n5016), .ZN(n2641) );
  INV_X1 U2956 ( .A(n4918), .ZN(n5039) );
  NOR2_X1 U2957 ( .A1(n4635), .A2(n4634), .ZN(n5036) );
  NAND2_X1 U2958 ( .A1(n2812), .A2(n2814), .ZN(n4848) );
  AOI21_X1 U2959 ( .B1(n2644), .B2(n2643), .A(n2645), .ZN(n4654) );
  INV_X1 U2960 ( .A(n2646), .ZN(n2645) );
  NOR2_X1 U2961 ( .A1(n4634), .A2(n2648), .ZN(n2643) );
  AND2_X1 U2962 ( .A1(n2920), .A2(n2919), .ZN(n5043) );
  NAND2_X1 U2963 ( .A1(n2605), .A2(n2603), .ZN(n4719) );
  INV_X1 U2964 ( .A(n2606), .ZN(n2603) );
  NAND2_X1 U2965 ( .A1(n4754), .A2(n2608), .ZN(n2605) );
  OAI21_X1 U2966 ( .B1(n4754), .B2(n4756), .A(n2712), .ZN(n4736) );
  NAND2_X1 U2967 ( .A1(n4816), .A2(n3601), .ZN(n4790) );
  INV_X1 U2968 ( .A(n2596), .ZN(n3433) );
  AND2_X1 U2969 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NAND2_X1 U2970 ( .A1(n3275), .A2(n3311), .ZN(n5125) );
  NOR2_X1 U2971 ( .A1(n2614), .A2(n2613), .ZN(n3242) );
  INV_X1 U2972 ( .A(n3240), .ZN(n2613) );
  INV_X1 U2973 ( .A(n3241), .ZN(n2614) );
  NAND2_X1 U2974 ( .A1(n3190), .A2(n3096), .ZN(n3098) );
  INV_X1 U2975 ( .A(n4806), .ZN(n4837) );
  OAI21_X1 U2976 ( .B1(n3038), .B2(n3063), .A(n3062), .ZN(n5072) );
  AND2_X1 U2977 ( .A1(n4843), .A2(n5304), .ZN(n5300) );
  OR2_X1 U2978 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  NAND2_X1 U2979 ( .A1(n2561), .A2(n2560), .ZN(n2585) );
  INV_X1 U2980 ( .A(n4851), .ZN(n2561) );
  AND2_X2 U2981 ( .A1(n4896), .A2(n4895), .ZN(n5312) );
  INV_X1 U2982 ( .A(IR_REG_29__SCAN_IN), .ZN(n2779) );
  INV_X1 U2983 ( .A(n2783), .ZN(n2780) );
  AND2_X1 U2984 ( .A1(n2729), .A2(n2761), .ZN(n4912) );
  AND2_X1 U2985 ( .A1(n2820), .A2(STATE_REG_SCAN_IN), .ZN(n2750) );
  XNOR2_X1 U2986 ( .A(n2765), .B(IR_REG_22__SCAN_IN), .ZN(n4915) );
  AND2_X1 U2987 ( .A1(n2697), .A2(n2734), .ZN(n2764) );
  XNOR2_X1 U2988 ( .A(n2767), .B(IR_REG_21__SCAN_IN), .ZN(n4916) );
  NOR2_X1 U2989 ( .A1(n2701), .A2(n2700), .ZN(n2699) );
  AND2_X1 U2990 ( .A1(n3493), .A2(n3423), .ZN(n4920) );
  OAI21_X1 U2991 ( .B1(n2735), .B2(n4151), .A(n2737), .ZN(n3328) );
  AND2_X1 U2992 ( .A1(n2863), .A2(n2862), .ZN(n4922) );
  AND2_X1 U2993 ( .A1(n2870), .A2(n2869), .ZN(n4923) );
  NOR2_X1 U2994 ( .A1(n2878), .A2(n2877), .ZN(n4924) );
  INV_X1 U2995 ( .A(n4558), .ZN(n4925) );
  NAND2_X1 U2996 ( .A1(n2549), .A2(n2526), .ZN(U3258) );
  NAND2_X1 U2997 ( .A1(n2551), .A2(n2550), .ZN(n2549) );
  NAND2_X2 U2998 ( .A1(n2794), .A2(n2821), .ZN(n3446) );
  INV_X2 U2999 ( .A(n3446), .ZN(n3127) );
  AND2_X1 U3000 ( .A1(n2685), .A2(n3520), .ZN(n2518) );
  INV_X1 U3001 ( .A(n2609), .ZN(n2608) );
  NAND2_X1 U3002 ( .A1(n2537), .A2(n2712), .ZN(n2609) );
  AND2_X1 U3003 ( .A1(n3389), .A2(n3390), .ZN(n2519) );
  INV_X1 U3004 ( .A(n3837), .ZN(n2667) );
  INV_X1 U3005 ( .A(n4408), .ZN(n2599) );
  AND2_X1 U3006 ( .A1(n2639), .A2(n4820), .ZN(n2520) );
  OR3_X1 U3007 ( .A1(n5145), .A2(n2632), .A3(n3413), .ZN(n2521) );
  AND2_X1 U3008 ( .A1(n4661), .A2(n4690), .ZN(n2522) );
  OR2_X1 U3009 ( .A1(n4727), .A2(n2636), .ZN(n2523) );
  NAND2_X1 U3010 ( .A1(n2723), .A2(n4174), .ZN(n2728) );
  NAND2_X1 U3011 ( .A1(n4431), .A2(n4428), .ZN(n3041) );
  NOR2_X1 U3012 ( .A1(n2860), .A2(IR_REG_9__SCAN_IN), .ZN(n2858) );
  OAI21_X1 U3013 ( .B1(n2667), .B2(n2666), .A(n4259), .ZN(n2665) );
  BUF_X1 U3014 ( .A(n3022), .Z(n3023) );
  INV_X1 U3015 ( .A(n4597), .ZN(n2544) );
  NAND4_X1 U3016 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n3039)
         );
  OAI21_X1 U3017 ( .B1(n4754), .B2(n2602), .A(n2601), .ZN(n3802) );
  OR2_X1 U3018 ( .A1(n2663), .A2(n2716), .ZN(n2524) );
  AND2_X1 U3019 ( .A1(n2697), .A2(n2622), .ZN(n2730) );
  AND2_X1 U3020 ( .A1(n4850), .A2(n5257), .ZN(n2525) );
  NAND2_X1 U3021 ( .A1(n2734), .A2(n2699), .ZN(n2766) );
  NOR2_X1 U3022 ( .A1(n4649), .A2(n4648), .ZN(n2526) );
  AND2_X1 U3023 ( .A1(n4641), .A2(n4642), .ZN(n2527) );
  AND2_X1 U3024 ( .A1(n4524), .A2(n3711), .ZN(n2528) );
  NOR2_X1 U3025 ( .A1(n3452), .A2(n3451), .ZN(n2529) );
  AND2_X1 U3026 ( .A1(n2757), .A2(n3983), .ZN(n2530) );
  NAND2_X1 U3027 ( .A1(n5003), .A2(n2621), .ZN(n2620) );
  NAND2_X1 U3028 ( .A1(n3519), .A2(n3518), .ZN(n2531) );
  OAI21_X1 U3029 ( .B1(n2687), .B2(n2684), .A(n2531), .ZN(n2683) );
  INV_X1 U3030 ( .A(n2665), .ZN(n2664) );
  AND3_X1 U3031 ( .A1(n2697), .A2(n2722), .A3(n2622), .ZN(n2723) );
  OR2_X1 U3032 ( .A1(n3316), .A2(n4307), .ZN(n2532) );
  INV_X1 U3033 ( .A(n2714), .ZN(n2675) );
  INV_X1 U3034 ( .A(IR_REG_26__SCAN_IN), .ZN(n2708) );
  INV_X1 U3035 ( .A(IR_REG_7__SCAN_IN), .ZN(n2866) );
  AND2_X1 U3036 ( .A1(n4797), .A2(n4783), .ZN(n4764) );
  AND2_X1 U3037 ( .A1(n3555), .A2(n2639), .ZN(n2533) );
  AND2_X1 U3038 ( .A1(n3564), .A2(n3562), .ZN(n2534) );
  AND2_X1 U3039 ( .A1(n2669), .A2(n2532), .ZN(n3789) );
  INV_X1 U3040 ( .A(n4978), .ZN(n2617) );
  OAI21_X1 U3041 ( .B1(n3352), .B2(n3351), .A(n3350), .ZN(n3445) );
  INV_X1 U3042 ( .A(IR_REG_25__SCAN_IN), .ZN(n4174) );
  AND2_X1 U3043 ( .A1(n4740), .A2(n3699), .ZN(n4756) );
  INV_X1 U3044 ( .A(n4756), .ZN(n2607) );
  OR2_X1 U3045 ( .A1(n4526), .A2(n3618), .ZN(n2535) );
  AND2_X1 U3046 ( .A1(n3841), .A2(n3840), .ZN(n2536) );
  AND4_X1 U3047 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n5201)
         );
  NAND2_X1 U3048 ( .A1(n4763), .A2(n3635), .ZN(n2537) );
  OR2_X1 U3049 ( .A1(n4530), .A2(n3453), .ZN(n2538) );
  NAND2_X1 U3050 ( .A1(n4726), .A2(n4279), .ZN(n2539) );
  OR2_X1 U3051 ( .A1(n5001), .A2(n2713), .ZN(n4999) );
  INV_X1 U3052 ( .A(n2705), .ZN(n2704) );
  NAND2_X1 U3053 ( .A1(n2706), .A2(n3818), .ZN(n2705) );
  NAND2_X2 U3054 ( .A1(n2841), .A2(n4848), .ZN(n3036) );
  AND2_X1 U3055 ( .A1(n4439), .A2(n4437), .ZN(n2540) );
  NAND2_X1 U3056 ( .A1(n3273), .A2(n3272), .ZN(n3299) );
  INV_X1 U3057 ( .A(n4820), .ZN(n4270) );
  NOR2_X1 U3058 ( .A1(n5145), .A2(n2629), .ZN(n2634) );
  OR2_X1 U3059 ( .A1(n3008), .A2(n2545), .ZN(n2541) );
  OR2_X1 U3060 ( .A1(n3372), .A2(n3371), .ZN(n2542) );
  INV_X1 U3061 ( .A(n3752), .ZN(n5262) );
  INV_X1 U3062 ( .A(n5016), .ZN(n2619) );
  INV_X1 U3063 ( .A(n3479), .ZN(n2633) );
  AND2_X1 U3064 ( .A1(n4917), .A2(REG1_REG_18__SCAN_IN), .ZN(n2543) );
  XNOR2_X1 U3065 ( .A(n2762), .B(n2757), .ZN(n2772) );
  INV_X1 U3066 ( .A(n4703), .ZN(n4711) );
  INV_X1 U3067 ( .A(n2648), .ZN(n2647) );
  OR2_X1 U3068 ( .A1(n4638), .A2(n2649), .ZN(n2648) );
  INV_X1 U3069 ( .A(n4921), .ZN(n2618) );
  NOR2_X1 U3070 ( .A1(n2554), .A2(n4919), .ZN(n4634) );
  XNOR2_X1 U3071 ( .A(n2554), .B(n4919), .ZN(n4623) );
  AND2_X1 U3072 ( .A1(n4920), .A2(REG1_REG_15__SCAN_IN), .ZN(n2555) );
  AND2_X1 U3073 ( .A1(n2558), .A2(n4958), .ZN(n2556) );
  XNOR2_X1 U3074 ( .A(n2558), .B(n2557), .ZN(n4959) );
  INV_X1 U3075 ( .A(n4958), .ZN(n2557) );
  NAND2_X1 U3076 ( .A1(n4564), .A2(n2884), .ZN(n2558) );
  AND3_X2 U3077 ( .A1(n4132), .A2(n3944), .A3(n2866), .ZN(n2719) );
  OAI21_X2 U3078 ( .B1(n4792), .B2(n4793), .A(n4487), .ZN(n4778) );
  NAND2_X1 U3079 ( .A1(n4562), .A2(n4563), .ZN(n4561) );
  NOR2_X1 U3080 ( .A1(n2880), .A2(n4908), .ZN(n2584) );
  NAND2_X2 U3081 ( .A1(n4682), .A2(n4688), .ZN(n4681) );
  MUX2_X1 U3082 ( .A(REG1_REG_29__SCAN_IN), .B(n2585), .S(n5308), .Z(U3547) );
  MUX2_X1 U3083 ( .A(REG0_REG_29__SCAN_IN), .B(n2585), .S(n5312), .Z(U3515) );
  MUX2_X1 U3084 ( .A(n2906), .B(n3894), .S(n2955), .Z(n3070) );
  XNOR2_X2 U3085 ( .A(n2586), .B(n3983), .ZN(n2763) );
  NAND3_X1 U3086 ( .A1(n3959), .A2(n4156), .A3(n4161), .ZN(n2587) );
  NAND4_X1 U3087 ( .A1(n2589), .A2(n2742), .A3(n4160), .A4(n2746), .ZN(n2588)
         );
  NAND2_X1 U3088 ( .A1(n4834), .A2(n2591), .ZN(n2590) );
  NAND3_X1 U3089 ( .A1(n3190), .A2(n3096), .A3(n3097), .ZN(n3181) );
  NOR2_X2 U3090 ( .A1(n2860), .A2(n2625), .ZN(n2734) );
  NOR2_X2 U3091 ( .A1(n2860), .A2(n2623), .ZN(n2622) );
  INV_X1 U3092 ( .A(n2634), .ZN(n3434) );
  INV_X1 U3093 ( .A(n4635), .ZN(n2644) );
  MUX2_X1 U3094 ( .A(n2882), .B(REG1_REG_1__SCAN_IN), .S(n2906), .Z(n4545) );
  AND2_X1 U3095 ( .A1(n2654), .A2(n2926), .ZN(n2927) );
  XNOR2_X1 U3096 ( .A(n2654), .B(n2925), .ZN(n2929) );
  NAND2_X1 U3097 ( .A1(n4350), .A2(n2656), .ZN(n2655) );
  OAI211_X1 U3098 ( .C1(n4350), .C2(n2662), .A(n2658), .B(n2655), .ZN(n3854)
         );
  OAI21_X1 U3099 ( .B1(n4350), .B2(n3838), .A(n3837), .ZN(n4258) );
  INV_X1 U3100 ( .A(n3221), .ZN(n2674) );
  OAI21_X1 U3101 ( .B1(n3146), .B2(n3145), .A(n2672), .ZN(n3222) );
  OAI211_X1 U3102 ( .C1(n3146), .C2(n2673), .A(n3317), .B(n2670), .ZN(n2669)
         );
  INV_X1 U3103 ( .A(n2671), .ZN(n2670) );
  OAI21_X1 U3104 ( .B1(n2674), .B2(n2672), .A(n2675), .ZN(n2671) );
  INV_X1 U3105 ( .A(n3352), .ZN(n2682) );
  NAND2_X1 U3106 ( .A1(n2734), .A2(n2720), .ZN(n2741) );
  OAI21_X1 U3107 ( .B1(n4322), .B2(n2705), .A(n2702), .ZN(n4297) );
  NAND2_X1 U3108 ( .A1(n2891), .A2(n2890), .ZN(n4575) );
  AOI211_X2 U3109 ( .C1(n4809), .C2(n4520), .A(n3710), .B(n3709), .ZN(n4861)
         );
  NAND2_X1 U3110 ( .A1(n3301), .A2(n3300), .ZN(n3372) );
  XNOR2_X1 U3111 ( .A(n3022), .B(n3070), .ZN(n3038) );
  OR2_X1 U3112 ( .A1(n2723), .A2(n4908), .ZN(n2709) );
  INV_X1 U3113 ( .A(n3310), .ZN(n3845) );
  AND2_X1 U3114 ( .A1(n3572), .A2(n3571), .ZN(n2711) );
  NAND2_X1 U3115 ( .A1(n3507), .A2(n3506), .ZN(n3554) );
  OR2_X1 U3116 ( .A1(n3765), .A2(n4765), .ZN(n2712) );
  AND4_X1 U3117 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3523)
         );
  OR2_X1 U3118 ( .A1(n4600), .A2(n4599), .ZN(n2713) );
  AND2_X1 U3119 ( .A1(n3220), .A2(n3219), .ZN(n2714) );
  AND2_X1 U3120 ( .A1(n3119), .A2(n3118), .ZN(n2715) );
  INV_X1 U3121 ( .A(n3456), .ZN(n2837) );
  XOR2_X1 U3122 ( .A(n3847), .B(n3846), .Z(n2716) );
  INV_X1 U3123 ( .A(n4601), .ZN(n4599) );
  AND2_X1 U3124 ( .A1(n3397), .A2(n3400), .ZN(n4450) );
  AND2_X1 U3125 ( .A1(n3695), .A2(n3690), .ZN(n4483) );
  INV_X1 U3126 ( .A(n5153), .ZN(n3413) );
  INV_X1 U3127 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4093) );
  AND2_X1 U3128 ( .A1(n3626), .A2(REG3_REG_23__SCAN_IN), .ZN(n3636) );
  NOR2_X1 U3129 ( .A1(n3373), .A2(n3905), .ZN(n3403) );
  INV_X1 U3130 ( .A(n2940), .ZN(n3666) );
  OR2_X1 U3131 ( .A1(n3131), .A2(n3916), .ZN(n3228) );
  NAND2_X1 U3132 ( .A1(n2937), .A2(REG3_REG_2__SCAN_IN), .ZN(n2852) );
  AND2_X1 U3133 ( .A1(n4908), .A2(n4174), .ZN(n2724) );
  OR2_X1 U3134 ( .A1(n3077), .A2(n4093), .ZN(n3131) );
  INV_X1 U3135 ( .A(n4525), .ZN(n3765) );
  INV_X1 U3136 ( .A(n3196), .ZN(n3200) );
  OAI22_X1 U3137 ( .A1(n2854), .A2(n3446), .B1(n5057), .B2(n3456), .ZN(n2845)
         );
  OR2_X1 U3138 ( .A1(n4350), .A2(n4349), .ZN(n4352) );
  OR2_X1 U3139 ( .A1(n4694), .A2(n3680), .ZN(n3669) );
  OR2_X1 U3140 ( .A1(n4731), .A2(n3680), .ZN(n3643) );
  INV_X1 U3141 ( .A(n4856), .ZN(n2832) );
  NOR2_X1 U3142 ( .A1(n2967), .A2(n4117), .ZN(n2995) );
  AND2_X1 U3143 ( .A1(n2831), .A2(n2824), .ZN(n4859) );
  AND2_X1 U3144 ( .A1(n3261), .A2(REG3_REG_10__SCAN_IN), .ZN(n3287) );
  INV_X1 U3145 ( .A(n5279), .ZN(n4317) );
  NAND2_X1 U3146 ( .A1(n3356), .A2(REG3_REG_13__SCAN_IN), .ZN(n3373) );
  AND2_X1 U3147 ( .A1(n3686), .A2(n3685), .ZN(n4405) );
  OR2_X1 U31480 ( .A1(n4768), .A2(n3680), .ZN(n3625) );
  AND4_X1 U31490 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3564)
         );
  OR2_X1 U3150 ( .A1(n2966), .A2(n2939), .ZN(n2944) );
  INV_X1 U3151 ( .A(n5009), .ZN(n5046) );
  INV_X1 U3152 ( .A(n5049), .ZN(n5033) );
  AND2_X1 U3153 ( .A1(n4849), .A2(n2815), .ZN(n5283) );
  NAND2_X1 U3154 ( .A1(n3047), .A2(n3046), .ZN(n5151) );
  AND2_X1 U3155 ( .A1(n5173), .A2(n4848), .ZN(n4843) );
  AND2_X1 U3156 ( .A1(n2763), .A2(n2853), .ZN(n4809) );
  INV_X1 U3157 ( .A(n5257), .ZN(n5111) );
  OR3_X1 U3158 ( .A1(n3270), .A2(n3269), .A3(n3268), .ZN(n5128) );
  OAI21_X1 U3159 ( .B1(n4855), .B2(D_REG_0__SCAN_IN), .A(n2796), .ZN(n4895) );
  INV_X1 U3160 ( .A(n2750), .ZN(n2754) );
  NAND2_X1 U3161 ( .A1(n2752), .A2(n4912), .ZN(n4855) );
  OR2_X1 U3162 ( .A1(n2876), .A2(IR_REG_6__SCAN_IN), .ZN(n2872) );
  AND2_X1 U3163 ( .A1(n2771), .A2(n2775), .ZN(n5053) );
  NAND2_X1 U3164 ( .A1(n2973), .A2(STATE_REG_SCAN_IN), .ZN(n5279) );
  NAND2_X1 U3165 ( .A1(n3679), .A2(n3678), .ZN(n4521) );
  OR2_X1 U3166 ( .A1(n2900), .A2(n4911), .ZN(n5049) );
  NAND2_X2 U3167 ( .A1(n3034), .A2(n5216), .ZN(n5173) );
  NAND2_X1 U3168 ( .A1(n5173), .A2(n5165), .ZN(n4806) );
  OR2_X1 U3169 ( .A1(n4894), .A2(n4895), .ZN(n5306) );
  INV_X2 U3170 ( .A(n5306), .ZN(n5308) );
  AND2_X1 U3171 ( .A1(n5116), .A2(n5115), .ZN(n5118) );
  INV_X1 U3172 ( .A(n5312), .ZN(n5309) );
  AND2_X1 U3173 ( .A1(n2873), .A2(n2872), .ZN(n4970) );
  INV_X2 U3174 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND4_X2 U3175 ( .A1(n2719), .A2(n2880), .A3(n2718), .A4(n2717), .ZN(n2860)
         );
  INV_X1 U3176 ( .A(n2809), .ZN(n4913) );
  NAND2_X1 U3177 ( .A1(n2728), .A2(IR_REG_31__SCAN_IN), .ZN(n2727) );
  MUX2_X1 U3178 ( .A(IR_REG_31__SCAN_IN), .B(n2727), .S(IR_REG_26__SCAN_IN), 
        .Z(n2729) );
  NAND2_X1 U3179 ( .A1(n2733), .A2(n3974), .ZN(n2731) );
  NAND2_X1 U3180 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2732) );
  INV_X1 U3181 ( .A(n2753), .ZN(n4914) );
  XNOR2_X1 U3182 ( .A(n2733), .B(n3974), .ZN(n2820) );
  NOR2_X4 U3183 ( .A1(n2821), .A2(n2754), .ZN(U4043) );
  OR2_X1 U3184 ( .A1(n2734), .A2(n4908), .ZN(n2735) );
  NAND2_X1 U3185 ( .A1(n2735), .A2(n4151), .ZN(n2737) );
  INV_X1 U3186 ( .A(DATAI_11_), .ZN(n3327) );
  MUX2_X1 U3187 ( .A(n3328), .B(n3327), .S(U3149), .Z(n2736) );
  INV_X1 U3188 ( .A(n2736), .ZN(U3341) );
  NAND2_X1 U3189 ( .A1(n2737), .A2(IR_REG_31__SCAN_IN), .ZN(n2738) );
  INV_X1 U3190 ( .A(IR_REG_12__SCAN_IN), .ZN(n4152) );
  XNOR2_X1 U3191 ( .A(n2738), .B(n4152), .ZN(n4596) );
  INV_X1 U3192 ( .A(DATAI_12_), .ZN(n4073) );
  MUX2_X1 U3193 ( .A(n4596), .B(n4073), .S(U3149), .Z(n2739) );
  INV_X1 U3194 ( .A(n2739), .ZN(U3340) );
  INV_X1 U3195 ( .A(DATAI_23_), .ZN(n2740) );
  AOI21_X1 U3196 ( .B1(n2740), .B2(U3149), .A(n2750), .ZN(U3329) );
  INV_X1 U3197 ( .A(DATAI_20_), .ZN(n2748) );
  NAND2_X1 U3198 ( .A1(n3379), .A2(n3959), .ZN(n3420) );
  NAND2_X1 U3199 ( .A1(n3421), .A2(n2742), .ZN(n2743) );
  NOR2_X2 U3200 ( .A1(n3420), .A2(n2743), .ZN(n3536) );
  NAND2_X1 U3201 ( .A1(n3536), .A2(n3537), .ZN(n3535) );
  INV_X1 U3202 ( .A(n3535), .ZN(n2744) );
  NAND2_X1 U3203 ( .A1(n2744), .A2(n4160), .ZN(n2745) );
  NAND2_X1 U3204 ( .A1(n2813), .A2(n4161), .ZN(n2812) );
  MUX2_X1 U3205 ( .A(n2748), .B(n2517), .S(STATE_REG_SCAN_IN), .Z(n2749) );
  INV_X1 U3206 ( .A(n2749), .ZN(U3332) );
  NAND2_X1 U3207 ( .A1(n2809), .A2(n2753), .ZN(n2751) );
  MUX2_X1 U3208 ( .A(n2753), .B(n2751), .S(B_REG_SCAN_IN), .Z(n2752) );
  NAND2_X1 U3209 ( .A1(n2831), .A2(n4855), .ZN(n4951) );
  INV_X1 U32100 ( .A(D_REG_0__SCAN_IN), .ZN(n2756) );
  INV_X1 U32110 ( .A(n4912), .ZN(n2808) );
  NAND2_X1 U32120 ( .A1(n2808), .A2(n2753), .ZN(n2796) );
  NOR2_X1 U32130 ( .A1(n2796), .A2(n2754), .ZN(n2755) );
  AOI21_X1 U32140 ( .B1(n4951), .B2(n2756), .A(n2755), .ZN(U3458) );
  INV_X1 U32150 ( .A(DATAI_28_), .ZN(n2759) );
  INV_X1 U32160 ( .A(IR_REG_27__SCAN_IN), .ZN(n2757) );
  INV_X1 U32170 ( .A(n2763), .ZN(n4553) );
  MUX2_X1 U32180 ( .A(n2759), .B(n2763), .S(STATE_REG_SCAN_IN), .Z(n2760) );
  INV_X1 U32190 ( .A(n2760), .ZN(U3324) );
  OR2_X1 U32200 ( .A1(n2764), .A2(n4908), .ZN(n2765) );
  NAND2_X1 U32210 ( .A1(n2766), .A2(IR_REG_31__SCAN_IN), .ZN(n2767) );
  NAND2_X1 U32220 ( .A1(n2820), .A2(n2853), .ZN(n2768) );
  AND2_X1 U32230 ( .A1(n4404), .A2(n2768), .ZN(n2774) );
  INV_X1 U32240 ( .A(n2774), .ZN(n2771) );
  INV_X1 U32250 ( .A(n2831), .ZN(n2770) );
  NOR2_X1 U32260 ( .A1(n2820), .A2(U3149), .ZN(n4517) );
  INV_X1 U32270 ( .A(n4517), .ZN(n2769) );
  NAND2_X1 U32280 ( .A1(n2770), .A2(n2769), .ZN(n2775) );
  NOR2_X1 U32290 ( .A1(n5053), .A2(U4043), .ZN(U3148) );
  INV_X1 U32300 ( .A(n2772), .ZN(n4911) );
  INV_X1 U32310 ( .A(REG2_REG_0__SCAN_IN), .ZN(n5070) );
  AOI21_X1 U32320 ( .B1(n4911), .B2(n5070), .A(n2763), .ZN(n4557) );
  OAI21_X1 U32330 ( .B1(n4911), .B2(REG1_REG_0__SCAN_IN), .A(n4557), .ZN(n2773) );
  XOR2_X1 U32340 ( .A(IR_REG_0__SCAN_IN), .B(n2773), .Z(n2777) );
  AND2_X1 U32350 ( .A1(n2775), .A2(n2774), .ZN(n2920) );
  INV_X1 U32360 ( .A(n2920), .ZN(n2900) );
  AOI22_X1 U32370 ( .A1(n5053), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2776) );
  OAI21_X1 U32380 ( .B1(n2777), .B2(n2900), .A(n2776), .ZN(U3240) );
  NAND2_X1 U32390 ( .A1(n2780), .A2(n2779), .ZN(n2782) );
  XNOR2_X2 U32400 ( .A(n2781), .B(IR_REG_30__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U32410 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  NOR2_X2 U32420 ( .A1(n4910), .A2(n2787), .ZN(n2938) );
  INV_X1 U32430 ( .A(n2787), .ZN(n2786) );
  NOR2_X2 U32440 ( .A1(n2786), .A2(n4910), .ZN(n2941) );
  NAND2_X1 U32450 ( .A1(n2941), .A2(REG0_REG_0__SCAN_IN), .ZN(n2790) );
  AND2_X4 U32460 ( .A1(n4910), .A2(n2787), .ZN(n2940) );
  NAND2_X1 U32470 ( .A1(n2940), .A2(REG2_REG_0__SCAN_IN), .ZN(n2789) );
  AND2_X2 U32480 ( .A1(n2786), .A2(n4910), .ZN(n2937) );
  NAND2_X1 U32490 ( .A1(n2937), .A2(REG3_REG_0__SCAN_IN), .ZN(n2788) );
  NAND2_X2 U32500 ( .A1(n2516), .A2(n4916), .ZN(n2842) );
  NAND2_X2 U32510 ( .A1(n2842), .A2(n2821), .ZN(n3456) );
  INV_X1 U32520 ( .A(n4915), .ZN(n4514) );
  INV_X1 U32530 ( .A(n4916), .ZN(n4426) );
  NAND2_X2 U32540 ( .A1(n2517), .A2(n2815), .ZN(n5229) );
  INV_X1 U32550 ( .A(n2842), .ZN(n2794) );
  INV_X1 U32560 ( .A(n2821), .ZN(n2795) );
  AOI222_X1 U32570 ( .A1(n3039), .A2(n3828), .B1(n4384), .B2(n3310), .C1(
        IR_REG_0__SCAN_IN), .C2(n2795), .ZN(n2846) );
  XNOR2_X1 U32580 ( .A(n2846), .B(n2847), .ZN(n4551) );
  INV_X1 U32590 ( .A(n4895), .ZN(n3032) );
  INV_X1 U32600 ( .A(n4855), .ZN(n4854) );
  NOR4_X1 U32610 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2800) );
  NOR4_X1 U32620 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2799) );
  NOR4_X1 U32630 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2798) );
  NOR4_X1 U32640 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2797) );
  AND4_X1 U32650 ( .A1(n2800), .A2(n2799), .A3(n2798), .A4(n2797), .ZN(n2806)
         );
  NOR2_X1 U32660 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_24__SCAN_IN), .ZN(n2804)
         );
  NOR4_X1 U32670 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2803) );
  NOR4_X1 U32680 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2802) );
  NOR4_X1 U32690 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2801) );
  AND4_X1 U32700 ( .A1(n2804), .A2(n2803), .A3(n2802), .A4(n2801), .ZN(n2805)
         );
  NAND2_X1 U32710 ( .A1(n2806), .A2(n2805), .ZN(n4853) );
  INV_X1 U32720 ( .A(n4853), .ZN(n2807) );
  NAND2_X1 U32730 ( .A1(n2807), .A2(D_REG_1__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U32740 ( .A1(n2809), .A2(n2808), .ZN(n4907) );
  INV_X1 U32750 ( .A(n4907), .ZN(n2810) );
  AOI21_X1 U32760 ( .B1(n4854), .B2(n2811), .A(n2810), .ZN(n2825) );
  NAND3_X1 U32770 ( .A1(n3032), .A2(n2831), .A3(n2825), .ZN(n2830) );
  INV_X1 U32780 ( .A(n2517), .ZN(n4849) );
  OR2_X1 U32790 ( .A1(n2813), .A2(n4161), .ZN(n2814) );
  INV_X1 U32800 ( .A(n2815), .ZN(n5056) );
  NOR2_X1 U32810 ( .A1(n4848), .A2(n5056), .ZN(n2816) );
  OR3_X1 U32820 ( .A1(n5283), .A2(n2853), .A3(n2816), .ZN(n2817) );
  NAND2_X1 U32830 ( .A1(n3032), .A2(n2825), .ZN(n2818) );
  NAND2_X1 U32840 ( .A1(n2818), .A2(n4856), .ZN(n2823) );
  NAND2_X1 U32850 ( .A1(n2517), .A2(n4848), .ZN(n2819) );
  NAND2_X1 U32860 ( .A1(n2819), .A2(n2853), .ZN(n2824) );
  AND3_X1 U32870 ( .A1(n2824), .A2(n2821), .A3(n2820), .ZN(n2822) );
  NAND2_X1 U32880 ( .A1(n2823), .A2(n2822), .ZN(n2973) );
  OR2_X1 U32890 ( .A1(n2973), .A2(U3149), .ZN(n4336) );
  NAND2_X1 U32900 ( .A1(n2825), .A2(n4859), .ZN(n3033) );
  INV_X1 U32910 ( .A(n2853), .ZN(n2848) );
  NOR2_X2 U32920 ( .A1(n4345), .A2(n4553), .ZN(n4358) );
  NAND2_X1 U32930 ( .A1(n2937), .A2(REG3_REG_1__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U32940 ( .A1(n2940), .A2(REG2_REG_1__SCAN_IN), .ZN(n2826) );
  OR2_X1 U32950 ( .A1(n2830), .A2(n5293), .ZN(n2833) );
  OAI22_X1 U32960 ( .A1(n5272), .A2(n5058), .B1(n4324), .B2(n5057), .ZN(n2834)
         );
  AOI21_X1 U32970 ( .B1(REG3_REG_0__SCAN_IN), .B2(n4336), .A(n2834), .ZN(n2835) );
  OAI21_X1 U32980 ( .B1(n4551), .B2(n4363), .A(n2835), .ZN(U3229) );
  NAND2_X1 U32990 ( .A1(n3023), .A2(n3310), .ZN(n2840) );
  INV_X1 U33000 ( .A(n2880), .ZN(n2836) );
  INV_X1 U33010 ( .A(DATAI_1_), .ZN(n3894) );
  NAND2_X1 U33020 ( .A1(n2840), .A2(n2839), .ZN(n2843) );
  NAND2_X4 U33030 ( .A1(n3036), .A2(n2842), .ZN(n3843) );
  NOR2_X1 U33040 ( .A1(n3070), .A2(n3446), .ZN(n2844) );
  OAI22_X1 U33050 ( .A1(n2847), .A2(n2846), .B1(n3843), .B2(n2845), .ZN(n2928)
         );
  XNOR2_X1 U33060 ( .A(n2929), .B(n2928), .ZN(n2857) );
  NAND2_X1 U33070 ( .A1(n2938), .A2(REG1_REG_2__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U33080 ( .A1(n2940), .A2(REG2_REG_2__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U33090 ( .A1(n2941), .A2(REG0_REG_2__SCAN_IN), .ZN(n2849) );
  OAI22_X1 U33100 ( .A1(n2854), .A2(n5154), .B1(n3102), .B2(n5200), .ZN(n3067)
         );
  INV_X1 U33110 ( .A(n4345), .ZN(n3798) );
  AOI22_X1 U33120 ( .A1(n3067), .A2(n3798), .B1(REG3_REG_1__SCAN_IN), .B2(
        n4336), .ZN(n2856) );
  NAND2_X1 U33130 ( .A1(n5263), .A2(n2838), .ZN(n2855) );
  OAI211_X1 U33140 ( .C1(n2857), .C2(n4363), .A(n2856), .B(n2855), .ZN(U3219)
         );
  OR2_X1 U33150 ( .A1(n2858), .A2(n4908), .ZN(n2859) );
  XNOR2_X1 U33160 ( .A(n2859), .B(IR_REG_10__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U33170 ( .A1(n2860), .A2(IR_REG_31__SCAN_IN), .ZN(n2861) );
  MUX2_X1 U33180 ( .A(IR_REG_31__SCAN_IN), .B(n2861), .S(IR_REG_9__SCAN_IN), 
        .Z(n2863) );
  INV_X1 U33190 ( .A(n2858), .ZN(n2862) );
  NAND2_X1 U33200 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4922), .ZN(n2899) );
  INV_X1 U33210 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2864) );
  MUX2_X1 U33220 ( .A(REG1_REG_9__SCAN_IN), .B(n2864), .S(n4922), .Z(n4986) );
  AND2_X1 U33230 ( .A1(n2880), .A2(n4132), .ZN(n2879) );
  NOR2_X1 U33240 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2865)
         );
  NAND2_X1 U33250 ( .A1(n2874), .A2(n4140), .ZN(n2876) );
  NAND2_X1 U33260 ( .A1(n2872), .A2(IR_REG_31__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U33270 ( .A1(n2868), .A2(n2866), .ZN(n2869) );
  NAND2_X1 U33280 ( .A1(n2869), .A2(IR_REG_31__SCAN_IN), .ZN(n2867) );
  XNOR2_X1 U33290 ( .A(n2867), .B(IR_REG_8__SCAN_IN), .ZN(n4978) );
  OR2_X1 U33300 ( .A1(n2868), .A2(n2866), .ZN(n2870) );
  NAND2_X1 U33310 ( .A1(n2876), .A2(IR_REG_31__SCAN_IN), .ZN(n2871) );
  MUX2_X1 U33320 ( .A(IR_REG_31__SCAN_IN), .B(n2871), .S(IR_REG_6__SCAN_IN), 
        .Z(n2873) );
  NOR2_X1 U33330 ( .A1(n2874), .A2(n4908), .ZN(n2875) );
  MUX2_X1 U33340 ( .A(n4908), .B(n2875), .S(IR_REG_5__SCAN_IN), .Z(n2878) );
  INV_X1 U33350 ( .A(n2876), .ZN(n2877) );
  NAND2_X1 U33360 ( .A1(n4924), .A2(REG1_REG_5__SCAN_IN), .ZN(n2893) );
  XNOR2_X1 U33370 ( .A(n2885), .B(IR_REG_3__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U33380 ( .A1(REG1_REG_2__SCAN_IN), .A2(n4925), .ZN(n2884) );
  INV_X1 U33390 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2881) );
  MUX2_X1 U33400 ( .A(REG1_REG_2__SCAN_IN), .B(n2881), .S(n4925), .Z(n4565) );
  INV_X1 U33410 ( .A(n2906), .ZN(n4926) );
  NAND2_X1 U33420 ( .A1(REG1_REG_1__SCAN_IN), .A2(n4926), .ZN(n2883) );
  INV_X1 U33430 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2882) );
  NAND3_X1 U33440 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .A3(
        n4545), .ZN(n4544) );
  NAND2_X1 U33450 ( .A1(n2883), .A2(n4544), .ZN(n4566) );
  NAND2_X1 U33460 ( .A1(n4565), .A2(n4566), .ZN(n4564) );
  INV_X1 U33470 ( .A(IR_REG_3__SCAN_IN), .ZN(n3936) );
  NAND2_X1 U33480 ( .A1(n2885), .A2(n3936), .ZN(n2886) );
  NAND2_X1 U33490 ( .A1(n2886), .A2(IR_REG_31__SCAN_IN), .ZN(n2887) );
  XNOR2_X1 U33500 ( .A(n2887), .B(IR_REG_4__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U33510 ( .A1(n5041), .A2(REG1_REG_4__SCAN_IN), .ZN(n2891) );
  INV_X1 U33520 ( .A(n5045), .ZN(n2888) );
  OR2_X1 U3353 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  INV_X1 U33540 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2892) );
  MUX2_X1 U3355 ( .A(REG1_REG_5__SCAN_IN), .B(n2892), .S(n4924), .Z(n4574) );
  NAND2_X1 U3356 ( .A1(n4575), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U3357 ( .A1(n2893), .A2(n4573), .ZN(n2894) );
  NAND2_X1 U3358 ( .A1(n4970), .A2(n2894), .ZN(n2895) );
  INV_X1 U3359 ( .A(n4970), .ZN(n2913) );
  XNOR2_X1 U3360 ( .A(n2913), .B(n2894), .ZN(n4969) );
  NAND2_X1 U3361 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4969), .ZN(n4968) );
  NAND2_X1 U3362 ( .A1(n4923), .A2(REG1_REG_7__SCAN_IN), .ZN(n2896) );
  NAND2_X1 U3363 ( .A1(n4978), .A2(n2897), .ZN(n2898) );
  NAND2_X1 U3364 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4977), .ZN(n4976) );
  XNOR2_X1 U3365 ( .A(n3007), .B(REG1_REG_10__SCAN_IN), .ZN(n2924) );
  AND2_X1 U3366 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U3367 ( .A1(n2920), .A2(n2763), .ZN(n5009) );
  NOR2_X1 U3368 ( .A1(n5009), .A2(n2618), .ZN(n2901) );
  AOI211_X1 U3369 ( .C1(n5053), .C2(ADDR_REG_10__SCAN_IN), .A(n3796), .B(n2901), .ZN(n2923) );
  NAND2_X1 U3370 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4922), .ZN(n2918) );
  INV_X1 U3371 ( .A(n4922), .ZN(n4993) );
  INV_X1 U3372 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U3373 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4922), .B1(n4993), .B2(n3277), .ZN(n4989) );
  NAND2_X1 U3374 ( .A1(n4923), .A2(REG2_REG_7__SCAN_IN), .ZN(n2915) );
  INV_X1 U3375 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2902) );
  MUX2_X1 U3376 ( .A(REG2_REG_7__SCAN_IN), .B(n2902), .S(n4923), .Z(n4589) );
  NAND2_X1 U3377 ( .A1(n4924), .A2(REG2_REG_5__SCAN_IN), .ZN(n2911) );
  INV_X1 U3378 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2903) );
  MUX2_X1 U3379 ( .A(n2903), .B(REG2_REG_5__SCAN_IN), .S(n4924), .Z(n2904) );
  INV_X1 U3380 ( .A(n2904), .ZN(n4571) );
  INV_X1 U3381 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2905) );
  AOI22_X1 U3382 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4925), .B1(n4558), .B2(n2905), .ZN(n4562) );
  NAND2_X1 U3383 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4926), .ZN(n2907) );
  AOI22_X1 U3384 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4926), .B1(n2906), .B2(n3072), .ZN(n4542) );
  NAND3_X1 U3385 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .A3(n4542), .ZN(n4541) );
  OAI21_X1 U3386 ( .B1(n2557), .B2(n2908), .A(n4956), .ZN(n2909) );
  NAND2_X1 U3387 ( .A1(n5045), .A2(n2909), .ZN(n2910) );
  NAND2_X1 U3388 ( .A1(n2911), .A2(n4570), .ZN(n2912) );
  NAND2_X1 U3389 ( .A1(n4970), .A2(n2912), .ZN(n2914) );
  XNOR2_X1 U3390 ( .A(n2913), .B(n2912), .ZN(n4967) );
  NAND2_X1 U3391 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4967), .ZN(n4966) );
  NAND2_X1 U3392 ( .A1(n4978), .A2(n2916), .ZN(n2917) );
  NOR2_X1 U3393 ( .A1(n2763), .A2(n2772), .ZN(n2919) );
  OAI211_X1 U3394 ( .C1(n2921), .C2(REG2_REG_10__SCAN_IN), .A(n5043), .B(n3012), .ZN(n2922) );
  OAI211_X1 U3395 ( .C1(n2924), .C2(n5049), .A(n2923), .B(n2922), .ZN(U3250)
         );
  INV_X1 U3396 ( .A(n2925), .ZN(n2926) );
  MUX2_X1 U3397 ( .A(n4925), .B(DATAI_2_), .S(n2955), .Z(n4335) );
  XNOR2_X1 U3398 ( .A(n2930), .B(n3843), .ZN(n2932) );
  INV_X2 U3399 ( .A(n3828), .ZN(n3842) );
  NAND2_X1 U3400 ( .A1(n4335), .A2(n3127), .ZN(n2931) );
  NOR2_X1 U3401 ( .A1(n2932), .A2(n2933), .ZN(n2935) );
  INV_X1 U3402 ( .A(n2935), .ZN(n2936) );
  NAND2_X1 U3403 ( .A1(n4331), .A2(n2936), .ZN(n2980) );
  INV_X1 U3404 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U3405 ( .A1(n2937), .A2(n4101), .ZN(n2945) );
  INV_X1 U3406 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2939) );
  NAND2_X1 U3407 ( .A1(n2940), .A2(REG2_REG_3__SCAN_IN), .ZN(n2943) );
  NAND2_X1 U3408 ( .A1(n2941), .A2(REG0_REG_3__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3409 ( .A1(n4540), .A2(n3127), .ZN(n2947) );
  MUX2_X1 U3410 ( .A(n4958), .B(DATAI_3_), .S(n4404), .Z(n3053) );
  NAND2_X1 U3411 ( .A1(n3053), .A2(n2837), .ZN(n2946) );
  INV_X1 U3412 ( .A(n3053), .ZN(n3109) );
  OAI22_X1 U3413 ( .A1(n3159), .A2(n3842), .B1(n3109), .B2(n3845), .ZN(n2949)
         );
  INV_X1 U3414 ( .A(n2949), .ZN(n2960) );
  NAND2_X1 U3415 ( .A1(n2980), .A2(n2981), .ZN(n2963) );
  NAND2_X1 U3416 ( .A1(n3130), .A2(REG1_REG_4__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U3417 ( .A1(n2940), .A2(REG2_REG_4__SCAN_IN), .ZN(n2953) );
  INV_X1 U3418 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4125) );
  NAND2_X1 U3419 ( .A1(n4125), .A2(n4101), .ZN(n2950) );
  NAND2_X1 U3420 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2967) );
  AND2_X1 U3421 ( .A1(n2950), .A2(n2967), .ZN(n2974) );
  NAND2_X1 U3422 ( .A1(n2937), .A2(n2974), .ZN(n2952) );
  NAND2_X1 U3423 ( .A1(n2941), .A2(REG0_REG_4__SCAN_IN), .ZN(n2951) );
  MUX2_X1 U3424 ( .A(n5045), .B(DATAI_4_), .S(n2955), .Z(n3090) );
  INV_X1 U3425 ( .A(n3090), .ZN(n3037) );
  XNOR2_X1 U3427 ( .A(n2956), .B(n3824), .ZN(n2987) );
  OR2_X1 U3428 ( .A1(n3030), .A2(n3842), .ZN(n2958) );
  NAND2_X1 U3429 ( .A1(n3090), .A2(n3127), .ZN(n2957) );
  NAND2_X1 U3430 ( .A1(n2958), .A2(n2957), .ZN(n2988) );
  XNOR2_X1 U3431 ( .A(n2987), .B(n2988), .ZN(n2964) );
  INV_X1 U3432 ( .A(n2959), .ZN(n2961) );
  NAND2_X1 U3433 ( .A1(n2961), .A2(n2960), .ZN(n2965) );
  AND2_X1 U3434 ( .A1(n2964), .A2(n2965), .ZN(n2962) );
  NAND2_X1 U3435 ( .A1(n2963), .A2(n2962), .ZN(n2991) );
  NAND2_X1 U3436 ( .A1(n2991), .A2(n5274), .ZN(n2979) );
  AOI21_X1 U3437 ( .B1(n2963), .B2(n2965), .A(n2964), .ZN(n2978) );
  NAND2_X1 U3438 ( .A1(n3130), .A2(REG1_REG_5__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U3439 ( .A1(n2940), .A2(REG2_REG_5__SCAN_IN), .ZN(n2971) );
  AND2_X1 U3440 ( .A1(n2967), .A2(n4117), .ZN(n2968) );
  NOR2_X1 U3441 ( .A1(n2995), .A2(n2968), .ZN(n3204) );
  NAND2_X1 U3442 ( .A1(n2937), .A2(n3204), .ZN(n2970) );
  NAND2_X1 U3443 ( .A1(n2941), .A2(REG0_REG_5__SCAN_IN), .ZN(n2969) );
  AOI22_X1 U3444 ( .A1(n4538), .A2(n4358), .B1(n3090), .B2(n5263), .ZN(n2977)
         );
  NOR2_X2 U3445 ( .A1(n4345), .A2(n2763), .ZN(n5265) );
  NOR2_X1 U3446 ( .A1(STATE_REG_SCAN_IN), .A2(n4125), .ZN(n5052) );
  INV_X1 U3447 ( .A(n2974), .ZN(n3056) );
  NOR2_X1 U3448 ( .A1(n5279), .A2(n3056), .ZN(n2975) );
  AOI211_X1 U3449 ( .C1(n5265), .C2(n4540), .A(n5052), .B(n2975), .ZN(n2976)
         );
  OAI211_X1 U3450 ( .C1(n2979), .C2(n2978), .A(n2977), .B(n2976), .ZN(U3227)
         );
  OAI21_X1 U3451 ( .B1(n2981), .B2(n2980), .A(n2963), .ZN(n2985) );
  OAI22_X1 U3452 ( .A1(n5272), .A2(n3030), .B1(n4324), .B2(n3109), .ZN(n2984)
         );
  INV_X1 U3453 ( .A(n3102), .ZN(n3025) );
  NAND2_X1 U3454 ( .A1(n3025), .A2(n5265), .ZN(n2982) );
  NAND2_X1 U3455 ( .A1(U3149), .A2(REG3_REG_3__SCAN_IN), .ZN(n4954) );
  OAI211_X1 U3456 ( .C1(REG3_REG_3__SCAN_IN), .C2(n5279), .A(n2982), .B(n4954), 
        .ZN(n2983) );
  AOI211_X1 U3457 ( .C1(n2985), .C2(n5274), .A(n2984), .B(n2983), .ZN(n2986)
         );
  INV_X1 U34580 ( .A(n2986), .ZN(U3215) );
  INV_X1 U34590 ( .A(n2987), .ZN(n2989) );
  NAND2_X1 U3460 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
  NAND2_X1 U3461 ( .A1(n2991), .A2(n2990), .ZN(n3121) );
  MUX2_X1 U3462 ( .A(n4924), .B(DATAI_5_), .S(n4404), .Z(n3196) );
  OAI22_X1 U3463 ( .A1(n3095), .A2(n3446), .B1(n3200), .B2(n3456), .ZN(n2992)
         );
  XNOR2_X1 U3464 ( .A(n2992), .B(n3824), .ZN(n3117) );
  OR2_X1 U3465 ( .A1(n3095), .A2(n3842), .ZN(n2994) );
  NAND2_X1 U3466 ( .A1(n3196), .A2(n3127), .ZN(n2993) );
  NAND2_X1 U34670 ( .A1(n2994), .A2(n2993), .ZN(n3118) );
  XNOR2_X1 U3468 ( .A(n3117), .B(n3118), .ZN(n3120) );
  XNOR2_X1 U34690 ( .A(n3121), .B(n3120), .ZN(n3006) );
  NAND2_X1 U3470 ( .A1(n3130), .A2(REG1_REG_6__SCAN_IN), .ZN(n3000) );
  NAND2_X1 U34710 ( .A1(n2941), .A2(REG0_REG_6__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3472 ( .A1(n2995), .A2(REG3_REG_6__SCAN_IN), .ZN(n3077) );
  OR2_X1 U34730 ( .A1(n2995), .A2(REG3_REG_6__SCAN_IN), .ZN(n2996) );
  AND2_X1 U3474 ( .A1(n3077), .A2(n2996), .ZN(n3087) );
  NAND2_X1 U34750 ( .A1(n2937), .A2(n3087), .ZN(n2998) );
  NAND2_X1 U3476 ( .A1(n2940), .A2(REG2_REG_6__SCAN_IN), .ZN(n2997) );
  OR2_X1 U34770 ( .A1(n3138), .A2(n5200), .ZN(n3002) );
  OR2_X1 U3478 ( .A1(n3030), .A2(n5154), .ZN(n3001) );
  NAND2_X1 U34790 ( .A1(n3002), .A2(n3001), .ZN(n3195) );
  NAND2_X1 U3480 ( .A1(n3195), .A2(n3798), .ZN(n3003) );
  NAND2_X1 U34810 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4576) );
  OAI211_X1 U3482 ( .C1(n4324), .C2(n3200), .A(n3003), .B(n4576), .ZN(n3004)
         );
  AOI21_X1 U34830 ( .B1(n3204), .B2(n4317), .A(n3004), .ZN(n3005) );
  OAI21_X1 U3484 ( .B1(n3006), .B2(n4363), .A(n3005), .ZN(U3224) );
  INV_X1 U34850 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U3486 ( .A(REG1_REG_11__SCAN_IN), .B(n5161), .S(n3328), .Z(n3009) );
  NOR2_X1 U34870 ( .A1(n3328), .A2(n5161), .ZN(n3008) );
  AOI211_X1 U3488 ( .C1(n3010), .C2(n3009), .A(n5049), .B(n3208), .ZN(n3021)
         );
  NAND2_X1 U34890 ( .A1(n4921), .A2(n3011), .ZN(n3013) );
  NAND2_X1 U3490 ( .A1(n3013), .A2(n3012), .ZN(n3016) );
  INV_X1 U34910 ( .A(REG2_REG_11__SCAN_IN), .ZN(n5172) );
  NOR2_X1 U3492 ( .A1(n3328), .A2(n5172), .ZN(n3014) );
  AOI21_X1 U34930 ( .B1(n5172), .B2(n3328), .A(n3014), .ZN(n3015) );
  NAND2_X1 U3494 ( .A1(n3015), .A2(n3016), .ZN(n3212) );
  OAI211_X1 U34950 ( .C1(n3016), .C2(n3015), .A(n5043), .B(n3212), .ZN(n3019)
         );
  NAND2_X1 U3496 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3343) );
  INV_X1 U34970 ( .A(n3343), .ZN(n3017) );
  AOI21_X1 U3498 ( .B1(n5053), .B2(ADDR_REG_11__SCAN_IN), .A(n3017), .ZN(n3018) );
  OAI211_X1 U34990 ( .C1(n5009), .C2(n3328), .A(n3019), .B(n3018), .ZN(n3020)
         );
  OR2_X1 U3500 ( .A1(n3021), .A2(n3020), .ZN(U3251) );
  AND2_X1 U35010 ( .A1(n3039), .A2(n4384), .ZN(n3063) );
  NAND2_X1 U3502 ( .A1(n3063), .A2(n3038), .ZN(n3062) );
  NAND2_X1 U35030 ( .A1(n3023), .A2(n2838), .ZN(n3024) );
  NAND2_X1 U3504 ( .A1(n3062), .A2(n3024), .ZN(n3154) );
  INV_X1 U35050 ( .A(n3154), .ZN(n3026) );
  NAND2_X1 U35060 ( .A1(n3025), .A2(n3165), .ZN(n4431) );
  NAND2_X1 U35070 ( .A1(n3026), .A2(n3041), .ZN(n3156) );
  NAND2_X1 U35080 ( .A1(n3102), .A2(n3165), .ZN(n3027) );
  NAND2_X1 U35090 ( .A1(n4540), .A2(n3053), .ZN(n3029) );
  NOR2_X1 U35100 ( .A1(n4540), .A2(n3053), .ZN(n3028) );
  NAND2_X1 U35110 ( .A1(n3030), .A2(n3090), .ZN(n4435) );
  NAND2_X1 U35120 ( .A1(n4539), .A2(n3037), .ZN(n3192) );
  NAND2_X1 U35130 ( .A1(n4435), .A2(n3192), .ZN(n3045) );
  NAND2_X1 U35140 ( .A1(n3031), .A2(n3045), .ZN(n3092) );
  OAI21_X1 U35150 ( .B1(n3031), .B2(n3045), .A(n3092), .ZN(n5090) );
  OR2_X1 U35160 ( .A1(n2842), .A2(n4848), .ZN(n3061) );
  INV_X1 U35170 ( .A(n3061), .ZN(n3035) );
  NAND2_X1 U35180 ( .A1(n5173), .A2(n3035), .ZN(n3419) );
  OAI22_X1 U35190 ( .A1(n3159), .A2(n5154), .B1(n3037), .B2(n5293), .ZN(n3051)
         );
  NOR2_X1 U35200 ( .A1(n3039), .A2(n5057), .ZN(n3065) );
  NAND2_X1 U35210 ( .A1(n5058), .A2(n2838), .ZN(n3040) );
  NAND2_X1 U35220 ( .A1(n3064), .A2(n3040), .ZN(n4433) );
  NAND2_X1 U35230 ( .A1(n4433), .A2(n4389), .ZN(n3157) );
  NAND2_X1 U35240 ( .A1(n3157), .A2(n4428), .ZN(n3042) );
  NAND2_X1 U35250 ( .A1(n3159), .A2(n3053), .ZN(n4434) );
  NAND2_X1 U35260 ( .A1(n4540), .A2(n3109), .ZN(n4430) );
  INV_X1 U35270 ( .A(n4434), .ZN(n3043) );
  NOR2_X1 U35280 ( .A1(n3045), .A2(n3043), .ZN(n3044) );
  NAND2_X1 U35290 ( .A1(n3105), .A2(n3044), .ZN(n3193) );
  INV_X1 U35300 ( .A(n3193), .ZN(n3049) );
  INV_X1 U35310 ( .A(n3045), .ZN(n4370) );
  AOI21_X1 U35320 ( .B1(n3105), .B2(n4434), .A(n4370), .ZN(n3048) );
  NAND2_X1 U35330 ( .A1(n4849), .A2(n4916), .ZN(n3047) );
  INV_X1 U35340 ( .A(n4848), .ZN(n5064) );
  NAND2_X1 U35350 ( .A1(n5064), .A2(n4915), .ZN(n3046) );
  NOR3_X1 U35360 ( .A1(n3049), .A2(n3048), .A3(n5206), .ZN(n3050) );
  AOI211_X1 U35370 ( .C1(n4809), .C2(n4538), .A(n3051), .B(n3050), .ZN(n3052)
         );
  OAI21_X1 U35380 ( .B1(n3036), .B2(n5090), .A(n3052), .ZN(n5091) );
  NAND2_X1 U35390 ( .A1(n5091), .A2(n5173), .ZN(n3060) );
  NAND2_X1 U35400 ( .A1(n3166), .A2(n3165), .ZN(n3164) );
  NAND2_X1 U35410 ( .A1(n3108), .A2(n3090), .ZN(n3054) );
  NAND2_X1 U35420 ( .A1(n3054), .A2(n5304), .ZN(n3055) );
  NOR2_X1 U35430 ( .A1(n3201), .A2(n3055), .ZN(n5092) );
  INV_X1 U35440 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3057) );
  OAI22_X1 U35450 ( .A1(n5173), .A2(n3057), .B1(n3056), .B2(n5216), .ZN(n3058)
         );
  AOI21_X1 U35460 ( .B1(n5092), .B2(n4843), .A(n3058), .ZN(n3059) );
  OAI211_X1 U35470 ( .C1(n5090), .C2(n3419), .A(n3060), .B(n3059), .ZN(U3286)
         );
  NAND2_X1 U35480 ( .A1(n3036), .A2(n3061), .ZN(n5165) );
  OAI21_X1 U35490 ( .B1(n4385), .B2(n3065), .A(n3064), .ZN(n3066) );
  NAND2_X1 U35500 ( .A1(n3066), .A2(n5151), .ZN(n3069) );
  INV_X1 U35510 ( .A(n3067), .ZN(n3068) );
  OAI211_X1 U35520 ( .C1(n5293), .C2(n3070), .A(n3069), .B(n3068), .ZN(n5073)
         );
  NAND2_X1 U35530 ( .A1(n5073), .A2(n5173), .ZN(n3075) );
  AOI21_X1 U35540 ( .B1(n4384), .B2(n2838), .A(n3166), .ZN(n5075) );
  INV_X1 U35550 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3072) );
  INV_X1 U35560 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3071) );
  OAI22_X1 U35570 ( .A1(n5173), .A2(n3072), .B1(n3071), .B2(n5216), .ZN(n3073)
         );
  AOI21_X1 U35580 ( .B1(n5300), .B2(n5075), .A(n3073), .ZN(n3074) );
  OAI211_X1 U35590 ( .C1(n4806), .C2(n5072), .A(n3075), .B(n3074), .ZN(U3289)
         );
  INV_X1 U35600 ( .A(n3138), .ZN(n4537) );
  MUX2_X1 U35610 ( .A(n4970), .B(DATAI_6_), .S(n4404), .Z(n3179) );
  INV_X1 U35620 ( .A(n3179), .ZN(n3123) );
  NAND2_X1 U35630 ( .A1(n4537), .A2(n3123), .ZN(n4439) );
  NAND2_X1 U35640 ( .A1(n3138), .A2(n3179), .ZN(n4437) );
  NAND2_X1 U35650 ( .A1(n4538), .A2(n3200), .ZN(n3093) );
  AND2_X1 U35660 ( .A1(n3093), .A2(n3192), .ZN(n4443) );
  NAND2_X1 U35670 ( .A1(n3193), .A2(n4443), .ZN(n3076) );
  NAND2_X1 U35680 ( .A1(n3095), .A2(n3196), .ZN(n4415) );
  NAND2_X1 U35690 ( .A1(n3076), .A2(n4415), .ZN(n3172) );
  XOR2_X1 U35700 ( .A(n2540), .B(n3172), .Z(n3085) );
  NAND2_X1 U35710 ( .A1(n3130), .A2(REG1_REG_7__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U35720 ( .A1(n2940), .A2(REG2_REG_7__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U35730 ( .A1(n3077), .A2(n4093), .ZN(n3078) );
  AND2_X1 U35740 ( .A1(n3131), .A2(n3078), .ZN(n3184) );
  NAND2_X1 U35750 ( .A1(n3612), .A2(n3184), .ZN(n3080) );
  NAND2_X1 U35760 ( .A1(n4375), .A2(REG0_REG_7__SCAN_IN), .ZN(n3079) );
  OAI22_X1 U35770 ( .A1(n3095), .A2(n5154), .B1(n3123), .B2(n5293), .ZN(n3083)
         );
  AOI21_X1 U35780 ( .B1(n4809), .B2(n4536), .A(n3083), .ZN(n3084) );
  OAI21_X1 U35790 ( .B1(n3085), .B2(n5206), .A(n3084), .ZN(n5106) );
  INV_X1 U35800 ( .A(n5106), .ZN(n3101) );
  NAND2_X1 U35810 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  NAND2_X1 U3582 ( .A1(n3202), .A2(n3179), .ZN(n3086) );
  AND2_X1 U3583 ( .A1(n2710), .A2(n3086), .ZN(n5107) );
  INV_X1 U3584 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3088) );
  INV_X1 U3585 ( .A(n3087), .ZN(n3150) );
  OAI22_X1 U3586 ( .A1(n5173), .A2(n3088), .B1(n3150), .B2(n5216), .ZN(n3089)
         );
  AOI21_X1 U3587 ( .B1(n5107), .B2(n5300), .A(n3089), .ZN(n3100) );
  NAND2_X1 U3588 ( .A1(n4539), .A2(n3090), .ZN(n3091) );
  NAND2_X1 U3589 ( .A1(n3095), .A2(n3200), .ZN(n3096) );
  INV_X1 U3590 ( .A(n2540), .ZN(n3097) );
  NAND2_X1 U3591 ( .A1(n3098), .A2(n2540), .ZN(n5104) );
  NAND3_X1 U3592 ( .A1(n3181), .A2(n5104), .A3(n4837), .ZN(n3099) );
  OAI211_X1 U3593 ( .C1(n3101), .C2(n4847), .A(n3100), .B(n3099), .ZN(U3284)
         );
  OAI22_X1 U3594 ( .A1(n3102), .A2(n5154), .B1(n5293), .B2(n3109), .ZN(n3107)
         );
  INV_X1 U3595 ( .A(n4388), .ZN(n3103) );
  NAND3_X1 U3596 ( .A1(n3157), .A2(n4428), .A3(n3103), .ZN(n3104) );
  AOI21_X1 U3597 ( .B1(n3105), .B2(n3104), .A(n5206), .ZN(n3106) );
  AOI211_X1 U3598 ( .C1(n4809), .C2(n4539), .A(n3107), .B(n3106), .ZN(n5084)
         );
  INV_X1 U3599 ( .A(n3164), .ZN(n3110) );
  OAI21_X1 U3600 ( .B1(n3110), .B2(n3109), .A(n3108), .ZN(n5085) );
  INV_X1 U3601 ( .A(n5085), .ZN(n3113) );
  INV_X1 U3602 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3111) );
  OAI22_X1 U3603 ( .A1(n5173), .A2(n3111), .B1(REG3_REG_3__SCAN_IN), .B2(n5216), .ZN(n3112) );
  AOI21_X1 U3604 ( .B1(n3113), .B2(n5300), .A(n3112), .ZN(n3116) );
  XOR2_X1 U3605 ( .A(n3114), .B(n4388), .Z(n5087) );
  NAND2_X1 U3606 ( .A1(n5087), .A2(n4837), .ZN(n3115) );
  OAI211_X1 U3607 ( .C1(n5084), .C2(n4847), .A(n3116), .B(n3115), .ZN(U3287)
         );
  INV_X1 U3608 ( .A(n3117), .ZN(n3119) );
  AOI21_X2 U3609 ( .B1(n3121), .B2(n3120), .A(n2715), .ZN(n3146) );
  OAI22_X1 U3610 ( .A1(n3138), .A2(n3446), .B1(n3123), .B2(n3719), .ZN(n3122)
         );
  XNOR2_X1 U3611 ( .A(n3122), .B(n3843), .ZN(n3125) );
  OAI22_X1 U3612 ( .A1(n3138), .A2(n3842), .B1(n3123), .B2(n3845), .ZN(n3124)
         );
  XNOR2_X1 U3613 ( .A(n3125), .B(n3124), .ZN(n3145) );
  MUX2_X1 U3614 ( .A(n4923), .B(DATAI_7_), .S(n4404), .Z(n3239) );
  INV_X1 U3615 ( .A(n3239), .ZN(n3176) );
  OAI22_X1 U3616 ( .A1(n3174), .A2(n3446), .B1(n3176), .B2(n3719), .ZN(n3126)
         );
  XNOR2_X1 U3617 ( .A(n3126), .B(n3824), .ZN(n3218) );
  OR2_X1 U3618 ( .A1(n3174), .A2(n3842), .ZN(n3129) );
  NAND2_X1 U3619 ( .A1(n3239), .A2(n3127), .ZN(n3128) );
  NAND2_X1 U3620 ( .A1(n3129), .A2(n3128), .ZN(n3219) );
  XNOR2_X1 U3621 ( .A(n3218), .B(n3219), .ZN(n3221) );
  XNOR2_X1 U3622 ( .A(n3222), .B(n3221), .ZN(n3144) );
  NAND2_X1 U3623 ( .A1(n3130), .A2(REG1_REG_8__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3624 ( .A1(n4375), .A2(REG0_REG_8__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3625 ( .A1(n3131), .A2(n3916), .ZN(n3132) );
  NAND2_X1 U3626 ( .A1(n3228), .A2(n3132), .ZN(n3253) );
  INV_X1 U3627 ( .A(n3253), .ZN(n3133) );
  NAND2_X1 U3628 ( .A1(n3612), .A2(n3133), .ZN(n3135) );
  NAND2_X1 U3629 ( .A1(n2940), .A2(REG2_REG_8__SCAN_IN), .ZN(n3134) );
  OR2_X1 U3630 ( .A1(n4314), .A2(n5200), .ZN(n3140) );
  OR2_X1 U3631 ( .A1(n3138), .A2(n5154), .ZN(n3139) );
  AND2_X1 U3632 ( .A1(n3140), .A2(n3139), .ZN(n3175) );
  NAND2_X1 U3633 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U3634 ( .A1(n5263), .A2(n3239), .ZN(n3141) );
  OAI211_X1 U3635 ( .C1(n3175), .C2(n4345), .A(n4586), .B(n3141), .ZN(n3142)
         );
  AOI21_X1 U3636 ( .B1(n3184), .B2(n4317), .A(n3142), .ZN(n3143) );
  OAI21_X1 U3637 ( .B1(n3144), .B2(n4363), .A(n3143), .ZN(U3210) );
  XOR2_X1 U3638 ( .A(n3146), .B(n3145), .Z(n3152) );
  AOI22_X1 U3639 ( .A1(n4536), .A2(n4358), .B1(n3179), .B2(n5263), .ZN(n3149)
         );
  INV_X1 U3640 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3147) );
  NOR2_X1 U3641 ( .A1(STATE_REG_SCAN_IN), .A2(n3147), .ZN(n4965) );
  AOI21_X1 U3642 ( .B1(n4538), .B2(n5265), .A(n4965), .ZN(n3148) );
  OAI211_X1 U3643 ( .C1(n3150), .C2(n5279), .A(n3149), .B(n3148), .ZN(n3151)
         );
  AOI21_X1 U3644 ( .B1(n3152), .B2(n5274), .A(n3151), .ZN(n3153) );
  INV_X1 U3645 ( .A(n3153), .ZN(U3236) );
  NAND2_X1 U3646 ( .A1(n3154), .A2(n4389), .ZN(n3155) );
  AND2_X1 U3647 ( .A1(n3156), .A2(n3155), .ZN(n3163) );
  OAI21_X1 U3648 ( .B1(n4389), .B2(n4433), .A(n3157), .ZN(n3161) );
  AOI22_X1 U3649 ( .A1(n3023), .A2(n5204), .B1(n4335), .B2(n5283), .ZN(n3158)
         );
  OAI21_X1 U3650 ( .B1(n3159), .B2(n5200), .A(n3158), .ZN(n3160) );
  AOI21_X1 U3651 ( .B1(n3161), .B2(n5151), .A(n3160), .ZN(n3162) );
  OAI21_X1 U3652 ( .B1(n3163), .B2(n3036), .A(n3162), .ZN(n5079) );
  INV_X1 U3653 ( .A(n5079), .ZN(n3170) );
  INV_X1 U3654 ( .A(n3163), .ZN(n5081) );
  INV_X1 U3655 ( .A(n3419), .ZN(n5222) );
  INV_X1 U3656 ( .A(n5300), .ZN(n3274) );
  OAI21_X1 U3657 ( .B1(n3166), .B2(n3165), .A(n3164), .ZN(n5078) );
  INV_X1 U3658 ( .A(n5216), .ZN(n5168) );
  AOI22_X1 U3659 ( .A1(n5285), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n5168), .ZN(n3167) );
  OAI21_X1 U3660 ( .B1(n3274), .B2(n5078), .A(n3167), .ZN(n3168) );
  AOI21_X1 U3661 ( .B1(n5081), .B2(n5222), .A(n3168), .ZN(n3169) );
  OAI21_X1 U3662 ( .B1(n3170), .B2(n4847), .A(n3169), .ZN(U3288) );
  INV_X1 U3663 ( .A(n4437), .ZN(n3171) );
  NAND2_X1 U3664 ( .A1(n3174), .A2(n3239), .ZN(n4438) );
  NAND2_X1 U3665 ( .A1(n4536), .A2(n3176), .ZN(n4441) );
  NAND2_X1 U3666 ( .A1(n4438), .A2(n4441), .ZN(n4387) );
  XNOR2_X1 U3667 ( .A(n3245), .B(n4387), .ZN(n3178) );
  OAI21_X1 U3668 ( .B1(n3176), .B2(n5293), .A(n3175), .ZN(n3177) );
  AOI21_X1 U3669 ( .B1(n3178), .B2(n5151), .A(n3177), .ZN(n5114) );
  NAND2_X1 U3670 ( .A1(n4537), .A2(n3179), .ZN(n3180) );
  NAND2_X1 U3671 ( .A1(n3181), .A2(n3180), .ZN(n3182) );
  OAI21_X1 U3672 ( .B1(n3182), .B2(n4387), .A(n3241), .ZN(n5112) );
  INV_X1 U3673 ( .A(n5112), .ZN(n3188) );
  AOI21_X1 U3674 ( .B1(n2710), .B2(n3239), .A(n5229), .ZN(n3183) );
  NAND2_X1 U3675 ( .A1(n3183), .A2(n3251), .ZN(n5113) );
  INV_X1 U3676 ( .A(n4843), .ZN(n4802) );
  NOR2_X1 U3677 ( .A1(n5113), .A2(n4802), .ZN(n3187) );
  INV_X1 U3678 ( .A(n3184), .ZN(n3185) );
  OAI22_X1 U3679 ( .A1(n5173), .A2(n2902), .B1(n3185), .B2(n5216), .ZN(n3186)
         );
  AOI211_X1 U3680 ( .C1(n3188), .C2(n4837), .A(n3187), .B(n3186), .ZN(n3189)
         );
  OAI21_X1 U3681 ( .B1(n4847), .B2(n5114), .A(n3189), .ZN(U3283) );
  OAI21_X1 U3682 ( .B1(n3191), .B2(n3094), .A(n3190), .ZN(n5101) );
  INV_X1 U3683 ( .A(n5101), .ZN(n3207) );
  NAND2_X1 U3684 ( .A1(n3193), .A2(n3192), .ZN(n3194) );
  XNOR2_X1 U3685 ( .A(n4368), .B(n3194), .ZN(n3198) );
  AOI21_X1 U3686 ( .B1(n3196), .B2(n5283), .A(n3195), .ZN(n3197) );
  OAI21_X1 U3687 ( .B1(n3198), .B2(n5206), .A(n3197), .ZN(n5099) );
  INV_X1 U3688 ( .A(n5099), .ZN(n3199) );
  MUX2_X1 U3689 ( .A(n2903), .B(n3199), .S(n5173), .Z(n3206) );
  NOR2_X1 U3690 ( .A1(n3201), .A2(n3200), .ZN(n5098) );
  INV_X1 U3691 ( .A(n3202), .ZN(n5097) );
  NOR3_X1 U3692 ( .A1(n5098), .A2(n5097), .A3(n3274), .ZN(n3203) );
  AOI21_X1 U3693 ( .B1(n5168), .B2(n3204), .A(n3203), .ZN(n3205) );
  OAI211_X1 U3694 ( .C1(n3207), .C2(n4806), .A(n3206), .B(n3205), .ZN(U3285)
         );
  INV_X1 U3695 ( .A(n3328), .ZN(n3209) );
  AOI21_X1 U3696 ( .B1(REG1_REG_11__SCAN_IN), .B2(n3209), .A(n3208), .ZN(n4597) );
  XNOR2_X1 U3697 ( .A(n4598), .B(REG1_REG_12__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U3698 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U3699 ( .A1(n5053), .A2(ADDR_REG_12__SCAN_IN), .ZN(n3210) );
  OAI211_X1 U3700 ( .C1(n5009), .C2(n4596), .A(n3365), .B(n3210), .ZN(n3211)
         );
  INV_X1 U3701 ( .A(n3211), .ZN(n3216) );
  OR2_X1 U3702 ( .A1(n3328), .A2(n5172), .ZN(n3213) );
  OAI211_X1 U3703 ( .C1(REG2_REG_12__SCAN_IN), .C2(n3214), .A(n5043), .B(n4608), .ZN(n3215) );
  OAI211_X1 U3704 ( .C1(n3217), .C2(n5049), .A(n3216), .B(n3215), .ZN(U3252)
         );
  INV_X1 U3705 ( .A(n3218), .ZN(n3220) );
  MUX2_X1 U3706 ( .A(n4978), .B(DATAI_8_), .S(n4404), .Z(n3252) );
  INV_X1 U3707 ( .A(n3252), .ZN(n3271) );
  OAI22_X1 U3708 ( .A1(n4314), .A2(n3446), .B1(n3271), .B2(n3456), .ZN(n3223)
         );
  XNOR2_X1 U3709 ( .A(n3223), .B(n3843), .ZN(n3227) );
  OR2_X1 U3710 ( .A1(n4314), .A2(n3842), .ZN(n3225) );
  NAND2_X1 U3711 ( .A1(n3252), .A2(n3127), .ZN(n3224) );
  NAND2_X1 U3712 ( .A1(n3225), .A2(n3224), .ZN(n3226) );
  NOR2_X1 U3713 ( .A1(n3227), .A2(n3226), .ZN(n3315) );
  AOI21_X1 U3714 ( .B1(n3227), .B2(n3226), .A(n3315), .ZN(n3314) );
  NAND2_X1 U3715 ( .A1(n3318), .A2(n3314), .ZN(n4308) );
  OAI21_X1 U3716 ( .B1(n3318), .B2(n3314), .A(n4308), .ZN(n3237) );
  NAND2_X1 U3717 ( .A1(n2938), .A2(REG1_REG_9__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U3718 ( .A1(n4375), .A2(REG0_REG_9__SCAN_IN), .ZN(n3232) );
  AND2_X1 U3719 ( .A1(n3228), .A2(n4313), .ZN(n3229) );
  NOR2_X1 U3720 ( .A1(n3261), .A2(n3229), .ZN(n4316) );
  NAND2_X1 U3721 ( .A1(n3612), .A2(n4316), .ZN(n3231) );
  NAND2_X1 U3722 ( .A1(n2940), .A2(REG2_REG_9__SCAN_IN), .ZN(n3230) );
  INV_X1 U3723 ( .A(n3312), .ZN(n4534) );
  AOI22_X1 U3724 ( .A1(n4534), .A2(n4358), .B1(n3252), .B2(n5263), .ZN(n3235)
         );
  NOR2_X1 U3725 ( .A1(STATE_REG_SCAN_IN), .A2(n3916), .ZN(n4975) );
  AOI21_X1 U3726 ( .B1(n4536), .B2(n5265), .A(n4975), .ZN(n3234) );
  OAI211_X1 U3727 ( .C1(n3253), .C2(n5279), .A(n3235), .B(n3234), .ZN(n3236)
         );
  AOI21_X1 U3728 ( .B1(n3237), .B2(n5274), .A(n3236), .ZN(n3238) );
  INV_X1 U3729 ( .A(n3238), .ZN(U3218) );
  NAND2_X1 U3730 ( .A1(n4536), .A2(n3239), .ZN(n3240) );
  NAND2_X1 U3731 ( .A1(n4314), .A2(n3252), .ZN(n3284) );
  INV_X1 U3732 ( .A(n4314), .ZN(n4535) );
  NAND2_X1 U3733 ( .A1(n4535), .A2(n3271), .ZN(n4416) );
  NAND2_X1 U3734 ( .A1(n3284), .A2(n4416), .ZN(n3243) );
  OAI21_X1 U3735 ( .B1(n3242), .B2(n3243), .A(n3273), .ZN(n5120) );
  INV_X1 U3736 ( .A(n3036), .ZN(n5209) );
  INV_X1 U3737 ( .A(n3243), .ZN(n4371) );
  INV_X1 U3738 ( .A(n4441), .ZN(n3244) );
  OAI21_X1 U3739 ( .B1(n4371), .B2(n3246), .A(n3259), .ZN(n3247) );
  NAND2_X1 U3740 ( .A1(n3247), .A2(n5151), .ZN(n3249) );
  AOI22_X1 U3741 ( .A1(n4536), .A2(n5204), .B1(n3252), .B2(n5283), .ZN(n3248)
         );
  OAI211_X1 U3742 ( .C1(n3312), .C2(n5200), .A(n3249), .B(n3248), .ZN(n3250)
         );
  AOI21_X1 U3743 ( .B1(n5120), .B2(n5209), .A(n3250), .ZN(n5122) );
  AOI21_X1 U3744 ( .B1(n3252), .B2(n3251), .A(n3275), .ZN(n5119) );
  INV_X1 U3745 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3254) );
  OAI22_X1 U3746 ( .A1(n5173), .A2(n3254), .B1(n3253), .B2(n5216), .ZN(n3255)
         );
  AOI21_X1 U3747 ( .B1(n5119), .B2(n5300), .A(n3255), .ZN(n3257) );
  NAND2_X1 U3748 ( .A1(n5120), .A2(n5222), .ZN(n3256) );
  OAI211_X1 U3749 ( .C1(n5122), .C2(n4847), .A(n3257), .B(n3256), .ZN(U3282)
         );
  NAND2_X1 U3750 ( .A1(n3259), .A2(n3284), .ZN(n3258) );
  MUX2_X1 U3751 ( .A(n4922), .B(DATAI_9_), .S(n4404), .Z(n4312) );
  NAND2_X1 U3752 ( .A1(n3312), .A2(n4312), .ZN(n3283) );
  NAND2_X1 U3753 ( .A1(n4534), .A2(n3311), .ZN(n4417) );
  NAND2_X1 U3754 ( .A1(n3283), .A2(n4417), .ZN(n3298) );
  INV_X1 U3755 ( .A(n3298), .ZN(n4367) );
  NAND2_X1 U3756 ( .A1(n3258), .A2(n4367), .ZN(n3286) );
  NAND3_X1 U3757 ( .A1(n3259), .A2(n3298), .A3(n3284), .ZN(n3260) );
  AOI21_X1 U3758 ( .B1(n3286), .B2(n3260), .A(n5206), .ZN(n3270) );
  NAND2_X1 U3759 ( .A1(n2938), .A2(REG1_REG_10__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U3760 ( .A1(n4375), .A2(REG0_REG_10__SCAN_IN), .ZN(n3266) );
  NOR2_X1 U3761 ( .A1(n3261), .A2(REG3_REG_10__SCAN_IN), .ZN(n3262) );
  OR2_X1 U3762 ( .A1(n3287), .A2(n3262), .ZN(n3801) );
  INV_X1 U3763 ( .A(n3801), .ZN(n3263) );
  NAND2_X1 U3764 ( .A1(n2937), .A2(n3263), .ZN(n3265) );
  NAND2_X1 U3765 ( .A1(n2940), .A2(REG2_REG_10__SCAN_IN), .ZN(n3264) );
  NOR2_X1 U3766 ( .A1(n5155), .A2(n5200), .ZN(n3269) );
  OAI22_X1 U3767 ( .A1(n4314), .A2(n5154), .B1(n3311), .B2(n5293), .ZN(n3268)
         );
  INV_X1 U3768 ( .A(n5128), .ZN(n3282) );
  NAND2_X1 U3769 ( .A1(n4314), .A2(n3271), .ZN(n3272) );
  XNOR2_X1 U3770 ( .A(n3299), .B(n3298), .ZN(n5130) );
  NAND2_X1 U3771 ( .A1(n5130), .A2(n4837), .ZN(n3281) );
  NOR2_X1 U3772 ( .A1(n3275), .A2(n3311), .ZN(n5127) );
  NOR2_X1 U3773 ( .A1(n5127), .A2(n3274), .ZN(n3279) );
  INV_X1 U3774 ( .A(n4316), .ZN(n3276) );
  OAI22_X1 U3775 ( .A1(n5173), .A2(n3277), .B1(n3276), .B2(n5216), .ZN(n3278)
         );
  AOI21_X1 U3776 ( .B1(n3279), .B2(n5125), .A(n3278), .ZN(n3280) );
  OAI211_X1 U3777 ( .C1(n4847), .C2(n3282), .A(n3281), .B(n3280), .ZN(U3281)
         );
  MUX2_X1 U3778 ( .A(n4921), .B(DATAI_10_), .S(n4404), .Z(n3382) );
  NAND2_X1 U3779 ( .A1(n5155), .A2(n3382), .ZN(n4419) );
  INV_X1 U3780 ( .A(n3382), .ZN(n3794) );
  NAND2_X1 U3781 ( .A1(n4533), .A2(n3794), .ZN(n3470) );
  NAND2_X1 U3782 ( .A1(n3284), .A2(n3283), .ZN(n3285) );
  NAND2_X1 U3783 ( .A1(n3285), .A2(n4417), .ZN(n4445) );
  NAND2_X1 U3784 ( .A1(n3286), .A2(n4445), .ZN(n3394) );
  XOR2_X1 U3785 ( .A(n4366), .B(n3394), .Z(n3294) );
  NAND2_X1 U3786 ( .A1(n4375), .A2(REG0_REG_11__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U3787 ( .A1(n3130), .A2(REG1_REG_11__SCAN_IN), .ZN(n3291) );
  OR2_X1 U3788 ( .A1(n3287), .A2(REG3_REG_11__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U3789 ( .A1(n3288), .A2(n3338), .ZN(n3345) );
  INV_X1 U3790 ( .A(n3345), .ZN(n5169) );
  NAND2_X1 U3791 ( .A1(n3612), .A2(n5169), .ZN(n3290) );
  NAND2_X1 U3792 ( .A1(n2940), .A2(REG2_REG_11__SCAN_IN), .ZN(n3289) );
  NAND4_X1 U3793 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n4532)
         );
  INV_X1 U3794 ( .A(n4532), .ZN(n3369) );
  OAI22_X1 U3795 ( .A1(n3369), .A2(n5200), .B1(n3312), .B2(n5154), .ZN(n3797)
         );
  AOI21_X1 U3796 ( .B1(n3382), .B2(n5283), .A(n3797), .ZN(n3293) );
  OAI21_X1 U3797 ( .B1(n3294), .B2(n5206), .A(n3293), .ZN(n5135) );
  INV_X1 U3798 ( .A(n5135), .ZN(n3304) );
  NAND2_X1 U3799 ( .A1(n5125), .A2(n3382), .ZN(n3295) );
  AND2_X1 U3800 ( .A1(n5145), .A2(n3295), .ZN(n5136) );
  INV_X1 U3801 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3296) );
  OAI22_X1 U3802 ( .A1(n5173), .A2(n3296), .B1(n3801), .B2(n5216), .ZN(n3297)
         );
  AOI21_X1 U3803 ( .B1(n5136), .B2(n5300), .A(n3297), .ZN(n3303) );
  NAND2_X1 U3804 ( .A1(n3312), .A2(n3311), .ZN(n3300) );
  OR2_X1 U3805 ( .A1(n3372), .A2(n4366), .ZN(n5142) );
  NAND2_X1 U3806 ( .A1(n3372), .A2(n4366), .ZN(n5133) );
  NAND3_X1 U3807 ( .A1(n5142), .A2(n5133), .A3(n4837), .ZN(n3302) );
  OAI211_X1 U3808 ( .C1(n3304), .C2(n4847), .A(n3303), .B(n3302), .ZN(U3280)
         );
  OR2_X1 U3809 ( .A1(n5155), .A2(n3842), .ZN(n3306) );
  NAND2_X1 U3810 ( .A1(n3382), .A2(n3127), .ZN(n3305) );
  NAND2_X1 U3811 ( .A1(n3306), .A2(n3305), .ZN(n3323) );
  INV_X1 U3812 ( .A(n3323), .ZN(n3326) );
  OAI22_X1 U3813 ( .A1(n5155), .A2(n3446), .B1(n3794), .B2(n3719), .ZN(n3307)
         );
  XNOR2_X1 U3814 ( .A(n3307), .B(n3824), .ZN(n3325) );
  OR2_X1 U3815 ( .A1(n3312), .A2(n3842), .ZN(n3309) );
  NAND2_X1 U3816 ( .A1(n4312), .A2(n3127), .ZN(n3308) );
  NAND2_X1 U3817 ( .A1(n3309), .A2(n3308), .ZN(n3320) );
  OAI22_X1 U3818 ( .A1(n3312), .A2(n3845), .B1(n3311), .B2(n3719), .ZN(n3313)
         );
  XNOR2_X1 U3819 ( .A(n3313), .B(n3843), .ZN(n3319) );
  XOR2_X1 U3820 ( .A(n3320), .B(n3319), .Z(n4310) );
  AND2_X1 U3821 ( .A1(n3314), .A2(n4310), .ZN(n3317) );
  INV_X1 U3822 ( .A(n4310), .ZN(n3316) );
  INV_X1 U3823 ( .A(n3315), .ZN(n4307) );
  INV_X1 U3824 ( .A(n3319), .ZN(n3322) );
  INV_X1 U3825 ( .A(n3320), .ZN(n3321) );
  NAND2_X1 U3826 ( .A1(n3322), .A2(n3321), .ZN(n3790) );
  XNOR2_X1 U3827 ( .A(n3325), .B(n3323), .ZN(n3792) );
  NAND2_X1 U3828 ( .A1(n4532), .A2(n3127), .ZN(n3330) );
  MUX2_X1 U3829 ( .A(n3328), .B(n3327), .S(n4404), .Z(n5153) );
  OR2_X1 U3830 ( .A1(n5153), .A2(n3719), .ZN(n3329) );
  NAND2_X1 U3831 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  XNOR2_X1 U3832 ( .A(n3331), .B(n3824), .ZN(n3334) );
  NOR2_X1 U3833 ( .A1(n5153), .A2(n3845), .ZN(n3332) );
  AOI21_X1 U3834 ( .B1(n4532), .B2(n3828), .A(n3332), .ZN(n3333) );
  NOR2_X1 U3835 ( .A1(n3334), .A2(n3333), .ZN(n3351) );
  INV_X1 U3836 ( .A(n3351), .ZN(n3335) );
  NAND2_X1 U3837 ( .A1(n3334), .A2(n3333), .ZN(n3350) );
  NAND2_X1 U3838 ( .A1(n3335), .A2(n3350), .ZN(n3336) );
  XNOR2_X1 U3839 ( .A(n3352), .B(n3336), .ZN(n3348) );
  AOI21_X1 U3840 ( .B1(n3338), .B2(n3337), .A(n3356), .ZN(n3482) );
  NAND2_X1 U3841 ( .A1(n3612), .A2(n3482), .ZN(n3342) );
  NAND2_X1 U3842 ( .A1(n3130), .A2(REG1_REG_12__SCAN_IN), .ZN(n3341) );
  NAND2_X1 U3843 ( .A1(n2940), .A2(REG2_REG_12__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U3844 ( .A1(n4375), .A2(REG0_REG_12__SCAN_IN), .ZN(n3339) );
  NAND4_X1 U3845 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n5203)
         );
  INV_X1 U3846 ( .A(n5203), .ZN(n5159) );
  OAI22_X1 U3847 ( .A1(n5272), .A2(n5159), .B1(n4324), .B2(n5153), .ZN(n3347)
         );
  NAND2_X1 U3848 ( .A1(n4533), .A2(n5265), .ZN(n3344) );
  OAI211_X1 U3849 ( .C1(n5279), .C2(n3345), .A(n3344), .B(n3343), .ZN(n3346)
         );
  AOI211_X1 U3850 ( .C1(n3348), .C2(n5274), .A(n3347), .B(n3346), .ZN(n3349)
         );
  INV_X1 U3851 ( .A(n3349), .ZN(U3233) );
  MUX2_X1 U3852 ( .A(n4596), .B(n4073), .S(n4404), .Z(n3479) );
  OAI22_X1 U3853 ( .A1(n5159), .A2(n3842), .B1(n3479), .B2(n3845), .ZN(n3440)
         );
  NAND2_X1 U3854 ( .A1(n5203), .A2(n3127), .ZN(n3354) );
  OR2_X1 U3855 ( .A1(n3479), .A2(n3456), .ZN(n3353) );
  NAND2_X1 U3856 ( .A1(n3354), .A2(n3353), .ZN(n3355) );
  XNOR2_X1 U3857 ( .A(n3355), .B(n3843), .ZN(n3441) );
  XOR2_X1 U3858 ( .A(n3440), .B(n3441), .Z(n3444) );
  XOR2_X1 U3859 ( .A(n3445), .B(n3444), .Z(n3368) );
  OAI21_X1 U3860 ( .B1(n3356), .B2(REG3_REG_13__SCAN_IN), .A(n3373), .ZN(n5217) );
  INV_X1 U3861 ( .A(n5217), .ZN(n3357) );
  NAND2_X1 U3862 ( .A1(n3612), .A2(n3357), .ZN(n3361) );
  NAND2_X1 U3863 ( .A1(n3130), .A2(REG1_REG_13__SCAN_IN), .ZN(n3360) );
  NAND2_X1 U3864 ( .A1(n2940), .A2(REG2_REG_13__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U3865 ( .A1(n4375), .A2(REG0_REG_13__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U3866 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n4531)
         );
  NAND2_X1 U3867 ( .A1(n4531), .A2(n4809), .ZN(n3363) );
  NAND2_X1 U3868 ( .A1(n4532), .A2(n5204), .ZN(n3362) );
  AND2_X1 U3869 ( .A1(n3363), .A2(n3362), .ZN(n3478) );
  NAND2_X1 U3870 ( .A1(n5263), .A2(n2633), .ZN(n3364) );
  OAI211_X1 U3871 ( .C1(n3478), .C2(n4345), .A(n3365), .B(n3364), .ZN(n3366)
         );
  AOI21_X1 U3872 ( .B1(n3482), .B2(n4317), .A(n3366), .ZN(n3367) );
  OAI21_X1 U3873 ( .B1(n3368), .B2(n4363), .A(n3367), .ZN(U3221) );
  NAND2_X1 U3874 ( .A1(n3369), .A2(n5153), .ZN(n3381) );
  INV_X1 U3875 ( .A(n3381), .ZN(n3383) );
  OR2_X1 U3876 ( .A1(n4366), .A2(n3383), .ZN(n3465) );
  AND2_X1 U3877 ( .A1(n5159), .A2(n3479), .ZN(n3385) );
  OR2_X1 U3878 ( .A1(n3465), .A2(n3385), .ZN(n5190) );
  NAND2_X1 U3879 ( .A1(n2741), .A2(IR_REG_31__SCAN_IN), .ZN(n3370) );
  XNOR2_X1 U3880 ( .A(n3370), .B(IR_REG_13__SCAN_IN), .ZN(n4998) );
  MUX2_X1 U3881 ( .A(n4998), .B(DATAI_13_), .S(n4404), .Z(n5182) );
  NOR2_X1 U3882 ( .A1(n4531), .A2(n5182), .ZN(n3386) );
  OR2_X1 U3883 ( .A1(n5190), .A2(n3386), .ZN(n3371) );
  NAND2_X1 U3884 ( .A1(n3130), .A2(REG1_REG_14__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U3885 ( .A1(n2940), .A2(REG2_REG_14__SCAN_IN), .ZN(n3377) );
  AND2_X1 U3886 ( .A1(n3373), .A2(n3905), .ZN(n3374) );
  NOR2_X1 U3887 ( .A1(n3403), .A2(n3374), .ZN(n3414) );
  NAND2_X1 U3888 ( .A1(n2937), .A2(n3414), .ZN(n3376) );
  NAND2_X1 U3889 ( .A1(n4375), .A2(REG0_REG_14__SCAN_IN), .ZN(n3375) );
  XNOR2_X1 U3890 ( .A(n3379), .B(IR_REG_14__SCAN_IN), .ZN(n5016) );
  MUX2_X1 U3891 ( .A(n5016), .B(DATAI_14_), .S(n4404), .Z(n3453) );
  NAND2_X1 U3892 ( .A1(n5201), .A2(n3453), .ZN(n4422) );
  INV_X1 U3893 ( .A(n5201), .ZN(n4530) );
  INV_X1 U3894 ( .A(n3453), .ZN(n3458) );
  NAND2_X1 U3895 ( .A1(n4530), .A2(n3458), .ZN(n4449) );
  INV_X1 U3896 ( .A(n4369), .ZN(n3389) );
  XNOR2_X1 U3897 ( .A(n5203), .B(n3479), .ZN(n4398) );
  NAND2_X1 U3898 ( .A1(n4532), .A2(n3413), .ZN(n3380) );
  NAND2_X1 U3899 ( .A1(n4533), .A2(n3382), .ZN(n5140) );
  AND2_X1 U3900 ( .A1(n5149), .A2(n5140), .ZN(n5141) );
  AND2_X1 U3901 ( .A1(n4398), .A2(n3466), .ZN(n3384) );
  OR2_X1 U3902 ( .A1(n3386), .A2(n5191), .ZN(n3388) );
  NAND2_X1 U3903 ( .A1(n4531), .A2(n5182), .ZN(n3387) );
  NAND2_X1 U3904 ( .A1(n2542), .A2(n3390), .ZN(n3391) );
  AND2_X1 U3905 ( .A1(n3391), .A2(n4369), .ZN(n3392) );
  NOR2_X1 U3906 ( .A1(n3433), .A2(n3392), .ZN(n5231) );
  INV_X1 U3907 ( .A(n4419), .ZN(n3393) );
  NAND2_X1 U3908 ( .A1(n4532), .A2(n5153), .ZN(n3474) );
  AND2_X1 U3909 ( .A1(n3474), .A2(n3470), .ZN(n3397) );
  NAND2_X1 U3910 ( .A1(n4531), .A2(n5199), .ZN(n3396) );
  NAND2_X1 U3911 ( .A1(n5203), .A2(n3479), .ZN(n3395) );
  AND2_X1 U3912 ( .A1(n3396), .A2(n3395), .ZN(n3400) );
  NAND2_X1 U3913 ( .A1(n3471), .A2(n4450), .ZN(n3402) );
  NOR2_X1 U3914 ( .A1(n5203), .A2(n3479), .ZN(n5196) );
  NOR2_X1 U3915 ( .A1(n4532), .A2(n5153), .ZN(n3398) );
  OR2_X1 U3916 ( .A1(n5196), .A2(n3398), .ZN(n3401) );
  NOR2_X1 U3917 ( .A1(n4531), .A2(n5199), .ZN(n3399) );
  AOI21_X1 U3918 ( .B1(n3401), .B2(n3400), .A(n3399), .ZN(n4423) );
  NAND2_X1 U3919 ( .A1(n3402), .A2(n4423), .ZN(n4482) );
  OAI21_X1 U3920 ( .B1(n4369), .B2(n4482), .A(n3491), .ZN(n3411) );
  NAND2_X1 U3921 ( .A1(n4375), .A2(REG0_REG_15__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U3922 ( .A1(n3130), .A2(REG1_REG_15__SCAN_IN), .ZN(n3407) );
  OR2_X1 U3923 ( .A1(n3403), .A2(REG3_REG_15__SCAN_IN), .ZN(n3404) );
  AND2_X1 U3924 ( .A1(n3425), .A2(n3404), .ZN(n3435) );
  NAND2_X1 U3925 ( .A1(n3612), .A2(n3435), .ZN(n3406) );
  NAND2_X1 U3926 ( .A1(n2940), .A2(REG2_REG_15__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U3927 ( .A1(n4531), .A2(n5204), .B1(n3453), .B2(n5283), .ZN(n3409)
         );
  OAI21_X1 U3928 ( .B1(n3523), .B2(n5200), .A(n3409), .ZN(n3410) );
  AOI21_X1 U3929 ( .B1(n3411), .B2(n5151), .A(n3410), .ZN(n3412) );
  OAI21_X1 U3930 ( .B1(n5231), .B2(n3036), .A(n3412), .ZN(n5233) );
  NAND2_X1 U3931 ( .A1(n5233), .A2(n5173), .ZN(n3418) );
  AOI21_X1 U3932 ( .B1(n3453), .B2(n2521), .A(n2634), .ZN(n5227) );
  INV_X1 U3933 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3415) );
  INV_X1 U3934 ( .A(n3414), .ZN(n3460) );
  OAI22_X1 U3935 ( .A1(n5173), .A2(n3415), .B1(n3460), .B2(n5216), .ZN(n3416)
         );
  AOI21_X1 U3936 ( .B1(n5227), .B2(n5300), .A(n3416), .ZN(n3417) );
  OAI211_X1 U3937 ( .C1(n5231), .C2(n3419), .A(n3418), .B(n3417), .ZN(U3276)
         );
  INV_X1 U3938 ( .A(n5173), .ZN(n4847) );
  NAND2_X1 U3939 ( .A1(n3491), .A2(n4422), .ZN(n3424) );
  NAND2_X1 U3940 ( .A1(n3420), .A2(IR_REG_31__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U3941 ( .A1(n3422), .A2(n3421), .ZN(n3493) );
  OR2_X1 U3942 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  MUX2_X1 U3943 ( .A(n4920), .B(DATAI_15_), .S(n4404), .Z(n3524) );
  NAND2_X1 U3944 ( .A1(n3523), .A2(n3524), .ZN(n4421) );
  INV_X1 U3945 ( .A(n3523), .ZN(n4529) );
  INV_X1 U3946 ( .A(n3524), .ZN(n3528) );
  NAND2_X1 U3947 ( .A1(n4529), .A2(n3528), .ZN(n4448) );
  NAND2_X1 U3948 ( .A1(n4421), .A2(n4448), .ZN(n3489) );
  XNOR2_X1 U3949 ( .A(n3424), .B(n3489), .ZN(n3432) );
  NAND2_X1 U3950 ( .A1(n4375), .A2(REG0_REG_16__SCAN_IN), .ZN(n3429) );
  NAND2_X1 U3951 ( .A1(n3130), .A2(REG1_REG_16__SCAN_IN), .ZN(n3428) );
  AOI21_X1 U3952 ( .B1(n3425), .B2(n4116), .A(n3495), .ZN(n3510) );
  NAND2_X1 U3953 ( .A1(n3612), .A2(n3510), .ZN(n3427) );
  NAND2_X1 U3954 ( .A1(n2940), .A2(REG2_REG_16__SCAN_IN), .ZN(n3426) );
  OAI22_X1 U3955 ( .A1(n5201), .A2(n5154), .B1(n3528), .B2(n5293), .ZN(n3430)
         );
  AOI21_X1 U3956 ( .B1(n4809), .B2(n4528), .A(n3430), .ZN(n3431) );
  OAI21_X1 U3957 ( .B1(n3432), .B2(n5206), .A(n3431), .ZN(n5237) );
  INV_X1 U3958 ( .A(n5237), .ZN(n3439) );
  INV_X1 U3959 ( .A(n3489), .ZN(n4391) );
  XNOR2_X1 U3960 ( .A(n3504), .B(n4391), .ZN(n5239) );
  NAND2_X1 U3961 ( .A1(n5239), .A2(n4837), .ZN(n3438) );
  AOI211_X1 U3962 ( .C1(n3524), .C2(n3434), .A(n5229), .B(n3508), .ZN(n5238)
         );
  INV_X1 U3963 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4611) );
  INV_X1 U3964 ( .A(n3435), .ZN(n3530) );
  OAI22_X1 U3965 ( .A1(n5173), .A2(n4611), .B1(n3530), .B2(n5216), .ZN(n3436)
         );
  AOI21_X1 U3966 ( .B1(n5238), .B2(n4843), .A(n3436), .ZN(n3437) );
  OAI211_X1 U3967 ( .C1(n4847), .C2(n3439), .A(n3438), .B(n3437), .ZN(U3275)
         );
  INV_X1 U3968 ( .A(n3440), .ZN(n3443) );
  INV_X1 U3969 ( .A(n3441), .ZN(n3442) );
  AOI22_X1 U3970 ( .A1(n4531), .A2(n3828), .B1(n5182), .B2(n3127), .ZN(n3450)
         );
  NAND2_X1 U3971 ( .A1(n4531), .A2(n3127), .ZN(n3448) );
  NAND2_X1 U3972 ( .A1(n5182), .A2(n2837), .ZN(n3447) );
  NAND2_X1 U3973 ( .A1(n3448), .A2(n3447), .ZN(n3449) );
  XNOR2_X1 U3974 ( .A(n3449), .B(n3843), .ZN(n3452) );
  XOR2_X1 U3975 ( .A(n3450), .B(n3452), .Z(n5183) );
  INV_X1 U3976 ( .A(n3450), .ZN(n3451) );
  OR2_X1 U3977 ( .A1(n5201), .A2(n3842), .ZN(n3455) );
  NAND2_X1 U3978 ( .A1(n3453), .A2(n3127), .ZN(n3454) );
  NAND2_X1 U3979 ( .A1(n3455), .A2(n3454), .ZN(n3517) );
  OAI22_X1 U3980 ( .A1(n5201), .A2(n3845), .B1(n3458), .B2(n3719), .ZN(n3457)
         );
  XNOR2_X1 U3981 ( .A(n3457), .B(n3843), .ZN(n3516) );
  XOR2_X1 U3982 ( .A(n3517), .B(n3516), .Z(n3520) );
  XNOR2_X1 U3983 ( .A(n3521), .B(n3520), .ZN(n3463) );
  OAI22_X1 U3984 ( .A1(n5272), .A2(n3523), .B1(n4324), .B2(n3458), .ZN(n3462)
         );
  NAND2_X1 U3985 ( .A1(n5265), .A2(n4531), .ZN(n3459) );
  NAND2_X1 U3986 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n5012) );
  OAI211_X1 U3987 ( .C1(n5279), .C2(n3460), .A(n3459), .B(n5012), .ZN(n3461)
         );
  AOI211_X1 U3988 ( .C1(n3463), .C2(n5274), .A(n3462), .B(n3461), .ZN(n3464)
         );
  INV_X1 U3989 ( .A(n3464), .ZN(U3212) );
  OR2_X1 U3990 ( .A1(n3372), .A2(n3465), .ZN(n3467) );
  AND2_X1 U3991 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  XNOR2_X1 U3992 ( .A(n3468), .B(n4398), .ZN(n5178) );
  INV_X1 U3993 ( .A(n5178), .ZN(n3487) );
  INV_X1 U3994 ( .A(n5194), .ZN(n3469) );
  OAI21_X1 U3995 ( .B1(n5146), .B2(n3479), .A(n3469), .ZN(n5176) );
  INV_X1 U3996 ( .A(n5176), .ZN(n3485) );
  INV_X1 U3997 ( .A(n5149), .ZN(n3472) );
  NAND2_X1 U3998 ( .A1(n3471), .A2(n3470), .ZN(n5150) );
  NAND2_X1 U3999 ( .A1(n3472), .A2(n5150), .ZN(n3473) );
  NAND2_X1 U4000 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  NAND2_X1 U4001 ( .A1(n4398), .A2(n3475), .ZN(n3477) );
  NOR2_X1 U4002 ( .A1(n4398), .A2(n3475), .ZN(n5195) );
  INV_X1 U4003 ( .A(n5195), .ZN(n3476) );
  NAND2_X1 U4004 ( .A1(n3477), .A2(n3476), .ZN(n3481) );
  OAI21_X1 U4005 ( .B1(n3479), .B2(n5293), .A(n3478), .ZN(n3480) );
  AOI21_X1 U4006 ( .B1(n3481), .B2(n5151), .A(n3480), .ZN(n5175) );
  AOI22_X1 U4007 ( .A1(n5285), .A2(REG2_REG_12__SCAN_IN), .B1(n3482), .B2(
        n5168), .ZN(n3483) );
  OAI21_X1 U4008 ( .B1(n5175), .B2(n4847), .A(n3483), .ZN(n3484) );
  AOI21_X1 U4009 ( .B1(n3485), .B2(n5300), .A(n3484), .ZN(n3486) );
  OAI21_X1 U4010 ( .B1(n3487), .B2(n4806), .A(n3486), .ZN(U3278) );
  INV_X1 U4011 ( .A(n4422), .ZN(n3488) );
  NOR2_X1 U4012 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND2_X1 U4013 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  NAND2_X1 U4014 ( .A1(n3492), .A2(n4448), .ZN(n3541) );
  NAND2_X1 U4015 ( .A1(n3493), .A2(IR_REG_31__SCAN_IN), .ZN(n3494) );
  XNOR2_X1 U4016 ( .A(n3494), .B(IR_REG_16__SCAN_IN), .ZN(n4919) );
  MUX2_X1 U4017 ( .A(n4919), .B(DATAI_16_), .S(n4404), .Z(n3582) );
  NAND2_X1 U4018 ( .A1(n3564), .A2(n3582), .ZN(n4485) );
  NAND2_X1 U4019 ( .A1(n4528), .A2(n3562), .ZN(n3689) );
  NAND2_X1 U4020 ( .A1(n4485), .A2(n3689), .ZN(n3553) );
  INV_X1 U4021 ( .A(n3553), .ZN(n4392) );
  XNOR2_X1 U4022 ( .A(n3541), .B(n4392), .ZN(n3502) );
  NAND2_X1 U4023 ( .A1(n3130), .A2(REG1_REG_17__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U4024 ( .A1(n2940), .A2(REG2_REG_17__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U4025 ( .A1(n4375), .A2(REG0_REG_17__SCAN_IN), .ZN(n3498) );
  NAND2_X1 U4026 ( .A1(n3495), .A2(REG3_REG_17__SCAN_IN), .ZN(n3545) );
  OAI21_X1 U4027 ( .B1(n3495), .B2(REG3_REG_17__SCAN_IN), .A(n3545), .ZN(n4295) );
  INV_X1 U4028 ( .A(n4295), .ZN(n3496) );
  NAND2_X1 U4029 ( .A1(n3612), .A2(n3496), .ZN(n3497) );
  NAND4_X1 U4030 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n4527)
         );
  INV_X1 U4031 ( .A(n4527), .ZN(n3692) );
  OAI22_X1 U4032 ( .A1(n3692), .A2(n5200), .B1(n3523), .B2(n5154), .ZN(n3578)
         );
  AOI21_X1 U4033 ( .B1(n3582), .B2(n5283), .A(n3578), .ZN(n3501) );
  OAI21_X1 U4034 ( .B1(n3502), .B2(n5206), .A(n3501), .ZN(n5243) );
  INV_X1 U4035 ( .A(n5243), .ZN(n3515) );
  NAND2_X1 U4036 ( .A1(n3504), .A2(n4529), .ZN(n3503) );
  NAND2_X1 U4037 ( .A1(n3503), .A2(n3528), .ZN(n3507) );
  NAND2_X1 U4038 ( .A1(n3505), .A2(n3523), .ZN(n3506) );
  XNOR2_X1 U4039 ( .A(n3554), .B(n3553), .ZN(n5245) );
  NAND2_X1 U4040 ( .A1(n5245), .A2(n4837), .ZN(n3514) );
  OAI21_X1 U4041 ( .B1(n3508), .B2(n3562), .A(n5304), .ZN(n3509) );
  NOR2_X1 U4042 ( .A1(n3509), .A2(n3555), .ZN(n5244) );
  INV_X1 U40430 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3511) );
  INV_X1 U4044 ( .A(n3510), .ZN(n3585) );
  OAI22_X1 U4045 ( .A1(n5173), .A2(n3511), .B1(n3585), .B2(n5216), .ZN(n3512)
         );
  AOI21_X1 U4046 ( .B1(n5244), .B2(n4843), .A(n3512), .ZN(n3513) );
  OAI211_X1 U4047 ( .C1(n4847), .C2(n3515), .A(n3514), .B(n3513), .ZN(U3274)
         );
  INV_X1 U4048 ( .A(n3516), .ZN(n3519) );
  INV_X1 U4049 ( .A(n3517), .ZN(n3518) );
  OAI22_X1 U4050 ( .A1(n3523), .A2(n3845), .B1(n3528), .B2(n3719), .ZN(n3522)
         );
  XNOR2_X1 U4051 ( .A(n3522), .B(n3824), .ZN(n3569) );
  OR2_X1 U4052 ( .A1(n3523), .A2(n3842), .ZN(n3526) );
  NAND2_X1 U4053 ( .A1(n3524), .A2(n3127), .ZN(n3525) );
  XNOR2_X1 U4054 ( .A(n3569), .B(n3570), .ZN(n3527) );
  XNOR2_X1 U4055 ( .A(n3574), .B(n3527), .ZN(n3533) );
  OAI22_X1 U4056 ( .A1(n5272), .A2(n3564), .B1(n4324), .B2(n3528), .ZN(n3532)
         );
  NAND2_X1 U4057 ( .A1(n4530), .A2(n5265), .ZN(n3529) );
  NAND2_X1 U4058 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4615) );
  OAI211_X1 U4059 ( .C1(n5279), .C2(n3530), .A(n3529), .B(n4615), .ZN(n3531)
         );
  AOI211_X1 U4060 ( .C1(n3533), .C2(n5274), .A(n3532), .B(n3531), .ZN(n3534)
         );
  INV_X1 U4061 ( .A(n3534), .ZN(U3238) );
  OR2_X1 U4062 ( .A1(n3536), .A2(n4908), .ZN(n3538) );
  MUX2_X1 U4063 ( .A(n3538), .B(IR_REG_31__SCAN_IN), .S(n3537), .Z(n3539) );
  AND2_X1 U4064 ( .A1(n3535), .A2(n3539), .ZN(n4918) );
  INV_X1 U4065 ( .A(DATAI_17_), .ZN(n3540) );
  MUX2_X1 U4066 ( .A(n5039), .B(n3540), .S(n4404), .Z(n3723) );
  NAND2_X1 U4067 ( .A1(n3541), .A2(n4392), .ZN(n3691) );
  INV_X1 U4068 ( .A(n3723), .ZN(n4292) );
  AND2_X1 U4069 ( .A1(n4527), .A2(n4292), .ZN(n3586) );
  INV_X1 U4070 ( .A(n3586), .ZN(n3542) );
  NAND2_X1 U4071 ( .A1(n3692), .A2(n3723), .ZN(n3587) );
  NAND2_X1 U4072 ( .A1(n3542), .A2(n3587), .ZN(n4365) );
  NAND3_X1 U4073 ( .A1(n3691), .A2(n3689), .A3(n4365), .ZN(n4827) );
  INV_X1 U4074 ( .A(n4827), .ZN(n3544) );
  AOI21_X1 U4075 ( .B1(n3691), .B2(n3689), .A(n4365), .ZN(n3543) );
  OAI21_X1 U4076 ( .B1(n3544), .B2(n3543), .A(n5151), .ZN(n3552) );
  NAND2_X1 U4077 ( .A1(n3130), .A2(REG1_REG_18__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4078 ( .A1(n2940), .A2(REG2_REG_18__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4079 ( .A1(n4375), .A2(REG0_REG_18__SCAN_IN), .ZN(n3549) );
  OAI21_X1 U4080 ( .B1(n3546), .B2(REG3_REG_18__SCAN_IN), .A(n3593), .ZN(n4840) );
  INV_X1 U4081 ( .A(n4840), .ZN(n3547) );
  NAND2_X1 U4082 ( .A1(n3612), .A2(n3547), .ZN(n3548) );
  NAND4_X1 U4083 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n4811)
         );
  AOI22_X1 U4084 ( .A1(n4528), .A2(n5204), .B1(n4809), .B2(n4811), .ZN(n4290)
         );
  OAI211_X1 U4085 ( .C1(n5293), .C2(n3723), .A(n3552), .B(n4290), .ZN(n5249)
         );
  INV_X1 U4086 ( .A(n5249), .ZN(n3561) );
  AOI21_X2 U4087 ( .B1(n3554), .B2(n3553), .A(n2534), .ZN(n3588) );
  XNOR2_X1 U4088 ( .A(n3588), .B(n4365), .ZN(n5251) );
  NAND2_X1 U4089 ( .A1(n5251), .A2(n4837), .ZN(n3560) );
  OR2_X1 U4090 ( .A1(n3555), .A2(n3723), .ZN(n3556) );
  AND3_X1 U4091 ( .A1(n4838), .A2(n3556), .A3(n5304), .ZN(n5250) );
  INV_X1 U4092 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3557) );
  OAI22_X1 U4093 ( .A1(n5173), .A2(n3557), .B1(n4295), .B2(n5216), .ZN(n3558)
         );
  AOI21_X1 U4094 ( .B1(n5250), .B2(n4843), .A(n3558), .ZN(n3559) );
  OAI211_X1 U4095 ( .C1(n4847), .C2(n3561), .A(n3560), .B(n3559), .ZN(U3273)
         );
  OAI22_X1 U4096 ( .A1(n3564), .A2(n3845), .B1(n3562), .B2(n3719), .ZN(n3563)
         );
  XNOR2_X1 U4097 ( .A(n3563), .B(n3843), .ZN(n3568) );
  OR2_X1 U4098 ( .A1(n3564), .A2(n3842), .ZN(n3566) );
  NAND2_X1 U4099 ( .A1(n3582), .A2(n3127), .ZN(n3565) );
  NAND2_X1 U4100 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  NOR2_X1 U4101 ( .A1(n3568), .A2(n3567), .ZN(n3718) );
  AOI21_X1 U4102 ( .B1(n3568), .B2(n3567), .A(n3718), .ZN(n3576) );
  NAND2_X1 U4103 ( .A1(n3569), .A2(n3570), .ZN(n3573) );
  INV_X1 U4104 ( .A(n3569), .ZN(n3572) );
  INV_X1 U4105 ( .A(n3570), .ZN(n3571) );
  AOI21_X1 U4106 ( .B1(n3574), .B2(n3573), .A(n2711), .ZN(n3575) );
  NAND2_X1 U4107 ( .A1(n3575), .A2(n3576), .ZN(n3730) );
  OAI21_X1 U4108 ( .B1(n3576), .B2(n3575), .A(n3730), .ZN(n3577) );
  NAND2_X1 U4109 ( .A1(n3577), .A2(n5274), .ZN(n3584) );
  INV_X1 U4110 ( .A(n3578), .ZN(n3580) );
  NOR2_X1 U4111 ( .A1(n4116), .A2(STATE_REG_SCAN_IN), .ZN(n4628) );
  INV_X1 U4112 ( .A(n4628), .ZN(n3579) );
  OAI21_X1 U4113 ( .B1(n3580), .B2(n4345), .A(n3579), .ZN(n3581) );
  AOI21_X1 U4114 ( .B1(n3582), .B2(n5263), .A(n3581), .ZN(n3583) );
  OAI211_X1 U4115 ( .C1(n5279), .C2(n3585), .A(n3584), .B(n3583), .ZN(U3223)
         );
  INV_X1 U4116 ( .A(n4811), .ZN(n3591) );
  NAND2_X1 U4117 ( .A1(n3535), .A2(IR_REG_31__SCAN_IN), .ZN(n3589) );
  XNOR2_X1 U4118 ( .A(n3589), .B(IR_REG_18__SCAN_IN), .ZN(n4917) );
  INV_X1 U4119 ( .A(n4917), .ZN(n4647) );
  INV_X1 U4120 ( .A(DATAI_18_), .ZN(n3590) );
  MUX2_X1 U4121 ( .A(n4647), .B(n3590), .S(n4404), .Z(n4833) );
  NAND2_X1 U4122 ( .A1(n3591), .A2(n4839), .ZN(n3693) );
  NAND2_X1 U4123 ( .A1(n4811), .A2(n4833), .ZN(n4807) );
  NAND2_X1 U4124 ( .A1(n3693), .A2(n4807), .ZN(n4835) );
  NAND2_X1 U4125 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U4126 ( .A1(n3130), .A2(REG1_REG_19__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4127 ( .A1(n4375), .A2(REG0_REG_19__SCAN_IN), .ZN(n3597) );
  INV_X1 U4128 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4271) );
  AND2_X1 U4129 ( .A1(n3593), .A2(n4271), .ZN(n3594) );
  NOR2_X1 U4130 ( .A1(n3602), .A2(n3594), .ZN(n4269) );
  NAND2_X1 U4131 ( .A1(n3612), .A2(n4269), .ZN(n3596) );
  NAND2_X1 U4132 ( .A1(n2940), .A2(REG2_REG_19__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4133 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n5264)
         );
  INV_X1 U4134 ( .A(n5264), .ZN(n3742) );
  INV_X1 U4135 ( .A(DATAI_19_), .ZN(n3599) );
  MUX2_X1 U4136 ( .A(n4848), .B(n3599), .S(n4404), .Z(n4820) );
  NAND2_X1 U4137 ( .A1(n3742), .A2(n4820), .ZN(n3601) );
  NAND2_X1 U4138 ( .A1(n5264), .A2(n4270), .ZN(n3600) );
  NAND2_X1 U4139 ( .A1(n3602), .A2(REG3_REG_20__SCAN_IN), .ZN(n3610) );
  OR2_X1 U4140 ( .A1(n3602), .A2(REG3_REG_20__SCAN_IN), .ZN(n3603) );
  NAND2_X1 U4141 ( .A1(n3610), .A2(n3603), .ZN(n5278) );
  INV_X1 U4142 ( .A(n5278), .ZN(n4800) );
  NAND2_X1 U4143 ( .A1(n4800), .A2(n3612), .ZN(n3607) );
  NAND2_X1 U4144 ( .A1(n4375), .A2(REG0_REG_20__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4145 ( .A1(n3130), .A2(REG1_REG_20__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4146 ( .A1(n2940), .A2(REG2_REG_20__SCAN_IN), .ZN(n3604) );
  INV_X1 U4147 ( .A(n4810), .ZN(n3608) );
  NAND2_X1 U4148 ( .A1(n4404), .A2(DATAI_20_), .ZN(n3752) );
  NAND2_X1 U4149 ( .A1(n3608), .A2(n5262), .ZN(n4411) );
  NAND2_X1 U4150 ( .A1(n4810), .A2(n3752), .ZN(n4487) );
  NAND2_X1 U4151 ( .A1(n4411), .A2(n4487), .ZN(n4793) );
  NAND2_X1 U4152 ( .A1(n4789), .A2(n3609), .ZN(n4775) );
  INV_X1 U4153 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4112) );
  NAND2_X1 U4154 ( .A1(n3610), .A2(n4112), .ZN(n3611) );
  AND2_X1 U4155 ( .A1(n3619), .A2(n3611), .ZN(n4784) );
  NAND2_X1 U4156 ( .A1(n4784), .A2(n3612), .ZN(n3616) );
  NAND2_X1 U4157 ( .A1(n4375), .A2(REG0_REG_21__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4158 ( .A1(n2938), .A2(REG1_REG_21__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4159 ( .A1(n2940), .A2(REG2_REG_21__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4160 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n4526)
         );
  NAND2_X1 U4161 ( .A1(n4404), .A2(DATAI_21_), .ZN(n4783) );
  AND2_X1 U4162 ( .A1(n4526), .A2(n4783), .ZN(n4757) );
  OR2_X1 U4163 ( .A1(n4526), .A2(n4783), .ZN(n3698) );
  INV_X1 U4164 ( .A(n3698), .ZN(n3617) );
  NAND2_X1 U4165 ( .A1(n4775), .A2(n4777), .ZN(n4774) );
  INV_X1 U4166 ( .A(n4783), .ZN(n3618) );
  INV_X1 U4167 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4325) );
  INV_X1 U4168 ( .A(n3626), .ZN(n3627) );
  NAND2_X1 U4169 ( .A1(n3619), .A2(n4325), .ZN(n3620) );
  NAND2_X1 U4170 ( .A1(n3627), .A2(n3620), .ZN(n4768) );
  INV_X1 U4171 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U4172 ( .A1(n3130), .A2(REG1_REG_22__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4173 ( .A1(n4375), .A2(REG0_REG_22__SCAN_IN), .ZN(n3621) );
  OAI211_X1 U4174 ( .C1(n4769), .C2(n3666), .A(n3622), .B(n3621), .ZN(n3623)
         );
  INV_X1 U4175 ( .A(n3623), .ZN(n3624) );
  NAND2_X1 U4176 ( .A1(n4404), .A2(DATAI_22_), .ZN(n4765) );
  OR2_X1 U4177 ( .A1(n4525), .A2(n4765), .ZN(n4740) );
  NAND2_X1 U4178 ( .A1(n4525), .A2(n4765), .ZN(n3699) );
  INV_X1 U4179 ( .A(n3636), .ZN(n3637) );
  INV_X1 U4180 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U4181 ( .A1(n3627), .A2(n4100), .ZN(n3628) );
  NAND2_X1 U4182 ( .A1(n4749), .A2(n3612), .ZN(n3634) );
  INV_X1 U4183 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3631) );
  NAND2_X1 U4184 ( .A1(n3130), .A2(REG1_REG_23__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4185 ( .A1(n4375), .A2(REG0_REG_23__SCAN_IN), .ZN(n3629) );
  OAI211_X1 U4186 ( .C1(n3631), .C2(n3666), .A(n3630), .B(n3629), .ZN(n3632)
         );
  INV_X1 U4187 ( .A(n3632), .ZN(n3633) );
  NAND2_X1 U4188 ( .A1(n4404), .A2(DATAI_23_), .ZN(n4748) );
  INV_X1 U4189 ( .A(n4748), .ZN(n3635) );
  INV_X1 U4190 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U4191 ( .A1(n3637), .A2(n4302), .ZN(n3638) );
  NAND2_X1 U4192 ( .A1(n3652), .A2(n3638), .ZN(n4731) );
  INV_X1 U4193 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U4194 ( .A1(n4375), .A2(REG0_REG_24__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U4195 ( .A1(n3130), .A2(REG1_REG_24__SCAN_IN), .ZN(n3639) );
  OAI211_X1 U4196 ( .C1(n4730), .C2(n3666), .A(n3640), .B(n3639), .ZN(n3641)
         );
  INV_X1 U4197 ( .A(n3641), .ZN(n3642) );
  AND2_X1 U4198 ( .A1(n4404), .A2(DATAI_24_), .ZN(n3711) );
  NOR2_X1 U4199 ( .A1(n4524), .A2(n3711), .ZN(n3644) );
  XNOR2_X1 U4200 ( .A(n3652), .B(REG3_REG_25__SCAN_IN), .ZN(n4280) );
  NAND2_X1 U4201 ( .A1(n4280), .A2(n3612), .ZN(n3649) );
  INV_X1 U4202 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4203 ( .A1(n4375), .A2(REG0_REG_25__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4204 ( .A1(n3130), .A2(REG1_REG_25__SCAN_IN), .ZN(n3645) );
  OAI211_X1 U4205 ( .C1(n3805), .C2(n3666), .A(n3646), .B(n3645), .ZN(n3647)
         );
  INV_X1 U4206 ( .A(n3647), .ZN(n3648) );
  NAND2_X1 U4207 ( .A1(n4404), .A2(DATAI_25_), .ZN(n3826) );
  OR2_X1 U4208 ( .A1(n4726), .A2(n3826), .ZN(n4707) );
  NAND2_X1 U4209 ( .A1(n4726), .A2(n3826), .ZN(n4461) );
  NAND2_X1 U4210 ( .A1(n4707), .A2(n4461), .ZN(n4408) );
  INV_X1 U4211 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3651) );
  INV_X1 U4212 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3650) );
  OAI21_X1 U4213 ( .B1(n3652), .B2(n3651), .A(n3650), .ZN(n3653) );
  AND2_X1 U4214 ( .A1(n3653), .A2(n3662), .ZN(n4357) );
  NAND2_X1 U4215 ( .A1(n4357), .A2(n3612), .ZN(n3658) );
  INV_X1 U4216 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U4217 ( .A1(n4375), .A2(REG0_REG_26__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4218 ( .A1(n3130), .A2(REG1_REG_26__SCAN_IN), .ZN(n3654) );
  OAI211_X1 U4219 ( .C1(n4704), .C2(n3666), .A(n3655), .B(n3654), .ZN(n3656)
         );
  INV_X1 U4220 ( .A(n3656), .ZN(n3657) );
  AND2_X1 U4221 ( .A1(n4404), .A2(DATAI_26_), .ZN(n4703) );
  NAND2_X1 U4222 ( .A1(n4523), .A2(n4703), .ZN(n3659) );
  INV_X1 U4223 ( .A(n3662), .ZN(n3660) );
  NAND2_X1 U4224 ( .A1(n3660), .A2(REG3_REG_27__SCAN_IN), .ZN(n3673) );
  INV_X1 U4225 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4226 ( .A1(n3662), .A2(n3661), .ZN(n3663) );
  NAND2_X1 U4227 ( .A1(n3673), .A2(n3663), .ZN(n4694) );
  INV_X1 U4228 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U4229 ( .A1(n3130), .A2(REG1_REG_27__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4230 ( .A1(n4375), .A2(REG0_REG_27__SCAN_IN), .ZN(n3664) );
  OAI211_X1 U4231 ( .C1(n4693), .C2(n3666), .A(n3665), .B(n3664), .ZN(n3667)
         );
  INV_X1 U4232 ( .A(n3667), .ZN(n3668) );
  NAND2_X1 U4233 ( .A1(n4404), .A2(DATAI_27_), .ZN(n4690) );
  NAND2_X1 U4234 ( .A1(n4712), .A2(n4690), .ZN(n3671) );
  NOR2_X1 U4235 ( .A1(n4712), .A2(n4690), .ZN(n3670) );
  INV_X1 U4236 ( .A(n3673), .ZN(n3672) );
  NAND2_X1 U4237 ( .A1(n3672), .A2(REG3_REG_28__SCAN_IN), .ZN(n4667) );
  INV_X1 U4238 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3912) );
  NAND2_X1 U4239 ( .A1(n3673), .A2(n3912), .ZN(n3674) );
  NAND2_X1 U4240 ( .A1(n4667), .A2(n3674), .ZN(n3851) );
  NAND2_X1 U4241 ( .A1(n2940), .A2(REG2_REG_28__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4242 ( .A1(n3130), .A2(REG1_REG_28__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4243 ( .A1(n4375), .A2(REG0_REG_28__SCAN_IN), .ZN(n3675) );
  AND2_X1 U4244 ( .A1(n4404), .A2(DATAI_28_), .ZN(n3848) );
  XNOR2_X1 U4245 ( .A(n4521), .B(n3848), .ZN(n4662) );
  XNOR2_X1 U4246 ( .A(n4663), .B(n4662), .ZN(n4862) );
  OR2_X1 U4247 ( .A1(n4667), .A2(n3680), .ZN(n3686) );
  INV_X1 U4248 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4249 ( .A1(n2940), .A2(REG2_REG_29__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4250 ( .A1(n4375), .A2(REG0_REG_29__SCAN_IN), .ZN(n3681) );
  OAI211_X1 U4251 ( .C1(n3683), .C2(n2966), .A(n3682), .B(n3681), .ZN(n3684)
         );
  INV_X1 U4252 ( .A(n3684), .ZN(n3685) );
  INV_X1 U4253 ( .A(n3848), .ZN(n4661) );
  OAI22_X1 U4254 ( .A1(n4712), .A2(n5154), .B1(n5293), .B2(n4661), .ZN(n3710)
         );
  NAND2_X1 U4255 ( .A1(n5264), .A2(n4820), .ZN(n3687) );
  AND2_X1 U4256 ( .A1(n4807), .A2(n3687), .ZN(n3695) );
  NAND2_X1 U4257 ( .A1(n4527), .A2(n3723), .ZN(n3688) );
  AND2_X1 U4258 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  NAND2_X1 U4259 ( .A1(n3691), .A2(n4483), .ZN(n3697) );
  NAND2_X1 U4260 ( .A1(n3692), .A2(n4292), .ZN(n4826) );
  NAND2_X1 U4261 ( .A1(n4826), .A2(n3693), .ZN(n3696) );
  NOR2_X1 U4262 ( .A1(n5264), .A2(n4820), .ZN(n3694) );
  AOI21_X1 U4263 ( .B1(n3696), .B2(n3695), .A(n3694), .ZN(n4412) );
  AND2_X1 U4264 ( .A1(n4740), .A2(n3698), .ZN(n4493) );
  NAND2_X1 U4265 ( .A1(n4763), .A2(n4748), .ZN(n3700) );
  AND2_X1 U4266 ( .A1(n3700), .A2(n3699), .ZN(n4459) );
  NAND2_X1 U4267 ( .A1(n4740), .A2(n4757), .ZN(n3701) );
  NAND2_X1 U4268 ( .A1(n4459), .A2(n3701), .ZN(n4494) );
  INV_X1 U4269 ( .A(n4494), .ZN(n3702) );
  NAND2_X1 U4270 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  OR2_X1 U4271 ( .A1(n4763), .A2(n4748), .ZN(n4456) );
  NAND2_X1 U4272 ( .A1(n3704), .A2(n4456), .ZN(n4722) );
  INV_X1 U4273 ( .A(n3711), .ZN(n4728) );
  NAND2_X1 U4274 ( .A1(n4524), .A2(n4728), .ZN(n4462) );
  NAND2_X1 U4275 ( .A1(n4407), .A2(n3711), .ZN(n4457) );
  NAND2_X1 U4276 ( .A1(n4684), .A2(n4703), .ZN(n4400) );
  NAND2_X1 U4277 ( .A1(n4400), .A2(n4707), .ZN(n4495) );
  INV_X1 U4278 ( .A(n4495), .ZN(n3705) );
  NOR2_X1 U4279 ( .A1(n4684), .A2(n4703), .ZN(n4465) );
  INV_X1 U4280 ( .A(n4690), .ZN(n4260) );
  NOR2_X1 U4281 ( .A1(n4712), .A2(n4260), .ZN(n4464) );
  NOR2_X1 U4282 ( .A1(n4522), .A2(n4690), .ZN(n3706) );
  NOR2_X1 U4283 ( .A1(n4464), .A2(n3706), .ZN(n4688) );
  INV_X1 U4284 ( .A(n3706), .ZN(n4473) );
  NAND3_X1 U4285 ( .A1(n4681), .A2(n4662), .A3(n4473), .ZN(n4670) );
  INV_X1 U4286 ( .A(n4670), .ZN(n3708) );
  AOI21_X1 U4287 ( .B1(n4681), .B2(n4473), .A(n4662), .ZN(n3707) );
  NOR3_X1 U4288 ( .A1(n3708), .A2(n3707), .A3(n5206), .ZN(n3709) );
  INV_X1 U4289 ( .A(n4861), .ZN(n3716) );
  NAND2_X1 U4290 ( .A1(n4767), .A2(n4748), .ZN(n4747) );
  INV_X1 U4291 ( .A(n4692), .ZN(n3712) );
  OAI211_X1 U4292 ( .C1(n3712), .C2(n4661), .A(n5304), .B(n2523), .ZN(n4860)
         );
  INV_X1 U4293 ( .A(n3851), .ZN(n3713) );
  INV_X1 U4294 ( .A(n5173), .ZN(n5285) );
  AOI22_X1 U4295 ( .A1(n3713), .A2(n5168), .B1(REG2_REG_28__SCAN_IN), .B2(
        n5285), .ZN(n3714) );
  OAI21_X1 U4296 ( .B1(n4860), .B2(n4802), .A(n3714), .ZN(n3715) );
  AOI21_X1 U4297 ( .B1(n3716), .B2(n5173), .A(n3715), .ZN(n3717) );
  OAI21_X1 U4298 ( .B1(n4862), .B2(n4806), .A(n3717), .ZN(U3262) );
  OAI22_X1 U4299 ( .A1(n4407), .A2(n5200), .B1(n3765), .B2(n5154), .ZN(n4744)
         );
  INV_X1 U4300 ( .A(n4744), .ZN(n3780) );
  INV_X1 U4301 ( .A(n3718), .ZN(n4288) );
  NAND2_X1 U4302 ( .A1(n4527), .A2(n3127), .ZN(n3721) );
  OR2_X1 U4303 ( .A1(n3723), .A2(n3719), .ZN(n3720) );
  NAND2_X1 U4304 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  XNOR2_X1 U4305 ( .A(n3722), .B(n3824), .ZN(n3725) );
  NOR2_X1 U4306 ( .A1(n3723), .A2(n3845), .ZN(n3724) );
  AOI21_X1 U4307 ( .B1(n4527), .B2(n3828), .A(n3724), .ZN(n3726) );
  NAND2_X1 U4308 ( .A1(n3725), .A2(n3726), .ZN(n3731) );
  INV_X1 U4309 ( .A(n3725), .ZN(n3728) );
  INV_X1 U4310 ( .A(n3726), .ZN(n3727) );
  NAND2_X1 U4311 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  NAND2_X1 U4312 ( .A1(n3731), .A2(n3729), .ZN(n4287) );
  INV_X1 U4313 ( .A(n3731), .ZN(n4342) );
  NAND2_X1 U4314 ( .A1(n4811), .A2(n3127), .ZN(n3733) );
  OR2_X1 U4315 ( .A1(n4833), .A2(n3719), .ZN(n3732) );
  NAND2_X1 U4316 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  XNOR2_X1 U4317 ( .A(n3734), .B(n3824), .ZN(n3736) );
  NOR2_X1 U4318 ( .A1(n4833), .A2(n3845), .ZN(n3735) );
  AOI21_X1 U4319 ( .B1(n4811), .B2(n3828), .A(n3735), .ZN(n3737) );
  NAND2_X1 U4320 ( .A1(n3736), .A2(n3737), .ZN(n3741) );
  INV_X1 U4321 ( .A(n3736), .ZN(n3739) );
  INV_X1 U4322 ( .A(n3737), .ZN(n3738) );
  NAND2_X1 U4323 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  AND2_X1 U4324 ( .A1(n3741), .A2(n3740), .ZN(n4341) );
  NAND2_X1 U4325 ( .A1(n4340), .A2(n3741), .ZN(n4267) );
  OAI22_X1 U4326 ( .A1(n3742), .A2(n3842), .B1(n4820), .B2(n3845), .ZN(n3746)
         );
  NAND2_X1 U4327 ( .A1(n5264), .A2(n3127), .ZN(n3744) );
  OR2_X1 U4328 ( .A1(n4820), .A2(n3719), .ZN(n3743) );
  NAND2_X1 U4329 ( .A1(n3744), .A2(n3743), .ZN(n3745) );
  XNOR2_X1 U4330 ( .A(n3745), .B(n3843), .ZN(n3747) );
  XOR2_X1 U4331 ( .A(n3746), .B(n3747), .Z(n4268) );
  NAND2_X1 U4332 ( .A1(n4810), .A2(n3127), .ZN(n3750) );
  OR2_X1 U4333 ( .A1(n3752), .A2(n3719), .ZN(n3749) );
  NAND2_X1 U4334 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  XNOR2_X1 U4335 ( .A(n3751), .B(n3824), .ZN(n3755) );
  NOR2_X1 U4336 ( .A1(n3752), .A2(n3845), .ZN(n3753) );
  AOI21_X1 U4337 ( .B1(n4810), .B2(n3828), .A(n3753), .ZN(n3754) );
  OR2_X1 U4338 ( .A1(n3755), .A2(n3754), .ZN(n5267) );
  NAND2_X1 U4339 ( .A1(n3755), .A2(n3754), .ZN(n5266) );
  NAND2_X1 U4340 ( .A1(n4526), .A2(n3310), .ZN(n3757) );
  OR2_X1 U4341 ( .A1(n4783), .A2(n3719), .ZN(n3756) );
  NAND2_X1 U4342 ( .A1(n3757), .A2(n3756), .ZN(n3758) );
  XNOR2_X1 U4343 ( .A(n3758), .B(n3843), .ZN(n3782) );
  NAND2_X1 U4344 ( .A1(n4526), .A2(n3828), .ZN(n3760) );
  OR2_X1 U4345 ( .A1(n3845), .A2(n4783), .ZN(n3759) );
  NAND2_X1 U4346 ( .A1(n3760), .A2(n3759), .ZN(n3781) );
  NOR2_X1 U4347 ( .A1(n3782), .A2(n3781), .ZN(n3763) );
  INV_X1 U4348 ( .A(n3782), .ZN(n3762) );
  INV_X1 U4349 ( .A(n3781), .ZN(n3761) );
  OAI22_X1 U4350 ( .A1(n3765), .A2(n3845), .B1(n3719), .B2(n4765), .ZN(n3764)
         );
  XNOR2_X1 U4351 ( .A(n3764), .B(n3843), .ZN(n3767) );
  OAI22_X1 U4352 ( .A1(n3765), .A2(n3842), .B1(n3845), .B2(n4765), .ZN(n3766)
         );
  XNOR2_X1 U4353 ( .A(n3767), .B(n3766), .ZN(n4323) );
  INV_X1 U4354 ( .A(n3775), .ZN(n4321) );
  NOR2_X1 U4355 ( .A1(n3767), .A2(n3766), .ZN(n3772) );
  NAND2_X1 U4356 ( .A1(n4763), .A2(n3127), .ZN(n3769) );
  OR2_X1 U4357 ( .A1(n4748), .A2(n3719), .ZN(n3768) );
  NAND2_X1 U4358 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  XNOR2_X1 U4359 ( .A(n3770), .B(n3824), .ZN(n3815) );
  NOR2_X1 U4360 ( .A1(n4748), .A2(n3845), .ZN(n3771) );
  AOI21_X1 U4361 ( .B1(n4763), .B2(n3828), .A(n3771), .ZN(n3814) );
  XNOR2_X1 U4362 ( .A(n3815), .B(n3814), .ZN(n3773) );
  OAI21_X1 U4363 ( .B1(n4321), .B2(n3772), .A(n3773), .ZN(n3776) );
  NOR2_X1 U4364 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  NAND3_X1 U4365 ( .A1(n3776), .A2(n5274), .A3(n3820), .ZN(n3779) );
  OAI22_X1 U4366 ( .A1(n4324), .A2(n4748), .B1(STATE_REG_SCAN_IN), .B2(n4100), 
        .ZN(n3777) );
  AOI21_X1 U4367 ( .B1(n4749), .B2(n4317), .A(n3777), .ZN(n3778) );
  OAI211_X1 U4368 ( .C1(n3780), .C2(n4345), .A(n3779), .B(n3778), .ZN(U3213)
         );
  XNOR2_X1 U4369 ( .A(n3782), .B(n3781), .ZN(n3783) );
  XNOR2_X1 U4370 ( .A(n3784), .B(n3783), .ZN(n3788) );
  OAI22_X1 U4371 ( .A1(n4324), .A2(n4783), .B1(STATE_REG_SCAN_IN), .B2(n4112), 
        .ZN(n3786) );
  AOI22_X1 U4372 ( .A1(n4525), .A2(n4809), .B1(n5204), .B2(n4810), .ZN(n4779)
         );
  NOR2_X1 U4373 ( .A1(n4779), .A2(n4345), .ZN(n3785) );
  AOI211_X1 U4374 ( .C1(n4317), .C2(n4784), .A(n3786), .B(n3785), .ZN(n3787)
         );
  OAI21_X1 U4375 ( .B1(n3788), .B2(n4363), .A(n3787), .ZN(U3220) );
  AND2_X1 U4376 ( .A1(n3789), .A2(n3790), .ZN(n3793) );
  OAI211_X1 U4377 ( .C1(n3793), .C2(n3792), .A(n5274), .B(n3791), .ZN(n3800)
         );
  NOR2_X1 U4378 ( .A1(n4324), .A2(n3794), .ZN(n3795) );
  AOI211_X1 U4379 ( .C1(n3798), .C2(n3797), .A(n3796), .B(n3795), .ZN(n3799)
         );
  OAI211_X1 U4380 ( .C1(n5279), .C2(n3801), .A(n3800), .B(n3799), .ZN(U3214)
         );
  XNOR2_X1 U4381 ( .A(n3802), .B(n4408), .ZN(n4874) );
  AND2_X1 U4382 ( .A1(n4727), .A2(n4279), .ZN(n3803) );
  NOR2_X1 U4383 ( .A1(n4700), .A2(n3803), .ZN(n4872) );
  NAND2_X1 U4384 ( .A1(n4280), .A2(n5168), .ZN(n3804) );
  OAI21_X1 U4385 ( .B1(n5173), .B2(n3805), .A(n3804), .ZN(n3806) );
  AOI21_X1 U4386 ( .B1(n4872), .B2(n5300), .A(n3806), .ZN(n3813) );
  OAI21_X1 U4387 ( .B1(n2599), .B2(n3807), .A(n4708), .ZN(n3808) );
  NAND2_X1 U4388 ( .A1(n3808), .A2(n5151), .ZN(n3811) );
  OAI22_X1 U4389 ( .A1(n4407), .A2(n5154), .B1(n3826), .B2(n5293), .ZN(n3809)
         );
  AOI21_X1 U4390 ( .B1(n4523), .B2(n4809), .A(n3809), .ZN(n3810) );
  NAND2_X1 U4391 ( .A1(n3811), .A2(n3810), .ZN(n4871) );
  NAND2_X1 U4392 ( .A1(n4871), .A2(n5173), .ZN(n3812) );
  OAI211_X1 U4393 ( .C1(n4874), .C2(n4806), .A(n3813), .B(n3812), .ZN(U3265)
         );
  OR2_X1 U4394 ( .A1(n3815), .A2(n3814), .ZN(n3818) );
  OAI22_X1 U4395 ( .A1(n4407), .A2(n3845), .B1(n3456), .B2(n4728), .ZN(n3816)
         );
  XNOR2_X1 U4396 ( .A(n3816), .B(n3824), .ZN(n3819) );
  OAI22_X1 U4397 ( .A1(n4407), .A2(n3842), .B1(n3446), .B2(n4728), .ZN(n4300)
         );
  INV_X1 U4398 ( .A(n4300), .ZN(n3817) );
  NAND2_X1 U4399 ( .A1(n4297), .A2(n3817), .ZN(n3821) );
  NAND3_X1 U4400 ( .A1(n3820), .A2(n3819), .A3(n3818), .ZN(n4296) );
  NAND2_X1 U4401 ( .A1(n3821), .A2(n4296), .ZN(n4350) );
  NAND2_X1 U4402 ( .A1(n4726), .A2(n3127), .ZN(n3823) );
  OR2_X1 U4403 ( .A1(n3826), .A2(n3719), .ZN(n3822) );
  NAND2_X1 U4404 ( .A1(n3823), .A2(n3822), .ZN(n3825) );
  XNOR2_X1 U4405 ( .A(n3825), .B(n3824), .ZN(n3830) );
  NOR2_X1 U4406 ( .A1(n3826), .A2(n3845), .ZN(n3827) );
  AOI21_X1 U4407 ( .B1(n4726), .B2(n3828), .A(n3827), .ZN(n3831) );
  AND2_X1 U4408 ( .A1(n3830), .A2(n3831), .ZN(n4349) );
  OAI22_X1 U4409 ( .A1(n4684), .A2(n3845), .B1(n3719), .B2(n4711), .ZN(n3829)
         );
  XNOR2_X1 U4410 ( .A(n3829), .B(n3843), .ZN(n4353) );
  OAI22_X1 U4411 ( .A1(n4684), .A2(n3842), .B1(n3845), .B2(n4711), .ZN(n4354)
         );
  NOR2_X1 U4412 ( .A1(n4353), .A2(n4354), .ZN(n3836) );
  OR2_X1 U4413 ( .A1(n4349), .A2(n3836), .ZN(n3838) );
  INV_X1 U4414 ( .A(n3830), .ZN(n3833) );
  INV_X1 U4415 ( .A(n3831), .ZN(n3832) );
  NAND2_X1 U4416 ( .A1(n3833), .A2(n3832), .ZN(n4351) );
  NAND2_X1 U4417 ( .A1(n4353), .A2(n4354), .ZN(n3834) );
  AND2_X1 U4418 ( .A1(n4351), .A2(n3834), .ZN(n3835) );
  OR2_X1 U4419 ( .A1(n3836), .A2(n3835), .ZN(n3837) );
  OAI22_X1 U4420 ( .A1(n4712), .A2(n3842), .B1(n3845), .B2(n4690), .ZN(n3840)
         );
  OAI22_X1 U4421 ( .A1(n4712), .A2(n3845), .B1(n3719), .B2(n4690), .ZN(n3839)
         );
  XNOR2_X1 U4422 ( .A(n3839), .B(n3843), .ZN(n3841) );
  XOR2_X1 U4423 ( .A(n3840), .B(n3841), .Z(n4259) );
  OAI22_X1 U4424 ( .A1(n4683), .A2(n3842), .B1(n4661), .B2(n3845), .ZN(n3844)
         );
  XNOR2_X1 U4425 ( .A(n3844), .B(n3843), .ZN(n3847) );
  OAI22_X1 U4426 ( .A1(n4683), .A2(n3845), .B1(n4661), .B2(n3456), .ZN(n3846)
         );
  NAND2_X1 U4427 ( .A1(n4522), .A2(n5265), .ZN(n3850) );
  AOI22_X1 U4428 ( .A1(n5263), .A2(n3848), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3849) );
  OAI211_X1 U4429 ( .C1(n3851), .C2(n5279), .A(n3850), .B(n3849), .ZN(n3852)
         );
  AOI21_X1 U4430 ( .B1(n4358), .B2(n4520), .A(n3852), .ZN(n3853) );
  OAI21_X1 U4431 ( .B1(n3854), .B2(n4363), .A(n3853), .ZN(n4257) );
  XOR2_X1 U4432 ( .A(DATAI_30_), .B(keyinput_1), .Z(n3858) );
  XOR2_X1 U4433 ( .A(DATAI_31_), .B(keyinput_0), .Z(n3857) );
  XNOR2_X1 U4434 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n3856) );
  XOR2_X1 U4435 ( .A(DATAI_28_), .B(keyinput_3), .Z(n3855) );
  AOI211_X1 U4436 ( .C1(n3858), .C2(n3857), .A(n3856), .B(n3855), .ZN(n3861)
         );
  XOR2_X1 U4437 ( .A(DATAI_27_), .B(keyinput_4), .Z(n3860) );
  XNOR2_X1 U4438 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n3859) );
  NOR3_X1 U4439 ( .A1(n3861), .A2(n3860), .A3(n3859), .ZN(n3864) );
  XOR2_X1 U4440 ( .A(DATAI_24_), .B(keyinput_7), .Z(n3863) );
  XNOR2_X1 U4441 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n3862) );
  NOR3_X1 U4442 ( .A1(n3864), .A2(n3863), .A3(n3862), .ZN(n3867) );
  XOR2_X1 U4443 ( .A(DATAI_23_), .B(keyinput_8), .Z(n3866) );
  XNOR2_X1 U4444 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n3865) );
  OAI21_X1 U4445 ( .B1(n3867), .B2(n3866), .A(n3865), .ZN(n3874) );
  XOR2_X1 U4446 ( .A(DATAI_21_), .B(keyinput_10), .Z(n3873) );
  XOR2_X1 U4447 ( .A(DATAI_20_), .B(keyinput_11), .Z(n3871) );
  XNOR2_X1 U4448 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n3870) );
  XNOR2_X1 U4449 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n3869) );
  XNOR2_X1 U4450 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n3868) );
  NAND4_X1 U4451 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3872)
         );
  AOI21_X1 U4452 ( .B1(n3874), .B2(n3873), .A(n3872), .ZN(n3877) );
  XOR2_X1 U4453 ( .A(DATAI_16_), .B(keyinput_15), .Z(n3876) );
  XNOR2_X1 U4454 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n3875) );
  OAI21_X1 U4455 ( .B1(n3877), .B2(n3876), .A(n3875), .ZN(n3880) );
  XNOR2_X1 U4456 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n3879) );
  XOR2_X1 U4457 ( .A(DATAI_13_), .B(keyinput_18), .Z(n3878) );
  AOI21_X1 U4458 ( .B1(n3880), .B2(n3879), .A(n3878), .ZN(n3883) );
  XNOR2_X1 U4459 ( .A(n4073), .B(keyinput_19), .ZN(n3882) );
  XNOR2_X1 U4460 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n3881) );
  OAI21_X1 U4461 ( .B1(n3883), .B2(n3882), .A(n3881), .ZN(n3886) );
  XOR2_X1 U4462 ( .A(DATAI_10_), .B(keyinput_21), .Z(n3885) );
  XOR2_X1 U4463 ( .A(DATAI_9_), .B(keyinput_22), .Z(n3884) );
  AOI21_X1 U4464 ( .B1(n3886), .B2(n3885), .A(n3884), .ZN(n3890) );
  XOR2_X1 U4465 ( .A(DATAI_8_), .B(keyinput_23), .Z(n3889) );
  XNOR2_X1 U4466 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n3888) );
  XNOR2_X1 U4467 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n3887) );
  OAI211_X1 U4468 ( .C1(n3890), .C2(n3889), .A(n3888), .B(n3887), .ZN(n3893)
         );
  XOR2_X1 U4469 ( .A(DATAI_5_), .B(keyinput_26), .Z(n3892) );
  XOR2_X1 U4470 ( .A(DATAI_4_), .B(keyinput_27), .Z(n3891) );
  AOI21_X1 U4471 ( .B1(n3893), .B2(n3892), .A(n3891), .ZN(n3901) );
  XOR2_X1 U4472 ( .A(DATAI_3_), .B(keyinput_28), .Z(n3900) );
  XOR2_X1 U4473 ( .A(DATAI_0_), .B(keyinput_31), .Z(n3898) );
  XNOR2_X1 U4474 ( .A(n3894), .B(keyinput_30), .ZN(n3897) );
  XNOR2_X1 U4475 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n3896) );
  XNOR2_X1 U4476 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n3895) );
  NOR4_X1 U4477 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  OAI21_X1 U4478 ( .B1(n3901), .B2(n3900), .A(n3899), .ZN(n3904) );
  XNOR2_X1 U4479 ( .A(n4093), .B(keyinput_33), .ZN(n3903) );
  XNOR2_X1 U4480 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_34), .ZN(n3902) );
  AOI21_X1 U4481 ( .B1(n3904), .B2(n3903), .A(n3902), .ZN(n3908) );
  XNOR2_X1 U4482 ( .A(n3905), .B(keyinput_35), .ZN(n3907) );
  XNOR2_X1 U4483 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_36), .ZN(n3906) );
  OAI21_X1 U4484 ( .B1(n3908), .B2(n3907), .A(n3906), .ZN(n3911) );
  XNOR2_X1 U4485 ( .A(n4101), .B(keyinput_38), .ZN(n3910) );
  XNOR2_X1 U4486 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .ZN(n3909) );
  NAND3_X1 U4487 ( .A1(n3911), .A2(n3910), .A3(n3909), .ZN(n3915) );
  XNOR2_X1 U4488 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n3914) );
  XNOR2_X1 U4489 ( .A(n3912), .B(keyinput_40), .ZN(n3913) );
  AOI21_X1 U4490 ( .B1(n3915), .B2(n3914), .A(n3913), .ZN(n3919) );
  XNOR2_X1 U4491 ( .A(n3916), .B(keyinput_41), .ZN(n3918) );
  XOR2_X1 U4492 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .Z(n3917) );
  NOR3_X1 U4493 ( .A1(n3919), .A2(n3918), .A3(n3917), .ZN(n3922) );
  XNOR2_X1 U4494 ( .A(n4112), .B(keyinput_43), .ZN(n3921) );
  XOR2_X1 U4495 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .Z(n3920) );
  OAI21_X1 U4496 ( .B1(n3922), .B2(n3921), .A(n3920), .ZN(n3926) );
  XNOR2_X1 U4497 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_45), .ZN(n3925) );
  XNOR2_X1 U4498 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_46), .ZN(n3924) );
  XNOR2_X1 U4499 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .ZN(n3923) );
  AOI211_X1 U4500 ( .C1(n3926), .C2(n3925), .A(n3924), .B(n3923), .ZN(n3929)
         );
  XOR2_X1 U4501 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .Z(n3928) );
  XNOR2_X1 U4502 ( .A(n4302), .B(keyinput_49), .ZN(n3927) );
  OAI21_X1 U4503 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3932) );
  XNOR2_X1 U4504 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .ZN(n3931) );
  XNOR2_X1 U4505 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_51), .ZN(n3930) );
  AOI21_X1 U4506 ( .B1(n3932), .B2(n3931), .A(n3930), .ZN(n3935) );
  XOR2_X1 U4507 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .Z(n3934) );
  XNOR2_X1 U4508 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .ZN(n3933) );
  NOR3_X1 U4509 ( .A1(n3935), .A2(n3934), .A3(n3933), .ZN(n3943) );
  XNOR2_X1 U4510 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n3942) );
  XOR2_X1 U4511 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .Z(n3940) );
  XNOR2_X1 U4512 ( .A(n3936), .B(keyinput_58), .ZN(n3939) );
  XNOR2_X1 U4513 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .ZN(n3938) );
  XNOR2_X1 U4514 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n3937) );
  NOR4_X1 U4515 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(n3941)
         );
  OAI21_X1 U4516 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3948) );
  XNOR2_X1 U4517 ( .A(n3944), .B(keyinput_59), .ZN(n3947) );
  XNOR2_X1 U4518 ( .A(n4140), .B(keyinput_60), .ZN(n3946) );
  XOR2_X1 U4519 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .Z(n3945) );
  AOI211_X1 U4520 ( .C1(n3948), .C2(n3947), .A(n3946), .B(n3945), .ZN(n3955)
         );
  XNOR2_X1 U4521 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n3954) );
  XNOR2_X1 U4522 ( .A(n3949), .B(keyinput_65), .ZN(n3952) );
  XNOR2_X1 U4523 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n3951) );
  XNOR2_X1 U4524 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n3950) );
  NOR3_X1 U4525 ( .A1(n3952), .A2(n3951), .A3(n3950), .ZN(n3953) );
  OAI21_X1 U4526 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3958) );
  XNOR2_X1 U4527 ( .A(n4151), .B(keyinput_66), .ZN(n3957) );
  XNOR2_X1 U4528 ( .A(n4152), .B(keyinput_67), .ZN(n3956) );
  AOI21_X1 U4529 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3962) );
  XNOR2_X1 U4530 ( .A(n4156), .B(keyinput_68), .ZN(n3961) );
  XNOR2_X1 U4531 ( .A(n3959), .B(keyinput_69), .ZN(n3960) );
  NOR3_X1 U4532 ( .A1(n3962), .A2(n3961), .A3(n3960), .ZN(n3970) );
  XNOR2_X1 U4533 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_72), .ZN(n3969) );
  XNOR2_X1 U4534 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_75), .ZN(n3968) );
  XNOR2_X1 U4535 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .ZN(n3966) );
  XNOR2_X1 U4536 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n3965) );
  XNOR2_X1 U4537 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .ZN(n3964) );
  XNOR2_X1 U4538 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n3963) );
  NAND4_X1 U4539 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  NOR4_X1 U4540 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3973)
         );
  XOR2_X1 U4541 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_76), .Z(n3972) );
  XNOR2_X1 U4542 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n3971) );
  NOR3_X1 U4543 ( .A1(n3973), .A2(n3972), .A3(n3971), .ZN(n3982) );
  XNOR2_X1 U4544 ( .A(n3974), .B(keyinput_78), .ZN(n3981) );
  XOR2_X1 U4545 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .Z(n3979) );
  XNOR2_X1 U4546 ( .A(n4174), .B(keyinput_80), .ZN(n3978) );
  XNOR2_X1 U4547 ( .A(n3975), .B(keyinput_79), .ZN(n3977) );
  XNOR2_X1 U4548 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_82), .ZN(n3976) );
  NOR4_X1 U4549 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  OAI21_X1 U4550 ( .B1(n3982), .B2(n3981), .A(n3980), .ZN(n3986) );
  XNOR2_X1 U4551 ( .A(n3983), .B(keyinput_83), .ZN(n3985) );
  XNOR2_X1 U4552 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .ZN(n3984) );
  NAND3_X1 U4553 ( .A1(n3986), .A2(n3985), .A3(n3984), .ZN(n3990) );
  XOR2_X1 U4554 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .Z(n3989) );
  XNOR2_X1 U4555 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .ZN(n3988) );
  XNOR2_X1 U4556 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_85), .ZN(n3987) );
  NAND4_X1 U4557 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3993)
         );
  XOR2_X1 U4558 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .Z(n3992) );
  XNOR2_X1 U4559 ( .A(D_REG_2__SCAN_IN), .B(keyinput_89), .ZN(n3991) );
  AOI21_X1 U4560 ( .B1(n3993), .B2(n3992), .A(n3991), .ZN(n3996) );
  INV_X1 U4561 ( .A(D_REG_4__SCAN_IN), .ZN(n4928) );
  XNOR2_X1 U4562 ( .A(n4928), .B(keyinput_91), .ZN(n3995) );
  XNOR2_X1 U4563 ( .A(D_REG_3__SCAN_IN), .B(keyinput_90), .ZN(n3994) );
  NOR3_X1 U4564 ( .A1(n3996), .A2(n3995), .A3(n3994), .ZN(n3999) );
  XNOR2_X1 U4565 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n3998) );
  XNOR2_X1 U4566 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .ZN(n3997) );
  OAI21_X1 U4567 ( .B1(n3999), .B2(n3998), .A(n3997), .ZN(n4005) );
  INV_X1 U4568 ( .A(D_REG_7__SCAN_IN), .ZN(n4931) );
  XNOR2_X1 U4569 ( .A(n4931), .B(keyinput_94), .ZN(n4004) );
  XOR2_X1 U4570 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .Z(n4002) );
  INV_X1 U4571 ( .A(D_REG_10__SCAN_IN), .ZN(n4933) );
  XNOR2_X1 U4572 ( .A(n4933), .B(keyinput_97), .ZN(n4001) );
  XNOR2_X1 U4573 ( .A(D_REG_9__SCAN_IN), .B(keyinput_96), .ZN(n4000) );
  NAND3_X1 U4574 ( .A1(n4002), .A2(n4001), .A3(n4000), .ZN(n4003) );
  AOI21_X1 U4575 ( .B1(n4005), .B2(n4004), .A(n4003), .ZN(n4008) );
  INV_X1 U4576 ( .A(D_REG_11__SCAN_IN), .ZN(n4934) );
  XNOR2_X1 U4577 ( .A(n4934), .B(keyinput_98), .ZN(n4007) );
  XNOR2_X1 U4578 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .ZN(n4006) );
  NOR3_X1 U4579 ( .A1(n4008), .A2(n4007), .A3(n4006), .ZN(n4014) );
  INV_X1 U4580 ( .A(D_REG_13__SCAN_IN), .ZN(n4936) );
  XNOR2_X1 U4581 ( .A(n4936), .B(keyinput_100), .ZN(n4013) );
  INV_X1 U4582 ( .A(D_REG_16__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U4583 ( .A(n4939), .B(keyinput_103), .ZN(n4011) );
  INV_X1 U4584 ( .A(D_REG_15__SCAN_IN), .ZN(n4938) );
  XNOR2_X1 U4585 ( .A(n4938), .B(keyinput_102), .ZN(n4010) );
  XNOR2_X1 U4586 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n4009) );
  NOR3_X1 U4587 ( .A1(n4011), .A2(n4010), .A3(n4009), .ZN(n4012) );
  OAI21_X1 U4588 ( .B1(n4014), .B2(n4013), .A(n4012), .ZN(n4017) );
  XNOR2_X1 U4589 ( .A(D_REG_17__SCAN_IN), .B(keyinput_104), .ZN(n4016) );
  INV_X1 U4590 ( .A(D_REG_18__SCAN_IN), .ZN(n4941) );
  XNOR2_X1 U4591 ( .A(n4941), .B(keyinput_105), .ZN(n4015) );
  AOI21_X1 U4592 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4021) );
  INV_X1 U4593 ( .A(D_REG_21__SCAN_IN), .ZN(n4943) );
  XNOR2_X1 U4594 ( .A(n4943), .B(keyinput_108), .ZN(n4020) );
  XNOR2_X1 U4595 ( .A(D_REG_19__SCAN_IN), .B(keyinput_106), .ZN(n4019) );
  XNOR2_X1 U4596 ( .A(D_REG_20__SCAN_IN), .B(keyinput_107), .ZN(n4018) );
  NOR4_X1 U4597 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4025)
         );
  XNOR2_X1 U4598 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4024) );
  XOR2_X1 U4599 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .Z(n4023) );
  XNOR2_X1 U4600 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .ZN(n4022) );
  OAI211_X1 U4601 ( .C1(n4025), .C2(n4024), .A(n4023), .B(n4022), .ZN(n4028)
         );
  XNOR2_X1 U4602 ( .A(D_REG_25__SCAN_IN), .B(keyinput_112), .ZN(n4027) );
  XNOR2_X1 U4603 ( .A(D_REG_26__SCAN_IN), .B(keyinput_113), .ZN(n4026) );
  AOI21_X1 U4604 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(n4034) );
  XNOR2_X1 U4605 ( .A(D_REG_27__SCAN_IN), .B(keyinput_114), .ZN(n4033) );
  INV_X1 U4606 ( .A(D_REG_28__SCAN_IN), .ZN(n4949) );
  XNOR2_X1 U4607 ( .A(n4949), .B(keyinput_115), .ZN(n4031) );
  INV_X1 U4608 ( .A(D_REG_29__SCAN_IN), .ZN(n4950) );
  XNOR2_X1 U4609 ( .A(n4950), .B(keyinput_116), .ZN(n4030) );
  XNOR2_X1 U4610 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n4029) );
  NOR3_X1 U4611 ( .A1(n4031), .A2(n4030), .A3(n4029), .ZN(n4032) );
  OAI21_X1 U4612 ( .B1(n4034), .B2(n4033), .A(n4032), .ZN(n4037) );
  XNOR2_X1 U4613 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n4036) );
  XNOR2_X1 U4614 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .ZN(n4035) );
  NAND3_X1 U4615 ( .A1(n4037), .A2(n4036), .A3(n4035), .ZN(n4043) );
  XOR2_X1 U4616 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .Z(n4042) );
  XOR2_X1 U4617 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .Z(n4040) );
  XNOR2_X1 U4618 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4039) );
  XNOR2_X1 U4619 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4038) );
  NAND3_X1 U4620 ( .A1(n4040), .A2(n4039), .A3(n4038), .ZN(n4041) );
  AOI21_X1 U4621 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4046) );
  XOR2_X1 U4622 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n4045) );
  XNOR2_X1 U4623 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n4044) );
  NOR3_X1 U4624 ( .A1(n4046), .A2(n4045), .A3(n4044), .ZN(n4255) );
  XOR2_X1 U4625 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .Z(n4254) );
  XOR2_X1 U4626 ( .A(DATAI_30_), .B(keyinput_129), .Z(n4050) );
  XOR2_X1 U4627 ( .A(keyinput_128), .B(DATAI_31_), .Z(n4049) );
  XOR2_X1 U4628 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4048) );
  XOR2_X1 U4629 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4047) );
  AOI211_X1 U4630 ( .C1(n4050), .C2(n4049), .A(n4048), .B(n4047), .ZN(n4053)
         );
  XOR2_X1 U4631 ( .A(DATAI_26_), .B(keyinput_133), .Z(n4052) );
  XNOR2_X1 U4632 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n4051) );
  NOR3_X1 U4633 ( .A1(n4053), .A2(n4052), .A3(n4051), .ZN(n4056) );
  XOR2_X1 U4634 ( .A(DATAI_25_), .B(keyinput_134), .Z(n4055) );
  XOR2_X1 U4635 ( .A(DATAI_24_), .B(keyinput_135), .Z(n4054) );
  NOR3_X1 U4636 ( .A1(n4056), .A2(n4055), .A3(n4054), .ZN(n4059) );
  XOR2_X1 U4637 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4058) );
  XOR2_X1 U4638 ( .A(DATAI_22_), .B(keyinput_137), .Z(n4057) );
  OAI21_X1 U4639 ( .B1(n4059), .B2(n4058), .A(n4057), .ZN(n4066) );
  XNOR2_X1 U4640 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n4065) );
  XNOR2_X1 U4641 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n4063) );
  XNOR2_X1 U4642 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4062) );
  XNOR2_X1 U4643 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n4061) );
  XNOR2_X1 U4644 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n4060) );
  NAND4_X1 U4645 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4064)
         );
  AOI21_X1 U4646 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4069) );
  XNOR2_X1 U4647 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n4068) );
  XOR2_X1 U4648 ( .A(DATAI_15_), .B(keyinput_144), .Z(n4067) );
  OAI21_X1 U4649 ( .B1(n4069), .B2(n4068), .A(n4067), .ZN(n4072) );
  XOR2_X1 U4650 ( .A(DATAI_14_), .B(keyinput_145), .Z(n4071) );
  XNOR2_X1 U4651 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n4070) );
  AOI21_X1 U4652 ( .B1(n4072), .B2(n4071), .A(n4070), .ZN(n4076) );
  XNOR2_X1 U4653 ( .A(n4073), .B(keyinput_147), .ZN(n4075) );
  XNOR2_X1 U4654 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n4074) );
  OAI21_X1 U4655 ( .B1(n4076), .B2(n4075), .A(n4074), .ZN(n4079) );
  XNOR2_X1 U4656 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n4078) );
  XOR2_X1 U4657 ( .A(DATAI_9_), .B(keyinput_150), .Z(n4077) );
  AOI21_X1 U4658 ( .B1(n4079), .B2(n4078), .A(n4077), .ZN(n4083) );
  XOR2_X1 U4659 ( .A(DATAI_8_), .B(keyinput_151), .Z(n4082) );
  XOR2_X1 U4660 ( .A(DATAI_7_), .B(keyinput_152), .Z(n4081) );
  XNOR2_X1 U4661 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n4080) );
  OAI211_X1 U4662 ( .C1(n4083), .C2(n4082), .A(n4081), .B(n4080), .ZN(n4086)
         );
  XNOR2_X1 U4663 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n4085) );
  XNOR2_X1 U4664 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n4084) );
  AOI21_X1 U4665 ( .B1(n4086), .B2(n4085), .A(n4084), .ZN(n4088) );
  XNOR2_X1 U4666 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n4087) );
  NOR2_X1 U4667 ( .A1(n4088), .A2(n4087), .ZN(n4096) );
  XNOR2_X1 U4668 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n4092) );
  XNOR2_X1 U4669 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n4091) );
  XNOR2_X1 U4670 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n4090) );
  XNOR2_X1 U4671 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n4089) );
  NAND4_X1 U4672 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4095)
         );
  XNOR2_X1 U4673 ( .A(n4093), .B(keyinput_161), .ZN(n4094) );
  OAI21_X1 U4674 ( .B1(n4096), .B2(n4095), .A(n4094), .ZN(n4099) );
  XNOR2_X1 U4675 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_162), .ZN(n4098) );
  XNOR2_X1 U4676 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .ZN(n4097) );
  AOI21_X1 U4677 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(n4105) );
  XNOR2_X1 U4678 ( .A(n4100), .B(keyinput_164), .ZN(n4104) );
  XOR2_X1 U4679 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .Z(n4103) );
  XNOR2_X1 U4680 ( .A(n4101), .B(keyinput_166), .ZN(n4102) );
  OAI211_X1 U4681 ( .C1(n4105), .C2(n4104), .A(n4103), .B(n4102), .ZN(n4108)
         );
  XNOR2_X1 U4682 ( .A(n4271), .B(keyinput_167), .ZN(n4107) );
  XNOR2_X1 U4683 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n4106) );
  AOI21_X1 U4684 ( .B1(n4108), .B2(n4107), .A(n4106), .ZN(n4111) );
  XOR2_X1 U4685 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .Z(n4110) );
  XNOR2_X1 U4686 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n4109) );
  NOR3_X1 U4687 ( .A1(n4111), .A2(n4110), .A3(n4109), .ZN(n4115) );
  XNOR2_X1 U4688 ( .A(n4112), .B(keyinput_171), .ZN(n4114) );
  XNOR2_X1 U4689 ( .A(keyinput_172), .B(REG3_REG_12__SCAN_IN), .ZN(n4113) );
  OAI21_X1 U4690 ( .B1(n4115), .B2(n4114), .A(n4113), .ZN(n4121) );
  XOR2_X1 U4691 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .Z(n4120) );
  XNOR2_X1 U4692 ( .A(n4116), .B(keyinput_174), .ZN(n4119) );
  XNOR2_X1 U4693 ( .A(n4117), .B(keyinput_175), .ZN(n4118) );
  AOI211_X1 U4694 ( .C1(n4121), .C2(n4120), .A(n4119), .B(n4118), .ZN(n4124)
         );
  XOR2_X1 U4695 ( .A(keyinput_176), .B(REG3_REG_17__SCAN_IN), .Z(n4123) );
  XNOR2_X1 U4696 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n4122) );
  OAI21_X1 U4697 ( .B1(n4124), .B2(n4123), .A(n4122), .ZN(n4128) );
  XNOR2_X1 U4698 ( .A(n4125), .B(keyinput_178), .ZN(n4127) );
  XNOR2_X1 U4699 ( .A(n4313), .B(keyinput_179), .ZN(n4126) );
  AOI21_X1 U4700 ( .B1(n4128), .B2(n4127), .A(n4126), .ZN(n4131) );
  XOR2_X1 U4701 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .Z(n4130) );
  XOR2_X1 U4702 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .Z(n4129) );
  NOR3_X1 U4703 ( .A1(n4131), .A2(n4130), .A3(n4129), .ZN(n4139) );
  INV_X1 U4704 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4997) );
  XNOR2_X1 U4705 ( .A(n4997), .B(keyinput_182), .ZN(n4138) );
  XOR2_X1 U4706 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .Z(n4136) );
  XNOR2_X1 U4707 ( .A(n4132), .B(keyinput_185), .ZN(n4135) );
  XNOR2_X1 U4708 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n4134) );
  XNOR2_X1 U4709 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_186), .ZN(n4133) );
  NOR4_X1 U4710 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4137)
         );
  OAI21_X1 U4711 ( .B1(n4139), .B2(n4138), .A(n4137), .ZN(n4144) );
  XNOR2_X1 U4712 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n4143) );
  XNOR2_X1 U4713 ( .A(n4140), .B(keyinput_188), .ZN(n4142) );
  XNOR2_X1 U4714 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n4141) );
  AOI211_X1 U4715 ( .C1(n4144), .C2(n4143), .A(n4142), .B(n4141), .ZN(n4150)
         );
  XNOR2_X1 U4716 ( .A(n2866), .B(keyinput_190), .ZN(n4149) );
  XNOR2_X1 U4717 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .ZN(n4147) );
  XNOR2_X1 U4718 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .ZN(n4146) );
  XNOR2_X1 U4719 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .ZN(n4145) );
  NOR3_X1 U4720 ( .A1(n4147), .A2(n4146), .A3(n4145), .ZN(n4148) );
  OAI21_X1 U4721 ( .B1(n4150), .B2(n4149), .A(n4148), .ZN(n4155) );
  XNOR2_X1 U4722 ( .A(n4151), .B(keyinput_194), .ZN(n4154) );
  XNOR2_X1 U4723 ( .A(n4152), .B(keyinput_195), .ZN(n4153) );
  AOI21_X1 U4724 ( .B1(n4155), .B2(n4154), .A(n4153), .ZN(n4159) );
  XNOR2_X1 U4725 ( .A(n4156), .B(keyinput_196), .ZN(n4158) );
  XNOR2_X1 U4726 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n4157) );
  NOR3_X1 U4727 ( .A1(n4159), .A2(n4158), .A3(n4157), .ZN(n4169) );
  XNOR2_X1 U4728 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4168) );
  XNOR2_X1 U4729 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .ZN(n4167) );
  XNOR2_X1 U4730 ( .A(n4160), .B(keyinput_201), .ZN(n4165) );
  XNOR2_X1 U4731 ( .A(n4161), .B(keyinput_202), .ZN(n4164) );
  XNOR2_X1 U4732 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_199), .ZN(n4163) );
  XNOR2_X1 U4733 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_203), .ZN(n4162) );
  NAND4_X1 U4734 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4166)
         );
  NOR4_X1 U4735 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4173)
         );
  XNOR2_X1 U4736 ( .A(n4170), .B(keyinput_205), .ZN(n4172) );
  XNOR2_X1 U4737 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4171) );
  NOR3_X1 U4738 ( .A1(n4173), .A2(n4172), .A3(n4171), .ZN(n4181) );
  XNOR2_X1 U4739 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4180) );
  XOR2_X1 U4740 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .Z(n4178) );
  XNOR2_X1 U4741 ( .A(n4174), .B(keyinput_208), .ZN(n4177) );
  XNOR2_X1 U4742 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4176) );
  XNOR2_X1 U4743 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4175) );
  NOR4_X1 U4744 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4179)
         );
  OAI21_X1 U4745 ( .B1(n4181), .B2(n4180), .A(n4179), .ZN(n4184) );
  XNOR2_X1 U4746 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n4183) );
  XNOR2_X1 U4747 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .ZN(n4182) );
  NAND3_X1 U4748 ( .A1(n4184), .A2(n4183), .A3(n4182), .ZN(n4189) );
  INV_X1 U4749 ( .A(keyinput_214), .ZN(n4185) );
  XNOR2_X1 U4750 ( .A(n4185), .B(IR_REG_31__SCAN_IN), .ZN(n4188) );
  XNOR2_X1 U4751 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .ZN(n4187) );
  XNOR2_X1 U4752 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n4186) );
  NAND4_X1 U4753 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4192)
         );
  XOR2_X1 U4754 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .Z(n4191) );
  XNOR2_X1 U4755 ( .A(keyinput_217), .B(D_REG_2__SCAN_IN), .ZN(n4190) );
  AOI21_X1 U4756 ( .B1(n4192), .B2(n4191), .A(n4190), .ZN(n4195) );
  XNOR2_X1 U4757 ( .A(n4928), .B(keyinput_219), .ZN(n4194) );
  XNOR2_X1 U4758 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .ZN(n4193) );
  NOR3_X1 U4759 ( .A1(n4195), .A2(n4194), .A3(n4193), .ZN(n4198) );
  INV_X1 U4760 ( .A(D_REG_5__SCAN_IN), .ZN(n4929) );
  XNOR2_X1 U4761 ( .A(n4929), .B(keyinput_220), .ZN(n4197) );
  INV_X1 U4762 ( .A(D_REG_6__SCAN_IN), .ZN(n4930) );
  XNOR2_X1 U4763 ( .A(n4930), .B(keyinput_221), .ZN(n4196) );
  OAI21_X1 U4764 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(n4204) );
  XNOR2_X1 U4765 ( .A(n4931), .B(keyinput_222), .ZN(n4203) );
  XNOR2_X1 U4766 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .ZN(n4202) );
  XNOR2_X1 U4767 ( .A(keyinput_224), .B(D_REG_9__SCAN_IN), .ZN(n4200) );
  XNOR2_X1 U4768 ( .A(keyinput_225), .B(D_REG_10__SCAN_IN), .ZN(n4199) );
  NAND2_X1 U4769 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  AOI211_X1 U4770 ( .C1(n4204), .C2(n4203), .A(n4202), .B(n4201), .ZN(n4207)
         );
  XNOR2_X1 U4771 ( .A(n4934), .B(keyinput_226), .ZN(n4206) );
  INV_X1 U4772 ( .A(D_REG_12__SCAN_IN), .ZN(n4935) );
  XNOR2_X1 U4773 ( .A(n4935), .B(keyinput_227), .ZN(n4205) );
  NOR3_X1 U4774 ( .A1(n4207), .A2(n4206), .A3(n4205), .ZN(n4213) );
  XNOR2_X1 U4775 ( .A(keyinput_228), .B(D_REG_13__SCAN_IN), .ZN(n4212) );
  XNOR2_X1 U4776 ( .A(n4939), .B(keyinput_231), .ZN(n4210) );
  XNOR2_X1 U4777 ( .A(n4938), .B(keyinput_230), .ZN(n4209) );
  INV_X1 U4778 ( .A(D_REG_14__SCAN_IN), .ZN(n4937) );
  XNOR2_X1 U4779 ( .A(n4937), .B(keyinput_229), .ZN(n4208) );
  NOR3_X1 U4780 ( .A1(n4210), .A2(n4209), .A3(n4208), .ZN(n4211) );
  OAI21_X1 U4781 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n4216) );
  INV_X1 U4782 ( .A(D_REG_17__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U4783 ( .A(n4940), .B(keyinput_232), .ZN(n4215) );
  XNOR2_X1 U4784 ( .A(keyinput_233), .B(D_REG_18__SCAN_IN), .ZN(n4214) );
  AOI21_X1 U4785 ( .B1(n4216), .B2(n4215), .A(n4214), .ZN(n4220) );
  INV_X1 U4786 ( .A(D_REG_19__SCAN_IN), .ZN(n4942) );
  XNOR2_X1 U4787 ( .A(n4942), .B(keyinput_234), .ZN(n4219) );
  XNOR2_X1 U4788 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .ZN(n4218) );
  XNOR2_X1 U4789 ( .A(keyinput_236), .B(D_REG_21__SCAN_IN), .ZN(n4217) );
  NOR4_X1 U4790 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4224)
         );
  XNOR2_X1 U4791 ( .A(keyinput_237), .B(D_REG_22__SCAN_IN), .ZN(n4223) );
  XOR2_X1 U4792 ( .A(D_REG_23__SCAN_IN), .B(keyinput_238), .Z(n4222) );
  XNOR2_X1 U4793 ( .A(keyinput_239), .B(D_REG_24__SCAN_IN), .ZN(n4221) );
  OAI211_X1 U4794 ( .C1(n4224), .C2(n4223), .A(n4222), .B(n4221), .ZN(n4227)
         );
  INV_X1 U4795 ( .A(D_REG_25__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U4796 ( .A(n4946), .B(keyinput_240), .ZN(n4226) );
  XNOR2_X1 U4797 ( .A(keyinput_241), .B(D_REG_26__SCAN_IN), .ZN(n4225) );
  AOI21_X1 U4798 ( .B1(n4227), .B2(n4226), .A(n4225), .ZN(n4233) );
  INV_X1 U4799 ( .A(D_REG_27__SCAN_IN), .ZN(n4948) );
  XNOR2_X1 U4800 ( .A(n4948), .B(keyinput_242), .ZN(n4232) );
  XNOR2_X1 U4801 ( .A(n4950), .B(keyinput_244), .ZN(n4230) );
  XNOR2_X1 U4802 ( .A(n4949), .B(keyinput_243), .ZN(n4229) );
  XNOR2_X1 U4803 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n4228) );
  NOR3_X1 U4804 ( .A1(n4230), .A2(n4229), .A3(n4228), .ZN(n4231) );
  OAI21_X1 U4805 ( .B1(n4233), .B2(n4232), .A(n4231), .ZN(n4236) );
  XNOR2_X1 U4806 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .ZN(n4235) );
  XNOR2_X1 U4807 ( .A(keyinput_246), .B(D_REG_31__SCAN_IN), .ZN(n4234) );
  NAND3_X1 U4808 ( .A1(n4236), .A2(n4235), .A3(n4234), .ZN(n4242) );
  XOR2_X1 U4809 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .Z(n4241) );
  XNOR2_X1 U4810 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .ZN(n4239) );
  XNOR2_X1 U4811 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .ZN(n4238) );
  XNOR2_X1 U4812 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .ZN(n4237) );
  NAND3_X1 U4813 ( .A1(n4239), .A2(n4238), .A3(n4237), .ZN(n4240) );
  AOI21_X1 U4814 ( .B1(n4242), .B2(n4241), .A(n4240), .ZN(n4245) );
  XOR2_X1 U4815 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .Z(n4244) );
  XOR2_X1 U4816 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .Z(n4243) );
  NOR3_X1 U4817 ( .A1(n4245), .A2(n4244), .A3(n4243), .ZN(n4247) );
  XOR2_X1 U4818 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4246) );
  NOR2_X1 U4819 ( .A1(n4247), .A2(n4246), .ZN(n4248) );
  NOR2_X1 U4820 ( .A1(n4248), .A2(keyinput_255), .ZN(n4251) );
  OAI21_X1 U4821 ( .B1(n4251), .B2(n4248), .A(keyinput_127), .ZN(n4249) );
  NAND2_X1 U4822 ( .A1(n4249), .A2(REG0_REG_8__SCAN_IN), .ZN(n4253) );
  INV_X1 U4823 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4250) );
  OAI21_X1 U4824 ( .B1(n4251), .B2(keyinput_127), .A(n4250), .ZN(n4252) );
  OAI211_X1 U4825 ( .C1(n4255), .C2(n4254), .A(n4253), .B(n4252), .ZN(n4256)
         );
  XNOR2_X1 U4826 ( .A(n4257), .B(n4256), .ZN(U3217) );
  XNOR2_X1 U4827 ( .A(n4258), .B(n4259), .ZN(n4265) );
  NAND2_X1 U4828 ( .A1(n4523), .A2(n5265), .ZN(n4262) );
  AOI22_X1 U4829 ( .A1(n5263), .A2(n4260), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4261) );
  OAI211_X1 U4830 ( .C1(n5279), .C2(n4694), .A(n4262), .B(n4261), .ZN(n4263)
         );
  AOI21_X1 U4831 ( .B1(n4358), .B2(n4521), .A(n4263), .ZN(n4264) );
  OAI21_X1 U4832 ( .B1(n4265), .B2(n4363), .A(n4264), .ZN(U3211) );
  OAI21_X1 U4833 ( .B1(n4268), .B2(n4267), .A(n4266), .ZN(n4275) );
  INV_X1 U4834 ( .A(n4269), .ZN(n4821) );
  AOI22_X1 U4835 ( .A1(n4358), .A2(n4810), .B1(n5263), .B2(n4270), .ZN(n4273)
         );
  NOR2_X1 U4836 ( .A1(STATE_REG_SCAN_IN), .A2(n4271), .ZN(n4658) );
  AOI21_X1 U4837 ( .B1(n5265), .B2(n4811), .A(n4658), .ZN(n4272) );
  OAI211_X1 U4838 ( .C1(n4821), .C2(n5279), .A(n4273), .B(n4272), .ZN(n4274)
         );
  AOI21_X1 U4839 ( .B1(n4275), .B2(n5274), .A(n4274), .ZN(n4276) );
  INV_X1 U4840 ( .A(n4276), .ZN(U3216) );
  INV_X1 U4841 ( .A(n4349), .ZN(n4277) );
  NAND2_X1 U4842 ( .A1(n4277), .A2(n4351), .ZN(n4278) );
  XNOR2_X1 U4843 ( .A(n4350), .B(n4278), .ZN(n4285) );
  INV_X1 U4844 ( .A(n5265), .ZN(n4326) );
  AOI22_X1 U4845 ( .A1(n5263), .A2(n4279), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n4282) );
  NAND2_X1 U4846 ( .A1(n4280), .A2(n4317), .ZN(n4281) );
  OAI211_X1 U4847 ( .C1(n4407), .C2(n4326), .A(n4282), .B(n4281), .ZN(n4283)
         );
  AOI21_X1 U4848 ( .B1(n4523), .B2(n4358), .A(n4283), .ZN(n4284) );
  OAI21_X1 U4849 ( .B1(n4285), .B2(n4363), .A(n4284), .ZN(U3222) );
  AND3_X1 U4850 ( .A1(n3730), .A2(n4288), .A3(n4287), .ZN(n4289) );
  OAI21_X1 U4851 ( .B1(n4286), .B2(n4289), .A(n5274), .ZN(n4294) );
  NAND2_X1 U4852 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n5030) );
  OAI21_X1 U4853 ( .B1(n4290), .B2(n4345), .A(n5030), .ZN(n4291) );
  AOI21_X1 U4854 ( .B1(n4292), .B2(n5263), .A(n4291), .ZN(n4293) );
  OAI211_X1 U4855 ( .C1(n4295), .C2(n5279), .A(n4294), .B(n4293), .ZN(U3225)
         );
  INV_X1 U4856 ( .A(n4296), .ZN(n4299) );
  INV_X1 U4857 ( .A(n4297), .ZN(n4298) );
  NOR2_X1 U4858 ( .A1(n4299), .A2(n4298), .ZN(n4301) );
  XNOR2_X1 U4859 ( .A(n4301), .B(n4300), .ZN(n4306) );
  OAI22_X1 U4860 ( .A1(n4324), .A2(n4728), .B1(STATE_REG_SCAN_IN), .B2(n4302), 
        .ZN(n4304) );
  INV_X1 U4861 ( .A(n4763), .ZN(n4720) );
  OAI22_X1 U4862 ( .A1(n4720), .A2(n4326), .B1(n4731), .B2(n5279), .ZN(n4303)
         );
  AOI211_X1 U4863 ( .C1(n4358), .C2(n4726), .A(n4304), .B(n4303), .ZN(n4305)
         );
  OAI21_X1 U4864 ( .B1(n4306), .B2(n4363), .A(n4305), .ZN(U3226) );
  NAND2_X1 U4865 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  OAI21_X1 U4866 ( .B1(n4310), .B2(n4309), .A(n3789), .ZN(n4311) );
  NAND2_X1 U4867 ( .A1(n4311), .A2(n5274), .ZN(n4320) );
  AOI22_X1 U4868 ( .A1(n4533), .A2(n4358), .B1(n4312), .B2(n5263), .ZN(n4319)
         );
  NOR2_X1 U4869 ( .A1(STATE_REG_SCAN_IN), .A2(n4313), .ZN(n4995) );
  NOR2_X1 U4870 ( .A1(n4326), .A2(n4314), .ZN(n4315) );
  AOI211_X1 U4871 ( .C1(n4317), .C2(n4316), .A(n4995), .B(n4315), .ZN(n4318)
         );
  NAND3_X1 U4872 ( .A1(n4320), .A2(n4319), .A3(n4318), .ZN(U3228) );
  AOI21_X1 U4873 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4330) );
  OAI22_X1 U4874 ( .A1(n4324), .A2(n4765), .B1(n5279), .B2(n4768), .ZN(n4328)
         );
  INV_X1 U4875 ( .A(n4526), .ZN(n5271) );
  OAI22_X1 U4876 ( .A1(n4326), .A2(n5271), .B1(STATE_REG_SCAN_IN), .B2(n4325), 
        .ZN(n4327) );
  AOI211_X1 U4877 ( .C1(n4358), .C2(n4763), .A(n4328), .B(n4327), .ZN(n4329)
         );
  OAI21_X1 U4878 ( .B1(n4330), .B2(n4363), .A(n4329), .ZN(U3232) );
  OAI21_X1 U4879 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(n4334) );
  NAND2_X1 U4880 ( .A1(n4334), .A2(n5274), .ZN(n4339) );
  AOI22_X1 U4881 ( .A1(n4358), .A2(n4540), .B1(n5265), .B2(n3023), .ZN(n4338)
         );
  AOI22_X1 U4882 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4336), .B1(n5263), .B2(n4335), .ZN(n4337) );
  NAND3_X1 U4883 ( .A1(n4339), .A2(n4338), .A3(n4337), .ZN(U3234) );
  INV_X1 U4884 ( .A(n4340), .ZN(n4344) );
  NOR3_X1 U4885 ( .A1(n4286), .A2(n4342), .A3(n4341), .ZN(n4343) );
  OAI21_X1 U4886 ( .B1(n4344), .B2(n4343), .A(n5274), .ZN(n4348) );
  AOI22_X1 U4887 ( .A1(n5204), .A2(n4527), .B1(n5264), .B2(n4809), .ZN(n4831)
         );
  NAND2_X1 U4888 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4646) );
  OAI21_X1 U4889 ( .B1(n4831), .B2(n4345), .A(n4646), .ZN(n4346) );
  AOI21_X1 U4890 ( .B1(n4839), .B2(n5263), .A(n4346), .ZN(n4347) );
  OAI211_X1 U4891 ( .C1(n4840), .C2(n5279), .A(n4348), .B(n4347), .ZN(U3235)
         );
  NAND2_X1 U4892 ( .A1(n4352), .A2(n4351), .ZN(n4356) );
  XOR2_X1 U4893 ( .A(n4354), .B(n4353), .Z(n4355) );
  XNOR2_X1 U4894 ( .A(n4356), .B(n4355), .ZN(n4364) );
  INV_X1 U4895 ( .A(n4357), .ZN(n4705) );
  NAND2_X1 U4896 ( .A1(n4522), .A2(n4358), .ZN(n4360) );
  AOI22_X1 U4897 ( .A1(n5263), .A2(n4703), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4359) );
  OAI211_X1 U4898 ( .C1(n5279), .C2(n4705), .A(n4360), .B(n4359), .ZN(n4361)
         );
  AOI21_X1 U4899 ( .B1(n5265), .B2(n4726), .A(n4361), .ZN(n4362) );
  OAI21_X1 U4900 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(U3237) );
  INV_X1 U4901 ( .A(n4835), .ZN(n4829) );
  NAND4_X1 U4902 ( .A1(n4829), .A2(n4367), .A3(n4366), .A4(n4365), .ZN(n4383)
         );
  NAND4_X1 U4903 ( .A1(n4371), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(n4382)
         );
  NAND2_X1 U4904 ( .A1(n3130), .A2(REG1_REG_30__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U4905 ( .A1(n2940), .A2(REG2_REG_30__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U4906 ( .A1(n4375), .A2(REG0_REG_30__SCAN_IN), .ZN(n4372) );
  NAND3_X1 U4907 ( .A1(n4374), .A2(n4373), .A3(n4372), .ZN(n4676) );
  NAND2_X1 U4908 ( .A1(n4404), .A2(DATAI_30_), .ZN(n5296) );
  OR2_X1 U4909 ( .A1(n4676), .A2(n5296), .ZN(n4379) );
  NAND2_X1 U4910 ( .A1(n3130), .A2(REG1_REG_31__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U4911 ( .A1(n2940), .A2(REG2_REG_31__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U4912 ( .A1(n4375), .A2(REG0_REG_31__SCAN_IN), .ZN(n4376) );
  NAND3_X1 U4913 ( .A1(n4378), .A2(n4377), .A3(n4376), .ZN(n5281) );
  NAND2_X1 U4914 ( .A1(n4404), .A2(DATAI_31_), .ZN(n5298) );
  NAND2_X1 U4915 ( .A1(n5281), .A2(n5298), .ZN(n4472) );
  AND2_X1 U4916 ( .A1(n4379), .A2(n4472), .ZN(n4474) );
  INV_X1 U4917 ( .A(n4474), .ZN(n4380) );
  OR4_X1 U4918 ( .A1(n5149), .A2(n4380), .A3(n4817), .A4(n4916), .ZN(n4381) );
  NOR4_X1 U4919 ( .A1(n4383), .A2(n4382), .A3(n4381), .A4(n4777), .ZN(n4386)
         );
  XNOR2_X1 U4920 ( .A(n3039), .B(n4384), .ZN(n5060) );
  NAND3_X1 U4921 ( .A1(n4386), .A2(n4385), .A3(n5060), .ZN(n4399) );
  INV_X1 U4922 ( .A(n4387), .ZN(n4390) );
  AND4_X1 U4923 ( .A1(n4390), .A2(n2540), .A3(n4389), .A4(n4388), .ZN(n4394)
         );
  INV_X1 U4924 ( .A(n4793), .ZN(n4393) );
  NAND4_X1 U4925 ( .A1(n4394), .A2(n4393), .A3(n4392), .A4(n4391), .ZN(n4397)
         );
  NAND2_X1 U4926 ( .A1(n2537), .A2(n4395), .ZN(n4741) );
  XNOR2_X1 U4927 ( .A(n4531), .B(n5182), .ZN(n5198) );
  NAND3_X1 U4928 ( .A1(n4741), .A2(n4756), .A3(n5198), .ZN(n4396) );
  NOR4_X1 U4929 ( .A1(n4399), .A2(n4398), .A3(n4397), .A4(n4396), .ZN(n4403)
         );
  INV_X1 U4930 ( .A(n4465), .ZN(n4401) );
  NAND2_X1 U4931 ( .A1(n4401), .A2(n4400), .ZN(n4709) );
  INV_X1 U4932 ( .A(n4709), .ZN(n4402) );
  NAND3_X1 U4933 ( .A1(n4403), .A2(n4688), .A3(n4402), .ZN(n4409) );
  AND2_X1 U4934 ( .A1(n4404), .A2(DATAI_29_), .ZN(n4675) );
  NAND2_X1 U4935 ( .A1(n4405), .A2(n4675), .ZN(n4475) );
  INV_X1 U4936 ( .A(n4675), .ZN(n4406) );
  NAND2_X1 U4937 ( .A1(n4520), .A2(n4406), .ZN(n4463) );
  INV_X1 U4938 ( .A(n4664), .ZN(n4671) );
  XNOR2_X1 U4939 ( .A(n4407), .B(n4728), .ZN(n4718) );
  INV_X1 U4940 ( .A(n4718), .ZN(n4721) );
  NOR4_X1 U4941 ( .A1(n4409), .A2(n4671), .A3(n4408), .A4(n4721), .ZN(n4410)
         );
  NAND2_X1 U4942 ( .A1(n4410), .A2(n4662), .ZN(n4469) );
  NAND2_X1 U4943 ( .A1(n4412), .A2(n4411), .ZN(n4488) );
  INV_X1 U4944 ( .A(n4449), .ZN(n4413) );
  NAND2_X1 U4945 ( .A1(n4421), .A2(n4413), .ZN(n4414) );
  NAND2_X1 U4946 ( .A1(n4414), .A2(n4448), .ZN(n4479) );
  INV_X1 U4947 ( .A(n4415), .ZN(n4418) );
  AND2_X1 U4948 ( .A1(n4417), .A2(n4416), .ZN(n4442) );
  NAND4_X1 U4949 ( .A1(n4418), .A2(n4442), .A3(n4441), .A4(n4439), .ZN(n4420)
         );
  NAND2_X1 U4950 ( .A1(n4420), .A2(n4419), .ZN(n4425) );
  NAND2_X1 U4951 ( .A1(n4422), .A2(n4421), .ZN(n4481) );
  INV_X1 U4952 ( .A(n4423), .ZN(n4424) );
  AOI211_X1 U4953 ( .C1(n4450), .C2(n4425), .A(n4481), .B(n4424), .ZN(n4453)
         );
  AOI21_X1 U4954 ( .B1(n3039), .B2(n5057), .A(n4426), .ZN(n4427) );
  OAI21_X1 U4955 ( .B1(n5058), .B2(n2838), .A(n4427), .ZN(n4429) );
  NAND2_X1 U4956 ( .A1(n4429), .A2(n4428), .ZN(n4432) );
  OAI211_X1 U4957 ( .C1(n4433), .C2(n4432), .A(n4431), .B(n4430), .ZN(n4436)
         );
  NAND3_X1 U4958 ( .A1(n4436), .A2(n4435), .A3(n4434), .ZN(n4440) );
  NAND2_X1 U4959 ( .A1(n4438), .A2(n4437), .ZN(n4444) );
  AOI21_X1 U4960 ( .B1(n4440), .B2(n4439), .A(n4444), .ZN(n4447) );
  OAI211_X1 U4961 ( .C1(n4444), .C2(n4443), .A(n4442), .B(n4441), .ZN(n4446)
         );
  OAI21_X1 U4962 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n4451) );
  NAND4_X1 U4963 ( .A1(n4451), .A2(n4450), .A3(n4449), .A4(n4448), .ZN(n4452)
         );
  OAI211_X1 U4964 ( .C1(n4479), .C2(n4453), .A(n4485), .B(n4452), .ZN(n4454)
         );
  OAI221_X1 U4965 ( .B1(n4488), .B2(n4483), .C1(n4488), .C2(n4454), .A(n4487), 
        .ZN(n4455) );
  OAI21_X1 U4966 ( .B1(n4757), .B2(n4455), .A(n4493), .ZN(n4458) );
  NAND2_X1 U4967 ( .A1(n4457), .A2(n4456), .ZN(n4490) );
  AOI21_X1 U4968 ( .B1(n4459), .B2(n4458), .A(n4490), .ZN(n4460) );
  INV_X1 U4969 ( .A(n4460), .ZN(n4467) );
  AND2_X1 U4970 ( .A1(n4462), .A2(n4461), .ZN(n4498) );
  NAND2_X1 U4971 ( .A1(n4521), .A2(n4661), .ZN(n4669) );
  AND2_X1 U4972 ( .A1(n4669), .A2(n4463), .ZN(n4476) );
  INV_X1 U4973 ( .A(n4476), .ZN(n4466) );
  NOR3_X1 U4974 ( .A1(n4466), .A2(n4465), .A3(n4464), .ZN(n4501) );
  OAI221_X1 U4975 ( .B1(n4467), .B2(n4495), .C1(n4498), .C2(n4495), .A(n4501), 
        .ZN(n4468) );
  MUX2_X1 U4976 ( .A(n4469), .B(n4468), .S(n2517), .Z(n4511) );
  INV_X1 U4977 ( .A(n5281), .ZN(n4471) );
  INV_X1 U4978 ( .A(n5298), .ZN(n4470) );
  AOI22_X1 U4979 ( .A1(n4471), .A2(n4470), .B1(n4676), .B2(n5296), .ZN(n4506)
         );
  INV_X1 U4980 ( .A(n4506), .ZN(n4510) );
  INV_X1 U4981 ( .A(n4472), .ZN(n4478) );
  OAI21_X1 U4982 ( .B1(n4521), .B2(n4661), .A(n4473), .ZN(n4496) );
  NAND2_X1 U4983 ( .A1(n4475), .A2(n4474), .ZN(n4502) );
  AOI21_X1 U4984 ( .B1(n4496), .B2(n4476), .A(n4502), .ZN(n4477) );
  INV_X1 U4985 ( .A(n4477), .ZN(n4500) );
  OAI21_X1 U4986 ( .B1(n4506), .B2(n4478), .A(n4500), .ZN(n4508) );
  INV_X1 U4987 ( .A(n4479), .ZN(n4480) );
  OAI21_X1 U4988 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n4486) );
  INV_X1 U4989 ( .A(n4483), .ZN(n4484) );
  AOI21_X1 U4990 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4489) );
  OAI21_X1 U4991 ( .B1(n4489), .B2(n4488), .A(n4487), .ZN(n4492) );
  INV_X1 U4992 ( .A(n4490), .ZN(n4491) );
  OAI221_X1 U4993 ( .B1(n4494), .B2(n4493), .C1(n4494), .C2(n4492), .A(n4491), 
        .ZN(n4497) );
  AOI211_X1 U4994 ( .C1(n4498), .C2(n4497), .A(n4496), .B(n4495), .ZN(n4499)
         );
  INV_X1 U4995 ( .A(n4499), .ZN(n4503) );
  OAI22_X1 U4996 ( .A1(n4503), .A2(n4502), .B1(n4501), .B2(n4500), .ZN(n4504)
         );
  OAI21_X1 U4997 ( .B1(n5296), .B2(n5281), .A(n4504), .ZN(n4505) );
  OAI211_X1 U4998 ( .C1(n4506), .C2(n5298), .A(n4505), .B(n4916), .ZN(n4507)
         );
  MUX2_X1 U4999 ( .A(n4508), .B(n4507), .S(n4849), .Z(n4509) );
  OAI21_X1 U5000 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n4512) );
  XNOR2_X1 U5001 ( .A(n4512), .B(n4848), .ZN(n4518) );
  INV_X1 U5002 ( .A(B_REG_SCAN_IN), .ZN(n4513) );
  AOI21_X1 U5003 ( .B1(n4517), .B2(n4514), .A(n4513), .ZN(n4516) );
  NAND3_X1 U5004 ( .A1(n4859), .A2(n4911), .A3(n5204), .ZN(n4515) );
  AOI22_X1 U5005 ( .A1(n4518), .A2(n4517), .B1(n4516), .B2(n4515), .ZN(n4519)
         );
  INV_X1 U5006 ( .A(n4519), .ZN(U3239) );
  MUX2_X1 U5007 ( .A(DATAO_REG_31__SCAN_IN), .B(n5281), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U5008 ( .A(DATAO_REG_30__SCAN_IN), .B(n4676), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U5009 ( .A(DATAO_REG_29__SCAN_IN), .B(n4520), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U5010 ( .A(DATAO_REG_28__SCAN_IN), .B(n4521), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U5011 ( .A(DATAO_REG_27__SCAN_IN), .B(n4522), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U5012 ( .A(DATAO_REG_26__SCAN_IN), .B(n4523), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U5013 ( .A(DATAO_REG_25__SCAN_IN), .B(n4726), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U5014 ( .A(DATAO_REG_24__SCAN_IN), .B(n4524), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U5015 ( .A(DATAO_REG_23__SCAN_IN), .B(n4763), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U5016 ( .A(DATAO_REG_22__SCAN_IN), .B(n4525), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U5017 ( .A(DATAO_REG_21__SCAN_IN), .B(n4526), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U5018 ( .A(DATAO_REG_20__SCAN_IN), .B(n4810), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U5019 ( .A(DATAO_REG_19__SCAN_IN), .B(n5264), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U5020 ( .A(DATAO_REG_18__SCAN_IN), .B(n4811), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U5021 ( .A(DATAO_REG_17__SCAN_IN), .B(n4527), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U5022 ( .A(DATAO_REG_16__SCAN_IN), .B(n4528), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U5023 ( .A(DATAO_REG_15__SCAN_IN), .B(n4529), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U5024 ( .A(DATAO_REG_14__SCAN_IN), .B(n4530), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U5025 ( .A(DATAO_REG_13__SCAN_IN), .B(n4531), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U5026 ( .A(DATAO_REG_12__SCAN_IN), .B(n5203), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U5027 ( .A(DATAO_REG_11__SCAN_IN), .B(n4532), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U5028 ( .A(DATAO_REG_10__SCAN_IN), .B(n4533), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U5029 ( .A(DATAO_REG_9__SCAN_IN), .B(n4534), .S(U4043), .Z(U3559) );
  MUX2_X1 U5030 ( .A(DATAO_REG_8__SCAN_IN), .B(n4535), .S(U4043), .Z(U3558) );
  MUX2_X1 U5031 ( .A(DATAO_REG_7__SCAN_IN), .B(n4536), .S(U4043), .Z(U3557) );
  MUX2_X1 U5032 ( .A(DATAO_REG_6__SCAN_IN), .B(n4537), .S(U4043), .Z(U3556) );
  MUX2_X1 U5033 ( .A(DATAO_REG_5__SCAN_IN), .B(n4538), .S(U4043), .Z(U3555) );
  MUX2_X1 U5034 ( .A(DATAO_REG_4__SCAN_IN), .B(n4539), .S(U4043), .Z(U3554) );
  MUX2_X1 U5035 ( .A(DATAO_REG_3__SCAN_IN), .B(n4540), .S(U4043), .Z(U3553) );
  MUX2_X1 U5036 ( .A(DATAO_REG_2__SCAN_IN), .B(n3025), .S(U4043), .Z(U3552) );
  MUX2_X1 U5037 ( .A(DATAO_REG_1__SCAN_IN), .B(n3023), .S(U4043), .Z(U3551) );
  MUX2_X1 U5038 ( .A(DATAO_REG_0__SCAN_IN), .B(n3039), .S(U4043), .Z(U3550) );
  NAND2_X1 U5039 ( .A1(n5046), .A2(n4926), .ZN(n4550) );
  INV_X1 U5040 ( .A(IR_REG_0__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5041 ( .A1(n4543), .A2(n5070), .ZN(n4552) );
  OAI211_X1 U5042 ( .C1(n4552), .C2(n4542), .A(n5043), .B(n4541), .ZN(n4549)
         );
  INV_X1 U5043 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U5044 ( .A1(n4543), .A2(n5061), .ZN(n4546) );
  OAI211_X1 U5045 ( .C1(n4546), .C2(n4545), .A(n5033), .B(n4544), .ZN(n4548)
         );
  AOI22_X1 U5046 ( .A1(n5053), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4547) );
  NAND4_X1 U5047 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n4547), .ZN(U3241)
         );
  MUX2_X1 U5048 ( .A(n4552), .B(n4551), .S(n2772), .Z(n4554) );
  NAND2_X1 U5049 ( .A1(n4554), .A2(n4553), .ZN(n4556) );
  OAI211_X1 U5050 ( .C1(IR_REG_0__SCAN_IN), .C2(n4557), .A(n4556), .B(U4043), 
        .ZN(n5054) );
  AOI22_X1 U5051 ( .A1(n5053), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4560) );
  OR2_X1 U5052 ( .A1(n5009), .A2(n4558), .ZN(n4559) );
  AND2_X1 U5053 ( .A1(n4560), .A2(n4559), .ZN(n4569) );
  OAI211_X1 U5054 ( .C1(n4563), .C2(n4562), .A(n5043), .B(n4561), .ZN(n4568)
         );
  OAI211_X1 U5055 ( .C1(n4566), .C2(n4565), .A(n5033), .B(n4564), .ZN(n4567)
         );
  NAND4_X1 U5056 ( .A1(n5054), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(U3242)
         );
  NAND2_X1 U5057 ( .A1(n5046), .A2(n4924), .ZN(n4581) );
  OAI211_X1 U5058 ( .C1(n4572), .C2(n4571), .A(n5043), .B(n4570), .ZN(n4580)
         );
  OAI211_X1 U5059 ( .C1(n4575), .C2(n4574), .A(n5033), .B(n4573), .ZN(n4579)
         );
  INV_X1 U5060 ( .A(n4576), .ZN(n4577) );
  AOI21_X1 U5061 ( .B1(n5053), .B2(ADDR_REG_5__SCAN_IN), .A(n4577), .ZN(n4578)
         );
  NAND4_X1 U5062 ( .A1(n4581), .A2(n4580), .A3(n4579), .A4(n4578), .ZN(U3245)
         );
  INV_X1 U5063 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4582) );
  MUX2_X1 U5064 ( .A(REG1_REG_7__SCAN_IN), .B(n4582), .S(n4923), .Z(n4584) );
  OAI211_X1 U5065 ( .C1(n4585), .C2(n4584), .A(n4583), .B(n5033), .ZN(n4595)
         );
  INV_X1 U5066 ( .A(n4586), .ZN(n4587) );
  AOI21_X1 U5067 ( .B1(n5053), .B2(ADDR_REG_7__SCAN_IN), .A(n4587), .ZN(n4594)
         );
  OAI211_X1 U5068 ( .C1(n4590), .C2(n4589), .A(n5043), .B(n4588), .ZN(n4593)
         );
  INV_X1 U5069 ( .A(n4923), .ZN(n4591) );
  OR2_X1 U5070 ( .A1(n5009), .A2(n4591), .ZN(n4592) );
  NAND4_X1 U5071 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(U3247)
         );
  INV_X1 U5072 ( .A(n4596), .ZN(n4607) );
  NOR2_X1 U5073 ( .A1(n4998), .A2(REG1_REG_13__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U5074 ( .A1(n4998), .A2(REG1_REG_13__SCAN_IN), .ZN(n4601) );
  INV_X1 U5075 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5240) );
  MUX2_X1 U5076 ( .A(n5240), .B(REG1_REG_15__SCAN_IN), .S(n4920), .Z(n4603) );
  NOR2_X1 U5077 ( .A1(n4920), .A2(REG1_REG_15__SCAN_IN), .ZN(n4602) );
  AOI211_X1 U5078 ( .C1(n4604), .C2(n4603), .A(n5049), .B(n4622), .ZN(n4621)
         );
  INV_X1 U5079 ( .A(n4920), .ZN(n4619) );
  NOR2_X1 U5080 ( .A1(n4998), .A2(REG2_REG_13__SCAN_IN), .ZN(n4605) );
  AOI21_X1 U5081 ( .B1(REG2_REG_13__SCAN_IN), .B2(n4998), .A(n4605), .ZN(n5004) );
  NAND2_X1 U5082 ( .A1(n4607), .A2(n4606), .ZN(n4609) );
  NAND2_X1 U5083 ( .A1(n5004), .A2(n5005), .ZN(n5003) );
  NAND2_X1 U5084 ( .A1(n2620), .A2(n5016), .ZN(n4610) );
  NAND2_X1 U5085 ( .A1(n4619), .A2(n4611), .ZN(n4612) );
  NAND2_X1 U5086 ( .A1(n4920), .A2(REG2_REG_15__SCAN_IN), .ZN(n4625) );
  AND2_X1 U5087 ( .A1(n4612), .A2(n4625), .ZN(n4613) );
  NAND2_X1 U5088 ( .A1(n4613), .A2(n4614), .ZN(n4624) );
  OAI211_X1 U5089 ( .C1(n4614), .C2(n4613), .A(n4624), .B(n5043), .ZN(n4618)
         );
  INV_X1 U5090 ( .A(n4615), .ZN(n4616) );
  AOI21_X1 U5091 ( .B1(n5053), .B2(ADDR_REG_15__SCAN_IN), .A(n4616), .ZN(n4617) );
  OAI211_X1 U5092 ( .C1(n5009), .C2(n4619), .A(n4618), .B(n4617), .ZN(n4620)
         );
  OR2_X1 U5093 ( .A1(n4621), .A2(n4620), .ZN(U3255) );
  INV_X1 U5094 ( .A(n4919), .ZN(n4642) );
  AOI21_X1 U5095 ( .B1(n4623), .B2(REG1_REG_16__SCAN_IN), .A(n4635), .ZN(n4633) );
  AND2_X1 U5096 ( .A1(n4626), .A2(REG2_REG_16__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5097 ( .B1(n4640), .B2(n4627), .A(n5043), .ZN(n4630) );
  AOI21_X1 U5098 ( .B1(n5053), .B2(ADDR_REG_16__SCAN_IN), .A(n4628), .ZN(n4629) );
  OAI211_X1 U5099 ( .C1(n4642), .C2(n5009), .A(n4630), .B(n4629), .ZN(n4631)
         );
  INV_X1 U5100 ( .A(n4631), .ZN(n4632) );
  OAI21_X1 U5101 ( .B1(n4633), .B2(n5049), .A(n4632), .ZN(U3256) );
  NOR2_X1 U5102 ( .A1(n5039), .A2(n5252), .ZN(n4636) );
  INV_X1 U5103 ( .A(REG1_REG_17__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U5104 ( .A1(n5039), .A2(n5252), .ZN(n5035) );
  INV_X1 U5105 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U5106 ( .A1(n4917), .A2(n5259), .ZN(n4637) );
  AOI21_X1 U5107 ( .B1(n4917), .B2(n5259), .A(n4637), .ZN(n4638) );
  INV_X1 U5108 ( .A(n4639), .ZN(n4641) );
  NAND2_X1 U5109 ( .A1(n3557), .A2(n5039), .ZN(n5028) );
  OAI221_X1 U5110 ( .B1(n5029), .B2(n4918), .C1(n5029), .C2(
        REG2_REG_17__SCAN_IN), .A(n5028), .ZN(n5027) );
  NAND2_X1 U5111 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4917), .ZN(n4643) );
  OAI21_X1 U5112 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4917), .A(n4643), .ZN(n4644) );
  NOR2_X1 U5113 ( .A1(n5027), .A2(n4644), .ZN(n4651) );
  INV_X1 U5114 ( .A(n5043), .ZN(n5024) );
  AOI211_X1 U5115 ( .C1(n5027), .C2(n4644), .A(n4651), .B(n5024), .ZN(n4649)
         );
  NAND2_X1 U5116 ( .A1(n5053), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4645) );
  OAI211_X1 U5117 ( .C1(n5009), .C2(n4647), .A(n4646), .B(n4645), .ZN(n4648)
         );
  INV_X1 U5118 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4650) );
  MUX2_X1 U5119 ( .A(n4650), .B(REG2_REG_19__SCAN_IN), .S(n4848), .Z(n4653) );
  AOI21_X1 U5120 ( .B1(n4917), .B2(REG2_REG_18__SCAN_IN), .A(n4651), .ZN(n4652) );
  XNOR2_X1 U5121 ( .A(n4653), .B(n4652), .ZN(n4657) );
  XNOR2_X1 U5122 ( .A(n4848), .B(REG1_REG_19__SCAN_IN), .ZN(n4655) );
  XNOR2_X1 U5123 ( .A(n4655), .B(n4654), .ZN(n4656) );
  AOI22_X1 U5124 ( .A1(n5043), .A2(n4657), .B1(n5033), .B2(n4656), .ZN(n4660)
         );
  AOI21_X1 U5125 ( .B1(n5053), .B2(ADDR_REG_19__SCAN_IN), .A(n4658), .ZN(n4659) );
  OAI211_X1 U5126 ( .C1(n4848), .C2(n5009), .A(n4660), .B(n4659), .ZN(U3259)
         );
  OAI22_X1 U5127 ( .A1(n4663), .A2(n4662), .B1(n4683), .B2(n4661), .ZN(n4665)
         );
  XNOR2_X1 U5128 ( .A(n4665), .B(n4664), .ZN(n4850) );
  INV_X1 U5129 ( .A(n4850), .ZN(n4680) );
  AOI211_X1 U5130 ( .C1(n4675), .C2(n2523), .A(n5229), .B(n5297), .ZN(n4852)
         );
  INV_X1 U5131 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4666) );
  OAI22_X1 U5132 ( .A1(n4667), .A2(n5216), .B1(n4666), .B2(n5173), .ZN(n4668)
         );
  AOI21_X1 U5133 ( .B1(n4852), .B2(n4843), .A(n4668), .ZN(n4679) );
  NAND2_X1 U5134 ( .A1(n4670), .A2(n4669), .ZN(n4672) );
  XNOR2_X1 U5135 ( .A(n4672), .B(n4671), .ZN(n4673) );
  NAND2_X1 U5136 ( .A1(n4911), .A2(B_REG_SCAN_IN), .ZN(n4674) );
  AND2_X1 U5137 ( .A1(n4809), .A2(n4674), .ZN(n5280) );
  AOI22_X1 U5138 ( .A1(n4676), .A2(n5280), .B1(n4675), .B2(n5283), .ZN(n4677)
         );
  NAND2_X1 U5139 ( .A1(n4851), .A2(n5173), .ZN(n4678) );
  OAI211_X1 U5140 ( .C1(n4680), .C2(n4806), .A(n4679), .B(n4678), .ZN(U3354)
         );
  OAI21_X1 U5141 ( .B1(n4682), .B2(n4688), .A(n4681), .ZN(n4687) );
  NOR2_X1 U5142 ( .A1(n4683), .A2(n5200), .ZN(n4686) );
  OAI22_X1 U5143 ( .A1(n4684), .A2(n5154), .B1(n4690), .B2(n5293), .ZN(n4685)
         );
  AOI211_X1 U5144 ( .C1(n4687), .C2(n5151), .A(n4686), .B(n4685), .ZN(n4864)
         );
  XNOR2_X1 U5145 ( .A(n4689), .B(n4688), .ZN(n4863) );
  NAND2_X1 U5146 ( .A1(n4863), .A2(n4837), .ZN(n4698) );
  OR2_X1 U5147 ( .A1(n4701), .A2(n4690), .ZN(n4691) );
  NAND2_X1 U5148 ( .A1(n4692), .A2(n4691), .ZN(n4866) );
  INV_X1 U5149 ( .A(n4866), .ZN(n4696) );
  OAI22_X1 U5150 ( .A1(n4694), .A2(n5216), .B1(n4693), .B2(n5173), .ZN(n4695)
         );
  AOI21_X1 U5151 ( .B1(n4696), .B2(n5300), .A(n4695), .ZN(n4697) );
  OAI211_X1 U5152 ( .C1(n4864), .C2(n4847), .A(n4698), .B(n4697), .ZN(U3263)
         );
  XOR2_X1 U5153 ( .A(n4709), .B(n4699), .Z(n4870) );
  INV_X1 U5154 ( .A(n4700), .ZN(n4702) );
  AOI21_X1 U5155 ( .B1(n4703), .B2(n4702), .A(n4701), .ZN(n4868) );
  OAI22_X1 U5156 ( .A1(n4705), .A2(n5216), .B1(n4704), .B2(n5173), .ZN(n4706)
         );
  AOI21_X1 U5157 ( .B1(n4868), .B2(n5300), .A(n4706), .ZN(n4717) );
  NAND2_X1 U5158 ( .A1(n4708), .A2(n4707), .ZN(n4710) );
  XNOR2_X1 U5159 ( .A(n4710), .B(n4709), .ZN(n4715) );
  OAI22_X1 U5160 ( .A1(n4712), .A2(n5200), .B1(n5293), .B2(n4711), .ZN(n4713)
         );
  AOI21_X1 U5161 ( .B1(n5204), .B2(n4726), .A(n4713), .ZN(n4714) );
  OAI21_X1 U5162 ( .B1(n4715), .B2(n5206), .A(n4714), .ZN(n4867) );
  NAND2_X1 U5163 ( .A1(n4867), .A2(n5173), .ZN(n4716) );
  OAI211_X1 U5164 ( .C1(n4870), .C2(n4806), .A(n4717), .B(n4716), .ZN(U3264)
         );
  XNOR2_X1 U5165 ( .A(n4719), .B(n4718), .ZN(n4877) );
  OAI22_X1 U5166 ( .A1(n4720), .A2(n5154), .B1(n4728), .B2(n5293), .ZN(n4725)
         );
  XNOR2_X1 U5167 ( .A(n4722), .B(n4721), .ZN(n4723) );
  NOR2_X1 U5168 ( .A1(n4723), .A2(n5206), .ZN(n4724) );
  AOI211_X1 U5169 ( .C1(n4809), .C2(n4726), .A(n4725), .B(n4724), .ZN(n4876)
         );
  INV_X1 U5170 ( .A(n4876), .ZN(n4734) );
  INV_X1 U5171 ( .A(n4747), .ZN(n4729) );
  OAI211_X1 U5172 ( .C1(n4729), .C2(n4728), .A(n5304), .B(n4727), .ZN(n4875)
         );
  NOR2_X1 U5173 ( .A1(n4875), .A2(n4802), .ZN(n4733) );
  OAI22_X1 U5174 ( .A1(n4731), .A2(n5216), .B1(n4730), .B2(n5173), .ZN(n4732)
         );
  AOI211_X1 U5175 ( .C1(n4734), .C2(n5173), .A(n4733), .B(n4732), .ZN(n4735)
         );
  OAI21_X1 U5176 ( .B1(n4877), .B2(n4806), .A(n4735), .ZN(U3266) );
  XOR2_X1 U5177 ( .A(n4741), .B(n4736), .Z(n4880) );
  INV_X1 U5178 ( .A(n4777), .ZN(n4737) );
  NAND2_X1 U5179 ( .A1(n4778), .A2(n4737), .ZN(n4755) );
  INV_X1 U5180 ( .A(n4757), .ZN(n4738) );
  AND2_X1 U5181 ( .A1(n4756), .A2(n4738), .ZN(n4739) );
  NAND2_X1 U5182 ( .A1(n4755), .A2(n4739), .ZN(n4759) );
  NAND2_X1 U5183 ( .A1(n4759), .A2(n4740), .ZN(n4742) );
  XNOR2_X1 U5184 ( .A(n4742), .B(n4741), .ZN(n4746) );
  NOR2_X1 U5185 ( .A1(n4748), .A2(n5293), .ZN(n4743) );
  OR2_X1 U5186 ( .A1(n4744), .A2(n4743), .ZN(n4745) );
  AOI21_X1 U5187 ( .B1(n4746), .B2(n5151), .A(n4745), .ZN(n4879) );
  INV_X1 U5188 ( .A(n4879), .ZN(n4752) );
  OAI211_X1 U5189 ( .C1(n4767), .C2(n4748), .A(n5304), .B(n4747), .ZN(n4878)
         );
  AOI22_X1 U5190 ( .A1(REG2_REG_23__SCAN_IN), .A2(n5285), .B1(n4749), .B2(
        n5168), .ZN(n4750) );
  OAI21_X1 U5191 ( .B1(n4878), .B2(n4802), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5192 ( .B1(n4752), .B2(n5173), .A(n4751), .ZN(n4753) );
  OAI21_X1 U5193 ( .B1(n4880), .B2(n4806), .A(n4753), .ZN(U3267) );
  XNOR2_X1 U5194 ( .A(n4754), .B(n4756), .ZN(n4883) );
  OAI22_X1 U5195 ( .A1(n5271), .A2(n5154), .B1(n4765), .B2(n5293), .ZN(n4762)
         );
  INV_X1 U5196 ( .A(n4755), .ZN(n4758) );
  OAI21_X1 U5197 ( .B1(n4758), .B2(n4757), .A(n2607), .ZN(n4760) );
  AOI21_X1 U5198 ( .B1(n4760), .B2(n4759), .A(n5206), .ZN(n4761) );
  AOI211_X1 U5199 ( .C1(n4809), .C2(n4763), .A(n4762), .B(n4761), .ZN(n4882)
         );
  INV_X1 U5200 ( .A(n4882), .ZN(n4772) );
  OAI21_X1 U5201 ( .B1(n4764), .B2(n4765), .A(n5304), .ZN(n4766) );
  OR2_X1 U5202 ( .A1(n4767), .A2(n4766), .ZN(n4881) );
  NOR2_X1 U5203 ( .A1(n4881), .A2(n4802), .ZN(n4771) );
  OAI22_X1 U5204 ( .A1(n5173), .A2(n4769), .B1(n4768), .B2(n5216), .ZN(n4770)
         );
  AOI211_X1 U5205 ( .C1(n4772), .C2(n5173), .A(n4771), .B(n4770), .ZN(n4773)
         );
  OAI21_X1 U5206 ( .B1(n4883), .B2(n4806), .A(n4773), .ZN(U3268) );
  OAI21_X1 U5207 ( .B1(n4775), .B2(n4777), .A(n4774), .ZN(n4776) );
  INV_X1 U5208 ( .A(n4776), .ZN(n4886) );
  XNOR2_X1 U5209 ( .A(n4778), .B(n4777), .ZN(n4781) );
  OAI21_X1 U5210 ( .B1(n4783), .B2(n5293), .A(n4779), .ZN(n4780) );
  AOI21_X1 U5211 ( .B1(n4781), .B2(n5151), .A(n4780), .ZN(n4885) );
  INV_X1 U5212 ( .A(n4885), .ZN(n4787) );
  INV_X1 U5213 ( .A(n4764), .ZN(n4782) );
  OAI211_X1 U5214 ( .C1(n4797), .C2(n4783), .A(n4782), .B(n5304), .ZN(n4884)
         );
  AOI22_X1 U5215 ( .A1(n5285), .A2(REG2_REG_21__SCAN_IN), .B1(n4784), .B2(
        n5168), .ZN(n4785) );
  OAI21_X1 U5216 ( .B1(n4884), .B2(n4802), .A(n4785), .ZN(n4786) );
  AOI21_X1 U5217 ( .B1(n4787), .B2(n5173), .A(n4786), .ZN(n4788) );
  OAI21_X1 U5218 ( .B1(n4886), .B2(n4806), .A(n4788), .ZN(U3269) );
  OAI21_X1 U5219 ( .B1(n4790), .B2(n4793), .A(n4789), .ZN(n4791) );
  INV_X1 U5220 ( .A(n4791), .ZN(n4889) );
  XOR2_X1 U5221 ( .A(n4793), .B(n4792), .Z(n4796) );
  AOI22_X1 U5222 ( .A1(n5264), .A2(n5204), .B1(n5262), .B2(n5283), .ZN(n4794)
         );
  OAI21_X1 U5223 ( .B1(n5271), .B2(n5200), .A(n4794), .ZN(n4795) );
  AOI21_X1 U5224 ( .B1(n4796), .B2(n5151), .A(n4795), .ZN(n4888) );
  INV_X1 U5225 ( .A(n4888), .ZN(n4804) );
  INV_X1 U5226 ( .A(n4797), .ZN(n4799) );
  AOI21_X1 U5227 ( .B1(n4819), .B2(n5262), .A(n5229), .ZN(n4798) );
  NAND2_X1 U5228 ( .A1(n4799), .A2(n4798), .ZN(n4887) );
  AOI22_X1 U5229 ( .A1(n5285), .A2(REG2_REG_20__SCAN_IN), .B1(n4800), .B2(
        n5168), .ZN(n4801) );
  OAI21_X1 U5230 ( .B1(n4887), .B2(n4802), .A(n4801), .ZN(n4803) );
  AOI21_X1 U5231 ( .B1(n4804), .B2(n5173), .A(n4803), .ZN(n4805) );
  OAI21_X1 U5232 ( .B1(n4889), .B2(n4806), .A(n4805), .ZN(U3270) );
  NAND3_X1 U5233 ( .A1(n4827), .A2(n4829), .A3(n4826), .ZN(n4828) );
  NAND2_X1 U5234 ( .A1(n4828), .A2(n4807), .ZN(n4808) );
  XNOR2_X1 U5235 ( .A(n4808), .B(n4817), .ZN(n4815) );
  NAND2_X1 U5236 ( .A1(n4810), .A2(n4809), .ZN(n4813) );
  NAND2_X1 U5237 ( .A1(n4811), .A2(n5204), .ZN(n4812) );
  OAI211_X1 U5238 ( .C1(n5293), .C2(n4820), .A(n4813), .B(n4812), .ZN(n4814)
         );
  AOI21_X1 U5239 ( .B1(n4815), .B2(n5151), .A(n4814), .ZN(n4891) );
  OAI21_X1 U5240 ( .B1(n4818), .B2(n4817), .A(n4816), .ZN(n4890) );
  NAND2_X1 U5241 ( .A1(n4890), .A2(n4837), .ZN(n4825) );
  OAI21_X1 U5242 ( .B1(n2533), .B2(n4820), .A(n4819), .ZN(n4893) );
  INV_X1 U5243 ( .A(n4893), .ZN(n4823) );
  OAI22_X1 U5244 ( .A1(n5173), .A2(n4650), .B1(n4821), .B2(n5216), .ZN(n4822)
         );
  AOI21_X1 U5245 ( .B1(n4823), .B2(n5300), .A(n4822), .ZN(n4824) );
  OAI211_X1 U5246 ( .C1(n4847), .C2(n4891), .A(n4825), .B(n4824), .ZN(U3271)
         );
  AND2_X1 U5247 ( .A1(n4827), .A2(n4826), .ZN(n4830) );
  OAI211_X1 U5248 ( .C1(n4830), .C2(n4829), .A(n4828), .B(n5151), .ZN(n4832)
         );
  OAI211_X1 U5249 ( .C1(n5293), .C2(n4833), .A(n4832), .B(n4831), .ZN(n5255)
         );
  INV_X1 U5250 ( .A(n5255), .ZN(n4846) );
  OAI21_X1 U5251 ( .B1(n4836), .B2(n4835), .A(n4834), .ZN(n5258) );
  NAND2_X1 U5252 ( .A1(n5258), .A2(n4837), .ZN(n4845) );
  AOI211_X1 U5253 ( .C1(n4839), .C2(n4838), .A(n5229), .B(n2533), .ZN(n5256)
         );
  INV_X1 U5254 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5255 ( .A1(n5173), .A2(n4841), .B1(n4840), .B2(n5216), .ZN(n4842)
         );
  AOI21_X1 U5256 ( .B1(n5256), .B2(n4843), .A(n4842), .ZN(n4844) );
  OAI211_X1 U5257 ( .C1(n4847), .C2(n4846), .A(n4845), .B(n4844), .ZN(U3272)
         );
  OR3_X1 U5258 ( .A1(n4849), .A2(n4848), .A3(n4915), .ZN(n5230) );
  NAND2_X1 U5259 ( .A1(n4854), .A2(n4853), .ZN(n4858) );
  OAI21_X1 U5260 ( .B1(n4855), .B2(D_REG_1__SCAN_IN), .A(n4907), .ZN(n4857) );
  NAND4_X1 U5261 ( .A1(n4859), .A2(n4858), .A3(n4857), .A4(n4856), .ZN(n4894)
         );
  OAI211_X1 U5262 ( .C1(n4862), .C2(n5111), .A(n4861), .B(n4860), .ZN(n4897)
         );
  MUX2_X1 U5263 ( .A(REG1_REG_28__SCAN_IN), .B(n4897), .S(n5308), .Z(U3546) );
  NAND2_X1 U5264 ( .A1(n4863), .A2(n5257), .ZN(n4865) );
  OAI211_X1 U5265 ( .C1(n5229), .C2(n4866), .A(n4865), .B(n4864), .ZN(n4898)
         );
  MUX2_X1 U5266 ( .A(REG1_REG_27__SCAN_IN), .B(n4898), .S(n5308), .Z(U3545) );
  AOI21_X1 U5267 ( .B1(n5304), .B2(n4868), .A(n4867), .ZN(n4869) );
  OAI21_X1 U5268 ( .B1(n4870), .B2(n5111), .A(n4869), .ZN(n4899) );
  MUX2_X1 U5269 ( .A(REG1_REG_26__SCAN_IN), .B(n4899), .S(n5308), .Z(U3544) );
  AOI21_X1 U5270 ( .B1(n5304), .B2(n4872), .A(n4871), .ZN(n4873) );
  OAI21_X1 U5271 ( .B1(n4874), .B2(n5111), .A(n4873), .ZN(n4900) );
  MUX2_X1 U5272 ( .A(REG1_REG_25__SCAN_IN), .B(n4900), .S(n5308), .Z(U3543) );
  OAI211_X1 U5273 ( .C1(n4877), .C2(n5111), .A(n4876), .B(n4875), .ZN(n4901)
         );
  MUX2_X1 U5274 ( .A(REG1_REG_24__SCAN_IN), .B(n4901), .S(n5308), .Z(U3542) );
  OAI211_X1 U5275 ( .C1(n4880), .C2(n5111), .A(n4879), .B(n4878), .ZN(n4902)
         );
  MUX2_X1 U5276 ( .A(REG1_REG_23__SCAN_IN), .B(n4902), .S(n5308), .Z(U3541) );
  OAI211_X1 U5277 ( .C1(n4883), .C2(n5111), .A(n4882), .B(n4881), .ZN(n4903)
         );
  MUX2_X1 U5278 ( .A(REG1_REG_22__SCAN_IN), .B(n4903), .S(n5308), .Z(U3540) );
  OAI211_X1 U5279 ( .C1(n4886), .C2(n5111), .A(n4885), .B(n4884), .ZN(n4904)
         );
  MUX2_X1 U5280 ( .A(REG1_REG_21__SCAN_IN), .B(n4904), .S(n5308), .Z(U3539) );
  OAI211_X1 U5281 ( .C1(n4889), .C2(n5111), .A(n4888), .B(n4887), .ZN(n4905)
         );
  MUX2_X1 U5282 ( .A(REG1_REG_20__SCAN_IN), .B(n4905), .S(n5308), .Z(U3538) );
  NAND2_X1 U5283 ( .A1(n4890), .A2(n5257), .ZN(n4892) );
  OAI211_X1 U5284 ( .C1(n5229), .C2(n4893), .A(n4892), .B(n4891), .ZN(n4906)
         );
  MUX2_X1 U5285 ( .A(REG1_REG_19__SCAN_IN), .B(n4906), .S(n5308), .Z(U3537) );
  INV_X1 U5286 ( .A(n4894), .ZN(n4896) );
  MUX2_X1 U5287 ( .A(REG0_REG_28__SCAN_IN), .B(n4897), .S(n5312), .Z(U3514) );
  MUX2_X1 U5288 ( .A(REG0_REG_27__SCAN_IN), .B(n4898), .S(n5312), .Z(U3513) );
  MUX2_X1 U5289 ( .A(REG0_REG_26__SCAN_IN), .B(n4899), .S(n5312), .Z(U3512) );
  MUX2_X1 U5290 ( .A(REG0_REG_25__SCAN_IN), .B(n4900), .S(n5312), .Z(U3511) );
  MUX2_X1 U5291 ( .A(REG0_REG_24__SCAN_IN), .B(n4901), .S(n5312), .Z(U3510) );
  MUX2_X1 U5292 ( .A(REG0_REG_23__SCAN_IN), .B(n4902), .S(n5312), .Z(U3509) );
  MUX2_X1 U5293 ( .A(REG0_REG_22__SCAN_IN), .B(n4903), .S(n5312), .Z(U3508) );
  MUX2_X1 U5294 ( .A(REG0_REG_21__SCAN_IN), .B(n4904), .S(n5312), .Z(U3507) );
  MUX2_X1 U5295 ( .A(REG0_REG_20__SCAN_IN), .B(n4905), .S(n5312), .Z(U3506) );
  MUX2_X1 U5296 ( .A(REG0_REG_19__SCAN_IN), .B(n4906), .S(n5312), .Z(U3505) );
  MUX2_X1 U5297 ( .A(n4907), .B(D_REG_1__SCAN_IN), .S(n4951), .Z(U3459) );
  NOR3_X1 U5298 ( .A1(n2782), .A2(IR_REG_30__SCAN_IN), .A3(n4908), .ZN(n4909)
         );
  MUX2_X1 U5299 ( .A(DATAI_31_), .B(n4909), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5300 ( .A(DATAI_30_), .B(n4910), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5301 ( .A(n2786), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5302 ( .A(n4911), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5303 ( .A(n4912), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5304 ( .A(n4913), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5305 ( .A(n4914), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5306 ( .A(n4915), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5307 ( .A(n4916), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5308 ( .A(DATAI_19_), .B(n5064), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5309 ( .A(DATAI_18_), .B(n4917), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5310 ( .A(n4918), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5311 ( .A(DATAI_16_), .B(n4919), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5312 ( .A(n4920), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5313 ( .A(n5016), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5314 ( .A(DATAI_13_), .B(n4998), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5315 ( .A(n4921), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5316 ( .A(n4922), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5317 ( .A(DATAI_8_), .B(n4978), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5318 ( .A(n4923), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5319 ( .A(n4970), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5320 ( .A(DATAI_5_), .B(n4924), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5321 ( .A(n5045), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5322 ( .A(n4958), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5323 ( .A(n4925), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5324 ( .A(n4926), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5325 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X2 U5326 ( .A(n4951), .ZN(n4953) );
  INV_X1 U5327 ( .A(D_REG_2__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U5328 ( .A1(n4953), .A2(n4927), .ZN(U3320) );
  AND2_X1 U5329 ( .A1(n4951), .A2(D_REG_3__SCAN_IN), .ZN(U3319) );
  NOR2_X1 U5330 ( .A1(n4953), .A2(n4928), .ZN(U3318) );
  NOR2_X1 U5331 ( .A1(n4953), .A2(n4929), .ZN(U3317) );
  NOR2_X1 U5332 ( .A1(n4953), .A2(n4930), .ZN(U3316) );
  NOR2_X1 U5333 ( .A1(n4953), .A2(n4931), .ZN(U3315) );
  AND2_X1 U5334 ( .A1(n4951), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  INV_X1 U5335 ( .A(D_REG_9__SCAN_IN), .ZN(n4932) );
  NOR2_X1 U5336 ( .A1(n4953), .A2(n4932), .ZN(U3313) );
  NOR2_X1 U5337 ( .A1(n4953), .A2(n4933), .ZN(U3312) );
  NOR2_X1 U5338 ( .A1(n4953), .A2(n4934), .ZN(U3311) );
  NOR2_X1 U5339 ( .A1(n4953), .A2(n4935), .ZN(U3310) );
  NOR2_X1 U5340 ( .A1(n4953), .A2(n4936), .ZN(U3309) );
  NOR2_X1 U5341 ( .A1(n4953), .A2(n4937), .ZN(U3308) );
  NOR2_X1 U5342 ( .A1(n4953), .A2(n4938), .ZN(U3307) );
  NOR2_X1 U5343 ( .A1(n4953), .A2(n4939), .ZN(U3306) );
  NOR2_X1 U5344 ( .A1(n4953), .A2(n4940), .ZN(U3305) );
  NOR2_X1 U5345 ( .A1(n4953), .A2(n4941), .ZN(U3304) );
  NOR2_X1 U5346 ( .A1(n4953), .A2(n4942), .ZN(U3303) );
  AND2_X1 U5347 ( .A1(n4951), .A2(D_REG_20__SCAN_IN), .ZN(U3302) );
  NOR2_X1 U5348 ( .A1(n4953), .A2(n4943), .ZN(U3301) );
  INV_X1 U5349 ( .A(D_REG_22__SCAN_IN), .ZN(n4944) );
  NOR2_X1 U5350 ( .A1(n4953), .A2(n4944), .ZN(U3300) );
  AND2_X1 U5351 ( .A1(n4951), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  INV_X1 U5352 ( .A(D_REG_24__SCAN_IN), .ZN(n4945) );
  NOR2_X1 U5353 ( .A1(n4953), .A2(n4945), .ZN(U3298) );
  NOR2_X1 U5354 ( .A1(n4953), .A2(n4946), .ZN(U3297) );
  INV_X1 U5355 ( .A(D_REG_26__SCAN_IN), .ZN(n4947) );
  NOR2_X1 U5356 ( .A1(n4953), .A2(n4947), .ZN(U3296) );
  NOR2_X1 U5357 ( .A1(n4953), .A2(n4948), .ZN(U3295) );
  NOR2_X1 U5358 ( .A1(n4953), .A2(n4949), .ZN(U3294) );
  NOR2_X1 U5359 ( .A1(n4953), .A2(n4950), .ZN(U3293) );
  AND2_X1 U5360 ( .A1(n4951), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  INV_X1 U5361 ( .A(D_REG_31__SCAN_IN), .ZN(n4952) );
  NOR2_X1 U5362 ( .A1(n4953), .A2(n4952), .ZN(U3291) );
  INV_X1 U5363 ( .A(n4954), .ZN(n4955) );
  AOI21_X1 U5364 ( .B1(n5053), .B2(ADDR_REG_3__SCAN_IN), .A(n4955), .ZN(n4964)
         );
  OAI211_X1 U5365 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4957), .A(n5043), .B(n4956), 
        .ZN(n4963) );
  NAND2_X1 U5366 ( .A1(n5046), .A2(n4958), .ZN(n4962) );
  XOR2_X1 U5367 ( .A(n4959), .B(REG1_REG_3__SCAN_IN), .Z(n4960) );
  NAND2_X1 U5368 ( .A1(n5033), .A2(n4960), .ZN(n4961) );
  NAND4_X1 U5369 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(U3243)
         );
  AOI21_X1 U5370 ( .B1(n5053), .B2(ADDR_REG_6__SCAN_IN), .A(n4965), .ZN(n4974)
         );
  OAI211_X1 U5371 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4967), .A(n5043), .B(n4966), 
        .ZN(n4973) );
  OAI211_X1 U5372 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4969), .A(n5033), .B(n4968), 
        .ZN(n4972) );
  NAND2_X1 U5373 ( .A1(n5046), .A2(n4970), .ZN(n4971) );
  NAND4_X1 U5374 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(U3246)
         );
  AOI21_X1 U5375 ( .B1(n5053), .B2(ADDR_REG_8__SCAN_IN), .A(n4975), .ZN(n4984)
         );
  OAI211_X1 U5376 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4977), .A(n5033), .B(n4976), 
        .ZN(n4983) );
  NAND2_X1 U5377 ( .A1(n5046), .A2(n4978), .ZN(n4982) );
  OAI211_X1 U5378 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4980), .A(n5043), .B(n4979), 
        .ZN(n4981) );
  NAND4_X1 U5379 ( .A1(n4984), .A2(n4983), .A3(n4982), .A4(n4981), .ZN(U3248)
         );
  OAI211_X1 U5380 ( .C1(n4987), .C2(n4986), .A(n5033), .B(n4985), .ZN(n4992)
         );
  OAI211_X1 U5381 ( .C1(n4990), .C2(n4989), .A(n5043), .B(n4988), .ZN(n4991)
         );
  OAI211_X1 U5382 ( .C1(n5009), .C2(n4993), .A(n4992), .B(n4991), .ZN(n4994)
         );
  AOI211_X1 U5383 ( .C1(n5053), .C2(ADDR_REG_9__SCAN_IN), .A(n4995), .B(n4994), 
        .ZN(n4996) );
  INV_X1 U5384 ( .A(n4996), .ZN(U3249) );
  NOR2_X1 U5385 ( .A1(STATE_REG_SCAN_IN), .A2(n4997), .ZN(n5186) );
  INV_X1 U5386 ( .A(n4998), .ZN(n5008) );
  NAND2_X1 U5387 ( .A1(n5008), .A2(REG1_REG_13__SCAN_IN), .ZN(n5000) );
  OAI211_X1 U5388 ( .C1(REG1_REG_13__SCAN_IN), .C2(n5008), .A(n5001), .B(n5000), .ZN(n5002) );
  NAND3_X1 U5389 ( .A1(n4999), .A2(n5033), .A3(n5002), .ZN(n5007) );
  OAI211_X1 U5390 ( .C1(n5005), .C2(n5004), .A(n5043), .B(n5003), .ZN(n5006)
         );
  OAI211_X1 U5391 ( .C1(n5009), .C2(n5008), .A(n5007), .B(n5006), .ZN(n5010)
         );
  AOI211_X1 U5392 ( .C1(n5053), .C2(ADDR_REG_13__SCAN_IN), .A(n5186), .B(n5010), .ZN(n5011) );
  INV_X1 U5393 ( .A(n5011), .ZN(U3253) );
  INV_X1 U5394 ( .A(n5012), .ZN(n5013) );
  AOI21_X1 U5395 ( .B1(n5053), .B2(ADDR_REG_14__SCAN_IN), .A(n5013), .ZN(n5022) );
  XOR2_X1 U5396 ( .A(REG1_REG_14__SCAN_IN), .B(n5014), .Z(n5015) );
  NAND2_X1 U5397 ( .A1(n5015), .A2(n5033), .ZN(n5021) );
  NAND2_X1 U5398 ( .A1(n5046), .A2(n5016), .ZN(n5020) );
  OAI211_X1 U5399 ( .C1(REG2_REG_14__SCAN_IN), .C2(n5018), .A(n5043), .B(n5017), .ZN(n5019) );
  NAND4_X1 U5400 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(U3254)
         );
  NOR2_X1 U5401 ( .A1(n5049), .A2(n5252), .ZN(n5026) );
  INV_X1 U5402 ( .A(n5029), .ZN(n5023) );
  NOR3_X1 U5403 ( .A1(n5024), .A2(n3557), .A3(n5023), .ZN(n5025) );
  AOI211_X1 U5404 ( .C1(n5036), .C2(n5026), .A(n5046), .B(n5025), .ZN(n5040)
         );
  OAI211_X1 U5405 ( .C1(n5029), .C2(n5028), .A(n5043), .B(n5027), .ZN(n5031)
         );
  NAND2_X1 U5406 ( .A1(n5031), .A2(n5030), .ZN(n5032) );
  AOI21_X1 U5407 ( .B1(n5053), .B2(ADDR_REG_17__SCAN_IN), .A(n5032), .ZN(n5038) );
  OAI211_X1 U5408 ( .C1(n5036), .C2(n5035), .A(n5034), .B(n5033), .ZN(n5037)
         );
  OAI211_X1 U5409 ( .C1(n5040), .C2(n5039), .A(n5038), .B(n5037), .ZN(U3257)
         );
  XNOR2_X1 U5410 ( .A(n5041), .B(REG1_REG_4__SCAN_IN), .ZN(n5050) );
  OAI211_X1 U5411 ( .C1(REG2_REG_4__SCAN_IN), .C2(n5044), .A(n5043), .B(n5042), 
        .ZN(n5048) );
  NAND2_X1 U5412 ( .A1(n5046), .A2(n5045), .ZN(n5047) );
  OAI211_X1 U5413 ( .C1(n5050), .C2(n5049), .A(n5048), .B(n5047), .ZN(n5051)
         );
  AOI211_X1 U5414 ( .C1(n5053), .C2(ADDR_REG_4__SCAN_IN), .A(n5052), .B(n5051), 
        .ZN(n5055) );
  NAND2_X1 U5415 ( .A1(n5055), .A2(n5054), .ZN(U3244) );
  INV_X1 U5416 ( .A(n5230), .ZN(n5212) );
  INV_X1 U5417 ( .A(n5060), .ZN(n5068) );
  NOR2_X1 U5418 ( .A1(n5057), .A2(n5056), .ZN(n5067) );
  NOR2_X1 U5419 ( .A1(n5209), .A2(n5151), .ZN(n5059) );
  OAI22_X1 U5420 ( .A1(n5060), .A2(n5059), .B1(n5058), .B2(n5200), .ZN(n5065)
         );
  AOI211_X1 U5421 ( .C1(n5212), .C2(n5068), .A(n5067), .B(n5065), .ZN(n5063)
         );
  AOI22_X1 U5422 ( .A1(n5308), .A2(n5063), .B1(n5061), .B2(n5306), .ZN(U3518)
         );
  INV_X1 U5423 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U5424 ( .A1(n5312), .A2(n5063), .B1(n5062), .B2(n5309), .ZN(U3467)
         );
  NAND2_X1 U5425 ( .A1(n2517), .A2(n5064), .ZN(n5066) );
  AOI21_X1 U5426 ( .B1(n5067), .B2(n5066), .A(n5065), .ZN(n5071) );
  AOI22_X1 U5427 ( .A1(n5068), .A2(n5222), .B1(REG3_REG_0__SCAN_IN), .B2(n5168), .ZN(n5069) );
  OAI221_X1 U5428 ( .B1(n4847), .B2(n5071), .C1(n5173), .C2(n5070), .A(n5069), 
        .ZN(U3290) );
  NOR2_X1 U5429 ( .A1(n5072), .A2(n5111), .ZN(n5074) );
  AOI211_X1 U5430 ( .C1(n5304), .C2(n5075), .A(n5074), .B(n5073), .ZN(n5077)
         );
  AOI22_X1 U5431 ( .A1(n5308), .A2(n5077), .B1(n2882), .B2(n5306), .ZN(U3519)
         );
  INV_X1 U5432 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U5433 ( .A1(n5312), .A2(n5077), .B1(n5076), .B2(n5309), .ZN(U3469)
         );
  NOR2_X1 U5434 ( .A1(n5078), .A2(n5229), .ZN(n5080) );
  AOI211_X1 U5435 ( .C1(n5212), .C2(n5081), .A(n5080), .B(n5079), .ZN(n5083)
         );
  AOI22_X1 U5436 ( .A1(n5308), .A2(n5083), .B1(n2881), .B2(n5306), .ZN(U3520)
         );
  INV_X1 U5437 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U5438 ( .A1(n5312), .A2(n5083), .B1(n5082), .B2(n5309), .ZN(U3471)
         );
  OAI21_X1 U5439 ( .B1(n5229), .B2(n5085), .A(n5084), .ZN(n5086) );
  AOI21_X1 U5440 ( .B1(n5257), .B2(n5087), .A(n5086), .ZN(n5089) );
  AOI22_X1 U5441 ( .A1(n5308), .A2(n5089), .B1(n2939), .B2(n5306), .ZN(U3521)
         );
  INV_X1 U5442 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U5443 ( .A1(n5312), .A2(n5089), .B1(n5088), .B2(n5309), .ZN(U3473)
         );
  INV_X1 U5444 ( .A(n5090), .ZN(n5093) );
  AOI211_X1 U5445 ( .C1(n5093), .C2(n5212), .A(n5092), .B(n5091), .ZN(n5096)
         );
  INV_X1 U5446 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U5447 ( .A1(n5308), .A2(n5096), .B1(n5094), .B2(n5306), .ZN(U3522)
         );
  INV_X1 U5448 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5095) );
  AOI22_X1 U5449 ( .A1(n5312), .A2(n5096), .B1(n5095), .B2(n5309), .ZN(U3475)
         );
  NOR3_X1 U5450 ( .A1(n5098), .A2(n5097), .A3(n5229), .ZN(n5100) );
  AOI211_X1 U5451 ( .C1(n5257), .C2(n5101), .A(n5100), .B(n5099), .ZN(n5103)
         );
  AOI22_X1 U5452 ( .A1(n5308), .A2(n5103), .B1(n2892), .B2(n5306), .ZN(U3523)
         );
  INV_X1 U5453 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5102) );
  AOI22_X1 U5454 ( .A1(n5312), .A2(n5103), .B1(n5102), .B2(n5309), .ZN(U3477)
         );
  AND3_X1 U5455 ( .A1(n3181), .A2(n5257), .A3(n5104), .ZN(n5105) );
  AOI211_X1 U5456 ( .C1(n5304), .C2(n5107), .A(n5106), .B(n5105), .ZN(n5110)
         );
  INV_X1 U5457 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5108) );
  AOI22_X1 U5458 ( .A1(n5308), .A2(n5110), .B1(n5108), .B2(n5306), .ZN(U3524)
         );
  INV_X1 U5459 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U5460 ( .A1(n5312), .A2(n5110), .B1(n5109), .B2(n5309), .ZN(U3479)
         );
  OR2_X1 U5461 ( .A1(n5112), .A2(n5111), .ZN(n5116) );
  AND2_X1 U5462 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  AOI22_X1 U5463 ( .A1(n5308), .A2(n5118), .B1(n4582), .B2(n5306), .ZN(U3525)
         );
  INV_X1 U5464 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U5465 ( .A1(n5312), .A2(n5118), .B1(n5117), .B2(n5309), .ZN(U3481)
         );
  AOI22_X1 U5466 ( .A1(n5120), .A2(n5212), .B1(n5304), .B2(n5119), .ZN(n5121)
         );
  AND2_X1 U5467 ( .A1(n5122), .A2(n5121), .ZN(n5124) );
  INV_X1 U5468 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5123) );
  AOI22_X1 U5469 ( .A1(n5308), .A2(n5124), .B1(n5123), .B2(n5306), .ZN(U3526)
         );
  AOI22_X1 U5470 ( .A1(n5312), .A2(n5124), .B1(n4250), .B2(n5309), .ZN(U3483)
         );
  INV_X1 U5471 ( .A(n5125), .ZN(n5126) );
  NOR3_X1 U5472 ( .A1(n5127), .A2(n5126), .A3(n5229), .ZN(n5129) );
  AOI211_X1 U5473 ( .C1(n5130), .C2(n5257), .A(n5129), .B(n5128), .ZN(n5132)
         );
  AOI22_X1 U5474 ( .A1(n5308), .A2(n5132), .B1(n2864), .B2(n5306), .ZN(U3527)
         );
  INV_X1 U5475 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5131) );
  AOI22_X1 U5476 ( .A1(n5312), .A2(n5132), .B1(n5131), .B2(n5309), .ZN(U3485)
         );
  AND3_X1 U5477 ( .A1(n5142), .A2(n5257), .A3(n5133), .ZN(n5134) );
  AOI211_X1 U5478 ( .C1(n5304), .C2(n5136), .A(n5135), .B(n5134), .ZN(n5139)
         );
  INV_X1 U5479 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5137) );
  AOI22_X1 U5480 ( .A1(n5308), .A2(n5139), .B1(n5137), .B2(n5306), .ZN(U3528)
         );
  INV_X1 U5481 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5138) );
  AOI22_X1 U5482 ( .A1(n5312), .A2(n5139), .B1(n5138), .B2(n5309), .ZN(U3487)
         );
  AND2_X1 U5483 ( .A1(n5142), .A2(n5140), .ZN(n5144) );
  NAND2_X1 U5484 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  OAI21_X1 U5485 ( .B1(n5144), .B2(n5149), .A(n5143), .ZN(n5166) );
  INV_X1 U5486 ( .A(n5145), .ZN(n5148) );
  INV_X1 U5487 ( .A(n5146), .ZN(n5147) );
  OAI21_X1 U5488 ( .B1(n5148), .B2(n5153), .A(n5147), .ZN(n5167) );
  NOR2_X1 U5489 ( .A1(n5167), .A2(n5229), .ZN(n5160) );
  XNOR2_X1 U5490 ( .A(n5150), .B(n5149), .ZN(n5152) );
  NAND2_X1 U5491 ( .A1(n5152), .A2(n5151), .ZN(n5158) );
  OAI22_X1 U5492 ( .A1(n5155), .A2(n5154), .B1(n5153), .B2(n5293), .ZN(n5156)
         );
  INV_X1 U5493 ( .A(n5156), .ZN(n5157) );
  OAI211_X1 U5494 ( .C1(n5159), .C2(n5200), .A(n5158), .B(n5157), .ZN(n5164)
         );
  AOI211_X1 U5495 ( .C1(n5166), .C2(n5257), .A(n5160), .B(n5164), .ZN(n5163)
         );
  AOI22_X1 U5496 ( .A1(n5308), .A2(n5163), .B1(n5161), .B2(n5306), .ZN(U3529)
         );
  INV_X1 U5497 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5162) );
  AOI22_X1 U5498 ( .A1(n5312), .A2(n5163), .B1(n5162), .B2(n5309), .ZN(U3489)
         );
  AOI21_X1 U5499 ( .B1(n5166), .B2(n5165), .A(n5164), .ZN(n5174) );
  INV_X1 U5500 ( .A(n5167), .ZN(n5170) );
  AOI22_X1 U5501 ( .A1(n5170), .A2(n5300), .B1(n5169), .B2(n5168), .ZN(n5171)
         );
  OAI221_X1 U5502 ( .B1(n4847), .B2(n5174), .C1(n5173), .C2(n5172), .A(n5171), 
        .ZN(U3279) );
  OAI21_X1 U5503 ( .B1(n5176), .B2(n5229), .A(n5175), .ZN(n5177) );
  AOI21_X1 U5504 ( .B1(n5178), .B2(n5257), .A(n5177), .ZN(n5181) );
  INV_X1 U5505 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5179) );
  AOI22_X1 U5506 ( .A1(n5308), .A2(n5181), .B1(n5179), .B2(n5306), .ZN(U3530)
         );
  INV_X1 U5507 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5180) );
  AOI22_X1 U5508 ( .A1(n5312), .A2(n5181), .B1(n5180), .B2(n5309), .ZN(U3491)
         );
  AOI22_X1 U5509 ( .A1(n5265), .A2(n5203), .B1(n5263), .B2(n5182), .ZN(n5189)
         );
  XNOR2_X1 U5510 ( .A(n5184), .B(n5183), .ZN(n5187) );
  NOR2_X1 U5511 ( .A1(n5272), .A2(n5201), .ZN(n5185) );
  AOI211_X1 U5512 ( .C1(n5187), .C2(n5274), .A(n5186), .B(n5185), .ZN(n5188)
         );
  OAI211_X1 U5513 ( .C1(n5279), .C2(n5217), .A(n5189), .B(n5188), .ZN(U3231)
         );
  OR2_X1 U5514 ( .A1(n3372), .A2(n5190), .ZN(n5192) );
  XOR2_X1 U5515 ( .A(n5198), .B(n5193), .Z(n5223) );
  OAI21_X1 U5516 ( .B1(n5194), .B2(n5199), .A(n2521), .ZN(n5220) );
  NOR2_X1 U5517 ( .A1(n5220), .A2(n5229), .ZN(n5211) );
  NOR2_X1 U5518 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  XNOR2_X1 U5519 ( .A(n5198), .B(n5197), .ZN(n5207) );
  OAI22_X1 U5520 ( .A1(n5201), .A2(n5200), .B1(n5293), .B2(n5199), .ZN(n5202)
         );
  AOI21_X1 U5521 ( .B1(n5204), .B2(n5203), .A(n5202), .ZN(n5205) );
  OAI21_X1 U5522 ( .B1(n5207), .B2(n5206), .A(n5205), .ZN(n5208) );
  AOI21_X1 U5523 ( .B1(n5223), .B2(n5209), .A(n5208), .ZN(n5226) );
  INV_X1 U5524 ( .A(n5226), .ZN(n5210) );
  AOI211_X1 U5525 ( .C1(n5212), .C2(n5223), .A(n5211), .B(n5210), .ZN(n5215)
         );
  INV_X1 U5526 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5213) );
  AOI22_X1 U5527 ( .A1(n5308), .A2(n5215), .B1(n5213), .B2(n5306), .ZN(U3531)
         );
  INV_X1 U5528 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5214) );
  AOI22_X1 U5529 ( .A1(n5312), .A2(n5215), .B1(n5214), .B2(n5309), .ZN(U3493)
         );
  INV_X1 U5530 ( .A(REG2_REG_13__SCAN_IN), .ZN(n5218) );
  OAI22_X1 U5531 ( .A1(n5173), .A2(n5218), .B1(n5217), .B2(n5216), .ZN(n5219)
         );
  INV_X1 U5532 ( .A(n5219), .ZN(n5225) );
  INV_X1 U5533 ( .A(n5220), .ZN(n5221) );
  AOI22_X1 U5534 ( .A1(n5223), .A2(n5222), .B1(n5300), .B2(n5221), .ZN(n5224)
         );
  OAI211_X1 U5535 ( .C1(n4847), .C2(n5226), .A(n5225), .B(n5224), .ZN(U3277)
         );
  INV_X1 U5536 ( .A(n5227), .ZN(n5228) );
  OAI22_X1 U5537 ( .A1(n5231), .A2(n5230), .B1(n5229), .B2(n5228), .ZN(n5232)
         );
  NOR2_X1 U5538 ( .A1(n5233), .A2(n5232), .ZN(n5236) );
  INV_X1 U5539 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5234) );
  AOI22_X1 U5540 ( .A1(n5308), .A2(n5236), .B1(n5234), .B2(n5306), .ZN(U3532)
         );
  INV_X1 U5541 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5235) );
  AOI22_X1 U5542 ( .A1(n5312), .A2(n5236), .B1(n5235), .B2(n5309), .ZN(U3495)
         );
  AOI211_X1 U5543 ( .C1(n5239), .C2(n5257), .A(n5238), .B(n5237), .ZN(n5242)
         );
  AOI22_X1 U5544 ( .A1(n5308), .A2(n5242), .B1(n5240), .B2(n5306), .ZN(U3533)
         );
  INV_X1 U5545 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5241) );
  AOI22_X1 U5546 ( .A1(n5312), .A2(n5242), .B1(n5241), .B2(n5309), .ZN(U3497)
         );
  AOI211_X1 U5547 ( .C1(n5245), .C2(n5257), .A(n5244), .B(n5243), .ZN(n5248)
         );
  INV_X1 U5548 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U5549 ( .A1(n5308), .A2(n5248), .B1(n5246), .B2(n5306), .ZN(U3534)
         );
  INV_X1 U5550 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5247) );
  AOI22_X1 U5551 ( .A1(n5312), .A2(n5248), .B1(n5247), .B2(n5309), .ZN(U3499)
         );
  AOI211_X1 U5552 ( .C1(n5251), .C2(n5257), .A(n5250), .B(n5249), .ZN(n5254)
         );
  AOI22_X1 U5553 ( .A1(n5308), .A2(n5254), .B1(n5252), .B2(n5306), .ZN(U3535)
         );
  INV_X1 U5554 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5253) );
  AOI22_X1 U5555 ( .A1(n5312), .A2(n5254), .B1(n5253), .B2(n5309), .ZN(U3501)
         );
  AOI211_X1 U5556 ( .C1(n5258), .C2(n5257), .A(n5256), .B(n5255), .ZN(n5261)
         );
  AOI22_X1 U5557 ( .A1(n5308), .A2(n5261), .B1(n5259), .B2(n5306), .ZN(U3536)
         );
  INV_X1 U5558 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5260) );
  AOI22_X1 U5559 ( .A1(n5312), .A2(n5261), .B1(n5260), .B2(n5309), .ZN(U3503)
         );
  AOI22_X1 U5560 ( .A1(n5265), .A2(n5264), .B1(n5263), .B2(n5262), .ZN(n5277)
         );
  NAND2_X1 U5561 ( .A1(n5267), .A2(n5266), .ZN(n5269) );
  XOR2_X1 U5562 ( .A(n5269), .B(n5268), .Z(n5275) );
  INV_X1 U5563 ( .A(REG3_REG_20__SCAN_IN), .ZN(n5270) );
  OAI22_X1 U5564 ( .A1(n5272), .A2(n5271), .B1(STATE_REG_SCAN_IN), .B2(n5270), 
        .ZN(n5273) );
  AOI21_X1 U5565 ( .B1(n5275), .B2(n5274), .A(n5273), .ZN(n5276) );
  OAI211_X1 U5566 ( .C1(n5279), .C2(n5278), .A(n5277), .B(n5276), .ZN(U3230)
         );
  INV_X1 U5567 ( .A(n5296), .ZN(n5284) );
  NAND2_X1 U5568 ( .A1(n5281), .A2(n5280), .ZN(n5295) );
  INV_X1 U5569 ( .A(n5295), .ZN(n5282) );
  AOI21_X1 U5570 ( .B1(n5284), .B2(n5283), .A(n5282), .ZN(n5287) );
  XOR2_X1 U5571 ( .A(n5296), .B(n5297), .Z(n5289) );
  AOI22_X1 U5572 ( .A1(n5289), .A2(n5300), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5285), .ZN(n5286) );
  OAI21_X1 U5573 ( .B1(n4847), .B2(n5287), .A(n5286), .ZN(U3261) );
  INV_X1 U5574 ( .A(n5287), .ZN(n5288) );
  AOI21_X1 U5575 ( .B1(n5289), .B2(n5304), .A(n5288), .ZN(n5292) );
  INV_X1 U5576 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5290) );
  AOI22_X1 U5577 ( .A1(n5308), .A2(n5292), .B1(n5290), .B2(n5306), .ZN(U3548)
         );
  INV_X1 U5578 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5291) );
  AOI22_X1 U5579 ( .A1(n5312), .A2(n5292), .B1(n5291), .B2(n5309), .ZN(U3516)
         );
  OR2_X1 U5580 ( .A1(n5298), .A2(n5293), .ZN(n5294) );
  AND2_X1 U5581 ( .A1(n5295), .A2(n5294), .ZN(n5302) );
  NAND2_X1 U5582 ( .A1(n5297), .A2(n5296), .ZN(n5299) );
  XNOR2_X1 U5583 ( .A(n5299), .B(n5298), .ZN(n5305) );
  AOI22_X1 U5584 ( .A1(n5305), .A2(n5300), .B1(n4847), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5301) );
  OAI21_X1 U5585 ( .B1(n4847), .B2(n5302), .A(n5301), .ZN(U3260) );
  INV_X1 U5586 ( .A(n5302), .ZN(n5303) );
  AOI21_X1 U5587 ( .B1(n5305), .B2(n5304), .A(n5303), .ZN(n5311) );
  INV_X1 U5588 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5307) );
  AOI22_X1 U5589 ( .A1(n5308), .A2(n5311), .B1(n5307), .B2(n5306), .ZN(U3549)
         );
  INV_X1 U5590 ( .A(REG0_REG_31__SCAN_IN), .ZN(n5310) );
  AOI22_X1 U5591 ( .A1(n5312), .A2(n5311), .B1(n5310), .B2(n5309), .ZN(U3517)
         );
  CLKBUF_X1 U2559 ( .A(n3456), .Z(n3719) );
  CLKBUF_X1 U3426 ( .A(n2792), .Z(n2516) );
endmodule

