

module b22_C_SARLock_k_128_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6593, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15648;

  NOR2_X1 U7317 ( .A1(n14806), .A2(n14805), .ZN(n15018) );
  OAI21_X1 U7318 ( .B1(n13418), .B2(n7342), .A(n7338), .ZN(n13474) );
  INV_X2 U7319 ( .A(n12370), .ZN(n12363) );
  XNOR2_X1 U7320 ( .A(n14730), .B(n15525), .ZN(n14772) );
  CLKBUF_X2 U7322 ( .A(n6603), .Z(n9294) );
  AND2_X1 U7323 ( .A1(n11693), .A2(n11701), .ZN(n11658) );
  INV_X1 U7324 ( .A(n8740), .ZN(n8724) );
  NAND2_X1 U7325 ( .A1(n9505), .A2(n14046), .ZN(n11955) );
  INV_X2 U7326 ( .A(n8428), .ZN(n9162) );
  XNOR2_X1 U7327 ( .A(n8322), .B(SI_1_), .ZN(n8443) );
  INV_X1 U7328 ( .A(n12178), .ZN(n12207) );
  NAND2_X1 U7329 ( .A1(n11692), .A2(n11700), .ZN(n8124) );
  NAND2_X1 U7330 ( .A1(n15155), .A2(n14171), .ZN(n11956) );
  BUF_X1 U7331 ( .A(n12303), .Z(n12327) );
  INV_X1 U7332 ( .A(n13512), .ZN(n6814) );
  INV_X1 U7333 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8412) );
  INV_X1 U7334 ( .A(n12369), .ZN(n12412) );
  INV_X1 U7335 ( .A(n9511), .ZN(n12219) );
  NAND2_X2 U7336 ( .A1(n12238), .A2(n11925), .ZN(n15091) );
  NAND2_X1 U7337 ( .A1(n7858), .A2(n11715), .ZN(n11040) );
  NAND2_X1 U7338 ( .A1(n11635), .A2(n11634), .ZN(n14947) );
  NAND2_X1 U7339 ( .A1(n13267), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7731) );
  OAI21_X2 U7340 ( .B1(n12124), .B2(n8802), .A(n8803), .ZN(n13925) );
  NAND2_X1 U7341 ( .A1(n8709), .A2(n8708), .ZN(n13957) );
  AND2_X1 U7342 ( .A1(n8249), .A2(n8250), .ZN(n10718) );
  NAND2_X1 U7343 ( .A1(n12146), .A2(n12145), .ZN(n14630) );
  XNOR2_X1 U7344 ( .A(n9446), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U7345 ( .A1(n7410), .A2(n14780), .ZN(n14781) );
  NAND2_X1 U7346 ( .A1(n8411), .A2(n8410), .ZN(n14014) );
  AND3_X1 U7347 ( .A1(n6788), .A2(n7762), .A3(n7763), .ZN(n6568) );
  INV_X1 U7348 ( .A(n12370), .ZN(n12329) );
  NAND2_X2 U7349 ( .A1(n8823), .A2(n8400), .ZN(n8824) );
  NAND2_X2 U7350 ( .A1(n6735), .A2(n7697), .ZN(n7954) );
  NOR2_X2 U7351 ( .A1(n6827), .A2(n7379), .ZN(n7378) );
  OAI21_X2 U7352 ( .B1(n11125), .B2(n9334), .A(n10606), .ZN(n10792) );
  NAND2_X2 U7353 ( .A1(n10608), .A2(n10607), .ZN(n10606) );
  AND2_X2 U7354 ( .A1(n12724), .A2(n11808), .ZN(n12707) );
  OAI21_X2 U7355 ( .B1(n10193), .B2(n10212), .A(n10320), .ZN(n10194) );
  NOR2_X1 U7356 ( .A1(n6699), .A2(n6746), .ZN(n6745) );
  NAND2_X2 U7357 ( .A1(n7376), .A2(n7375), .ZN(n8669) );
  NAND2_X2 U7358 ( .A1(n7734), .A2(n7737), .ZN(n8082) );
  NAND2_X1 U7359 ( .A1(n7738), .A2(n7737), .ZN(n11639) );
  AOI21_X2 U7360 ( .B1(n6948), .B2(n6950), .A(n6677), .ZN(n6946) );
  XNOR2_X2 U7361 ( .A(n7258), .B(n6854), .ZN(n7257) );
  OAI21_X2 U7362 ( .B1(n14372), .B2(n7149), .A(n7147), .ZN(n14519) );
  NAND2_X2 U7363 ( .A1(n14565), .A2(n14369), .ZN(n14372) );
  XNOR2_X2 U7364 ( .A(n14726), .B(n15489), .ZN(n14769) );
  OAI211_X2 U7365 ( .C1(n11388), .C2(n7508), .A(n7510), .B(1'b1), .ZN(n11582)
         );
  OR2_X2 U7366 ( .A1(n8875), .A2(n8957), .ZN(n13879) );
  AOI21_X2 U7367 ( .B1(n10589), .B2(n10588), .A(n10587), .ZN(n10747) );
  XNOR2_X1 U7368 ( .A(n10586), .B(n7545), .ZN(n10589) );
  NAND2_X1 U7369 ( .A1(n6802), .A2(n14771), .ZN(n14774) );
  CLKBUF_X1 U7370 ( .A(n11639), .Z(n6569) );
  BUF_X4 U7371 ( .A(n11639), .Z(n6570) );
  NOR2_X1 U7372 ( .A1(n6859), .A2(n6702), .ZN(n6799) );
  OR2_X2 U7373 ( .A1(n8362), .A2(n6614), .ZN(n7376) );
  OR2_X2 U7374 ( .A1(n12601), .A2(n15550), .ZN(n11692) );
  XNOR2_X2 U7375 ( .A(n7395), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14761) );
  INV_X2 U7376 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7395) );
  OR2_X2 U7377 ( .A1(n11348), .A2(n9759), .ZN(n9496) );
  CLKBUF_X2 U7378 ( .A(n10244), .Z(n6590) );
  NAND2_X2 U7379 ( .A1(n12113), .A2(n12112), .ZN(n14645) );
  XNOR2_X2 U7380 ( .A(n13925), .B(n13410), .ZN(n13646) );
  AOI21_X2 U7381 ( .B1(n8113), .B2(n6739), .A(n11821), .ZN(n6738) );
  NAND2_X2 U7382 ( .A1(n12706), .A2(n7138), .ZN(n8113) );
  NOR2_X2 U7383 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8106), .ZN(n8169) );
  CLKBUF_X1 U7384 ( .A(n9629), .Z(n6571) );
  BUF_X2 U7385 ( .A(n9629), .Z(n6572) );
  XNOR2_X1 U7386 ( .A(n7771), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9629) );
  XNOR2_X2 U7388 ( .A(n8179), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8194) );
  NAND2_X2 U7389 ( .A1(n8214), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8179) );
  XNOR2_X2 U7390 ( .A(n7696), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7941) );
  XNOR2_X2 U7391 ( .A(n11620), .B(n11677), .ZN(n12685) );
  OAI21_X2 U7392 ( .B1(n8056), .B2(n7219), .A(n7217), .ZN(n7223) );
  INV_X2 U7393 ( .A(n6796), .ZN(n8056) );
  AND2_X1 U7394 ( .A1(n9486), .A2(n12234), .ZN(n9490) );
  INV_X1 U7395 ( .A(n12234), .ZN(n12123) );
  INV_X4 U7396 ( .A(n7170), .ZN(n12234) );
  XNOR2_X2 U7397 ( .A(n7706), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8091) );
  MUX2_X1 U7398 ( .A(n13213), .B(n13212), .S(n15613), .Z(n13214) );
  OR2_X1 U7399 ( .A1(n9099), .A2(n9098), .ZN(n7638) );
  OR2_X1 U7400 ( .A1(n9088), .A2(n9087), .ZN(n7653) );
  NAND2_X1 U7401 ( .A1(n14058), .A2(n12368), .ZN(n14117) );
  OR2_X1 U7402 ( .A1(n13709), .A2(n13710), .ZN(n13707) );
  NAND2_X1 U7403 ( .A1(n8827), .A2(n8826), .ZN(n13913) );
  NAND2_X1 U7404 ( .A1(n14130), .A2(n14129), .ZN(n7544) );
  OR2_X1 U7405 ( .A1(n13724), .A2(n8901), .ZN(n8903) );
  OAI21_X1 U7406 ( .B1(n14108), .B2(n7533), .A(n7532), .ZN(n14148) );
  NAND2_X1 U7407 ( .A1(n8895), .A2(n8894), .ZN(n11382) );
  NAND2_X1 U7408 ( .A1(n12054), .A2(n12053), .ZN(n14677) );
  OAI211_X1 U7409 ( .C1(n8705), .C2(n8375), .A(n8374), .B(n8373), .ZN(n8379)
         );
  OAI21_X1 U7410 ( .B1(n10987), .B2(n11660), .A(n11698), .ZN(n11119) );
  OR2_X1 U7411 ( .A1(n8973), .A2(n8972), .ZN(n8979) );
  INV_X1 U7412 ( .A(n11959), .ZN(n11961) );
  CLKBUF_X2 U7413 ( .A(n8108), .Z(n8072) );
  INV_X2 U7414 ( .A(n14172), .ZN(n6855) );
  INV_X1 U7415 ( .A(n14174), .ZN(n6817) );
  INV_X1 U7416 ( .A(n13514), .ZN(n6854) );
  INV_X1 U7417 ( .A(n12241), .ZN(n12178) );
  INV_X1 U7418 ( .A(n6569), .ZN(n6798) );
  NAND2_X4 U7419 ( .A1(n10035), .A2(n15091), .ZN(n12369) );
  INV_X2 U7420 ( .A(n6577), .ZN(n8613) );
  CLKBUF_X2 U7421 ( .A(P1_U4016), .Z(n6576) );
  INV_X1 U7422 ( .A(n15224), .ZN(n10712) );
  INV_X1 U7423 ( .A(n8432), .ZN(n6577) );
  NAND2_X2 U7424 ( .A1(n11682), .A2(n11841), .ZN(n8226) );
  INV_X2 U7425 ( .A(n9194), .ZN(n9057) );
  NAND2_X1 U7428 ( .A1(n8313), .A2(n8311), .ZN(n8432) );
  NAND2_X1 U7429 ( .A1(n15134), .A2(n12222), .ZN(n10032) );
  INV_X2 U7430 ( .A(n9477), .ZN(n12066) );
  NAND2_X4 U7431 ( .A1(n12302), .A2(n13279), .ZN(n9625) );
  INV_X1 U7432 ( .A(n11925), .ZN(n15134) );
  INV_X2 U7433 ( .A(n14445), .ZN(n9547) );
  MUX2_X1 U7434 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8409), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8411) );
  OR2_X1 U7435 ( .A1(n7925), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7946) );
  INV_X8 U7436 ( .A(n9681), .ZN(n11919) );
  INV_X4 U7437 ( .A(n8324), .ZN(n9681) );
  INV_X2 U7438 ( .A(n9603), .ZN(n15485) );
  NOR2_X1 U7439 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  NOR2_X1 U7440 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7301) );
  OR2_X1 U7441 ( .A1(n14616), .A2(n15199), .ZN(n6913) );
  AND2_X1 U7442 ( .A1(n14425), .A2(n14424), .ZN(n14627) );
  NAND2_X1 U7443 ( .A1(n14385), .A2(n6872), .ZN(n14423) );
  OR2_X1 U7444 ( .A1(n13918), .A2(n13917), .ZN(n13989) );
  NOR2_X1 U7445 ( .A1(n14613), .A2(n14612), .ZN(n14614) );
  CLKBUF_X1 U7446 ( .A(n12466), .Z(n12468) );
  NAND2_X1 U7447 ( .A1(n13629), .A2(n8821), .ZN(n13613) );
  NAND2_X1 U7448 ( .A1(n13631), .A2(n13630), .ZN(n13629) );
  NAND2_X1 U7449 ( .A1(n7275), .A2(n6597), .ZN(n13904) );
  NAND2_X1 U7450 ( .A1(n8797), .A2(n8796), .ZN(n13647) );
  OR2_X1 U7451 ( .A1(n13618), .A2(n8914), .ZN(n7275) );
  OAI21_X1 U7452 ( .B1(n12428), .B2(n11624), .A(n11623), .ZN(n14951) );
  NAND2_X1 U7453 ( .A1(n9296), .A2(n9295), .ZN(n11645) );
  AND2_X2 U7454 ( .A1(n11812), .A2(n11813), .ZN(n12708) );
  NAND2_X1 U7455 ( .A1(n8929), .A2(n8928), .ZN(n12691) );
  NAND2_X1 U7456 ( .A1(n8417), .A2(n8416), .ZN(n13899) );
  NAND2_X1 U7457 ( .A1(n14099), .A2(n14098), .ZN(n14097) );
  AND2_X1 U7458 ( .A1(n7226), .A2(n7225), .ZN(n11626) );
  NAND2_X1 U7459 ( .A1(n8104), .A2(n8103), .ZN(n12701) );
  NAND2_X1 U7460 ( .A1(n9149), .A2(n9148), .ZN(n9187) );
  OR2_X1 U7461 ( .A1(n12715), .A2(n12492), .ZN(n11812) );
  AOI21_X1 U7462 ( .B1(n7284), .B2(n7286), .A(n6673), .ZN(n7283) );
  NAND2_X1 U7463 ( .A1(n13464), .A2(n13327), .ZN(n13330) );
  XNOR2_X1 U7464 ( .A(n8855), .B(n8854), .ZN(n14009) );
  NAND2_X1 U7465 ( .A1(n7544), .A2(n7542), .ZN(n14052) );
  NAND2_X1 U7466 ( .A1(n12177), .A2(n12176), .ZN(n14430) );
  OR2_X1 U7467 ( .A1(n13669), .A2(n7285), .ZN(n7281) );
  NOR2_X2 U7468 ( .A1(n14630), .A2(n14461), .ZN(n14436) );
  NAND2_X1 U7469 ( .A1(n8717), .A2(n8716), .ZN(n13726) );
  MUX2_X1 U7470 ( .A(n13567), .B(n13566), .S(n13565), .Z(n13570) );
  INV_X1 U7471 ( .A(n12892), .ZN(n12757) );
  XNOR2_X1 U7472 ( .A(n8841), .B(n8840), .ZN(n14013) );
  NAND2_X1 U7473 ( .A1(n8070), .A2(n8069), .ZN(n12768) );
  NAND2_X1 U7474 ( .A1(n8815), .A2(n8814), .ZN(n13920) );
  OAI21_X1 U7475 ( .B1(n13706), .B2(n8905), .A(n8904), .ZN(n13694) );
  NAND2_X1 U7476 ( .A1(n8801), .A2(n8800), .ZN(n12124) );
  XNOR2_X1 U7477 ( .A(n7056), .B(n7055), .ZN(n14884) );
  CLKBUF_X1 U7478 ( .A(n13418), .Z(n6782) );
  NAND2_X1 U7479 ( .A1(n12309), .A2(n7639), .ZN(n6583) );
  NAND2_X1 U7480 ( .A1(n11600), .A2(n6659), .ZN(n12309) );
  NAND2_X1 U7481 ( .A1(n8770), .A2(n8769), .ZN(n13937) );
  NAND2_X1 U7482 ( .A1(n14720), .A2(n11922), .ZN(n14651) );
  AOI21_X1 U7483 ( .B1(n11473), .B2(n12593), .A(n11474), .ZN(n11507) );
  NAND2_X1 U7484 ( .A1(n12086), .A2(n12085), .ZN(n14540) );
  NAND2_X1 U7485 ( .A1(n12603), .A2(n12602), .ZN(n7053) );
  NAND2_X1 U7486 ( .A1(n7704), .A2(n7703), .ZN(n8037) );
  AND2_X1 U7487 ( .A1(n8387), .A2(n7644), .ZN(n6957) );
  NAND2_X1 U7488 ( .A1(n11333), .A2(n11332), .ZN(n11388) );
  NAND2_X1 U7489 ( .A1(n12068), .A2(n12067), .ZN(n14670) );
  NAND2_X1 U7490 ( .A1(n11135), .A2(n6661), .ZN(n11333) );
  NAND2_X1 U7491 ( .A1(n10894), .A2(n10893), .ZN(n11135) );
  NAND2_X1 U7492 ( .A1(n6941), .A2(n6725), .ZN(n7171) );
  NAND4_X1 U7493 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n12580)
         );
  NAND2_X1 U7494 ( .A1(n11214), .A2(n6848), .ZN(n11897) );
  OR2_X1 U7495 ( .A1(n10763), .A2(n10762), .ZN(n6941) );
  NAND2_X1 U7496 ( .A1(n8890), .A2(n8889), .ZN(n13848) );
  NAND2_X1 U7497 ( .A1(n6621), .A2(n6849), .ZN(n11857) );
  NAND2_X1 U7498 ( .A1(n8574), .A2(n8573), .ZN(n13845) );
  INV_X2 U7499 ( .A(n15566), .ZN(n14943) );
  AOI21_X1 U7500 ( .B1(n8620), .B2(n8361), .A(n8360), .ZN(n8362) );
  AND2_X1 U7501 ( .A1(n10286), .A2(n11959), .ZN(n10117) );
  OR2_X1 U7502 ( .A1(n10192), .A2(n10191), .ZN(n10193) );
  BUF_X1 U7503 ( .A(n9326), .Z(n9328) );
  INV_X1 U7504 ( .A(n9326), .ZN(n12440) );
  NOR2_X1 U7505 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  NAND2_X2 U7506 ( .A1(n11955), .A2(n11956), .ZN(n10279) );
  INV_X1 U7507 ( .A(n9321), .ZN(n6574) );
  NAND2_X1 U7508 ( .A1(n8510), .A2(n8509), .ZN(n15396) );
  OR2_X1 U7509 ( .A1(n15464), .A2(n10734), .ZN(n11688) );
  NAND4_X2 U7510 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n12600)
         );
  NAND4_X2 U7511 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n13513)
         );
  XNOR2_X1 U7512 ( .A(n9620), .B(n9636), .ZN(n15514) );
  NAND2_X1 U7513 ( .A1(n8959), .A2(n10721), .ZN(n9237) );
  INV_X2 U7514 ( .A(n8166), .ZN(n11637) );
  INV_X2 U7515 ( .A(n10061), .ZN(n6575) );
  INV_X2 U7516 ( .A(n8167), .ZN(n11636) );
  XNOR2_X1 U7517 ( .A(n13515), .B(n8968), .ZN(n10250) );
  NAND4_X1 U7518 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n14169)
         );
  AND2_X1 U7519 ( .A1(n9510), .A2(n9509), .ZN(n11959) );
  NOR2_X1 U7520 ( .A1(n15493), .A2(n6634), .ZN(n9620) );
  INV_X1 U7521 ( .A(n14046), .ZN(n15155) );
  CLKBUF_X1 U7522 ( .A(n14173), .Z(n6776) );
  NAND2_X1 U7523 ( .A1(n9504), .A2(n7032), .ZN(n14046) );
  NAND4_X1 U7524 ( .A1(n9472), .A2(n9471), .A3(n9470), .A4(n9469), .ZN(n14174)
         );
  NAND4_X1 U7525 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n13514)
         );
  NOR2_X2 U7526 ( .A1(n8226), .A2(n8175), .ZN(n8165) );
  INV_X2 U7527 ( .A(n11624), .ZN(n11633) );
  NAND2_X1 U7528 ( .A1(n7669), .A2(n8114), .ZN(n12673) );
  INV_X1 U7529 ( .A(n10035), .ZN(n12371) );
  INV_X4 U7530 ( .A(n9162), .ZN(n8859) );
  AND2_X1 U7531 ( .A1(n9269), .A2(n9272), .ZN(n6585) );
  INV_X4 U7532 ( .A(n9057), .ZN(n9137) );
  OAI211_X1 U7533 ( .C1(n8437), .C2(n9984), .A(n8471), .B(n8470), .ZN(n15224)
         );
  INV_X1 U7534 ( .A(n10032), .ZN(n11929) );
  NAND3_X1 U7535 ( .A1(n6991), .A2(n6990), .A3(n6992), .ZN(n11682) );
  INV_X4 U7536 ( .A(n11168), .ZN(n12223) );
  AND3_X1 U7537 ( .A1(n7175), .A2(n7173), .A3(P3_REG2_REG_3__SCAN_IN), .ZN(
        n15473) );
  INV_X2 U7538 ( .A(n8802), .ZN(n9188) );
  NAND2_X1 U7539 ( .A1(n9477), .A2(n9681), .ZN(n7170) );
  NOR2_X2 U7541 ( .A1(n11035), .A2(n10718), .ZN(n10647) );
  NAND2_X4 U7542 ( .A1(n14014), .A2(n9855), .ZN(n8437) );
  NAND2_X1 U7543 ( .A1(n9539), .A2(n9543), .ZN(n12222) );
  XNOR2_X1 U7544 ( .A(n7733), .B(P3_IR_REG_29__SCAN_IN), .ZN(n13273) );
  XNOR2_X1 U7545 ( .A(n7674), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11841) );
  NOR2_X1 U7546 ( .A1(n15476), .A2(n15618), .ZN(n15475) );
  CLKBUF_X1 U7547 ( .A(n9554), .Z(n11866) );
  OR2_X1 U7548 ( .A1(n11035), .A2(n10718), .ZN(n8960) );
  AOI21_X1 U7549 ( .B1(n9881), .B2(n14821), .A(n14822), .ZN(n15639) );
  XNOR2_X1 U7550 ( .A(n9545), .B(n9544), .ZN(n10042) );
  NAND2_X1 U7551 ( .A1(n14002), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U7552 ( .A1(n6753), .A2(n6752), .ZN(n7718) );
  NAND2_X1 U7553 ( .A1(n8253), .A2(n8274), .ZN(n11035) );
  NAND2_X1 U7554 ( .A1(n7256), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7733) );
  XNOR2_X1 U7555 ( .A(n9536), .B(n9535), .ZN(n11925) );
  MUX2_X1 U7556 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9538), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9539) );
  OAI21_X1 U7557 ( .B1(n9543), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U7558 ( .A1(n8189), .A2(n7715), .ZN(n7729) );
  NAND2_X1 U7559 ( .A1(n7679), .A2(n7678), .ZN(n7822) );
  MUX2_X1 U7560 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8251), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8253) );
  NAND2_X1 U7561 ( .A1(n7449), .A2(n7447), .ZN(n14445) );
  XNOR2_X1 U7562 ( .A(n8254), .B(n8256), .ZN(n11319) );
  OR2_X1 U7563 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  NAND2_X1 U7564 ( .A1(n9445), .A2(n6671), .ZN(n6805) );
  NAND2_X1 U7565 ( .A1(n9543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U7566 ( .A1(n14709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9446) );
  XNOR2_X1 U7567 ( .A(n9450), .B(n9449), .ZN(n14714) );
  NOR2_X1 U7568 ( .A1(n9680), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14835) );
  NAND2_X1 U7569 ( .A1(n7632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U7570 ( .A1(n9541), .A2(n9426), .ZN(n9543) );
  NAND2_X1 U7571 ( .A1(n9680), .A2(P1_U3086), .ZN(n12296) );
  AND2_X1 U7572 ( .A1(n9440), .A2(n9427), .ZN(n9435) );
  CLKBUF_X1 U7573 ( .A(n8269), .Z(n6589) );
  NOR2_X1 U7574 ( .A1(n10257), .A2(n7547), .ZN(n9440) );
  NAND2_X2 U7575 ( .A1(n9681), .A2(P1_U3086), .ZN(n12426) );
  INV_X1 U7576 ( .A(n8252), .ZN(n8250) );
  NAND2_X1 U7577 ( .A1(n8252), .A2(n8255), .ZN(n8274) );
  NOR2_X1 U7578 ( .A1(n8259), .A2(n8258), .ZN(n8269) );
  AND2_X1 U7579 ( .A1(n7046), .A2(n7045), .ZN(n7044) );
  AND2_X1 U7580 ( .A1(n6920), .A2(n6706), .ZN(n14726) );
  NAND2_X1 U7581 ( .A1(n8441), .A2(n8440), .ZN(n15228) );
  AND2_X1 U7582 ( .A1(n6828), .A2(n7656), .ZN(n7659) );
  NOR2_X2 U7583 ( .A1(n7844), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7875) );
  AND4_X1 U7584 ( .A1(n9537), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(n9432)
         );
  AND2_X1 U7585 ( .A1(n9537), .A2(n9428), .ZN(n9426) );
  OR2_X1 U7586 ( .A1(n7826), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7844) );
  AND4_X1 U7587 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n9423)
         );
  AND4_X1 U7588 ( .A1(n7800), .A2(n7816), .A3(n7657), .A4(n7837), .ZN(n7658)
         );
  NAND2_X1 U7589 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7715), .ZN(n6752) );
  AND3_X1 U7590 ( .A1(n9425), .A2(n9424), .A3(n9540), .ZN(n9537) );
  AND2_X1 U7591 ( .A1(n8260), .A2(n7507), .ZN(n6602) );
  NAND2_X1 U7592 ( .A1(n6830), .A2(n6829), .ZN(n7077) );
  NOR2_X1 U7593 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n9424) );
  INV_X1 U7594 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9535) );
  NOR2_X1 U7595 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9425) );
  NOR2_X2 U7596 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9462) );
  INV_X1 U7597 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9428) );
  INV_X4 U7598 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X2 U7599 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7308) );
  INV_X1 U7600 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9501) );
  INV_X4 U7601 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7602 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9415) );
  NOR2_X1 U7603 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9416) );
  INV_X1 U7604 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7816) );
  INV_X4 U7605 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7606 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9544) );
  INV_X1 U7607 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9692) );
  NOR2_X1 U7608 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7307) );
  INV_X1 U7609 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9540) );
  NOR2_X1 U7610 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8240) );
  INV_X1 U7611 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U7613 ( .A1(n14075), .A2(n6582), .ZN(n6579) );
  AND2_X1 U7614 ( .A1(n6579), .A2(n6580), .ZN(n12340) );
  OR2_X1 U7615 ( .A1(n6581), .A2(n12336), .ZN(n6580) );
  INV_X1 U7616 ( .A(n14084), .ZN(n6581) );
  AND2_X1 U7617 ( .A1(n14074), .A2(n14084), .ZN(n6582) );
  CLKBUF_X1 U7618 ( .A(n10752), .Z(n6584) );
  NAND2_X1 U7619 ( .A1(n12309), .A2(n7639), .ZN(n14108) );
  NOR2_X1 U7620 ( .A1(n10040), .A2(n10039), .ZN(n10066) );
  NAND3_X1 U7621 ( .A1(n9270), .A2(n6585), .A3(n9278), .ZN(n9287) );
  AND2_X1 U7622 ( .A1(n8980), .A2(n6663), .ZN(n6586) );
  INV_X1 U7623 ( .A(n13565), .ZN(n6587) );
  OR2_X1 U7624 ( .A1(n8979), .A2(n8978), .ZN(n6663) );
  NAND2_X1 U7625 ( .A1(n7325), .A2(n7324), .ZN(n8957) );
  NOR2_X2 U7626 ( .A1(n14670), .A2(n14575), .ZN(n14554) );
  NAND2_X1 U7627 ( .A1(n8572), .A2(n8246), .ZN(n6588) );
  NAND2_X1 U7628 ( .A1(n8572), .A2(n8246), .ZN(n8259) );
  OR2_X1 U7629 ( .A1(n9045), .A2(n9044), .ZN(n7650) );
  NOR2_X1 U7630 ( .A1(n9068), .A2(n9067), .ZN(n6775) );
  OAI22_X1 U7631 ( .A1(n9130), .A2(n9129), .B1(n9135), .B2(n9136), .ZN(n9146)
         );
  AOI21_X2 U7632 ( .B1(n7223), .B2(n6856), .A(n6733), .ZN(n7706) );
  XNOR2_X2 U7633 ( .A(n13330), .B(n13328), .ZN(n13360) );
  OR2_X1 U7634 ( .A1(n9081), .A2(n9080), .ZN(n6680) );
  NOR2_X2 U7635 ( .A1(n14930), .A2(n12630), .ZN(n12632) );
  NOR2_X1 U7636 ( .A1(n6588), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8252) );
  NOR2_X1 U7637 ( .A1(n7397), .A2(n7396), .ZN(n15017) );
  OAI22_X2 U7638 ( .A1(n13726), .A2(n8735), .B1(n13713), .B2(n13951), .ZN(
        n13709) );
  OAI21_X2 U7639 ( .B1(n13647), .B2(n13646), .A(n8811), .ZN(n13631) );
  NAND2_X1 U7640 ( .A1(n8519), .A2(n8518), .ZN(n10664) );
  XNOR2_X1 U7641 ( .A(n7759), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10244) );
  OAI21_X2 U7642 ( .B1(n8996), .B2(n7621), .A(n6779), .ZN(n9002) );
  NOR2_X2 U7643 ( .A1(n14584), .A2(n14682), .ZN(n7104) );
  OR2_X1 U7644 ( .A1(n8312), .A2(n8313), .ZN(n6591) );
  NOR2_X2 U7645 ( .A1(n10623), .A2(n15170), .ZN(n10626) );
  OR2_X4 U7647 ( .A1(n8312), .A2(n8313), .ZN(n8430) );
  OAI222_X1 U7648 ( .A1(n8312), .A2(P2_U3088), .B1(n14022), .B2(n12439), .C1(
        n12438), .C2(n14024), .ZN(P2_U3297) );
  NAND2_X1 U7649 ( .A1(n8312), .A2(n8313), .ZN(n8429) );
  XNOR2_X2 U7650 ( .A(n8310), .B(n14003), .ZN(n8312) );
  NAND2_X1 U7651 ( .A1(n6749), .A2(n6747), .ZN(n11703) );
  AND2_X1 U7652 ( .A1(n6748), .A2(n11702), .ZN(n6747) );
  AND2_X1 U7653 ( .A1(n11701), .A2(n11700), .ZN(n6748) );
  INV_X1 U7654 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7837) );
  INV_X1 U7655 ( .A(n13273), .ZN(n7737) );
  INV_X1 U7656 ( .A(n7738), .ZN(n7734) );
  AND2_X1 U7657 ( .A1(n6936), .A2(n6692), .ZN(n14785) );
  OR2_X1 U7658 ( .A1(n14782), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U7659 ( .A1(n12762), .A2(n8154), .ZN(n8156) );
  NOR2_X1 U7660 ( .A1(n7462), .A2(n8665), .ZN(n7461) );
  XNOR2_X1 U7661 ( .A(n12250), .B(n14379), .ZN(n14474) );
  INV_X1 U7662 ( .A(n11705), .ZN(n6744) );
  AND2_X1 U7663 ( .A1(n11703), .A2(n6842), .ZN(n6841) );
  MUX2_X1 U7664 ( .A(n14526), .B(n14540), .S(n12228), .Z(n12087) );
  AND2_X1 U7665 ( .A1(n12766), .A2(n11798), .ZN(n6840) );
  AOI21_X1 U7666 ( .B1(n7612), .B2(n7609), .A(n9119), .ZN(n7608) );
  OR2_X1 U7667 ( .A1(n12194), .A2(n12191), .ZN(n7016) );
  NAND2_X1 U7668 ( .A1(n12191), .A2(n12194), .ZN(n7018) );
  NAND2_X1 U7669 ( .A1(n14420), .A2(n7380), .ZN(n7379) );
  AND3_X1 U7670 ( .A1(n14441), .A2(n14451), .A3(n12278), .ZN(n7380) );
  OR4_X1 U7671 ( .A1(n14491), .A2(n14522), .A3(n14509), .A4(n12276), .ZN(
        n12277) );
  INV_X1 U7672 ( .A(n10966), .ZN(n7418) );
  AOI21_X1 U7673 ( .B1(n10798), .B2(n6897), .A(n10797), .ZN(n6893) );
  NAND2_X1 U7674 ( .A1(n10493), .A2(n10494), .ZN(n6897) );
  AOI21_X1 U7675 ( .B1(n7370), .B2(n7371), .A(n6678), .ZN(n7368) );
  INV_X1 U7676 ( .A(n8343), .ZN(n7371) );
  NOR2_X1 U7677 ( .A1(n11900), .A2(n11899), .ZN(n6982) );
  NAND2_X1 U7678 ( .A1(n11900), .A2(n11899), .ZN(n6983) );
  AND2_X1 U7679 ( .A1(n12476), .A2(n6976), .ZN(n6975) );
  NAND2_X1 U7680 ( .A1(n11846), .A2(n9357), .ZN(n6976) );
  NAND2_X1 U7681 ( .A1(n6961), .A2(n9320), .ZN(n9326) );
  NAND4_X1 U7682 ( .A1(n6962), .A2(n10789), .A3(n8196), .A4(n8945), .ZN(n6961)
         );
  NAND3_X1 U7683 ( .A1(n7936), .A2(n6601), .A3(n7139), .ZN(n8187) );
  AND2_X1 U7684 ( .A1(n7713), .A2(n7662), .ZN(n7139) );
  NOR2_X1 U7685 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7656) );
  NOR2_X1 U7686 ( .A1(n9124), .A2(n9125), .ZN(n9123) );
  INV_X1 U7687 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U7688 ( .A1(n13834), .A2(n9244), .ZN(n8584) );
  INV_X1 U7689 ( .A(n14019), .ZN(n8288) );
  NAND2_X1 U7690 ( .A1(n7332), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7331) );
  INV_X1 U7691 ( .A(n7333), .ZN(n7332) );
  NAND2_X1 U7692 ( .A1(n11396), .A2(n7515), .ZN(n7514) );
  INV_X1 U7693 ( .A(n11389), .ZN(n7515) );
  OR2_X1 U7694 ( .A1(n10536), .A2(n10537), .ZN(n7546) );
  OR2_X1 U7695 ( .A1(n11926), .A2(n12222), .ZN(n11927) );
  NOR2_X1 U7696 ( .A1(n11987), .A2(n15191), .ZN(n7096) );
  OR2_X1 U7697 ( .A1(n10614), .A2(n6893), .ZN(n6890) );
  NAND2_X1 U7698 ( .A1(n7388), .A2(n8856), .ZN(n9149) );
  NAND2_X1 U7699 ( .A1(n7387), .A2(n7385), .ZN(n7388) );
  NOR2_X1 U7700 ( .A1(n7386), .A2(n8854), .ZN(n7385) );
  INV_X1 U7701 ( .A(n8404), .ZN(n7386) );
  NAND2_X1 U7702 ( .A1(n9541), .A2(n9432), .ZN(n9445) );
  OR2_X1 U7703 ( .A1(n8585), .A2(n8586), .ZN(n8588) );
  CLKBUF_X1 U7704 ( .A(n8552), .Z(n8554) );
  XNOR2_X1 U7705 ( .A(n8342), .B(SI_7_), .ZN(n8521) );
  CLKBUF_X1 U7706 ( .A(n8520), .Z(n8522) );
  NOR2_X1 U7707 ( .A1(n14737), .A2(n6940), .ZN(n14755) );
  AND2_X1 U7708 ( .A1(n14738), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n6940) );
  NOR2_X1 U7709 ( .A1(n14785), .A2(n14786), .ZN(n14737) );
  NOR2_X1 U7710 ( .A1(n14744), .A2(n6795), .ZN(n14753) );
  AND2_X1 U7711 ( .A1(n14745), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n6795) );
  NOR2_X1 U7712 ( .A1(n12484), .A2(n7231), .ZN(n7230) );
  INV_X1 U7713 ( .A(n9361), .ZN(n7231) );
  INV_X1 U7714 ( .A(n11677), .ZN(n7200) );
  AND4_X1 U7715 ( .A1(n7753), .A2(n7752), .A3(n7751), .A4(n7750), .ZN(n12523)
         );
  AND4_X1 U7716 ( .A1(n7987), .A2(n7986), .A3(n7985), .A4(n7984), .ZN(n11563)
         );
  NAND2_X1 U7717 ( .A1(n12656), .A2(n7179), .ZN(n7178) );
  OR2_X1 U7718 ( .A1(n14915), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U7719 ( .A1(n7179), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7177) );
  INV_X1 U7720 ( .A(n6622), .ZN(n11624) );
  AND2_X2 U7721 ( .A1(n11818), .A2(n9290), .ZN(n12441) );
  NAND2_X1 U7722 ( .A1(n6792), .A2(n6791), .ZN(n8932) );
  AND2_X1 U7723 ( .A1(n11815), .A2(n11812), .ZN(n7138) );
  NAND2_X1 U7724 ( .A1(n12752), .A2(n8157), .ZN(n12736) );
  INV_X1 U7725 ( .A(n7124), .ZN(n7123) );
  AND2_X1 U7726 ( .A1(n7121), .A2(n12741), .ZN(n7120) );
  NAND2_X1 U7727 ( .A1(n7124), .A2(n7122), .ZN(n7121) );
  OAI21_X1 U7728 ( .B1(n12775), .B2(n8153), .A(n11655), .ZN(n12762) );
  NAND2_X1 U7729 ( .A1(n10734), .A2(n8123), .ZN(n15554) );
  AND2_X1 U7730 ( .A1(n8192), .A2(n8213), .ZN(n9899) );
  OR2_X1 U7731 ( .A1(n8183), .A2(n8198), .ZN(n8192) );
  NAND2_X1 U7732 ( .A1(n11626), .A2(n11625), .ZN(n11628) );
  NAND2_X1 U7733 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n10786), .ZN(n7703) );
  AND2_X1 U7734 ( .A1(n7839), .A2(n7850), .ZN(n10207) );
  INV_X1 U7735 ( .A(n8657), .ZN(n8299) );
  AOI21_X1 U7736 ( .B1(n6597), .B2(n8914), .A(n6655), .ZN(n7271) );
  XNOR2_X1 U7737 ( .A(n13905), .B(n13499), .ZN(n13608) );
  NAND2_X1 U7738 ( .A1(n6674), .A2(n7300), .ZN(n7297) );
  AOI21_X1 U7739 ( .B1(n7468), .B2(n7467), .A(n6654), .ZN(n7466) );
  INV_X1 U7740 ( .A(n8651), .ZN(n7468) );
  NOR2_X1 U7741 ( .A1(n8636), .A2(n7469), .ZN(n7467) );
  OR2_X1 U7742 ( .A1(n11454), .A2(n13797), .ZN(n7300) );
  NAND2_X1 U7743 ( .A1(n13800), .A2(n8618), .ZN(n11374) );
  NAND2_X1 U7744 ( .A1(n8584), .A2(n7503), .ZN(n13818) );
  NOR2_X1 U7745 ( .A1(n13815), .A2(n7504), .ZN(n7503) );
  INV_X1 U7746 ( .A(n8583), .ZN(n7504) );
  AND2_X1 U7747 ( .A1(n8866), .A2(n10173), .ZN(n13854) );
  AND2_X1 U7748 ( .A1(n7629), .A2(n8414), .ZN(n7628) );
  AND2_X1 U7749 ( .A1(n6602), .A2(n8261), .ZN(n7506) );
  INV_X1 U7750 ( .A(n8262), .ZN(n8267) );
  AOI21_X1 U7751 ( .B1(n7150), .B2(n7148), .A(n6658), .ZN(n7147) );
  INV_X1 U7752 ( .A(n7150), .ZN(n7149) );
  INV_X1 U7753 ( .A(n14352), .ZN(n6908) );
  NAND2_X1 U7754 ( .A1(n14350), .A2(n14349), .ZN(n14551) );
  NAND2_X1 U7755 ( .A1(n14567), .A2(n14566), .ZN(n14350) );
  OR2_X1 U7756 ( .A1(n14156), .A2(n14984), .ZN(n12031) );
  AND2_X1 U7757 ( .A1(n11795), .A2(n8175), .ZN(n12849) );
  NOR2_X1 U7758 ( .A1(n14927), .A2(n13194), .ZN(n14930) );
  NAND2_X1 U7759 ( .A1(n13905), .A2(n15223), .ZN(n13354) );
  OAI21_X1 U7760 ( .B1(n7490), .B2(n15313), .A(n15457), .ZN(n7488) );
  OR2_X1 U7761 ( .A1(n12124), .A2(n12123), .ZN(n12126) );
  NAND2_X1 U7762 ( .A1(n14393), .A2(n14556), .ZN(n14547) );
  INV_X1 U7763 ( .A(n8995), .ZN(n7623) );
  NOR2_X1 U7764 ( .A1(n11940), .A2(n11939), .ZN(n11941) );
  NAND2_X1 U7765 ( .A1(n11935), .A2(n12241), .ZN(n11936) );
  AND2_X1 U7766 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  NAND2_X1 U7767 ( .A1(n11947), .A2(n12241), .ZN(n11951) );
  MUX2_X1 U7768 ( .A(n11945), .B(n11944), .S(n12241), .Z(n11953) );
  NAND2_X1 U7769 ( .A1(n7031), .A2(n6633), .ZN(n11969) );
  NOR2_X1 U7770 ( .A1(n9011), .A2(n7601), .ZN(n7600) );
  INV_X1 U7771 ( .A(n9012), .ZN(n7601) );
  NAND2_X1 U7772 ( .A1(n6751), .A2(n6750), .ZN(n11699) );
  INV_X1 U7773 ( .A(n11694), .ZN(n6750) );
  OR2_X1 U7774 ( .A1(n9030), .A2(n9031), .ZN(n7624) );
  OAI21_X1 U7775 ( .B1(n9027), .B2(n9026), .A(n7626), .ZN(n7625) );
  INV_X1 U7776 ( .A(n11993), .ZN(n11996) );
  NOR2_X1 U7777 ( .A1(n6743), .A2(n11713), .ZN(n6742) );
  AND2_X1 U7778 ( .A1(n11704), .A2(n11795), .ZN(n6743) );
  INV_X1 U7779 ( .A(n7825), .ZN(n11704) );
  AND2_X1 U7780 ( .A1(n12253), .A2(n12008), .ZN(n6768) );
  NAND2_X1 U7781 ( .A1(n7026), .A2(n12114), .ZN(n7025) );
  INV_X1 U7782 ( .A(n12115), .ZN(n7026) );
  AND2_X1 U7783 ( .A1(n12128), .A2(n12129), .ZN(n7651) );
  MUX2_X1 U7784 ( .A(n14488), .B(n12250), .S(n12241), .Z(n12129) );
  INV_X1 U7785 ( .A(n9115), .ZN(n7615) );
  AOI22_X1 U7786 ( .A1(n11801), .A2(n12759), .B1(n11800), .B2(n12757), .ZN(
        n11807) );
  INV_X1 U7787 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8177) );
  AOI21_X1 U7788 ( .B1(n9116), .B2(n7605), .A(n7602), .ZN(n9124) );
  NAND2_X1 U7789 ( .A1(n7607), .A2(n7606), .ZN(n7605) );
  NAND2_X1 U7790 ( .A1(n7604), .A2(n7603), .ZN(n7602) );
  OAI21_X1 U7791 ( .B1(n10675), .B2(n7265), .A(n8888), .ZN(n7264) );
  NOR2_X1 U7792 ( .A1(n13889), .A2(n13865), .ZN(n7039) );
  INV_X1 U7793 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7631) );
  INV_X1 U7794 ( .A(n6602), .ZN(n7047) );
  NAND2_X1 U7795 ( .A1(n7017), .A2(n7016), .ZN(n7011) );
  AND2_X1 U7796 ( .A1(n7018), .A2(n7013), .ZN(n6825) );
  AOI21_X1 U7797 ( .B1(n7014), .B2(n7018), .A(n7013), .ZN(n7012) );
  INV_X1 U7798 ( .A(n11955), .ZN(n6862) );
  INV_X1 U7799 ( .A(n6949), .ZN(n6948) );
  OAI21_X1 U7800 ( .B1(n8345), .B2(n6950), .A(n8349), .ZN(n6949) );
  INV_X1 U7801 ( .A(n8347), .ZN(n6950) );
  INV_X1 U7802 ( .A(n8336), .ZN(n7366) );
  NOR2_X1 U7803 ( .A1(n14727), .A2(n14728), .ZN(n14729) );
  AOI21_X1 U7804 ( .B1(n6987), .B2(n11081), .A(n6688), .ZN(n6985) );
  AOI211_X1 U7805 ( .C1(n12441), .C2(n11822), .A(n11821), .B(n11820), .ZN(
        n11827) );
  INV_X1 U7806 ( .A(n9633), .ZN(n7085) );
  NOR2_X1 U7807 ( .A1(n7059), .A2(n7058), .ZN(n7057) );
  AOI21_X1 U7808 ( .B1(n12648), .B2(n12636), .A(n12635), .ZN(n12637) );
  AND2_X1 U7809 ( .A1(n7649), .A2(n11790), .ZN(n7118) );
  AOI21_X1 U7810 ( .B1(n8150), .B2(n7559), .A(n7558), .ZN(n7557) );
  INV_X1 U7811 ( .A(n12787), .ZN(n7558) );
  OAI21_X1 U7812 ( .B1(n11775), .B2(n7117), .A(n11785), .ZN(n7116) );
  INV_X1 U7813 ( .A(n11776), .ZN(n7117) );
  NOR2_X1 U7814 ( .A1(n7552), .A2(n12842), .ZN(n7549) );
  AND2_X1 U7815 ( .A1(n12842), .A2(n7110), .ZN(n7109) );
  NAND2_X1 U7816 ( .A1(n8145), .A2(n11762), .ZN(n7110) );
  INV_X1 U7817 ( .A(n7646), .ZN(n7583) );
  AND2_X1 U7818 ( .A1(n6695), .A2(n8144), .ZN(n7585) );
  NAND2_X1 U7819 ( .A1(n8143), .A2(n7646), .ZN(n7586) );
  NOR2_X1 U7820 ( .A1(n11725), .A2(n7571), .ZN(n7570) );
  INV_X1 U7821 ( .A(n11038), .ZN(n7571) );
  AND2_X1 U7822 ( .A1(n11728), .A2(n11727), .ZN(n11725) );
  NAND2_X1 U7823 ( .A1(n10153), .A2(n7767), .ZN(n8121) );
  INV_X1 U7824 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8185) );
  INV_X1 U7825 ( .A(n8187), .ZN(n8189) );
  NOR2_X1 U7826 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7672) );
  NOR2_X1 U7827 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n7671) );
  AND2_X1 U7828 ( .A1(n7665), .A2(n7670), .ZN(n6999) );
  NAND2_X1 U7829 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7693), .ZN(n7694) );
  OAI21_X1 U7830 ( .B1(n7903), .B2(n6714), .A(n7914), .ZN(n7210) );
  NOR2_X1 U7831 ( .A1(n6714), .A2(n7207), .ZN(n7206) );
  INV_X1 U7832 ( .A(n7688), .ZN(n7207) );
  AND2_X1 U7833 ( .A1(n6638), .A2(n7658), .ZN(n6858) );
  NAND2_X1 U7834 ( .A1(n7886), .A2(n7885), .ZN(n7689) );
  INV_X1 U7835 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7899) );
  INV_X1 U7836 ( .A(n7680), .ZN(n7215) );
  INV_X1 U7837 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6830) );
  INV_X1 U7838 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U7839 ( .A1(n7359), .A2(n7357), .ZN(n7356) );
  INV_X1 U7840 ( .A(n11877), .ZN(n7357) );
  INV_X1 U7841 ( .A(n11590), .ZN(n7345) );
  NAND2_X1 U7842 ( .A1(n13608), .A2(n7474), .ZN(n7471) );
  NAND2_X1 U7843 ( .A1(n7475), .A2(n8838), .ZN(n7474) );
  INV_X1 U7844 ( .A(n8837), .ZN(n7475) );
  OAI21_X1 U7845 ( .B1(n13657), .B2(n6959), .A(n6690), .ZN(n7285) );
  NAND2_X1 U7846 ( .A1(n7288), .A2(n8911), .ZN(n6959) );
  INV_X1 U7847 ( .A(n8782), .ZN(n7478) );
  OR2_X1 U7848 ( .A1(n13937), .A2(n8780), .ZN(n8782) );
  AND2_X1 U7849 ( .A1(n13747), .A2(n7280), .ZN(n7279) );
  NAND2_X1 U7850 ( .A1(n8899), .A2(n8900), .ZN(n7280) );
  INV_X1 U7851 ( .A(n13504), .ZN(n13374) );
  NOR2_X1 U7852 ( .A1(n13973), .A2(n7296), .ZN(n7293) );
  INV_X1 U7853 ( .A(n7298), .ZN(n7291) );
  NOR2_X1 U7854 ( .A1(n13967), .A2(n7050), .ZN(n7049) );
  INV_X1 U7855 ( .A(n7051), .ZN(n7050) );
  INV_X1 U7856 ( .A(n7269), .ZN(n7268) );
  OAI21_X1 U7857 ( .B1(n13855), .B2(n7270), .A(n13833), .ZN(n7269) );
  INV_X1 U7858 ( .A(n8891), .ZN(n7270) );
  INV_X1 U7859 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8239) );
  AND2_X1 U7860 ( .A1(n13885), .A2(n6697), .ZN(n13825) );
  INV_X1 U7861 ( .A(n15435), .ZN(n7036) );
  NOR2_X1 U7862 ( .A1(n7047), .A2(n7630), .ZN(n7045) );
  INV_X1 U7863 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8257) );
  INV_X1 U7864 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8260) );
  INV_X1 U7865 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8256) );
  INV_X1 U7866 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U7867 ( .A1(n8236), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U7868 ( .A1(n7306), .A2(n7307), .ZN(n7303) );
  NOR2_X1 U7869 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7306) );
  NAND2_X1 U7870 ( .A1(n7378), .A2(n6636), .ZN(n12281) );
  INV_X1 U7871 ( .A(n12282), .ZN(n7381) );
  NAND2_X1 U7872 ( .A1(n11871), .A2(n14714), .ZN(n7654) );
  NAND2_X1 U7873 ( .A1(n7101), .A2(n14623), .ZN(n7100) );
  NOR2_X1 U7874 ( .A1(n12279), .A2(n7100), .ZN(n7099) );
  NOR2_X1 U7875 ( .A1(n14474), .A2(n7415), .ZN(n7414) );
  INV_X1 U7876 ( .A(n14358), .ZN(n7415) );
  NOR2_X1 U7877 ( .A1(n14553), .A2(n7153), .ZN(n7152) );
  INV_X1 U7878 ( .A(n14371), .ZN(n7153) );
  NOR2_X1 U7879 ( .A1(n14346), .A2(n7428), .ZN(n7427) );
  INV_X1 U7880 ( .A(n12031), .ZN(n7428) );
  NAND2_X1 U7881 ( .A1(n12272), .A2(n11430), .ZN(n7156) );
  NOR2_X1 U7882 ( .A1(n12253), .A2(n7158), .ZN(n7157) );
  INV_X1 U7883 ( .A(n11362), .ZN(n7158) );
  OAI21_X1 U7884 ( .B1(n7419), .B2(n7418), .A(n12267), .ZN(n7417) );
  NOR2_X1 U7885 ( .A1(n10902), .A2(n7418), .ZN(n6888) );
  NOR2_X1 U7886 ( .A1(n10819), .A2(n7420), .ZN(n7419) );
  INV_X1 U7887 ( .A(n10805), .ZN(n7420) );
  INV_X1 U7888 ( .A(n6893), .ZN(n6892) );
  NAND2_X1 U7889 ( .A1(n14529), .A2(n14651), .ZN(n14511) );
  NAND2_X1 U7890 ( .A1(n12017), .A2(n11436), .ZN(n11529) );
  INV_X1 U7891 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7432) );
  INV_X1 U7892 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9458) );
  INV_X1 U7893 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U7894 ( .A1(n8393), .A2(n8394), .ZN(n7390) );
  INV_X1 U7895 ( .A(n8378), .ZN(n6952) );
  NOR2_X1 U7896 ( .A1(n8381), .A2(SI_20_), .ZN(n6955) );
  INV_X1 U7897 ( .A(n8736), .ZN(n8381) );
  INV_X1 U7898 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9419) );
  AND2_X1 U7899 ( .A1(n8652), .A2(n7377), .ZN(n7375) );
  INV_X1 U7900 ( .A(n8603), .ZN(n7374) );
  XNOR2_X1 U7901 ( .A(n8344), .B(SI_8_), .ZN(n8537) );
  NAND2_X1 U7902 ( .A1(n6918), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14723) );
  OAI21_X1 U7903 ( .B1(n14723), .B2(n14761), .A(n7394), .ZN(n7393) );
  NAND2_X1 U7904 ( .A1(n14724), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7394) );
  XNOR2_X1 U7905 ( .A(n14729), .B(n7413), .ZN(n14757) );
  INV_X1 U7906 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14734) );
  AND2_X1 U7907 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14792), .ZN(n14741) );
  INV_X1 U7908 ( .A(n6938), .ZN(n14740) );
  NAND2_X1 U7909 ( .A1(n14859), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6925) );
  INV_X1 U7910 ( .A(n14859), .ZN(n6926) );
  NAND2_X1 U7911 ( .A1(n6719), .A2(n6978), .ZN(n6977) );
  INV_X1 U7912 ( .A(n6982), .ZN(n6978) );
  OR2_X1 U7913 ( .A1(n10791), .A2(n10928), .ZN(n9335) );
  NAND2_X1 U7914 ( .A1(n6970), .A2(n6968), .ZN(n7232) );
  AND2_X1 U7915 ( .A1(n12536), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U7916 ( .A1(n6971), .A2(n6973), .ZN(n6969) );
  AOI21_X1 U7917 ( .B1(n12507), .B2(n7254), .A(n6681), .ZN(n7253) );
  INV_X1 U7918 ( .A(n9351), .ZN(n7254) );
  NAND2_X1 U7919 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  INV_X1 U7920 ( .A(n9650), .ZN(n6965) );
  AOI21_X1 U7921 ( .B1(n9335), .B2(n7243), .A(n7242), .ZN(n7241) );
  INV_X1 U7922 ( .A(n10923), .ZN(n7242) );
  INV_X1 U7923 ( .A(n10791), .ZN(n7243) );
  INV_X1 U7924 ( .A(n9335), .ZN(n7244) );
  OR2_X1 U7925 ( .A1(n11080), .A2(n11081), .ZN(n6988) );
  NAND2_X1 U7926 ( .A1(n10153), .A2(n10349), .ZN(n11685) );
  OR2_X1 U7927 ( .A1(n9342), .A2(n9341), .ZN(n11473) );
  AND2_X1 U7928 ( .A1(n9342), .A2(n9341), .ZN(n11474) );
  INV_X1 U7929 ( .A(n8121), .ZN(n10294) );
  INV_X1 U7930 ( .A(n7253), .ZN(n7251) );
  INV_X1 U7931 ( .A(n12507), .ZN(n7255) );
  XNOR2_X1 U7932 ( .A(n10292), .B(n15585), .ZN(n9331) );
  AND2_X1 U7933 ( .A1(n12555), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U7934 ( .A1(n7236), .A2(n9382), .ZN(n7235) );
  NAND2_X1 U7935 ( .A1(n10789), .A2(n8945), .ZN(n11836) );
  INV_X1 U7936 ( .A(n11831), .ZN(n6845) );
  OAI21_X1 U7937 ( .B1(n6598), .B2(n11649), .A(n11830), .ZN(n11650) );
  NAND2_X1 U7938 ( .A1(n8213), .A2(n8212), .ZN(n9594) );
  AND4_X1 U7939 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(n12567)
         );
  AND4_X1 U7940 ( .A1(n7930), .A2(n7929), .A3(n7928), .A4(n7927), .ZN(n11517)
         );
  NAND4_X1 U7941 ( .A1(n7758), .A2(n7757), .A3(n7756), .A4(n7755), .ZN(n15464)
         );
  OR2_X1 U7942 ( .A1(n6570), .A2(n7754), .ZN(n7758) );
  OR2_X1 U7943 ( .A1(n8082), .A2(n10744), .ZN(n7755) );
  NAND2_X1 U7944 ( .A1(n6572), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7087) );
  OR2_X1 U7945 ( .A1(n6572), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7086) );
  NOR2_X1 U7946 ( .A1(n15517), .A2(n15622), .ZN(n15516) );
  OAI21_X1 U7947 ( .B1(n7189), .B2(n15514), .A(n7188), .ZN(n10192) );
  OR2_X1 U7948 ( .A1(n9622), .A2(n15515), .ZN(n7189) );
  NAND2_X1 U7949 ( .A1(n9621), .A2(n7193), .ZN(n7188) );
  NAND2_X1 U7950 ( .A1(n7190), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7192) );
  INV_X1 U7951 ( .A(n15514), .ZN(n7190) );
  AND2_X1 U7952 ( .A1(n10945), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7089) );
  XNOR2_X1 U7953 ( .A(n7053), .B(n15530), .ZN(n15533) );
  AND2_X1 U7954 ( .A1(n7183), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7181) );
  NOR2_X1 U7955 ( .A1(n15533), .A2(n15534), .ZN(n15532) );
  NAND2_X1 U7956 ( .A1(n6943), .A2(n6942), .ZN(n14892) );
  INV_X1 U7957 ( .A(n14894), .ZN(n6942) );
  INV_X1 U7958 ( .A(n6738), .ZN(n11620) );
  INV_X1 U7959 ( .A(n11819), .ZN(n6739) );
  INV_X1 U7960 ( .A(n12445), .ZN(n12688) );
  NAND2_X1 U7961 ( .A1(n8163), .A2(n11815), .ZN(n6790) );
  NAND2_X1 U7962 ( .A1(n12718), .A2(n8159), .ZN(n12709) );
  AND2_X1 U7963 ( .A1(n11802), .A2(n11679), .ZN(n7125) );
  OR2_X1 U7964 ( .A1(n7126), .A2(n8090), .ZN(n7124) );
  AND2_X1 U7965 ( .A1(n12759), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U7966 ( .A1(n8077), .A2(n11679), .ZN(n7127) );
  NAND2_X1 U7967 ( .A1(n8156), .A2(n7553), .ZN(n12752) );
  INV_X1 U7968 ( .A(n8155), .ZN(n7554) );
  CLKBUF_X1 U7969 ( .A(n12767), .Z(n6787) );
  NAND2_X1 U7970 ( .A1(n12790), .A2(n8152), .ZN(n12775) );
  AND2_X1 U7971 ( .A1(n11655), .A2(n11654), .ZN(n12779) );
  NAND2_X1 U7972 ( .A1(n12844), .A2(n8148), .ZN(n12829) );
  NAND2_X1 U7973 ( .A1(n12862), .A2(n8147), .ZN(n12846) );
  NAND2_X1 U7974 ( .A1(n12846), .A2(n12845), .ZN(n12844) );
  CLKBUF_X1 U7975 ( .A(n12867), .Z(n6786) );
  NAND2_X1 U7976 ( .A1(n6786), .A2(n12866), .ZN(n12865) );
  NAND2_X1 U7977 ( .A1(n8138), .A2(n7570), .ZN(n7569) );
  OAI21_X1 U7978 ( .B1(n11040), .B2(n7873), .A(n7874), .ZN(n11093) );
  INV_X1 U7979 ( .A(n11725), .ZN(n11092) );
  NOR2_X1 U7980 ( .A1(n8135), .A2(n7563), .ZN(n7562) );
  INV_X1 U7981 ( .A(n8130), .ZN(n7563) );
  AND2_X1 U7982 ( .A1(n11715), .A2(n11714), .ZN(n11708) );
  AND2_X1 U7983 ( .A1(n10877), .A2(n10874), .ZN(n10875) );
  AND3_X1 U7984 ( .A1(n7804), .A2(n7803), .A3(n7802), .ZN(n10413) );
  OR2_X1 U7985 ( .A1(n15461), .A2(n15577), .ZN(n11693) );
  NAND2_X1 U7986 ( .A1(n8120), .A2(n8227), .ZN(n11097) );
  OR2_X1 U7987 ( .A1(n11682), .A2(n11841), .ZN(n15606) );
  OR2_X1 U7988 ( .A1(n11097), .A2(n15611), .ZN(n15600) );
  NOR2_X1 U7989 ( .A1(n11833), .A2(n11841), .ZN(n15611) );
  INV_X1 U7990 ( .A(n15606), .ZN(n14950) );
  NAND2_X1 U7991 ( .A1(n9899), .A2(n8193), .ZN(n6962) );
  NAND2_X1 U7992 ( .A1(n14713), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7225) );
  NAND2_X1 U7993 ( .A1(n8181), .A2(n8180), .ZN(n8184) );
  NAND2_X1 U7994 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11034), .ZN(n7224) );
  INV_X1 U7995 ( .A(n6993), .ZN(n6992) );
  OR2_X1 U7996 ( .A1(n7666), .A2(n6995), .ZN(n6991) );
  NAND2_X1 U7997 ( .A1(n7666), .A2(n6994), .ZN(n6990) );
  OAI21_X1 U7998 ( .B1(n8048), .B2(n10872), .A(n6683), .ZN(n6796) );
  NAND2_X1 U7999 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U8000 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n6832), .ZN(n6831) );
  XNOR2_X1 U8001 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7903) );
  NAND2_X1 U8002 ( .A1(n7689), .A2(n7688), .ZN(n7904) );
  XNOR2_X1 U8003 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7820) );
  INV_X1 U8004 ( .A(n7659), .ZN(n7799) );
  NOR2_X1 U8005 ( .A1(n11497), .A2(n7349), .ZN(n7348) );
  INV_X1 U8006 ( .A(n11495), .ZN(n7349) );
  NAND2_X1 U8007 ( .A1(n13399), .A2(n13337), .ZN(n7319) );
  OR2_X1 U8008 ( .A1(n6782), .A2(n13419), .ZN(n13416) );
  NAND3_X1 U8009 ( .A1(n13312), .A2(n13313), .A3(n7362), .ZN(n13455) );
  AND2_X1 U8010 ( .A1(n13459), .A2(n13370), .ZN(n7362) );
  OR2_X1 U8011 ( .A1(n8696), .A2(n8300), .ZN(n8710) );
  NAND2_X1 U8012 ( .A1(n13419), .A2(n13300), .ZN(n7343) );
  INV_X1 U8013 ( .A(n6593), .ZN(n9159) );
  NOR2_X1 U8014 ( .A1(n15249), .A2(n15248), .ZN(n15247) );
  NAND2_X1 U8015 ( .A1(n15292), .A2(n11008), .ZN(n11009) );
  AND2_X1 U8016 ( .A1(n13535), .A2(n13534), .ZN(n13536) );
  NAND2_X1 U8017 ( .A1(n13536), .A2(n13539), .ZN(n6813) );
  NAND2_X1 U8018 ( .A1(n9157), .A2(n9156), .ZN(n13571) );
  NAND2_X1 U8019 ( .A1(n13613), .A2(n8837), .ZN(n7473) );
  NAND2_X1 U8020 ( .A1(n7274), .A2(n13411), .ZN(n7273) );
  INV_X1 U8021 ( .A(n7285), .ZN(n7286) );
  OR2_X1 U8022 ( .A1(n13669), .A2(n8911), .ZN(n7289) );
  NAND2_X1 U8023 ( .A1(n8787), .A2(n8786), .ZN(n13673) );
  NAND2_X1 U8024 ( .A1(n13670), .A2(n8920), .ZN(n13671) );
  AND2_X1 U8025 ( .A1(n7482), .A2(n8765), .ZN(n7481) );
  INV_X1 U8026 ( .A(n13679), .ZN(n7482) );
  NAND2_X1 U8027 ( .A1(n13696), .A2(n8764), .ZN(n7483) );
  NAND2_X1 U8028 ( .A1(n7483), .A2(n8765), .ZN(n13680) );
  OR2_X1 U8029 ( .A1(n8756), .A2(n13395), .ZN(n8772) );
  NOR2_X1 U8030 ( .A1(n13754), .A2(n13957), .ZN(n13729) );
  AOI21_X1 U8031 ( .B1(n7498), .B2(n7497), .A(n6672), .ZN(n7496) );
  INV_X1 U8032 ( .A(n6625), .ZN(n7497) );
  NAND2_X1 U8033 ( .A1(n13765), .A2(n7498), .ZN(n7495) );
  NAND2_X1 U8034 ( .A1(n7500), .A2(n6625), .ZN(n7499) );
  INV_X1 U8035 ( .A(n13765), .ZN(n7500) );
  NOR2_X1 U8036 ( .A1(n8896), .A2(n7299), .ZN(n7298) );
  INV_X1 U8037 ( .A(n7300), .ZN(n7299) );
  NAND2_X1 U8038 ( .A1(n13813), .A2(n8892), .ZN(n13796) );
  NAND2_X1 U8039 ( .A1(n13818), .A2(n6610), .ZN(n13800) );
  INV_X1 U8040 ( .A(n9244), .ZN(n13833) );
  NAND2_X1 U8041 ( .A1(n13848), .A2(n13855), .ZN(n13850) );
  NOR2_X1 U8042 ( .A1(n15322), .A2(n15224), .ZN(n10701) );
  OR2_X1 U8043 ( .A1(n8802), .A2(n9707), .ZN(n8459) );
  NAND2_X1 U8044 ( .A1(n8446), .A2(n8445), .ZN(n15311) );
  OR2_X1 U8045 ( .A1(n15321), .A2(n15318), .ZN(n15322) );
  AND2_X1 U8046 ( .A1(n11319), .A2(n11035), .ZN(n10719) );
  NAND2_X1 U8047 ( .A1(n8858), .A2(n8857), .ZN(n12429) );
  XNOR2_X1 U8048 ( .A(n8917), .B(n8864), .ZN(n12434) );
  NAND2_X1 U8049 ( .A1(n8656), .A2(n8655), .ZN(n13981) );
  NAND2_X1 U8050 ( .A1(n10181), .A2(n10719), .ZN(n15428) );
  INV_X1 U8051 ( .A(n8410), .ZN(n8413) );
  NAND2_X1 U8052 ( .A1(n8677), .A2(n7329), .ZN(n7324) );
  NAND2_X1 U8053 ( .A1(n7328), .A2(n7327), .ZN(n7326) );
  INV_X1 U8054 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8478) );
  NOR2_X1 U8055 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7305) );
  AND2_X1 U8056 ( .A1(n10053), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9584) );
  AND2_X1 U8057 ( .A1(n14139), .A2(n7529), .ZN(n7528) );
  OR2_X1 U8058 ( .A1(n14068), .A2(n7530), .ZN(n7529) );
  INV_X1 U8059 ( .A(n12398), .ZN(n7530) );
  AND2_X1 U8060 ( .A1(n11388), .A2(n11387), .ZN(n7518) );
  NAND2_X1 U8061 ( .A1(n11390), .A2(n11389), .ZN(n7513) );
  NAND2_X1 U8062 ( .A1(n14097), .A2(n6660), .ZN(n14058) );
  AND2_X1 U8063 ( .A1(n14036), .A2(n7522), .ZN(n7521) );
  NAND2_X1 U8064 ( .A1(n7523), .A2(n12377), .ZN(n7522) );
  INV_X1 U8065 ( .A(n14118), .ZN(n7523) );
  INV_X1 U8066 ( .A(n7514), .ZN(n7509) );
  OAI21_X1 U8067 ( .B1(n7514), .B2(n11387), .A(n7636), .ZN(n7511) );
  OR2_X1 U8068 ( .A1(n11577), .A2(n11576), .ZN(n7636) );
  NAND2_X1 U8069 ( .A1(n11580), .A2(n11579), .ZN(n11600) );
  AOI21_X1 U8070 ( .B1(n7534), .B2(n7537), .A(n6600), .ZN(n7532) );
  INV_X1 U8071 ( .A(n7534), .ZN(n7533) );
  NAND2_X1 U8072 ( .A1(n7531), .A2(n6834), .ZN(n14147) );
  AND2_X1 U8073 ( .A1(n7534), .A2(n6600), .ZN(n6834) );
  XNOR2_X1 U8074 ( .A(n14336), .B(n7382), .ZN(n12282) );
  INV_X1 U8075 ( .A(n14335), .ZN(n7382) );
  AND2_X1 U8076 ( .A1(n7005), .A2(n7004), .ZN(n12245) );
  INV_X1 U8077 ( .A(n12219), .ZN(n12199) );
  INV_X1 U8079 ( .A(n12149), .ZN(n12218) );
  NOR2_X1 U8080 ( .A1(n10304), .A2(n7453), .ZN(n7448) );
  INV_X1 U8081 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U8082 ( .A1(n14485), .A2(n7414), .ZN(n14471) );
  AND2_X1 U8083 ( .A1(n14360), .A2(n12249), .ZN(n14451) );
  AND2_X1 U8084 ( .A1(n14546), .A2(n14373), .ZN(n7150) );
  NAND2_X1 U8085 ( .A1(n14372), .A2(n7152), .ZN(n7151) );
  OR2_X1 U8086 ( .A1(n12084), .A2(n12123), .ZN(n12086) );
  INV_X1 U8087 ( .A(n14551), .ZN(n6910) );
  OR2_X1 U8088 ( .A1(n11538), .A2(n11537), .ZN(n12069) );
  NAND2_X1 U8089 ( .A1(n7426), .A2(n14345), .ZN(n14590) );
  AND2_X1 U8090 ( .A1(n7429), .A2(n14345), .ZN(n7425) );
  INV_X1 U8091 ( .A(n14589), .ZN(n7429) );
  NAND2_X1 U8092 ( .A1(n11530), .A2(n7427), .ZN(n7426) );
  NAND2_X1 U8093 ( .A1(n11529), .A2(n11532), .ZN(n11530) );
  NAND2_X1 U8094 ( .A1(n11363), .A2(n7157), .ZN(n11431) );
  NAND2_X1 U8095 ( .A1(n10905), .A2(n7419), .ZN(n10967) );
  NAND2_X1 U8096 ( .A1(n6890), .A2(n6886), .ZN(n10905) );
  NOR2_X1 U8097 ( .A1(n6887), .A2(n10902), .ZN(n6886) );
  INV_X1 U8098 ( .A(n6889), .ZN(n6887) );
  NAND2_X1 U8099 ( .A1(n10489), .A2(n10488), .ZN(n10614) );
  INV_X1 U8100 ( .A(n10911), .ZN(n15084) );
  CLKBUF_X2 U8101 ( .A(n9477), .Z(n11922) );
  NAND2_X1 U8102 ( .A1(n6689), .A2(n6905), .ZN(n14523) );
  NAND2_X1 U8103 ( .A1(n6907), .A2(n14551), .ZN(n6905) );
  NAND2_X1 U8104 ( .A1(n8386), .A2(SI_22_), .ZN(n8387) );
  OR2_X1 U8105 ( .A1(n11920), .A2(n8766), .ZN(n8768) );
  NAND2_X1 U8106 ( .A1(n8387), .A2(n6762), .ZN(n11920) );
  OR2_X1 U8107 ( .A1(n8386), .A2(SI_22_), .ZN(n6762) );
  OR2_X1 U8108 ( .A1(n6956), .A2(n10554), .ZN(n8382) );
  NAND2_X1 U8109 ( .A1(n6956), .A2(n10554), .ZN(n8380) );
  INV_X1 U8110 ( .A(n8382), .ZN(n7383) );
  NAND2_X1 U8111 ( .A1(n8380), .A2(n8381), .ZN(n7384) );
  AND4_X1 U8112 ( .A1(n9502), .A2(n9423), .A3(n15648), .A4(n9540), .ZN(n10301)
         );
  OR2_X1 U8113 ( .A1(n10005), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n10006) );
  INV_X1 U8114 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U8115 ( .A1(n8588), .A2(n8354), .ZN(n8604) );
  NAND2_X1 U8116 ( .A1(n6947), .A2(n8347), .ZN(n8571) );
  NAND2_X1 U8117 ( .A1(n8554), .A2(n8345), .ZN(n6947) );
  INV_X1 U8118 ( .A(n14723), .ZN(n14762) );
  XNOR2_X1 U8119 ( .A(n14757), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14758) );
  NOR2_X1 U8120 ( .A1(n14775), .A2(n14776), .ZN(n14777) );
  NAND2_X1 U8121 ( .A1(n7391), .A2(n14789), .ZN(n14791) );
  NAND2_X1 U8122 ( .A1(n14841), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7391) );
  XNOR2_X1 U8123 ( .A(n6938), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14792) );
  OAI21_X1 U8124 ( .B1(n15016), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6644), .ZN(
        n7397) );
  OAI22_X1 U8125 ( .A1(n14753), .A2(n14746), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n15528), .ZN(n14809) );
  XNOR2_X1 U8126 ( .A(n9329), .B(n15461), .ZN(n9652) );
  NAND2_X1 U8127 ( .A1(n6974), .A2(n9357), .ZN(n12475) );
  OR2_X1 U8128 ( .A1(n11845), .A2(n11846), .ZN(n6974) );
  INV_X1 U8129 ( .A(n8122), .ZN(n10734) );
  OAI211_X1 U8130 ( .C1(n7132), .C2(n7131), .A(n7133), .B(n7130), .ZN(n8122)
         );
  OR2_X1 U8131 ( .A1(n12302), .A2(n7136), .ZN(n7130) );
  NAND2_X1 U8132 ( .A1(n7238), .A2(n12499), .ZN(n12496) );
  NAND2_X1 U8133 ( .A1(n10410), .A2(n7246), .ZN(n10546) );
  NAND2_X1 U8134 ( .A1(n9330), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U8135 ( .A1(n6966), .A2(n6963), .ZN(n10410) );
  AND2_X1 U8136 ( .A1(n6639), .A2(n10412), .ZN(n6963) );
  NAND2_X1 U8137 ( .A1(n6967), .A2(n6971), .ZN(n12535) );
  OR2_X1 U8138 ( .A1(n11845), .A2(n6973), .ZN(n6967) );
  AND2_X1 U8139 ( .A1(n9594), .A2(n10151), .ZN(n11839) );
  OR3_X1 U8140 ( .A1(n8035), .A2(n8034), .A3(n8033), .ZN(n12830) );
  OAI22_X1 U8141 ( .A1(n15491), .A2(n15490), .B1(n9606), .B2(n15504), .ZN(
        n15510) );
  NOR2_X1 U8142 ( .A1(n10194), .A2(n10981), .ZN(n10321) );
  INV_X1 U8143 ( .A(n7171), .ZN(n11050) );
  NOR2_X1 U8144 ( .A1(n14914), .A2(n12656), .ZN(n12659) );
  AOI21_X1 U8145 ( .B1(n6758), .B2(n6757), .A(n14920), .ZN(n12645) );
  NAND2_X1 U8146 ( .A1(n12643), .A2(n12644), .ZN(n6757) );
  INV_X1 U8147 ( .A(n12665), .ZN(n6758) );
  INV_X1 U8148 ( .A(n15547), .ZN(n7196) );
  NOR2_X1 U8149 ( .A1(n15541), .A2(n6734), .ZN(n7065) );
  NOR2_X1 U8150 ( .A1(n6732), .A2(n15541), .ZN(n7069) );
  NAND2_X1 U8151 ( .A1(n14929), .A2(n7068), .ZN(n7067) );
  INV_X1 U8152 ( .A(n7070), .ZN(n7068) );
  OAI21_X1 U8153 ( .B1(n7072), .B2(n7076), .A(n7071), .ZN(n7070) );
  NAND2_X1 U8154 ( .A1(n7076), .A2(n12664), .ZN(n7071) );
  AND2_X1 U8155 ( .A1(P3_U3897), .A2(n12302), .ZN(n15538) );
  XNOR2_X1 U8156 ( .A(n8930), .B(n12441), .ZN(n12692) );
  OAI21_X1 U8157 ( .B1(n8935), .B2(n6628), .A(n8941), .ZN(n8942) );
  AND3_X1 U8158 ( .A1(n7842), .A2(n7841), .A3(n7840), .ZN(n15589) );
  AND2_X1 U8159 ( .A1(n15566), .A2(n15565), .ZN(n12872) );
  INV_X1 U8160 ( .A(n14938), .ZN(n15553) );
  INV_X1 U8161 ( .A(n12870), .ZN(n14944) );
  NAND2_X1 U8162 ( .A1(n15631), .A2(n14950), .ZN(n13211) );
  NAND2_X1 U8163 ( .A1(n15613), .A2(n14950), .ZN(n13263) );
  INV_X1 U8164 ( .A(n7315), .ZN(n7314) );
  INV_X1 U8165 ( .A(n13382), .ZN(n13356) );
  INV_X1 U8166 ( .A(n13632), .ZN(n13410) );
  NAND2_X1 U8167 ( .A1(n10559), .A2(n11859), .ZN(n11865) );
  OAI211_X1 U8168 ( .C1(n8437), .C2(n9955), .A(n8484), .B(n8483), .ZN(n15383)
         );
  NAND2_X1 U8169 ( .A1(n8742), .A2(n8741), .ZN(n13948) );
  NAND2_X1 U8170 ( .A1(n8628), .A2(n8627), .ZN(n11454) );
  NAND2_X1 U8171 ( .A1(n8820), .A2(n8819), .ZN(n13500) );
  NAND2_X1 U8172 ( .A1(n8794), .A2(n8793), .ZN(n13466) );
  INV_X1 U8173 ( .A(n12434), .ZN(n6820) );
  NAND2_X1 U8174 ( .A1(n14013), .A2(n9188), .ZN(n8843) );
  NAND2_X1 U8175 ( .A1(n8643), .A2(n8642), .ZN(n13792) );
  NAND2_X1 U8176 ( .A1(n13883), .A2(n10657), .ZN(n14957) );
  XNOR2_X1 U8177 ( .A(n6772), .B(n8864), .ZN(n7491) );
  NAND2_X1 U8178 ( .A1(n6774), .A2(n13498), .ZN(n6773) );
  INV_X1 U8179 ( .A(n8873), .ZN(n7490) );
  AOI21_X1 U8180 ( .B1(n7491), .B2(n15313), .A(n7490), .ZN(n12437) );
  NAND2_X1 U8181 ( .A1(n8294), .A2(n8293), .ZN(n15366) );
  INV_X1 U8182 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14003) );
  NAND2_X1 U8183 ( .A1(n10492), .A2(n10491), .ZN(n15170) );
  NAND2_X1 U8184 ( .A1(n7033), .A2(n12234), .ZN(n7032) );
  INV_X1 U8185 ( .A(n9702), .ZN(n7033) );
  NOR2_X1 U8186 ( .A1(n14050), .A2(n7543), .ZN(n7542) );
  INV_X1 U8187 ( .A(n12347), .ZN(n7543) );
  NAND2_X1 U8188 ( .A1(n12024), .A2(n12023), .ZN(n14682) );
  NAND2_X1 U8189 ( .A1(n11434), .A2(n11433), .ZN(n14156) );
  AND2_X1 U8190 ( .A1(n12237), .A2(n14190), .ZN(n14569) );
  XNOR2_X1 U8191 ( .A(n6808), .B(n6807), .ZN(n14607) );
  NAND2_X1 U8192 ( .A1(n7161), .A2(n7159), .ZN(n6808) );
  NAND2_X1 U8193 ( .A1(n7160), .A2(n6632), .ZN(n7159) );
  AOI21_X1 U8194 ( .B1(n14617), .B2(n15094), .A(n14415), .ZN(n6811) );
  AOI21_X1 U8195 ( .B1(n14408), .B2(n6917), .A(n14407), .ZN(n14620) );
  NAND2_X1 U8196 ( .A1(n10304), .A2(n7452), .ZN(n7449) );
  NOR2_X1 U8197 ( .A1(n7448), .A2(n7450), .ZN(n7447) );
  NAND2_X1 U8198 ( .A1(n7455), .A2(n7451), .ZN(n7450) );
  NAND2_X1 U8199 ( .A1(n7146), .A2(n7145), .ZN(n14468) );
  AND2_X1 U8200 ( .A1(n7146), .A2(n6624), .ZN(n14467) );
  NAND2_X1 U8201 ( .A1(n10912), .A2(n11337), .ZN(n10821) );
  OR2_X1 U8202 ( .A1(n15098), .A2(n10363), .ZN(n14601) );
  XNOR2_X1 U8203 ( .A(n6756), .B(n6807), .ZN(n14615) );
  NAND2_X1 U8204 ( .A1(n6867), .A2(n6869), .ZN(n6756) );
  OAI21_X1 U8205 ( .B1(n14614), .B2(n15199), .A(n6915), .ZN(n6912) );
  OR2_X1 U8206 ( .A1(n15200), .A2(n6916), .ZN(n6915) );
  INV_X1 U8207 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6916) );
  AND2_X1 U8208 ( .A1(n14791), .A2(n14790), .ZN(n14842) );
  NOR2_X1 U8209 ( .A1(n14790), .A2(n14791), .ZN(n14843) );
  INV_X1 U8210 ( .A(n14843), .ZN(n7408) );
  XNOR2_X1 U8211 ( .A(n14804), .B(n14803), .ZN(n15016) );
  NAND2_X1 U8212 ( .A1(n6935), .A2(n6620), .ZN(n6931) );
  AOI21_X1 U8213 ( .B1(n6931), .B2(n6612), .A(n6929), .ZN(n15024) );
  NAND2_X1 U8214 ( .A1(n6933), .A2(n6930), .ZN(n6929) );
  INV_X1 U8215 ( .A(n6642), .ZN(n6930) );
  OR2_X1 U8216 ( .A1(n15024), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U8217 ( .A1(n6804), .A2(n6642), .ZN(n7403) );
  INV_X1 U8218 ( .A(n14812), .ZN(n6804) );
  OAI21_X1 U8219 ( .B1(n6932), .B2(n15018), .A(n6612), .ZN(n14812) );
  NAND2_X1 U8220 ( .A1(n6620), .A2(n6933), .ZN(n6932) );
  AOI21_X1 U8221 ( .B1(n7400), .B2(n7399), .A(P2_ADDR_REG_16__SCAN_IN), .ZN(
        n7402) );
  AND2_X1 U8222 ( .A1(n7403), .A2(n15029), .ZN(n7399) );
  NAND2_X1 U8223 ( .A1(n11933), .A2(n11932), .ZN(n11937) );
  NOR2_X1 U8224 ( .A1(n11931), .A2(n12241), .ZN(n11932) );
  INV_X1 U8225 ( .A(n11928), .ZN(n11933) );
  AND2_X1 U8226 ( .A1(n11930), .A2(n11929), .ZN(n11931) );
  OR2_X1 U8227 ( .A1(n8994), .A2(n8995), .ZN(n6779) );
  NOR2_X1 U8228 ( .A1(n7623), .A2(n7622), .ZN(n7621) );
  NAND2_X1 U8229 ( .A1(n11962), .A2(n11963), .ZN(n7030) );
  NAND2_X1 U8230 ( .A1(n7436), .A2(n7435), .ZN(n11977) );
  OR2_X1 U8231 ( .A1(n11974), .A2(n7437), .ZN(n7435) );
  INV_X1 U8232 ( .A(n7599), .ZN(n7598) );
  AOI21_X1 U8233 ( .B1(n7600), .B2(n6595), .A(n6675), .ZN(n7599) );
  NAND2_X1 U8234 ( .A1(n9030), .A2(n9031), .ZN(n7626) );
  NOR2_X1 U8235 ( .A1(n7024), .A2(n6596), .ZN(n6767) );
  NOR2_X1 U8236 ( .A1(n11990), .A2(n11988), .ZN(n7024) );
  NAND2_X1 U8237 ( .A1(n6766), .A2(n6765), .ZN(n11993) );
  OR2_X1 U8238 ( .A1(n7023), .A2(n11989), .ZN(n6765) );
  NAND2_X1 U8239 ( .A1(n7433), .A2(n6767), .ZN(n6766) );
  INV_X1 U8240 ( .A(n11988), .ZN(n7023) );
  INV_X1 U8241 ( .A(n6843), .ZN(n6842) );
  OAI21_X1 U8242 ( .B1(n11698), .B2(n8226), .A(n11710), .ZN(n6843) );
  NAND2_X1 U8243 ( .A1(n12001), .A2(n11999), .ZN(n7440) );
  OR2_X1 U8244 ( .A1(n12001), .A2(n11999), .ZN(n7439) );
  NAND2_X1 U8245 ( .A1(n6741), .A2(n11712), .ZN(n6784) );
  AND2_X1 U8246 ( .A1(n9061), .A2(n9055), .ZN(n7593) );
  AND2_X1 U8247 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  OR2_X1 U8248 ( .A1(n11751), .A2(n11750), .ZN(n11758) );
  AND2_X1 U8249 ( .A1(n7444), .A2(n12088), .ZN(n7443) );
  INV_X1 U8250 ( .A(n12087), .ZN(n7444) );
  NAND2_X1 U8251 ( .A1(n7442), .A2(n12087), .ZN(n7441) );
  INV_X1 U8252 ( .A(n12088), .ZN(n7442) );
  NAND2_X1 U8253 ( .A1(n7620), .A2(n6617), .ZN(n7619) );
  OAI21_X1 U8254 ( .B1(n12103), .B2(n7020), .A(n7019), .ZN(n12108) );
  NAND2_X1 U8255 ( .A1(n12105), .A2(n12102), .ZN(n7019) );
  NOR2_X1 U8256 ( .A1(n12105), .A2(n12102), .ZN(n7020) );
  OAI21_X1 U8257 ( .B1(n7445), .B2(n7443), .A(n7441), .ZN(n12103) );
  NAND2_X1 U8258 ( .A1(n7029), .A2(n12115), .ZN(n7028) );
  OAI21_X1 U8259 ( .B1(n11789), .B2(n11788), .A(n12788), .ZN(n11793) );
  NAND2_X1 U8260 ( .A1(n9093), .A2(n6605), .ZN(n7634) );
  INV_X1 U8261 ( .A(n12141), .ZN(n7022) );
  NOR2_X1 U8262 ( .A1(n12144), .A2(n12141), .ZN(n7021) );
  MUX2_X1 U8263 ( .A(n14630), .B(n14452), .S(n12178), .Z(n12162) );
  NAND2_X1 U8264 ( .A1(n7616), .A2(n7614), .ZN(n7613) );
  AND2_X1 U8265 ( .A1(n9114), .A2(n9115), .ZN(n7616) );
  NOR2_X1 U8266 ( .A1(n9120), .A2(n7609), .ZN(n7611) );
  AND2_X1 U8267 ( .A1(n12708), .A2(n11810), .ZN(n6838) );
  NAND2_X1 U8268 ( .A1(n7608), .A2(n7610), .ZN(n7604) );
  INV_X1 U8269 ( .A(n7612), .ZN(n7610) );
  NAND2_X1 U8270 ( .A1(n7611), .A2(n7616), .ZN(n7603) );
  INV_X1 U8271 ( .A(n7608), .ZN(n7607) );
  INV_X1 U8272 ( .A(n7611), .ZN(n7606) );
  NAND2_X1 U8273 ( .A1(n12181), .A2(n12179), .ZN(n7446) );
  AOI21_X1 U8274 ( .B1(n8521), .B2(n8343), .A(n8537), .ZN(n7370) );
  AND2_X1 U8275 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  INV_X1 U8276 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n6996) );
  NOR2_X1 U8277 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7561) );
  NOR2_X1 U8278 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7661) );
  NOR2_X1 U8279 ( .A1(n13730), .A2(n13948), .ZN(n7035) );
  NOR2_X1 U8280 ( .A1(n13845), .A2(n7038), .ZN(n7037) );
  INV_X1 U8281 ( .A(n7039), .ZN(n7038) );
  NAND2_X1 U8282 ( .A1(n8242), .A2(n7334), .ZN(n7333) );
  INV_X1 U8283 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7334) );
  INV_X1 U8284 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8235) );
  NOR2_X1 U8285 ( .A1(n14553), .A2(n14522), .ZN(n6901) );
  INV_X1 U8286 ( .A(n14354), .ZN(n6903) );
  NOR2_X1 U8287 ( .A1(n6982), .A2(n6981), .ZN(n6980) );
  INV_X1 U8288 ( .A(n11505), .ZN(n6981) );
  INV_X1 U8289 ( .A(n11828), .ZN(n6847) );
  NOR2_X1 U8290 ( .A1(n6570), .A2(n7768), .ZN(n6746) );
  OR2_X1 U8291 ( .A1(n8108), .A2(n10300), .ZN(n7757) );
  OR2_X1 U8292 ( .A1(n10435), .A2(n10434), .ZN(n10436) );
  OR2_X1 U8293 ( .A1(n10329), .A2(n10328), .ZN(n7054) );
  NAND2_X1 U8294 ( .A1(n10436), .A2(n10441), .ZN(n10758) );
  NOR2_X1 U8295 ( .A1(n12641), .A2(n7063), .ZN(n7061) );
  INV_X1 U8296 ( .A(n12638), .ZN(n7063) );
  INV_X1 U8297 ( .A(n12658), .ZN(n7179) );
  NAND2_X1 U8298 ( .A1(n12691), .A2(n12579), .ZN(n7579) );
  BUF_X1 U8299 ( .A(n11677), .Z(n7572) );
  INV_X1 U8300 ( .A(n7579), .ZN(n7578) );
  NAND2_X1 U8301 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  INV_X1 U8302 ( .A(n7125), .ZN(n7122) );
  OR2_X1 U8303 ( .A1(n12598), .A2(n15589), .ZN(n11710) );
  AND2_X1 U8304 ( .A1(n11710), .A2(n11706), .ZN(n11662) );
  NAND2_X1 U8305 ( .A1(n6737), .A2(n6736), .ZN(n7825) );
  INV_X1 U8306 ( .A(n10293), .ZN(n11659) );
  NAND2_X1 U8307 ( .A1(n11688), .A2(n11686), .ZN(n10293) );
  OR2_X1 U8308 ( .A1(n8226), .A2(n11838), .ZN(n10310) );
  OAI21_X1 U8309 ( .B1(n8211), .B2(n8210), .A(n9899), .ZN(n8947) );
  AND4_X1 U8310 ( .A1(n7712), .A2(n8180), .A3(n8177), .A4(n7711), .ZN(n7713)
         );
  INV_X1 U8311 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7711) );
  INV_X1 U8312 ( .A(n7224), .ZN(n7221) );
  AND2_X1 U8313 ( .A1(n6997), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8314 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6996), .ZN(n6995) );
  OAI22_X1 U8315 ( .A1(n6997), .A2(n6995), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        n6996), .ZN(n6993) );
  NAND2_X1 U8316 ( .A1(n7213), .A2(n7211), .ZN(n7705) );
  NAND2_X1 U8317 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7212), .ZN(n7211) );
  AND2_X1 U8318 ( .A1(n7664), .A2(n8020), .ZN(n7665) );
  INV_X1 U8319 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U8320 ( .A1(n7956), .A2(n7561), .ZN(n7991) );
  INV_X1 U8321 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7657) );
  INV_X1 U8322 ( .A(n13384), .ZN(n13336) );
  NOR2_X1 U8323 ( .A1(n13913), .A2(n13920), .ZN(n7042) );
  INV_X1 U8324 ( .A(n7287), .ZN(n7284) );
  NOR2_X1 U8325 ( .A1(n13699), .A2(n13937), .ZN(n13670) );
  INV_X1 U8326 ( .A(n7466), .ZN(n7462) );
  NOR2_X1 U8327 ( .A1(n13792), .A2(n13981), .ZN(n7051) );
  INV_X1 U8328 ( .A(n8637), .ZN(n7469) );
  INV_X1 U8329 ( .A(n10697), .ZN(n9239) );
  INV_X1 U8330 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U8331 ( .A1(n13621), .A2(n7041), .ZN(n13591) );
  NOR2_X1 U8332 ( .A1(n13905), .A2(n13899), .ZN(n7041) );
  NAND2_X1 U8333 ( .A1(n7035), .A2(n7034), .ZN(n13699) );
  INV_X1 U8334 ( .A(n7035), .ZN(n13715) );
  NAND2_X1 U8335 ( .A1(n13885), .A2(n7037), .ZN(n13842) );
  NAND2_X1 U8336 ( .A1(n13885), .A2(n15415), .ZN(n13884) );
  INV_X1 U8337 ( .A(n11035), .ZN(n9163) );
  INV_X1 U8338 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7507) );
  AND2_X1 U8339 ( .A1(n7330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7329) );
  INV_X1 U8340 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U8341 ( .A1(n7333), .A2(n7329), .ZN(n7328) );
  NAND2_X1 U8342 ( .A1(n8412), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7327) );
  OR3_X1 U8343 ( .A1(n8538), .A2(P2_IR_REG_6__SCAN_IN), .A3(
        P2_IR_REG_7__SCAN_IN), .ZN(n8555) );
  OR2_X1 U8344 ( .A1(n8493), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8503) );
  OR2_X1 U8345 ( .A1(n12321), .A2(n7535), .ZN(n7534) );
  INV_X1 U8346 ( .A(n12325), .ZN(n7535) );
  NAND2_X1 U8347 ( .A1(n7011), .A2(n6825), .ZN(n12212) );
  INV_X1 U8348 ( .A(n12229), .ZN(n7010) );
  INV_X1 U8349 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U8350 ( .A1(n7458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7457) );
  INV_X1 U8351 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7459) );
  INV_X1 U8352 ( .A(n7152), .ZN(n7148) );
  NOR2_X1 U8353 ( .A1(n12069), .A2(n9992), .ZN(n12077) );
  INV_X1 U8354 ( .A(n7421), .ZN(n6875) );
  AOI21_X1 U8355 ( .B1(n7425), .B2(n7423), .A(n7422), .ZN(n7421) );
  INV_X1 U8356 ( .A(n14348), .ZN(n7422) );
  INV_X1 U8357 ( .A(n7427), .ZN(n7423) );
  NOR2_X1 U8358 ( .A1(n7424), .A2(n12272), .ZN(n6879) );
  INV_X1 U8359 ( .A(n7425), .ZN(n7424) );
  INV_X1 U8360 ( .A(n12017), .ZN(n6876) );
  NOR2_X1 U8361 ( .A1(n11446), .A2(n14156), .ZN(n7106) );
  NOR2_X1 U8362 ( .A1(n12002), .A2(n7094), .ZN(n7092) );
  NAND2_X1 U8363 ( .A1(n6892), .A2(n6895), .ZN(n6889) );
  NAND2_X1 U8364 ( .A1(n6860), .A2(n6866), .ZN(n9550) );
  NAND2_X1 U8365 ( .A1(n11959), .A2(n14170), .ZN(n6866) );
  NOR2_X1 U8366 ( .A1(n9549), .A2(n6862), .ZN(n6861) );
  NAND2_X1 U8367 ( .A1(n6865), .A2(n6864), .ZN(n10459) );
  INV_X1 U8368 ( .A(n9550), .ZN(n6865) );
  NAND2_X1 U8369 ( .A1(n6776), .A2(n6575), .ZN(n11942) );
  NAND2_X1 U8370 ( .A1(n14538), .A2(n14445), .ZN(n10050) );
  AND3_X1 U8371 ( .A1(n6904), .A2(n6902), .A3(n6900), .ZN(n14502) );
  AOI21_X1 U8372 ( .B1(n6903), .B2(n14520), .A(n14356), .ZN(n6902) );
  NAND2_X1 U8373 ( .A1(n6907), .A2(n6901), .ZN(n6900) );
  NAND2_X1 U8374 ( .A1(n14551), .A2(n6606), .ZN(n6904) );
  OR2_X1 U8375 ( .A1(n6906), .A2(n14553), .ZN(n6899) );
  NAND2_X1 U8376 ( .A1(n7104), .A2(n7103), .ZN(n14575) );
  AND2_X1 U8377 ( .A1(n10042), .A2(n12222), .ZN(n12238) );
  NAND2_X1 U8378 ( .A1(n9541), .A2(n7102), .ZN(n9460) );
  AND2_X1 U8379 ( .A1(n9432), .A2(n7432), .ZN(n7102) );
  NAND2_X1 U8380 ( .A1(n8395), .A2(n7390), .ZN(n8813) );
  OR2_X1 U8381 ( .A1(n8705), .A2(n10081), .ZN(n8719) );
  INV_X1 U8382 ( .A(n8670), .ZN(n8368) );
  AND2_X1 U8383 ( .A1(n8668), .A2(n8671), .ZN(n8369) );
  NAND2_X1 U8384 ( .A1(n8638), .A2(SI_14_), .ZN(n7377) );
  NAND2_X1 U8385 ( .A1(n8333), .A2(n8332), .ZN(n8496) );
  OAI21_X1 U8386 ( .B1(n8324), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6824), .ZN(
        n8322) );
  NAND2_X1 U8387 ( .A1(n8324), .A2(n9659), .ZN(n6824) );
  INV_X1 U8388 ( .A(n14759), .ZN(n6921) );
  AND2_X1 U8389 ( .A1(n14734), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6937) );
  OAI21_X1 U8390 ( .B1(n14755), .B2(n14756), .A(n6939), .ZN(n6938) );
  NAND2_X1 U8391 ( .A1(n14739), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6939) );
  AOI21_X1 U8392 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n15045), .A(n14743), .ZN(
        n14801) );
  AND2_X1 U8393 ( .A1(n11268), .A2(n6703), .ZN(n6987) );
  NOR2_X1 U8394 ( .A1(n8027), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8044) );
  OR2_X1 U8395 ( .A1(n14939), .A2(n8170), .ZN(n12445) );
  NAND2_X1 U8396 ( .A1(n7134), .A2(n7135), .ZN(n7133) );
  NAND2_X1 U8397 ( .A1(n6793), .A2(n12545), .ZN(n12529) );
  INV_X1 U8398 ( .A(n12468), .ZN(n6793) );
  INV_X1 U8399 ( .A(n6975), .ZN(n6973) );
  AOI21_X1 U8400 ( .B1(n6975), .B2(n6972), .A(n6635), .ZN(n6971) );
  INV_X1 U8401 ( .A(n9357), .ZN(n6972) );
  AND2_X1 U8402 ( .A1(n8044), .A2(n8043), .ZN(n8050) );
  NAND2_X1 U8403 ( .A1(n8050), .A2(n12537), .ZN(n8059) );
  NAND2_X1 U8404 ( .A1(n9365), .A2(n9364), .ZN(n7229) );
  AND2_X1 U8405 ( .A1(n7981), .A2(n12570), .ZN(n7995) );
  AND4_X1 U8406 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n12492)
         );
  AND4_X1 U8407 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(n12566)
         );
  AND4_X1 U8408 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n11899)
         );
  OR2_X1 U8409 ( .A1(n10238), .A2(n10744), .ZN(n10240) );
  NAND2_X1 U8410 ( .A1(n10134), .A2(n10135), .ZN(n10133) );
  NAND2_X1 U8411 ( .A1(n7175), .A2(n7173), .ZN(n15474) );
  NOR2_X1 U8412 ( .A1(n15473), .A2(n7174), .ZN(n15495) );
  NOR2_X1 U8413 ( .A1(n15495), .A2(n15494), .ZN(n15493) );
  NAND2_X1 U8414 ( .A1(n7083), .A2(n7084), .ZN(n9634) );
  NAND2_X1 U8415 ( .A1(n7080), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7079) );
  INV_X1 U8416 ( .A(n9638), .ZN(n7080) );
  AOI21_X1 U8417 ( .B1(n9613), .B2(n15509), .A(n9612), .ZN(n10203) );
  INV_X1 U8418 ( .A(n7054), .ZN(n10420) );
  NOR2_X1 U8419 ( .A1(n10766), .A2(n10767), .ZN(n10770) );
  XNOR2_X1 U8420 ( .A(n7171), .B(n14838), .ZN(n10946) );
  NOR2_X1 U8421 ( .A1(n10946), .A2(n11313), .ZN(n11051) );
  INV_X1 U8422 ( .A(n7088), .ZN(n11057) );
  NOR2_X1 U8423 ( .A1(n10940), .A2(n10939), .ZN(n11071) );
  INV_X1 U8424 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15528) );
  AND2_X1 U8425 ( .A1(n7185), .A2(n7184), .ZN(n12622) );
  INV_X1 U8426 ( .A(n7056), .ZN(n12628) );
  OR2_X1 U8427 ( .A1(n14876), .A2(n12651), .ZN(n6943) );
  AND2_X1 U8428 ( .A1(n14892), .A2(n12654), .ZN(n12655) );
  OAI211_X1 U8429 ( .C1(n14906), .C2(n7064), .A(n7062), .B(n7060), .ZN(n14927)
         );
  INV_X1 U8430 ( .A(n12641), .ZN(n7064) );
  NAND2_X1 U8431 ( .A1(n12641), .A2(n7063), .ZN(n7062) );
  NAND2_X1 U8432 ( .A1(n14906), .A2(n7061), .ZN(n7060) );
  OAI21_X1 U8433 ( .B1(n14899), .B2(n12640), .A(n14897), .ZN(n14921) );
  OR2_X1 U8434 ( .A1(n14908), .A2(n14909), .ZN(n14906) );
  INV_X1 U8435 ( .A(n12631), .ZN(n7074) );
  INV_X1 U8436 ( .A(n12664), .ZN(n7073) );
  NOR2_X1 U8437 ( .A1(n7074), .A2(n7073), .ZN(n7072) );
  INV_X1 U8438 ( .A(n12668), .ZN(n7076) );
  OAI21_X1 U8439 ( .B1(n7572), .B2(n7577), .A(n7575), .ZN(n7574) );
  NAND2_X1 U8440 ( .A1(n11677), .A2(n7579), .ZN(n7575) );
  NOR2_X1 U8441 ( .A1(n7580), .A2(n7578), .ZN(n7577) );
  NAND2_X1 U8442 ( .A1(n7557), .A2(n7560), .ZN(n7555) );
  INV_X1 U8443 ( .A(n8150), .ZN(n7560) );
  AOI21_X1 U8444 ( .B1(n7115), .B2(n7117), .A(n11787), .ZN(n7113) );
  INV_X1 U8445 ( .A(n7116), .ZN(n7115) );
  NAND2_X1 U8446 ( .A1(n12816), .A2(n8150), .ZN(n12803) );
  AOI21_X1 U8447 ( .B1(n12828), .B2(n7551), .A(n6646), .ZN(n7550) );
  INV_X1 U8448 ( .A(n8148), .ZN(n7551) );
  NAND2_X1 U8449 ( .A1(n8149), .A2(n11777), .ZN(n12816) );
  AOI21_X1 U8450 ( .B1(n7109), .B2(n7111), .A(n11769), .ZN(n7107) );
  INV_X1 U8451 ( .A(n11762), .ZN(n7111) );
  INV_X1 U8452 ( .A(n7585), .ZN(n7584) );
  AOI21_X1 U8453 ( .B1(n7585), .B2(n7583), .A(n6686), .ZN(n7582) );
  NAND2_X1 U8454 ( .A1(n7586), .A2(n7585), .ZN(n11559) );
  AND2_X1 U8455 ( .A1(n7965), .A2(n7964), .ZN(n7981) );
  NAND2_X1 U8456 ( .A1(n7586), .A2(n8144), .ZN(n11515) );
  AND2_X1 U8457 ( .A1(n11757), .A2(n11752), .ZN(n11748) );
  OAI21_X1 U8458 ( .B1(n8138), .B2(n7568), .A(n7565), .ZN(n11306) );
  AOI21_X1 U8459 ( .B1(n7567), .B2(n7566), .A(n6637), .ZN(n7565) );
  INV_X1 U8460 ( .A(n7570), .ZN(n7566) );
  AND2_X1 U8461 ( .A1(n11039), .A2(n11038), .ZN(n11718) );
  INV_X1 U8462 ( .A(n11662), .ZN(n10877) );
  NAND2_X1 U8463 ( .A1(n8131), .A2(n8130), .ZN(n11123) );
  AND2_X1 U8464 ( .A1(n11707), .A2(n7825), .ZN(n11657) );
  INV_X1 U8465 ( .A(n11702), .ZN(n11660) );
  CLKBUF_X1 U8466 ( .A(n10987), .Z(n11146) );
  NAND2_X1 U8467 ( .A1(n7129), .A2(n11688), .ZN(n15549) );
  INV_X1 U8468 ( .A(n12849), .ZN(n15561) );
  NAND2_X1 U8469 ( .A1(n7128), .A2(n11688), .ZN(n10735) );
  INV_X1 U8470 ( .A(n7129), .ZN(n7128) );
  AND2_X1 U8471 ( .A1(n8081), .A2(n8080), .ZN(n12892) );
  INV_X1 U8472 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U8473 ( .A1(n8214), .A2(n8218), .ZN(n9403) );
  AND2_X1 U8474 ( .A1(n8925), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8475 ( .A1(n8187), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6754) );
  AND2_X1 U8476 ( .A1(n8191), .A2(n8190), .ZN(n8213) );
  NOR2_X1 U8477 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  NOR2_X1 U8478 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n8188) );
  AND2_X1 U8479 ( .A1(n12987), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7228) );
  INV_X1 U8480 ( .A(n7220), .ZN(n7219) );
  AOI21_X1 U8481 ( .B1(n7220), .B2(n7218), .A(n6618), .ZN(n7217) );
  NOR2_X1 U8482 ( .A1(n8067), .A2(n7221), .ZN(n7220) );
  INV_X1 U8483 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U8484 ( .A1(n7701), .A2(n7700), .ZN(n8002) );
  INV_X1 U8485 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8003) );
  INV_X1 U8486 ( .A(n7991), .ZN(n8004) );
  NAND2_X1 U8487 ( .A1(n7198), .A2(n7698), .ZN(n7977) );
  CLKBUF_X1 U8488 ( .A(n7955), .Z(n7956) );
  INV_X1 U8489 ( .A(n7210), .ZN(n7209) );
  OR2_X1 U8490 ( .A1(n7916), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7918) );
  XNOR2_X1 U8491 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7885) );
  NAND2_X1 U8492 ( .A1(n7658), .A2(n7659), .ZN(n7852) );
  XNOR2_X1 U8493 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7868) );
  NOR2_X1 U8494 ( .A1(n6626), .A2(n7215), .ZN(n7214) );
  XNOR2_X1 U8495 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7854) );
  NOR2_X1 U8496 ( .A1(n7799), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7817) );
  OAI21_X1 U8497 ( .B1(n7204), .B2(n7203), .A(n7201), .ZN(n7798) );
  AOI21_X1 U8498 ( .B1(n7202), .B2(n7785), .A(n6685), .ZN(n7201) );
  INV_X1 U8499 ( .A(n7677), .ZN(n7202) );
  XNOR2_X1 U8500 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7796) );
  NAND2_X1 U8501 ( .A1(n7187), .A2(n7186), .ZN(n7783) );
  INV_X1 U8502 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7186) );
  NAND2_X1 U8503 ( .A1(n7077), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7771) );
  AND2_X1 U8504 ( .A1(n8423), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7765) );
  NOR2_X1 U8505 ( .A1(n7316), .A2(n7321), .ZN(n7311) );
  INV_X1 U8506 ( .A(n13343), .ZN(n7316) );
  AND2_X1 U8507 ( .A1(n13343), .A2(n6623), .ZN(n7315) );
  INV_X1 U8508 ( .A(n13337), .ZN(n7313) );
  INV_X1 U8509 ( .A(n13344), .ZN(n7322) );
  OR2_X1 U8510 ( .A1(n8645), .A2(n8644), .ZN(n8657) );
  NAND2_X1 U8511 ( .A1(n11299), .A2(n11490), .ZN(n7350) );
  INV_X1 U8512 ( .A(n13853), .ZN(n11873) );
  OR2_X1 U8513 ( .A1(n8630), .A2(n8629), .ZN(n8645) );
  NAND2_X1 U8514 ( .A1(n13392), .A2(n13322), .ZN(n13326) );
  INV_X1 U8515 ( .A(n7359), .ZN(n7358) );
  AND2_X1 U8516 ( .A1(n11228), .A2(n7356), .ZN(n7355) );
  NOR2_X1 U8517 ( .A1(n11263), .A2(n7360), .ZN(n7359) );
  INV_X1 U8518 ( .A(n11222), .ZN(n7360) );
  NAND2_X1 U8519 ( .A1(n11865), .A2(n7335), .ZN(n10637) );
  NOR2_X1 U8520 ( .A1(n10640), .A2(n7336), .ZN(n7335) );
  INV_X1 U8521 ( .A(n10563), .ZN(n7336) );
  AOI21_X1 U8522 ( .B1(n7348), .B2(n7346), .A(n7345), .ZN(n7344) );
  INV_X1 U8523 ( .A(n7348), .ZN(n7347) );
  INV_X1 U8524 ( .A(n11490), .ZN(n7346) );
  AND2_X1 U8525 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  XNOR2_X1 U8526 ( .A(n8276), .B(n8275), .ZN(n9840) );
  OAI21_X1 U8527 ( .B1(n8274), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8276) );
  AOI21_X1 U8528 ( .B1(n9942), .B2(n9931), .A(n9930), .ZN(n9933) );
  NOR2_X1 U8529 ( .A1(n10013), .A2(n10014), .ZN(n11004) );
  AOI21_X1 U8530 ( .B1(n13522), .B2(n13824), .A(n13519), .ZN(n15262) );
  OAI21_X1 U8531 ( .B1(n11002), .B2(n15273), .A(n15275), .ZN(n11007) );
  XOR2_X1 U8532 ( .A(n15299), .B(n11009), .Z(n15303) );
  INV_X1 U8533 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U8534 ( .A1(n7352), .A2(n8239), .ZN(n7351) );
  INV_X1 U8535 ( .A(n7353), .ZN(n7352) );
  INV_X1 U8536 ( .A(n6813), .ZN(n13550) );
  NAND2_X1 U8537 ( .A1(n9190), .A2(n9189), .ZN(n13575) );
  NOR2_X1 U8538 ( .A1(n12429), .A2(n13591), .ZN(n13579) );
  OR2_X1 U8539 ( .A1(n8846), .A2(n8306), .ZN(n12430) );
  NAND2_X1 U8540 ( .A1(n8838), .A2(n7476), .ZN(n7472) );
  NAND2_X1 U8541 ( .A1(n7471), .A2(n7476), .ZN(n7470) );
  NAND2_X1 U8542 ( .A1(n13905), .A2(n8852), .ZN(n7476) );
  INV_X1 U8543 ( .A(n13608), .ZN(n8915) );
  AND2_X1 U8544 ( .A1(n8830), .A2(n8844), .ZN(n13622) );
  NAND2_X1 U8545 ( .A1(n13652), .A2(n13641), .ZN(n13636) );
  OR2_X1 U8546 ( .A1(n8788), .A2(n13365), .ZN(n8804) );
  INV_X1 U8547 ( .A(n7481), .ZN(n7480) );
  AOI21_X1 U8548 ( .B1(n7481), .B2(n7479), .A(n7478), .ZN(n7477) );
  INV_X1 U8549 ( .A(n8764), .ZN(n7479) );
  NAND2_X1 U8550 ( .A1(n8301), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8728) );
  AOI21_X1 U8551 ( .B1(n7279), .B2(n7277), .A(n6670), .ZN(n7276) );
  INV_X1 U8552 ( .A(n7279), .ZN(n7278) );
  INV_X1 U8553 ( .A(n8900), .ZN(n7277) );
  NAND2_X1 U8554 ( .A1(n13788), .A2(n6608), .ZN(n13754) );
  AOI21_X1 U8555 ( .B1(n7293), .B2(n7291), .A(n6669), .ZN(n7290) );
  INV_X1 U8556 ( .A(n7293), .ZN(n7292) );
  NAND2_X1 U8557 ( .A1(n13788), .A2(n7049), .ZN(n13774) );
  NAND2_X1 U8558 ( .A1(n13788), .A2(n14967), .ZN(n13980) );
  AND2_X1 U8559 ( .A1(n11376), .A2(n11380), .ZN(n13788) );
  NAND2_X1 U8560 ( .A1(n7267), .A2(n7266), .ZN(n13811) );
  AOI21_X1 U8561 ( .B1(n7268), .B2(n7270), .A(n6651), .ZN(n7266) );
  NAND2_X1 U8562 ( .A1(n8584), .A2(n8583), .ZN(n13816) );
  INV_X1 U8563 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8560) );
  OR2_X1 U8564 ( .A1(n8561), .A2(n8560), .ZN(n8576) );
  INV_X1 U8565 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8542) );
  OR2_X1 U8566 ( .A1(n8543), .A2(n8542), .ZN(n8561) );
  AND2_X1 U8567 ( .A1(n7260), .A2(n6709), .ZN(n7259) );
  INV_X1 U8568 ( .A(n13870), .ZN(n13868) );
  INV_X1 U8569 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8528) );
  OR2_X1 U8570 ( .A1(n8529), .A2(n8528), .ZN(n8543) );
  AND2_X1 U8571 ( .A1(n10689), .A2(n10671), .ZN(n13885) );
  NOR2_X1 U8572 ( .A1(n10686), .A2(n15396), .ZN(n10689) );
  OR2_X1 U8573 ( .A1(n10702), .A2(n15390), .ZN(n10686) );
  NAND2_X1 U8574 ( .A1(n10701), .A2(n10706), .ZN(n10702) );
  CLKBUF_X1 U8575 ( .A(n13879), .Z(n6801) );
  INV_X1 U8576 ( .A(n7257), .ZN(n15320) );
  NAND2_X1 U8577 ( .A1(n8437), .A2(n7485), .ZN(n7484) );
  OAI21_X1 U8578 ( .B1(n9709), .B2(n9681), .A(n7486), .ZN(n7485) );
  NAND2_X1 U8579 ( .A1(n9681), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7486) );
  INV_X1 U8580 ( .A(n15428), .ZN(n15434) );
  AND2_X1 U8581 ( .A1(n15438), .A2(n6801), .ZN(n15407) );
  OR2_X1 U8582 ( .A1(n15438), .A2(n9163), .ZN(n10183) );
  INV_X1 U8583 ( .A(n8258), .ZN(n7046) );
  NAND2_X1 U8584 ( .A1(n8274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8254) );
  NOR2_X1 U8585 ( .A1(n8605), .A2(n7353), .ZN(n8640) );
  AND2_X1 U8586 ( .A1(n8523), .A2(n8508), .ZN(n9852) );
  AND2_X1 U8587 ( .A1(n7308), .A2(n7309), .ZN(n8439) );
  INV_X1 U8588 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7309) );
  INV_X1 U8589 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8423) );
  AND2_X1 U8590 ( .A1(n14985), .A2(n14986), .ZN(n12321) );
  OR2_X1 U8591 ( .A1(n10465), .A2(n10464), .ZN(n10501) );
  XNOR2_X1 U8592 ( .A(n6778), .B(n6777), .ZN(n10038) );
  INV_X1 U8593 ( .A(n12413), .ZN(n6777) );
  OAI22_X1 U8594 ( .A1(n6575), .A2(n12371), .B1(n11938), .B2(n12370), .ZN(
        n6778) );
  NOR2_X1 U8595 ( .A1(n9681), .A2(n9710), .ZN(n7166) );
  INV_X1 U8596 ( .A(n10585), .ZN(n7545) );
  AOI22_X1 U8597 ( .A1(n10033), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n10035), .B2(
        n10371), .ZN(n6816) );
  NAND2_X1 U8598 ( .A1(n14117), .A2(n14118), .ZN(n14116) );
  NOR2_X1 U8599 ( .A1(n11186), .A2(n9991), .ZN(n11345) );
  AND2_X1 U8600 ( .A1(n11345), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11437) );
  INV_X1 U8601 ( .A(n11348), .ZN(n12147) );
  NAND2_X1 U8602 ( .A1(n12092), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U8603 ( .A1(n9451), .A2(n14714), .ZN(n9494) );
  INV_X1 U8604 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14724) );
  NAND2_X1 U8605 ( .A1(n12236), .A2(n12235), .ZN(n14336) );
  AND2_X1 U8606 ( .A1(n14436), .A2(n6698), .ZN(n14339) );
  INV_X1 U8607 ( .A(n7100), .ZN(n7098) );
  AND2_X1 U8608 ( .A1(n6632), .A2(n6872), .ZN(n7162) );
  INV_X1 U8609 ( .A(n7163), .ZN(n7160) );
  NAND2_X1 U8610 ( .A1(n6631), .A2(n6827), .ZN(n14401) );
  NOR2_X1 U8611 ( .A1(n14413), .A2(n7164), .ZN(n7163) );
  INV_X1 U8612 ( .A(n14386), .ZN(n7164) );
  NAND2_X1 U8613 ( .A1(n14417), .A2(n14420), .ZN(n14416) );
  XNOR2_X1 U8614 ( .A(n14630), .B(n14452), .ZN(n14441) );
  OAI21_X1 U8615 ( .B1(n6884), .B2(n14485), .A(n6880), .ZN(n14442) );
  AOI21_X1 U8616 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(n6880) );
  INV_X1 U8617 ( .A(n14360), .ZN(n6881) );
  INV_X1 U8618 ( .A(n7414), .ZN(n6882) );
  INV_X1 U8619 ( .A(n7457), .ZN(n7452) );
  NAND2_X1 U8620 ( .A1(n7452), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7451) );
  INV_X1 U8621 ( .A(n7456), .ZN(n7455) );
  OAI22_X1 U8622 ( .A1(n7457), .A2(n7459), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        n7458), .ZN(n7456) );
  NAND2_X1 U8623 ( .A1(n14380), .A2(n14491), .ZN(n7144) );
  OR2_X1 U8624 ( .A1(n7145), .A2(n7143), .ZN(n7142) );
  INV_X1 U8625 ( .A(n14380), .ZN(n7143) );
  AND2_X1 U8626 ( .A1(n14474), .A2(n6624), .ZN(n7145) );
  XNOR2_X1 U8627 ( .A(n14677), .B(n14370), .ZN(n14566) );
  NAND2_X1 U8628 ( .A1(n6877), .A2(n6874), .ZN(n14567) );
  OR2_X1 U8629 ( .A1(n11436), .A2(n6878), .ZN(n6877) );
  AOI21_X1 U8630 ( .B1(n6879), .B2(n6876), .A(n6875), .ZN(n6874) );
  INV_X1 U8631 ( .A(n6879), .ZN(n6878) );
  NAND2_X1 U8632 ( .A1(n7106), .A2(n7105), .ZN(n14584) );
  INV_X1 U8633 ( .A(n7106), .ZN(n11535) );
  INV_X1 U8634 ( .A(n7155), .ZN(n7154) );
  OAI21_X1 U8635 ( .B1(n7156), .B2(n7157), .A(n11531), .ZN(n7155) );
  OR2_X1 U8636 ( .A1(n10960), .A2(n10959), .ZN(n11186) );
  INV_X1 U8637 ( .A(n7417), .ZN(n7416) );
  NAND2_X1 U8638 ( .A1(n10912), .A2(n7096), .ZN(n10969) );
  OR2_X1 U8639 ( .A1(n10501), .A2(n10500), .ZN(n10514) );
  NOR2_X1 U8640 ( .A1(n10514), .A2(n10513), .ZN(n10822) );
  NAND2_X1 U8641 ( .A1(n6891), .A2(n6892), .ZN(n10906) );
  NAND2_X1 U8642 ( .A1(n10614), .A2(n6894), .ZN(n6891) );
  NAND2_X1 U8643 ( .A1(n7091), .A2(n7090), .ZN(n10623) );
  NAND2_X1 U8644 ( .A1(n10459), .A2(n10458), .ZN(n10486) );
  AND2_X1 U8645 ( .A1(n6652), .A2(n9506), .ZN(n7140) );
  INV_X1 U8646 ( .A(n15091), .ZN(n14538) );
  INV_X1 U8647 ( .A(n15077), .ZN(n15080) );
  NAND2_X1 U8648 ( .A1(n9586), .A2(n10123), .ZN(n14393) );
  OR2_X1 U8649 ( .A1(n14174), .A2(n15135), .ZN(n11934) );
  INV_X1 U8650 ( .A(n14364), .ZN(n6868) );
  INV_X1 U8651 ( .A(n14363), .ZN(n6873) );
  AND2_X1 U8652 ( .A1(n6871), .A2(n14413), .ZN(n6870) );
  NAND2_X1 U8653 ( .A1(n6872), .A2(n14363), .ZN(n6871) );
  NAND2_X1 U8654 ( .A1(n10044), .A2(n10043), .ZN(n15169) );
  INV_X1 U8655 ( .A(n15169), .ZN(n15194) );
  AND2_X1 U8656 ( .A1(n10041), .A2(n10054), .ZN(n10123) );
  INV_X1 U8657 ( .A(n15198), .ZN(n15131) );
  XNOR2_X1 U8658 ( .A(n9155), .B(n9154), .ZN(n12224) );
  AND2_X1 U8659 ( .A1(n7432), .A2(n9458), .ZN(n7431) );
  INV_X1 U8660 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9449) );
  XNOR2_X1 U8661 ( .A(n9459), .B(n9458), .ZN(n9554) );
  NAND2_X1 U8662 ( .A1(n9460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9459) );
  AND2_X1 U8663 ( .A1(n8825), .A2(n8824), .ZN(n12295) );
  OR2_X1 U8664 ( .A1(n8823), .A2(n8400), .ZN(n8825) );
  NAND2_X1 U8665 ( .A1(n9444), .A2(n9443), .ZN(n10053) );
  NAND2_X1 U8666 ( .A1(n8381), .A2(SI_20_), .ZN(n6953) );
  NOR2_X1 U8667 ( .A1(n6955), .A2(n6952), .ZN(n6951) );
  XNOR2_X1 U8668 ( .A(n8721), .B(n8718), .ZN(n12052) );
  INV_X1 U8669 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U8670 ( .A1(n7369), .A2(n8343), .ZN(n8536) );
  NAND2_X1 U8671 ( .A1(n8522), .A2(n8341), .ZN(n7369) );
  INV_X1 U8672 ( .A(n8521), .ZN(n8341) );
  OR2_X1 U8673 ( .A1(n9518), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9691) );
  AND2_X2 U8674 ( .A1(n9462), .A2(n9487), .ZN(n9502) );
  INV_X1 U8675 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U8676 ( .A1(n15643), .A2(n15644), .ZN(n14765) );
  INV_X1 U8677 ( .A(n7393), .ZN(n14760) );
  NAND2_X1 U8678 ( .A1(n14840), .A2(n14839), .ZN(n7410) );
  NAND2_X1 U8679 ( .A1(n7404), .A2(n7406), .ZN(n14797) );
  NAND2_X1 U8680 ( .A1(n6934), .A2(n15296), .ZN(n6933) );
  INV_X1 U8681 ( .A(n15022), .ZN(n6934) );
  NAND2_X1 U8682 ( .A1(n15027), .A2(n6925), .ZN(n6924) );
  NAND2_X1 U8683 ( .A1(n14859), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8684 ( .A1(n14752), .A2(n14751), .ZN(n14868) );
  NAND2_X1 U8685 ( .A1(n10792), .A2(n10791), .ZN(n10790) );
  AND2_X1 U8686 ( .A1(n6988), .A2(n6703), .ZN(n11269) );
  NAND2_X1 U8687 ( .A1(n6988), .A2(n6987), .ZN(n11267) );
  NAND2_X1 U8688 ( .A1(n9389), .A2(n9388), .ZN(n12455) );
  NAND2_X1 U8689 ( .A1(n10790), .A2(n9335), .ZN(n10924) );
  OAI21_X1 U8690 ( .B1(n10792), .B2(n7244), .A(n7241), .ZN(n10922) );
  NAND2_X1 U8691 ( .A1(n7232), .A2(n9361), .ZN(n12483) );
  NAND2_X1 U8692 ( .A1(n8058), .A2(n8057), .ZN(n12781) );
  NAND2_X1 U8693 ( .A1(n7747), .A2(n7746), .ZN(n12727) );
  INV_X1 U8694 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n14900) );
  NAND2_X1 U8695 ( .A1(n12508), .A2(n12507), .ZN(n12506) );
  NAND2_X1 U8696 ( .A1(n12563), .A2(n9351), .ZN(n12508) );
  NAND2_X1 U8697 ( .A1(n7252), .A2(n7253), .ZN(n12516) );
  OR2_X1 U8698 ( .A1(n12563), .A2(n7255), .ZN(n7252) );
  AND2_X1 U8699 ( .A1(n6966), .A2(n6639), .ZN(n10411) );
  AOI21_X1 U8700 ( .B1(n7241), .B2(n7244), .A(n6684), .ZN(n7240) );
  INV_X1 U8701 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U8702 ( .A1(n6984), .A2(n11504), .ZN(n11902) );
  OAI21_X1 U8703 ( .B1(n15554), .B2(n9328), .A(n11688), .ZN(n9324) );
  INV_X1 U8704 ( .A(n12576), .ZN(n15463) );
  AOI21_X1 U8705 ( .B1(n7250), .B2(n7255), .A(n6724), .ZN(n7248) );
  NOR2_X1 U8706 ( .A1(n12514), .A2(n7251), .ZN(n7250) );
  AND2_X1 U8707 ( .A1(n9332), .A2(n6737), .ZN(n7245) );
  NAND2_X1 U8708 ( .A1(n12554), .A2(n6989), .ZN(n12556) );
  NAND2_X1 U8709 ( .A1(n12496), .A2(n6609), .ZN(n6989) );
  NAND2_X1 U8710 ( .A1(n9406), .A2(n9405), .ZN(n12571) );
  AND2_X1 U8711 ( .A1(n9393), .A2(n11839), .ZN(n15469) );
  NAND2_X1 U8712 ( .A1(n10152), .A2(n11843), .ZN(n12573) );
  OR2_X1 U8713 ( .A1(n7652), .A2(n11836), .ZN(n6836) );
  OAI21_X1 U8714 ( .B1(n11652), .B2(n7640), .A(n11651), .ZN(n11653) );
  INV_X1 U8715 ( .A(n11650), .ZN(n11651) );
  INV_X1 U8716 ( .A(n12523), .ZN(n12582) );
  INV_X1 U8717 ( .A(n11563), .ZN(n12848) );
  INV_X1 U8718 ( .A(n12566), .ZN(n12590) );
  OR2_X1 U8719 ( .A1(n8108), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n6794) );
  CLKBUF_X1 U8720 ( .A(n12601), .Z(n6822) );
  NOR2_X1 U8721 ( .A1(n10356), .A2(n9616), .ZN(n10355) );
  INV_X1 U8722 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15489) );
  INV_X1 U8723 ( .A(n7192), .ZN(n15513) );
  INV_X1 U8724 ( .A(n15538), .ZN(n14920) );
  INV_X1 U8725 ( .A(n9621), .ZN(n7191) );
  AOI21_X1 U8726 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(n10433) );
  NOR2_X1 U8727 ( .A1(n10321), .A2(n10322), .ZN(n10324) );
  NOR2_X1 U8728 ( .A1(n10422), .A2(n15629), .ZN(n10766) );
  INV_X1 U8729 ( .A(n6941), .ZN(n10944) );
  XNOR2_X1 U8730 ( .A(n7088), .B(n14838), .ZN(n10934) );
  NOR2_X1 U8731 ( .A1(n10934), .A2(n11323), .ZN(n11059) );
  NAND2_X1 U8732 ( .A1(n12618), .A2(n6723), .ZN(n7180) );
  NOR2_X1 U8733 ( .A1(n15532), .A2(n12605), .ZN(n12606) );
  INV_X1 U8734 ( .A(n7053), .ZN(n12604) );
  XNOR2_X1 U8735 ( .A(n12650), .B(n12649), .ZN(n14877) );
  INV_X1 U8736 ( .A(n6943), .ZN(n14895) );
  XNOR2_X1 U8737 ( .A(n12655), .B(n14925), .ZN(n14915) );
  NOR2_X1 U8738 ( .A1(n14915), .A2(n14916), .ZN(n14914) );
  OAI21_X1 U8739 ( .B1(n6682), .B2(n15560), .A(n9408), .ZN(n6852) );
  AND2_X1 U8740 ( .A1(n12739), .A2(n12738), .ZN(n12886) );
  NAND2_X1 U8741 ( .A1(n7119), .A2(n7124), .ZN(n12740) );
  NAND2_X1 U8742 ( .A1(n6787), .A2(n7125), .ZN(n7119) );
  NAND2_X1 U8743 ( .A1(n8156), .A2(n8155), .ZN(n12750) );
  NAND2_X1 U8744 ( .A1(n11790), .A2(n12793), .ZN(n12780) );
  NAND2_X1 U8745 ( .A1(n7114), .A2(n11776), .ZN(n12802) );
  NAND2_X1 U8746 ( .A1(n12820), .A2(n11775), .ZN(n7114) );
  NAND2_X1 U8747 ( .A1(n12829), .A2(n12828), .ZN(n12827) );
  NAND2_X1 U8748 ( .A1(n12865), .A2(n11762), .ZN(n12843) );
  NAND2_X1 U8749 ( .A1(n7569), .A2(n7567), .ZN(n11202) );
  NAND2_X1 U8750 ( .A1(n8138), .A2(n11038), .ZN(n11091) );
  AND2_X1 U8751 ( .A1(n7564), .A2(n8134), .ZN(n10977) );
  INV_X1 U8752 ( .A(n10413), .ZN(n15581) );
  OR2_X1 U8753 ( .A1(n10316), .A2(n10315), .ZN(n12870) );
  AND2_X1 U8754 ( .A1(n10307), .A2(n15552), .ZN(n14938) );
  INV_X1 U8755 ( .A(n12715), .ZN(n13219) );
  INV_X1 U8756 ( .A(n12744), .ZN(n13227) );
  NAND2_X1 U8757 ( .A1(n8040), .A2(n8039), .ZN(n13244) );
  OR3_X1 U8758 ( .A1(n12913), .A2(n12912), .A3(n12911), .ZN(n13245) );
  NAND2_X1 U8759 ( .A1(n7962), .A2(n7961), .ZN(n13260) );
  NAND2_X1 U8760 ( .A1(n9403), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13266) );
  XNOR2_X1 U8761 ( .A(n11632), .B(n11631), .ZN(n13269) );
  NAND2_X1 U8762 ( .A1(n11628), .A2(n11627), .ZN(n11632) );
  INV_X1 U8763 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13268) );
  INV_X1 U8764 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7730) );
  INV_X1 U8765 ( .A(n11625), .ZN(n6797) );
  INV_X1 U8766 ( .A(n8213), .ZN(n13285) );
  NAND2_X1 U8767 ( .A1(n8184), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U8768 ( .A1(n7222), .A2(n7224), .ZN(n8068) );
  NAND2_X1 U8769 ( .A1(n8056), .A2(n8055), .ZN(n7222) );
  NAND2_X1 U8770 ( .A1(n7673), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7674) );
  INV_X1 U8771 ( .A(n11682), .ZN(n10789) );
  XNOR2_X1 U8772 ( .A(n7667), .B(n6998), .ZN(n10555) );
  INV_X1 U8773 ( .A(SI_19_), .ZN(n10158) );
  INV_X1 U8774 ( .A(SI_15_), .ZN(n9873) );
  INV_X1 U8775 ( .A(SI_13_), .ZN(n9745) );
  INV_X1 U8776 ( .A(SI_12_), .ZN(n9689) );
  INV_X1 U8777 ( .A(n7208), .ZN(n7915) );
  AOI21_X1 U8778 ( .B1(n7904), .B2(n7903), .A(n6714), .ZN(n7208) );
  INV_X1 U8779 ( .A(SI_10_), .ZN(n9668) );
  XNOR2_X1 U8780 ( .A(n7902), .B(n7901), .ZN(n10945) );
  INV_X1 U8781 ( .A(n10424), .ZN(n10441) );
  INV_X1 U8782 ( .A(n10197), .ZN(n10212) );
  NAND2_X1 U8783 ( .A1(n7216), .A2(n7680), .ZN(n7834) );
  NAND2_X1 U8784 ( .A1(n7799), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U8785 ( .A1(n7204), .A2(n7677), .ZN(n7786) );
  NAND2_X1 U8786 ( .A1(n11919), .A2(P3_U3151), .ZN(n13284) );
  NAND2_X1 U8787 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7759) );
  NAND2_X1 U8788 ( .A1(n7350), .A2(n11495), .ZN(n11496) );
  NAND2_X1 U8789 ( .A1(n11883), .A2(n11222), .ZN(n11262) );
  OR2_X1 U8790 ( .A1(n8740), .A2(n9660), .ZN(n8471) );
  NOR2_X1 U8791 ( .A1(n13382), .A2(n13381), .ZN(n13387) );
  AND2_X1 U8792 ( .A1(n11892), .A2(n11213), .ZN(n6848) );
  NAND2_X1 U8793 ( .A1(n13455), .A2(n7361), .ZN(n13392) );
  AND2_X1 U8794 ( .A1(n13393), .A2(n13317), .ZN(n7361) );
  AND2_X1 U8795 ( .A1(n13455), .A2(n13317), .ZN(n13394) );
  NAND2_X1 U8796 ( .A1(n7319), .A2(n6623), .ZN(n7318) );
  NAND2_X1 U8797 ( .A1(n7337), .A2(n7341), .ZN(n13427) );
  NAND2_X1 U8798 ( .A1(n13416), .A2(n13300), .ZN(n13428) );
  NAND2_X1 U8799 ( .A1(n6782), .A2(n13300), .ZN(n7337) );
  NAND2_X1 U8800 ( .A1(n13360), .A2(n13359), .ZN(n13400) );
  AND2_X1 U8801 ( .A1(n10405), .A2(n10398), .ZN(n6849) );
  NAND2_X1 U8802 ( .A1(n11218), .A2(n11877), .ZN(n11883) );
  MUX2_X1 U8803 ( .A(n7308), .B(n14025), .S(n8437), .Z(n10721) );
  NAND2_X1 U8804 ( .A1(n13312), .A2(n13370), .ZN(n13450) );
  AOI21_X1 U8805 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(n7338) );
  INV_X1 U8806 ( .A(n13306), .ZN(n7339) );
  INV_X1 U8807 ( .A(n13300), .ZN(n7340) );
  NAND2_X1 U8808 ( .A1(n11865), .A2(n10563), .ZN(n10639) );
  NAND2_X1 U8809 ( .A1(n8810), .A2(n8809), .ZN(n13632) );
  NAND2_X1 U8810 ( .A1(n8779), .A2(n8778), .ZN(n13461) );
  NAND2_X1 U8811 ( .A1(n8763), .A2(n8762), .ZN(n13501) );
  NAND2_X1 U8812 ( .A1(n11014), .A2(n6759), .ZN(n11106) );
  AND2_X1 U8813 ( .A1(n11012), .A2(n11107), .ZN(n6759) );
  NAND2_X1 U8814 ( .A1(n11106), .A2(n11107), .ZN(n11108) );
  OAI21_X1 U8815 ( .B1(n13536), .B2(n13539), .A(n6813), .ZN(n13537) );
  INV_X1 U8816 ( .A(n13571), .ZN(n13897) );
  NAND2_X1 U8817 ( .A1(n7473), .A2(n8838), .ZN(n13599) );
  NAND2_X1 U8818 ( .A1(n7275), .A2(n7273), .ZN(n13609) );
  NAND2_X1 U8819 ( .A1(n7282), .A2(n7286), .ZN(n13628) );
  NAND2_X1 U8820 ( .A1(n13669), .A2(n7287), .ZN(n7282) );
  NAND2_X1 U8821 ( .A1(n7289), .A2(n7288), .ZN(n13656) );
  NAND2_X1 U8822 ( .A1(n7289), .A2(n7287), .ZN(n13927) );
  NAND2_X1 U8823 ( .A1(n7483), .A2(n7481), .ZN(n13683) );
  NAND2_X1 U8824 ( .A1(n8726), .A2(n8725), .ZN(n13951) );
  NAND2_X1 U8825 ( .A1(n7495), .A2(n7496), .ZN(n13738) );
  NAND2_X1 U8826 ( .A1(n7499), .A2(n7501), .ZN(n13751) );
  NAND2_X1 U8827 ( .A1(n7294), .A2(n7295), .ZN(n13972) );
  NAND2_X1 U8828 ( .A1(n11382), .A2(n7298), .ZN(n7294) );
  NAND2_X1 U8829 ( .A1(n7463), .A2(n7466), .ZN(n13974) );
  NAND2_X1 U8830 ( .A1(n7465), .A2(n8637), .ZN(n13783) );
  NAND2_X1 U8831 ( .A1(n11374), .A2(n8636), .ZN(n7465) );
  OAI21_X1 U8832 ( .B1(n11382), .B2(n6674), .A(n7300), .ZN(n13787) );
  NAND2_X1 U8833 ( .A1(n8608), .A2(n8607), .ZN(n13808) );
  NAND2_X1 U8834 ( .A1(n8594), .A2(n8593), .ZN(n15435) );
  NAND2_X1 U8835 ( .A1(n13850), .A2(n8891), .ZN(n13832) );
  NAND2_X1 U8836 ( .A1(n8558), .A2(n8557), .ZN(n13865) );
  NAND2_X1 U8837 ( .A1(n7263), .A2(n8887), .ZN(n10662) );
  NAND2_X1 U8838 ( .A1(n10676), .A2(n10675), .ZN(n7263) );
  OR2_X1 U8839 ( .A1(n10183), .A2(n15364), .ZN(n13880) );
  NAND2_X1 U8840 ( .A1(n6771), .A2(n9849), .ZN(n6770) );
  XNOR2_X1 U8841 ( .A(n15311), .B(n7257), .ZN(n15314) );
  INV_X1 U8842 ( .A(n14957), .ZN(n15317) );
  INV_X1 U8843 ( .A(n8968), .ZN(n10864) );
  NOR2_X2 U8844 ( .A1(n15316), .A2(n6587), .ZN(n15326) );
  OR2_X1 U8845 ( .A1(n13935), .A2(n13934), .ZN(n13992) );
  AND2_X1 U8846 ( .A1(n10176), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15367) );
  INV_X1 U8847 ( .A(n15367), .ZN(n15364) );
  INV_X1 U8848 ( .A(n8313), .ZN(n11869) );
  INV_X1 U8849 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14012) );
  INV_X1 U8850 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U8851 ( .A1(n8408), .A2(n8264), .ZN(n14019) );
  INV_X1 U8852 ( .A(n6589), .ZN(n8270) );
  INV_X1 U8853 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11320) );
  CLKBUF_X1 U8854 ( .A(n11319), .Z(n6783) );
  INV_X1 U8855 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10027) );
  INV_X1 U8856 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9753) );
  INV_X1 U8857 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9687) );
  INV_X1 U8858 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9686) );
  INV_X1 U8859 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9662) );
  INV_X1 U8860 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8479) );
  INV_X1 U8861 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U8862 ( .A1(n7525), .A2(n7526), .ZN(n14027) );
  AOI21_X1 U8863 ( .B1(n7528), .B2(n7530), .A(n6665), .ZN(n7526) );
  NAND2_X1 U8864 ( .A1(n14987), .A2(n12321), .ZN(n14990) );
  AND2_X1 U8865 ( .A1(n7513), .A2(n7512), .ZN(n11397) );
  INV_X1 U8866 ( .A(n7518), .ZN(n7512) );
  NAND2_X1 U8867 ( .A1(n7516), .A2(n7513), .ZN(n11578) );
  AND2_X1 U8868 ( .A1(n10533), .A2(n10532), .ZN(n10534) );
  NAND2_X1 U8869 ( .A1(n7544), .A2(n12347), .ZN(n14051) );
  AND2_X1 U8870 ( .A1(n10123), .A2(n10058), .ZN(n14152) );
  NAND2_X1 U8871 ( .A1(n11135), .A2(n11134), .ZN(n11138) );
  NAND2_X1 U8872 ( .A1(n14097), .A2(n12362), .ZN(n14060) );
  NAND2_X1 U8873 ( .A1(n12101), .A2(n12100), .ZN(n14657) );
  OR2_X1 U8874 ( .A1(n12099), .A2(n12123), .ZN(n12101) );
  NAND2_X1 U8875 ( .A1(n11600), .A2(n11599), .ZN(n11606) );
  AOI21_X1 U8876 ( .B1(n7521), .B2(n7524), .A(n6666), .ZN(n7520) );
  INV_X1 U8877 ( .A(n12377), .ZN(n7524) );
  INV_X1 U8878 ( .A(n14540), .ZN(n14663) );
  OR2_X1 U8879 ( .A1(n12308), .A2(n12307), .ZN(n7639) );
  NAND2_X1 U8880 ( .A1(n6583), .A2(n14107), .ZN(n14987) );
  INV_X1 U8881 ( .A(n7511), .ZN(n7510) );
  AOI21_X1 U8882 ( .B1(n11396), .B2(n11386), .A(n7509), .ZN(n7508) );
  NAND2_X1 U8883 ( .A1(n12340), .A2(n6806), .ZN(n14130) );
  NAND2_X1 U8884 ( .A1(n12338), .A2(n12339), .ZN(n6806) );
  INV_X1 U8885 ( .A(n14989), .ZN(n14119) );
  AND2_X1 U8886 ( .A1(n11342), .A2(n15169), .ZN(n14995) );
  AND2_X1 U8887 ( .A1(n6648), .A2(n7655), .ZN(n7009) );
  INV_X1 U8888 ( .A(n14376), .ZN(n14525) );
  OAI21_X1 U8889 ( .B1(n14100), .B2(n12202), .A(n12083), .ZN(n14526) );
  OAI211_X1 U8890 ( .C1(n14585), .C2(n12202), .A(n11545), .B(n11544), .ZN(
        n14568) );
  INV_X1 U8891 ( .A(n14385), .ZN(n14421) );
  NAND2_X1 U8892 ( .A1(n14471), .A2(n6883), .ZN(n14450) );
  NAND2_X1 U8893 ( .A1(n14485), .A2(n14358), .ZN(n14473) );
  NAND2_X1 U8894 ( .A1(n7151), .A2(n14373), .ZN(n14535) );
  NAND2_X1 U8895 ( .A1(n6909), .A2(n14352), .ZN(n14545) );
  NAND2_X1 U8896 ( .A1(n6910), .A2(n14553), .ZN(n6909) );
  NAND2_X1 U8897 ( .A1(n7426), .A2(n7425), .ZN(n14596) );
  NAND2_X1 U8898 ( .A1(n11530), .A2(n12031), .ZN(n14347) );
  NAND2_X1 U8899 ( .A1(n11431), .A2(n11430), .ZN(n11533) );
  NAND2_X1 U8900 ( .A1(n11363), .A2(n11362), .ZN(n11365) );
  NAND2_X1 U8901 ( .A1(n11172), .A2(n11171), .ZN(n12311) );
  NAND2_X1 U8902 ( .A1(n10967), .A2(n10966), .ZN(n11180) );
  NAND2_X1 U8903 ( .A1(n10905), .A2(n10805), .ZN(n10814) );
  NAND2_X1 U8904 ( .A1(n10808), .A2(n10807), .ZN(n15191) );
  NAND2_X1 U8905 ( .A1(n6896), .A2(n10494), .ZN(n10799) );
  OR2_X1 U8906 ( .A1(n10614), .A2(n10493), .ZN(n6896) );
  NAND2_X1 U8907 ( .A1(n6863), .A2(n11955), .ZN(n10112) );
  NAND2_X1 U8908 ( .A1(n7141), .A2(n9506), .ZN(n10111) );
  INV_X1 U8909 ( .A(n15093), .ZN(n15148) );
  NAND2_X1 U8910 ( .A1(n10052), .A2(n10108), .ZN(n14556) );
  AND2_X1 U8911 ( .A1(n11934), .A2(n11930), .ZN(n15130) );
  AND3_X2 U8912 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n15213) );
  XNOR2_X1 U8913 ( .A(n9434), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U8914 ( .A1(n9433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9434) );
  XNOR2_X1 U8915 ( .A(n9437), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U8916 ( .A1(n9443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9437) );
  INV_X1 U8917 ( .A(n9451), .ZN(n11871) );
  INV_X1 U8918 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14713) );
  NOR2_X1 U8919 ( .A1(n7540), .A2(n7539), .ZN(n7538) );
  OAI21_X1 U8920 ( .B1(n9433), .B2(P1_IR_REG_25__SCAN_IN), .A(n6687), .ZN(
        n7541) );
  NOR2_X1 U8921 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7539) );
  INV_X1 U8922 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U8923 ( .A1(n7389), .A2(n8395), .ZN(n8801) );
  INV_X1 U8924 ( .A(n9438), .ZN(n11617) );
  XNOR2_X1 U8925 ( .A(n8785), .B(n8784), .ZN(n12111) );
  NAND2_X1 U8926 ( .A1(n8387), .A2(n8768), .ZN(n8785) );
  INV_X1 U8927 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10872) );
  OR2_X1 U8928 ( .A1(n7384), .A2(n7383), .ZN(n8739) );
  NAND2_X1 U8929 ( .A1(n8382), .A2(n8380), .ZN(n8737) );
  INV_X1 U8930 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n12990) );
  INV_X1 U8931 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11167) );
  INV_X1 U8932 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9743) );
  INV_X1 U8933 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9719) );
  INV_X1 U8934 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9697) );
  CLKBUF_X1 U8935 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14721) );
  INV_X1 U8936 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14763) );
  XNOR2_X1 U8937 ( .A(n14764), .B(n6803), .ZN(n15643) );
  INV_X1 U8938 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6803) );
  XNOR2_X1 U8939 ( .A(n14758), .B(n7412), .ZN(n15633) );
  INV_X1 U8940 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7412) );
  XNOR2_X1 U8941 ( .A(n14777), .B(n7411), .ZN(n14840) );
  INV_X1 U8942 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7411) );
  INV_X1 U8943 ( .A(n14788), .ZN(n7392) );
  INV_X1 U8944 ( .A(n7397), .ZN(n14805) );
  XNOR2_X1 U8945 ( .A(n6928), .B(n6927), .ZN(n14862) );
  INV_X1 U8946 ( .A(n14863), .ZN(n6927) );
  OR2_X1 U8947 ( .A1(n12660), .A2(n15547), .ZN(n12661) );
  AOI21_X1 U8948 ( .B1(n12680), .B2(n15538), .A(n12679), .ZN(n7194) );
  NAND2_X1 U8949 ( .A1(n7197), .A2(n7196), .ZN(n7195) );
  INV_X1 U8950 ( .A(n8942), .ZN(n12695) );
  AOI21_X1 U8951 ( .B1(n11645), .B2(n9316), .A(n9315), .ZN(n9317) );
  OR2_X1 U8952 ( .A1(n8955), .A2(n13211), .ZN(n7641) );
  AOI21_X1 U8953 ( .B1(n11645), .B2(n9310), .A(n9309), .ZN(n9311) );
  OR2_X1 U8954 ( .A1(n8955), .A2(n13263), .ZN(n7642) );
  NAND2_X1 U8955 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n9657) );
  AOI21_X1 U8956 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13358) );
  NAND2_X1 U8957 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  OAI211_X1 U8958 ( .C1(n12437), .C2(n15316), .A(n6821), .B(n6819), .ZN(
        P2_U3236) );
  NOR2_X1 U8959 ( .A1(n6604), .A2(n12435), .ZN(n6821) );
  NAND2_X1 U8960 ( .A1(n6820), .A2(n15327), .ZN(n6819) );
  OAI21_X1 U8961 ( .B1(n7491), .B2(n7490), .A(n7487), .ZN(n7489) );
  INV_X1 U8962 ( .A(n7488), .ZN(n7487) );
  NAND2_X1 U8963 ( .A1(n6679), .A2(n6809), .ZN(P1_U3265) );
  INV_X1 U8964 ( .A(n6810), .ZN(n6809) );
  OAI21_X1 U8965 ( .B1(n14620), .B2(n15098), .A(n6811), .ZN(n6810) );
  NAND2_X1 U8966 ( .A1(n15200), .A2(n6917), .ZN(n6914) );
  INV_X1 U8967 ( .A(n6912), .ZN(n6911) );
  NOR2_X1 U8968 ( .A1(n14848), .A2(n14847), .ZN(n14846) );
  AND2_X1 U8969 ( .A1(n7409), .A2(n7408), .ZN(n14848) );
  NOR2_X1 U8970 ( .A1(n15021), .A2(n15022), .ZN(n15020) );
  INV_X1 U8971 ( .A(n6931), .ZN(n15021) );
  INV_X1 U8972 ( .A(n7403), .ZN(n15025) );
  AND2_X1 U8973 ( .A1(n7400), .A2(n7403), .ZN(n15028) );
  NOR2_X1 U8974 ( .A1(n7402), .A2(n15027), .ZN(n14860) );
  OR2_X1 U8975 ( .A1(n9010), .A2(n9012), .ZN(n6595) );
  AND2_X1 U8976 ( .A1(n11984), .A2(n11986), .ZN(n6596) );
  AND2_X1 U8977 ( .A1(n8915), .A2(n7273), .ZN(n6597) );
  INV_X2 U8978 ( .A(n9057), .ZN(n9132) );
  INV_X1 U8979 ( .A(n15585), .ZN(n6736) );
  INV_X1 U8980 ( .A(n11396), .ZN(n7517) );
  INV_X2 U8981 ( .A(n8437), .ZN(n6771) );
  OR2_X1 U8982 ( .A1(n14951), .A2(n11647), .ZN(n6598) );
  NAND2_X1 U8983 ( .A1(n7187), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6599) );
  INV_X1 U8984 ( .A(n12828), .ZN(n7552) );
  XNOR2_X1 U8985 ( .A(n12327), .B(n12326), .ZN(n6600) );
  AND2_X1 U8986 ( .A1(n6650), .A2(n7561), .ZN(n6601) );
  AND2_X1 U8987 ( .A1(n9625), .A2(n9680), .ZN(n6603) );
  INV_X1 U8988 ( .A(n13913), .ZN(n7274) );
  AND2_X1 U8989 ( .A1(n12436), .A2(n15326), .ZN(n6604) );
  AND2_X1 U8990 ( .A1(n9091), .A2(n9090), .ZN(n6605) );
  AND2_X1 U8991 ( .A1(n14520), .A2(n6907), .ZN(n6606) );
  INV_X1 U8992 ( .A(n13899), .ZN(n6774) );
  AND2_X1 U8993 ( .A1(n6909), .A2(n6907), .ZN(n6607) );
  AND2_X1 U8994 ( .A1(n8312), .A2(n11869), .ZN(n8428) );
  NAND2_X1 U8995 ( .A1(n7229), .A2(n9368), .ZN(n12542) );
  MUX2_X1 U8996 ( .A(n14394), .B(n14618), .S(n12241), .Z(n12193) );
  AND4_X1 U8997 ( .A1(n9515), .A2(n9514), .A3(n9513), .A4(n9512), .ZN(n11960)
         );
  NAND2_X1 U8998 ( .A1(n11164), .A2(n11163), .ZN(n12002) );
  AND2_X1 U8999 ( .A1(n7049), .A2(n7048), .ZN(n6608) );
  NOR2_X1 U9000 ( .A1(n12555), .A2(n7237), .ZN(n6609) );
  NOR2_X1 U9001 ( .A1(n8704), .A2(n7502), .ZN(n7498) );
  AND2_X1 U9002 ( .A1(n7505), .A2(n8602), .ZN(n6610) );
  OR2_X1 U9003 ( .A1(n11101), .A2(n12595), .ZN(n6611) );
  INV_X1 U9004 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U9005 ( .A1(n15022), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6612) );
  INV_X1 U9006 ( .A(n12211), .ZN(n7013) );
  AND2_X1 U9007 ( .A1(n7322), .A2(n13341), .ZN(n6613) );
  NOR2_X1 U9008 ( .A1(n8638), .A2(SI_14_), .ZN(n6614) );
  AND2_X1 U9009 ( .A1(n6926), .A2(n14818), .ZN(n6615) );
  NAND2_X1 U9010 ( .A1(n7956), .A2(n7663), .ZN(n7959) );
  OR2_X1 U9011 ( .A1(n8605), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6616) );
  AND2_X1 U9012 ( .A1(n9072), .A2(n9071), .ZN(n6617) );
  INV_X2 U9013 ( .A(n15455), .ZN(n15457) );
  NAND2_X1 U9014 ( .A1(n13885), .A2(n7039), .ZN(n7040) );
  AND2_X1 U9015 ( .A1(n11320), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6618) );
  INV_X1 U9016 ( .A(n11972), .ZN(n7090) );
  INV_X1 U9017 ( .A(n9032), .ZN(n9121) );
  OAI21_X2 U9018 ( .B1(n8437), .B2(n15228), .A(n7484), .ZN(n8968) );
  OR2_X1 U9019 ( .A1(n8059), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n6619) );
  OR2_X1 U9020 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n15017), .ZN(n6620) );
  INV_X1 U9021 ( .A(n12599), .ZN(n6737) );
  OR2_X1 U9022 ( .A1(n15220), .A2(n15219), .ZN(n6621) );
  INV_X1 U9023 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9436) );
  AND2_X1 U9024 ( .A1(n9625), .A2(n9681), .ZN(n6622) );
  OR2_X1 U9025 ( .A1(n13404), .A2(n13401), .ZN(n6623) );
  INV_X1 U9026 ( .A(n14387), .ZN(n6807) );
  INV_X1 U9027 ( .A(n7785), .ZN(n7203) );
  NAND2_X1 U9028 ( .A1(n14645), .A2(n14378), .ZN(n6624) );
  NAND4_X1 U9029 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n14172)
         );
  NOR2_X1 U9030 ( .A1(n10347), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9630) );
  OR2_X1 U9031 ( .A1(n13967), .A2(n9077), .ZN(n6625) );
  AND2_X1 U9032 ( .A1(n9687), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6626) );
  OR2_X1 U9033 ( .A1(n14511), .A2(n14645), .ZN(n6627) );
  INV_X1 U9034 ( .A(n6907), .ZN(n6906) );
  NOR2_X1 U9035 ( .A1(n14546), .A2(n6908), .ZN(n6907) );
  AND2_X1 U9036 ( .A1(n8932), .A2(n7580), .ZN(n6628) );
  XNOR2_X1 U9037 ( .A(n12701), .B(n12580), .ZN(n11815) );
  INV_X1 U9038 ( .A(n11815), .ZN(n6791) );
  AND2_X1 U9039 ( .A1(n8459), .A2(n6770), .ZN(n6629) );
  AND2_X1 U9040 ( .A1(n10134), .A2(n15485), .ZN(n6630) );
  AND2_X1 U9041 ( .A1(n14416), .A2(n14363), .ZN(n6631) );
  NAND2_X1 U9042 ( .A1(n14116), .A2(n12377), .ZN(n14035) );
  NAND2_X1 U9043 ( .A1(n14618), .A2(n14394), .ZN(n6632) );
  AND2_X1 U9044 ( .A1(n12247), .A2(n14364), .ZN(n14413) );
  INV_X1 U9045 ( .A(n14413), .ZN(n6827) );
  AND2_X1 U9046 ( .A1(n7305), .A2(n7308), .ZN(n8454) );
  OR2_X1 U9047 ( .A1(n11962), .A2(n11963), .ZN(n6633) );
  AND2_X1 U9048 ( .A1(n15504), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U9049 ( .A1(n14372), .A2(n14371), .ZN(n14552) );
  AND2_X1 U9050 ( .A1(n9358), .A2(n12588), .ZN(n6635) );
  INV_X1 U9051 ( .A(n14618), .ZN(n7101) );
  NAND2_X2 U9052 ( .A1(n8460), .A2(n6629), .ZN(n15318) );
  INV_X1 U9053 ( .A(n15318), .ZN(n7258) );
  AND3_X1 U9054 ( .A1(n7381), .A2(n12280), .A3(n14387), .ZN(n6636) );
  AND2_X1 U9055 ( .A1(n12594), .A2(n11273), .ZN(n6637) );
  AND4_X1 U9056 ( .A1(n7661), .A2(n7899), .A3(n7864), .A4(n7660), .ZN(n6638)
         );
  NAND2_X1 U9057 ( .A1(n9329), .A2(n15461), .ZN(n6639) );
  OR2_X1 U9058 ( .A1(n7043), .A2(n13905), .ZN(n6640) );
  OR2_X1 U9059 ( .A1(n13957), .A2(n13374), .ZN(n6641) );
  XNOR2_X1 U9060 ( .A(n14811), .B(n14810), .ZN(n6642) );
  NAND2_X1 U9061 ( .A1(n8541), .A2(n8540), .ZN(n13889) );
  NOR2_X1 U9062 ( .A1(n12584), .A2(n12528), .ZN(n6643) );
  NAND2_X1 U9063 ( .A1(n8680), .A2(n8679), .ZN(n13967) );
  OR2_X1 U9064 ( .A1(n14804), .A2(n14803), .ZN(n6644) );
  AND2_X1 U9065 ( .A1(n15504), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6645) );
  AND2_X1 U9066 ( .A1(n12835), .A2(n12847), .ZN(n6646) );
  OR2_X1 U9067 ( .A1(n9037), .A2(n9038), .ZN(n6647) );
  NAND2_X1 U9068 ( .A1(n12243), .A2(n12242), .ZN(n6648) );
  AND2_X1 U9069 ( .A1(n13482), .A2(n13343), .ZN(n6649) );
  AND4_X1 U9070 ( .A1(n7672), .A2(n7671), .A3(n7670), .A4(n8003), .ZN(n6650)
         );
  INV_X1 U9071 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7413) );
  AND2_X1 U9072 ( .A1(n13845), .A2(n13852), .ZN(n6651) );
  NAND2_X1 U9073 ( .A1(n11959), .A2(n11960), .ZN(n6652) );
  AND3_X1 U9074 ( .A1(n6944), .A2(n7066), .A3(n7067), .ZN(n6653) );
  AND2_X1 U9075 ( .A1(n13792), .A2(n11300), .ZN(n6654) );
  INV_X1 U9076 ( .A(n12279), .ZN(n14611) );
  AND2_X1 U9077 ( .A1(n13905), .A2(n13499), .ZN(n6655) );
  NOR2_X1 U9078 ( .A1(n12632), .A2(n12631), .ZN(n6656) );
  NAND2_X1 U9079 ( .A1(n12248), .A2(n14363), .ZN(n6872) );
  INV_X1 U9080 ( .A(n6872), .ZN(n14420) );
  INV_X1 U9081 ( .A(n12788), .ZN(n12796) );
  AND2_X1 U9082 ( .A1(n11790), .A2(n11791), .ZN(n12788) );
  AND2_X1 U9083 ( .A1(n14906), .A2(n12638), .ZN(n6657) );
  AND2_X1 U9084 ( .A1(n14540), .A2(n14526), .ZN(n6658) );
  AND2_X1 U9085 ( .A1(n11608), .A2(n11599), .ZN(n6659) );
  AND2_X1 U9086 ( .A1(n12365), .A2(n12362), .ZN(n6660) );
  AND2_X1 U9087 ( .A1(n11136), .A2(n11134), .ZN(n6661) );
  NOR2_X1 U9088 ( .A1(n14682), .A2(n14568), .ZN(n6662) );
  INV_X1 U9089 ( .A(n7537), .ZN(n7536) );
  NAND2_X1 U9090 ( .A1(n12325), .A2(n14107), .ZN(n7537) );
  OR2_X1 U9091 ( .A1(n14490), .A2(n14486), .ZN(n7146) );
  AND2_X1 U9092 ( .A1(n12017), .A2(n12011), .ZN(n12253) );
  AND2_X1 U9093 ( .A1(n7715), .A2(n7716), .ZN(n6664) );
  AND2_X1 U9094 ( .A1(n12404), .A2(n12403), .ZN(n6665) );
  AND2_X1 U9095 ( .A1(n12383), .A2(n12382), .ZN(n6666) );
  AND2_X1 U9096 ( .A1(n11767), .A2(n11768), .ZN(n12842) );
  OR2_X1 U9097 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6667) );
  INV_X1 U9098 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7715) );
  INV_X1 U9099 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7716) );
  OR2_X1 U9100 ( .A1(n12691), .A2(n9304), .ZN(n11818) );
  OR2_X1 U9101 ( .A1(n12109), .A2(n12108), .ZN(n6668) );
  NOR2_X1 U9102 ( .A1(n13981), .A2(n13784), .ZN(n6669) );
  NOR2_X1 U9103 ( .A1(n13957), .A2(n13504), .ZN(n6670) );
  AND2_X1 U9104 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6671) );
  NOR2_X1 U9105 ( .A1(n13962), .A2(n13475), .ZN(n6672) );
  NOR2_X1 U9106 ( .A1(n13920), .A2(n13500), .ZN(n6673) );
  INV_X1 U9107 ( .A(n7502), .ZN(n7501) );
  NOR2_X1 U9108 ( .A1(n13779), .A2(n13505), .ZN(n7502) );
  INV_X1 U9109 ( .A(n7296), .ZN(n7295) );
  OAI21_X1 U9110 ( .B1(n8896), .B2(n7297), .A(n8897), .ZN(n7296) );
  INV_X1 U9111 ( .A(n6895), .ZN(n6894) );
  NAND2_X1 U9112 ( .A1(n6898), .A2(n10494), .ZN(n6895) );
  AND2_X1 U9113 ( .A1(n11454), .A2(n13797), .ZN(n6674) );
  AND2_X1 U9114 ( .A1(n9015), .A2(n9014), .ZN(n6675) );
  OR2_X1 U9115 ( .A1(n14615), .A2(n15178), .ZN(n6676) );
  AND2_X1 U9116 ( .A1(n8569), .A2(SI_10_), .ZN(n6677) );
  AND2_X1 U9117 ( .A1(n8344), .A2(SI_8_), .ZN(n6678) );
  OR2_X1 U9118 ( .A1(n14621), .A2(n14601), .ZN(n6679) );
  AND2_X1 U9119 ( .A1(n9353), .A2(n12831), .ZN(n6681) );
  INV_X1 U9120 ( .A(n12499), .ZN(n7236) );
  AND2_X1 U9121 ( .A1(n8932), .A2(n6790), .ZN(n6682) );
  AND2_X1 U9122 ( .A1(n11761), .A2(n11762), .ZN(n12866) );
  INV_X1 U9123 ( .A(n7094), .ZN(n7093) );
  NAND2_X1 U9124 ( .A1(n7096), .A2(n7095), .ZN(n7094) );
  INV_X1 U9125 ( .A(n7321), .ZN(n7320) );
  NAND2_X1 U9126 ( .A1(n6623), .A2(n13359), .ZN(n7321) );
  INV_X1 U9127 ( .A(n7630), .ZN(n7629) );
  NAND2_X1 U9128 ( .A1(n8261), .A2(n7631), .ZN(n7630) );
  INV_X1 U9129 ( .A(n12272), .ZN(n11532) );
  INV_X1 U9130 ( .A(n7568), .ZN(n7567) );
  NAND2_X1 U9131 ( .A1(n11731), .A2(n6611), .ZN(n7568) );
  INV_X1 U9132 ( .A(n7342), .ZN(n7341) );
  NAND2_X1 U9133 ( .A1(n13429), .A2(n7343), .ZN(n7342) );
  OR2_X1 U9134 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7705), .ZN(n6683) );
  AND2_X1 U9135 ( .A1(n9337), .A2(n12596), .ZN(n6684) );
  AND2_X1 U9136 ( .A1(n9660), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U9137 ( .A1(n12858), .A2(n11558), .ZN(n6686) );
  AND2_X1 U9138 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n6687) );
  INV_X1 U9139 ( .A(n6884), .ZN(n6883) );
  NAND2_X1 U9140 ( .A1(n14451), .A2(n14359), .ZN(n6884) );
  AND2_X1 U9141 ( .A1(n9340), .A2(n12594), .ZN(n6688) );
  AND2_X1 U9142 ( .A1(n6899), .A2(n14354), .ZN(n6689) );
  NAND2_X1 U9143 ( .A1(n13925), .A2(n13632), .ZN(n6690) );
  INV_X1 U9144 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8242) );
  MUX2_X1 U9145 ( .A(n14394), .B(n14618), .S(n12228), .Z(n12191) );
  INV_X1 U9146 ( .A(n7288), .ZN(n6960) );
  OR2_X1 U9147 ( .A1(n13673), .A2(n13466), .ZN(n7288) );
  AND3_X1 U9148 ( .A1(n11830), .A2(n11676), .A3(n7200), .ZN(n6691) );
  OR2_X1 U9149 ( .A1(n14736), .A2(n14735), .ZN(n6692) );
  OR2_X1 U9150 ( .A1(n14729), .A2(n7413), .ZN(n6693) );
  INV_X1 U9151 ( .A(n8994), .ZN(n7622) );
  AND2_X1 U9152 ( .A1(n7376), .A2(n7377), .ZN(n6694) );
  NOR2_X1 U9153 ( .A1(n11748), .A2(n11756), .ZN(n6695) );
  INV_X1 U9154 ( .A(n9114), .ZN(n7617) );
  NOR2_X1 U9155 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6696) );
  AND2_X1 U9156 ( .A1(n7037), .A2(n7036), .ZN(n6697) );
  INV_X1 U9157 ( .A(n8887), .ZN(n7265) );
  AND2_X1 U9158 ( .A1(n7099), .A2(n14606), .ZN(n6698) );
  AND2_X1 U9159 ( .A1(n7778), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6699) );
  AND2_X1 U9160 ( .A1(n7778), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6700) );
  INV_X1 U9161 ( .A(n9382), .ZN(n7237) );
  NOR2_X1 U9162 ( .A1(n14860), .A2(n14859), .ZN(n6701) );
  AND2_X1 U9163 ( .A1(n7778), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U9164 ( .A1(n9339), .A2(n10927), .ZN(n6703) );
  AND2_X1 U9165 ( .A1(n7713), .A2(n6664), .ZN(n6704) );
  AND2_X1 U9166 ( .A1(n14471), .A2(n14359), .ZN(n6705) );
  NAND2_X1 U9167 ( .A1(n14725), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6706) );
  AND2_X1 U9168 ( .A1(n6889), .A2(n6888), .ZN(n6707) );
  NOR2_X1 U9169 ( .A1(n8651), .A2(n7469), .ZN(n6708) );
  INV_X1 U9170 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8414) );
  OR2_X1 U9171 ( .A1(n15404), .A2(n13509), .ZN(n6709) );
  INV_X1 U9172 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8261) );
  OR2_X1 U9173 ( .A1(n9093), .A2(n6605), .ZN(n6710) );
  INV_X1 U9174 ( .A(n7136), .ZN(n7135) );
  AOI22_X1 U9175 ( .A1(n9680), .A2(SI_1_), .B1(n9681), .B2(n9665), .ZN(n7136)
         );
  NAND2_X1 U9176 ( .A1(n11985), .A2(n7434), .ZN(n6711) );
  NAND2_X1 U9177 ( .A1(n11974), .A2(n7437), .ZN(n6712) );
  OR2_X1 U9178 ( .A1(n13570), .A2(n13569), .ZN(P2_U3233) );
  NAND2_X2 U9179 ( .A1(n8437), .A2(n9681), .ZN(n8740) );
  AND2_X1 U9180 ( .A1(n7690), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6714) );
  INV_X1 U9181 ( .A(n11777), .ZN(n7559) );
  INV_X1 U9182 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U9183 ( .A1(n10301), .A2(n9542), .ZN(n10304) );
  OR2_X1 U9184 ( .A1(n8677), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U9185 ( .A1(n13498), .A2(n13854), .B1(n13573), .B2(n13496), .ZN(
        n8873) );
  INV_X1 U9186 ( .A(SI_14_), .ZN(n9749) );
  NOR2_X1 U9187 ( .A1(n8605), .A2(n7351), .ZN(n8653) );
  INV_X1 U9188 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7354) );
  NAND2_X1 U9189 ( .A1(n8836), .A2(n8835), .ZN(n13633) );
  OR2_X1 U9190 ( .A1(n14842), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7409) );
  INV_X1 U9191 ( .A(n7104), .ZN(n14583) );
  NAND2_X1 U9192 ( .A1(n8319), .A2(n8318), .ZN(n13498) );
  NAND2_X1 U9193 ( .A1(n13788), .A2(n7051), .ZN(n7052) );
  AND2_X1 U9194 ( .A1(n7350), .A2(n7348), .ZN(n6716) );
  NAND2_X1 U9195 ( .A1(n7615), .A2(n7617), .ZN(n7614) );
  INV_X1 U9196 ( .A(n7614), .ZN(n7609) );
  AND2_X1 U9197 ( .A1(n8004), .A2(n8003), .ZN(n7666) );
  AND2_X1 U9198 ( .A1(n7151), .A2(n7150), .ZN(n6717) );
  AND2_X1 U9199 ( .A1(n13818), .A2(n8602), .ZN(n6718) );
  NAND2_X1 U9200 ( .A1(n6589), .A2(n8260), .ZN(n8265) );
  INV_X1 U9201 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8236) );
  INV_X1 U9202 ( .A(n9073), .ZN(n7620) );
  NAND2_X1 U9203 ( .A1(n11504), .A2(n6983), .ZN(n6719) );
  INV_X1 U9204 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U9205 ( .A1(n14832), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6720) );
  OR2_X1 U9206 ( .A1(n7620), .A2(n6617), .ZN(n6721) );
  NAND2_X2 U9207 ( .A1(n10316), .A2(n15553), .ZN(n15566) );
  INV_X1 U9208 ( .A(n14959), .ZN(n15327) );
  XNOR2_X1 U9209 ( .A(n8182), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8198) );
  INV_X1 U9210 ( .A(n8430), .ZN(n9158) );
  INV_X1 U9211 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6851) );
  INV_X1 U9212 ( .A(n13799), .ZN(n7505) );
  NAND2_X1 U9213 ( .A1(n8693), .A2(n8692), .ZN(n13962) );
  INV_X1 U9214 ( .A(n13962), .ZN(n7048) );
  NAND2_X1 U9215 ( .A1(n8755), .A2(n8754), .ZN(n13943) );
  INV_X1 U9216 ( .A(n13943), .ZN(n7034) );
  OR2_X1 U9217 ( .A1(n9640), .A2(n7134), .ZN(n15541) );
  AND2_X1 U9218 ( .A1(n11883), .A2(n7359), .ZN(n6722) );
  INV_X1 U9219 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U9220 ( .A1(n7541), .A2(n7538), .ZN(n12298) );
  INV_X1 U9221 ( .A(n12298), .ZN(n6818) );
  INV_X1 U9222 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11036) );
  AND2_X1 U9223 ( .A1(n6962), .A2(n8196), .ZN(n9319) );
  INV_X1 U9224 ( .A(n14677), .ZN(n7103) );
  AND2_X1 U9225 ( .A1(n12617), .A2(n12619), .ZN(n6723) );
  NAND2_X1 U9226 ( .A1(n11528), .A2(n11527), .ZN(n14686) );
  INV_X1 U9227 ( .A(n14686), .ZN(n7105) );
  AND2_X1 U9228 ( .A1(n9354), .A2(n12509), .ZN(n6724) );
  NAND2_X1 U9229 ( .A1(n10912), .A2(n7093), .ZN(n7097) );
  NAND2_X1 U9230 ( .A1(n10945), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6725) );
  AND2_X1 U9231 ( .A1(n7569), .A2(n6611), .ZN(n6726) );
  AND2_X1 U9232 ( .A1(n7714), .A2(n8177), .ZN(n8215) );
  INV_X1 U9233 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13072) );
  INV_X1 U9234 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10277) );
  INV_X1 U9235 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10919) );
  OR2_X1 U9236 ( .A1(n15457), .A2(n12978), .ZN(n6727) );
  INV_X1 U9237 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U9238 ( .A1(n8398), .A2(n8397), .ZN(n6728) );
  OR2_X1 U9239 ( .A1(n10304), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6729) );
  AND2_X1 U9240 ( .A1(n9553), .A2(n9552), .ZN(n15178) );
  INV_X1 U9241 ( .A(n13279), .ZN(n7134) );
  INV_X1 U9242 ( .A(n12600), .ZN(n7247) );
  INV_X1 U9243 ( .A(n8055), .ZN(n7218) );
  CLKBUF_X1 U9244 ( .A(n15464), .Z(n6800) );
  NAND2_X1 U9245 ( .A1(n10955), .A2(n10954), .ZN(n15005) );
  INV_X1 U9246 ( .A(n15005), .ZN(n7095) );
  OAI22_X1 U9247 ( .A1(n15460), .A2(n15459), .B1(n6822), .B2(n9327), .ZN(n9650) );
  NAND2_X1 U9248 ( .A1(n10458), .A2(n9531), .ZN(n12256) );
  INV_X1 U9249 ( .A(n12256), .ZN(n6864) );
  NOR2_X1 U9250 ( .A1(n15516), .A2(n9637), .ZN(n6730) );
  NAND2_X1 U9251 ( .A1(n10117), .A2(n10593), .ZN(n10476) );
  INV_X1 U9252 ( .A(n10476), .ZN(n7091) );
  AND2_X1 U9253 ( .A1(n7192), .A2(n7191), .ZN(n6731) );
  OR2_X1 U9254 ( .A1(n7076), .A2(n7073), .ZN(n6732) );
  AND2_X1 U9255 ( .A1(n11429), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U9256 ( .A1(n7076), .A2(n7074), .ZN(n6734) );
  INV_X1 U9257 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11618) );
  INV_X1 U9258 ( .A(n12649), .ZN(n7055) );
  INV_X1 U9259 ( .A(n12648), .ZN(n7059) );
  INV_X1 U9260 ( .A(n12673), .ZN(n8115) );
  INV_X1 U9261 ( .A(n15178), .ZN(n6917) );
  INV_X1 U9262 ( .A(n6590), .ZN(n7137) );
  INV_X1 U9263 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14870) );
  INV_X1 U9264 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6918) );
  INV_X1 U9265 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14725) );
  INV_X1 U9266 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n7058) );
  AND2_X1 U9267 ( .A1(n9163), .A2(n8874), .ZN(n10173) );
  AOI21_X1 U9268 ( .B1(n12618), .B2(n12617), .A(n12619), .ZN(n12620) );
  OR2_X1 U9269 ( .A1(n12618), .A2(n12619), .ZN(n7182) );
  OR2_X1 U9270 ( .A1(n12617), .A2(n12619), .ZN(n7183) );
  INV_X1 U9271 ( .A(n8078), .ZN(n6856) );
  NAND2_X2 U9272 ( .A1(n9681), .A2(P2_U3088), .ZN(n14024) );
  INV_X1 U9273 ( .A(n15326), .ZN(n13886) );
  AND2_X2 U9274 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  OAI21_X2 U9275 ( .B1(n14490), .B2(n7144), .A(n7142), .ZN(n14456) );
  NAND2_X1 U9276 ( .A1(n14052), .A2(n12355), .ZN(n14099) );
  NAND2_X1 U9277 ( .A1(n10752), .A2(n10751), .ZN(n10889) );
  NAND2_X2 U9278 ( .A1(n12391), .A2(n12390), .ZN(n14067) );
  NAND2_X1 U9279 ( .A1(n14044), .A2(n14043), .ZN(n14042) );
  NAND2_X1 U9280 ( .A1(n10038), .A2(n10037), .ZN(n10064) );
  NAND2_X1 U9281 ( .A1(n7941), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U9282 ( .A1(n12720), .A2(n12719), .ZN(n12718) );
  NAND2_X2 U9283 ( .A1(n11929), .A2(n10056), .ZN(n12370) );
  NAND2_X1 U9284 ( .A1(n7774), .A2(n7772), .ZN(n7204) );
  NAND3_X1 U9285 ( .A1(n7556), .A2(n7555), .A3(n12796), .ZN(n12790) );
  NAND2_X1 U9286 ( .A1(n8054), .A2(n12788), .ZN(n12793) );
  NAND2_X1 U9287 ( .A1(n11521), .A2(n11748), .ZN(n11568) );
  AND2_X2 U9288 ( .A1(n7936), .A2(n7662), .ZN(n7955) );
  AND2_X2 U9289 ( .A1(n6858), .A2(n7659), .ZN(n7936) );
  NAND2_X1 U9290 ( .A1(n6740), .A2(n11710), .ZN(n10976) );
  NAND2_X1 U9291 ( .A1(n11206), .A2(n11734), .ZN(n11312) );
  NAND2_X1 U9292 ( .A1(n12743), .A2(n11803), .ZN(n12725) );
  NAND2_X1 U9293 ( .A1(n10873), .A2(n11662), .ZN(n6740) );
  NAND2_X1 U9294 ( .A1(n6823), .A2(n6791), .ZN(n7635) );
  OAI21_X1 U9295 ( .B1(n6744), .B2(n11704), .A(n6742), .ZN(n6741) );
  NAND3_X1 U9296 ( .A1(n7770), .A2(n7769), .A3(n6745), .ZN(n12601) );
  MUX2_X1 U9297 ( .A(n11755), .B(n11754), .S(n8226), .Z(n11760) );
  INV_X1 U9298 ( .A(n11699), .ZN(n6749) );
  INV_X1 U9299 ( .A(n11695), .ZN(n6751) );
  OAI21_X1 U9300 ( .B1(n11684), .B2(n11683), .A(n11686), .ZN(n11691) );
  OAI22_X1 U9301 ( .A1(n11743), .A2(n11742), .B1(n11795), .B2(n11741), .ZN(
        n11747) );
  NAND2_X1 U9302 ( .A1(n6754), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6753) );
  INV_X2 U9303 ( .A(n8124), .ZN(n15555) );
  OAI21_X2 U9304 ( .B1(n12767), .B2(n7123), .A(n7120), .ZN(n12743) );
  NAND2_X1 U9305 ( .A1(n11570), .A2(n11755), .ZN(n12867) );
  NAND2_X1 U9306 ( .A1(n7782), .A2(n7781), .ZN(n6859) );
  AOI22_X1 U9307 ( .A1(n14027), .A2(n14028), .B1(n12410), .B2(n12409), .ZN(
        n12418) );
  INV_X2 U9308 ( .A(n7654), .ZN(n12198) );
  NAND2_X1 U9309 ( .A1(n8015), .A2(n11778), .ZN(n12820) );
  INV_X2 U9310 ( .A(n9625), .ZN(n8038) );
  NAND2_X1 U9311 ( .A1(n8841), .A2(n8403), .ZN(n7387) );
  NAND2_X1 U9312 ( .A1(n6945), .A2(n6946), .ZN(n8585) );
  OAI21_X1 U9313 ( .B1(n8689), .B2(n8370), .A(n8687), .ZN(n8372) );
  NAND2_X1 U9314 ( .A1(n7765), .A2(n7760), .ZN(n7676) );
  NAND3_X1 U9315 ( .A1(n6691), .A2(n6845), .A3(n6598), .ZN(n7199) );
  NOR2_X1 U9316 ( .A1(n10074), .A2(n10034), .ZN(n10040) );
  NOR2_X1 U9317 ( .A1(n10535), .A2(n10534), .ZN(n14044) );
  NAND2_X1 U9318 ( .A1(n7699), .A2(n6831), .ZN(n7990) );
  NAND2_X1 U9319 ( .A1(n7702), .A2(n6850), .ZN(n8018) );
  NAND2_X1 U9320 ( .A1(n14042), .A2(n7546), .ZN(n10586) );
  NOR2_X1 U9321 ( .A1(n10066), .A2(n10065), .ZN(n10069) );
  NAND2_X1 U9322 ( .A1(n6798), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U9323 ( .A1(n8066), .A2(n8065), .ZN(n12767) );
  OAI21_X2 U9324 ( .B1(n14582), .B2(n6662), .A(n14368), .ZN(n14565) );
  NAND2_X1 U9325 ( .A1(n9492), .A2(n9491), .ZN(n10278) );
  NAND2_X1 U9326 ( .A1(n10817), .A2(n10816), .ZN(n10903) );
  NAND2_X1 U9327 ( .A1(n11249), .A2(n11165), .ZN(n11179) );
  NAND2_X1 U9328 ( .A1(n14456), .A2(n14455), .ZN(n14454) );
  NAND2_X1 U9329 ( .A1(n10952), .A2(n10951), .ZN(n10957) );
  NAND2_X1 U9330 ( .A1(n10473), .A2(n10472), .ZN(n10475) );
  OAI21_X1 U9331 ( .B1(n11363), .B2(n7156), .A(n7154), .ZN(n11534) );
  NAND2_X1 U9332 ( .A1(n11250), .A2(n12270), .ZN(n11249) );
  NAND2_X1 U9333 ( .A1(n10957), .A2(n10956), .ZN(n11160) );
  INV_X1 U9334 ( .A(n6812), .ZN(n14621) );
  AOI22_X1 U9335 ( .A1(n9876), .A2(n9875), .B1(n9849), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n9973) );
  AOI21_X1 U9336 ( .B1(n9853), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9956), .ZN(
        n9860) );
  NAND2_X1 U9337 ( .A1(n14517), .A2(n14375), .ZN(n14510) );
  NAND2_X1 U9338 ( .A1(n10278), .A2(n10279), .ZN(n7141) );
  NAND2_X1 U9339 ( .A1(n6760), .A2(n14522), .ZN(n14517) );
  NAND2_X1 U9340 ( .A1(n8379), .A2(n8378), .ZN(n6956) );
  INV_X1 U9341 ( .A(n14519), .ZN(n6760) );
  NAND2_X1 U9342 ( .A1(n14454), .A2(n14382), .ZN(n14435) );
  INV_X1 U9343 ( .A(n14490), .ZN(n14492) );
  NAND2_X1 U9344 ( .A1(n9532), .A2(n12256), .ZN(n10473) );
  NAND2_X1 U9345 ( .A1(n9547), .A2(n15133), .ZN(n11924) );
  NAND2_X1 U9346 ( .A1(n10393), .A2(n10392), .ZN(n15220) );
  NAND2_X1 U9347 ( .A1(n13294), .A2(n13293), .ZN(n13418) );
  NAND2_X1 U9348 ( .A1(n11290), .A2(n11232), .ZN(n11298) );
  OAI21_X2 U9349 ( .B1(n13474), .B2(n13473), .A(n13311), .ZN(n13448) );
  NAND2_X1 U9350 ( .A1(n8750), .A2(n8385), .ZN(n8386) );
  OAI21_X1 U9351 ( .B1(n8813), .B2(n8812), .A(n6728), .ZN(n6826) );
  NAND2_X1 U9352 ( .A1(n8390), .A2(n8389), .ZN(n8392) );
  NAND2_X1 U9353 ( .A1(n7272), .A2(n7271), .ZN(n13590) );
  NAND2_X1 U9354 ( .A1(n6761), .A2(n12210), .ZN(n12213) );
  NAND2_X1 U9355 ( .A1(n7012), .A2(n7015), .ZN(n6761) );
  OAI21_X2 U9356 ( .B1(n8458), .B2(n8457), .A(n8326), .ZN(n8469) );
  INV_X1 U9357 ( .A(n7016), .ZN(n7014) );
  NAND2_X1 U9358 ( .A1(n8752), .A2(n8751), .ZN(n8750) );
  INV_X1 U9359 ( .A(n6826), .ZN(n8823) );
  NAND2_X2 U9360 ( .A1(n12190), .A2(n12189), .ZN(n14618) );
  NAND3_X1 U9361 ( .A1(n6764), .A2(n6763), .A3(n7446), .ZN(n12192) );
  NAND3_X1 U9362 ( .A1(n12166), .A2(n12165), .A3(n12181), .ZN(n6763) );
  NAND3_X1 U9363 ( .A1(n12166), .A2(n12165), .A3(n12179), .ZN(n6764) );
  NAND3_X1 U9364 ( .A1(n12010), .A2(n12009), .A3(n6768), .ZN(n12021) );
  AOI21_X1 U9365 ( .B1(n12108), .B2(n12109), .A(n12106), .ZN(n12107) );
  NAND2_X1 U9366 ( .A1(n8568), .A2(n8567), .ZN(n13834) );
  NAND2_X1 U9367 ( .A1(n7464), .A2(n6708), .ZN(n7463) );
  NAND2_X1 U9368 ( .A1(n13583), .A2(n6773), .ZN(n6772) );
  OAI22_X1 U9369 ( .A1(n10664), .A2(n8535), .B1(n13875), .B2(n15404), .ZN(
        n13871) );
  NAND2_X1 U9370 ( .A1(n15311), .A2(n7257), .ZN(n8462) );
  NAND2_X1 U9371 ( .A1(n6769), .A2(n15444), .ZN(n6958) );
  NAND2_X1 U9372 ( .A1(n12437), .A2(n7492), .ZN(n6769) );
  XNOR2_X1 U9373 ( .A(n13513), .B(n10712), .ZN(n9238) );
  INV_X1 U9374 ( .A(n6775), .ZN(n9069) );
  NAND2_X1 U9375 ( .A1(n9022), .A2(n9021), .ZN(n9027) );
  OAI21_X1 U9376 ( .B1(n7627), .B2(n7625), .A(n7624), .ZN(n9037) );
  AND2_X2 U9377 ( .A1(n9502), .A2(n15648), .ZN(n9714) );
  NAND2_X1 U9378 ( .A1(n9548), .A2(n11942), .ZN(n10447) );
  NAND2_X1 U9379 ( .A1(n10618), .A2(n10510), .ZN(n10511) );
  INV_X1 U9380 ( .A(n14173), .ZN(n11938) );
  NAND4_X1 U9381 ( .A1(n9456), .A2(n9457), .A3(n9455), .A4(n9454), .ZN(n14173)
         );
  NAND2_X1 U9383 ( .A1(n10616), .A2(n10615), .ZN(n10618) );
  NAND2_X1 U9384 ( .A1(n12092), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U9385 ( .A1(n9235), .A2(n7648), .ZN(n9270) );
  NAND2_X1 U9386 ( .A1(n8980), .A2(n6663), .ZN(n8987) );
  NAND2_X1 U9387 ( .A1(n8965), .A2(n8964), .ZN(n8971) );
  NAND2_X1 U9388 ( .A1(n9111), .A2(n9110), .ZN(n9116) );
  OAI21_X1 U9389 ( .B1(n9013), .B2(n7600), .A(n6595), .ZN(n9019) );
  INV_X1 U9390 ( .A(n7168), .ZN(n7167) );
  NAND2_X1 U9391 ( .A1(n7527), .A2(n12398), .ZN(n14138) );
  OAI21_X2 U9392 ( .B1(n10747), .B2(n10746), .A(n10745), .ZN(n10752) );
  NAND2_X1 U9393 ( .A1(n14367), .A2(n14366), .ZN(n14582) );
  NAND2_X1 U9394 ( .A1(n7587), .A2(n7590), .ZN(n9068) );
  AOI21_X1 U9395 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n7627) );
  NAND2_X1 U9396 ( .A1(n6630), .A2(n10135), .ZN(n7083) );
  AOI21_X1 U9397 ( .B1(n9088), .B2(n9087), .A(n9085), .ZN(n9086) );
  NAND2_X1 U9398 ( .A1(n6680), .A2(n9082), .ZN(n9088) );
  NAND2_X1 U9399 ( .A1(n9002), .A2(n9003), .ZN(n9001) );
  OR2_X2 U9400 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U9401 ( .A1(n6780), .A2(n6647), .ZN(n9045) );
  INV_X1 U9402 ( .A(n6781), .ZN(n6780) );
  AOI21_X1 U9403 ( .B1(n9037), .B2(n9038), .A(n9039), .ZN(n6781) );
  NOR2_X1 U9404 ( .A1(n14883), .A2(n12629), .ZN(n14908) );
  NOR2_X1 U9405 ( .A1(n11059), .A2(n11060), .ZN(n11063) );
  NAND2_X1 U9406 ( .A1(n7054), .A2(n6720), .ZN(n10421) );
  NAND2_X1 U9407 ( .A1(n11179), .A2(n12269), .ZN(n11363) );
  NAND2_X1 U9408 ( .A1(n10889), .A2(n10888), .ZN(n10894) );
  INV_X1 U9409 ( .A(n7081), .ZN(n9635) );
  NAND2_X1 U9410 ( .A1(n12632), .A2(n7069), .ZN(n6944) );
  NAND2_X1 U9411 ( .A1(n7618), .A2(n7619), .ZN(n9081) );
  NOR2_X1 U9412 ( .A1(n10211), .A2(n10196), .ZN(n10326) );
  NOR2_X1 U9413 ( .A1(n15475), .A2(n9634), .ZN(n15498) );
  NAND2_X1 U9414 ( .A1(n9637), .A2(n7080), .ZN(n7078) );
  NAND2_X2 U9415 ( .A1(n8913), .A2(n8912), .ZN(n13618) );
  NAND2_X2 U9416 ( .A1(n13769), .A2(n8898), .ZN(n13760) );
  NAND2_X2 U9417 ( .A1(n8910), .A2(n8909), .ZN(n13669) );
  OAI21_X1 U9418 ( .B1(n11218), .B2(n7358), .A(n7355), .ZN(n11290) );
  OAI21_X1 U9419 ( .B1(n11298), .B2(n11297), .A(n11296), .ZN(n11491) );
  NAND2_X4 U9420 ( .A1(n13879), .A2(n8960), .ZN(n13384) );
  NAND3_X1 U9421 ( .A1(n6676), .A2(n14616), .A3(n14614), .ZN(n14695) );
  NAND2_X1 U9422 ( .A1(n10698), .A2(n10697), .ZN(n7460) );
  AOI21_X1 U9423 ( .B1(n8443), .B2(n8442), .A(n8323), .ZN(n8458) );
  NAND2_X1 U9424 ( .A1(n6784), .A2(n11720), .ZN(n11726) );
  NAND2_X1 U9425 ( .A1(n6785), .A2(n6840), .ZN(n6839) );
  NAND3_X1 U9426 ( .A1(n11793), .A2(n11794), .A3(n11792), .ZN(n6785) );
  NAND2_X1 U9427 ( .A1(n6844), .A2(n11830), .ZN(n11832) );
  OAI21_X1 U9428 ( .B1(n11697), .B2(n11795), .A(n6841), .ZN(n11705) );
  NAND2_X1 U9429 ( .A1(n12706), .A2(n11812), .ZN(n6823) );
  NOR2_X1 U9430 ( .A1(n6569), .A2(n7761), .ZN(n6789) );
  NAND2_X1 U9431 ( .A1(n6568), .A2(n7767), .ZN(n9321) );
  INV_X1 U9432 ( .A(n11405), .ZN(n8143) );
  INV_X1 U9433 ( .A(n8163), .ZN(n6792) );
  NAND2_X1 U9434 ( .A1(n8128), .A2(n8127), .ZN(n10992) );
  NOR2_X1 U9435 ( .A1(n6700), .A2(n6789), .ZN(n6788) );
  NAND2_X1 U9436 ( .A1(n7548), .A2(n7550), .ZN(n12814) );
  INV_X1 U9437 ( .A(n6852), .ZN(n7643) );
  NAND3_X1 U9438 ( .A1(n8134), .A2(n10975), .A3(n7564), .ZN(n8137) );
  NAND2_X1 U9439 ( .A1(n7239), .A2(n7240), .ZN(n11080) );
  NAND2_X1 U9440 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NAND2_X1 U9441 ( .A1(n6574), .A2(n11686), .ZN(n7129) );
  NAND2_X2 U9442 ( .A1(n6799), .A2(n6794), .ZN(n15461) );
  NAND2_X2 U9443 ( .A1(n12565), .A2(n12564), .ZN(n12563) );
  NAND2_X1 U9444 ( .A1(n6986), .A2(n6985), .ZN(n9342) );
  AOI21_X1 U9445 ( .B1(n10546), .B2(n10545), .A(n7245), .ZN(n10608) );
  NAND2_X1 U9446 ( .A1(n7393), .A2(n6921), .ZN(n6920) );
  INV_X1 U9447 ( .A(n6919), .ZN(n14730) );
  NAND2_X1 U9448 ( .A1(n6924), .A2(n6922), .ZN(n6928) );
  NOR2_X1 U9449 ( .A1(n14732), .A2(n14731), .ZN(n14779) );
  NOR2_X1 U9450 ( .A1(n14733), .A2(n6937), .ZN(n14736) );
  XNOR2_X1 U9451 ( .A(n14736), .B(n14735), .ZN(n14782) );
  NAND2_X1 U9452 ( .A1(n7933), .A2(n7931), .ZN(n7695) );
  NAND2_X1 U9453 ( .A1(n7692), .A2(n7691), .ZN(n7933) );
  NAND2_X1 U9454 ( .A1(n7822), .A2(n7820), .ZN(n7216) );
  AOI21_X2 U9455 ( .B1(n7745), .B2(n7708), .A(n7228), .ZN(n8100) );
  XNOR2_X1 U9456 ( .A(n7199), .B(n12673), .ZN(n7652) );
  OAI22_X1 U9457 ( .A1(n9291), .A2(n9292), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(
        n14012), .ZN(n11621) );
  NAND2_X1 U9458 ( .A1(n8018), .A2(n8016), .ZN(n7704) );
  AOI21_X1 U9459 ( .B1(n8923), .B2(n8924), .A(n7227), .ZN(n9291) );
  XNOR2_X1 U9460 ( .A(n11626), .B(n6797), .ZN(n12428) );
  NAND2_X1 U9461 ( .A1(n11621), .A2(n11622), .ZN(n7226) );
  NAND2_X1 U9462 ( .A1(n11312), .A2(n11311), .ZN(n11310) );
  NAND2_X1 U9463 ( .A1(n10577), .A2(n10576), .ZN(n11214) );
  AOI21_X1 U9464 ( .B1(n7402), .B2(n6923), .A(n6615), .ZN(n6922) );
  NAND2_X1 U9465 ( .A1(n15632), .A2(n15633), .ZN(n6802) );
  XNOR2_X1 U9466 ( .A(n14787), .B(n7392), .ZN(n14841) );
  OAI21_X1 U9467 ( .B1(n12370), .B2(n6817), .A(n6816), .ZN(n6815) );
  NOR2_X1 U9468 ( .A1(n10069), .A2(n10068), .ZN(n10535) );
  NAND3_X2 U9469 ( .A1(n6805), .A2(n9460), .A3(n6667), .ZN(n14187) );
  NAND2_X1 U9470 ( .A1(n12328), .A2(n14147), .ZN(n14075) );
  OAI21_X1 U9471 ( .B1(n10038), .B2(n10037), .A(n10064), .ZN(n10039) );
  AOI21_X1 U9472 ( .B1(n14423), .B2(n14386), .A(n6827), .ZN(n14414) );
  INV_X1 U9473 ( .A(n9494), .ZN(n9511) );
  AOI21_X1 U9474 ( .B1(n14423), .B2(n7163), .A(n14414), .ZN(n6812) );
  NAND2_X1 U9475 ( .A1(n9480), .A2(n9479), .ZN(n15078) );
  NAND2_X1 U9476 ( .A1(n15293), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15292) );
  XNOR2_X1 U9477 ( .A(n10706), .B(n6814), .ZN(n10697) );
  INV_X1 U9478 ( .A(n6815), .ZN(n10076) );
  NAND3_X2 U9479 ( .A1(n6818), .A2(n9439), .A3(n9438), .ZN(n10056) );
  OAI21_X2 U9480 ( .B1(n13613), .B2(n7472), .A(n7470), .ZN(n13585) );
  NAND2_X1 U9481 ( .A1(n7463), .A2(n7461), .ZN(n8667) );
  NAND2_X1 U9482 ( .A1(n8933), .A2(n12441), .ZN(n8934) );
  NAND2_X1 U9483 ( .A1(n7990), .A2(n7988), .ZN(n7701) );
  NAND2_X2 U9484 ( .A1(n13707), .A2(n8749), .ZN(n13696) );
  NAND2_X1 U9485 ( .A1(n11310), .A2(n11740), .ZN(n11411) );
  NAND2_X1 U9486 ( .A1(n7890), .A2(n11728), .ZN(n11207) );
  NAND2_X4 U9487 ( .A1(n7718), .A2(n7729), .ZN(n13279) );
  INV_X1 U9488 ( .A(n7077), .ZN(n6828) );
  NAND2_X1 U9489 ( .A1(n8113), .A2(n7635), .ZN(n12696) );
  OR4_X1 U9490 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12273) );
  INV_X1 U9491 ( .A(n12288), .ZN(n7008) );
  XNOR2_X1 U9492 ( .A(n8362), .B(n9749), .ZN(n8639) );
  INV_X1 U9493 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7719) );
  AOI21_X1 U9494 ( .B1(n6870), .B2(n6873), .A(n6868), .ZN(n6867) );
  AOI21_X2 U9495 ( .B1(n8669), .B2(n8369), .A(n8368), .ZN(n8689) );
  NAND2_X1 U9496 ( .A1(n7373), .A2(n7372), .ZN(n8620) );
  NAND2_X1 U9497 ( .A1(n6954), .A2(n6953), .ZN(n8752) );
  NAND2_X1 U9498 ( .A1(n15078), .A2(n15077), .ZN(n9492) );
  INV_X1 U9499 ( .A(n10454), .ZN(n9478) );
  OAI21_X1 U9500 ( .B1(n11829), .B2(n6846), .A(n6845), .ZN(n6844) );
  OAI21_X1 U9501 ( .B1(n11811), .B2(n12719), .A(n6838), .ZN(n6837) );
  NAND2_X1 U9502 ( .A1(n6837), .A2(n11814), .ZN(n11816) );
  NAND2_X1 U9503 ( .A1(n7695), .A2(n7694), .ZN(n7696) );
  XNOR2_X1 U9504 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7760) );
  NOR2_X1 U9505 ( .A1(n14877), .A2(n14878), .ZN(n14876) );
  NAND2_X1 U9506 ( .A1(n7178), .A2(n7176), .ZN(n12676) );
  NOR2_X1 U9507 ( .A1(n11051), .A2(n11052), .ZN(n11056) );
  NOR2_X1 U9508 ( .A1(n10759), .A2(n10760), .ZN(n10763) );
  XNOR2_X1 U9509 ( .A(n12678), .B(n12677), .ZN(n7197) );
  XNOR2_X2 U9510 ( .A(n7801), .B(n7800), .ZN(n15504) );
  NAND3_X1 U9511 ( .A1(n7195), .A2(n7194), .A3(n6653), .ZN(P3_U3201) );
  AOI21_X1 U9512 ( .B1(n6833), .B2(n11837), .A(n6835), .ZN(n11844) );
  XNOR2_X1 U9513 ( .A(n11653), .B(n8115), .ZN(n6833) );
  OR2_X2 U9514 ( .A1(n15496), .A2(n6645), .ZN(n7081) );
  OAI21_X1 U9515 ( .B1(n15517), .B2(n7079), .A(n7078), .ZN(n10209) );
  NOR2_X1 U9516 ( .A1(n14884), .A2(n14885), .ZN(n14883) );
  NOR2_X1 U9517 ( .A1(n10326), .A2(n10327), .ZN(n10329) );
  NOR2_X1 U9518 ( .A1(n12606), .A2(n12611), .ZN(n12627) );
  NOR2_X1 U9519 ( .A1(n10770), .A2(n10769), .ZN(n10933) );
  NAND2_X1 U9520 ( .A1(n11835), .A2(n6836), .ZN(n6835) );
  NAND2_X1 U9521 ( .A1(n6839), .A2(n11799), .ZN(n11801) );
  NAND2_X1 U9522 ( .A1(n6598), .A2(n6847), .ZN(n6846) );
  NAND2_X1 U9523 ( .A1(n12161), .A2(n12162), .ZN(n12160) );
  INV_X1 U9524 ( .A(n12192), .ZN(n7017) );
  NAND2_X1 U9525 ( .A1(n12245), .A2(n7009), .ZN(n7003) );
  NAND2_X1 U9526 ( .A1(n7003), .A2(n7008), .ZN(n7006) );
  NAND2_X1 U9527 ( .A1(n8469), .A2(n8468), .ZN(n8329) );
  OAI22_X1 U9528 ( .A1(n7651), .A2(n12130), .B1(n12129), .B2(n12128), .ZN(
        n12142) );
  NOR2_X1 U9529 ( .A1(n12759), .A2(n7554), .ZN(n7553) );
  XNOR2_X2 U9530 ( .A(n12757), .B(n12584), .ZN(n12759) );
  XNOR2_X1 U9531 ( .A(n6853), .B(n13552), .ZN(n13564) );
  OR2_X1 U9532 ( .A1(n13551), .A2(n13550), .ZN(n6853) );
  XNOR2_X2 U9533 ( .A(n8467), .B(n8478), .ZN(n9984) );
  OAI21_X2 U9534 ( .B1(n13696), .B2(n7480), .A(n7477), .ZN(n13661) );
  NAND2_X1 U9535 ( .A1(n7460), .A2(n8485), .ZN(n10651) );
  NAND2_X1 U9536 ( .A1(n8473), .A2(n8472), .ZN(n10698) );
  NAND2_X1 U9537 ( .A1(n13585), .A2(n13584), .ZN(n13583) );
  XNOR2_X1 U9538 ( .A(n15093), .B(n6855), .ZN(n15077) );
  NAND2_X1 U9539 ( .A1(n12725), .A2(n12726), .ZN(n12724) );
  NAND2_X1 U9540 ( .A1(n8002), .A2(n8000), .ZN(n7702) );
  NAND2_X1 U9541 ( .A1(n8037), .A2(n8036), .ZN(n7213) );
  OAI21_X1 U9542 ( .B1(n11832), .B2(n11838), .A(n6857), .ZN(n11835) );
  NAND2_X1 U9543 ( .A1(n11832), .A2(n11833), .ZN(n6857) );
  XNOR2_X1 U9544 ( .A(n7705), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8048) );
  OAI21_X2 U9545 ( .B1(n8091), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7707), .ZN(
        n7745) );
  NAND2_X1 U9546 ( .A1(n12696), .A2(n11097), .ZN(n8176) );
  NAND2_X2 U9547 ( .A1(n12707), .A2(n12708), .ZN(n12706) );
  NAND2_X1 U9548 ( .A1(n7108), .A2(n7107), .ZN(n12834) );
  INV_X1 U9549 ( .A(n11093), .ZN(n7889) );
  NAND2_X2 U9550 ( .A1(n9714), .A2(n9423), .ZN(n10257) );
  NAND2_X1 U9551 ( .A1(n6863), .A2(n6861), .ZN(n6860) );
  NAND2_X1 U9552 ( .A1(n10280), .A2(n12254), .ZN(n6863) );
  OAI21_X1 U9553 ( .B1(n14417), .B2(n6873), .A(n6870), .ZN(n14402) );
  NAND2_X1 U9554 ( .A1(n14417), .A2(n6870), .ZN(n6869) );
  NAND2_X1 U9555 ( .A1(n7416), .A2(n6885), .ZN(n11182) );
  NAND2_X1 U9556 ( .A1(n6707), .A2(n6890), .ZN(n6885) );
  INV_X1 U9557 ( .A(n10797), .ZN(n6898) );
  OAI211_X1 U9558 ( .C1(n6914), .C2(n14615), .A(n6913), .B(n6911), .ZN(
        P1_U3525) );
  NOR2_X2 U9559 ( .A1(n14799), .A2(n14800), .ZN(n14804) );
  OAI21_X1 U9560 ( .B1(n14757), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6693), .ZN(
        n6919) );
  INV_X1 U9561 ( .A(n6928), .ZN(n14864) );
  INV_X1 U9562 ( .A(n15018), .ZN(n6935) );
  MUX2_X1 U9563 ( .A(n7789), .B(P3_REG2_REG_4__SCAN_IN), .S(n15504), .Z(n15494) );
  MUX2_X1 U9564 ( .A(n15620), .B(P3_REG1_REG_4__SCAN_IN), .S(n15504), .Z(
        n15497) );
  OR2_X2 U9565 ( .A1(n11056), .A2(n11055), .ZN(n12618) );
  NAND2_X1 U9566 ( .A1(n8552), .A2(n6948), .ZN(n6945) );
  NAND2_X1 U9567 ( .A1(n8379), .A2(n6951), .ZN(n6954) );
  INV_X4 U9568 ( .A(n9681), .ZN(n9680) );
  MUX2_X1 U9569 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9681), .Z(n8342) );
  NAND2_X1 U9570 ( .A1(n8768), .A2(n6957), .ZN(n8390) );
  INV_X1 U9571 ( .A(n7493), .ZN(n7492) );
  NAND2_X1 U9572 ( .A1(n6958), .A2(n8922), .ZN(P2_U3496) );
  NOR2_X1 U9573 ( .A1(n13657), .A2(n6960), .ZN(n7287) );
  INV_X1 U9574 ( .A(n9652), .ZN(n6964) );
  INV_X1 U9575 ( .A(n6966), .ZN(n9651) );
  NAND2_X1 U9576 ( .A1(n11845), .A2(n6971), .ZN(n6970) );
  NAND2_X1 U9577 ( .A1(n11507), .A2(n11505), .ZN(n6984) );
  NAND2_X1 U9578 ( .A1(n6979), .A2(n6977), .ZN(n12457) );
  NAND2_X1 U9579 ( .A1(n11507), .A2(n6980), .ZN(n6979) );
  NAND2_X1 U9580 ( .A1(n11080), .A2(n6987), .ZN(n6986) );
  INV_X1 U9581 ( .A(n6988), .ZN(n11079) );
  NAND2_X1 U9582 ( .A1(n7666), .A2(n7665), .ZN(n8023) );
  NAND2_X1 U9583 ( .A1(n7666), .A2(n6999), .ZN(n8114) );
  NAND2_X1 U9584 ( .A1(n12076), .A2(n7000), .ZN(n7445) );
  NAND2_X1 U9585 ( .A1(n7001), .A2(n14553), .ZN(n7000) );
  NAND2_X1 U9586 ( .A1(n7002), .A2(n12064), .ZN(n7001) );
  NAND2_X1 U9587 ( .A1(n12061), .A2(n14566), .ZN(n7002) );
  NAND2_X1 U9588 ( .A1(n12233), .A2(n12232), .ZN(n7004) );
  NAND2_X1 U9589 ( .A1(n7007), .A2(n7010), .ZN(n7005) );
  NOR2_X1 U9590 ( .A1(n12289), .A2(n7006), .ZN(n12294) );
  NAND2_X1 U9591 ( .A1(n12231), .A2(n12230), .ZN(n7007) );
  NAND2_X1 U9592 ( .A1(n12192), .A2(n7018), .ZN(n7015) );
  OAI22_X1 U9593 ( .A1(n12142), .A2(n7021), .B1(n12143), .B2(n7022), .ZN(
        n12161) );
  NAND2_X1 U9594 ( .A1(n7027), .A2(n7025), .ZN(n12128) );
  NAND3_X1 U9595 ( .A1(n12110), .A2(n6668), .A3(n7028), .ZN(n7027) );
  INV_X1 U9596 ( .A(n12114), .ZN(n7029) );
  NAND3_X1 U9597 ( .A1(n11958), .A2(n11957), .A3(n7030), .ZN(n7031) );
  NAND3_X1 U9598 ( .A1(n7031), .A2(n6633), .A3(n11967), .ZN(n11966) );
  NAND2_X2 U9599 ( .A1(n8437), .A2(n9680), .ZN(n8802) );
  XNOR2_X2 U9600 ( .A(n8415), .B(n8414), .ZN(n9855) );
  INV_X1 U9601 ( .A(n7040), .ZN(n13841) );
  NAND2_X1 U9602 ( .A1(n13652), .A2(n7042), .ZN(n7043) );
  INV_X1 U9603 ( .A(n7043), .ZN(n13621) );
  NAND2_X1 U9604 ( .A1(n8248), .A2(n7044), .ZN(n8410) );
  NOR3_X2 U9605 ( .A1(n6588), .A2(n8258), .A3(n7047), .ZN(n8262) );
  INV_X1 U9606 ( .A(n7052), .ZN(n13978) );
  OR2_X2 U9607 ( .A1(n11063), .A2(n11062), .ZN(n12603) );
  OR2_X2 U9608 ( .A1(n12627), .A2(n7057), .ZN(n7056) );
  NAND2_X1 U9609 ( .A1(n7075), .A2(n7065), .ZN(n7066) );
  INV_X1 U9610 ( .A(n12632), .ZN(n7075) );
  XNOR2_X2 U9611 ( .A(n7081), .B(n15512), .ZN(n15517) );
  NAND3_X1 U9612 ( .A1(n7083), .A2(n7084), .A3(n7082), .ZN(n15476) );
  NAND3_X1 U9613 ( .A1(n10133), .A2(n9633), .A3(n9603), .ZN(n7082) );
  NAND2_X1 U9614 ( .A1(n7085), .A2(n15485), .ZN(n7084) );
  NAND2_X1 U9615 ( .A1(n7087), .A2(n7086), .ZN(n10135) );
  OR2_X2 U9616 ( .A1(n10933), .A2(n7089), .ZN(n7088) );
  NAND2_X1 U9617 ( .A1(n7092), .A2(n10912), .ZN(n11197) );
  INV_X1 U9618 ( .A(n7097), .ZN(n11245) );
  NOR2_X2 U9619 ( .A1(n6627), .A2(n12250), .ZN(n14477) );
  NOR2_X2 U9620 ( .A1(n14537), .A2(n14657), .ZN(n14529) );
  AND2_X1 U9621 ( .A1(n14436), .A2(n7098), .ZN(n14409) );
  NAND2_X1 U9622 ( .A1(n14436), .A2(n7099), .ZN(n14388) );
  NAND2_X1 U9623 ( .A1(n14436), .A2(n14623), .ZN(n14426) );
  NAND2_X1 U9624 ( .A1(n12867), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U9625 ( .A1(n12820), .A2(n7115), .ZN(n7112) );
  NAND2_X1 U9626 ( .A1(n7112), .A2(n7113), .ZN(n12795) );
  NAND2_X1 U9627 ( .A1(n12793), .A2(n7118), .ZN(n8066) );
  OAI21_X1 U9628 ( .B1(n6787), .B2(n8077), .A(n11679), .ZN(n12758) );
  INV_X1 U9629 ( .A(n12302), .ZN(n7131) );
  NAND2_X1 U9630 ( .A1(n13279), .A2(n6590), .ZN(n7132) );
  NAND2_X1 U9631 ( .A1(n8113), .A2(n9289), .ZN(n8930) );
  AND2_X2 U9632 ( .A1(n7955), .A2(n6601), .ZN(n7714) );
  NAND2_X1 U9633 ( .A1(n7141), .A2(n7140), .ZN(n9517) );
  NAND2_X1 U9634 ( .A1(n14385), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U9635 ( .A1(n12066), .A2(n14177), .ZN(n7169) );
  NAND2_X1 U9636 ( .A1(n9477), .A2(n9680), .ZN(n11168) );
  OAI21_X1 U9637 ( .B1(n7170), .B2(n9709), .A(n7165), .ZN(n7168) );
  NAND2_X1 U9638 ( .A1(n11922), .A2(n7166), .ZN(n7165) );
  NAND2_X2 U9639 ( .A1(n7167), .A2(n7169), .ZN(n10061) );
  INV_X1 U9640 ( .A(n9619), .ZN(n7172) );
  NAND2_X1 U9641 ( .A1(n7172), .A2(n9603), .ZN(n7173) );
  INV_X1 U9642 ( .A(n7175), .ZN(n7174) );
  NAND2_X1 U9643 ( .A1(n9619), .A2(n15485), .ZN(n7175) );
  INV_X1 U9644 ( .A(n12620), .ZN(n7184) );
  NAND3_X1 U9645 ( .A1(n7182), .A2(n7183), .A3(n7180), .ZN(n15527) );
  NAND3_X1 U9646 ( .A1(n7182), .A2(n7181), .A3(n7180), .ZN(n7185) );
  INV_X1 U9647 ( .A(n7185), .ZN(n15526) );
  NOR2_X1 U9648 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7187) );
  MUX2_X1 U9649 ( .A(n10357), .B(n15531), .S(P3_IR_REG_0__SCAN_IN), .Z(n10358)
         );
  INV_X1 U9650 ( .A(n9622), .ZN(n7193) );
  NAND2_X1 U9651 ( .A1(n7977), .A2(n7975), .ZN(n7699) );
  NAND2_X1 U9652 ( .A1(n7954), .A2(n7953), .ZN(n7198) );
  NAND2_X1 U9653 ( .A1(n7205), .A2(n7209), .ZN(n7692) );
  NAND2_X1 U9654 ( .A1(n7689), .A2(n7206), .ZN(n7205) );
  NAND2_X1 U9655 ( .A1(n7216), .A2(n7214), .ZN(n7682) );
  INV_X1 U9656 ( .A(n7223), .ZN(n8079) );
  INV_X1 U9657 ( .A(n6568), .ZN(n10153) );
  OAI22_X1 U9658 ( .A1(n15561), .A2(n6568), .B1(n10737), .B2(n15563), .ZN(
        n10740) );
  NAND3_X1 U9659 ( .A1(n7229), .A2(n12485), .A3(n9368), .ZN(n12543) );
  NAND2_X1 U9660 ( .A1(n7232), .A2(n7230), .ZN(n12481) );
  NAND2_X1 U9661 ( .A1(n9378), .A2(n12498), .ZN(n7238) );
  NAND2_X1 U9662 ( .A1(n7233), .A2(n7234), .ZN(n12554) );
  NAND3_X1 U9663 ( .A1(n9378), .A2(n12498), .A3(n9382), .ZN(n7233) );
  NAND2_X1 U9664 ( .A1(n10792), .A2(n7241), .ZN(n7239) );
  NAND2_X1 U9665 ( .A1(n12563), .A2(n7250), .ZN(n7249) );
  NAND2_X2 U9666 ( .A1(n7249), .A2(n7248), .ZN(n11845) );
  NAND2_X1 U9667 ( .A1(n7714), .A2(n6704), .ZN(n7256) );
  INV_X1 U9668 ( .A(n7256), .ZN(n7732) );
  OAI22_X1 U9669 ( .A1(n9325), .A2(n9324), .B1(n9323), .B2(n9328), .ZN(n15460)
         );
  INV_X4 U9670 ( .A(n12440), .ZN(n10292) );
  NAND2_X1 U9671 ( .A1(n9346), .A2(n9345), .ZN(n12459) );
  NAND4_X1 U9672 ( .A1(n7257), .A2(n15369), .A3(n6573), .A4(n10718), .ZN(n9240) );
  NAND2_X1 U9673 ( .A1(n7261), .A2(n7259), .ZN(n13869) );
  OR2_X1 U9674 ( .A1(n7264), .A2(n8887), .ZN(n7260) );
  NAND2_X1 U9675 ( .A1(n10676), .A2(n7262), .ZN(n7261) );
  INV_X1 U9676 ( .A(n7264), .ZN(n7262) );
  NAND2_X1 U9677 ( .A1(n13848), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U9678 ( .A1(n13618), .A2(n6597), .ZN(n7272) );
  OAI21_X1 U9679 ( .B1(n13760), .B2(n7278), .A(n7276), .ZN(n13724) );
  OAI21_X1 U9680 ( .B1(n13760), .B2(n8899), .A(n8900), .ZN(n13746) );
  NAND2_X1 U9681 ( .A1(n7281), .A2(n7283), .ZN(n8913) );
  OAI21_X1 U9682 ( .B1(n11382), .B2(n7292), .A(n7290), .ZN(n13767) );
  NAND4_X1 U9683 ( .A1(n7301), .A2(n7302), .A3(n8235), .A4(n7308), .ZN(n7304)
         );
  NOR2_X2 U9684 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7302) );
  NOR2_X2 U9685 ( .A1(n7304), .A2(n7303), .ZN(n8572) );
  OAI211_X1 U9686 ( .C1(n13399), .C2(n7314), .A(n7310), .B(n7312), .ZN(n13348)
         );
  NAND2_X1 U9687 ( .A1(n13360), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U9688 ( .A1(n13360), .A2(n7320), .ZN(n7317) );
  AOI21_X1 U9689 ( .B1(n7315), .B2(n7313), .A(n6613), .ZN(n7312) );
  NAND2_X1 U9690 ( .A1(n7317), .A2(n7318), .ZN(n13482) );
  NOR2_X1 U9691 ( .A1(n8677), .A2(n7331), .ZN(n7323) );
  NOR2_X1 U9692 ( .A1(n7323), .A2(n7326), .ZN(n7325) );
  OAI21_X1 U9693 ( .B1(n11491), .B2(n7347), .A(n7344), .ZN(n13292) );
  OAI211_X1 U9694 ( .C1(n8334), .C2(n7366), .A(n7363), .B(n8337), .ZN(n8340)
         );
  NAND2_X1 U9695 ( .A1(n8333), .A2(n7364), .ZN(n7363) );
  AND2_X1 U9696 ( .A1(n8336), .A2(n8332), .ZN(n7364) );
  NAND2_X1 U9697 ( .A1(n7365), .A2(n8336), .ZN(n8501) );
  NAND2_X1 U9698 ( .A1(n8496), .A2(n8334), .ZN(n7365) );
  NAND2_X1 U9699 ( .A1(n7367), .A2(n7368), .ZN(n8552) );
  NAND2_X1 U9700 ( .A1(n8520), .A2(n7370), .ZN(n7367) );
  AOI21_X1 U9701 ( .B1(n8586), .B2(n8354), .A(n7374), .ZN(n7372) );
  NAND2_X1 U9702 ( .A1(n8585), .A2(n8354), .ZN(n7373) );
  NAND2_X1 U9703 ( .A1(n7387), .A2(n8404), .ZN(n8855) );
  INV_X1 U9704 ( .A(n7390), .ZN(n7389) );
  NAND2_X1 U9705 ( .A1(n8395), .A2(n8393), .ZN(n8799) );
  NOR2_X2 U9706 ( .A1(n14783), .A2(n14784), .ZN(n14787) );
  INV_X1 U9707 ( .A(n14806), .ZN(n7396) );
  OR2_X1 U9708 ( .A1(n15024), .A2(n7401), .ZN(n7398) );
  OAI21_X1 U9709 ( .B1(n7403), .B2(n15029), .A(n7398), .ZN(n15027) );
  OR2_X1 U9710 ( .A1(n15029), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U9711 ( .A1(n7405), .A2(n14847), .ZN(n7404) );
  NAND2_X1 U9712 ( .A1(n7407), .A2(n14794), .ZN(n7405) );
  NAND2_X1 U9713 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  NAND3_X1 U9714 ( .A1(n7409), .A2(n7408), .A3(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7406) );
  NAND2_X1 U9715 ( .A1(n9432), .A2(n7431), .ZN(n7430) );
  NOR2_X2 U9716 ( .A1(n7430), .A2(n10257), .ZN(n9448) );
  OAI21_X1 U9717 ( .B1(n15077), .B2(n15079), .A(n11946), .ZN(n10280) );
  NAND3_X1 U9718 ( .A1(n11982), .A2(n11981), .A3(n6711), .ZN(n7433) );
  INV_X1 U9719 ( .A(n11984), .ZN(n7434) );
  NAND3_X1 U9720 ( .A1(n11971), .A2(n11970), .A3(n6712), .ZN(n7436) );
  INV_X1 U9721 ( .A(n11973), .ZN(n7437) );
  NAND2_X1 U9722 ( .A1(n7438), .A2(n7440), .ZN(n12006) );
  NAND3_X1 U9723 ( .A1(n11998), .A2(n7439), .A3(n11997), .ZN(n7438) );
  NAND3_X1 U9724 ( .A1(n7459), .A2(n7454), .A3(P1_IR_REG_19__SCAN_IN), .ZN(
        n7453) );
  INV_X2 U9725 ( .A(n10257), .ZN(n9541) );
  NAND2_X1 U9726 ( .A1(n10651), .A2(n10650), .ZN(n8500) );
  INV_X1 U9727 ( .A(n11374), .ZN(n7464) );
  OAI211_X1 U9728 ( .C1(n7492), .C2(n15455), .A(n7489), .B(n6727), .ZN(
        P2_U3528) );
  OAI21_X1 U9729 ( .B1(n12434), .B2(n15407), .A(n8921), .ZN(n7493) );
  NAND2_X1 U9730 ( .A1(n7495), .A2(n7494), .ZN(n8717) );
  AND2_X1 U9731 ( .A1(n6641), .A2(n7496), .ZN(n7494) );
  NAND2_X1 U9732 ( .A1(n8269), .A2(n7506), .ZN(n8408) );
  NOR2_X1 U9733 ( .A1(n7518), .A2(n7517), .ZN(n7516) );
  XNOR2_X1 U9734 ( .A(n11388), .B(n11386), .ZN(n11390) );
  NAND2_X1 U9735 ( .A1(n7519), .A2(n7520), .ZN(n14090) );
  NAND2_X1 U9736 ( .A1(n14117), .A2(n7521), .ZN(n7519) );
  NAND2_X1 U9737 ( .A1(n14067), .A2(n7528), .ZN(n7525) );
  NAND2_X1 U9738 ( .A1(n14067), .A2(n14068), .ZN(n7527) );
  NAND2_X1 U9739 ( .A1(n6583), .A2(n7536), .ZN(n7531) );
  INV_X1 U9740 ( .A(n9439), .ZN(n12425) );
  INV_X1 U9741 ( .A(n9445), .ZN(n7540) );
  NAND2_X1 U9742 ( .A1(n9426), .A2(n6696), .ZN(n7547) );
  NAND2_X1 U9743 ( .A1(n12846), .A2(n7549), .ZN(n7548) );
  NAND2_X1 U9744 ( .A1(n8121), .A2(n10293), .ZN(n15556) );
  NAND2_X1 U9745 ( .A1(n15464), .A2(n10734), .ZN(n11686) );
  NAND2_X1 U9746 ( .A1(n8149), .A2(n7557), .ZN(n7556) );
  NAND2_X1 U9747 ( .A1(n8131), .A2(n7562), .ZN(n7564) );
  OAI211_X1 U9748 ( .C1(n7576), .C2(n8932), .A(n7574), .B(n7573), .ZN(n9307)
         );
  NAND3_X1 U9749 ( .A1(n8932), .A2(n7572), .A3(n7580), .ZN(n7573) );
  OR2_X1 U9750 ( .A1(n11677), .A2(n7578), .ZN(n7576) );
  NAND2_X1 U9751 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NOR2_X2 U9752 ( .A1(n12441), .A2(n7581), .ZN(n7580) );
  INV_X1 U9753 ( .A(n8931), .ZN(n7581) );
  OAI21_X1 U9754 ( .B1(n8143), .B2(n7584), .A(n7582), .ZN(n8146) );
  NAND3_X1 U9755 ( .A1(n7589), .A2(n7588), .A3(n7595), .ZN(n7587) );
  NAND2_X1 U9756 ( .A1(n9056), .A2(n9055), .ZN(n7588) );
  NAND2_X1 U9757 ( .A1(n9052), .A2(n9051), .ZN(n7589) );
  NAND3_X1 U9758 ( .A1(n7592), .A2(n7591), .A3(n7596), .ZN(n7590) );
  NAND2_X1 U9759 ( .A1(n9056), .A2(n7593), .ZN(n7591) );
  NAND2_X1 U9760 ( .A1(n9052), .A2(n7594), .ZN(n7592) );
  AND2_X1 U9761 ( .A1(n9061), .A2(n9051), .ZN(n7594) );
  INV_X1 U9762 ( .A(n9061), .ZN(n7595) );
  INV_X1 U9763 ( .A(n9060), .ZN(n7596) );
  AOI21_X1 U9764 ( .B1(n9013), .B2(n6595), .A(n7598), .ZN(n7597) );
  INV_X1 U9765 ( .A(n7597), .ZN(n9018) );
  AND2_X1 U9766 ( .A1(n9120), .A2(n7613), .ZN(n7612) );
  NAND3_X1 U9767 ( .A1(n9069), .A2(n9070), .A3(n6721), .ZN(n7618) );
  NAND2_X1 U9768 ( .A1(n8262), .A2(n7628), .ZN(n7632) );
  NAND3_X1 U9769 ( .A1(n9089), .A2(n7653), .A3(n6710), .ZN(n7633) );
  NAND2_X1 U9770 ( .A1(n7633), .A2(n7634), .ZN(n9099) );
  AOI21_X1 U9771 ( .B1(n9099), .B2(n9098), .A(n9096), .ZN(n9097) );
  AND2_X1 U9772 ( .A1(n12497), .A2(n12500), .ZN(n9378) );
  NAND2_X1 U9773 ( .A1(n9377), .A2(n9376), .ZN(n12497) );
  NAND2_X1 U9774 ( .A1(n10447), .A2(n9478), .ZN(n9480) );
  AND2_X1 U9775 ( .A1(n10249), .A2(n9237), .ZN(n15369) );
  CLKBUF_X1 U9776 ( .A(n11214), .Z(n11888) );
  INV_X1 U9777 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7722) );
  INV_X1 U9778 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7721) );
  INV_X1 U9779 ( .A(n12209), .ZN(n12210) );
  NAND2_X1 U9780 ( .A1(n11937), .A2(n11936), .ZN(n11943) );
  NAND2_X1 U9781 ( .A1(n9375), .A2(n6643), .ZN(n12498) );
  NAND2_X2 U9782 ( .A1(n12126), .A2(n12125), .ZN(n12250) );
  NAND2_X1 U9783 ( .A1(n14402), .A2(n14401), .ZN(n14408) );
  NAND2_X1 U9784 ( .A1(n8176), .A2(n7643), .ZN(n12697) );
  INV_X1 U9785 ( .A(n8957), .ZN(n13565) );
  XNOR2_X1 U9786 ( .A(n13292), .B(n13290), .ZN(n13289) );
  CLKBUF_X1 U9787 ( .A(n11491), .Z(n11299) );
  MUX2_X1 U9788 ( .A(n14630), .B(n14452), .S(n12241), .Z(n12159) );
  INV_X1 U9789 ( .A(n12143), .ZN(n12144) );
  OAI211_X1 U9790 ( .C1(n9187), .C2(n9186), .A(n9185), .B(n9184), .ZN(n14001)
         );
  NAND2_X1 U9791 ( .A1(n8957), .A2(n11319), .ZN(n8963) );
  NAND2_X1 U9792 ( .A1(n7720), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U9793 ( .A1(n9370), .A2(n9369), .ZN(n12527) );
  NAND2_X1 U9794 ( .A1(n7889), .A2(n11725), .ZN(n7890) );
  NAND4_X4 U9795 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n14171)
         );
  OR2_X2 U9796 ( .A1(n12202), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9498) );
  AND2_X1 U9797 ( .A1(n10056), .A2(n9584), .ZN(n10052) );
  NAND2_X1 U9798 ( .A1(n8462), .A2(n8461), .ZN(n10163) );
  NAND2_X1 U9799 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  XNOR2_X1 U9800 ( .A(n12600), .B(n10413), .ZN(n11702) );
  AOI21_X2 U9801 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12648), .A(n12647), .ZN(
        n12650) );
  NOR2_X1 U9802 ( .A1(n11620), .A2(n11828), .ZN(n11652) );
  INV_X1 U9803 ( .A(n9019), .ZN(n9020) );
  NAND2_X1 U9804 ( .A1(n11938), .A2(n6575), .ZN(n9479) );
  AND2_X1 U9805 ( .A1(n10076), .A2(n12327), .ZN(n10034) );
  INV_X1 U9806 ( .A(n9053), .ZN(n9056) );
  AND2_X1 U9807 ( .A1(n9855), .A2(n10173), .ZN(n13851) );
  INV_X1 U9808 ( .A(n9106), .ZN(n9109) );
  AOI21_X1 U9809 ( .B1(n12692), .B2(n15600), .A(n8942), .ZN(n8954) );
  NAND2_X2 U9810 ( .A1(n13880), .A2(n10646), .ZN(n13883) );
  NAND2_X1 U9811 ( .A1(n13880), .A2(n10185), .ZN(n15223) );
  AND3_X2 U9812 ( .A1(n10645), .A2(n10183), .A3(n15366), .ZN(n15444) );
  NAND2_X1 U9813 ( .A1(n9541), .A2(n9537), .ZN(n7637) );
  AND2_X2 U9814 ( .A1(n10313), .A2(n8232), .ZN(n15631) );
  NAND2_X1 U9815 ( .A1(n6845), .A2(n11646), .ZN(n7640) );
  OR2_X1 U9816 ( .A1(n8388), .A2(n11090), .ZN(n7644) );
  OR2_X1 U9817 ( .A1(n13215), .A2(n13211), .ZN(n7645) );
  OR2_X1 U9818 ( .A1(n11557), .A2(n11517), .ZN(n7646) );
  INV_X1 U9819 ( .A(n12485), .ZN(n12585) );
  INV_X1 U9820 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13176) );
  INV_X1 U9821 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10786) );
  INV_X1 U9822 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7693) );
  OR2_X1 U9823 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9632), .ZN(n7647) );
  INV_X1 U9824 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15525) );
  INV_X1 U9825 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10084) );
  INV_X1 U9826 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10360) );
  AND2_X1 U9827 ( .A1(n9234), .A2(n9233), .ZN(n7648) );
  INV_X1 U9828 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10835) );
  INV_X1 U9829 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7883) );
  INV_X1 U9830 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10004) );
  INV_X1 U9831 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10306) );
  CLKBUF_X3 U9832 ( .A(n13331), .Z(n13318) );
  OR2_X1 U9833 ( .A1(n12781), .A2(n12546), .ZN(n7649) );
  INV_X1 U9834 ( .A(n11645), .ZN(n12683) );
  INV_X1 U9835 ( .A(n9254), .ZN(n8864) );
  INV_X1 U9836 ( .A(n13845), .ZN(n8918) );
  INV_X1 U9837 ( .A(n13729), .ZN(n13741) );
  AND2_X2 U9838 ( .A1(n8952), .A2(n11839), .ZN(n15613) );
  AND2_X1 U9839 ( .A1(n12284), .A2(n12286), .ZN(n7655) );
  NAND2_X1 U9840 ( .A1(n11949), .A2(n12178), .ZN(n11950) );
  NAND2_X1 U9841 ( .A1(n8975), .A2(n8974), .ZN(n8978) );
  NAND2_X1 U9842 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  INV_X1 U9843 ( .A(n9010), .ZN(n9011) );
  OAI21_X1 U9844 ( .B1(n11287), .B2(n9264), .A(n9035), .ZN(n9036) );
  INV_X1 U9845 ( .A(n9036), .ZN(n9039) );
  AND2_X1 U9846 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  NAND2_X1 U9847 ( .A1(n9046), .A2(n7650), .ZN(n9053) );
  INV_X1 U9848 ( .A(n9054), .ZN(n9055) );
  INV_X1 U9849 ( .A(n12127), .ZN(n12130) );
  OAI21_X1 U9850 ( .B1(n13374), .B2(n9264), .A(n9092), .ZN(n9093) );
  INV_X1 U9851 ( .A(n12162), .ZN(n12163) );
  INV_X1 U9852 ( .A(n9107), .ZN(n9108) );
  INV_X1 U9853 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7660) );
  INV_X1 U9854 ( .A(SI_17_), .ZN(n8370) );
  INV_X1 U9855 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7670) );
  INV_X1 U9856 ( .A(n9220), .ZN(n9211) );
  INV_X1 U9857 ( .A(n8783), .ZN(n8388) );
  INV_X1 U9858 ( .A(n6800), .ZN(n8123) );
  INV_X1 U9859 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9860 ( .A1(n9212), .A2(n9211), .ZN(n9213) );
  INV_X1 U9861 ( .A(n13951), .ZN(n8919) );
  INV_X1 U9862 ( .A(n10279), .ZN(n12254) );
  INV_X1 U9863 ( .A(n8621), .ZN(n8360) );
  INV_X1 U9864 ( .A(n12528), .ZN(n9376) );
  INV_X1 U9865 ( .A(n12814), .ZN(n8149) );
  INV_X1 U9866 ( .A(n11658), .ZN(n8127) );
  OR2_X1 U9867 ( .A1(n12673), .A2(n8221), .ZN(n8946) );
  INV_X1 U9868 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8178) );
  INV_X1 U9869 ( .A(n8710), .ZN(n8301) );
  INV_X1 U9870 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U9871 ( .A1(n13729), .A2(n8919), .ZN(n13730) );
  INV_X1 U9872 ( .A(SI_11_), .ZN(n8350) );
  INV_X1 U9873 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7964) );
  INV_X1 U9874 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8043) );
  INV_X1 U9875 ( .A(n9336), .ZN(n9337) );
  OR2_X1 U9876 ( .A1(n8946), .A2(n11836), .ZN(n9391) );
  OAI22_X1 U9877 ( .A1(n9304), .A2(n15561), .B1(n14935), .B2(n11647), .ZN(
        n9305) );
  NOR2_X1 U9878 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8095), .ZN(n8094) );
  NOR2_X1 U9879 ( .A1(n8084), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8083) );
  OR2_X1 U9880 ( .A1(n7908), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7925) );
  INV_X1 U9881 ( .A(n15512), .ZN(n9636) );
  NAND2_X1 U9882 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12438), .ZN(n11627) );
  NAND2_X1 U9883 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10306), .ZN(n7700) );
  NOR2_X1 U9884 ( .A1(n9216), .A2(n9215), .ZN(n9217) );
  OR2_X1 U9885 ( .A1(n8829), .A2(n8304), .ZN(n8844) );
  INV_X1 U9886 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U9887 ( .A1(n8299), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8696) );
  INV_X1 U9888 ( .A(n13673), .ZN(n8920) );
  OR2_X1 U9889 ( .A1(n8728), .A2(n8727), .ZN(n8744) );
  INV_X1 U9890 ( .A(n11319), .ZN(n8874) );
  OR2_X1 U9891 ( .A1(n8596), .A2(n8595), .ZN(n8611) );
  INV_X1 U9892 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10959) );
  INV_X1 U9893 ( .A(n11139), .ZN(n11136) );
  NAND2_X1 U9894 ( .A1(n11597), .A2(n11598), .ZN(n11599) );
  AND2_X1 U9895 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  INV_X1 U9896 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11537) );
  OR2_X1 U9897 ( .A1(n11923), .A2(n15134), .ZN(n10044) );
  INV_X1 U9898 ( .A(n12261), .ZN(n10615) );
  INV_X1 U9899 ( .A(n10447), .ZN(n12255) );
  INV_X1 U9900 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7891) );
  AND2_X1 U9901 ( .A1(n7875), .A2(n7735), .ZN(n7892) );
  INV_X1 U9902 ( .A(n12830), .ZN(n12517) );
  INV_X1 U9903 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12570) );
  INV_X1 U9904 ( .A(n8082), .ZN(n8166) );
  AND2_X1 U9905 ( .A1(n8198), .A2(n8194), .ZN(n8212) );
  INV_X1 U9906 ( .A(n11680), .ZN(n12766) );
  INV_X1 U9907 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13162) );
  AND2_X1 U9908 ( .A1(n11746), .A2(n11749), .ZN(n11410) );
  INV_X1 U9909 ( .A(n15560), .ZN(n12861) );
  INV_X1 U9910 ( .A(n11731), .ZN(n11664) );
  NOR2_X2 U9911 ( .A1(n11837), .A2(n8164), .ZN(n15560) );
  INV_X1 U9912 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7864) );
  INV_X1 U9913 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13365) );
  INV_X1 U9914 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U9915 ( .A1(n8303), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8829) );
  AND2_X1 U9916 ( .A1(n12430), .A2(n8307), .ZN(n13593) );
  OR2_X1 U9917 ( .A1(n8744), .A2(n8743), .ZN(n8756) );
  INV_X1 U9918 ( .A(n13501), .ZN(n13714) );
  INV_X1 U9919 ( .A(n9246), .ZN(n13815) );
  INV_X1 U9920 ( .A(n9243), .ZN(n13855) );
  INV_X1 U9921 ( .A(n13851), .ZN(n13872) );
  AND2_X1 U9922 ( .A1(n10177), .A2(n10176), .ZN(n10178) );
  AND2_X1 U9923 ( .A1(n9164), .A2(n8865), .ZN(n13712) );
  NAND2_X1 U9924 ( .A1(n10885), .A2(n10887), .ZN(n10888) );
  NAND2_X1 U9925 ( .A1(n11133), .A2(n11132), .ZN(n11134) );
  INV_X1 U9926 ( .A(n11607), .ZN(n11608) );
  OR2_X1 U9927 ( .A1(n12335), .A2(n12334), .ZN(n12336) );
  NAND2_X2 U9928 ( .A1(n9554), .A2(n14187), .ZN(n9477) );
  INV_X1 U9929 ( .A(n14568), .ZN(n14132) );
  INV_X1 U9930 ( .A(n9495), .ZN(n9522) );
  AND2_X1 U9931 ( .A1(n12077), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12089) );
  INV_X1 U9932 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10513) );
  INV_X1 U9933 ( .A(n15070), .ZN(n15046) );
  AND2_X1 U9934 ( .A1(n10110), .A2(n10109), .ZN(n9586) );
  NAND2_X1 U9935 ( .A1(n14404), .A2(n14569), .ZN(n14405) );
  AND2_X1 U9936 ( .A1(n15134), .A2(n15133), .ZN(n12237) );
  AND2_X1 U9937 ( .A1(n9546), .A2(n12327), .ZN(n10362) );
  INV_X1 U9938 ( .A(n14451), .ZN(n14455) );
  INV_X1 U9939 ( .A(n14161), .ZN(n14981) );
  INV_X1 U9940 ( .A(n14569), .ZN(n14591) );
  INV_X1 U9941 ( .A(n12265), .ZN(n10819) );
  INV_X1 U9942 ( .A(n12259), .ZN(n10474) );
  NAND2_X1 U9943 ( .A1(n8824), .A2(n8401), .ZN(n8841) );
  AND2_X1 U9944 ( .A1(n8668), .A2(n8365), .ZN(n8652) );
  AND2_X1 U9945 ( .A1(n8619), .A2(n8357), .ZN(n8603) );
  NOR2_X1 U9946 ( .A1(n14742), .A2(n14741), .ZN(n14795) );
  OR2_X1 U9947 ( .A1(n12571), .A2(n15561), .ZN(n11083) );
  INV_X1 U9948 ( .A(n11083), .ZN(n15465) );
  INV_X1 U9949 ( .A(n13266), .ZN(n10151) );
  AND2_X1 U9950 ( .A1(n11839), .A2(n14950), .ZN(n10307) );
  OR2_X1 U9951 ( .A1(n8072), .A2(n8936), .ZN(n11643) );
  AND4_X1 U9952 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(n12485)
         );
  AND4_X1 U9953 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(n12509)
         );
  INV_X1 U9954 ( .A(n15531), .ZN(n14926) );
  AND2_X1 U9955 ( .A1(n8169), .A2(n8168), .ZN(n14939) );
  OR2_X1 U9956 ( .A1(n11097), .A2(n11037), .ZN(n15565) );
  NOR2_X1 U9957 ( .A1(n15631), .A2(n9314), .ZN(n9315) );
  NOR2_X1 U9958 ( .A1(n8220), .A2(n8219), .ZN(n10313) );
  AND2_X1 U9959 ( .A1(n14937), .A2(n14936), .ZN(n14949) );
  NOR2_X1 U9960 ( .A1(n9899), .A2(n13266), .ZN(n9908) );
  AND2_X1 U9961 ( .A1(n7938), .A2(n7937), .ZN(n11068) );
  INV_X1 U9962 ( .A(n13284), .ZN(n14834) );
  AOI21_X1 U9963 ( .B1(n13348), .B2(n13347), .A(n13480), .ZN(n13357) );
  INV_X1 U9964 ( .A(n15216), .ZN(n13476) );
  INV_X1 U9965 ( .A(n13480), .ZN(n13492) );
  AND3_X1 U9966 ( .A1(n8872), .A2(n8871), .A3(n8870), .ZN(n9166) );
  OR2_X1 U9967 ( .A1(n13645), .A2(n8613), .ZN(n8810) );
  OR2_X1 U9968 ( .A1(n9854), .A2(n9845), .ZN(n15265) );
  INV_X1 U9969 ( .A(n15263), .ZN(n15302) );
  INV_X1 U9970 ( .A(n13979), .ZN(n15323) );
  NAND2_X1 U9971 ( .A1(n10179), .A2(n10178), .ZN(n10255) );
  OR2_X1 U9972 ( .A1(n8963), .A2(n10718), .ZN(n15438) );
  INV_X1 U9973 ( .A(n15407), .ZN(n15379) );
  AND2_X1 U9974 ( .A1(n8288), .A2(n8287), .ZN(n15330) );
  AND2_X1 U9975 ( .A1(n9592), .A2(n9840), .ZN(n10176) );
  INV_X1 U9976 ( .A(n14998), .ZN(n14134) );
  AND2_X1 U9977 ( .A1(n10122), .A2(n10109), .ZN(n10058) );
  AND4_X1 U9978 ( .A1(n11918), .A2(n11917), .A3(n11916), .A4(n11915), .ZN(
        n14376) );
  AND2_X1 U9979 ( .A1(n9796), .A2(n9795), .ZN(n15070) );
  INV_X1 U9980 ( .A(n15053), .ZN(n15071) );
  NAND2_X1 U9981 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  AND2_X1 U9982 ( .A1(n12237), .A2(n11866), .ZN(n14570) );
  INV_X1 U9983 ( .A(n14601), .ZN(n14562) );
  OR2_X1 U9984 ( .A1(n15098), .A2(n10043), .ZN(n15088) );
  INV_X1 U9985 ( .A(n14543), .ZN(n15094) );
  INV_X1 U9986 ( .A(n15088), .ZN(n14558) );
  AND2_X1 U9987 ( .A1(n9570), .A2(n9569), .ZN(n10122) );
  NAND2_X1 U9988 ( .A1(n12238), .A2(n14445), .ZN(n15184) );
  NAND2_X1 U9989 ( .A1(n10911), .A2(n15184), .ZN(n15198) );
  NAND2_X1 U9990 ( .A1(n9568), .A2(n6818), .ZN(n9731) );
  AND2_X1 U9991 ( .A1(n9741), .A2(n9740), .ZN(n10801) );
  AND2_X1 U9992 ( .A1(n9643), .A2(n9642), .ZN(n15458) );
  INV_X1 U9993 ( .A(n9412), .ZN(n9413) );
  INV_X1 U9994 ( .A(n15469), .ZN(n12552) );
  NAND2_X1 U9995 ( .A1(n9395), .A2(n10307), .ZN(n12576) );
  INV_X1 U9996 ( .A(n12492), .ZN(n12581) );
  OR2_X1 U9997 ( .A1(n9594), .A2(n13266), .ZN(n12589) );
  MUX2_X1 U9998 ( .A(n9640), .B(n12589), .S(n7131), .Z(n15531) );
  OR2_X1 U9999 ( .A1(n9640), .A2(n9627), .ZN(n15547) );
  INV_X1 U10000 ( .A(n12872), .ZN(n12857) );
  INV_X1 U10001 ( .A(n15631), .ZN(n15628) );
  INV_X1 U10002 ( .A(n12701), .ZN(n13215) );
  INV_X1 U10003 ( .A(n8142), .ZN(n11557) );
  INV_X1 U10004 ( .A(n15613), .ZN(n15612) );
  AND2_X1 U10005 ( .A1(n8201), .A2(n8200), .ZN(n13265) );
  INV_X1 U10006 ( .A(SI_20_), .ZN(n10554) );
  INV_X1 U10007 ( .A(SI_16_), .ZN(n10001) );
  NAND2_X1 U10008 ( .A1(n10254), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15226) );
  NAND3_X1 U10009 ( .A1(n10184), .A2(n15428), .A3(n10174), .ZN(n13480) );
  INV_X1 U10010 ( .A(n15223), .ZN(n13447) );
  NAND2_X1 U10011 ( .A1(n8851), .A2(n8850), .ZN(n13499) );
  OR2_X1 U10012 ( .A1(n9842), .A2(P2_U3088), .ZN(n13507) );
  OR2_X1 U10013 ( .A1(n9861), .A2(P2_U3088), .ZN(n15297) );
  OR2_X1 U10014 ( .A1(n9854), .A2(n14014), .ZN(n15263) );
  NAND2_X1 U10015 ( .A1(n13883), .A2(n10648), .ZN(n14959) );
  OR2_X1 U10016 ( .A1(n15226), .A2(n10255), .ZN(n15455) );
  AND3_X1 U10017 ( .A1(n15411), .A2(n15410), .A3(n15409), .ZN(n15450) );
  INV_X1 U10018 ( .A(n15444), .ZN(n15442) );
  INV_X1 U10019 ( .A(n10718), .ZN(n10920) );
  INV_X1 U10020 ( .A(n12002), .ZN(n14852) );
  NAND2_X1 U10021 ( .A1(n10528), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14998) );
  NAND2_X1 U10022 ( .A1(n10058), .A2(n10048), .ZN(n14989) );
  INV_X1 U10023 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11429) );
  OR2_X1 U10024 ( .A1(n9782), .A2(n14333), .ZN(n15053) );
  INV_X1 U10025 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U10026 ( .A1(n9726), .A2(n9724), .ZN(n15075) );
  OR2_X1 U10027 ( .A1(n14393), .A2(n14445), .ZN(n14543) );
  INV_X1 U10028 ( .A(n14547), .ZN(n15086) );
  OR2_X1 U10029 ( .A1(n15098), .A2(n12239), .ZN(n10918) );
  INV_X2 U10030 ( .A(n14547), .ZN(n15098) );
  INV_X1 U10031 ( .A(n15213), .ZN(n15210) );
  INV_X1 U10032 ( .A(n15200), .ZN(n15199) );
  AND3_X2 U10033 ( .A1(n10124), .A2(n10123), .A3(n10110), .ZN(n15200) );
  AND2_X2 U10034 ( .A1(n10052), .A2(n9731), .ZN(n15129) );
  INV_X1 U10035 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11868) );
  INV_X1 U10036 ( .A(n10042), .ZN(n15133) );
  INV_X1 U10037 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9758) );
  INV_X2 U10038 ( .A(n12589), .ZN(P3_U3897) );
  INV_X1 U10039 ( .A(n13507), .ZN(P2_U3947) );
  OR4_X1 U10040 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(P1_U3288) );
  INV_X1 U10041 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8233) );
  INV_X2 U10042 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10043 ( .A1(n8114), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U10044 ( .A1(n8023), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7668) );
  MUX2_X1 U10045 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7668), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n7669) );
  NAND2_X1 U10046 ( .A1(n10555), .A2(n8115), .ZN(n11833) );
  INV_X1 U10047 ( .A(n7714), .ZN(n7673) );
  AOI22_X1 U10048 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10919), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7212), .ZN(n8036) );
  AOI22_X1 U10049 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n13072), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6851), .ZN(n8000) );
  XNOR2_X1 U10050 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n7975) );
  XNOR2_X1 U10051 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n7931) );
  INV_X1 U10052 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U10053 ( .A1(n9659), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U10054 ( .A1(n7676), .A2(n7675), .ZN(n7774) );
  XNOR2_X1 U10055 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7772) );
  INV_X1 U10056 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U10057 ( .A1(n9661), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7677) );
  XNOR2_X1 U10058 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7785) );
  NAND2_X1 U10059 ( .A1(n7798), .A2(n7796), .ZN(n7679) );
  NAND2_X1 U10060 ( .A1(n9662), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U10061 ( .A1(n9686), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U10062 ( .A1(n9697), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U10063 ( .A1(n7682), .A2(n7681), .ZN(n7855) );
  NAND2_X1 U10064 ( .A1(n7855), .A2(n7854), .ZN(n7685) );
  INV_X1 U10065 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U10066 ( .A1(n7683), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U10067 ( .A1(n7685), .A2(n7684), .ZN(n7870) );
  NAND2_X1 U10068 ( .A1(n7870), .A2(n7868), .ZN(n7687) );
  NAND2_X1 U10069 ( .A1(n9719), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U10070 ( .A1(n7687), .A2(n7686), .ZN(n7886) );
  NAND2_X1 U10071 ( .A1(n9743), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7688) );
  INV_X1 U10072 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7690) );
  XNOR2_X1 U10073 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7914) );
  NAND2_X1 U10074 ( .A1(n9758), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U10075 ( .A1(n11167), .A2(n7696), .ZN(n7697) );
  XNOR2_X1 U10076 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7953) );
  NAND2_X1 U10077 ( .A1(n12990), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7698) );
  AOI22_X1 U10078 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n10360), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n10306), .ZN(n7988) );
  AOI22_X1 U10079 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10835), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n10786), .ZN(n8016) );
  INV_X1 U10080 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U10081 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11036), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n11034), .ZN(n8055) );
  AOI22_X1 U10082 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11320), .B2(n10084), .ZN(n8067) );
  INV_X1 U10083 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U10084 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11429), .B2(n10160), .ZN(n8078) );
  NAND2_X1 U10085 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7706), .ZN(n7707) );
  INV_X1 U10086 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14023) );
  NAND2_X1 U10087 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n14023), .ZN(n7708) );
  INV_X1 U10088 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U10089 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n14017), .B2(n12297), .ZN(n7709) );
  INV_X1 U10090 ( .A(n7709), .ZN(n7710) );
  XNOR2_X1 U10091 ( .A(n8100), .B(n7710), .ZN(n13280) );
  NOR2_X1 U10092 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n7712) );
  NAND2_X1 U10093 ( .A1(n7729), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7717) );
  XNOR2_X2 U10094 ( .A(n7717), .B(n7716), .ZN(n12302) );
  NAND3_X1 U10095 ( .A1(n14870), .A2(n7719), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7720) );
  NAND3_X1 U10096 ( .A1(n7722), .A2(n7721), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7724) );
  NAND2_X2 U10097 ( .A1(n7726), .A2(n7725), .ZN(n8324) );
  NAND2_X1 U10098 ( .A1(n13280), .A2(n11633), .ZN(n7728) );
  NAND2_X1 U10099 ( .A1(n9294), .A2(SI_26_), .ZN(n7727) );
  NAND2_X2 U10100 ( .A1(n7728), .A2(n7727), .ZN(n12715) );
  NAND2_X1 U10101 ( .A1(n7732), .A2(n7730), .ZN(n13267) );
  XNOR2_X2 U10102 ( .A(n7731), .B(n13268), .ZN(n7738) );
  AND2_X2 U10103 ( .A1(n7738), .A2(n6755), .ZN(n7778) );
  INV_X1 U10104 ( .A(n7778), .ZN(n8167) );
  NAND2_X1 U10105 ( .A1(n11636), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7742) );
  INV_X1 U10106 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12713) );
  OR2_X1 U10107 ( .A1(n8082), .A2(n12713), .ZN(n7741) );
  NAND2_X2 U10108 ( .A1(n6755), .A2(n7734), .ZN(n8108) );
  NOR2_X1 U10109 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7807) );
  INV_X1 U10110 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10111 ( .A1(n7807), .A2(n7808), .ZN(n7826) );
  NOR2_X1 U10112 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .ZN(n7735) );
  NAND2_X1 U10113 ( .A1(n7892), .A2(n7891), .ZN(n7908) );
  NOR2_X2 U10114 ( .A1(n7946), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10115 ( .A1(n7995), .A2(n14900), .ZN(n8008) );
  OR2_X2 U10116 ( .A1(n8008), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8027) );
  NOR2_X2 U10117 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n6619), .ZN(n8071) );
  INV_X1 U10118 ( .A(n8071), .ZN(n8084) );
  INV_X1 U10119 ( .A(n8083), .ZN(n8095) );
  INV_X1 U10120 ( .A(n8094), .ZN(n7749) );
  NOR2_X2 U10121 ( .A1(n7749), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7748) );
  INV_X1 U10122 ( .A(n7748), .ZN(n7736) );
  NOR2_X2 U10123 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n7736), .ZN(n8105) );
  AOI21_X1 U10124 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n7736), .A(n8105), .ZN(
        n12712) );
  OR2_X1 U10125 ( .A1(n8072), .A2(n12712), .ZN(n7740) );
  INV_X1 U10126 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13217) );
  OR2_X1 U10127 ( .A1(n6570), .A2(n13217), .ZN(n7739) );
  NAND2_X1 U10128 ( .A1(n12715), .A2(n12492), .ZN(n11813) );
  AOI22_X1 U10129 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n14023), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n12987), .ZN(n7743) );
  INV_X1 U10130 ( .A(n7743), .ZN(n7744) );
  XNOR2_X1 U10131 ( .A(n7745), .B(n7744), .ZN(n13286) );
  NAND2_X1 U10132 ( .A1(n13286), .A2(n11633), .ZN(n7747) );
  NAND2_X1 U10133 ( .A1(n9294), .A2(SI_25_), .ZN(n7746) );
  NAND2_X1 U10134 ( .A1(n11636), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7753) );
  INV_X1 U10135 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12729) );
  OR2_X1 U10136 ( .A1(n8082), .A2(n12729), .ZN(n7752) );
  AOI21_X1 U10137 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n7749), .A(n7748), .ZN(
        n12728) );
  OR2_X1 U10138 ( .A1(n8072), .A2(n12728), .ZN(n7751) );
  INV_X1 U10139 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13221) );
  OR2_X1 U10140 ( .A1(n6570), .A2(n13221), .ZN(n7750) );
  OR2_X1 U10141 ( .A1(n12727), .A2(n12523), .ZN(n11809) );
  NAND2_X1 U10142 ( .A1(n12727), .A2(n12523), .ZN(n11808) );
  NAND2_X1 U10143 ( .A1(n11809), .A2(n11808), .ZN(n12719) );
  INV_X1 U10144 ( .A(n12719), .ZN(n12726) );
  INV_X1 U10145 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7754) );
  INV_X1 U10146 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U10147 ( .A1(n7778), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7756) );
  XNOR2_X1 U10148 ( .A(n7760), .B(n7765), .ZN(n9665) );
  INV_X1 U10149 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10319) );
  OR2_X1 U10150 ( .A1(n8108), .A2(n10319), .ZN(n7763) );
  INV_X1 U10151 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10314) );
  OR2_X1 U10152 ( .A1(n8082), .A2(n10314), .ZN(n7762) );
  INV_X1 U10153 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n7761) );
  INV_X1 U10154 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9473) );
  AND2_X1 U10155 ( .A1(n9473), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7764) );
  NOR2_X1 U10156 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  INV_X1 U10157 ( .A(SI_0_), .ZN(n9474) );
  MUX2_X1 U10158 ( .A(n7766), .B(n9474), .S(n9680), .Z(n9658) );
  MUX2_X1 U10159 ( .A(n9616), .B(n9658), .S(n9625), .Z(n10349) );
  INV_X1 U10160 ( .A(n10349), .ZN(n7767) );
  INV_X1 U10161 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10136) );
  OR2_X1 U10162 ( .A1(n8108), .A2(n10136), .ZN(n7770) );
  INV_X1 U10163 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7768) );
  INV_X1 U10164 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15568) );
  OR2_X1 U10165 ( .A1(n8082), .A2(n15568), .ZN(n7769) );
  INV_X1 U10166 ( .A(SI_2_), .ZN(n9674) );
  NAND2_X1 U10167 ( .A1(n6603), .A2(n9674), .ZN(n7776) );
  INV_X1 U10168 ( .A(n7772), .ZN(n7773) );
  XNOR2_X1 U10169 ( .A(n7774), .B(n7773), .ZN(n9675) );
  NAND2_X1 U10170 ( .A1(n6622), .A2(n9675), .ZN(n7775) );
  OAI211_X1 U10171 ( .C1(n6572), .C2(n9625), .A(n7776), .B(n7775), .ZN(n15550)
         );
  NAND2_X1 U10172 ( .A1(n12601), .A2(n15550), .ZN(n11700) );
  NAND2_X1 U10173 ( .A1(n15549), .A2(n15555), .ZN(n7777) );
  NAND2_X1 U10174 ( .A1(n7777), .A2(n11692), .ZN(n10988) );
  INV_X1 U10175 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7779) );
  INV_X1 U10176 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7780) );
  OR2_X1 U10177 ( .A1(n8082), .A2(n7780), .ZN(n7781) );
  NAND2_X1 U10178 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7783), .ZN(n7784) );
  XNOR2_X1 U10179 ( .A(n7784), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9603) );
  INV_X1 U10180 ( .A(SI_3_), .ZN(n9672) );
  NAND2_X1 U10181 ( .A1(n6603), .A2(n9672), .ZN(n7788) );
  XNOR2_X1 U10182 ( .A(n7786), .B(n7203), .ZN(n9673) );
  NAND2_X1 U10183 ( .A1(n6622), .A2(n9673), .ZN(n7787) );
  OAI211_X1 U10184 ( .C1(n9603), .C2(n9625), .A(n7788), .B(n7787), .ZN(n15577)
         );
  NAND2_X1 U10185 ( .A1(n15461), .A2(n15577), .ZN(n11701) );
  NAND2_X1 U10186 ( .A1(n10988), .A2(n11658), .ZN(n10987) );
  NAND2_X1 U10187 ( .A1(n7778), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7795) );
  INV_X1 U10188 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7789) );
  OR2_X1 U10189 ( .A1(n8082), .A2(n7789), .ZN(n7794) );
  AND2_X1 U10190 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7790) );
  NOR2_X1 U10191 ( .A1(n7807), .A2(n7790), .ZN(n11148) );
  OR2_X1 U10192 ( .A1(n8108), .A2(n11148), .ZN(n7793) );
  INV_X1 U10193 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7791) );
  OR2_X1 U10194 ( .A1(n6569), .A2(n7791), .ZN(n7792) );
  INV_X1 U10195 ( .A(SI_4_), .ZN(n8330) );
  NAND2_X1 U10196 ( .A1(n6603), .A2(n8330), .ZN(n7804) );
  INV_X1 U10197 ( .A(n11624), .ZN(n8927) );
  INV_X1 U10198 ( .A(n7796), .ZN(n7797) );
  XNOR2_X1 U10199 ( .A(n7798), .B(n7797), .ZN(n14824) );
  NAND2_X1 U10200 ( .A1(n6622), .A2(n14824), .ZN(n7803) );
  NAND2_X1 U10201 ( .A1(n8038), .A2(n15504), .ZN(n7802) );
  INV_X1 U10202 ( .A(n11693), .ZN(n7806) );
  NOR2_X1 U10203 ( .A1(n12600), .A2(n15581), .ZN(n7805) );
  AOI21_X1 U10204 ( .B1(n11702), .B2(n7806), .A(n7805), .ZN(n11698) );
  NAND2_X1 U10205 ( .A1(n7778), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7814) );
  INV_X1 U10206 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15515) );
  OR2_X1 U10207 ( .A1(n8082), .A2(n15515), .ZN(n7813) );
  OR2_X1 U10208 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  AND2_X1 U10209 ( .A1(n7826), .A2(n7809), .ZN(n11120) );
  OR2_X1 U10210 ( .A1(n8108), .A2(n11120), .ZN(n7812) );
  INV_X1 U10211 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n7810) );
  OR2_X1 U10212 ( .A1(n6570), .A2(n7810), .ZN(n7811) );
  NAND4_X1 U10213 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n12599) );
  OR2_X1 U10214 ( .A1(n7817), .A2(n7883), .ZN(n7815) );
  MUX2_X1 U10215 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7815), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7818) );
  NAND2_X1 U10216 ( .A1(n7817), .A2(n7816), .ZN(n7836) );
  NAND2_X1 U10217 ( .A1(n7818), .A2(n7836), .ZN(n15512) );
  INV_X1 U10218 ( .A(SI_5_), .ZN(n7819) );
  NAND2_X1 U10219 ( .A1(n6603), .A2(n7819), .ZN(n7824) );
  INV_X1 U10220 ( .A(n7820), .ZN(n7821) );
  XNOR2_X1 U10221 ( .A(n7822), .B(n7821), .ZN(n14827) );
  NAND2_X1 U10222 ( .A1(n8927), .A2(n14827), .ZN(n7823) );
  OAI211_X1 U10223 ( .C1(n9636), .C2(n9625), .A(n7824), .B(n7823), .ZN(n15585)
         );
  NAND2_X1 U10224 ( .A1(n12599), .A2(n15585), .ZN(n11707) );
  NAND2_X1 U10225 ( .A1(n11119), .A2(n11657), .ZN(n11118) );
  NAND2_X1 U10226 ( .A1(n11118), .A2(n7825), .ZN(n10873) );
  NAND2_X1 U10227 ( .A1(n7778), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7832) );
  INV_X1 U10228 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10190) );
  OR2_X1 U10229 ( .A1(n11637), .A2(n10190), .ZN(n7831) );
  NAND2_X1 U10230 ( .A1(n7826), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7827) );
  AND2_X1 U10231 ( .A1(n7844), .A2(n7827), .ZN(n10881) );
  OR2_X1 U10232 ( .A1(n8108), .A2(n10881), .ZN(n7830) );
  INV_X1 U10233 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7828) );
  OR2_X1 U10234 ( .A1(n6570), .A2(n7828), .ZN(n7829) );
  NAND4_X1 U10235 ( .A1(n7832), .A2(n7831), .A3(n7830), .A4(n7829), .ZN(n12598) );
  NAND2_X1 U10236 ( .A1(n9294), .A2(SI_6_), .ZN(n7842) );
  XNOR2_X1 U10237 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7833) );
  XNOR2_X1 U10238 ( .A(n7834), .B(n7833), .ZN(n9676) );
  NAND2_X1 U10239 ( .A1(n8927), .A2(n9676), .ZN(n7841) );
  NAND2_X1 U10240 ( .A1(n7836), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7835) );
  MUX2_X1 U10241 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7835), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n7839) );
  INV_X1 U10242 ( .A(n7836), .ZN(n7838) );
  NAND2_X1 U10243 ( .A1(n7838), .A2(n7837), .ZN(n7850) );
  NAND2_X1 U10244 ( .A1(n8038), .A2(n10207), .ZN(n7840) );
  NAND2_X1 U10245 ( .A1(n12598), .A2(n15589), .ZN(n11706) );
  NAND2_X1 U10246 ( .A1(n11636), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7849) );
  INV_X1 U10247 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n7843) );
  OR2_X1 U10248 ( .A1(n6570), .A2(n7843), .ZN(n7848) );
  AND2_X1 U10249 ( .A1(n7844), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7845) );
  NOR2_X1 U10250 ( .A1(n7875), .A2(n7845), .ZN(n10982) );
  OR2_X1 U10251 ( .A1(n8072), .A2(n10982), .ZN(n7847) );
  INV_X1 U10252 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10981) );
  OR2_X1 U10253 ( .A1(n11637), .A2(n10981), .ZN(n7846) );
  NAND4_X1 U10254 ( .A1(n7849), .A2(n7848), .A3(n7847), .A4(n7846), .ZN(n12597) );
  NAND2_X1 U10255 ( .A1(n7850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7851) );
  MUX2_X1 U10256 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7851), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n7853) );
  AND2_X1 U10257 ( .A1(n7853), .A2(n7852), .ZN(n10197) );
  XNOR2_X1 U10258 ( .A(n7855), .B(n7854), .ZN(n9664) );
  NAND2_X1 U10259 ( .A1(n11633), .A2(n9664), .ZN(n7857) );
  INV_X1 U10260 ( .A(SI_7_), .ZN(n9663) );
  NAND2_X1 U10261 ( .A1(n9294), .A2(n9663), .ZN(n7856) );
  OAI211_X1 U10262 ( .C1(n10197), .C2(n9625), .A(n7857), .B(n7856), .ZN(n15594) );
  OR2_X1 U10263 ( .A1(n12597), .A2(n15594), .ZN(n11715) );
  NAND2_X1 U10264 ( .A1(n12597), .A2(n15594), .ZN(n11714) );
  NAND2_X1 U10265 ( .A1(n10976), .A2(n11708), .ZN(n7858) );
  NAND2_X1 U10266 ( .A1(n11636), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7863) );
  INV_X1 U10267 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n7859) );
  OR2_X1 U10268 ( .A1(n6570), .A2(n7859), .ZN(n7862) );
  XNOR2_X1 U10269 ( .A(n7875), .B(P3_REG3_REG_8__SCAN_IN), .ZN(n10925) );
  OR2_X1 U10270 ( .A1(n8072), .A2(n10925), .ZN(n7861) );
  INV_X1 U10271 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11046) );
  OR2_X1 U10272 ( .A1(n11637), .A2(n11046), .ZN(n7860) );
  NAND4_X1 U10273 ( .A1(n7863), .A2(n7862), .A3(n7861), .A4(n7860), .ZN(n12596) );
  NAND2_X1 U10274 ( .A1(n7852), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U10275 ( .A(n7865), .B(P3_IR_REG_31__SCAN_IN), .S(n7864), .Z(n7867)
         );
  NOR2_X1 U10276 ( .A1(n7852), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7900) );
  INV_X1 U10277 ( .A(n7900), .ZN(n7866) );
  NAND2_X1 U10278 ( .A1(n7867), .A2(n7866), .ZN(n14832) );
  NAND2_X1 U10279 ( .A1(n9294), .A2(SI_8_), .ZN(n7872) );
  INV_X1 U10280 ( .A(n7868), .ZN(n7869) );
  XNOR2_X1 U10281 ( .A(n7870), .B(n7869), .ZN(n14830) );
  NAND2_X1 U10282 ( .A1(n11633), .A2(n14830), .ZN(n7871) );
  OAI211_X1 U10283 ( .C1(n9625), .C2(n14832), .A(n7872), .B(n7871), .ZN(n11721) );
  INV_X1 U10284 ( .A(n11721), .ZN(n15601) );
  NOR2_X1 U10285 ( .A1(n12596), .A2(n15601), .ZN(n7873) );
  NAND2_X1 U10286 ( .A1(n12596), .A2(n15601), .ZN(n7874) );
  NAND2_X1 U10287 ( .A1(n11636), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7882) );
  INV_X1 U10288 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10423) );
  OR2_X1 U10289 ( .A1(n11637), .A2(n10423), .ZN(n7881) );
  INV_X1 U10290 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10926) );
  INV_X1 U10291 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11082) );
  AOI21_X1 U10292 ( .B1(n7875), .B2(n10926), .A(n11082), .ZN(n7876) );
  OR2_X1 U10293 ( .A1(n7892), .A2(n7876), .ZN(n11100) );
  INV_X1 U10294 ( .A(n11100), .ZN(n7877) );
  OR2_X1 U10295 ( .A1(n8072), .A2(n7877), .ZN(n7880) );
  INV_X1 U10296 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n7878) );
  OR2_X1 U10297 ( .A1(n6570), .A2(n7878), .ZN(n7879) );
  NAND4_X1 U10298 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n12595) );
  OR2_X1 U10299 ( .A1(n7900), .A2(n7883), .ZN(n7884) );
  XNOR2_X1 U10300 ( .A(n7884), .B(P3_IR_REG_9__SCAN_IN), .ZN(n10424) );
  INV_X1 U10301 ( .A(SI_9_), .ZN(n9670) );
  NAND2_X1 U10302 ( .A1(n9294), .A2(n9670), .ZN(n7888) );
  XNOR2_X1 U10303 ( .A(n7886), .B(n7885), .ZN(n9671) );
  NAND2_X1 U10304 ( .A1(n11633), .A2(n9671), .ZN(n7887) );
  OAI211_X1 U10305 ( .C1(n10424), .C2(n9625), .A(n7888), .B(n7887), .ZN(n15607) );
  OR2_X1 U10306 ( .A1(n12595), .A2(n15607), .ZN(n11728) );
  NAND2_X1 U10307 ( .A1(n12595), .A2(n15607), .ZN(n11727) );
  NAND2_X1 U10308 ( .A1(n11636), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7898) );
  INV_X1 U10309 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11208) );
  OR2_X1 U10310 ( .A1(n8082), .A2(n11208), .ZN(n7897) );
  OR2_X1 U10311 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  AND2_X1 U10312 ( .A1(n7908), .A2(n7893), .ZN(n11276) );
  OR2_X1 U10313 ( .A1(n8072), .A2(n11276), .ZN(n7896) );
  INV_X1 U10314 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n7894) );
  OR2_X1 U10315 ( .A1(n6570), .A2(n7894), .ZN(n7895) );
  NAND4_X1 U10316 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n12594) );
  NAND2_X1 U10317 ( .A1(n7900), .A2(n7899), .ZN(n7916) );
  NAND2_X1 U10318 ( .A1(n7916), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7902) );
  INV_X1 U10319 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7901) );
  INV_X1 U10320 ( .A(n10945), .ZN(n10773) );
  NAND2_X1 U10321 ( .A1(n9294), .A2(n9668), .ZN(n7906) );
  XNOR2_X1 U10322 ( .A(n7904), .B(n7903), .ZN(n9669) );
  NAND2_X1 U10323 ( .A1(n11633), .A2(n9669), .ZN(n7905) );
  OAI211_X1 U10324 ( .C1(n10773), .C2(n9625), .A(n7906), .B(n7905), .ZN(n11281) );
  OR2_X1 U10325 ( .A1(n12594), .A2(n11281), .ZN(n11734) );
  NAND2_X1 U10326 ( .A1(n12594), .A2(n11281), .ZN(n11733) );
  NAND2_X1 U10327 ( .A1(n11734), .A2(n11733), .ZN(n11731) );
  NAND2_X1 U10328 ( .A1(n11207), .A2(n11664), .ZN(n11206) );
  NAND2_X1 U10329 ( .A1(n7778), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7913) );
  INV_X1 U10330 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n7907) );
  OR2_X1 U10331 ( .A1(n6570), .A2(n7907), .ZN(n7912) );
  NAND2_X1 U10332 ( .A1(n7908), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7909) );
  AND2_X1 U10333 ( .A1(n7925), .A2(n7909), .ZN(n11479) );
  OR2_X1 U10334 ( .A1(n8072), .A2(n11479), .ZN(n7911) );
  INV_X1 U10335 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11313) );
  OR2_X1 U10336 ( .A1(n8082), .A2(n11313), .ZN(n7910) );
  NAND4_X1 U10337 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n12593) );
  XNOR2_X1 U10338 ( .A(n7915), .B(n7914), .ZN(n14833) );
  NAND2_X1 U10339 ( .A1(n14833), .A2(n11633), .ZN(n7923) );
  NAND2_X1 U10340 ( .A1(n7918), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7917) );
  MUX2_X1 U10341 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7917), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n7921) );
  INV_X1 U10342 ( .A(n7918), .ZN(n7920) );
  INV_X1 U10343 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10344 ( .A1(n7920), .A2(n7919), .ZN(n7934) );
  NAND2_X1 U10345 ( .A1(n7921), .A2(n7934), .ZN(n14838) );
  AOI22_X1 U10346 ( .A1(n9294), .A2(n8350), .B1(n8038), .B2(n14838), .ZN(n7922) );
  NAND2_X1 U10347 ( .A1(n7923), .A2(n7922), .ZN(n11326) );
  OR2_X1 U10348 ( .A1(n12593), .A2(n11326), .ZN(n11740) );
  NAND2_X1 U10349 ( .A1(n12593), .A2(n11326), .ZN(n11744) );
  NAND2_X1 U10350 ( .A1(n11740), .A2(n11744), .ZN(n11742) );
  INV_X1 U10351 ( .A(n11742), .ZN(n11311) );
  NAND2_X1 U10352 ( .A1(n7778), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7930) );
  INV_X1 U10353 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n7924) );
  OR2_X1 U10354 ( .A1(n6570), .A2(n7924), .ZN(n7929) );
  NAND2_X1 U10355 ( .A1(n7925), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7926) );
  AND2_X1 U10356 ( .A1(n7946), .A2(n7926), .ZN(n11412) );
  OR2_X1 U10357 ( .A1(n8072), .A2(n11412), .ZN(n7928) );
  INV_X1 U10358 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11053) );
  OR2_X1 U10359 ( .A1(n11637), .A2(n11053), .ZN(n7927) );
  INV_X1 U10360 ( .A(n7931), .ZN(n7932) );
  XNOR2_X1 U10361 ( .A(n7933), .B(n7932), .ZN(n9688) );
  NAND2_X1 U10362 ( .A1(n9688), .A2(n11633), .ZN(n7940) );
  NAND2_X1 U10363 ( .A1(n7934), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7935) );
  MUX2_X1 U10364 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7935), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7938) );
  INV_X1 U10365 ( .A(n7936), .ZN(n7937) );
  AOI22_X1 U10366 ( .A1(n9294), .A2(SI_12_), .B1(n8038), .B2(n11068), .ZN(
        n7939) );
  NAND2_X1 U10367 ( .A1(n7940), .A2(n7939), .ZN(n8142) );
  OR2_X1 U10368 ( .A1(n11517), .A2(n8142), .ZN(n11746) );
  NAND2_X1 U10369 ( .A1(n11517), .A2(n8142), .ZN(n11749) );
  NAND2_X1 U10370 ( .A1(n11411), .A2(n11410), .ZN(n11409) );
  NAND2_X1 U10371 ( .A1(n11409), .A2(n11749), .ZN(n11521) );
  XNOR2_X1 U10372 ( .A(n7941), .B(n10027), .ZN(n9744) );
  NAND2_X1 U10373 ( .A1(n9744), .A2(n11633), .ZN(n7944) );
  OR2_X1 U10374 ( .A1(n7936), .A2(n7883), .ZN(n7942) );
  XNOR2_X1 U10375 ( .A(n7942), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U10376 ( .A1(n9294), .A2(SI_13_), .B1(n8038), .B2(n12619), .ZN(
        n7943) );
  NAND2_X1 U10377 ( .A1(n7944), .A2(n7943), .ZN(n11908) );
  NAND2_X1 U10378 ( .A1(n7778), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7952) );
  INV_X1 U10379 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n7945) );
  OR2_X1 U10380 ( .A1(n11637), .A2(n7945), .ZN(n7951) );
  AND2_X1 U10381 ( .A1(n7946), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7947) );
  NOR2_X1 U10382 ( .A1(n7965), .A2(n7947), .ZN(n11906) );
  OR2_X1 U10383 ( .A1(n8072), .A2(n11906), .ZN(n7950) );
  INV_X1 U10384 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n7948) );
  OR2_X1 U10385 ( .A1(n6570), .A2(n7948), .ZN(n7949) );
  OR2_X1 U10386 ( .A1(n11908), .A2(n11899), .ZN(n11757) );
  NAND2_X1 U10387 ( .A1(n11908), .A2(n11899), .ZN(n11752) );
  NAND2_X1 U10388 ( .A1(n11568), .A2(n11752), .ZN(n7974) );
  XNOR2_X1 U10389 ( .A(n7954), .B(n7953), .ZN(n9750) );
  NAND2_X1 U10390 ( .A1(n9750), .A2(n11633), .ZN(n7962) );
  NOR2_X1 U10391 ( .A1(n7956), .A2(n7883), .ZN(n7957) );
  MUX2_X1 U10392 ( .A(n7883), .B(n7957), .S(P3_IR_REG_14__SCAN_IN), .Z(n7958)
         );
  INV_X1 U10393 ( .A(n7958), .ZN(n7960) );
  NAND2_X1 U10394 ( .A1(n7960), .A2(n7959), .ZN(n12648) );
  AOI22_X1 U10395 ( .A1(n9294), .A2(n9749), .B1(n8038), .B2(n12648), .ZN(n7961) );
  NAND2_X1 U10396 ( .A1(n11636), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7972) );
  INV_X1 U10397 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n7963) );
  OR2_X1 U10398 ( .A1(n11637), .A2(n7963), .ZN(n7971) );
  NOR2_X1 U10399 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  OR2_X1 U10400 ( .A1(n7981), .A2(n7966), .ZN(n12463) );
  INV_X1 U10401 ( .A(n12463), .ZN(n7967) );
  OR2_X1 U10402 ( .A1(n8072), .A2(n7967), .ZN(n7970) );
  INV_X1 U10403 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n7968) );
  OR2_X1 U10404 ( .A1(n6570), .A2(n7968), .ZN(n7969) );
  OR2_X1 U10405 ( .A1(n13260), .A2(n12566), .ZN(n12858) );
  NAND2_X1 U10406 ( .A1(n13260), .A2(n12566), .ZN(n7973) );
  NAND2_X1 U10407 ( .A1(n12858), .A2(n7973), .ZN(n11756) );
  NAND2_X1 U10408 ( .A1(n7974), .A2(n11756), .ZN(n11570) );
  OR2_X1 U10409 ( .A1(n13260), .A2(n12590), .ZN(n11755) );
  INV_X1 U10410 ( .A(n7975), .ZN(n7976) );
  XNOR2_X1 U10411 ( .A(n7977), .B(n7976), .ZN(n9872) );
  NAND2_X1 U10412 ( .A1(n9872), .A2(n11633), .ZN(n7980) );
  NAND2_X1 U10413 ( .A1(n7959), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7978) );
  XNOR2_X1 U10414 ( .A(n7978), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U10415 ( .A1(n9294), .A2(SI_15_), .B1(n8038), .B2(n12649), .ZN(
        n7979) );
  NAND2_X1 U10416 ( .A1(n7980), .A2(n7979), .ZN(n12562) );
  NAND2_X1 U10417 ( .A1(n7778), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7987) );
  INV_X1 U10418 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14878) );
  OR2_X1 U10419 ( .A1(n11637), .A2(n14878), .ZN(n7986) );
  NOR2_X1 U10420 ( .A1(n7981), .A2(n12570), .ZN(n7982) );
  OR2_X1 U10421 ( .A1(n7995), .A2(n7982), .ZN(n12868) );
  INV_X1 U10422 ( .A(n12868), .ZN(n7983) );
  OR2_X1 U10423 ( .A1(n8108), .A2(n7983), .ZN(n7985) );
  INV_X1 U10424 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13255) );
  OR2_X1 U10425 ( .A1(n6570), .A2(n13255), .ZN(n7984) );
  OR2_X1 U10426 ( .A1(n12562), .A2(n11563), .ZN(n11761) );
  NAND2_X1 U10427 ( .A1(n12562), .A2(n11563), .ZN(n11762) );
  INV_X1 U10428 ( .A(n7988), .ZN(n7989) );
  XNOR2_X1 U10429 ( .A(n7990), .B(n7989), .ZN(n10000) );
  NAND2_X1 U10430 ( .A1(n10000), .A2(n11633), .ZN(n7994) );
  NAND2_X1 U10431 ( .A1(n7991), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7992) );
  XNOR2_X1 U10432 ( .A(n7992), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U10433 ( .A1(n9294), .A2(SI_16_), .B1(n8038), .B2(n12652), .ZN(
        n7993) );
  NAND2_X1 U10434 ( .A1(n7994), .A2(n7993), .ZN(n12505) );
  NAND2_X1 U10435 ( .A1(n7778), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7999) );
  OR2_X1 U10436 ( .A1(n11637), .A2(n13162), .ZN(n7998) );
  XNOR2_X1 U10437 ( .A(n7995), .B(P3_REG3_REG_16__SCAN_IN), .ZN(n12852) );
  OR2_X1 U10438 ( .A1(n8072), .A2(n12852), .ZN(n7997) );
  INV_X1 U10439 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13251) );
  OR2_X1 U10440 ( .A1(n6570), .A2(n13251), .ZN(n7996) );
  OR2_X1 U10441 ( .A1(n12505), .A2(n12567), .ZN(n11767) );
  NAND2_X1 U10442 ( .A1(n12505), .A2(n12567), .ZN(n11768) );
  INV_X1 U10443 ( .A(n8000), .ZN(n8001) );
  XNOR2_X1 U10444 ( .A(n8002), .B(n8001), .ZN(n10029) );
  NAND2_X1 U10445 ( .A1(n10029), .A2(n11633), .ZN(n8007) );
  NAND2_X1 U10446 ( .A1(n8004), .A2(n8003), .ZN(n8019) );
  NAND2_X1 U10447 ( .A1(n8019), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8005) );
  XNOR2_X1 U10448 ( .A(n8005), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U10449 ( .A1(n9294), .A2(SI_17_), .B1(n8038), .B2(n14925), .ZN(
        n8006) );
  NAND2_X1 U10450 ( .A1(n8007), .A2(n8006), .ZN(n12835) );
  NAND2_X1 U10451 ( .A1(n7778), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10452 ( .A1(n8008), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8009) );
  AND2_X1 U10453 ( .A1(n8027), .A2(n8009), .ZN(n12836) );
  OR2_X1 U10454 ( .A1(n12836), .A2(n8072), .ZN(n8012) );
  INV_X1 U10455 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14916) );
  OR2_X1 U10456 ( .A1(n11637), .A2(n14916), .ZN(n8011) );
  INV_X1 U10457 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13247) );
  OR2_X1 U10458 ( .A1(n6570), .A2(n13247), .ZN(n8010) );
  NOR2_X1 U10459 ( .A1(n12835), .A2(n12509), .ZN(n11773) );
  INV_X1 U10460 ( .A(n11773), .ZN(n8014) );
  NAND2_X1 U10461 ( .A1(n12835), .A2(n12509), .ZN(n11778) );
  NAND2_X1 U10462 ( .A1(n8014), .A2(n11778), .ZN(n12828) );
  NAND2_X1 U10463 ( .A1(n12834), .A2(n7552), .ZN(n8015) );
  INV_X1 U10464 ( .A(n8016), .ZN(n8017) );
  XNOR2_X1 U10465 ( .A(n8018), .B(n8017), .ZN(n10080) );
  NAND2_X1 U10466 ( .A1(n10080), .A2(n11633), .ZN(n8026) );
  NAND2_X1 U10467 ( .A1(n7666), .A2(n8020), .ZN(n8021) );
  NAND2_X1 U10468 ( .A1(n8021), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8022) );
  MUX2_X1 U10469 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8022), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8024) );
  NAND2_X1 U10470 ( .A1(n8024), .A2(n8023), .ZN(n12657) );
  INV_X1 U10471 ( .A(n12657), .ZN(n12666) );
  AOI22_X1 U10472 ( .A1(n9294), .A2(SI_18_), .B1(n8038), .B2(n12666), .ZN(
        n8025) );
  NAND2_X1 U10473 ( .A1(n8026), .A2(n8025), .ZN(n12910) );
  INV_X1 U10474 ( .A(n8072), .ZN(n8061) );
  INV_X1 U10475 ( .A(n8044), .ZN(n8029) );
  NAND2_X1 U10476 ( .A1(n8027), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10477 ( .A1(n8029), .A2(n8028), .ZN(n12821) );
  AND2_X1 U10478 ( .A1(n8061), .A2(n12821), .ZN(n8035) );
  INV_X1 U10479 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8030) );
  NOR2_X1 U10480 ( .A1(n6570), .A2(n8030), .ZN(n8034) );
  INV_X1 U10481 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10482 ( .A1(n11636), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8031) );
  OAI21_X1 U10483 ( .B1(n8032), .B2(n11637), .A(n8031), .ZN(n8033) );
  OR2_X1 U10484 ( .A1(n12910), .A2(n12517), .ZN(n11775) );
  NAND2_X1 U10485 ( .A1(n12910), .A2(n12517), .ZN(n11776) );
  XNOR2_X1 U10486 ( .A(n8037), .B(n8036), .ZN(n10157) );
  NAND2_X1 U10487 ( .A1(n10157), .A2(n11633), .ZN(n8040) );
  AOI22_X1 U10488 ( .A1(n9294), .A2(n10158), .B1(n8038), .B2(n12673), .ZN(
        n8039) );
  INV_X1 U10489 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13242) );
  NAND2_X1 U10490 ( .A1(n11636), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8042) );
  INV_X1 U10491 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13049) );
  OR2_X1 U10492 ( .A1(n11637), .A2(n13049), .ZN(n8041) );
  AND2_X1 U10493 ( .A1(n8042), .A2(n8041), .ZN(n8047) );
  NOR2_X1 U10494 ( .A1(n8044), .A2(n8043), .ZN(n8045) );
  OR2_X1 U10495 ( .A1(n8050), .A2(n8045), .ZN(n12809) );
  NAND2_X1 U10496 ( .A1(n12809), .A2(n8061), .ZN(n8046) );
  OAI211_X1 U10497 ( .C1(n6570), .C2(n13242), .A(n8047), .B(n8046), .ZN(n12588) );
  NAND2_X1 U10498 ( .A1(n13244), .A2(n12588), .ZN(n11785) );
  OR2_X1 U10499 ( .A1(n13244), .A2(n12588), .ZN(n11784) );
  INV_X1 U10500 ( .A(n12795), .ZN(n8054) );
  XNOR2_X1 U10501 ( .A(n8048), .B(n10872), .ZN(n10552) );
  AND2_X1 U10502 ( .A1(n9294), .A2(SI_20_), .ZN(n8049) );
  AOI21_X2 U10503 ( .B1(n10552), .B2(n11633), .A(n8049), .ZN(n13240) );
  INV_X1 U10504 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13238) );
  OR2_X1 U10505 ( .A1(n8050), .A2(n12537), .ZN(n8051) );
  NAND2_X1 U10506 ( .A1(n8059), .A2(n8051), .ZN(n12797) );
  NAND2_X1 U10507 ( .A1(n12797), .A2(n8061), .ZN(n8053) );
  AOI22_X1 U10508 ( .A1(n8166), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n11636), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8052) );
  OAI211_X1 U10509 ( .C1(n6570), .C2(n13238), .A(n8053), .B(n8052), .ZN(n12587) );
  NAND2_X1 U10510 ( .A1(n13240), .A2(n12587), .ZN(n11790) );
  INV_X1 U10511 ( .A(n13240), .ZN(n8151) );
  INV_X1 U10512 ( .A(n12587), .ZN(n12486) );
  NAND2_X1 U10513 ( .A1(n8151), .A2(n12486), .ZN(n11791) );
  XNOR2_X1 U10514 ( .A(n8056), .B(n7218), .ZN(n10787) );
  NAND2_X1 U10515 ( .A1(n10787), .A2(n11633), .ZN(n8058) );
  NAND2_X1 U10516 ( .A1(n9294), .A2(SI_21_), .ZN(n8057) );
  INV_X1 U10517 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10518 ( .A1(n8059), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10519 ( .A1(n8060), .A2(n6619), .ZN(n12782) );
  NAND2_X1 U10520 ( .A1(n12782), .A2(n8061), .ZN(n8063) );
  AOI22_X1 U10521 ( .A1(n6798), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n11636), 
        .B2(P3_REG1_REG_21__SCAN_IN), .ZN(n8062) );
  OAI211_X1 U10522 ( .C1(n11637), .C2(n8064), .A(n8063), .B(n8062), .ZN(n12586) );
  INV_X1 U10523 ( .A(n12586), .ZN(n12546) );
  NAND2_X1 U10524 ( .A1(n12781), .A2(n12546), .ZN(n8065) );
  XNOR2_X1 U10525 ( .A(n8068), .B(n8067), .ZN(n10869) );
  NAND2_X1 U10526 ( .A1(n10869), .A2(n11633), .ZN(n8070) );
  NAND2_X1 U10527 ( .A1(n9294), .A2(SI_22_), .ZN(n8069) );
  NAND2_X1 U10528 ( .A1(n11636), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8076) );
  INV_X1 U10529 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12770) );
  OR2_X1 U10530 ( .A1(n8082), .A2(n12770), .ZN(n8075) );
  AOI21_X1 U10531 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(n6619), .A(n8071), .ZN(
        n12769) );
  OR2_X1 U10532 ( .A1(n8072), .A2(n12769), .ZN(n8074) );
  INV_X1 U10533 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13230) );
  OR2_X1 U10534 ( .A1(n6570), .A2(n13230), .ZN(n8073) );
  NAND2_X1 U10535 ( .A1(n12768), .A2(n12485), .ZN(n11678) );
  INV_X1 U10536 ( .A(n11678), .ZN(n8077) );
  OR2_X1 U10537 ( .A1(n12768), .A2(n12485), .ZN(n11679) );
  XNOR2_X1 U10538 ( .A(n8079), .B(n8078), .ZN(n11088) );
  NAND2_X1 U10539 ( .A1(n11088), .A2(n11633), .ZN(n8081) );
  NAND2_X1 U10540 ( .A1(n9294), .A2(SI_23_), .ZN(n8080) );
  NAND2_X1 U10541 ( .A1(n11636), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8089) );
  INV_X1 U10542 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12755) );
  OR2_X1 U10543 ( .A1(n8082), .A2(n12755), .ZN(n8088) );
  AOI21_X1 U10544 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(n8084), .A(n8083), .ZN(
        n12754) );
  OR2_X1 U10545 ( .A1(n8072), .A2(n12754), .ZN(n8087) );
  INV_X1 U10546 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n8085) );
  OR2_X1 U10547 ( .A1(n6570), .A2(n8085), .ZN(n8086) );
  NAND4_X1 U10548 ( .A1(n8089), .A2(n8088), .A3(n8087), .A4(n8086), .ZN(n12584) );
  NAND2_X1 U10549 ( .A1(n12892), .A2(n12584), .ZN(n11802) );
  INV_X1 U10550 ( .A(n11802), .ZN(n8090) );
  XOR2_X1 U10551 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8091), .Z(n11462) );
  NAND2_X1 U10552 ( .A1(n11462), .A2(n11633), .ZN(n8093) );
  NAND2_X1 U10553 ( .A1(n9294), .A2(SI_24_), .ZN(n8092) );
  NAND2_X2 U10554 ( .A1(n8093), .A2(n8092), .ZN(n12744) );
  NAND2_X1 U10555 ( .A1(n11636), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8099) );
  INV_X1 U10556 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12746) );
  OR2_X1 U10557 ( .A1(n11637), .A2(n12746), .ZN(n8098) );
  AOI21_X1 U10558 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n8095), .A(n8094), .ZN(
        n12745) );
  OR2_X1 U10559 ( .A1(n8072), .A2(n12745), .ZN(n8097) );
  INV_X1 U10560 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13225) );
  OR2_X1 U10561 ( .A1(n6570), .A2(n13225), .ZN(n8096) );
  NAND4_X1 U10562 ( .A1(n8099), .A2(n8098), .A3(n8097), .A4(n8096), .ZN(n12583) );
  XNOR2_X1 U10563 ( .A(n12744), .B(n12583), .ZN(n12741) );
  INV_X1 U10564 ( .A(n12583), .ZN(n9371) );
  NAND2_X1 U10565 ( .A1(n12744), .A2(n9371), .ZN(n11803) );
  NOR2_X1 U10566 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n12297), .ZN(n8101) );
  OAI22_X1 U10567 ( .A1(n8101), .A2(n8100), .B1(P2_DATAO_REG_26__SCAN_IN), 
        .B2(n14017), .ZN(n8923) );
  INV_X1 U10568 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14016) );
  INV_X1 U10569 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8925) );
  AOI22_X1 U10570 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n14016), .B2(n8925), .ZN(n8102) );
  XNOR2_X1 U10571 ( .A(n8923), .B(n8102), .ZN(n13276) );
  NAND2_X1 U10572 ( .A1(n13276), .A2(n11633), .ZN(n8104) );
  NAND2_X1 U10573 ( .A1(n9294), .A2(SI_27_), .ZN(n8103) );
  NAND2_X1 U10574 ( .A1(n11636), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8112) );
  INV_X1 U10575 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12699) );
  OR2_X1 U10576 ( .A1(n11637), .A2(n12699), .ZN(n8111) );
  INV_X1 U10577 ( .A(n8105), .ZN(n8106) );
  AND2_X1 U10578 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8106), .ZN(n8107) );
  NOR2_X1 U10579 ( .A1(n8169), .A2(n8107), .ZN(n12698) );
  OR2_X1 U10580 ( .A1(n8072), .A2(n12698), .ZN(n8110) );
  INV_X1 U10581 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13213) );
  OR2_X1 U10582 ( .A1(n6570), .A2(n13213), .ZN(n8109) );
  INV_X1 U10583 ( .A(n10555), .ZN(n8945) );
  OR2_X1 U10584 ( .A1(n8945), .A2(n11682), .ZN(n8222) );
  XNOR2_X1 U10585 ( .A(n8222), .B(n11841), .ZN(n8117) );
  OR2_X1 U10586 ( .A1(n11682), .A2(n8115), .ZN(n8116) );
  NAND2_X1 U10587 ( .A1(n8117), .A2(n8116), .ZN(n9396) );
  NAND2_X1 U10588 ( .A1(n10555), .A2(n12673), .ZN(n11834) );
  INV_X1 U10589 ( .A(n11834), .ZN(n11838) );
  AND2_X1 U10590 ( .A1(n15606), .A2(n11838), .ZN(n8118) );
  NAND2_X1 U10591 ( .A1(n9396), .A2(n8118), .ZN(n8120) );
  AND2_X1 U10592 ( .A1(n12673), .A2(n11841), .ZN(n8119) );
  NAND2_X1 U10593 ( .A1(n11834), .A2(n8119), .ZN(n8227) );
  NAND2_X1 U10594 ( .A1(n15556), .A2(n15554), .ZN(n8125) );
  NAND2_X1 U10595 ( .A1(n8125), .A2(n8124), .ZN(n15558) );
  INV_X1 U10596 ( .A(n15550), .ZN(n15462) );
  OR2_X1 U10597 ( .A1(n6822), .A2(n15462), .ZN(n8126) );
  NAND2_X1 U10598 ( .A1(n15558), .A2(n8126), .ZN(n10990) );
  INV_X1 U10599 ( .A(n10990), .ZN(n8128) );
  INV_X1 U10600 ( .A(n15577), .ZN(n10999) );
  NAND2_X1 U10601 ( .A1(n15461), .A2(n10999), .ZN(n8129) );
  NAND2_X1 U10602 ( .A1(n10992), .A2(n8129), .ZN(n11149) );
  NAND2_X1 U10603 ( .A1(n11149), .A2(n11660), .ZN(n8131) );
  NAND2_X1 U10604 ( .A1(n12600), .A2(n10413), .ZN(n8130) );
  INV_X1 U10605 ( .A(n15589), .ZN(n8132) );
  AND2_X1 U10606 ( .A1(n12598), .A2(n8132), .ZN(n8133) );
  OR2_X1 U10607 ( .A1(n11657), .A2(n8133), .ZN(n8135) );
  OR2_X1 U10608 ( .A1(n12599), .A2(n6736), .ZN(n10874) );
  OR2_X1 U10609 ( .A1(n8133), .A2(n10875), .ZN(n8134) );
  INV_X1 U10610 ( .A(n11708), .ZN(n10975) );
  INV_X1 U10611 ( .A(n15594), .ZN(n10984) );
  NAND2_X1 U10612 ( .A1(n12597), .A2(n10984), .ZN(n8136) );
  NAND2_X1 U10613 ( .A1(n8137), .A2(n8136), .ZN(n11042) );
  OR2_X1 U10614 ( .A1(n12596), .A2(n11721), .ZN(n11039) );
  NAND2_X1 U10615 ( .A1(n11042), .A2(n11039), .ZN(n8138) );
  NAND2_X1 U10616 ( .A1(n12596), .A2(n11721), .ZN(n11038) );
  INV_X1 U10617 ( .A(n15607), .ZN(n11101) );
  INV_X1 U10618 ( .A(n11281), .ZN(n11273) );
  INV_X1 U10619 ( .A(n11326), .ZN(n11482) );
  OR2_X1 U10620 ( .A1(n12593), .A2(n11482), .ZN(n8139) );
  NAND2_X1 U10621 ( .A1(n11306), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U10622 ( .A1(n12593), .A2(n11482), .ZN(n8140) );
  NAND2_X1 U10623 ( .A1(n8141), .A2(n8140), .ZN(n11405) );
  NAND2_X1 U10624 ( .A1(n11557), .A2(n11517), .ZN(n8144) );
  INV_X1 U10625 ( .A(n11899), .ZN(n12591) );
  NAND2_X1 U10626 ( .A1(n11908), .A2(n12591), .ZN(n11560) );
  OR2_X1 U10627 ( .A1(n11756), .A2(n11560), .ZN(n11558) );
  INV_X1 U10628 ( .A(n12866), .ZN(n8145) );
  NAND2_X1 U10629 ( .A1(n8146), .A2(n8145), .ZN(n12862) );
  NAND2_X1 U10630 ( .A1(n12562), .A2(n12848), .ZN(n8147) );
  INV_X1 U10631 ( .A(n12842), .ZN(n12845) );
  INV_X1 U10632 ( .A(n12567), .ZN(n12831) );
  NAND2_X1 U10633 ( .A1(n12505), .A2(n12831), .ZN(n8148) );
  INV_X1 U10634 ( .A(n12509), .ZN(n12847) );
  NAND2_X1 U10635 ( .A1(n11775), .A2(n11776), .ZN(n11777) );
  NAND2_X1 U10636 ( .A1(n11784), .A2(n11785), .ZN(n12804) );
  OR2_X1 U10637 ( .A1(n12910), .A2(n12830), .ZN(n12805) );
  AND2_X1 U10638 ( .A1(n12804), .A2(n12805), .ZN(n8150) );
  INV_X1 U10639 ( .A(n12588), .ZN(n9359) );
  OR2_X1 U10640 ( .A1(n13244), .A2(n9359), .ZN(n12787) );
  NAND2_X1 U10641 ( .A1(n8151), .A2(n12587), .ZN(n8152) );
  NAND2_X1 U10642 ( .A1(n12781), .A2(n12586), .ZN(n11654) );
  INV_X1 U10643 ( .A(n11654), .ZN(n8153) );
  OR2_X1 U10644 ( .A1(n12781), .A2(n12586), .ZN(n11655) );
  NAND2_X1 U10645 ( .A1(n12768), .A2(n12585), .ZN(n8154) );
  OR2_X1 U10646 ( .A1(n12768), .A2(n12585), .ZN(n8155) );
  NAND2_X1 U10647 ( .A1(n12757), .A2(n12584), .ZN(n8157) );
  INV_X1 U10648 ( .A(n12741), .ZN(n12735) );
  NAND2_X1 U10649 ( .A1(n12736), .A2(n12735), .ZN(n12734) );
  NAND2_X1 U10650 ( .A1(n12744), .A2(n12583), .ZN(n8158) );
  NAND2_X1 U10651 ( .A1(n12734), .A2(n8158), .ZN(n12720) );
  NAND2_X1 U10652 ( .A1(n12727), .A2(n12582), .ZN(n8159) );
  OR2_X1 U10653 ( .A1(n12715), .A2(n12581), .ZN(n8160) );
  NAND2_X1 U10654 ( .A1(n12709), .A2(n8160), .ZN(n8162) );
  NAND2_X1 U10655 ( .A1(n12715), .A2(n12581), .ZN(n8161) );
  AND2_X1 U10656 ( .A1(n11682), .A2(n8945), .ZN(n11837) );
  INV_X1 U10657 ( .A(n11841), .ZN(n8221) );
  INV_X1 U10658 ( .A(n8946), .ZN(n8164) );
  INV_X2 U10659 ( .A(n8226), .ZN(n11795) );
  NAND2_X1 U10660 ( .A1(n7131), .A2(n7134), .ZN(n9627) );
  AND2_X1 U10661 ( .A1(n9625), .A2(n9627), .ZN(n8175) );
  NAND2_X1 U10662 ( .A1(n8166), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8174) );
  INV_X1 U10663 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8943) );
  OR2_X1 U10664 ( .A1(n8167), .A2(n8943), .ZN(n8173) );
  INV_X1 U10665 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8168) );
  NOR2_X1 U10666 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  OR2_X1 U10667 ( .A1(n8072), .A2(n12688), .ZN(n8172) );
  INV_X1 U10668 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8953) );
  OR2_X1 U10669 ( .A1(n6570), .A2(n8953), .ZN(n8171) );
  AND4_X2 U10670 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .ZN(n9304)
         );
  INV_X1 U10671 ( .A(n9304), .ZN(n12579) );
  AOI22_X1 U10672 ( .A1(n8165), .A2(n12579), .B1(n12581), .B2(n12849), .ZN(
        n9408) );
  AOI21_X1 U10673 ( .B1(n15611), .B2(n12696), .A(n12697), .ZN(n13212) );
  NAND2_X1 U10674 ( .A1(n8215), .A2(n8178), .ZN(n8214) );
  XNOR2_X1 U10675 ( .A(n8194), .B(P3_B_REG_SCAN_IN), .ZN(n8183) );
  INV_X1 U10676 ( .A(n8214), .ZN(n8181) );
  INV_X1 U10677 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8180) );
  OAI21_X1 U10678 ( .B1(n8184), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8186) );
  OR2_X1 U10679 ( .A1(n8186), .A2(n8185), .ZN(n8191) );
  INV_X1 U10680 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8193) );
  INV_X1 U10681 ( .A(n8194), .ZN(n8195) );
  NAND2_X1 U10682 ( .A1(n13285), .A2(n8195), .ZN(n8196) );
  INV_X1 U10683 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10684 ( .A1(n9899), .A2(n8197), .ZN(n8201) );
  INV_X1 U10685 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10686 ( .A1(n13285), .A2(n8199), .ZN(n8200) );
  XNOR2_X1 U10687 ( .A(n9319), .B(n13265), .ZN(n8220) );
  NOR2_X1 U10688 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .ZN(
        n8205) );
  NOR4_X1 U10689 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8204) );
  NOR4_X1 U10690 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8203) );
  NOR4_X1 U10691 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8202) );
  NAND4_X1 U10692 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n8211)
         );
  NOR4_X1 U10693 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8209) );
  NOR4_X1 U10694 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8208) );
  NOR4_X1 U10695 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8207) );
  NOR4_X1 U10696 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8206) );
  NAND4_X1 U10697 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8210)
         );
  INV_X1 U10698 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U10699 ( .A1(n8216), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8217) );
  MUX2_X1 U10700 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8217), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8218) );
  NAND2_X1 U10701 ( .A1(n8947), .A2(n11839), .ZN(n8219) );
  NAND2_X1 U10702 ( .A1(n8222), .A2(n8221), .ZN(n8225) );
  NAND2_X1 U10703 ( .A1(n11834), .A2(n8946), .ZN(n8223) );
  NAND2_X1 U10704 ( .A1(n10789), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U10705 ( .A1(n8225), .A2(n8224), .ZN(n8230) );
  NAND2_X1 U10706 ( .A1(n8226), .A2(n8227), .ZN(n10308) );
  NAND2_X1 U10707 ( .A1(n10310), .A2(n10308), .ZN(n8228) );
  NAND2_X1 U10708 ( .A1(n13265), .A2(n8228), .ZN(n8229) );
  OAI21_X1 U10709 ( .B1(n13265), .B2(n8230), .A(n8229), .ZN(n8231) );
  INV_X1 U10710 ( .A(n8231), .ZN(n8232) );
  MUX2_X1 U10711 ( .A(n8233), .B(n13212), .S(n15631), .Z(n8234) );
  NAND2_X1 U10712 ( .A1(n8234), .A2(n7645), .ZN(P3_U3486) );
  NOR2_X2 U10713 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n8243) );
  NAND2_X1 U10714 ( .A1(n8572), .A2(n8243), .ZN(n8605) );
  NOR2_X1 U10715 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8237) );
  NAND2_X1 U10716 ( .A1(n8653), .A2(n8237), .ZN(n8677) );
  NOR2_X1 U10717 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8241) );
  NAND4_X1 U10718 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n8245)
         );
  NAND3_X1 U10719 ( .A1(n8243), .A2(n8242), .A3(n8674), .ZN(n8244) );
  NAND2_X1 U10720 ( .A1(n6588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8247) );
  MUX2_X1 U10721 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8247), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8249) );
  INV_X1 U10722 ( .A(n8259), .ZN(n8248) );
  NAND2_X1 U10723 ( .A1(n13565), .A2(n10920), .ZN(n10181) );
  NAND2_X1 U10724 ( .A1(n8250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U10725 ( .A1(n10181), .A2(n10173), .ZN(n10177) );
  NAND4_X1 U10726 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8275), .ZN(n8258)
         );
  NAND2_X1 U10727 ( .A1(n8267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8263) );
  MUX2_X1 U10728 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8263), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8264) );
  NAND2_X1 U10729 ( .A1(n8265), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8266) );
  MUX2_X1 U10730 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8266), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8268) );
  NAND2_X1 U10731 ( .A1(n8268), .A2(n8267), .ZN(n14020) );
  NAND2_X1 U10732 ( .A1(n8270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8271) );
  MUX2_X1 U10733 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8271), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8272) );
  NAND2_X1 U10734 ( .A1(n8272), .A2(n8265), .ZN(n11619) );
  NOR2_X1 U10735 ( .A1(n14020), .A2(n11619), .ZN(n8273) );
  NAND2_X1 U10736 ( .A1(n8288), .A2(n8273), .ZN(n9592) );
  NOR4_X1 U10737 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8285) );
  INV_X1 U10738 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15331) );
  INV_X1 U10739 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15334) );
  INV_X1 U10740 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15355) );
  INV_X1 U10741 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15338) );
  NAND4_X1 U10742 ( .A1(n15331), .A2(n15334), .A3(n15355), .A4(n15338), .ZN(
        n8282) );
  NOR4_X1 U10743 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8280) );
  NOR4_X1 U10744 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8279) );
  NOR4_X1 U10745 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n8278) );
  NOR4_X1 U10746 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8277) );
  NAND4_X1 U10747 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), .ZN(n8281)
         );
  NOR4_X1 U10748 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n8282), .A4(n8281), .ZN(n8284) );
  NOR4_X1 U10749 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8283) );
  NAND3_X1 U10750 ( .A1(n8285), .A2(n8284), .A3(n8283), .ZN(n8289) );
  XNOR2_X1 U10751 ( .A(n11619), .B(P2_B_REG_SCAN_IN), .ZN(n8286) );
  NAND2_X1 U10752 ( .A1(n14020), .A2(n8286), .ZN(n8287) );
  NAND2_X1 U10753 ( .A1(n8289), .A2(n15330), .ZN(n10171) );
  INV_X1 U10754 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U10755 ( .A1(n15330), .A2(n15362), .ZN(n8291) );
  NAND2_X1 U10756 ( .A1(n14019), .A2(n11619), .ZN(n8290) );
  NAND2_X1 U10757 ( .A1(n8291), .A2(n8290), .ZN(n15363) );
  AND3_X1 U10758 ( .A1(n15367), .A2(n10171), .A3(n15363), .ZN(n8292) );
  AND2_X1 U10759 ( .A1(n10177), .A2(n8292), .ZN(n10645) );
  INV_X1 U10760 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15365) );
  NAND2_X1 U10761 ( .A1(n15330), .A2(n15365), .ZN(n8294) );
  NAND2_X1 U10762 ( .A1(n14019), .A2(n14020), .ZN(n8293) );
  NAND2_X1 U10763 ( .A1(n15442), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U10764 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8487) );
  INV_X1 U10765 ( .A(n8487), .ZN(n8295) );
  NAND2_X1 U10766 ( .A1(n8295), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8512) );
  INV_X1 U10767 ( .A(n8512), .ZN(n8296) );
  NAND2_X1 U10768 ( .A1(n8296), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8529) );
  INV_X1 U10769 ( .A(n8576), .ZN(n8297) );
  NAND2_X1 U10770 ( .A1(n8297), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8596) );
  INV_X1 U10771 ( .A(n8611), .ZN(n8298) );
  NAND2_X1 U10772 ( .A1(n8298), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8630) );
  INV_X1 U10773 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8629) );
  INV_X1 U10774 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10775 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n8300) );
  INV_X1 U10776 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8727) );
  INV_X1 U10777 ( .A(n8772), .ZN(n8302) );
  NAND2_X1 U10778 ( .A1(n8302), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8788) );
  INV_X1 U10779 ( .A(n8804), .ZN(n8303) );
  NAND2_X1 U10780 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8304) );
  INV_X1 U10781 ( .A(n8844), .ZN(n8305) );
  NAND2_X1 U10782 ( .A1(n8305), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8846) );
  INV_X1 U10783 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10784 ( .A1(n8846), .A2(n8306), .ZN(n8307) );
  XNOR2_X2 U10785 ( .A(n8308), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8313) );
  NOR2_X1 U10786 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .ZN(n8309) );
  NAND2_X1 U10787 ( .A1(n8413), .A2(n8309), .ZN(n14002) );
  INV_X1 U10788 ( .A(n8312), .ZN(n8311) );
  NAND2_X1 U10789 ( .A1(n13593), .A2(n6577), .ZN(n8319) );
  INV_X1 U10790 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10791 ( .A1(n9159), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10792 ( .A1(n8859), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8314) );
  OAI211_X1 U10793 ( .C1(n8316), .C2(n8430), .A(n8315), .B(n8314), .ZN(n8317)
         );
  INV_X1 U10794 ( .A(n8317), .ZN(n8318) );
  INV_X1 U10795 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9710) );
  AND2_X1 U10796 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8320) );
  NAND2_X1 U10797 ( .A1(n9681), .A2(n8320), .ZN(n9476) );
  AND2_X1 U10798 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10799 ( .A1(n8324), .A2(n8321), .ZN(n8425) );
  NAND2_X1 U10800 ( .A1(n9476), .A2(n8425), .ZN(n8442) );
  INV_X1 U10801 ( .A(SI_1_), .ZN(n9667) );
  NOR2_X1 U10802 ( .A1(n8322), .A2(n9667), .ZN(n8323) );
  MUX2_X1 U10803 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8324), .Z(n8325) );
  XNOR2_X1 U10804 ( .A(n8325), .B(SI_2_), .ZN(n8457) );
  NAND2_X1 U10805 ( .A1(n8325), .A2(SI_2_), .ZN(n8326) );
  MUX2_X1 U10806 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8324), .Z(n8327) );
  XNOR2_X1 U10807 ( .A(n8327), .B(n9672), .ZN(n8468) );
  NAND2_X1 U10808 ( .A1(n8327), .A2(SI_3_), .ZN(n8328) );
  NAND2_X1 U10809 ( .A1(n8329), .A2(n8328), .ZN(n8481) );
  MUX2_X1 U10810 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8324), .Z(n8331) );
  XNOR2_X1 U10811 ( .A(n8331), .B(n8330), .ZN(n8482) );
  NAND2_X1 U10812 ( .A1(n8481), .A2(n8482), .ZN(n8333) );
  NAND2_X1 U10813 ( .A1(n8331), .A2(SI_4_), .ZN(n8332) );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n11919), .Z(n8335) );
  XNOR2_X1 U10815 ( .A(n8335), .B(SI_5_), .ZN(n8495) );
  INV_X1 U10816 ( .A(n8495), .ZN(n8334) );
  NAND2_X1 U10817 ( .A1(n8335), .A2(SI_5_), .ZN(n8336) );
  MUX2_X1 U10818 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11919), .Z(n8338) );
  XNOR2_X1 U10819 ( .A(n8338), .B(SI_6_), .ZN(n8502) );
  INV_X1 U10820 ( .A(n8502), .ZN(n8337) );
  NAND2_X1 U10821 ( .A1(n8338), .A2(SI_6_), .ZN(n8339) );
  NAND2_X1 U10822 ( .A1(n8340), .A2(n8339), .ZN(n8520) );
  NAND2_X1 U10823 ( .A1(n8342), .A2(SI_7_), .ZN(n8343) );
  MUX2_X1 U10824 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11919), .Z(n8344) );
  MUX2_X1 U10825 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9680), .Z(n8346) );
  XNOR2_X1 U10826 ( .A(n8346), .B(SI_9_), .ZN(n8553) );
  INV_X1 U10827 ( .A(n8553), .ZN(n8345) );
  NAND2_X1 U10828 ( .A1(n8346), .A2(SI_9_), .ZN(n8347) );
  MUX2_X1 U10829 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9680), .Z(n8569) );
  INV_X1 U10830 ( .A(n8569), .ZN(n8348) );
  NAND2_X1 U10831 ( .A1(n8348), .A2(n9668), .ZN(n8349) );
  MUX2_X1 U10832 ( .A(n9758), .B(n9753), .S(n9680), .Z(n8351) );
  NAND2_X1 U10833 ( .A1(n8351), .A2(n8350), .ZN(n8354) );
  INV_X1 U10834 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U10835 ( .A1(n8352), .A2(SI_11_), .ZN(n8353) );
  NAND2_X1 U10836 ( .A1(n8354), .A2(n8353), .ZN(n8586) );
  MUX2_X1 U10837 ( .A(n7693), .B(n10004), .S(n9680), .Z(n8355) );
  NAND2_X1 U10838 ( .A1(n8355), .A2(n9689), .ZN(n8619) );
  INV_X1 U10839 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U10840 ( .A1(n8356), .A2(SI_12_), .ZN(n8357) );
  MUX2_X1 U10841 ( .A(n11167), .B(n10027), .S(n9680), .Z(n8358) );
  NAND2_X1 U10842 ( .A1(n8358), .A2(n9745), .ZN(n8622) );
  AND2_X1 U10843 ( .A1(n8619), .A2(n8622), .ZN(n8361) );
  INV_X1 U10844 ( .A(n8358), .ZN(n8359) );
  NAND2_X1 U10845 ( .A1(n8359), .A2(SI_13_), .ZN(n8621) );
  MUX2_X1 U10846 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9680), .Z(n8638) );
  MUX2_X1 U10847 ( .A(n6832), .B(n10277), .S(n9680), .Z(n8363) );
  NAND2_X1 U10848 ( .A1(n8363), .A2(n9873), .ZN(n8668) );
  INV_X1 U10849 ( .A(n8363), .ZN(n8364) );
  NAND2_X1 U10850 ( .A1(n8364), .A2(SI_15_), .ZN(n8365) );
  MUX2_X1 U10851 ( .A(n10306), .B(n10360), .S(n9680), .Z(n8366) );
  NAND2_X1 U10852 ( .A1(n8366), .A2(n10001), .ZN(n8671) );
  INV_X1 U10853 ( .A(n8366), .ZN(n8367) );
  NAND2_X1 U10854 ( .A1(n8367), .A2(SI_16_), .ZN(n8670) );
  MUX2_X1 U10855 ( .A(n6851), .B(n13072), .S(n11919), .Z(n8687) );
  NAND2_X1 U10856 ( .A1(n8689), .A2(n8370), .ZN(n8371) );
  NAND2_X1 U10857 ( .A1(n8372), .A2(n8371), .ZN(n8705) );
  MUX2_X1 U10858 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9680), .Z(n8718) );
  NOR2_X1 U10859 ( .A1(n8718), .A2(SI_18_), .ZN(n8375) );
  MUX2_X1 U10860 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9680), .Z(n8376) );
  XNOR2_X1 U10861 ( .A(n8376), .B(SI_19_), .ZN(n8722) );
  INV_X1 U10862 ( .A(n8722), .ZN(n8374) );
  NAND2_X1 U10863 ( .A1(n8718), .A2(SI_18_), .ZN(n8373) );
  INV_X1 U10864 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U10865 ( .A1(n8377), .A2(n10158), .ZN(n8378) );
  MUX2_X1 U10866 ( .A(n10872), .B(n10921), .S(n9680), .Z(n8736) );
  MUX2_X1 U10867 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11919), .Z(n8383) );
  NAND2_X1 U10868 ( .A1(n8383), .A2(SI_21_), .ZN(n8385) );
  OAI21_X1 U10869 ( .B1(SI_21_), .B2(n8383), .A(n8385), .ZN(n8384) );
  INV_X1 U10870 ( .A(n8384), .ZN(n8751) );
  MUX2_X1 U10871 ( .A(n10084), .B(n11320), .S(n9680), .Z(n8766) );
  MUX2_X1 U10872 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11919), .Z(n8783) );
  INV_X1 U10873 ( .A(SI_23_), .ZN(n11090) );
  NAND2_X1 U10874 ( .A1(n8388), .A2(n11090), .ZN(n8389) );
  INV_X1 U10875 ( .A(SI_24_), .ZN(n8391) );
  OR2_X2 U10876 ( .A1(n8392), .A2(n8391), .ZN(n8395) );
  NAND2_X1 U10877 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  INV_X1 U10878 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11616) );
  MUX2_X1 U10879 ( .A(n11616), .B(n11618), .S(n9680), .Z(n8798) );
  INV_X1 U10880 ( .A(n8798), .ZN(n8394) );
  MUX2_X1 U10881 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11919), .Z(n8396) );
  XNOR2_X1 U10882 ( .A(n8396), .B(SI_25_), .ZN(n8812) );
  INV_X1 U10883 ( .A(n8396), .ZN(n8398) );
  INV_X1 U10884 ( .A(SI_25_), .ZN(n8397) );
  MUX2_X1 U10885 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n11919), .Z(n8399) );
  NAND2_X1 U10886 ( .A1(n8399), .A2(SI_26_), .ZN(n8401) );
  OAI21_X1 U10887 ( .B1(SI_26_), .B2(n8399), .A(n8401), .ZN(n8822) );
  INV_X1 U10888 ( .A(n8822), .ZN(n8400) );
  MUX2_X1 U10889 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9680), .Z(n8839) );
  INV_X1 U10890 ( .A(n8839), .ZN(n8402) );
  INV_X1 U10891 ( .A(SI_27_), .ZN(n13277) );
  NAND2_X1 U10892 ( .A1(n8402), .A2(n13277), .ZN(n8403) );
  NAND2_X1 U10893 ( .A1(n8839), .A2(SI_27_), .ZN(n8404) );
  MUX2_X1 U10894 ( .A(n11868), .B(n14012), .S(n11919), .Z(n8405) );
  INV_X1 U10895 ( .A(SI_28_), .ZN(n12300) );
  NAND2_X1 U10896 ( .A1(n8405), .A2(n12300), .ZN(n8856) );
  INV_X1 U10897 ( .A(n8405), .ZN(n8406) );
  NAND2_X1 U10898 ( .A1(n8406), .A2(SI_28_), .ZN(n8407) );
  NAND2_X1 U10899 ( .A1(n8856), .A2(n8407), .ZN(n8854) );
  NAND2_X1 U10900 ( .A1(n8408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10901 ( .A1(n14009), .A2(n9188), .ZN(n8417) );
  OR2_X1 U10902 ( .A1(n8740), .A2(n14012), .ZN(n8416) );
  INV_X1 U10903 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10722) );
  OR2_X1 U10904 ( .A1(n8432), .A2(n10722), .ZN(n8422) );
  NAND2_X1 U10905 ( .A1(n8428), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8421) );
  INV_X1 U10906 ( .A(n8429), .ZN(n8418) );
  NAND2_X1 U10907 ( .A1(n8418), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8420) );
  INV_X1 U10908 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10723) );
  OR2_X1 U10909 ( .A1(n6591), .A2(n10723), .ZN(n8419) );
  NAND4_X2 U10910 ( .A1(n8421), .A2(n8422), .A3(n8420), .A4(n8419), .ZN(n8959)
         );
  INV_X1 U10911 ( .A(n8959), .ZN(n8427) );
  NAND2_X1 U10912 ( .A1(n9680), .A2(SI_0_), .ZN(n8424) );
  NAND2_X1 U10913 ( .A1(n8424), .A2(n8423), .ZN(n8426) );
  NAND2_X1 U10914 ( .A1(n8426), .A2(n8425), .ZN(n14025) );
  INV_X1 U10915 ( .A(n10721), .ZN(n8876) );
  NAND2_X1 U10916 ( .A1(n8427), .A2(n8876), .ZN(n10249) );
  INV_X1 U10917 ( .A(n10249), .ZN(n8444) );
  NAND2_X1 U10918 ( .A1(n8428), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8436) );
  INV_X1 U10919 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9831) );
  OR2_X1 U10920 ( .A1(n8429), .A2(n9831), .ZN(n8435) );
  INV_X1 U10921 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9846) );
  OR2_X1 U10922 ( .A1(n8430), .A2(n9846), .ZN(n8434) );
  INV_X1 U10923 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8431) );
  OR2_X1 U10924 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  NAND4_X2 U10925 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n13515) );
  NAND2_X1 U10926 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8438) );
  MUX2_X1 U10927 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8438), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8441) );
  INV_X1 U10928 ( .A(n8439), .ZN(n8440) );
  XNOR2_X1 U10929 ( .A(n8443), .B(n8442), .ZN(n9709) );
  NAND2_X1 U10930 ( .A1(n8444), .A2(n6573), .ZN(n8446) );
  INV_X1 U10931 ( .A(n13515), .ZN(n10270) );
  NAND2_X1 U10932 ( .A1(n10270), .A2(n8968), .ZN(n8445) );
  NAND2_X1 U10933 ( .A1(n8428), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8451) );
  INV_X1 U10934 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10234) );
  OR2_X1 U10935 ( .A1(n8432), .A2(n10234), .ZN(n8450) );
  INV_X1 U10936 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9833) );
  OR2_X1 U10937 ( .A1(n8429), .A2(n9833), .ZN(n8449) );
  INV_X1 U10938 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8447) );
  OR2_X1 U10939 ( .A1(n8430), .A2(n8447), .ZN(n8448) );
  NOR2_X1 U10940 ( .A1(n8439), .A2(n8412), .ZN(n8452) );
  MUX2_X1 U10941 ( .A(n8412), .B(n8452), .S(P2_IR_REG_2__SCAN_IN), .Z(n8453)
         );
  INV_X1 U10942 ( .A(n8453), .ZN(n8456) );
  INV_X1 U10943 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U10944 ( .A1(n8456), .A2(n8455), .ZN(n9878) );
  OR2_X1 U10945 ( .A1(n8740), .A2(n9661), .ZN(n8460) );
  XNOR2_X1 U10946 ( .A(n8458), .B(n8457), .ZN(n9707) );
  NAND2_X1 U10947 ( .A1(n6854), .A2(n15318), .ZN(n8461) );
  NAND2_X1 U10948 ( .A1(n8859), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8466) );
  OR2_X1 U10949 ( .A1(n8613), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8465) );
  INV_X1 U10950 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10711) );
  OR2_X1 U10951 ( .A1(n8430), .A2(n10711), .ZN(n8464) );
  INV_X1 U10952 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9834) );
  OR2_X1 U10953 ( .A1(n6593), .A2(n9834), .ZN(n8463) );
  OR2_X1 U10954 ( .A1(n8454), .A2(n8412), .ZN(n8467) );
  XNOR2_X1 U10955 ( .A(n8469), .B(n8468), .ZN(n9702) );
  OR2_X1 U10956 ( .A1(n8802), .A2(n9702), .ZN(n8470) );
  INV_X1 U10957 ( .A(n9238), .ZN(n10162) );
  NAND2_X1 U10958 ( .A1(n10163), .A2(n10162), .ZN(n8473) );
  INV_X1 U10959 ( .A(n13513), .ZN(n10402) );
  NAND2_X1 U10960 ( .A1(n10402), .A2(n15224), .ZN(n8472) );
  NAND2_X1 U10961 ( .A1(n8859), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8477) );
  INV_X1 U10962 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9837) );
  OR2_X1 U10963 ( .A1(n6593), .A2(n9837), .ZN(n8476) );
  OAI21_X1 U10964 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8487), .ZN(n10705) );
  OR2_X1 U10965 ( .A1(n8613), .A2(n10705), .ZN(n8475) );
  INV_X1 U10966 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10700) );
  OR2_X1 U10967 ( .A1(n8430), .A2(n10700), .ZN(n8474) );
  NAND4_X1 U10968 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n13512) );
  NAND2_X1 U10969 ( .A1(n8454), .A2(n8478), .ZN(n8493) );
  NAND2_X1 U10970 ( .A1(n8493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U10971 ( .A(n8480), .B(n8479), .ZN(n9955) );
  OR2_X1 U10972 ( .A1(n8740), .A2(n9662), .ZN(n8484) );
  XNOR2_X1 U10973 ( .A(n8481), .B(n8482), .ZN(n9683) );
  OR2_X1 U10974 ( .A1(n8802), .A2(n9683), .ZN(n8483) );
  INV_X1 U10975 ( .A(n15383), .ZN(n10706) );
  NAND2_X1 U10976 ( .A1(n6814), .A2(n15383), .ZN(n8485) );
  NAND2_X1 U10977 ( .A1(n8859), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8492) );
  INV_X1 U10978 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10655) );
  OR2_X1 U10979 ( .A1(n8430), .A2(n10655), .ZN(n8491) );
  INV_X1 U10980 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10981 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  NAND2_X1 U10982 ( .A1(n8512), .A2(n8488), .ZN(n11856) );
  OR2_X1 U10983 ( .A1(n8613), .A2(n11856), .ZN(n8490) );
  INV_X1 U10984 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9838) );
  OR2_X1 U10985 ( .A1(n6593), .A2(n9838), .ZN(n8489) );
  NAND4_X1 U10986 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n13511) );
  NAND2_X1 U10987 ( .A1(n8503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8494) );
  XNOR2_X1 U10988 ( .A(n8494), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10989 ( .A1(n8724), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6771), .B2(
        n9851), .ZN(n8498) );
  XNOR2_X1 U10990 ( .A(n8495), .B(n8496), .ZN(n9685) );
  NAND2_X1 U10991 ( .A1(n9685), .A2(n9188), .ZN(n8497) );
  NAND2_X1 U10992 ( .A1(n8498), .A2(n8497), .ZN(n15390) );
  XNOR2_X1 U10993 ( .A(n13511), .B(n15390), .ZN(n10650) );
  INV_X1 U10994 ( .A(n13511), .ZN(n8884) );
  NAND2_X1 U10995 ( .A1(n8884), .A2(n15390), .ZN(n8499) );
  NAND2_X1 U10996 ( .A1(n8500), .A2(n8499), .ZN(n10680) );
  XNOR2_X1 U10997 ( .A(n8501), .B(n8502), .ZN(n10460) );
  NAND2_X1 U10998 ( .A1(n10460), .A2(n9188), .ZN(n8510) );
  INV_X1 U10999 ( .A(n8503), .ZN(n8505) );
  INV_X1 U11000 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U11001 ( .A1(n8505), .A2(n8504), .ZN(n8538) );
  NAND2_X1 U11002 ( .A1(n8538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8507) );
  INV_X1 U11003 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U11004 ( .A1(n8507), .A2(n8506), .ZN(n8523) );
  OR2_X1 U11005 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  AOI22_X1 U11006 ( .A1(n8724), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6771), .B2(
        n9852), .ZN(n8509) );
  NAND2_X1 U11007 ( .A1(n8859), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8517) );
  INV_X1 U11008 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9839) );
  OR2_X1 U11009 ( .A1(n6593), .A2(n9839), .ZN(n8516) );
  INV_X1 U11010 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U11011 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  NAND2_X1 U11012 ( .A1(n8529), .A2(n8513), .ZN(n10690) );
  OR2_X1 U11013 ( .A1(n8613), .A2(n10690), .ZN(n8515) );
  INV_X1 U11014 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10685) );
  OR2_X1 U11015 ( .A1(n8430), .A2(n10685), .ZN(n8514) );
  NAND4_X1 U11016 ( .A1(n8517), .A2(n8516), .A3(n8515), .A4(n8514), .ZN(n13510) );
  XNOR2_X1 U11017 ( .A(n15396), .B(n13510), .ZN(n10679) );
  NAND2_X1 U11018 ( .A1(n10680), .A2(n10679), .ZN(n8519) );
  INV_X1 U11019 ( .A(n13510), .ZN(n10573) );
  NAND2_X1 U11020 ( .A1(n10573), .A2(n15396), .ZN(n8518) );
  XNOR2_X1 U11021 ( .A(n8522), .B(n8521), .ZN(n10490) );
  NAND2_X1 U11022 ( .A1(n10490), .A2(n9188), .ZN(n8526) );
  NAND2_X1 U11023 ( .A1(n8523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8524) );
  XNOR2_X1 U11024 ( .A(n8524), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U11025 ( .A1(n8724), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6771), .B2(
        n9895), .ZN(n8525) );
  NAND2_X1 U11026 ( .A1(n8526), .A2(n8525), .ZN(n15404) );
  NAND2_X1 U11027 ( .A1(n8859), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8534) );
  INV_X1 U11028 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8527) );
  OR2_X1 U11029 ( .A1(n6593), .A2(n8527), .ZN(n8533) );
  NAND2_X1 U11030 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U11031 ( .A1(n8543), .A2(n8530), .ZN(n10670) );
  OR2_X1 U11032 ( .A1(n8613), .A2(n10670), .ZN(n8532) );
  INV_X1 U11033 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10668) );
  OR2_X1 U11034 ( .A1(n8430), .A2(n10668), .ZN(n8531) );
  NAND4_X1 U11035 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n13509) );
  INV_X1 U11036 ( .A(n13509), .ZN(n13875) );
  AND2_X1 U11037 ( .A1(n15404), .A2(n13875), .ZN(n8535) );
  XNOR2_X1 U11038 ( .A(n8536), .B(n8537), .ZN(n10495) );
  NAND2_X1 U11039 ( .A1(n10495), .A2(n9188), .ZN(n8541) );
  NAND2_X1 U11040 ( .A1(n8555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U11041 ( .A(n8539), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U11042 ( .A1(n8724), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6771), .B2(
        n9853), .ZN(n8540) );
  NAND2_X1 U11043 ( .A1(n8859), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8549) );
  INV_X1 U11044 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n13882) );
  OR2_X1 U11045 ( .A1(n8430), .A2(n13882), .ZN(n8548) );
  NAND2_X1 U11046 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U11047 ( .A1(n8561), .A2(n8544), .ZN(n13881) );
  OR2_X1 U11048 ( .A1(n8613), .A2(n13881), .ZN(n8547) );
  INV_X1 U11049 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8545) );
  OR2_X1 U11050 ( .A1(n6593), .A2(n8545), .ZN(n8546) );
  NAND4_X1 U11051 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n13853) );
  XNOR2_X1 U11052 ( .A(n13889), .B(n11873), .ZN(n13870) );
  NAND2_X1 U11053 ( .A1(n13871), .A2(n13868), .ZN(n8551) );
  OR2_X1 U11054 ( .A1(n13889), .A2(n11873), .ZN(n8550) );
  NAND2_X1 U11055 ( .A1(n8551), .A2(n8550), .ZN(n13856) );
  XNOR2_X1 U11056 ( .A(n8554), .B(n8553), .ZN(n10800) );
  NAND2_X1 U11057 ( .A1(n10800), .A2(n9188), .ZN(n8558) );
  OAI21_X1 U11058 ( .B1(n8555), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8556) );
  XNOR2_X1 U11059 ( .A(n8556), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11060 ( .A1(n8724), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6771), .B2(
        n10012), .ZN(n8557) );
  NAND2_X1 U11061 ( .A1(n9159), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8566) );
  INV_X1 U11062 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8559) );
  OR2_X1 U11063 ( .A1(n9162), .A2(n8559), .ZN(n8565) );
  NAND2_X1 U11064 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U11065 ( .A1(n8576), .A2(n8562), .ZN(n13860) );
  OR2_X1 U11066 ( .A1(n8613), .A2(n13860), .ZN(n8564) );
  INV_X1 U11067 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13861) );
  OR2_X1 U11068 ( .A1(n8430), .A2(n13861), .ZN(n8563) );
  NAND4_X1 U11069 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n13508) );
  XNOR2_X1 U11070 ( .A(n13865), .B(n13508), .ZN(n9243) );
  NAND2_X1 U11071 ( .A1(n13856), .A2(n9243), .ZN(n8568) );
  INV_X1 U11072 ( .A(n13508), .ZN(n13873) );
  OR2_X1 U11073 ( .A1(n13865), .A2(n13873), .ZN(n8567) );
  XNOR2_X1 U11074 ( .A(n8569), .B(SI_10_), .ZN(n8570) );
  XNOR2_X1 U11075 ( .A(n8571), .B(n8570), .ZN(n10806) );
  NAND2_X1 U11076 ( .A1(n10806), .A2(n9188), .ZN(n8574) );
  OR2_X1 U11077 ( .A1(n8572), .A2(n8412), .ZN(n8590) );
  XNOR2_X1 U11078 ( .A(n8590), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U11079 ( .A1(n8724), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6771), 
        .B2(n11005), .ZN(n8573) );
  NAND2_X1 U11080 ( .A1(n8859), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8582) );
  INV_X1 U11081 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n13840) );
  OR2_X1 U11082 ( .A1(n8430), .A2(n13840), .ZN(n8581) );
  INV_X1 U11083 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U11084 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  NAND2_X1 U11085 ( .A1(n8596), .A2(n8577), .ZN(n13839) );
  OR2_X1 U11086 ( .A1(n8613), .A2(n13839), .ZN(n8580) );
  INV_X1 U11087 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8578) );
  OR2_X1 U11088 ( .A1(n6593), .A2(n8578), .ZN(n8579) );
  NAND4_X1 U11089 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n13852) );
  XNOR2_X1 U11090 ( .A(n13845), .B(n13852), .ZN(n9244) );
  INV_X1 U11091 ( .A(n13852), .ZN(n11287) );
  OR2_X1 U11092 ( .A1(n13845), .A2(n11287), .ZN(n8583) );
  NAND2_X1 U11093 ( .A1(n8585), .A2(n8586), .ZN(n8587) );
  NAND2_X1 U11094 ( .A1(n8588), .A2(n8587), .ZN(n10953) );
  NAND2_X1 U11095 ( .A1(n10953), .A2(n9188), .ZN(n8594) );
  INV_X1 U11096 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U11097 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  NAND2_X1 U11098 ( .A1(n8591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8592) );
  XNOR2_X1 U11099 ( .A(n8592), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U11100 ( .A1(n8724), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6771), 
        .B2(n11019), .ZN(n8593) );
  NAND2_X1 U11101 ( .A1(n8859), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8601) );
  INV_X1 U11102 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13824) );
  OR2_X1 U11103 ( .A1(n8430), .A2(n13824), .ZN(n8600) );
  NAND2_X1 U11104 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  NAND2_X1 U11105 ( .A1(n8611), .A2(n8597), .ZN(n13823) );
  OR2_X1 U11106 ( .A1(n8613), .A2(n13823), .ZN(n8599) );
  INV_X1 U11107 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11020) );
  OR2_X1 U11108 ( .A1(n6593), .A2(n11020), .ZN(n8598) );
  NAND4_X1 U11109 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n13798) );
  XNOR2_X1 U11110 ( .A(n15435), .B(n13798), .ZN(n9246) );
  INV_X1 U11111 ( .A(n13798), .ZN(n13835) );
  NAND2_X1 U11112 ( .A1(n15435), .A2(n13835), .ZN(n8602) );
  XNOR2_X1 U11113 ( .A(n8604), .B(n8603), .ZN(n11161) );
  NAND2_X1 U11114 ( .A1(n11161), .A2(n9188), .ZN(n8608) );
  NAND2_X1 U11115 ( .A1(n8605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U11116 ( .A(n8606), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15268) );
  AOI22_X1 U11117 ( .A1(n8724), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6771), 
        .B2(n15268), .ZN(n8607) );
  NAND2_X1 U11118 ( .A1(n9159), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8617) );
  INV_X1 U11119 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8609) );
  OR2_X1 U11120 ( .A1(n9162), .A2(n8609), .ZN(n8616) );
  INV_X1 U11121 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U11122 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  NAND2_X1 U11123 ( .A1(n8630), .A2(n8612), .ZN(n13803) );
  OR2_X1 U11124 ( .A1(n8613), .A2(n13803), .ZN(n8615) );
  INV_X1 U11125 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13804) );
  OR2_X1 U11126 ( .A1(n8430), .A2(n13804), .ZN(n8614) );
  NAND4_X1 U11127 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n13814) );
  INV_X1 U11128 ( .A(n13814), .ZN(n9050) );
  XNOR2_X1 U11129 ( .A(n13808), .B(n9050), .ZN(n13799) );
  OR2_X1 U11130 ( .A1(n13808), .A2(n9050), .ZN(n8618) );
  NAND2_X1 U11131 ( .A1(n8620), .A2(n8619), .ZN(n8624) );
  AND2_X1 U11132 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  XNOR2_X1 U11133 ( .A(n8624), .B(n8623), .ZN(n11166) );
  NAND2_X1 U11134 ( .A1(n11166), .A2(n9188), .ZN(n8628) );
  NAND2_X1 U11135 ( .A1(n6616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8625) );
  XNOR2_X1 U11136 ( .A(n8625), .B(n7354), .ZN(n15273) );
  INV_X1 U11137 ( .A(n15273), .ZN(n8626) );
  AOI22_X1 U11138 ( .A1(n8724), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6771), 
        .B2(n8626), .ZN(n8627) );
  NAND2_X1 U11139 ( .A1(n8859), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8635) );
  INV_X1 U11140 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11023) );
  OR2_X1 U11141 ( .A1(n6593), .A2(n11023), .ZN(n8634) );
  NAND2_X1 U11142 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND2_X1 U11143 ( .A1(n8645), .A2(n8631), .ZN(n11377) );
  OR2_X1 U11144 ( .A1(n8613), .A2(n11377), .ZN(n8633) );
  INV_X1 U11145 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11002) );
  OR2_X1 U11146 ( .A1(n8430), .A2(n11002), .ZN(n8632) );
  NAND4_X1 U11147 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n13797) );
  INV_X1 U11148 ( .A(n13797), .ZN(n11239) );
  XNOR2_X1 U11149 ( .A(n11454), .B(n11239), .ZN(n11381) );
  INV_X1 U11150 ( .A(n11381), .ZN(n8636) );
  OR2_X1 U11151 ( .A1(n11454), .A2(n11239), .ZN(n8637) );
  XNOR2_X1 U11152 ( .A(n8639), .B(n8638), .ZN(n11358) );
  NAND2_X1 U11153 ( .A1(n11358), .A2(n9188), .ZN(n8643) );
  OR2_X1 U11154 ( .A1(n8640), .A2(n8412), .ZN(n8641) );
  XNOR2_X1 U11155 ( .A(n8641), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U11156 ( .A1(n8724), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6771), 
        .B2(n11006), .ZN(n8642) );
  NAND2_X1 U11157 ( .A1(n8859), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8650) );
  INV_X1 U11158 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11016) );
  OR2_X1 U11159 ( .A1(n6593), .A2(n11016), .ZN(n8649) );
  NAND2_X1 U11160 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U11161 ( .A1(n8657), .A2(n8646), .ZN(n13789) );
  OR2_X1 U11162 ( .A1(n8613), .A2(n13789), .ZN(n8648) );
  INV_X1 U11163 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13790) );
  OR2_X1 U11164 ( .A1(n8430), .A2(n13790), .ZN(n8647) );
  NAND4_X1 U11165 ( .A1(n8650), .A2(n8649), .A3(n8648), .A4(n8647), .ZN(n13506) );
  INV_X1 U11166 ( .A(n13506), .ZN(n11300) );
  NOR2_X1 U11167 ( .A1(n13792), .A2(n11300), .ZN(n8651) );
  XNOR2_X1 U11168 ( .A(n6694), .B(n8652), .ZN(n11432) );
  NAND2_X1 U11169 ( .A1(n11432), .A2(n9188), .ZN(n8656) );
  OR2_X1 U11170 ( .A1(n8653), .A2(n8412), .ZN(n8654) );
  XNOR2_X1 U11171 ( .A(n8654), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U11172 ( .A1(n8724), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6771), 
        .B2(n15299), .ZN(n8655) );
  NAND2_X1 U11173 ( .A1(n8859), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8664) );
  INV_X1 U11174 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U11175 ( .A1(n8657), .A2(n13166), .ZN(n8658) );
  NAND2_X1 U11176 ( .A1(n8696), .A2(n8658), .ZN(n11593) );
  OR2_X1 U11177 ( .A1(n8613), .A2(n11593), .ZN(n8663) );
  INV_X1 U11178 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8659) );
  OR2_X1 U11179 ( .A1(n8430), .A2(n8659), .ZN(n8662) );
  INV_X1 U11180 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8660) );
  OR2_X1 U11181 ( .A1(n6593), .A2(n8660), .ZN(n8661) );
  NAND4_X1 U11182 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n13784) );
  INV_X1 U11183 ( .A(n13784), .ZN(n11498) );
  AND2_X1 U11184 ( .A1(n13981), .A2(n11498), .ZN(n8665) );
  OR2_X1 U11185 ( .A1(n13981), .A2(n11498), .ZN(n8666) );
  NAND2_X2 U11186 ( .A1(n8667), .A2(n8666), .ZN(n13765) );
  NAND2_X1 U11187 ( .A1(n8669), .A2(n8668), .ZN(n8673) );
  AND2_X1 U11188 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U11189 ( .A(n8673), .B(n8672), .ZN(n11526) );
  NAND2_X1 U11190 ( .A1(n11526), .A2(n9188), .ZN(n8680) );
  NAND2_X1 U11191 ( .A1(n8653), .A2(n8674), .ZN(n8675) );
  NAND2_X1 U11192 ( .A1(n8675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8676) );
  MUX2_X1 U11193 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8676), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8678) );
  AND2_X1 U11194 ( .A1(n8678), .A2(n8677), .ZN(n11110) );
  AOI22_X1 U11195 ( .A1(n8724), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6771), 
        .B2(n11110), .ZN(n8679) );
  NAND2_X1 U11196 ( .A1(n9159), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8686) );
  INV_X1 U11197 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8681) );
  OR2_X1 U11198 ( .A1(n9162), .A2(n8681), .ZN(n8685) );
  INV_X1 U11199 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8695) );
  XNOR2_X1 U11200 ( .A(n8696), .B(n8695), .ZN(n13776) );
  OR2_X1 U11201 ( .A1(n8613), .A2(n13776), .ZN(n8684) );
  INV_X1 U11202 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8682) );
  OR2_X1 U11203 ( .A1(n8430), .A2(n8682), .ZN(n8683) );
  NAND4_X1 U11204 ( .A1(n8686), .A2(n8685), .A3(n8684), .A4(n8683), .ZN(n13505) );
  INV_X1 U11205 ( .A(n13505), .ZN(n9077) );
  INV_X1 U11206 ( .A(n13967), .ZN(n13779) );
  XNOR2_X1 U11207 ( .A(n8687), .B(SI_17_), .ZN(n8688) );
  XNOR2_X1 U11208 ( .A(n8689), .B(n8688), .ZN(n12022) );
  NAND2_X1 U11209 ( .A1(n12022), .A2(n9188), .ZN(n8693) );
  NAND2_X1 U11210 ( .A1(n8677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8690) );
  MUX2_X1 U11211 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8690), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8691) );
  NAND2_X1 U11212 ( .A1(n8691), .A2(n6715), .ZN(n13543) );
  INV_X1 U11213 ( .A(n13543), .ZN(n13533) );
  AOI22_X1 U11214 ( .A1(n8724), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6771), 
        .B2(n13533), .ZN(n8692) );
  INV_X1 U11215 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8694) );
  OAI21_X1 U11216 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  NAND2_X1 U11217 ( .A1(n8697), .A2(n8710), .ZN(n13756) );
  OR2_X1 U11218 ( .A1(n13756), .A2(n8613), .ZN(n8703) );
  INV_X1 U11219 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13542) );
  OR2_X1 U11220 ( .A1(n6593), .A2(n13542), .ZN(n8702) );
  INV_X1 U11221 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8698) );
  OR2_X1 U11222 ( .A1(n9162), .A2(n8698), .ZN(n8701) );
  INV_X1 U11223 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8699) );
  OR2_X1 U11224 ( .A1(n8430), .A2(n8699), .ZN(n8700) );
  NAND4_X1 U11225 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n13770) );
  INV_X1 U11226 ( .A(n13770), .ZN(n13475) );
  AND2_X1 U11227 ( .A1(n13962), .A2(n13475), .ZN(n8704) );
  INV_X1 U11228 ( .A(SI_18_), .ZN(n10081) );
  NAND2_X1 U11229 ( .A1(n8705), .A2(n10081), .ZN(n8706) );
  NAND2_X1 U11230 ( .A1(n8719), .A2(n8706), .ZN(n8721) );
  NAND2_X1 U11231 ( .A1(n12052), .A2(n9188), .ZN(n8709) );
  NAND2_X1 U11232 ( .A1(n6715), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U11233 ( .A(n8707), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U11234 ( .A1(n8724), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6771), 
        .B2(n13555), .ZN(n8708) );
  INV_X1 U11235 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U11236 ( .A1(n8710), .A2(n13538), .ZN(n8711) );
  NAND2_X1 U11237 ( .A1(n8728), .A2(n8711), .ZN(n13742) );
  OR2_X1 U11238 ( .A1(n13742), .A2(n8613), .ZN(n8715) );
  NAND2_X1 U11239 ( .A1(n8859), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11240 ( .A1(n9159), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11241 ( .A1(n9158), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8712) );
  NAND4_X1 U11242 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n13504) );
  NAND2_X1 U11243 ( .A1(n13957), .A2(n13374), .ZN(n8716) );
  INV_X1 U11244 ( .A(n8718), .ZN(n8720) );
  OAI21_X1 U11245 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8723) );
  XNOR2_X1 U11246 ( .A(n8723), .B(n8722), .ZN(n12065) );
  NAND2_X1 U11247 ( .A1(n12065), .A2(n9188), .ZN(n8726) );
  AOI22_X1 U11248 ( .A1(n8724), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8957), 
        .B2(n6771), .ZN(n8725) );
  INV_X1 U11249 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U11250 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND2_X1 U11251 ( .A1(n8744), .A2(n8729), .ZN(n13734) );
  OR2_X1 U11252 ( .A1(n13734), .A2(n8613), .ZN(n8734) );
  INV_X1 U11253 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13559) );
  OR2_X1 U11254 ( .A1(n6593), .A2(n13559), .ZN(n8732) );
  INV_X1 U11255 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8730) );
  OR2_X1 U11256 ( .A1(n9162), .A2(n8730), .ZN(n8731) );
  AND2_X1 U11257 ( .A1(n8732), .A2(n8731), .ZN(n8733) );
  OAI211_X1 U11258 ( .C1(n8430), .C2(n13552), .A(n8734), .B(n8733), .ZN(n13503) );
  INV_X1 U11259 ( .A(n13503), .ZN(n13713) );
  AND2_X1 U11260 ( .A1(n13951), .A2(n13713), .ZN(n8735) );
  NAND2_X1 U11261 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11262 ( .A1(n8739), .A2(n8738), .ZN(n12084) );
  OR2_X1 U11263 ( .A1(n12084), .A2(n8802), .ZN(n8742) );
  OR2_X1 U11264 ( .A1(n8740), .A2(n10921), .ZN(n8741) );
  NAND2_X1 U11265 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U11266 ( .A1(n8756), .A2(n8745), .ZN(n13717) );
  AOI22_X1 U11267 ( .A1(n9159), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n8859), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11268 ( .A1(n9158), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8746) );
  OAI211_X1 U11269 ( .C1(n13717), .C2(n8613), .A(n8747), .B(n8746), .ZN(n13502) );
  INV_X1 U11270 ( .A(n13502), .ZN(n13375) );
  NAND2_X1 U11271 ( .A1(n13948), .A2(n13375), .ZN(n8749) );
  OR2_X1 U11272 ( .A1(n13948), .A2(n13375), .ZN(n8748) );
  NAND2_X1 U11273 ( .A1(n8749), .A2(n8748), .ZN(n13710) );
  OR2_X1 U11274 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11275 ( .A1(n8750), .A2(n8753), .ZN(n12099) );
  OR2_X1 U11276 ( .A1(n12099), .A2(n8802), .ZN(n8755) );
  OR2_X1 U11277 ( .A1(n8740), .A2(n11036), .ZN(n8754) );
  NAND2_X1 U11278 ( .A1(n8756), .A2(n13395), .ZN(n8757) );
  AND2_X1 U11279 ( .A1(n8772), .A2(n8757), .ZN(n13701) );
  NAND2_X1 U11280 ( .A1(n13701), .A2(n6577), .ZN(n8763) );
  INV_X1 U11281 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11282 ( .A1(n9159), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11283 ( .A1(n8859), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8758) );
  OAI211_X1 U11284 ( .C1(n8760), .C2(n8430), .A(n8759), .B(n8758), .ZN(n8761)
         );
  INV_X1 U11285 ( .A(n8761), .ZN(n8762) );
  OR2_X1 U11286 ( .A1(n13943), .A2(n13714), .ZN(n8764) );
  NAND2_X1 U11287 ( .A1(n13943), .A2(n13714), .ZN(n8765) );
  NAND2_X1 U11288 ( .A1(n11920), .A2(n8766), .ZN(n8767) );
  NAND2_X1 U11289 ( .A1(n8768), .A2(n8767), .ZN(n11318) );
  OR2_X1 U11290 ( .A1(n11318), .A2(n8802), .ZN(n8770) );
  OR2_X1 U11291 ( .A1(n8740), .A2(n11320), .ZN(n8769) );
  INV_X1 U11292 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11293 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U11294 ( .A1(n8788), .A2(n8773), .ZN(n13467) );
  OR2_X1 U11295 ( .A1(n13467), .A2(n8613), .ZN(n8779) );
  INV_X1 U11296 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11297 ( .A1(n8859), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11298 ( .A1(n9159), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8774) );
  OAI211_X1 U11299 ( .C1(n8776), .C2(n8430), .A(n8775), .B(n8774), .ZN(n8777)
         );
  INV_X1 U11300 ( .A(n8777), .ZN(n8778) );
  INV_X1 U11301 ( .A(n13461), .ZN(n8780) );
  NAND2_X1 U11302 ( .A1(n13937), .A2(n8780), .ZN(n8781) );
  NAND2_X1 U11303 ( .A1(n8782), .A2(n8781), .ZN(n13679) );
  XNOR2_X1 U11304 ( .A(n8783), .B(SI_23_), .ZN(n8784) );
  NAND2_X1 U11305 ( .A1(n12111), .A2(n9188), .ZN(n8787) );
  OR2_X1 U11306 ( .A1(n8740), .A2(n11429), .ZN(n8786) );
  NAND2_X1 U11307 ( .A1(n8788), .A2(n13365), .ZN(n8789) );
  AND2_X1 U11308 ( .A1(n8804), .A2(n8789), .ZN(n13666) );
  NAND2_X1 U11309 ( .A1(n13666), .A2(n6577), .ZN(n8794) );
  INV_X1 U11310 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U11311 ( .A1(n8859), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8791) );
  INV_X1 U11312 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13060) );
  OR2_X1 U11313 ( .A1(n6593), .A2(n13060), .ZN(n8790) );
  OAI211_X1 U11314 ( .C1(n13093), .C2(n8430), .A(n8791), .B(n8790), .ZN(n8792)
         );
  INV_X1 U11315 ( .A(n8792), .ZN(n8793) );
  INV_X1 U11316 ( .A(n13466), .ZN(n9236) );
  NAND2_X1 U11317 ( .A1(n13673), .A2(n9236), .ZN(n8795) );
  NAND2_X1 U11318 ( .A1(n13661), .A2(n8795), .ZN(n8797) );
  OR2_X1 U11319 ( .A1(n13673), .A2(n9236), .ZN(n8796) );
  NAND2_X1 U11320 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  OR2_X1 U11321 ( .A1(n8740), .A2(n11618), .ZN(n8803) );
  INV_X1 U11322 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U11323 ( .A1(n8804), .A2(n13443), .ZN(n8805) );
  NAND2_X1 U11324 ( .A1(n8829), .A2(n8805), .ZN(n13645) );
  INV_X1 U11325 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13653) );
  NAND2_X1 U11326 ( .A1(n8859), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11327 ( .A1(n9159), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8806) );
  OAI211_X1 U11328 ( .C1(n13653), .C2(n8430), .A(n8807), .B(n8806), .ZN(n8808)
         );
  INV_X1 U11329 ( .A(n8808), .ZN(n8809) );
  NAND2_X1 U11330 ( .A1(n13925), .A2(n13410), .ZN(n8811) );
  XNOR2_X1 U11331 ( .A(n8813), .B(n8812), .ZN(n12424) );
  NAND2_X1 U11332 ( .A1(n12424), .A2(n9188), .ZN(n8815) );
  OR2_X1 U11333 ( .A1(n8740), .A2(n14023), .ZN(n8814) );
  XNOR2_X1 U11334 ( .A(n8829), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13638) );
  NAND2_X1 U11335 ( .A1(n13638), .A2(n6577), .ZN(n8820) );
  INV_X1 U11336 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13089) );
  NAND2_X1 U11337 ( .A1(n9158), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11338 ( .A1(n8859), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8816) );
  OAI211_X1 U11339 ( .C1(n6593), .C2(n13089), .A(n8817), .B(n8816), .ZN(n8818)
         );
  INV_X1 U11340 ( .A(n8818), .ZN(n8819) );
  XNOR2_X1 U11341 ( .A(n13920), .B(n13500), .ZN(n13630) );
  INV_X1 U11342 ( .A(n13500), .ZN(n13484) );
  NAND2_X1 U11343 ( .A1(n13920), .A2(n13484), .ZN(n8821) );
  NAND2_X1 U11344 ( .A1(n12295), .A2(n9188), .ZN(n8827) );
  OR2_X1 U11345 ( .A1(n8740), .A2(n14017), .ZN(n8826) );
  INV_X1 U11346 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13408) );
  INV_X1 U11347 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8828) );
  OAI21_X1 U11348 ( .B1(n8829), .B2(n13408), .A(n8828), .ZN(n8830) );
  NAND2_X1 U11349 ( .A1(n13622), .A2(n6577), .ZN(n8836) );
  INV_X1 U11350 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U11351 ( .A1(n9159), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11352 ( .A1(n8859), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8831) );
  OAI211_X1 U11353 ( .C1(n8833), .C2(n8430), .A(n8832), .B(n8831), .ZN(n8834)
         );
  INV_X1 U11354 ( .A(n8834), .ZN(n8835) );
  INV_X1 U11355 ( .A(n13633), .ZN(n13411) );
  OR2_X1 U11356 ( .A1(n13913), .A2(n13411), .ZN(n8837) );
  NAND2_X1 U11357 ( .A1(n13913), .A2(n13411), .ZN(n8838) );
  XNOR2_X1 U11358 ( .A(n8839), .B(SI_27_), .ZN(n8840) );
  OR2_X1 U11359 ( .A1(n8740), .A2(n14016), .ZN(n8842) );
  NAND2_X2 U11360 ( .A1(n8843), .A2(n8842), .ZN(n13905) );
  INV_X1 U11361 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U11362 ( .A1(n8844), .A2(n13069), .ZN(n8845) );
  NAND2_X1 U11363 ( .A1(n8846), .A2(n8845), .ZN(n13604) );
  OR2_X1 U11364 ( .A1(n13604), .A2(n8613), .ZN(n8851) );
  INV_X1 U11365 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U11366 ( .A1(n9159), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U11367 ( .A1(n8859), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8847) );
  OAI211_X1 U11368 ( .C1(n13603), .C2(n8430), .A(n8848), .B(n8847), .ZN(n8849)
         );
  INV_X1 U11369 ( .A(n8849), .ZN(n8850) );
  INV_X1 U11370 ( .A(n13499), .ZN(n8852) );
  NAND2_X1 U11371 ( .A1(n13899), .A2(n13498), .ZN(n8916) );
  OR2_X1 U11372 ( .A1(n13899), .A2(n13498), .ZN(n8853) );
  NAND2_X1 U11373 ( .A1(n8916), .A2(n8853), .ZN(n13584) );
  INV_X1 U11374 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11870) );
  MUX2_X1 U11375 ( .A(n14713), .B(n11870), .S(n11919), .Z(n9151) );
  XNOR2_X1 U11376 ( .A(n9151), .B(SI_29_), .ZN(n9148) );
  XNOR2_X1 U11377 ( .A(n9149), .B(n9148), .ZN(n12195) );
  NAND2_X1 U11378 ( .A1(n12195), .A2(n9188), .ZN(n8858) );
  OR2_X1 U11379 ( .A1(n8740), .A2(n11870), .ZN(n8857) );
  INV_X1 U11380 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U11381 ( .A1(n9158), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11382 ( .A1(n8859), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8860) );
  OAI211_X1 U11383 ( .C1(n12978), .C2(n6593), .A(n8861), .B(n8860), .ZN(n8862)
         );
  INV_X1 U11384 ( .A(n8862), .ZN(n8863) );
  OAI21_X1 U11385 ( .B1(n12430), .B2(n8613), .A(n8863), .ZN(n13497) );
  XNOR2_X1 U11386 ( .A(n12429), .B(n13497), .ZN(n9254) );
  NAND2_X1 U11387 ( .A1(n6587), .A2(n8874), .ZN(n9164) );
  NAND2_X1 U11388 ( .A1(n9163), .A2(n10718), .ZN(n8865) );
  INV_X2 U11389 ( .A(n13712), .ZN(n15313) );
  INV_X1 U11390 ( .A(n9855), .ZN(n8866) );
  INV_X1 U11391 ( .A(n14014), .ZN(n9845) );
  AOI21_X1 U11392 ( .B1(n9845), .B2(P2_B_REG_SCAN_IN), .A(n13872), .ZN(n13573)
         );
  INV_X1 U11393 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8867) );
  OR2_X1 U11394 ( .A1(n6593), .A2(n8867), .ZN(n8872) );
  INV_X1 U11395 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8868) );
  OR2_X1 U11396 ( .A1(n8430), .A2(n8868), .ZN(n8871) );
  INV_X1 U11397 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8869) );
  OR2_X1 U11398 ( .A1(n9162), .A2(n8869), .ZN(n8870) );
  INV_X1 U11399 ( .A(n9166), .ZN(n13496) );
  XNOR2_X1 U11400 ( .A(n8874), .B(n10647), .ZN(n8875) );
  AND2_X1 U11401 ( .A1(n8959), .A2(n8876), .ZN(n10248) );
  OAI22_X1 U11402 ( .A1(n6573), .A2(n10248), .B1(n13515), .B2(n8968), .ZN(
        n15319) );
  NAND2_X1 U11403 ( .A1(n15319), .A2(n15320), .ZN(n8878) );
  NAND2_X1 U11404 ( .A1(n6854), .A2(n7258), .ZN(n8877) );
  NAND2_X1 U11405 ( .A1(n8878), .A2(n8877), .ZN(n10161) );
  NAND2_X1 U11406 ( .A1(n10161), .A2(n9238), .ZN(n8880) );
  NAND2_X1 U11407 ( .A1(n10402), .A2(n10712), .ZN(n8879) );
  NAND2_X1 U11408 ( .A1(n8880), .A2(n8879), .ZN(n10696) );
  NAND2_X1 U11409 ( .A1(n10696), .A2(n9239), .ZN(n8882) );
  NAND2_X1 U11410 ( .A1(n6814), .A2(n10706), .ZN(n8881) );
  NAND2_X1 U11411 ( .A1(n8882), .A2(n8881), .ZN(n10649) );
  INV_X1 U11412 ( .A(n10650), .ZN(n8883) );
  NAND2_X1 U11413 ( .A1(n10649), .A2(n8883), .ZN(n8886) );
  INV_X1 U11414 ( .A(n15390), .ZN(n10658) );
  NAND2_X1 U11415 ( .A1(n8884), .A2(n10658), .ZN(n8885) );
  NAND2_X1 U11416 ( .A1(n8886), .A2(n8885), .ZN(n10676) );
  INV_X1 U11417 ( .A(n10679), .ZN(n10675) );
  INV_X1 U11418 ( .A(n15396), .ZN(n10691) );
  NAND2_X1 U11419 ( .A1(n10691), .A2(n10573), .ZN(n8887) );
  XNOR2_X1 U11420 ( .A(n15404), .B(n13509), .ZN(n10663) );
  INV_X1 U11421 ( .A(n10663), .ZN(n8888) );
  OR2_X1 U11422 ( .A1(n13869), .A2(n13868), .ZN(n8890) );
  NAND2_X1 U11423 ( .A1(n13889), .A2(n13853), .ZN(n8889) );
  NAND2_X1 U11424 ( .A1(n13865), .A2(n13508), .ZN(n8891) );
  NAND2_X1 U11425 ( .A1(n13811), .A2(n13815), .ZN(n13813) );
  NAND2_X1 U11426 ( .A1(n15435), .A2(n13798), .ZN(n8892) );
  OR2_X1 U11427 ( .A1(n13808), .A2(n13814), .ZN(n8893) );
  NAND2_X1 U11428 ( .A1(n13796), .A2(n8893), .ZN(n8895) );
  NAND2_X1 U11429 ( .A1(n13808), .A2(n13814), .ZN(n8894) );
  NOR2_X1 U11430 ( .A1(n13792), .A2(n13506), .ZN(n8896) );
  NAND2_X1 U11431 ( .A1(n13792), .A2(n13506), .ZN(n8897) );
  XNOR2_X1 U11432 ( .A(n13981), .B(n11498), .ZN(n13971) );
  INV_X1 U11433 ( .A(n13971), .ZN(n13973) );
  XNOR2_X1 U11434 ( .A(n13967), .B(n9077), .ZN(n13764) );
  INV_X1 U11435 ( .A(n13764), .ZN(n13766) );
  OR2_X2 U11436 ( .A1(n13767), .A2(n13766), .ZN(n13769) );
  NAND2_X1 U11437 ( .A1(n13967), .A2(n13505), .ZN(n8898) );
  AND2_X1 U11438 ( .A1(n13962), .A2(n13770), .ZN(n8899) );
  OR2_X1 U11439 ( .A1(n13962), .A2(n13770), .ZN(n8900) );
  XNOR2_X1 U11440 ( .A(n13957), .B(n13374), .ZN(n13747) );
  NOR2_X1 U11441 ( .A1(n13951), .A2(n13503), .ZN(n8901) );
  NAND2_X1 U11442 ( .A1(n13951), .A2(n13503), .ZN(n8902) );
  NAND2_X1 U11443 ( .A1(n8903), .A2(n8902), .ZN(n13706) );
  AND2_X1 U11444 ( .A1(n13948), .A2(n13502), .ZN(n8905) );
  OR2_X1 U11445 ( .A1(n13948), .A2(n13502), .ZN(n8904) );
  NOR2_X1 U11446 ( .A1(n13943), .A2(n13501), .ZN(n8906) );
  OR2_X1 U11447 ( .A1(n13694), .A2(n8906), .ZN(n8908) );
  NAND2_X1 U11448 ( .A1(n13943), .A2(n13501), .ZN(n8907) );
  NAND2_X1 U11449 ( .A1(n8908), .A2(n8907), .ZN(n13678) );
  NAND2_X1 U11450 ( .A1(n13678), .A2(n13679), .ZN(n8910) );
  NAND2_X1 U11451 ( .A1(n13937), .A2(n13461), .ZN(n8909) );
  AND2_X1 U11452 ( .A1(n13673), .A2(n13466), .ZN(n8911) );
  INV_X1 U11453 ( .A(n13646), .ZN(n13657) );
  NAND2_X1 U11454 ( .A1(n13920), .A2(n13500), .ZN(n8912) );
  AND2_X1 U11455 ( .A1(n13913), .A2(n13633), .ZN(n8914) );
  INV_X1 U11456 ( .A(n13584), .ZN(n13589) );
  NAND2_X1 U11457 ( .A1(n13590), .A2(n13589), .ZN(n13588) );
  NAND2_X1 U11458 ( .A1(n13588), .A2(n8916), .ZN(n8917) );
  INV_X1 U11459 ( .A(n13905), .ZN(n13605) );
  INV_X1 U11460 ( .A(n13920), .ZN(n13641) );
  NAND2_X1 U11461 ( .A1(n10864), .A2(n10721), .ZN(n15321) );
  INV_X1 U11462 ( .A(n15404), .ZN(n10671) );
  INV_X1 U11463 ( .A(n13889), .ZN(n15415) );
  INV_X1 U11464 ( .A(n13808), .ZN(n14974) );
  AND2_X1 U11465 ( .A1(n13825), .A2(n14974), .ZN(n11376) );
  INV_X1 U11466 ( .A(n11454), .ZN(n11380) );
  INV_X1 U11467 ( .A(n13792), .ZN(n14967) );
  NOR2_X1 U11468 ( .A1(n13925), .A2(n13671), .ZN(n13652) );
  NAND2_X2 U11469 ( .A1(n10719), .A2(n10920), .ZN(n13979) );
  AOI211_X1 U11470 ( .C1(n12429), .C2(n13591), .A(n13979), .B(n13579), .ZN(
        n12436) );
  AOI21_X1 U11471 ( .B1(n15434), .B2(n12429), .A(n12436), .ZN(n8921) );
  INV_X1 U11472 ( .A(n12580), .ZN(n11817) );
  NAND2_X1 U11473 ( .A1(n12701), .A2(n11817), .ZN(n9289) );
  NAND2_X1 U11474 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n14016), .ZN(n8924) );
  AOI22_X1 U11475 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14012), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11868), .ZN(n8926) );
  XNOR2_X1 U11476 ( .A(n9291), .B(n8926), .ZN(n12299) );
  NAND2_X1 U11477 ( .A1(n12299), .A2(n8927), .ZN(n8929) );
  NAND2_X1 U11478 ( .A1(n9294), .A2(SI_28_), .ZN(n8928) );
  NAND2_X1 U11479 ( .A1(n12691), .A2(n9304), .ZN(n9290) );
  OR2_X1 U11480 ( .A1(n12701), .A2(n12580), .ZN(n8931) );
  NAND2_X1 U11481 ( .A1(n8934), .A2(n12861), .ZN(n8935) );
  INV_X1 U11482 ( .A(n14939), .ZN(n8936) );
  NAND2_X1 U11483 ( .A1(n11636), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8940) );
  INV_X1 U11484 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9308) );
  OR2_X1 U11485 ( .A1(n6570), .A2(n9308), .ZN(n8939) );
  INV_X1 U11486 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n8937) );
  OR2_X1 U11487 ( .A1(n11637), .A2(n8937), .ZN(n8938) );
  NAND4_X1 U11488 ( .A1(n11643), .A2(n8940), .A3(n8939), .A4(n8938), .ZN(
        n12578) );
  AOI22_X1 U11489 ( .A1(n8165), .A2(n12578), .B1(n12580), .B2(n12849), .ZN(
        n8941) );
  MUX2_X1 U11490 ( .A(n8954), .B(n8943), .S(n15628), .Z(n8944) );
  INV_X1 U11491 ( .A(n12691), .ZN(n8955) );
  NAND2_X1 U11492 ( .A1(n8944), .A2(n7641), .ZN(P3_U3487) );
  NAND3_X1 U11493 ( .A1(n13265), .A2(n9319), .A3(n8947), .ZN(n9397) );
  NOR2_X1 U11494 ( .A1(n8226), .A2(n11834), .ZN(n10221) );
  INV_X1 U11495 ( .A(n9391), .ZN(n9398) );
  NOR2_X1 U11496 ( .A1(n10221), .A2(n9398), .ZN(n8951) );
  INV_X1 U11497 ( .A(n13265), .ZN(n8949) );
  INV_X1 U11498 ( .A(n9319), .ZN(n8948) );
  NAND3_X1 U11499 ( .A1(n8949), .A2(n8948), .A3(n8947), .ZN(n9404) );
  INV_X1 U11500 ( .A(n9396), .ZN(n8950) );
  OAI22_X1 U11501 ( .A1(n9397), .A2(n8951), .B1(n9404), .B2(n8950), .ZN(n8952)
         );
  MUX2_X1 U11502 ( .A(n8954), .B(n8953), .S(n15612), .Z(n8956) );
  NAND2_X1 U11503 ( .A1(n8956), .A2(n7642), .ZN(P3_U3455) );
  AND2_X1 U11504 ( .A1(n8957), .A2(n11319), .ZN(n8958) );
  AND2_X1 U11505 ( .A1(n8958), .A2(n10647), .ZN(n9192) );
  OAI21_X1 U11506 ( .B1(n9192), .B2(n10721), .A(n9237), .ZN(n8962) );
  OR2_X1 U11507 ( .A1(n8960), .A2(n8963), .ZN(n9194) );
  NAND2_X1 U11508 ( .A1(n8959), .A2(n9194), .ZN(n8961) );
  NAND2_X1 U11509 ( .A1(n8962), .A2(n8961), .ZN(n8965) );
  NAND3_X1 U11510 ( .A1(n9237), .A2(n10647), .A3(n8963), .ZN(n8964) );
  NAND2_X1 U11511 ( .A1(n13515), .A2(n9192), .ZN(n8967) );
  NAND2_X1 U11512 ( .A1(n9194), .A2(n8968), .ZN(n8966) );
  NAND2_X1 U11513 ( .A1(n8967), .A2(n8966), .ZN(n8970) );
  AOI22_X1 U11514 ( .A1(n13515), .A2(n9194), .B1(n9192), .B2(n8968), .ZN(n8969) );
  AOI21_X1 U11515 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n8973) );
  NOR2_X1 U11516 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  NAND2_X1 U11517 ( .A1(n13514), .A2(n9137), .ZN(n8975) );
  NAND2_X1 U11518 ( .A1(n9192), .A2(n15318), .ZN(n8974) );
  AOI22_X1 U11519 ( .A1(n13514), .A2(n9121), .B1(n9137), .B2(n15318), .ZN(
        n8976) );
  AOI21_X1 U11520 ( .B1(n8979), .B2(n8978), .A(n8976), .ZN(n8977) );
  INV_X1 U11521 ( .A(n8977), .ZN(n8980) );
  INV_X1 U11522 ( .A(n9192), .ZN(n9032) );
  INV_X1 U11523 ( .A(n9032), .ZN(n9207) );
  NAND2_X1 U11524 ( .A1(n13513), .A2(n9207), .ZN(n8982) );
  NAND2_X1 U11525 ( .A1(n9194), .A2(n15224), .ZN(n8981) );
  NAND2_X1 U11526 ( .A1(n8982), .A2(n8981), .ZN(n8988) );
  NAND2_X1 U11527 ( .A1(n8987), .A2(n8988), .ZN(n8986) );
  NAND2_X1 U11528 ( .A1(n13513), .A2(n9137), .ZN(n8984) );
  NAND2_X1 U11529 ( .A1(n9207), .A2(n15224), .ZN(n8983) );
  NAND2_X1 U11530 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NAND2_X1 U11531 ( .A1(n8986), .A2(n8985), .ZN(n8991) );
  INV_X1 U11532 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U11533 ( .A1(n6586), .A2(n8989), .ZN(n8990) );
  NAND2_X1 U11534 ( .A1(n8991), .A2(n8990), .ZN(n8996) );
  NAND2_X1 U11535 ( .A1(n13512), .A2(n9137), .ZN(n8993) );
  NAND2_X1 U11536 ( .A1(n9192), .A2(n15383), .ZN(n8992) );
  NAND2_X1 U11537 ( .A1(n8993), .A2(n8992), .ZN(n8995) );
  AOI22_X1 U11538 ( .A1(n13512), .A2(n9121), .B1(n9194), .B2(n15383), .ZN(
        n8994) );
  NAND2_X1 U11539 ( .A1(n13511), .A2(n9207), .ZN(n8998) );
  NAND2_X1 U11540 ( .A1(n9194), .A2(n15390), .ZN(n8997) );
  NAND2_X1 U11541 ( .A1(n8998), .A2(n8997), .ZN(n9003) );
  INV_X1 U11542 ( .A(n9121), .ZN(n9264) );
  NAND2_X1 U11543 ( .A1(n13511), .A2(n9137), .ZN(n8999) );
  OAI21_X1 U11544 ( .B1(n10658), .B2(n9264), .A(n8999), .ZN(n9000) );
  NAND2_X1 U11545 ( .A1(n9001), .A2(n9000), .ZN(n9007) );
  INV_X1 U11546 ( .A(n9002), .ZN(n9005) );
  INV_X1 U11547 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U11548 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U11549 ( .A1(n9007), .A2(n9006), .ZN(n9013) );
  NAND2_X1 U11550 ( .A1(n15396), .A2(n9207), .ZN(n9009) );
  NAND2_X1 U11551 ( .A1(n13510), .A2(n9132), .ZN(n9008) );
  NAND2_X1 U11552 ( .A1(n9009), .A2(n9008), .ZN(n9012) );
  AOI22_X1 U11553 ( .A1(n15396), .A2(n9194), .B1(n13510), .B2(n9195), .ZN(
        n9010) );
  NAND2_X1 U11554 ( .A1(n15404), .A2(n9137), .ZN(n9015) );
  NAND2_X1 U11555 ( .A1(n13509), .A2(n9121), .ZN(n9014) );
  NAND2_X1 U11556 ( .A1(n15404), .A2(n9207), .ZN(n9016) );
  OAI21_X1 U11557 ( .B1(n13875), .B2(n9057), .A(n9016), .ZN(n9017) );
  NAND2_X1 U11558 ( .A1(n9018), .A2(n9017), .ZN(n9022) );
  NAND2_X1 U11559 ( .A1(n9020), .A2(n6675), .ZN(n9021) );
  NAND2_X1 U11560 ( .A1(n13889), .A2(n9207), .ZN(n9024) );
  NAND2_X1 U11561 ( .A1(n13853), .A2(n9132), .ZN(n9023) );
  NAND2_X1 U11562 ( .A1(n9024), .A2(n9023), .ZN(n9026) );
  AOI22_X1 U11563 ( .A1(n13889), .A2(n9137), .B1(n9192), .B2(n13853), .ZN(
        n9025) );
  NAND2_X1 U11564 ( .A1(n13865), .A2(n9132), .ZN(n9029) );
  NAND2_X1 U11565 ( .A1(n13508), .A2(n9207), .ZN(n9028) );
  NAND2_X1 U11566 ( .A1(n9029), .A2(n9028), .ZN(n9031) );
  AOI22_X1 U11567 ( .A1(n13865), .A2(n9121), .B1(n13508), .B2(n9132), .ZN(
        n9030) );
  INV_X1 U11568 ( .A(n9032), .ZN(n9195) );
  NAND2_X1 U11569 ( .A1(n13845), .A2(n9195), .ZN(n9034) );
  NAND2_X1 U11570 ( .A1(n13852), .A2(n9132), .ZN(n9033) );
  NAND2_X1 U11571 ( .A1(n9034), .A2(n9033), .ZN(n9038) );
  NAND2_X1 U11572 ( .A1(n13845), .A2(n9132), .ZN(n9035) );
  NAND2_X1 U11573 ( .A1(n15435), .A2(n9132), .ZN(n9041) );
  NAND2_X1 U11574 ( .A1(n13798), .A2(n9195), .ZN(n9040) );
  NAND2_X1 U11575 ( .A1(n9041), .A2(n9040), .ZN(n9044) );
  AOI22_X1 U11576 ( .A1(n15435), .A2(n9121), .B1(n13798), .B2(n9132), .ZN(
        n9042) );
  AOI21_X1 U11577 ( .B1(n9045), .B2(n9044), .A(n9042), .ZN(n9043) );
  INV_X1 U11578 ( .A(n9043), .ZN(n9046) );
  NAND2_X1 U11579 ( .A1(n13808), .A2(n9195), .ZN(n9048) );
  NAND2_X1 U11580 ( .A1(n13814), .A2(n9132), .ZN(n9047) );
  NAND2_X1 U11581 ( .A1(n9048), .A2(n9047), .ZN(n9054) );
  NAND2_X1 U11582 ( .A1(n9053), .A2(n9054), .ZN(n9052) );
  NAND2_X1 U11583 ( .A1(n13808), .A2(n9132), .ZN(n9049) );
  OAI21_X1 U11584 ( .B1(n9050), .B2(n9264), .A(n9049), .ZN(n9051) );
  NAND2_X1 U11585 ( .A1(n11454), .A2(n9132), .ZN(n9059) );
  NAND2_X1 U11586 ( .A1(n13797), .A2(n9207), .ZN(n9058) );
  NAND2_X1 U11587 ( .A1(n9059), .A2(n9058), .ZN(n9061) );
  AOI22_X1 U11588 ( .A1(n11454), .A2(n9121), .B1(n13797), .B2(n9132), .ZN(
        n9060) );
  NAND2_X1 U11589 ( .A1(n13792), .A2(n9195), .ZN(n9063) );
  NAND2_X1 U11590 ( .A1(n13506), .A2(n9132), .ZN(n9062) );
  NAND2_X1 U11591 ( .A1(n9063), .A2(n9062), .ZN(n9067) );
  NAND2_X1 U11592 ( .A1(n9068), .A2(n9067), .ZN(n9066) );
  NAND2_X1 U11593 ( .A1(n13792), .A2(n9132), .ZN(n9064) );
  OAI21_X1 U11594 ( .B1(n11300), .B2(n9264), .A(n9064), .ZN(n9065) );
  NAND2_X1 U11595 ( .A1(n9066), .A2(n9065), .ZN(n9070) );
  NAND2_X1 U11596 ( .A1(n13981), .A2(n9132), .ZN(n9072) );
  NAND2_X1 U11597 ( .A1(n13784), .A2(n9195), .ZN(n9071) );
  AOI22_X1 U11598 ( .A1(n13981), .A2(n9121), .B1(n13784), .B2(n9132), .ZN(
        n9073) );
  NAND2_X1 U11599 ( .A1(n13967), .A2(n9195), .ZN(n9075) );
  NAND2_X1 U11600 ( .A1(n13505), .A2(n9132), .ZN(n9074) );
  NAND2_X1 U11601 ( .A1(n9075), .A2(n9074), .ZN(n9080) );
  NAND2_X1 U11602 ( .A1(n9081), .A2(n9080), .ZN(n9079) );
  NAND2_X1 U11603 ( .A1(n13967), .A2(n9132), .ZN(n9076) );
  OAI21_X1 U11604 ( .B1(n9077), .B2(n9264), .A(n9076), .ZN(n9078) );
  NAND2_X1 U11605 ( .A1(n9079), .A2(n9078), .ZN(n9082) );
  NAND2_X1 U11606 ( .A1(n13962), .A2(n9137), .ZN(n9084) );
  NAND2_X1 U11607 ( .A1(n13770), .A2(n9195), .ZN(n9083) );
  NAND2_X1 U11608 ( .A1(n9084), .A2(n9083), .ZN(n9087) );
  AOI22_X1 U11609 ( .A1(n13962), .A2(n9121), .B1(n13770), .B2(n9132), .ZN(
        n9085) );
  INV_X1 U11610 ( .A(n9086), .ZN(n9089) );
  NAND2_X1 U11611 ( .A1(n13957), .A2(n9195), .ZN(n9091) );
  NAND2_X1 U11612 ( .A1(n13504), .A2(n9132), .ZN(n9090) );
  NAND2_X1 U11613 ( .A1(n13957), .A2(n9137), .ZN(n9092) );
  NAND2_X1 U11614 ( .A1(n13951), .A2(n9137), .ZN(n9095) );
  NAND2_X1 U11615 ( .A1(n13503), .A2(n9195), .ZN(n9094) );
  NAND2_X1 U11616 ( .A1(n9095), .A2(n9094), .ZN(n9098) );
  AOI22_X1 U11617 ( .A1(n13951), .A2(n9207), .B1(n13503), .B2(n9132), .ZN(
        n9096) );
  INV_X1 U11618 ( .A(n9097), .ZN(n9100) );
  NAND2_X1 U11619 ( .A1(n9100), .A2(n7638), .ZN(n9106) );
  NAND2_X1 U11620 ( .A1(n13948), .A2(n9195), .ZN(n9102) );
  NAND2_X1 U11621 ( .A1(n13502), .A2(n9137), .ZN(n9101) );
  NAND2_X1 U11622 ( .A1(n9102), .A2(n9101), .ZN(n9107) );
  NAND2_X1 U11623 ( .A1(n9106), .A2(n9107), .ZN(n9105) );
  NAND2_X1 U11624 ( .A1(n13948), .A2(n9137), .ZN(n9103) );
  OAI21_X1 U11625 ( .B1(n13375), .B2(n9264), .A(n9103), .ZN(n9104) );
  NAND2_X1 U11626 ( .A1(n9105), .A2(n9104), .ZN(n9111) );
  NAND2_X1 U11627 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U11628 ( .A1(n13943), .A2(n9137), .ZN(n9113) );
  NAND2_X1 U11629 ( .A1(n13501), .A2(n9195), .ZN(n9112) );
  NAND2_X1 U11630 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  AOI22_X1 U11631 ( .A1(n13943), .A2(n9207), .B1(n13501), .B2(n9132), .ZN(
        n9114) );
  NAND2_X1 U11632 ( .A1(n13937), .A2(n9195), .ZN(n9118) );
  NAND2_X1 U11633 ( .A1(n13461), .A2(n9137), .ZN(n9117) );
  NAND2_X1 U11634 ( .A1(n9118), .A2(n9117), .ZN(n9120) );
  AOI22_X1 U11635 ( .A1(n13937), .A2(n9194), .B1(n9192), .B2(n13461), .ZN(
        n9119) );
  AOI22_X1 U11636 ( .A1(n13673), .A2(n9194), .B1(n9121), .B2(n13466), .ZN(
        n9125) );
  AOI22_X1 U11637 ( .A1(n13673), .A2(n9121), .B1(n13466), .B2(n9132), .ZN(
        n9122) );
  NOR2_X1 U11638 ( .A1(n9123), .A2(n9122), .ZN(n9147) );
  INV_X1 U11639 ( .A(n9124), .ZN(n9130) );
  INV_X1 U11640 ( .A(n9125), .ZN(n9129) );
  NAND2_X1 U11641 ( .A1(n13925), .A2(n9137), .ZN(n9127) );
  NAND2_X1 U11642 ( .A1(n13632), .A2(n9195), .ZN(n9126) );
  NAND2_X1 U11643 ( .A1(n9127), .A2(n9126), .ZN(n9135) );
  AND2_X1 U11644 ( .A1(n13632), .A2(n9137), .ZN(n9128) );
  AOI21_X1 U11645 ( .B1(n13925), .B2(n9121), .A(n9128), .ZN(n9136) );
  AND2_X1 U11646 ( .A1(n13633), .A2(n9132), .ZN(n9131) );
  AOI21_X1 U11647 ( .B1(n13913), .B2(n9207), .A(n9131), .ZN(n9199) );
  NAND2_X1 U11648 ( .A1(n13913), .A2(n9132), .ZN(n9134) );
  NAND2_X1 U11649 ( .A1(n13633), .A2(n9195), .ZN(n9133) );
  NAND2_X1 U11650 ( .A1(n9134), .A2(n9133), .ZN(n9202) );
  AOI22_X1 U11651 ( .A1(n9199), .A2(n9202), .B1(n9136), .B2(n9135), .ZN(n9144)
         );
  NAND2_X1 U11652 ( .A1(n13920), .A2(n9207), .ZN(n9139) );
  NAND2_X1 U11653 ( .A1(n13500), .A2(n9137), .ZN(n9138) );
  NAND2_X1 U11654 ( .A1(n9139), .A2(n9138), .ZN(n9200) );
  INV_X1 U11655 ( .A(n9200), .ZN(n9142) );
  AND2_X1 U11656 ( .A1(n13500), .A2(n9192), .ZN(n9140) );
  AOI21_X1 U11657 ( .B1(n13920), .B2(n9194), .A(n9140), .ZN(n9201) );
  INV_X1 U11658 ( .A(n9201), .ZN(n9141) );
  NAND2_X1 U11659 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  OAI21_X1 U11660 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9218) );
  INV_X1 U11661 ( .A(SI_29_), .ZN(n9150) );
  NAND2_X1 U11662 ( .A1(n9151), .A2(n9150), .ZN(n9176) );
  NAND2_X1 U11663 ( .A1(n9187), .A2(n9176), .ZN(n9155) );
  MUX2_X1 U11664 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9680), .Z(n9152) );
  NAND2_X1 U11665 ( .A1(n9152), .A2(SI_30_), .ZN(n9179) );
  INV_X1 U11666 ( .A(n9152), .ZN(n9153) );
  INV_X1 U11667 ( .A(SI_30_), .ZN(n12427) );
  NAND2_X1 U11668 ( .A1(n9153), .A2(n12427), .ZN(n9177) );
  AND2_X1 U11669 ( .A1(n9179), .A2(n9177), .ZN(n9154) );
  NAND2_X1 U11670 ( .A1(n12224), .A2(n9188), .ZN(n9157) );
  INV_X1 U11671 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12438) );
  OR2_X1 U11672 ( .A1(n8740), .A2(n12438), .ZN(n9156) );
  INV_X1 U11673 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U11674 ( .A1(n9158), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11675 ( .A1(n9159), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9160) );
  OAI211_X1 U11676 ( .C1(n9162), .C2(n13076), .A(n9161), .B(n9160), .ZN(n13574) );
  NAND2_X1 U11677 ( .A1(n13574), .A2(n9137), .ZN(n9265) );
  OAI211_X1 U11678 ( .C1(n9164), .C2(n10718), .A(n9163), .B(n10181), .ZN(n9165) );
  INV_X1 U11679 ( .A(n9165), .ZN(n9167) );
  AOI21_X1 U11680 ( .B1(n9265), .B2(n9167), .A(n9166), .ZN(n9168) );
  AOI21_X1 U11681 ( .B1(n13571), .B2(n9207), .A(n9168), .ZN(n9230) );
  NAND2_X1 U11682 ( .A1(n13571), .A2(n9137), .ZN(n9170) );
  NAND2_X1 U11683 ( .A1(n13496), .A2(n9195), .ZN(n9169) );
  NAND2_X1 U11684 ( .A1(n9170), .A2(n9169), .ZN(n9229) );
  AND2_X1 U11685 ( .A1(n13497), .A2(n9137), .ZN(n9171) );
  AOI21_X1 U11686 ( .B1(n12429), .B2(n9207), .A(n9171), .ZN(n9227) );
  NAND2_X1 U11687 ( .A1(n12429), .A2(n9137), .ZN(n9173) );
  NAND2_X1 U11688 ( .A1(n13497), .A2(n9195), .ZN(n9172) );
  NAND2_X1 U11689 ( .A1(n9173), .A2(n9172), .ZN(n9226) );
  OAI22_X1 U11690 ( .A1(n9230), .A2(n9229), .B1(n9227), .B2(n9226), .ZN(n9191)
         );
  MUX2_X1 U11691 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11919), .Z(n9175) );
  INV_X1 U11692 ( .A(SI_31_), .ZN(n9174) );
  XNOR2_X1 U11693 ( .A(n9175), .B(n9174), .ZN(n9180) );
  NAND2_X1 U11694 ( .A1(n9180), .A2(n9179), .ZN(n9186) );
  NAND2_X1 U11695 ( .A1(n9177), .A2(n9176), .ZN(n9182) );
  NOR2_X1 U11696 ( .A1(n9182), .A2(n9180), .ZN(n9178) );
  NAND2_X1 U11697 ( .A1(n9187), .A2(n9178), .ZN(n9185) );
  INV_X1 U11698 ( .A(n9180), .ZN(n9183) );
  XNOR2_X1 U11699 ( .A(n9180), .B(n9179), .ZN(n9181) );
  OAI21_X1 U11700 ( .B1(n9183), .B2(n9182), .A(n9181), .ZN(n9184) );
  NAND2_X1 U11701 ( .A1(n14001), .A2(n9188), .ZN(n9190) );
  INV_X1 U11702 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14004) );
  OR2_X1 U11703 ( .A1(n8740), .A2(n14004), .ZN(n9189) );
  XNOR2_X1 U11704 ( .A(n13575), .B(n13574), .ZN(n9257) );
  NAND2_X1 U11705 ( .A1(n9191), .A2(n9257), .ZN(n9232) );
  AND2_X1 U11706 ( .A1(n13498), .A2(n9192), .ZN(n9193) );
  AOI21_X1 U11707 ( .B1(n13899), .B2(n9194), .A(n9193), .ZN(n9223) );
  NAND2_X1 U11708 ( .A1(n13899), .A2(n9195), .ZN(n9197) );
  NAND2_X1 U11709 ( .A1(n13498), .A2(n9137), .ZN(n9196) );
  NAND2_X1 U11710 ( .A1(n9197), .A2(n9196), .ZN(n9222) );
  NAND2_X1 U11711 ( .A1(n9223), .A2(n9222), .ZN(n9198) );
  AND2_X1 U11712 ( .A1(n9232), .A2(n9198), .ZN(n9221) );
  INV_X1 U11713 ( .A(n9221), .ZN(n9216) );
  INV_X1 U11714 ( .A(n9199), .ZN(n9204) );
  AND2_X1 U11715 ( .A1(n9201), .A2(n9200), .ZN(n9203) );
  OR2_X1 U11716 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  INV_X1 U11717 ( .A(n9202), .ZN(n9205) );
  AOI22_X1 U11718 ( .A1(n9206), .A2(n9205), .B1(n9204), .B2(n9203), .ZN(n9214)
         );
  NAND2_X1 U11719 ( .A1(n13905), .A2(n9137), .ZN(n9209) );
  NAND2_X1 U11720 ( .A1(n13499), .A2(n9207), .ZN(n9208) );
  NAND2_X1 U11721 ( .A1(n9209), .A2(n9208), .ZN(n9219) );
  INV_X1 U11722 ( .A(n9219), .ZN(n9212) );
  AND2_X1 U11723 ( .A1(n13499), .A2(n9137), .ZN(n9210) );
  AOI21_X1 U11724 ( .B1(n13905), .B2(n9207), .A(n9210), .ZN(n9220) );
  NAND2_X1 U11725 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  NAND2_X1 U11726 ( .A1(n9218), .A2(n9217), .ZN(n9235) );
  NAND3_X1 U11727 ( .A1(n9221), .A2(n9220), .A3(n9219), .ZN(n9234) );
  INV_X1 U11728 ( .A(n9222), .ZN(n9225) );
  INV_X1 U11729 ( .A(n9223), .ZN(n9224) );
  AOI22_X1 U11730 ( .A1(n9227), .A2(n9226), .B1(n9225), .B2(n9224), .ZN(n9228)
         );
  NAND2_X1 U11731 ( .A1(n9228), .A2(n9257), .ZN(n9231) );
  AOI22_X1 U11732 ( .A1(n9232), .A2(n9231), .B1(n9230), .B2(n9229), .ZN(n9233)
         );
  INV_X1 U11733 ( .A(n9270), .ZN(n9263) );
  XNOR2_X1 U11734 ( .A(n13571), .B(n13496), .ZN(n9256) );
  XNOR2_X1 U11735 ( .A(n13913), .B(n13633), .ZN(n13617) );
  XNOR2_X1 U11736 ( .A(n13673), .B(n9236), .ZN(n13667) );
  XNOR2_X1 U11737 ( .A(n13943), .B(n13714), .ZN(n13695) );
  XNOR2_X1 U11738 ( .A(n13951), .B(n13713), .ZN(n13725) );
  XNOR2_X1 U11739 ( .A(n13962), .B(n13475), .ZN(n13759) );
  XNOR2_X1 U11740 ( .A(n13792), .B(n11300), .ZN(n13786) );
  NOR3_X1 U11741 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(n9241) );
  NAND4_X1 U11742 ( .A1(n9241), .A2(n10663), .A3(n10679), .A4(n10650), .ZN(
        n9242) );
  NOR2_X1 U11743 ( .A1(n9242), .A2(n13870), .ZN(n9245) );
  NAND4_X1 U11744 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n9247)
         );
  OR4_X1 U11745 ( .A1(n13786), .A2(n11381), .A3(n13799), .A4(n9247), .ZN(n9248) );
  OR4_X1 U11746 ( .A1(n13759), .A2(n13764), .A3(n13971), .A4(n9248), .ZN(n9249) );
  OR4_X1 U11747 ( .A1(n13710), .A2(n13747), .A3(n13725), .A4(n9249), .ZN(n9250) );
  OR4_X1 U11748 ( .A1(n13667), .A2(n13695), .A3(n13679), .A4(n9250), .ZN(n9251) );
  NOR2_X1 U11749 ( .A1(n13646), .A2(n9251), .ZN(n9252) );
  AND2_X1 U11750 ( .A1(n13617), .A2(n9252), .ZN(n9253) );
  AND4_X1 U11751 ( .A1(n13584), .A2(n9253), .A3(n13608), .A4(n13630), .ZN(
        n9255) );
  NAND4_X1 U11752 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n9284)
         );
  INV_X1 U11753 ( .A(n9840), .ZN(n9258) );
  AND2_X1 U11754 ( .A1(n9258), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9272) );
  AND2_X1 U11755 ( .A1(n9272), .A2(n11035), .ZN(n9271) );
  AND2_X1 U11756 ( .A1(n6587), .A2(n9271), .ZN(n9279) );
  INV_X1 U11757 ( .A(n9272), .ZN(n11427) );
  MUX2_X1 U11758 ( .A(n11035), .B(n6783), .S(n10920), .Z(n9259) );
  NOR2_X1 U11759 ( .A1(n11427), .A2(n9259), .ZN(n9260) );
  AND2_X1 U11760 ( .A1(n6587), .A2(n9260), .ZN(n9276) );
  AOI21_X1 U11761 ( .B1(n9284), .B2(n9279), .A(n9276), .ZN(n9261) );
  INV_X1 U11762 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11763 ( .A1(n9263), .A2(n9262), .ZN(n9288) );
  NAND2_X1 U11764 ( .A1(n9057), .A2(n13574), .ZN(n9267) );
  NAND2_X1 U11765 ( .A1(n9265), .A2(n9264), .ZN(n9266) );
  MUX2_X1 U11766 ( .A(n9267), .B(n9266), .S(n13575), .Z(n9278) );
  NAND2_X1 U11767 ( .A1(n10647), .A2(n6783), .ZN(n9268) );
  OAI211_X1 U11768 ( .C1(n6587), .C2(n11035), .A(n10181), .B(n9268), .ZN(n9269) );
  NAND2_X1 U11769 ( .A1(n13565), .A2(n9271), .ZN(n9283) );
  INV_X1 U11770 ( .A(n9278), .ZN(n9277) );
  INV_X1 U11771 ( .A(P2_B_REG_SCAN_IN), .ZN(n12992) );
  AOI21_X1 U11772 ( .B1(n9272), .B2(n6783), .A(n12992), .ZN(n9275) );
  INV_X1 U11773 ( .A(n10181), .ZN(n9273) );
  NAND4_X1 U11774 ( .A1(n9273), .A2(n9845), .A3(n13854), .A4(n15367), .ZN(
        n9274) );
  AOI22_X1 U11775 ( .A1(n9277), .A2(n9276), .B1(n9275), .B2(n9274), .ZN(n9282)
         );
  NAND2_X1 U11776 ( .A1(n9278), .A2(n10920), .ZN(n9280) );
  NAND3_X1 U11777 ( .A1(n9280), .A2(n9284), .A3(n9279), .ZN(n9281) );
  OAI211_X1 U11778 ( .C1(n9284), .C2(n9283), .A(n9282), .B(n9281), .ZN(n9285)
         );
  INV_X1 U11779 ( .A(n9285), .ZN(n9286) );
  NAND3_X1 U11780 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(P2_U3328) );
  NAND2_X1 U11781 ( .A1(n9290), .A2(n9289), .ZN(n11819) );
  NOR2_X1 U11782 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n11868), .ZN(n9292) );
  OAI22_X1 U11783 ( .A1(n11870), .A2(n14713), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11622) );
  INV_X1 U11784 ( .A(n11622), .ZN(n9293) );
  XNOR2_X1 U11785 ( .A(n11621), .B(n9293), .ZN(n13274) );
  NAND2_X1 U11786 ( .A1(n13274), .A2(n11633), .ZN(n9296) );
  NAND2_X1 U11787 ( .A1(n9294), .A2(SI_29_), .ZN(n9295) );
  INV_X1 U11788 ( .A(n12578), .ZN(n12448) );
  XNOR2_X1 U11789 ( .A(n11645), .B(n12448), .ZN(n11677) );
  INV_X1 U11790 ( .A(P3_B_REG_SCAN_IN), .ZN(n9297) );
  OR2_X1 U11791 ( .A1(n12302), .A2(n9297), .ZN(n9298) );
  NAND2_X1 U11792 ( .A1(n8165), .A2(n9298), .ZN(n14935) );
  NAND2_X1 U11793 ( .A1(n11636), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9303) );
  INV_X1 U11794 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9299) );
  OR2_X1 U11795 ( .A1(n11637), .A2(n9299), .ZN(n9302) );
  INV_X1 U11796 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n9300) );
  OR2_X1 U11797 ( .A1(n6570), .A2(n9300), .ZN(n9301) );
  NAND4_X1 U11798 ( .A1(n11643), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(
        n12577) );
  INV_X1 U11799 ( .A(n12577), .ZN(n11647) );
  INV_X1 U11800 ( .A(n9305), .ZN(n9306) );
  OAI21_X1 U11801 ( .B1(n9307), .B2(n15560), .A(n9306), .ZN(n12681) );
  AOI21_X1 U11802 ( .B1(n12685), .B2(n15600), .A(n12681), .ZN(n9313) );
  OR2_X1 U11803 ( .A1(n9313), .A2(n15612), .ZN(n9312) );
  INV_X1 U11804 ( .A(n13263), .ZN(n9310) );
  NOR2_X1 U11805 ( .A1(n15613), .A2(n9308), .ZN(n9309) );
  NAND2_X1 U11806 ( .A1(n9312), .A2(n9311), .ZN(P3_U3456) );
  OR2_X1 U11807 ( .A1(n9313), .A2(n15628), .ZN(n9318) );
  INV_X1 U11808 ( .A(n13211), .ZN(n9316) );
  INV_X1 U11809 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11810 ( .A1(n9318), .A2(n9317), .ZN(P3_U3488) );
  INV_X1 U11811 ( .A(n12594), .ZN(n11094) );
  OAI21_X1 U11812 ( .B1(n11682), .B2(n12673), .A(n10555), .ZN(n9320) );
  XNOR2_X1 U11813 ( .A(n10292), .B(n11281), .ZN(n9340) );
  XNOR2_X1 U11814 ( .A(n10292), .B(n15607), .ZN(n9338) );
  INV_X1 U11815 ( .A(n9338), .ZN(n9339) );
  INV_X1 U11816 ( .A(n12595), .ZN(n10927) );
  INV_X1 U11817 ( .A(n12598), .ZN(n11125) );
  XNOR2_X1 U11818 ( .A(n10292), .B(n15589), .ZN(n9333) );
  INV_X1 U11819 ( .A(n9333), .ZN(n9334) );
  XNOR2_X1 U11820 ( .A(n9328), .B(n10413), .ZN(n9330) );
  NAND3_X1 U11821 ( .A1(n6574), .A2(n9326), .A3(n11686), .ZN(n9322) );
  OAI21_X1 U11822 ( .B1(n11686), .B2(n9328), .A(n9322), .ZN(n9325) );
  NAND2_X1 U11823 ( .A1(n10294), .A2(n15554), .ZN(n9323) );
  XNOR2_X1 U11824 ( .A(n15550), .B(n9326), .ZN(n9327) );
  XNOR2_X1 U11825 ( .A(n9327), .B(n6822), .ZN(n15459) );
  XNOR2_X1 U11826 ( .A(n9328), .B(n15577), .ZN(n9329) );
  XNOR2_X1 U11827 ( .A(n9330), .B(n12600), .ZN(n10412) );
  XOR2_X1 U11828 ( .A(n12599), .B(n9331), .Z(n10545) );
  INV_X1 U11829 ( .A(n9331), .ZN(n9332) );
  XOR2_X1 U11830 ( .A(n12598), .B(n9333), .Z(n10607) );
  XNOR2_X1 U11831 ( .A(n11708), .B(n10292), .ZN(n10791) );
  INV_X1 U11832 ( .A(n12597), .ZN(n10928) );
  XNOR2_X1 U11833 ( .A(n10292), .B(n11721), .ZN(n9336) );
  XNOR2_X1 U11834 ( .A(n9336), .B(n12596), .ZN(n10923) );
  INV_X1 U11835 ( .A(n12596), .ZN(n11095) );
  XNOR2_X1 U11836 ( .A(n9338), .B(n12595), .ZN(n11081) );
  XOR2_X1 U11837 ( .A(n12594), .B(n9340), .Z(n11268) );
  XNOR2_X1 U11838 ( .A(n10292), .B(n11326), .ZN(n9341) );
  XNOR2_X1 U11839 ( .A(n11557), .B(n10292), .ZN(n9343) );
  INV_X1 U11840 ( .A(n11517), .ZN(n12592) );
  NAND2_X1 U11841 ( .A1(n9343), .A2(n12592), .ZN(n11505) );
  INV_X1 U11842 ( .A(n9343), .ZN(n9344) );
  NAND2_X1 U11843 ( .A1(n9344), .A2(n11517), .ZN(n11504) );
  XNOR2_X1 U11844 ( .A(n11908), .B(n10292), .ZN(n11900) );
  INV_X1 U11845 ( .A(n12457), .ZN(n9346) );
  XNOR2_X1 U11846 ( .A(n13260), .B(n10292), .ZN(n9347) );
  XNOR2_X1 U11847 ( .A(n9347), .B(n12590), .ZN(n12458) );
  INV_X1 U11848 ( .A(n12458), .ZN(n9345) );
  NAND2_X1 U11849 ( .A1(n9347), .A2(n12590), .ZN(n9348) );
  NAND2_X1 U11850 ( .A1(n12459), .A2(n9348), .ZN(n12565) );
  XNOR2_X1 U11851 ( .A(n12562), .B(n10292), .ZN(n9349) );
  XOR2_X1 U11852 ( .A(n11563), .B(n9349), .Z(n12564) );
  INV_X1 U11853 ( .A(n9349), .ZN(n9350) );
  NAND2_X1 U11854 ( .A1(n9350), .A2(n12848), .ZN(n9351) );
  XNOR2_X1 U11855 ( .A(n12505), .B(n10292), .ZN(n9352) );
  XOR2_X1 U11856 ( .A(n12567), .B(n9352), .Z(n12507) );
  INV_X1 U11857 ( .A(n9352), .ZN(n9353) );
  XNOR2_X1 U11858 ( .A(n12835), .B(n10292), .ZN(n9354) );
  NOR2_X1 U11859 ( .A1(n9354), .A2(n12509), .ZN(n12514) );
  XNOR2_X1 U11860 ( .A(n12910), .B(n10292), .ZN(n9355) );
  XNOR2_X1 U11861 ( .A(n9355), .B(n12517), .ZN(n11846) );
  INV_X1 U11862 ( .A(n9355), .ZN(n9356) );
  NAND2_X1 U11863 ( .A1(n9356), .A2(n12830), .ZN(n9357) );
  XNOR2_X1 U11864 ( .A(n13244), .B(n10292), .ZN(n9358) );
  XOR2_X1 U11865 ( .A(n12588), .B(n9358), .Z(n12476) );
  XNOR2_X1 U11866 ( .A(n13240), .B(n10292), .ZN(n9360) );
  XNOR2_X1 U11867 ( .A(n9360), .B(n12486), .ZN(n12536) );
  NAND2_X1 U11868 ( .A1(n9360), .A2(n12587), .ZN(n9361) );
  XNOR2_X1 U11869 ( .A(n12781), .B(n10292), .ZN(n9362) );
  NAND2_X1 U11870 ( .A1(n9362), .A2(n12546), .ZN(n9363) );
  OAI21_X1 U11871 ( .B1(n9362), .B2(n12546), .A(n9363), .ZN(n12484) );
  NAND2_X1 U11872 ( .A1(n12481), .A2(n9363), .ZN(n9367) );
  INV_X1 U11873 ( .A(n9367), .ZN(n9365) );
  XNOR2_X1 U11874 ( .A(n12768), .B(n10292), .ZN(n9366) );
  INV_X1 U11875 ( .A(n9366), .ZN(n9364) );
  NAND2_X1 U11876 ( .A1(n12543), .A2(n9368), .ZN(n9370) );
  XNOR2_X1 U11877 ( .A(n12757), .B(n10292), .ZN(n9369) );
  OAI21_X1 U11878 ( .B1(n9370), .B2(n9369), .A(n12527), .ZN(n12466) );
  INV_X1 U11879 ( .A(n12466), .ZN(n9375) );
  XNOR2_X1 U11880 ( .A(n12744), .B(n10292), .ZN(n9372) );
  NAND2_X1 U11881 ( .A1(n9372), .A2(n9371), .ZN(n12500) );
  INV_X1 U11882 ( .A(n9372), .ZN(n9373) );
  NAND2_X1 U11883 ( .A1(n9373), .A2(n12583), .ZN(n9374) );
  NAND2_X1 U11884 ( .A1(n12500), .A2(n9374), .ZN(n12528) );
  INV_X1 U11885 ( .A(n12527), .ZN(n9377) );
  XNOR2_X1 U11886 ( .A(n12727), .B(n10292), .ZN(n9379) );
  NAND2_X1 U11887 ( .A1(n9379), .A2(n12523), .ZN(n9382) );
  INV_X1 U11888 ( .A(n9379), .ZN(n9380) );
  NAND2_X1 U11889 ( .A1(n9380), .A2(n12582), .ZN(n9381) );
  AND2_X1 U11890 ( .A1(n9382), .A2(n9381), .ZN(n12499) );
  XNOR2_X1 U11891 ( .A(n12715), .B(n12440), .ZN(n9383) );
  NOR2_X1 U11892 ( .A1(n9383), .A2(n12581), .ZN(n9384) );
  AOI21_X1 U11893 ( .B1(n9383), .B2(n12581), .A(n9384), .ZN(n12555) );
  INV_X1 U11894 ( .A(n9384), .ZN(n9385) );
  NAND2_X1 U11895 ( .A1(n12554), .A2(n9385), .ZN(n9389) );
  INV_X1 U11896 ( .A(n9389), .ZN(n9387) );
  XNOR2_X1 U11897 ( .A(n12701), .B(n12440), .ZN(n12449) );
  NOR2_X1 U11898 ( .A1(n12449), .A2(n12580), .ZN(n12443) );
  AOI21_X1 U11899 ( .B1(n12449), .B2(n12580), .A(n12443), .ZN(n9388) );
  INV_X1 U11900 ( .A(n9388), .ZN(n9386) );
  NAND2_X1 U11901 ( .A1(n9387), .A2(n9386), .ZN(n9390) );
  NAND2_X1 U11902 ( .A1(n9390), .A2(n12455), .ZN(n9394) );
  NAND2_X1 U11903 ( .A1(n9396), .A2(n15606), .ZN(n9392) );
  OAI22_X1 U11904 ( .A1(n9397), .A2(n9392), .B1(n9404), .B2(n9391), .ZN(n9393)
         );
  NAND2_X1 U11905 ( .A1(n9394), .A2(n15469), .ZN(n9414) );
  NAND2_X1 U11906 ( .A1(n9397), .A2(n11833), .ZN(n9395) );
  INV_X1 U11907 ( .A(n12698), .ZN(n9410) );
  NAND2_X1 U11908 ( .A1(n9397), .A2(n9396), .ZN(n9400) );
  NAND2_X1 U11909 ( .A1(n9404), .A2(n9398), .ZN(n9399) );
  NAND4_X1 U11910 ( .A1(n9400), .A2(n9594), .A3(n9399), .A4(n10310), .ZN(n9402) );
  AND3_X1 U11911 ( .A1(n9404), .A2(n11839), .A3(n10221), .ZN(n9401) );
  AOI21_X1 U11912 ( .B1(n9402), .B2(P3_STATE_REG_SCAN_IN), .A(n9401), .ZN(
        n10152) );
  INV_X1 U11913 ( .A(n9403), .ZN(n9624) );
  NAND2_X1 U11914 ( .A1(n9624), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11843) );
  INV_X1 U11915 ( .A(n9404), .ZN(n9406) );
  AND2_X1 U11916 ( .A1(n11839), .A2(n11838), .ZN(n9405) );
  INV_X1 U11917 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9407) );
  OAI22_X1 U11918 ( .A1(n9408), .A2(n12571), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9407), .ZN(n9409) );
  AOI21_X1 U11919 ( .B1(n9410), .B2(n12573), .A(n9409), .ZN(n9411) );
  OAI21_X1 U11920 ( .B1(n13215), .B2(n12576), .A(n9411), .ZN(n9412) );
  NAND2_X1 U11921 ( .A1(n9414), .A2(n9413), .ZN(P3_U3154) );
  NOR2_X1 U11923 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n9422) );
  NOR2_X1 U11924 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9421) );
  NOR2_X1 U11925 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9420) );
  NAND2_X1 U11926 ( .A1(n9435), .A2(n9436), .ZN(n9433) );
  AND3_X1 U11927 ( .A1(n9544), .A2(n9428), .A3(n9535), .ZN(n9431) );
  NOR2_X1 U11928 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n9430) );
  NOR2_X1 U11929 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9429) );
  INV_X1 U11930 ( .A(n9435), .ZN(n9443) );
  INV_X1 U11931 ( .A(n9440), .ZN(n9441) );
  NAND2_X1 U11932 ( .A1(n9441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9442) );
  MUX2_X1 U11933 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9442), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9444) );
  INV_X1 U11934 ( .A(n9584), .ZN(n9732) );
  NOR2_X1 U11935 ( .A1(n10056), .A2(n9732), .ZN(P1_U4016) );
  NAND2_X1 U11936 ( .A1(n9448), .A2(n9449), .ZN(n14709) );
  INV_X1 U11937 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9447) );
  OR2_X1 U11938 ( .A1(n9448), .A2(n9447), .ZN(n9450) );
  NAND2_X1 U11939 ( .A1(n9511), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9457) );
  INV_X1 U11940 ( .A(n14714), .ZN(n9452) );
  NAND2_X1 U11941 ( .A1(n9451), .A2(n9452), .ZN(n9466) );
  INV_X2 U11942 ( .A(n9466), .ZN(n12092) );
  INV_X1 U11943 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U11944 ( .A1(n11871), .A2(n9452), .ZN(n9495) );
  INV_X1 U11945 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9760) );
  OR2_X1 U11946 ( .A1(n9495), .A2(n9760), .ZN(n9455) );
  INV_X1 U11947 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9453) );
  OR2_X1 U11948 ( .A1(n7654), .A2(n9453), .ZN(n9454) );
  NAND2_X1 U11949 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14721), .ZN(n9461) );
  MUX2_X1 U11950 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9461), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9464) );
  INV_X1 U11951 ( .A(n9462), .ZN(n9463) );
  NAND2_X1 U11952 ( .A1(n9464), .A2(n9463), .ZN(n14180) );
  INV_X1 U11953 ( .A(n14180), .ZN(n14177) );
  NAND2_X1 U11954 ( .A1(n11938), .A2(n10061), .ZN(n9548) );
  NAND2_X1 U11955 ( .A1(n12198), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9472) );
  INV_X1 U11956 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9465) );
  OR2_X1 U11957 ( .A1(n9466), .A2(n9465), .ZN(n9471) );
  INV_X1 U11958 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9467) );
  OR2_X1 U11959 ( .A1(n9494), .A2(n9467), .ZN(n9470) );
  INV_X1 U11960 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9468) );
  OR2_X1 U11961 ( .A1(n9495), .A2(n9468), .ZN(n9469) );
  OAI21_X1 U11962 ( .B1(n9680), .B2(n9474), .A(n9473), .ZN(n9475) );
  AND2_X1 U11963 ( .A1(n9476), .A2(n9475), .ZN(n14722) );
  MUX2_X1 U11964 ( .A(n14721), .B(n14722), .S(n11922), .Z(n10371) );
  AND2_X1 U11965 ( .A1(n14174), .A2(n10371), .ZN(n10454) );
  NAND2_X1 U11966 ( .A1(n12198), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9485) );
  INV_X1 U11967 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14194) );
  INV_X1 U11968 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9481) );
  OR2_X1 U11969 ( .A1(n9494), .A2(n9481), .ZN(n9483) );
  INV_X1 U11970 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9763) );
  OR2_X1 U11971 ( .A1(n9495), .A2(n9763), .ZN(n9482) );
  INV_X1 U11972 ( .A(n9707), .ZN(n9486) );
  INV_X1 U11973 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9708) );
  OR2_X1 U11974 ( .A1(n9462), .A2(n9447), .ZN(n9488) );
  XNOR2_X1 U11975 ( .A(n9488), .B(n9487), .ZN(n14197) );
  OAI22_X1 U11976 ( .A1(n11168), .A2(n9708), .B1(n11922), .B2(n14197), .ZN(
        n9489) );
  OR2_X2 U11977 ( .A1(n9490), .A2(n9489), .ZN(n15093) );
  OR2_X1 U11978 ( .A1(n14172), .A2(n15093), .ZN(n9491) );
  NAND2_X1 U11979 ( .A1(n12198), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9499) );
  INV_X2 U11980 ( .A(n12092), .ZN(n12202) );
  INV_X1 U11981 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9493) );
  OR2_X1 U11982 ( .A1(n9494), .A2(n9493), .ZN(n9497) );
  INV_X2 U11983 ( .A(n9522), .ZN(n11348) );
  INV_X1 U11984 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9759) );
  INV_X1 U11985 ( .A(n14171), .ZN(n9505) );
  NOR2_X1 U11986 ( .A1(n9502), .A2(n9447), .ZN(n9500) );
  MUX2_X1 U11987 ( .A(n9447), .B(n9500), .S(P1_IR_REG_3__SCAN_IN), .Z(n9503)
         );
  AND2_X1 U11988 ( .A1(n9502), .A2(n9501), .ZN(n9507) );
  NOR2_X1 U11989 ( .A1(n9503), .A2(n9507), .ZN(n14214) );
  AOI22_X1 U11990 ( .A1(n12223), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n12066), 
        .B2(n14214), .ZN(n9504) );
  NAND2_X1 U11991 ( .A1(n9505), .A2(n15155), .ZN(n9506) );
  OR2_X1 U11992 ( .A1(n9683), .A2(n12123), .ZN(n9510) );
  INV_X1 U11993 ( .A(n9507), .ZN(n9518) );
  NAND2_X1 U11994 ( .A1(n9518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9508) );
  XNOR2_X1 U11995 ( .A(n9508), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U11996 ( .A1(n12223), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12066), 
        .B2(n14228), .ZN(n9509) );
  NAND2_X1 U11997 ( .A1(n12218), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9515) );
  INV_X1 U11998 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10366) );
  OR2_X1 U11999 ( .A1(n12219), .A2(n10366), .ZN(n9514) );
  NAND2_X1 U12000 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9524) );
  OAI21_X1 U12001 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9524), .ZN(n10544) );
  OR2_X1 U12002 ( .A1(n12202), .A2(n10544), .ZN(n9513) );
  INV_X1 U12003 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9768) );
  OR2_X1 U12004 ( .A1(n11348), .A2(n9768), .ZN(n9512) );
  INV_X1 U12005 ( .A(n11960), .ZN(n14170) );
  NAND2_X1 U12006 ( .A1(n11961), .A2(n14170), .ZN(n9516) );
  NAND2_X1 U12007 ( .A1(n9517), .A2(n9516), .ZN(n9533) );
  INV_X1 U12008 ( .A(n9533), .ZN(n9532) );
  NAND2_X1 U12009 ( .A1(n9685), .A2(n12234), .ZN(n9521) );
  NAND2_X1 U12010 ( .A1(n9691), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U12011 ( .A(n9519), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U12012 ( .A1(n12223), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12066), 
        .B2(n9824), .ZN(n9520) );
  NAND2_X1 U12013 ( .A1(n9521), .A2(n9520), .ZN(n11964) );
  NAND2_X1 U12014 ( .A1(n12198), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9530) );
  INV_X1 U12015 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9772) );
  OR2_X1 U12016 ( .A1(n11348), .A2(n9772), .ZN(n9529) );
  INV_X1 U12017 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9523) );
  AND2_X1 U12018 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  NOR2_X1 U12019 ( .A1(n9524), .A2(n9523), .ZN(n9555) );
  OR2_X1 U12020 ( .A1(n9525), .A2(n9555), .ZN(n10601) );
  OR2_X1 U12021 ( .A1(n12202), .A2(n10601), .ZN(n9528) );
  INV_X1 U12022 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9526) );
  OR2_X1 U12023 ( .A1(n12219), .A2(n9526), .ZN(n9527) );
  INV_X1 U12024 ( .A(n14169), .ZN(n10594) );
  NAND2_X1 U12025 ( .A1(n11964), .A2(n10594), .ZN(n10458) );
  OR2_X1 U12026 ( .A1(n11964), .A2(n10594), .ZN(n9531) );
  NAND2_X1 U12027 ( .A1(n9533), .A2(n6864), .ZN(n9534) );
  NAND2_X1 U12028 ( .A1(n10473), .A2(n9534), .ZN(n10381) );
  NAND2_X1 U12029 ( .A1(n7637), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9538) );
  OR2_X1 U12030 ( .A1(n10032), .A2(n11924), .ZN(n9546) );
  NAND2_X1 U12031 ( .A1(n11924), .A2(n10032), .ZN(n12303) );
  NAND2_X1 U12032 ( .A1(n10362), .A2(n9547), .ZN(n10911) );
  NAND2_X1 U12033 ( .A1(n10381), .A2(n15084), .ZN(n9566) );
  INV_X1 U12034 ( .A(n10371), .ZN(n15135) );
  NAND2_X1 U12035 ( .A1(n9548), .A2(n11934), .ZN(n11928) );
  NAND2_X1 U12036 ( .A1(n11928), .A2(n11942), .ZN(n15079) );
  OR2_X1 U12037 ( .A1(n14172), .A2(n15148), .ZN(n11946) );
  NOR2_X1 U12038 ( .A1(n14170), .A2(n11959), .ZN(n9549) );
  NAND2_X1 U12039 ( .A1(n9550), .A2(n12256), .ZN(n9551) );
  NAND2_X1 U12040 ( .A1(n10459), .A2(n9551), .ZN(n9564) );
  NAND2_X1 U12041 ( .A1(n14445), .A2(n15133), .ZN(n9553) );
  INV_X1 U12042 ( .A(n12222), .ZN(n9587) );
  NAND2_X1 U12043 ( .A1(n15134), .A2(n9587), .ZN(n9552) );
  INV_X1 U12044 ( .A(n11866), .ZN(n14190) );
  OR2_X1 U12045 ( .A1(n11960), .A2(n14591), .ZN(n9562) );
  NAND2_X1 U12046 ( .A1(n12218), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9560) );
  INV_X1 U12047 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9791) );
  OR2_X1 U12048 ( .A1(n12219), .A2(n9791), .ZN(n9559) );
  NAND2_X1 U12049 ( .A1(n9555), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10465) );
  OR2_X1 U12050 ( .A1(n9555), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12051 ( .A1(n10465), .A2(n9556), .ZN(n10477) );
  OR2_X1 U12052 ( .A1(n12202), .A2(n10477), .ZN(n9558) );
  INV_X1 U12053 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9774) );
  OR2_X1 U12054 ( .A1(n11348), .A2(n9774), .ZN(n9557) );
  NAND4_X1 U12055 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n14168) );
  NAND2_X1 U12056 ( .A1(n14168), .A2(n14570), .ZN(n9561) );
  AND2_X1 U12057 ( .A1(n9562), .A2(n9561), .ZN(n10600) );
  INV_X1 U12058 ( .A(n10600), .ZN(n9563) );
  AOI21_X1 U12059 ( .B1(n9564), .B2(n6917), .A(n9563), .ZN(n9565) );
  NAND2_X1 U12060 ( .A1(n9566), .A2(n9565), .ZN(n10379) );
  NAND2_X1 U12061 ( .A1(n12425), .A2(P1_B_REG_SCAN_IN), .ZN(n9567) );
  MUX2_X1 U12062 ( .A(P1_B_REG_SCAN_IN), .B(n9567), .S(n11617), .Z(n9568) );
  OR2_X1 U12063 ( .A1(n9731), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U12064 ( .A1(n12298), .A2(n11617), .ZN(n9569) );
  INV_X1 U12065 ( .A(n10122), .ZN(n10110) );
  OR2_X1 U12066 ( .A1(n9731), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U12067 ( .A1(n12298), .A2(n12425), .ZN(n9571) );
  AND2_X1 U12068 ( .A1(n9572), .A2(n9571), .ZN(n10109) );
  NOR4_X1 U12069 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9576) );
  NOR4_X1 U12070 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9575) );
  NOR4_X1 U12071 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9574) );
  NOR4_X1 U12072 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9573) );
  NAND4_X1 U12073 ( .A1(n9576), .A2(n9575), .A3(n9574), .A4(n9573), .ZN(n9582)
         );
  NOR2_X1 U12074 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n9580) );
  NOR4_X1 U12075 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9579) );
  NOR4_X1 U12076 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9578) );
  NOR4_X1 U12077 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9577) );
  NAND4_X1 U12078 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n9581)
         );
  NOR2_X1 U12079 ( .A1(n9582), .A2(n9581), .ZN(n9583) );
  OR2_X1 U12080 ( .A1(n9731), .A2(n9583), .ZN(n10049) );
  AND2_X1 U12081 ( .A1(n10049), .A2(n10052), .ZN(n10041) );
  NAND2_X1 U12082 ( .A1(n9547), .A2(n12222), .ZN(n9585) );
  NAND2_X1 U12083 ( .A1(n9585), .A2(n12237), .ZN(n10054) );
  INV_X1 U12084 ( .A(n10050), .ZN(n10108) );
  MUX2_X1 U12085 ( .A(n10379), .B(P1_REG2_REG_5__SCAN_IN), .S(n15098), .Z(
        n9591) );
  NAND2_X1 U12086 ( .A1(n14445), .A2(n11929), .ZN(n12239) );
  INV_X1 U12087 ( .A(n10918), .ZN(n15095) );
  AND2_X1 U12088 ( .A1(n10381), .A2(n15095), .ZN(n9590) );
  NAND2_X1 U12089 ( .A1(n6575), .A2(n15135), .ZN(n15092) );
  NOR2_X1 U12090 ( .A1(n15092), .A2(n15093), .ZN(n15090) );
  AND2_X1 U12091 ( .A1(n15090), .A2(n15155), .ZN(n10286) );
  INV_X1 U12092 ( .A(n11964), .ZN(n10593) );
  OAI211_X1 U12093 ( .C1(n10117), .C2(n10593), .A(n14538), .B(n10476), .ZN(
        n10378) );
  NOR2_X1 U12094 ( .A1(n14543), .A2(n10378), .ZN(n9589) );
  AND2_X1 U12095 ( .A1(n11925), .A2(n9587), .ZN(n12244) );
  NAND2_X1 U12096 ( .A1(n12244), .A2(n10042), .ZN(n10043) );
  OAI22_X1 U12097 ( .A1(n15088), .A2(n10593), .B1(n10601), .B2(n14556), .ZN(
        n9588) );
  INV_X1 U12098 ( .A(n9592), .ZN(n9593) );
  NAND2_X1 U12099 ( .A1(n9593), .A2(n9840), .ZN(n9842) );
  MUX2_X1 U12100 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13279), .Z(n9595) );
  XNOR2_X1 U12101 ( .A(n9595), .B(n6590), .ZN(n10235) );
  MUX2_X1 U12102 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13279), .Z(n10356) );
  NAND2_X1 U12103 ( .A1(n10235), .A2(n10355), .ZN(n9598) );
  INV_X1 U12104 ( .A(n9595), .ZN(n9596) );
  NAND2_X1 U12105 ( .A1(n9596), .A2(n6590), .ZN(n9597) );
  NAND2_X1 U12106 ( .A1(n9598), .A2(n9597), .ZN(n10146) );
  MUX2_X1 U12107 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13279), .Z(n9599) );
  XNOR2_X1 U12108 ( .A(n9599), .B(n6572), .ZN(n10145) );
  NAND2_X1 U12109 ( .A1(n10146), .A2(n10145), .ZN(n9602) );
  INV_X1 U12110 ( .A(n9599), .ZN(n9600) );
  NAND2_X1 U12111 ( .A1(n9600), .A2(n6572), .ZN(n9601) );
  NAND2_X1 U12112 ( .A1(n9602), .A2(n9601), .ZN(n15481) );
  MUX2_X1 U12113 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13279), .Z(n9604) );
  XNOR2_X1 U12114 ( .A(n9604), .B(n9603), .ZN(n15480) );
  NOR2_X1 U12115 ( .A1(n9604), .A2(n15485), .ZN(n9605) );
  AOI21_X1 U12116 ( .B1(n15481), .B2(n15480), .A(n9605), .ZN(n15491) );
  MUX2_X1 U12117 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13279), .Z(n9606) );
  XNOR2_X1 U12118 ( .A(n9606), .B(n15504), .ZN(n15490) );
  MUX2_X1 U12119 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13279), .Z(n9607) );
  NAND2_X1 U12120 ( .A1(n9607), .A2(n15512), .ZN(n15508) );
  NAND2_X1 U12121 ( .A1(n15510), .A2(n15508), .ZN(n9613) );
  INV_X1 U12122 ( .A(n9607), .ZN(n9608) );
  NAND2_X1 U12123 ( .A1(n9608), .A2(n9636), .ZN(n15509) );
  INV_X1 U12124 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10206) );
  MUX2_X1 U12125 ( .A(n10190), .B(n10206), .S(n13279), .Z(n9609) );
  NAND2_X1 U12126 ( .A1(n9609), .A2(n10207), .ZN(n10195) );
  INV_X1 U12127 ( .A(n9609), .ZN(n9610) );
  INV_X1 U12128 ( .A(n10207), .ZN(n9679) );
  NAND2_X1 U12129 ( .A1(n9610), .A2(n9679), .ZN(n9611) );
  NAND2_X1 U12130 ( .A1(n10195), .A2(n9611), .ZN(n9612) );
  INV_X1 U12131 ( .A(n10203), .ZN(n9615) );
  NAND3_X1 U12132 ( .A1(n9613), .A2(n15509), .A3(n9612), .ZN(n9614) );
  AOI21_X1 U12133 ( .B1(n9615), .B2(n9614), .A(n14920), .ZN(n9649) );
  XNOR2_X1 U12134 ( .A(n6571), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U12135 ( .A1(n9616), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12136 ( .A1(n10244), .A2(n10352), .ZN(n9617) );
  NAND2_X1 U12137 ( .A1(n9617), .A2(n6599), .ZN(n10238) );
  INV_X1 U12138 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U12139 ( .A1(n10240), .A2(n6599), .ZN(n10138) );
  NAND2_X1 U12140 ( .A1(n10139), .A2(n10138), .ZN(n10141) );
  INV_X1 U12141 ( .A(n6572), .ZN(n10150) );
  NAND2_X1 U12142 ( .A1(n10150), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12143 ( .A1(n10141), .A2(n9618), .ZN(n9619) );
  NOR2_X1 U12144 ( .A1(n9636), .A2(n9620), .ZN(n9621) );
  AOI22_X1 U12145 ( .A1(n10207), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10190), 
        .B2(n9679), .ZN(n9622) );
  AOI21_X1 U12146 ( .B1(n6731), .B2(n9622), .A(n10192), .ZN(n9628) );
  INV_X1 U12147 ( .A(n11839), .ZN(n9623) );
  NAND2_X1 U12148 ( .A1(n9623), .A2(n11843), .ZN(n9643) );
  OR2_X1 U12149 ( .A1(n8226), .A2(n9624), .ZN(n9626) );
  AND2_X1 U12150 ( .A1(n9626), .A2(n9625), .ZN(n9641) );
  NAND2_X1 U12151 ( .A1(n9643), .A2(n9641), .ZN(n9640) );
  NOR2_X1 U12152 ( .A1(n9628), .A2(n15547), .ZN(n9648) );
  INV_X1 U12153 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15616) );
  INV_X1 U12154 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10347) );
  INV_X1 U12155 ( .A(n9630), .ZN(n9632) );
  NAND2_X1 U12156 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9630), .ZN(n9631) );
  OAI21_X1 U12157 ( .B1(n6590), .B2(n9630), .A(n9631), .ZN(n10237) );
  NAND2_X1 U12158 ( .A1(n10237), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U12159 ( .A1(n10236), .A2(n7647), .ZN(n10134) );
  NAND2_X1 U12160 ( .A1(n10150), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9633) );
  INV_X1 U12161 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15618) );
  INV_X1 U12162 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15620) );
  NOR2_X1 U12163 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  NOR2_X1 U12164 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  INV_X1 U12165 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U12166 ( .A1(n10207), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n10206), 
        .B2(n9679), .ZN(n9638) );
  AOI21_X1 U12167 ( .B1(n6730), .B2(n9638), .A(n10209), .ZN(n9639) );
  NOR2_X1 U12168 ( .A1(n9639), .A2(n15541), .ZN(n9647) );
  INV_X1 U12169 ( .A(n9641), .ZN(n9642) );
  INV_X1 U12170 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U12171 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10609), .ZN(n9644) );
  AOI21_X1 U12172 ( .B1(n15458), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n9644), .ZN(
        n9645) );
  OAI21_X1 U12173 ( .B1(n15531), .B2(n9679), .A(n9645), .ZN(n9646) );
  OR4_X1 U12174 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(P3_U3188) );
  AOI211_X1 U12175 ( .C1(n9652), .C2(n9650), .A(n12552), .B(n9651), .ZN(n9656)
         );
  INV_X1 U12176 ( .A(n12573), .ZN(n12549) );
  INV_X1 U12177 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10998) );
  NOR2_X1 U12178 ( .A1(n12549), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9655) );
  OAI22_X1 U12179 ( .A1(n12576), .A2(n15577), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10998), .ZN(n9654) );
  INV_X1 U12180 ( .A(n6822), .ZN(n10737) );
  INV_X1 U12181 ( .A(n8165), .ZN(n15563) );
  OR2_X1 U12182 ( .A1(n12571), .A2(n15563), .ZN(n15467) );
  OAI22_X1 U12183 ( .A1(n10737), .A2(n11083), .B1(n15467), .B2(n7247), .ZN(
        n9653) );
  OR4_X1 U12184 ( .A1(n9656), .A2(n9655), .A3(n9654), .A4(n9653), .ZN(P3_U3158) );
  OAI21_X1 U12185 ( .B1(n9658), .B2(P3_STATE_REG_SCAN_IN), .A(n9657), .ZN(
        P3_U3295) );
  NAND2_X2 U12186 ( .A1(n9680), .A2(P2_U3088), .ZN(n14022) );
  OAI222_X1 U12187 ( .A1(n14024), .A2(n9659), .B1(n14022), .B2(n9709), .C1(
        P2_U3088), .C2(n15228), .ZN(P2_U3326) );
  OAI222_X1 U12188 ( .A1(n14024), .A2(n9660), .B1(n14022), .B2(n9702), .C1(
        P2_U3088), .C2(n9984), .ZN(P2_U3324) );
  OAI222_X1 U12189 ( .A1(n14024), .A2(n9661), .B1(n14022), .B2(n9707), .C1(
        P2_U3088), .C2(n9878), .ZN(P2_U3325) );
  OAI222_X1 U12190 ( .A1(n14024), .A2(n9662), .B1(n14022), .B2(n9683), .C1(
        P2_U3088), .C2(n9955), .ZN(P2_U3323) );
  INV_X1 U12191 ( .A(n14835), .ZN(n13282) );
  OAI222_X1 U12192 ( .A1(n13282), .A2(n9664), .B1(n13284), .B2(n9663), .C1(
        n10212), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12193 ( .A(n9665), .ZN(n9666) );
  OAI222_X1 U12194 ( .A1(P3_U3151), .A2(n7137), .B1(n13284), .B2(n9667), .C1(
        n13282), .C2(n9666), .ZN(P3_U3294) );
  OAI222_X1 U12195 ( .A1(n13282), .A2(n9669), .B1(n13284), .B2(n9668), .C1(
        n10945), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12196 ( .A1(n13282), .A2(n9671), .B1(n13284), .B2(n9670), .C1(
        n10441), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12197 ( .A1(n15485), .A2(P3_U3151), .B1(n13282), .B2(n9673), .C1(
        n9672), .C2(n13284), .ZN(P3_U3292) );
  OAI222_X1 U12198 ( .A1(n10150), .A2(P3_U3151), .B1(n13282), .B2(n9675), .C1(
        n9674), .C2(n13284), .ZN(P3_U3293) );
  INV_X1 U12199 ( .A(n9676), .ZN(n9678) );
  INV_X1 U12200 ( .A(SI_6_), .ZN(n9677) );
  OAI222_X1 U12201 ( .A1(n9679), .A2(P3_U3151), .B1(n13282), .B2(n9678), .C1(
        n9677), .C2(n13284), .ZN(P3_U3289) );
  INV_X1 U12202 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9684) );
  INV_X1 U12203 ( .A(n14228), .ZN(n9682) );
  OAI222_X1 U12204 ( .A1(n12296), .A2(n9684), .B1(n12426), .B2(n9683), .C1(
        P1_U3086), .C2(n9682), .ZN(P1_U3351) );
  INV_X1 U12205 ( .A(n9685), .ZN(n9699) );
  INV_X1 U12206 ( .A(n9851), .ZN(n9941) );
  OAI222_X1 U12207 ( .A1(n14024), .A2(n9686), .B1(n14022), .B2(n9699), .C1(
        P2_U3088), .C2(n9941), .ZN(P2_U3322) );
  INV_X1 U12208 ( .A(n10460), .ZN(n9696) );
  INV_X1 U12209 ( .A(n9852), .ZN(n15241) );
  OAI222_X1 U12210 ( .A1(n14024), .A2(n9687), .B1(n14022), .B2(n9696), .C1(
        P2_U3088), .C2(n15241), .ZN(P2_U3321) );
  INV_X1 U12211 ( .A(n9688), .ZN(n9690) );
  INV_X1 U12212 ( .A(n11068), .ZN(n12616) );
  OAI222_X1 U12213 ( .A1(n13282), .A2(n9690), .B1(n13284), .B2(n9689), .C1(
        n12616), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12214 ( .A(n9691), .ZN(n9693) );
  NAND2_X1 U12215 ( .A1(n9693), .A2(n9692), .ZN(n9704) );
  NAND2_X1 U12216 ( .A1(n9704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9694) );
  XNOR2_X1 U12217 ( .A(n9694), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14245) );
  INV_X1 U12218 ( .A(n14245), .ZN(n9695) );
  OAI222_X1 U12219 ( .A1(n12296), .A2(n9697), .B1(n12426), .B2(n9696), .C1(
        P1_U3086), .C2(n9695), .ZN(P1_U3349) );
  INV_X1 U12220 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9700) );
  INV_X1 U12221 ( .A(n9824), .ZN(n9698) );
  OAI222_X1 U12222 ( .A1(n12296), .A2(n9700), .B1(n12426), .B2(n9699), .C1(
        P1_U3086), .C2(n9698), .ZN(P1_U3350) );
  INV_X1 U12223 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9703) );
  INV_X1 U12224 ( .A(n14214), .ZN(n9701) );
  OAI222_X1 U12225 ( .A1(n12296), .A2(n9703), .B1(n12426), .B2(n9702), .C1(
        P1_U3086), .C2(n9701), .ZN(P1_U3352) );
  INV_X1 U12226 ( .A(n10490), .ZN(n9712) );
  OAI21_X1 U12227 ( .B1(n9704), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9705) );
  XNOR2_X1 U12228 ( .A(n9705), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14258) );
  INV_X1 U12229 ( .A(n12296), .ZN(n14717) );
  AOI22_X1 U12230 ( .A1(n14258), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14717), .ZN(n9706) );
  OAI21_X1 U12231 ( .B1(n9712), .B2(n12426), .A(n9706), .ZN(P1_U3348) );
  OAI222_X1 U12232 ( .A1(n12296), .A2(n9708), .B1(n12426), .B2(n9707), .C1(
        P1_U3086), .C2(n14197), .ZN(P1_U3353) );
  OAI222_X1 U12233 ( .A1(n12296), .A2(n9710), .B1(n12426), .B2(n9709), .C1(
        P1_U3086), .C2(n14180), .ZN(P1_U3354) );
  INV_X1 U12234 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9713) );
  INV_X1 U12235 ( .A(n9895), .ZN(n9711) );
  OAI222_X1 U12236 ( .A1(n14024), .A2(n9713), .B1(n14022), .B2(n9712), .C1(
        P2_U3088), .C2(n9711), .ZN(P2_U3320) );
  INV_X1 U12237 ( .A(n10495), .ZN(n9720) );
  NOR2_X1 U12238 ( .A1(n9714), .A2(n9447), .ZN(n9715) );
  MUX2_X1 U12239 ( .A(n9447), .B(n9715), .S(P1_IR_REG_8__SCAN_IN), .Z(n9718)
         );
  INV_X1 U12240 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U12241 ( .A1(n9714), .A2(n9716), .ZN(n9738) );
  INV_X1 U12242 ( .A(n9738), .ZN(n9717) );
  NOR2_X1 U12243 ( .A1(n9718), .A2(n9717), .ZN(n10496) );
  INV_X1 U12244 ( .A(n10496), .ZN(n9783) );
  OAI222_X1 U12245 ( .A1(n12296), .A2(n9719), .B1(n12426), .B2(n9720), .C1(
        P1_U3086), .C2(n9783), .ZN(P1_U3347) );
  INV_X1 U12246 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9721) );
  INV_X1 U12247 ( .A(n9853), .ZN(n9970) );
  OAI222_X1 U12248 ( .A1(n14024), .A2(n9721), .B1(n14022), .B2(n9720), .C1(
        P2_U3088), .C2(n9970), .ZN(P2_U3319) );
  INV_X1 U12249 ( .A(n10052), .ZN(n9722) );
  OR2_X1 U12250 ( .A1(n10053), .A2(P1_U3086), .ZN(n12293) );
  NAND2_X1 U12251 ( .A1(n9722), .A2(n12293), .ZN(n9726) );
  NAND2_X1 U12252 ( .A1(n10053), .A2(n12237), .ZN(n9723) );
  NAND2_X1 U12253 ( .A1(n9723), .A2(n11922), .ZN(n9724) );
  INV_X1 U12254 ( .A(n9724), .ZN(n9725) );
  NAND2_X1 U12255 ( .A1(n9726), .A2(n9725), .ZN(n9782) );
  INV_X1 U12256 ( .A(n9782), .ZN(n9796) );
  INV_X1 U12257 ( .A(n14187), .ZN(n14333) );
  NOR2_X1 U12258 ( .A1(n14187), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U12259 ( .A1(n9727), .A2(n11866), .ZN(n14193) );
  OAI21_X1 U12260 ( .B1(n14333), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14193), .ZN(
        n9728) );
  XNOR2_X1 U12261 ( .A(n9728), .B(n14721), .ZN(n9729) );
  AOI22_X1 U12262 ( .A1(n9796), .A2(n9729), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9730) );
  OAI21_X1 U12263 ( .B1(n6918), .B2(n15075), .A(n9730), .ZN(P1_U3243) );
  OR2_X1 U12264 ( .A1(n6818), .A2(n9732), .ZN(n9734) );
  OAI22_X1 U12265 ( .A1(n15129), .A2(P1_D_REG_1__SCAN_IN), .B1(n9439), .B2(
        n9734), .ZN(n9733) );
  INV_X1 U12266 ( .A(n9733), .ZN(P1_U3446) );
  OAI22_X1 U12267 ( .A1(n15129), .A2(P1_D_REG_0__SCAN_IN), .B1(n9438), .B2(
        n9734), .ZN(n9735) );
  INV_X1 U12268 ( .A(n9735), .ZN(P1_U3445) );
  INV_X1 U12269 ( .A(n15075), .ZN(n14269) );
  NOR2_X1 U12270 ( .A1(n14269), .A2(n6576), .ZN(P1_U3085) );
  INV_X1 U12271 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U12272 ( .A1(n13574), .A2(P2_U3947), .ZN(n9736) );
  OAI21_X1 U12273 ( .B1(P2_U3947), .B2(n11629), .A(n9736), .ZN(P2_U3562) );
  INV_X1 U12274 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9737) );
  INV_X1 U12275 ( .A(n10800), .ZN(n9742) );
  INV_X1 U12276 ( .A(n10012), .ZN(n9870) );
  OAI222_X1 U12277 ( .A1(n14024), .A2(n9737), .B1(n14022), .B2(n9742), .C1(
        P2_U3088), .C2(n9870), .ZN(P2_U3318) );
  NOR2_X1 U12278 ( .A1(n9738), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9755) );
  INV_X1 U12279 ( .A(n9755), .ZN(n9741) );
  NAND2_X1 U12280 ( .A1(n9738), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U12281 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9739), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9740) );
  INV_X1 U12282 ( .A(n10801), .ZN(n10085) );
  OAI222_X1 U12283 ( .A1(n12296), .A2(n9743), .B1(n12426), .B2(n9742), .C1(
        P1_U3086), .C2(n10085), .ZN(P1_U3346) );
  INV_X1 U12284 ( .A(n12619), .ZN(n15530) );
  INV_X1 U12285 ( .A(n9744), .ZN(n9746) );
  OAI222_X1 U12286 ( .A1(n15530), .A2(P3_U3151), .B1(n13282), .B2(n9746), .C1(
        n9745), .C2(n13284), .ZN(P3_U3282) );
  INV_X1 U12287 ( .A(n10806), .ZN(n9751) );
  OR2_X1 U12288 ( .A1(n9755), .A2(n9447), .ZN(n9747) );
  XNOR2_X1 U12289 ( .A(n9747), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14273) );
  AOI22_X1 U12290 ( .A1(n14273), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14717), .ZN(n9748) );
  OAI21_X1 U12291 ( .B1(n9751), .B2(n12426), .A(n9748), .ZN(P1_U3345) );
  OAI222_X1 U12292 ( .A1(n13282), .A2(n9750), .B1(n13284), .B2(n9749), .C1(
        n12648), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12293 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9752) );
  INV_X1 U12294 ( .A(n11005), .ZN(n11018) );
  OAI222_X1 U12295 ( .A1(n14024), .A2(n9752), .B1(n14022), .B2(n9751), .C1(
        P2_U3088), .C2(n11018), .ZN(P2_U3317) );
  INV_X1 U12296 ( .A(n10953), .ZN(n9757) );
  INV_X1 U12297 ( .A(n11019), .ZN(n13522) );
  OAI222_X1 U12298 ( .A1(n14024), .A2(n9753), .B1(n14022), .B2(n9757), .C1(
        P2_U3088), .C2(n13522), .ZN(P2_U3316) );
  INV_X1 U12299 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U12300 ( .A1(n9755), .A2(n9754), .ZN(n9985) );
  NAND2_X1 U12301 ( .A1(n9985), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9756) );
  XNOR2_X1 U12302 ( .A(n9756), .B(P1_IR_REG_11__SCAN_IN), .ZN(n15037) );
  INV_X1 U12303 ( .A(n15037), .ZN(n10089) );
  OAI222_X1 U12304 ( .A1(n12296), .A2(n9758), .B1(n12426), .B2(n9757), .C1(
        P1_U3086), .C2(n10089), .ZN(P1_U3344) );
  INV_X1 U12305 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10499) );
  MUX2_X1 U12306 ( .A(n10499), .B(P1_REG1_REG_8__SCAN_IN), .S(n10496), .Z(
        n9781) );
  MUX2_X1 U12307 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9759), .S(n14214), .Z(n9767) );
  MUX2_X1 U12308 ( .A(n9760), .B(P1_REG1_REG_1__SCAN_IN), .S(n14180), .Z(n9762) );
  AND2_X1 U12309 ( .A1(n14721), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12310 ( .A1(n9762), .A2(n9761), .ZN(n14200) );
  NAND2_X1 U12311 ( .A1(n14177), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U12312 ( .A1(n14200), .A2(n14199), .ZN(n9765) );
  MUX2_X1 U12313 ( .A(n9763), .B(P1_REG1_REG_2__SCAN_IN), .S(n14197), .Z(n9764) );
  NAND2_X1 U12314 ( .A1(n9765), .A2(n9764), .ZN(n14216) );
  INV_X1 U12315 ( .A(n14197), .ZN(n14196) );
  NAND2_X1 U12316 ( .A1(n14196), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14215) );
  NAND2_X1 U12317 ( .A1(n14216), .A2(n14215), .ZN(n9766) );
  NAND2_X1 U12318 ( .A1(n9767), .A2(n9766), .ZN(n14231) );
  NAND2_X1 U12319 ( .A1(n14214), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14230) );
  NAND2_X1 U12320 ( .A1(n14231), .A2(n14230), .ZN(n9770) );
  MUX2_X1 U12321 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9768), .S(n14228), .Z(n9769) );
  NAND2_X1 U12322 ( .A1(n9770), .A2(n9769), .ZN(n14233) );
  NAND2_X1 U12323 ( .A1(n14228), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U12324 ( .A1(n14233), .A2(n9771), .ZN(n9820) );
  MUX2_X1 U12325 ( .A(n9772), .B(P1_REG1_REG_5__SCAN_IN), .S(n9824), .Z(n9821)
         );
  OR2_X1 U12326 ( .A1(n9820), .A2(n9821), .ZN(n9818) );
  OR2_X1 U12327 ( .A1(n9824), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9773) );
  AND2_X1 U12328 ( .A1(n9818), .A2(n9773), .ZN(n14239) );
  MUX2_X1 U12329 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9774), .S(n14245), .Z(
        n14238) );
  NAND2_X1 U12330 ( .A1(n14239), .A2(n14238), .ZN(n14255) );
  NAND2_X1 U12331 ( .A1(n14245), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U12332 ( .A1(n14255), .A2(n14254), .ZN(n9777) );
  INV_X1 U12333 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9775) );
  MUX2_X1 U12334 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9775), .S(n14258), .Z(n9776) );
  NAND2_X1 U12335 ( .A1(n9777), .A2(n9776), .ZN(n14257) );
  NAND2_X1 U12336 ( .A1(n14258), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12337 ( .A1(n14257), .A2(n9778), .ZN(n9780) );
  OR2_X1 U12338 ( .A1(n9780), .A2(n9781), .ZN(n9806) );
  INV_X1 U12339 ( .A(n9806), .ZN(n9779) );
  AOI21_X1 U12340 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9801) );
  AND2_X1 U12341 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9785) );
  OR2_X1 U12342 ( .A1(n9782), .A2(n14190), .ZN(n14320) );
  NOR2_X1 U12343 ( .A1(n14320), .A2(n9783), .ZN(n9784) );
  AOI211_X1 U12344 ( .C1(n14269), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9785), .B(
        n9784), .ZN(n9800) );
  INV_X1 U12345 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10503) );
  XNOR2_X1 U12346 ( .A(n10496), .B(n10503), .ZN(n9798) );
  MUX2_X1 U12347 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9493), .S(n14214), .Z(
        n14213) );
  XNOR2_X1 U12348 ( .A(n14180), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14179) );
  AND2_X1 U12349 ( .A1(n14721), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U12350 ( .A1(n14179), .A2(n14189), .ZN(n14178) );
  NAND2_X1 U12351 ( .A1(n14177), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U12352 ( .A1(n14178), .A2(n9786), .ZN(n14203) );
  MUX2_X1 U12353 ( .A(n9481), .B(P1_REG2_REG_2__SCAN_IN), .S(n14197), .Z(
        n14204) );
  NAND2_X1 U12354 ( .A1(n14203), .A2(n14204), .ZN(n14202) );
  NAND2_X1 U12355 ( .A1(n14196), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U12356 ( .A1(n14202), .A2(n9787), .ZN(n14212) );
  NAND2_X1 U12357 ( .A1(n14213), .A2(n14212), .ZN(n14211) );
  NAND2_X1 U12358 ( .A1(n14214), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12359 ( .A1(n14211), .A2(n9788), .ZN(n14226) );
  MUX2_X1 U12360 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10366), .S(n14228), .Z(
        n14227) );
  NAND2_X1 U12361 ( .A1(n14226), .A2(n14227), .ZN(n14225) );
  NAND2_X1 U12362 ( .A1(n14228), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U12363 ( .A1(n14225), .A2(n9789), .ZN(n9826) );
  MUX2_X1 U12364 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9526), .S(n9824), .Z(n9827)
         );
  NAND2_X1 U12365 ( .A1(n9826), .A2(n9827), .ZN(n9825) );
  NAND2_X1 U12366 ( .A1(n9824), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U12367 ( .A1(n9825), .A2(n9790), .ZN(n14241) );
  XNOR2_X1 U12368 ( .A(n14245), .B(n9791), .ZN(n14242) );
  NAND2_X1 U12369 ( .A1(n14241), .A2(n14242), .ZN(n14240) );
  NAND2_X1 U12370 ( .A1(n14245), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U12371 ( .A1(n14240), .A2(n9792), .ZN(n14251) );
  INV_X1 U12372 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U12373 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9793), .S(n14258), .Z(
        n14252) );
  NAND2_X1 U12374 ( .A1(n14251), .A2(n14252), .ZN(n14250) );
  NAND2_X1 U12375 ( .A1(n14258), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U12376 ( .A1(n14250), .A2(n9794), .ZN(n9797) );
  NOR2_X1 U12377 ( .A1(n11866), .A2(n14187), .ZN(n9795) );
  NAND2_X1 U12378 ( .A1(n9797), .A2(n9798), .ZN(n9812) );
  OAI211_X1 U12379 ( .C1(n9798), .C2(n9797), .A(n15070), .B(n9812), .ZN(n9799)
         );
  OAI211_X1 U12380 ( .C1(n9801), .C2(n15053), .A(n9800), .B(n9799), .ZN(
        P1_U3251) );
  OR2_X1 U12381 ( .A1(n10496), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U12382 ( .A1(n9806), .A2(n9804), .ZN(n9802) );
  INV_X1 U12383 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15208) );
  MUX2_X1 U12384 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15208), .S(n10801), .Z(
        n9803) );
  NAND2_X1 U12385 ( .A1(n9802), .A2(n9803), .ZN(n10087) );
  INV_X1 U12386 ( .A(n9803), .ZN(n9805) );
  NAND3_X1 U12387 ( .A1(n9806), .A2(n9805), .A3(n9804), .ZN(n9807) );
  AND2_X1 U12388 ( .A1(n10087), .A2(n9807), .ZN(n9817) );
  NOR2_X1 U12389 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10513), .ZN(n9809) );
  NOR2_X1 U12390 ( .A1(n14320), .A2(n10085), .ZN(n9808) );
  AOI211_X1 U12391 ( .C1(n14269), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9809), .B(
        n9808), .ZN(n9816) );
  INV_X1 U12392 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9810) );
  MUX2_X1 U12393 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9810), .S(n10801), .Z(n9814) );
  NAND2_X1 U12394 ( .A1(n10496), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U12395 ( .A1(n9812), .A2(n9811), .ZN(n9813) );
  NAND2_X1 U12396 ( .A1(n9813), .A2(n9814), .ZN(n10094) );
  OAI211_X1 U12397 ( .C1(n9814), .C2(n9813), .A(n15070), .B(n10094), .ZN(n9815) );
  OAI211_X1 U12398 ( .C1(n9817), .C2(n15053), .A(n9816), .B(n9815), .ZN(
        P1_U3252) );
  INV_X1 U12399 ( .A(n9818), .ZN(n9819) );
  AOI21_X1 U12400 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9830) );
  INV_X1 U12401 ( .A(n14320), .ZN(n15067) );
  INV_X1 U12402 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U12403 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10599) );
  OAI21_X1 U12404 ( .B1(n15075), .B2(n9822), .A(n10599), .ZN(n9823) );
  AOI21_X1 U12405 ( .B1(n9824), .B2(n15067), .A(n9823), .ZN(n9829) );
  OAI211_X1 U12406 ( .C1(n9827), .C2(n9826), .A(n15070), .B(n9825), .ZN(n9828)
         );
  OAI211_X1 U12407 ( .C1(n9830), .C2(n15053), .A(n9829), .B(n9828), .ZN(
        P1_U3248) );
  INV_X1 U12408 ( .A(n15228), .ZN(n9832) );
  XNOR2_X1 U12409 ( .A(n15228), .B(n9831), .ZN(n15231) );
  INV_X1 U12410 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10020) );
  NOR3_X1 U12411 ( .A1(n15231), .A2(n7308), .A3(n10020), .ZN(n15230) );
  AOI21_X1 U12412 ( .B1(n9832), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15230), .ZN(
        n9880) );
  MUX2_X1 U12413 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9833), .S(n9878), .Z(n9879)
         );
  NOR2_X1 U12414 ( .A1(n9880), .A2(n9879), .ZN(n9981) );
  NOR2_X1 U12415 ( .A1(n9878), .A2(n9833), .ZN(n9976) );
  MUX2_X1 U12416 ( .A(n9834), .B(P2_REG1_REG_3__SCAN_IN), .S(n9984), .Z(n9835)
         );
  OAI21_X1 U12417 ( .B1(n9981), .B2(n9976), .A(n9835), .ZN(n9979) );
  INV_X1 U12418 ( .A(n9984), .ZN(n9836) );
  NAND2_X1 U12419 ( .A1(n9836), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9950) );
  MUX2_X1 U12420 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9837), .S(n9955), .Z(n9949)
         );
  AOI21_X1 U12421 ( .B1(n9979), .B2(n9950), .A(n9949), .ZN(n9948) );
  NOR2_X1 U12422 ( .A1(n9955), .A2(n9837), .ZN(n9936) );
  MUX2_X1 U12423 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9838), .S(n9851), .Z(n9935)
         );
  OAI21_X1 U12424 ( .B1(n9948), .B2(n9936), .A(n9935), .ZN(n9938) );
  OAI21_X1 U12425 ( .B1(n9838), .B2(n9941), .A(n9938), .ZN(n15246) );
  MUX2_X1 U12426 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9839), .S(n9852), .Z(n15245) );
  NAND2_X1 U12427 ( .A1(n15246), .A2(n15245), .ZN(n15244) );
  NAND2_X1 U12428 ( .A1(n9852), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9886) );
  MUX2_X1 U12429 ( .A(n8527), .B(P2_REG1_REG_7__SCAN_IN), .S(n9895), .Z(n9885)
         );
  AOI21_X1 U12430 ( .B1(n15244), .B2(n9886), .A(n9885), .ZN(n9898) );
  AOI21_X1 U12431 ( .B1(n9895), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9898), .ZN(
        n9964) );
  MUX2_X1 U12432 ( .A(n8545), .B(P2_REG1_REG_8__SCAN_IN), .S(n9853), .Z(n9963)
         );
  NOR2_X1 U12433 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  AOI21_X1 U12434 ( .B1(n9853), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9962), .ZN(
        n9865) );
  INV_X1 U12435 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U12436 ( .A1(n10173), .A2(n9840), .ZN(n9841) );
  NAND2_X1 U12437 ( .A1(n8437), .A2(n9841), .ZN(n9843) );
  NAND2_X1 U12438 ( .A1(n9843), .A2(n9842), .ZN(n9861) );
  OR2_X1 U12439 ( .A1(n9855), .A2(P2_U3088), .ZN(n14010) );
  INV_X1 U12440 ( .A(n14010), .ZN(n9844) );
  NAND2_X1 U12441 ( .A1(n9861), .A2(n9844), .ZN(n9854) );
  NOR3_X1 U12442 ( .A1(n9865), .A2(n15452), .A3(n15265), .ZN(n9857) );
  NOR2_X1 U12443 ( .A1(n15228), .A2(n9846), .ZN(n9847) );
  AOI21_X1 U12444 ( .B1(n9846), .B2(n15228), .A(n9847), .ZN(n15236) );
  NAND3_X1 U12445 ( .A1(n15236), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n15234) );
  INV_X1 U12446 ( .A(n9847), .ZN(n9848) );
  NAND2_X1 U12447 ( .A1(n15234), .A2(n9848), .ZN(n9876) );
  XNOR2_X1 U12448 ( .A(n9878), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9875) );
  INV_X1 U12449 ( .A(n9878), .ZN(n9849) );
  MUX2_X1 U12450 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10711), .S(n9984), .Z(n9972) );
  NOR2_X1 U12451 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  NOR2_X1 U12452 ( .A1(n9984), .A2(n10711), .ZN(n9944) );
  MUX2_X1 U12453 ( .A(n10700), .B(P2_REG2_REG_4__SCAN_IN), .S(n9955), .Z(n9943) );
  OAI21_X1 U12454 ( .B1(n9971), .B2(n9944), .A(n9943), .ZN(n9942) );
  INV_X1 U12455 ( .A(n9955), .ZN(n9850) );
  NAND2_X1 U12456 ( .A1(n9850), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9931) );
  MUX2_X1 U12457 ( .A(n10655), .B(P2_REG2_REG_5__SCAN_IN), .S(n9851), .Z(n9930) );
  AOI21_X1 U12458 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n9851), .A(n9933), .ZN(
        n15249) );
  MUX2_X1 U12459 ( .A(n10685), .B(P2_REG2_REG_6__SCAN_IN), .S(n9852), .Z(
        n15248) );
  NOR2_X1 U12460 ( .A1(n15241), .A2(n10685), .ZN(n9890) );
  MUX2_X1 U12461 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10668), .S(n9895), .Z(n9889) );
  OAI21_X1 U12462 ( .B1(n15247), .B2(n9890), .A(n9889), .ZN(n9959) );
  NAND2_X1 U12463 ( .A1(n9895), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9958) );
  MUX2_X1 U12464 ( .A(n13882), .B(P2_REG2_REG_8__SCAN_IN), .S(n9853), .Z(n9957) );
  AOI21_X1 U12465 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9956) );
  NOR3_X1 U12466 ( .A1(n9860), .A2(n13861), .A3(n15263), .ZN(n9856) );
  AND2_X1 U12467 ( .A1(n9855), .A2(n9861), .ZN(n15227) );
  AND2_X1 U12468 ( .A1(n15227), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15300) );
  NOR3_X1 U12469 ( .A1(n9857), .A2(n9856), .A3(n15300), .ZN(n9871) );
  NAND2_X1 U12470 ( .A1(n9870), .A2(n13861), .ZN(n9859) );
  MUX2_X1 U12471 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13861), .S(n10012), .Z(
        n9858) );
  NAND2_X1 U12472 ( .A1(n9860), .A2(n9858), .ZN(n10011) );
  OAI21_X1 U12473 ( .B1(n9860), .B2(n9859), .A(n10011), .ZN(n9863) );
  INV_X1 U12474 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14845) );
  NAND2_X1 U12475 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11872) );
  OAI21_X1 U12476 ( .B1(n15297), .B2(n14845), .A(n11872), .ZN(n9862) );
  AOI21_X1 U12477 ( .B1(n9863), .B2(n15302), .A(n9862), .ZN(n9869) );
  NOR3_X1 U12478 ( .A1(n9865), .A2(n10012), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9867) );
  MUX2_X1 U12479 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15452), .S(n10012), .Z(
        n9864) );
  NAND2_X1 U12480 ( .A1(n9865), .A2(n9864), .ZN(n10007) );
  INV_X1 U12481 ( .A(n10007), .ZN(n9866) );
  INV_X1 U12482 ( .A(n15265), .ZN(n15305) );
  OAI21_X1 U12483 ( .B1(n9867), .B2(n9866), .A(n15305), .ZN(n9868) );
  OAI211_X1 U12484 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9868), .ZN(
        P2_U3223) );
  INV_X1 U12485 ( .A(n9872), .ZN(n9874) );
  OAI222_X1 U12486 ( .A1(n13282), .A2(n9874), .B1(n13284), .B2(n9873), .C1(
        n7055), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12487 ( .A(n15300), .ZN(n15290) );
  XNOR2_X1 U12488 ( .A(n9876), .B(n9875), .ZN(n9877) );
  OAI22_X1 U12489 ( .A1(n15290), .A2(n9878), .B1(n9877), .B2(n15263), .ZN(
        n9884) );
  AOI211_X1 U12490 ( .C1(n9880), .C2(n9879), .A(n9981), .B(n15265), .ZN(n9883)
         );
  INV_X1 U12491 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9881) );
  OAI22_X1 U12492 ( .A1(n15297), .A2(n9881), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10234), .ZN(n9882) );
  OR3_X1 U12493 ( .A1(n9884), .A2(n9883), .A3(n9882), .ZN(P2_U3216) );
  NAND3_X1 U12494 ( .A1(n15244), .A2(n9886), .A3(n9885), .ZN(n9887) );
  NAND2_X1 U12495 ( .A1(n9887), .A2(n15305), .ZN(n9897) );
  INV_X1 U12496 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9888) );
  NAND2_X1 U12497 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10580) );
  OAI21_X1 U12498 ( .B1(n15297), .B2(n9888), .A(n10580), .ZN(n9894) );
  INV_X1 U12499 ( .A(n9959), .ZN(n9892) );
  NOR3_X1 U12500 ( .A1(n15247), .A2(n9890), .A3(n9889), .ZN(n9891) );
  NOR3_X1 U12501 ( .A1(n9892), .A2(n9891), .A3(n15263), .ZN(n9893) );
  AOI211_X1 U12502 ( .C1(n15300), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9896)
         );
  OAI21_X1 U12503 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(P2_U3221) );
  CLKBUF_X1 U12504 ( .A(n9908), .Z(n9927) );
  INV_X1 U12505 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U12506 ( .A1(n9927), .A2(n9900), .ZN(P3_U3247) );
  INV_X1 U12507 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U12508 ( .A1(n9927), .A2(n9901), .ZN(P3_U3250) );
  INV_X1 U12509 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9902) );
  NOR2_X1 U12510 ( .A1(n9927), .A2(n9902), .ZN(P3_U3254) );
  INV_X1 U12511 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U12512 ( .A1(n9927), .A2(n9903), .ZN(P3_U3251) );
  INV_X1 U12513 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U12514 ( .A1(n9927), .A2(n9904), .ZN(P3_U3249) );
  INV_X1 U12515 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U12516 ( .A1(n9927), .A2(n9905), .ZN(P3_U3257) );
  INV_X1 U12517 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9906) );
  NOR2_X1 U12518 ( .A1(n9927), .A2(n9906), .ZN(P3_U3261) );
  INV_X1 U12519 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U12520 ( .A1(n9927), .A2(n9907), .ZN(P3_U3259) );
  INV_X1 U12521 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U12522 ( .A1(n9927), .A2(n9909), .ZN(P3_U3260) );
  INV_X1 U12523 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U12524 ( .A1(n9908), .A2(n9910), .ZN(P3_U3242) );
  INV_X1 U12525 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U12526 ( .A1(n9908), .A2(n9911), .ZN(P3_U3258) );
  INV_X1 U12527 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U12528 ( .A1(n9927), .A2(n9912), .ZN(P3_U3263) );
  INV_X1 U12529 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U12530 ( .A1(n9908), .A2(n9913), .ZN(P3_U3245) );
  INV_X1 U12531 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U12532 ( .A1(n9927), .A2(n9914), .ZN(P3_U3246) );
  INV_X1 U12533 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U12534 ( .A1(n9908), .A2(n9915), .ZN(P3_U3244) );
  INV_X1 U12535 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U12536 ( .A1(n9927), .A2(n9916), .ZN(P3_U3253) );
  INV_X1 U12537 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U12538 ( .A1(n9908), .A2(n9917), .ZN(P3_U3239) );
  INV_X1 U12539 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U12540 ( .A1(n9927), .A2(n9918), .ZN(P3_U3248) );
  INV_X1 U12541 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U12542 ( .A1(n9927), .A2(n9919), .ZN(P3_U3256) );
  INV_X1 U12543 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U12544 ( .A1(n9908), .A2(n9920), .ZN(P3_U3235) );
  INV_X1 U12545 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U12546 ( .A1(n9908), .A2(n9921), .ZN(P3_U3236) );
  INV_X1 U12547 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U12548 ( .A1(n9908), .A2(n9922), .ZN(P3_U3237) );
  INV_X1 U12549 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n13091) );
  NOR2_X1 U12550 ( .A1(n9908), .A2(n13091), .ZN(P3_U3238) );
  INV_X1 U12551 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n13173) );
  NOR2_X1 U12552 ( .A1(n9908), .A2(n13173), .ZN(P3_U3234) );
  INV_X1 U12553 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9923) );
  NOR2_X1 U12554 ( .A1(n9927), .A2(n9923), .ZN(P3_U3252) );
  INV_X1 U12555 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9924) );
  NOR2_X1 U12556 ( .A1(n9908), .A2(n9924), .ZN(P3_U3241) );
  INV_X1 U12557 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12558 ( .A1(n9927), .A2(n9925), .ZN(P3_U3262) );
  INV_X1 U12559 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U12560 ( .A1(n9927), .A2(n9926), .ZN(P3_U3255) );
  INV_X1 U12561 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U12562 ( .A1(n9927), .A2(n9928), .ZN(P3_U3240) );
  INV_X1 U12563 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U12564 ( .A1(n9927), .A2(n9929), .ZN(P3_U3243) );
  INV_X1 U12565 ( .A(n15297), .ZN(n15298) );
  AND2_X1 U12566 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n11853) );
  AND3_X1 U12567 ( .A1(n9942), .A2(n9931), .A3(n9930), .ZN(n9932) );
  NOR3_X1 U12568 ( .A1(n15263), .A2(n9933), .A3(n9932), .ZN(n9934) );
  AOI211_X1 U12569 ( .C1(n15298), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n11853), .B(
        n9934), .ZN(n9940) );
  OR3_X1 U12570 ( .A1(n9948), .A2(n9936), .A3(n9935), .ZN(n9937) );
  NAND3_X1 U12571 ( .A1(n15305), .A2(n9938), .A3(n9937), .ZN(n9939) );
  OAI211_X1 U12572 ( .C1(n15290), .C2(n9941), .A(n9940), .B(n9939), .ZN(
        P2_U3219) );
  AND2_X1 U12573 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10399) );
  INV_X1 U12574 ( .A(n9942), .ZN(n9946) );
  NOR3_X1 U12575 ( .A1(n9971), .A2(n9944), .A3(n9943), .ZN(n9945) );
  NOR3_X1 U12576 ( .A1(n15263), .A2(n9946), .A3(n9945), .ZN(n9947) );
  AOI211_X1 U12577 ( .C1(n15298), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10399), .B(
        n9947), .ZN(n9954) );
  INV_X1 U12578 ( .A(n9948), .ZN(n9952) );
  NAND3_X1 U12579 ( .A1(n9979), .A2(n9950), .A3(n9949), .ZN(n9951) );
  NAND3_X1 U12580 ( .A1(n15305), .A2(n9952), .A3(n9951), .ZN(n9953) );
  OAI211_X1 U12581 ( .C1(n15290), .C2(n9955), .A(n9954), .B(n9953), .ZN(
        P2_U3218) );
  INV_X1 U12582 ( .A(n9956), .ZN(n9961) );
  NAND3_X1 U12583 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n9960) );
  NAND3_X1 U12584 ( .A1(n9961), .A2(n15302), .A3(n9960), .ZN(n9969) );
  NAND2_X1 U12585 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11884) );
  AOI211_X1 U12586 ( .C1(n9964), .C2(n9963), .A(n9962), .B(n15265), .ZN(n9965)
         );
  INV_X1 U12587 ( .A(n9965), .ZN(n9966) );
  NAND2_X1 U12588 ( .A1(n11884), .A2(n9966), .ZN(n9967) );
  AOI21_X1 U12589 ( .B1(n15298), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9967), .ZN(
        n9968) );
  OAI211_X1 U12590 ( .C1(n15290), .C2(n9970), .A(n9969), .B(n9968), .ZN(
        P2_U3222) );
  AND2_X1 U12591 ( .A1(n15298), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n9975) );
  AOI211_X1 U12592 ( .C1(n9973), .C2(n9972), .A(n9971), .B(n15263), .ZN(n9974)
         );
  AOI211_X1 U12593 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n9975), 
        .B(n9974), .ZN(n9983) );
  INV_X1 U12594 ( .A(n9976), .ZN(n9978) );
  MUX2_X1 U12595 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9834), .S(n9984), .Z(n9977)
         );
  NAND2_X1 U12596 ( .A1(n9978), .A2(n9977), .ZN(n9980) );
  OAI211_X1 U12597 ( .C1(n9981), .C2(n9980), .A(n15305), .B(n9979), .ZN(n9982)
         );
  OAI211_X1 U12598 ( .C1(n15290), .C2(n9984), .A(n9983), .B(n9982), .ZN(
        P2_U3217) );
  INV_X1 U12599 ( .A(n11161), .ZN(n10003) );
  INV_X1 U12600 ( .A(n9985), .ZN(n9987) );
  INV_X1 U12601 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12602 ( .A1(n9987), .A2(n9986), .ZN(n10005) );
  NAND2_X1 U12603 ( .A1(n10005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9988) );
  XNOR2_X1 U12604 ( .A(n9988), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U12605 ( .A1(n11162), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14717), .ZN(n9989) );
  OAI21_X1 U12606 ( .B1(n10003), .B2(n12426), .A(n9989), .ZN(P1_U3343) );
  NAND2_X1 U12607 ( .A1(n12218), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9998) );
  INV_X1 U12608 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n13063) );
  OR2_X1 U12609 ( .A1(n11348), .A2(n13063), .ZN(n9997) );
  INV_X1 U12610 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10464) );
  INV_X1 U12611 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10500) );
  AND2_X1 U12612 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n9990) );
  NAND2_X1 U12613 ( .A1(n10822), .A2(n9990), .ZN(n10960) );
  NAND2_X1 U12614 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n9991) );
  NAND2_X1 U12615 ( .A1(n11437), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11538) );
  NAND2_X1 U12616 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n9992) );
  NAND2_X1 U12617 ( .A1(n12089), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12090) );
  INV_X1 U12618 ( .A(n12090), .ZN(n11913) );
  NAND2_X1 U12619 ( .A1(n11913), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11912) );
  INV_X1 U12620 ( .A(n11912), .ZN(n9993) );
  NAND2_X1 U12621 ( .A1(n9993), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12117) );
  OAI21_X1 U12622 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9993), .A(n12117), .ZN(
        n14494) );
  OR2_X1 U12623 ( .A1(n12202), .A2(n14494), .ZN(n9996) );
  INV_X1 U12624 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9994) );
  OR2_X1 U12625 ( .A1(n12219), .A2(n9994), .ZN(n9995) );
  NAND4_X1 U12626 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n14378) );
  NAND2_X1 U12627 ( .A1(n6576), .A2(n14378), .ZN(n9999) );
  OAI21_X1 U12628 ( .B1(n6576), .B2(n11429), .A(n9999), .ZN(P1_U3583) );
  INV_X1 U12629 ( .A(n10000), .ZN(n10002) );
  INV_X1 U12630 ( .A(n12652), .ZN(n14903) );
  OAI222_X1 U12631 ( .A1(n13282), .A2(n10002), .B1(n13284), .B2(n10001), .C1(
        n14903), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12632 ( .A(n15268), .ZN(n11022) );
  OAI222_X1 U12633 ( .A1(n14024), .A2(n10004), .B1(n14022), .B2(n10003), .C1(
        n11022), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12634 ( .A(n11166), .ZN(n10028) );
  NAND2_X1 U12635 ( .A1(n10006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10128) );
  XNOR2_X1 U12636 ( .A(n10128), .B(n10127), .ZN(n11169) );
  OAI222_X1 U12637 ( .A1(n12426), .A2(n10028), .B1(n11169), .B2(P1_U3086), 
        .C1(n11167), .C2(n12296), .ZN(P1_U3342) );
  OAI21_X1 U12638 ( .B1(n10012), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10007), .ZN(
        n10009) );
  MUX2_X1 U12639 ( .A(n8578), .B(P2_REG1_REG_10__SCAN_IN), .S(n11005), .Z(
        n10008) );
  NOR2_X1 U12640 ( .A1(n10009), .A2(n10008), .ZN(n13527) );
  AOI211_X1 U12641 ( .C1(n10009), .C2(n10008), .A(n15265), .B(n13527), .ZN(
        n10010) );
  INV_X1 U12642 ( .A(n10010), .ZN(n10019) );
  NAND2_X1 U12643 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11259)
         );
  MUX2_X1 U12644 ( .A(n13840), .B(P2_REG2_REG_10__SCAN_IN), .S(n11005), .Z(
        n10014) );
  OAI21_X1 U12645 ( .B1(n10012), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10011), .ZN(
        n10013) );
  AOI211_X1 U12646 ( .C1(n10014), .C2(n10013), .A(n11004), .B(n15263), .ZN(
        n10015) );
  INV_X1 U12647 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U12648 ( .A1(n11259), .A2(n10016), .ZN(n10017) );
  AOI21_X1 U12649 ( .B1(n15298), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10017), 
        .ZN(n10018) );
  OAI211_X1 U12650 ( .C1(n15290), .C2(n11018), .A(n10019), .B(n10018), .ZN(
        P2_U3224) );
  OAI22_X1 U12651 ( .A1(n10723), .A2(n15263), .B1(n15265), .B2(n10020), .ZN(
        n10023) );
  NAND2_X1 U12652 ( .A1(n15302), .A2(n10723), .ZN(n10021) );
  OAI211_X1 U12653 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15265), .A(n15290), .B(
        n10021), .ZN(n10022) );
  MUX2_X1 U12654 ( .A(n10023), .B(n10022), .S(P2_IR_REG_0__SCAN_IN), .Z(n10026) );
  INV_X1 U12655 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10024) );
  OAI22_X1 U12656 ( .A1(n15297), .A2(n10024), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10722), .ZN(n10025) );
  OR2_X1 U12657 ( .A1(n10026), .A2(n10025), .ZN(P2_U3214) );
  OAI222_X1 U12658 ( .A1(P2_U3088), .A2(n15273), .B1(n14022), .B2(n10028), 
        .C1(n10027), .C2(n14024), .ZN(P2_U3314) );
  INV_X1 U12659 ( .A(n10029), .ZN(n10031) );
  OAI22_X1 U12660 ( .A1(n14925), .A2(P3_U3151), .B1(SI_17_), .B2(n13284), .ZN(
        n10030) );
  AOI21_X1 U12661 ( .B1(n10031), .B2(n14835), .A(n10030), .ZN(P3_U3278) );
  AND2_X2 U12662 ( .A1(n10056), .A2(n10032), .ZN(n10035) );
  INV_X1 U12663 ( .A(n10056), .ZN(n10033) );
  INV_X1 U12664 ( .A(n14721), .ZN(n14182) );
  OAI222_X1 U12665 ( .A1(n12370), .A2(n15135), .B1(n12369), .B2(n6817), .C1(
        n10056), .C2(n14182), .ZN(n10075) );
  OAI22_X1 U12666 ( .A1(n12369), .A2(n11938), .B1(n6575), .B2(n12370), .ZN(
        n10036) );
  INV_X1 U12667 ( .A(n10036), .ZN(n10037) );
  AOI21_X1 U12668 ( .B1(n10040), .B2(n10039), .A(n10066), .ZN(n10063) );
  INV_X1 U12669 ( .A(n10041), .ZN(n10047) );
  NAND2_X1 U12670 ( .A1(n14445), .A2(n10042), .ZN(n11923) );
  INV_X1 U12671 ( .A(n12237), .ZN(n10045) );
  NAND2_X1 U12672 ( .A1(n15194), .A2(n10045), .ZN(n10046) );
  NOR2_X1 U12673 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  NAND2_X1 U12674 ( .A1(n10058), .A2(n10049), .ZN(n10051) );
  NAND2_X1 U12675 ( .A1(n10051), .A2(n10050), .ZN(n10057) );
  AND2_X1 U12676 ( .A1(n10057), .A2(n10052), .ZN(n11342) );
  AND2_X1 U12677 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  AND2_X1 U12678 ( .A1(n10056), .A2(n10055), .ZN(n12290) );
  NAND2_X1 U12679 ( .A1(n10057), .A2(n12290), .ZN(n10528) );
  NOR2_X1 U12680 ( .A1(n10528), .A2(P1_U3086), .ZN(n10073) );
  AND2_X1 U12681 ( .A1(n14152), .A2(n14569), .ZN(n14140) );
  INV_X1 U12682 ( .A(n14570), .ZN(n14593) );
  NOR2_X1 U12683 ( .A1(n6855), .A2(n14593), .ZN(n10450) );
  AOI22_X1 U12684 ( .A1(n14140), .A2(n14174), .B1(n10450), .B2(n14152), .ZN(
        n10059) );
  OAI21_X1 U12685 ( .B1(n10073), .B2(n14175), .A(n10059), .ZN(n10060) );
  AOI21_X1 U12686 ( .B1(n14995), .B2(n10061), .A(n10060), .ZN(n10062) );
  OAI21_X1 U12687 ( .B1(n10063), .B2(n14989), .A(n10062), .ZN(P1_U3222) );
  INV_X1 U12688 ( .A(n10064), .ZN(n10065) );
  OAI22_X1 U12689 ( .A1(n12369), .A2(n6855), .B1(n15148), .B2(n12370), .ZN(
        n10531) );
  AOI22_X1 U12690 ( .A1(n12329), .A2(n14172), .B1(n10035), .B2(n15093), .ZN(
        n10067) );
  XNOR2_X1 U12691 ( .A(n10067), .B(n12413), .ZN(n10533) );
  XOR2_X1 U12692 ( .A(n10531), .B(n10533), .Z(n10068) );
  AOI21_X1 U12693 ( .B1(n10069), .B2(n10068), .A(n10535), .ZN(n10072) );
  AOI22_X1 U12694 ( .A1(n6776), .A2(n14569), .B1(n14570), .B2(n14171), .ZN(
        n15081) );
  INV_X1 U12695 ( .A(n14152), .ZN(n14124) );
  OAI22_X1 U12696 ( .A1(n10073), .A2(n14194), .B1(n15081), .B2(n14124), .ZN(
        n10070) );
  AOI21_X1 U12697 ( .B1(n14995), .B2(n15093), .A(n10070), .ZN(n10071) );
  OAI21_X1 U12698 ( .B1(n10072), .B2(n14989), .A(n10071), .ZN(P1_U3237) );
  INV_X1 U12699 ( .A(n14995), .ZN(n14128) );
  INV_X1 U12700 ( .A(n10073), .ZN(n10078) );
  AOI21_X1 U12701 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n14188) );
  AND2_X1 U12702 ( .A1(n14152), .A2(n14570), .ZN(n14141) );
  INV_X1 U12703 ( .A(n14141), .ZN(n14983) );
  OAI22_X1 U12704 ( .A1(n14188), .A2(n14989), .B1(n11938), .B2(n14983), .ZN(
        n10077) );
  AOI21_X1 U12705 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10078), .A(n10077), .ZN(
        n10079) );
  OAI21_X1 U12706 ( .B1(n15135), .B2(n14128), .A(n10079), .ZN(P1_U3232) );
  INV_X1 U12707 ( .A(n10080), .ZN(n10082) );
  OAI222_X1 U12708 ( .A1(n13282), .A2(n10082), .B1(n13284), .B2(n10081), .C1(
        n12657), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U12709 ( .A1(n13461), .A2(P2_U3947), .ZN(n10083) );
  OAI21_X1 U12710 ( .B1(P2_U3947), .B2(n10084), .A(n10083), .ZN(P2_U3553) );
  INV_X1 U12711 ( .A(n11162), .ZN(n10107) );
  INV_X1 U12712 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14857) );
  MUX2_X1 U12713 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14857), .S(n11162), .Z(
        n10092) );
  INV_X1 U12714 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U12715 ( .A1(n10085), .A2(n15208), .ZN(n10086) );
  NAND2_X1 U12716 ( .A1(n10087), .A2(n10086), .ZN(n14265) );
  INV_X1 U12717 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15211) );
  MUX2_X1 U12718 ( .A(n15211), .B(P1_REG1_REG_10__SCAN_IN), .S(n14273), .Z(
        n14264) );
  OR2_X1 U12719 ( .A1(n14265), .A2(n14264), .ZN(n14266) );
  NAND2_X1 U12720 ( .A1(n14273), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U12721 ( .A1(n14266), .A2(n10088), .ZN(n15034) );
  MUX2_X1 U12722 ( .A(n15010), .B(P1_REG1_REG_11__SCAN_IN), .S(n15037), .Z(
        n15033) );
  NOR2_X1 U12723 ( .A1(n15034), .A2(n15033), .ZN(n15036) );
  AOI21_X1 U12724 ( .B1(n15010), .B2(n10089), .A(n15036), .ZN(n10090) );
  INV_X1 U12725 ( .A(n10090), .ZN(n10091) );
  NAND2_X1 U12726 ( .A1(n10092), .A2(n10091), .ZN(n10259) );
  OAI21_X1 U12727 ( .B1(n10092), .B2(n10091), .A(n10259), .ZN(n10103) );
  NAND2_X1 U12728 ( .A1(n10801), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U12729 ( .A1(n10094), .A2(n10093), .ZN(n14271) );
  INV_X1 U12730 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n13179) );
  MUX2_X1 U12731 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n13179), .S(n14273), .Z(
        n14272) );
  NAND2_X1 U12732 ( .A1(n14271), .A2(n14272), .ZN(n14270) );
  NAND2_X1 U12733 ( .A1(n14273), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12734 ( .A1(n14270), .A2(n10095), .ZN(n15032) );
  OR2_X1 U12735 ( .A1(n15037), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U12736 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n15037), .ZN(n10096) );
  AND2_X1 U12737 ( .A1(n10097), .A2(n10096), .ZN(n15031) );
  AND2_X1 U12738 ( .A1(n15032), .A2(n15031), .ZN(n15041) );
  AOI21_X1 U12739 ( .B1(n15037), .B2(P1_REG2_REG_11__SCAN_IN), .A(n15041), 
        .ZN(n10101) );
  INV_X1 U12740 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U12741 ( .A(n10098), .B(P1_REG2_REG_12__SCAN_IN), .S(n11162), .Z(
        n10099) );
  INV_X1 U12742 ( .A(n10099), .ZN(n10100) );
  NAND2_X1 U12743 ( .A1(n10100), .A2(n10101), .ZN(n10262) );
  OAI21_X1 U12744 ( .B1(n10101), .B2(n10100), .A(n10262), .ZN(n10102) );
  AOI22_X1 U12745 ( .A1(n15071), .A2(n10103), .B1(n15070), .B2(n10102), .ZN(
        n10106) );
  NAND2_X1 U12746 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11611)
         );
  INV_X1 U12747 ( .A(n11611), .ZN(n10104) );
  AOI21_X1 U12748 ( .B1(n14269), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10104), 
        .ZN(n10105) );
  OAI211_X1 U12749 ( .C1(n10107), .C2(n14320), .A(n10106), .B(n10105), .ZN(
        P1_U3255) );
  NOR2_X1 U12750 ( .A1(n10109), .A2(n10108), .ZN(n10124) );
  INV_X1 U12751 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10121) );
  XNOR2_X1 U12752 ( .A(n11959), .B(n11960), .ZN(n12258) );
  XNOR2_X1 U12753 ( .A(n10111), .B(n12258), .ZN(n10370) );
  XNOR2_X1 U12754 ( .A(n10112), .B(n12258), .ZN(n10115) );
  NAND2_X1 U12755 ( .A1(n14171), .A2(n14569), .ZN(n10114) );
  NAND2_X1 U12756 ( .A1(n14169), .A2(n14570), .ZN(n10113) );
  NAND2_X1 U12757 ( .A1(n10114), .A2(n10113), .ZN(n10539) );
  AOI21_X1 U12758 ( .B1(n10115), .B2(n6917), .A(n10539), .ZN(n10367) );
  OAI21_X1 U12759 ( .B1(n10286), .B2(n11959), .A(n14538), .ZN(n10116) );
  OR2_X1 U12760 ( .A1(n10117), .A2(n10116), .ZN(n10364) );
  INV_X1 U12761 ( .A(n10364), .ZN(n10118) );
  AOI21_X1 U12762 ( .B1(n11961), .B2(n15169), .A(n10118), .ZN(n10119) );
  OAI211_X1 U12763 ( .C1(n10370), .C2(n15131), .A(n10367), .B(n10119), .ZN(
        n10125) );
  NAND2_X1 U12764 ( .A1(n10125), .A2(n15200), .ZN(n10120) );
  OAI21_X1 U12765 ( .B1(n15200), .B2(n10121), .A(n10120), .ZN(P1_U3471) );
  NAND2_X1 U12766 ( .A1(n10125), .A2(n15213), .ZN(n10126) );
  OAI21_X1 U12767 ( .B1(n15213), .B2(n9768), .A(n10126), .ZN(P1_U3532) );
  INV_X1 U12768 ( .A(n11358), .ZN(n10131) );
  NAND2_X1 U12769 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  NAND2_X1 U12770 ( .A1(n10129), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10130) );
  XNOR2_X1 U12771 ( .A(n10130), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15057) );
  INV_X1 U12772 ( .A(n15057), .ZN(n10852) );
  OAI222_X1 U12773 ( .A1(n12426), .A2(n10131), .B1(n10852), .B2(P1_U3086), 
        .C1(n12990), .C2(n12296), .ZN(P1_U3341) );
  INV_X1 U12774 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10132) );
  INV_X1 U12775 ( .A(n11006), .ZN(n15289) );
  OAI222_X1 U12776 ( .A1(n14024), .A2(n10132), .B1(n14022), .B2(n10131), .C1(
        n15289), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12777 ( .A(n15541), .ZN(n14929) );
  OAI21_X1 U12778 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10144) );
  INV_X1 U12779 ( .A(n15458), .ZN(n15529) );
  INV_X1 U12780 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10137) );
  OAI22_X1 U12781 ( .A1(n15529), .A2(n10137), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10136), .ZN(n10143) );
  OR2_X1 U12782 ( .A1(n10139), .A2(n10138), .ZN(n10140) );
  AOI21_X1 U12783 ( .B1(n10141), .B2(n10140), .A(n15547), .ZN(n10142) );
  AOI211_X1 U12784 ( .C1(n14929), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10149) );
  XNOR2_X1 U12785 ( .A(n10146), .B(n10145), .ZN(n10147) );
  NAND2_X1 U12786 ( .A1(n10147), .A2(n15538), .ZN(n10148) );
  OAI211_X1 U12787 ( .C1(n15531), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        P3_U3184) );
  AND2_X1 U12788 ( .A1(n10152), .A2(n10151), .ZN(n15472) );
  AND2_X1 U12789 ( .A1(n9321), .A2(n11685), .ZN(n11656) );
  INV_X1 U12790 ( .A(n11656), .ZN(n10155) );
  OAI22_X1 U12791 ( .A1(n15467), .A2(n8123), .B1(n12576), .B2(n10349), .ZN(
        n10154) );
  AOI21_X1 U12792 ( .B1(n15469), .B2(n10155), .A(n10154), .ZN(n10156) );
  OAI21_X1 U12793 ( .B1(n15472), .B2(n10319), .A(n10156), .ZN(P3_U3172) );
  OAI222_X1 U12794 ( .A1(P3_U3151), .A2(n12673), .B1(n13284), .B2(n10158), 
        .C1(n13282), .C2(n10157), .ZN(P3_U3276) );
  NAND2_X1 U12795 ( .A1(n13466), .A2(P2_U3947), .ZN(n10159) );
  OAI21_X1 U12796 ( .B1(P2_U3947), .B2(n10160), .A(n10159), .ZN(P2_U3554) );
  INV_X1 U12797 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10167) );
  XNOR2_X1 U12798 ( .A(n10161), .B(n10162), .ZN(n10717) );
  AOI211_X1 U12799 ( .C1(n15224), .C2(n15322), .A(n13979), .B(n10701), .ZN(
        n10714) );
  AOI21_X1 U12800 ( .B1(n15434), .B2(n15224), .A(n10714), .ZN(n10165) );
  XNOR2_X1 U12801 ( .A(n10163), .B(n10162), .ZN(n10164) );
  INV_X1 U12802 ( .A(n13854), .ZN(n13874) );
  OAI22_X1 U12803 ( .A1(n6854), .A2(n13874), .B1(n6814), .B2(n13872), .ZN(
        n15214) );
  AOI21_X1 U12804 ( .B1(n10164), .B2(n15313), .A(n15214), .ZN(n10710) );
  OAI211_X1 U12805 ( .C1(n15407), .C2(n10717), .A(n10165), .B(n10710), .ZN(
        n10483) );
  NAND2_X1 U12806 ( .A1(n10483), .A2(n15444), .ZN(n10166) );
  OAI21_X1 U12807 ( .B1(n15444), .B2(n10167), .A(n10166), .ZN(P2_U3439) );
  XNOR2_X1 U12808 ( .A(n8968), .B(n13384), .ZN(n10226) );
  OR2_X2 U12809 ( .A1(n8957), .A2(n13979), .ZN(n13331) );
  NAND2_X1 U12810 ( .A1(n13515), .A2(n13331), .ZN(n10228) );
  XNOR2_X1 U12811 ( .A(n10226), .B(n10228), .ZN(n10225) );
  OR2_X1 U12812 ( .A1(n10721), .A2(n13331), .ZN(n10168) );
  NAND2_X1 U12813 ( .A1(n10249), .A2(n10168), .ZN(n10273) );
  AND2_X1 U12814 ( .A1(n13384), .A2(n10721), .ZN(n10169) );
  OR2_X1 U12815 ( .A1(n10273), .A2(n10169), .ZN(n10224) );
  XOR2_X1 U12816 ( .A(n10225), .B(n10224), .Z(n10189) );
  INV_X1 U12817 ( .A(n15363), .ZN(n10170) );
  NAND2_X1 U12818 ( .A1(n10171), .A2(n10170), .ZN(n10175) );
  NOR2_X1 U12819 ( .A1(n15366), .A2(n10175), .ZN(n10172) );
  NAND2_X1 U12820 ( .A1(n10172), .A2(n15367), .ZN(n10182) );
  INV_X1 U12821 ( .A(n10182), .ZN(n10184) );
  INV_X1 U12822 ( .A(n10173), .ZN(n10174) );
  AND2_X1 U12823 ( .A1(n10183), .A2(n15366), .ZN(n10180) );
  NAND2_X1 U12824 ( .A1(n10183), .A2(n10175), .ZN(n10179) );
  OR2_X1 U12825 ( .A1(n10180), .A2(n10255), .ZN(n10254) );
  NOR2_X1 U12826 ( .A1(n10254), .A2(P2_U3088), .ZN(n10275) );
  INV_X1 U12827 ( .A(n10275), .ZN(n10187) );
  AOI22_X1 U12828 ( .A1(n13854), .A2(n8959), .B1(n13514), .B2(n13851), .ZN(
        n10251) );
  OR2_X1 U12829 ( .A1(n10182), .A2(n10181), .ZN(n15216) );
  AND2_X1 U12830 ( .A1(n10719), .A2(n10718), .ZN(n10657) );
  NAND2_X1 U12831 ( .A1(n10184), .A2(n10657), .ZN(n10185) );
  OAI22_X1 U12832 ( .A1(n10251), .A2(n15216), .B1(n13447), .B2(n10864), .ZN(
        n10186) );
  AOI21_X1 U12833 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10187), .A(n10186), .ZN(
        n10188) );
  OAI21_X1 U12834 ( .B1(n10189), .B2(n13480), .A(n10188), .ZN(P2_U3194) );
  NOR2_X1 U12835 ( .A1(n10207), .A2(n10190), .ZN(n10191) );
  NAND2_X1 U12836 ( .A1(n10193), .A2(n10212), .ZN(n10320) );
  AOI21_X1 U12837 ( .B1(n10194), .B2(n10981), .A(n10321), .ZN(n10220) );
  INV_X1 U12838 ( .A(n10195), .ZN(n10202) );
  INV_X1 U12839 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10196) );
  MUX2_X1 U12840 ( .A(n10981), .B(n10196), .S(n13279), .Z(n10198) );
  NAND2_X1 U12841 ( .A1(n10198), .A2(n10197), .ZN(n10340) );
  INV_X1 U12842 ( .A(n10198), .ZN(n10199) );
  NAND2_X1 U12843 ( .A1(n10199), .A2(n10212), .ZN(n10200) );
  AND2_X1 U12844 ( .A1(n10340), .A2(n10200), .ZN(n10201) );
  OAI21_X1 U12845 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(n10341) );
  INV_X1 U12846 ( .A(n10341), .ZN(n10205) );
  NOR3_X1 U12847 ( .A1(n10203), .A2(n10202), .A3(n10201), .ZN(n10204) );
  OAI21_X1 U12848 ( .B1(n10205), .B2(n10204), .A(n15538), .ZN(n10219) );
  NOR2_X1 U12849 ( .A1(n10207), .A2(n10206), .ZN(n10208) );
  NAND2_X1 U12850 ( .A1(n10210), .A2(n10212), .ZN(n10325) );
  OAI21_X1 U12851 ( .B1(n10210), .B2(n10212), .A(n10325), .ZN(n10211) );
  AOI21_X1 U12852 ( .B1(n10211), .B2(n10196), .A(n10326), .ZN(n10216) );
  AND2_X1 U12853 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12854 ( .A1(n15531), .A2(n10212), .ZN(n10213) );
  AOI211_X1 U12855 ( .C1(n15458), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n10214), .B(
        n10213), .ZN(n10215) );
  OAI21_X1 U12856 ( .B1(n10216), .B2(n15541), .A(n10215), .ZN(n10217) );
  INV_X1 U12857 ( .A(n10217), .ZN(n10218) );
  OAI211_X1 U12858 ( .C1(n10220), .C2(n15547), .A(n10219), .B(n10218), .ZN(
        P3_U3189) );
  NOR3_X1 U12859 ( .A1(n11656), .A2(n14950), .A3(n10221), .ZN(n10222) );
  AOI21_X1 U12860 ( .B1(n8165), .B2(n6800), .A(n10222), .ZN(n10346) );
  MUX2_X1 U12861 ( .A(n7761), .B(n10346), .S(n15613), .Z(n10223) );
  OAI21_X1 U12862 ( .B1(n10349), .B2(n13263), .A(n10223), .ZN(P3_U3390) );
  NAND2_X1 U12863 ( .A1(n10225), .A2(n10224), .ZN(n10230) );
  INV_X1 U12864 ( .A(n10226), .ZN(n10227) );
  NAND2_X1 U12865 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  NAND2_X1 U12866 ( .A1(n10230), .A2(n10229), .ZN(n10388) );
  NAND2_X1 U12867 ( .A1(n13514), .A2(n13318), .ZN(n10391) );
  XNOR2_X1 U12868 ( .A(n15318), .B(n13384), .ZN(n10389) );
  XNOR2_X1 U12869 ( .A(n10391), .B(n10389), .ZN(n10387) );
  XNOR2_X1 U12870 ( .A(n10388), .B(n10387), .ZN(n10231) );
  NAND2_X1 U12871 ( .A1(n10231), .A2(n13492), .ZN(n10233) );
  OAI22_X1 U12872 ( .A1(n10270), .A2(n13874), .B1(n10402), .B2(n13872), .ZN(
        n15312) );
  AOI22_X1 U12873 ( .A1(n15312), .A2(n13476), .B1(n15318), .B2(n15223), .ZN(
        n10232) );
  OAI211_X1 U12874 ( .C1(n10275), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        P2_U3209) );
  XOR2_X1 U12875 ( .A(n10235), .B(n10355), .Z(n10247) );
  OAI21_X1 U12876 ( .B1(n10237), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10236), .ZN(
        n10243) );
  OAI22_X1 U12877 ( .A1(n15529), .A2(n7395), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10300), .ZN(n10242) );
  NAND2_X1 U12878 ( .A1(n10238), .A2(n10744), .ZN(n10239) );
  AOI21_X1 U12879 ( .B1(n10240), .B2(n10239), .A(n15547), .ZN(n10241) );
  AOI211_X1 U12880 ( .C1(n14929), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10246) );
  NAND2_X1 U12881 ( .A1(n14926), .A2(n6590), .ZN(n10245) );
  OAI211_X1 U12882 ( .C1(n10247), .C2(n14920), .A(n10246), .B(n10245), .ZN(
        P3_U3183) );
  XNOR2_X1 U12883 ( .A(n6573), .B(n10248), .ZN(n10866) );
  OAI211_X1 U12884 ( .C1(n10864), .C2(n10721), .A(n15323), .B(n15321), .ZN(
        n10860) );
  OAI21_X1 U12885 ( .B1(n10864), .B2(n15428), .A(n10860), .ZN(n10253) );
  XNOR2_X1 U12886 ( .A(n6573), .B(n10249), .ZN(n10252) );
  OAI21_X1 U12887 ( .B1(n10252), .B2(n13712), .A(n10251), .ZN(n10859) );
  AOI211_X1 U12888 ( .C1(n10866), .C2(n15379), .A(n10253), .B(n10859), .ZN(
        n15374) );
  NAND2_X1 U12889 ( .A1(n15455), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U12890 ( .B1(n15374), .B2(n15455), .A(n10256), .ZN(P2_U3500) );
  INV_X1 U12891 ( .A(n11432), .ZN(n10276) );
  NAND2_X1 U12892 ( .A1(n10257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10258) );
  XNOR2_X1 U12893 ( .A(n10258), .B(P1_IR_REG_15__SCAN_IN), .ZN(n15068) );
  INV_X1 U12894 ( .A(n15068), .ZN(n10842) );
  OAI222_X1 U12895 ( .A1(n12426), .A2(n10276), .B1(n10842), .B2(P1_U3086), 
        .C1(n6832), .C2(n12296), .ZN(P1_U3340) );
  MUX2_X1 U12896 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11173), .S(n11169), .Z(
        n10850) );
  OAI21_X1 U12897 ( .B1(n11162), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10259), 
        .ZN(n10849) );
  XOR2_X1 U12898 ( .A(n10850), .B(n10849), .Z(n10266) );
  INV_X1 U12899 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10260) );
  MUX2_X1 U12900 ( .A(n10260), .B(P1_REG2_REG_13__SCAN_IN), .S(n11169), .Z(
        n10261) );
  INV_X1 U12901 ( .A(n10261), .ZN(n10264) );
  OAI21_X1 U12902 ( .B1(n11162), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10262), 
        .ZN(n10263) );
  NOR2_X1 U12903 ( .A1(n10263), .A2(n10264), .ZN(n10838) );
  AOI211_X1 U12904 ( .C1(n10264), .C2(n10263), .A(n10838), .B(n15046), .ZN(
        n10265) );
  AOI21_X1 U12905 ( .B1(n15071), .B2(n10266), .A(n10265), .ZN(n10269) );
  NAND2_X1 U12906 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14110)
         );
  INV_X1 U12907 ( .A(n14110), .ZN(n10267) );
  AOI21_X1 U12908 ( .B1(n14269), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10267), 
        .ZN(n10268) );
  OAI211_X1 U12909 ( .C1(n11169), .C2(n14320), .A(n10269), .B(n10268), .ZN(
        P1_U3256) );
  NAND2_X1 U12910 ( .A1(n13476), .A2(n13851), .ZN(n13421) );
  INV_X1 U12911 ( .A(n13331), .ZN(n13732) );
  OR2_X1 U12912 ( .A1(n13480), .A2(n13732), .ZN(n13483) );
  OAI22_X1 U12913 ( .A1(n10270), .A2(n13421), .B1(n9237), .B2(n13483), .ZN(
        n10272) );
  NOR2_X1 U12914 ( .A1(n13447), .A2(n10721), .ZN(n10271) );
  AOI211_X1 U12915 ( .C1(n13492), .C2(n10273), .A(n10272), .B(n10271), .ZN(
        n10274) );
  OAI21_X1 U12916 ( .B1(n10275), .B2(n10722), .A(n10274), .ZN(P2_U3204) );
  INV_X1 U12917 ( .A(n15299), .ZN(n11026) );
  OAI222_X1 U12918 ( .A1(n14024), .A2(n10277), .B1(n14022), .B2(n10276), .C1(
        n11026), .C2(P2_U3088), .ZN(P2_U3312) );
  XNOR2_X1 U12919 ( .A(n10278), .B(n10279), .ZN(n15158) );
  XNOR2_X1 U12920 ( .A(n10280), .B(n10279), .ZN(n10284) );
  OR2_X1 U12921 ( .A1(n11960), .A2(n14593), .ZN(n10282) );
  NAND2_X1 U12922 ( .A1(n14172), .A2(n14569), .ZN(n10281) );
  NAND2_X1 U12923 ( .A1(n10282), .A2(n10281), .ZN(n14045) );
  INV_X1 U12924 ( .A(n14045), .ZN(n10283) );
  OAI21_X1 U12925 ( .B1(n10284), .B2(n15178), .A(n10283), .ZN(n10285) );
  AOI21_X1 U12926 ( .B1(n15158), .B2(n15084), .A(n10285), .ZN(n15160) );
  OAI21_X1 U12927 ( .B1(n15090), .B2(n15155), .A(n14538), .ZN(n10287) );
  OR2_X1 U12928 ( .A1(n10287), .A2(n10286), .ZN(n15154) );
  OAI22_X1 U12929 ( .A1(n14543), .A2(n15154), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14556), .ZN(n10289) );
  NOR2_X1 U12930 ( .A1(n15088), .A2(n15155), .ZN(n10288) );
  AOI211_X1 U12931 ( .C1(n15098), .C2(P1_REG2_REG_3__SCAN_IN), .A(n10289), .B(
        n10288), .ZN(n10291) );
  NAND2_X1 U12932 ( .A1(n15095), .A2(n15158), .ZN(n10290) );
  OAI211_X1 U12933 ( .C1(n15098), .C2(n15160), .A(n10291), .B(n10290), .ZN(
        P1_U3290) );
  OAI22_X1 U12934 ( .A1(n15467), .A2(n10737), .B1(n12576), .B2(n10734), .ZN(
        n10298) );
  MUX2_X1 U12935 ( .A(n15556), .B(n10735), .S(n10292), .Z(n10296) );
  NAND2_X1 U12936 ( .A1(n10293), .A2(n9321), .ZN(n10736) );
  NAND2_X1 U12937 ( .A1(n11659), .A2(n10294), .ZN(n10738) );
  MUX2_X1 U12938 ( .A(n10736), .B(n10738), .S(n12440), .Z(n10295) );
  AOI21_X1 U12939 ( .B1(n10296), .B2(n10295), .A(n12552), .ZN(n10297) );
  AOI211_X1 U12940 ( .C1(n15465), .C2(n10153), .A(n10298), .B(n10297), .ZN(
        n10299) );
  OAI21_X1 U12941 ( .B1(n15472), .B2(n10300), .A(n10299), .ZN(P3_U3162) );
  INV_X1 U12942 ( .A(n11526), .ZN(n10361) );
  INV_X1 U12943 ( .A(n10301), .ZN(n10302) );
  NAND2_X1 U12944 ( .A1(n10302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10303) );
  MUX2_X1 U12945 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10303), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10305) );
  NAND2_X1 U12946 ( .A1(n10305), .A2(n10304), .ZN(n14289) );
  OAI222_X1 U12947 ( .A1(n12426), .A2(n10361), .B1(n14289), .B2(P1_U3086), 
        .C1(n10306), .C2(n12296), .ZN(P1_U3339) );
  INV_X1 U12948 ( .A(n11833), .ZN(n15552) );
  INV_X1 U12949 ( .A(n10308), .ZN(n10309) );
  XNOR2_X1 U12950 ( .A(n13265), .B(n10309), .ZN(n10311) );
  AND2_X1 U12951 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  NAND2_X1 U12952 ( .A1(n10313), .A2(n10312), .ZN(n10316) );
  MUX2_X1 U12953 ( .A(n10314), .B(n10346), .S(n15566), .Z(n10318) );
  NAND2_X1 U12954 ( .A1(n14950), .A2(n11833), .ZN(n10315) );
  NAND2_X1 U12955 ( .A1(n14944), .A2(n7767), .ZN(n10317) );
  OAI211_X1 U12956 ( .C1(n15553), .C2(n10319), .A(n10318), .B(n10317), .ZN(
        P3_U3233) );
  INV_X1 U12957 ( .A(n10320), .ZN(n10322) );
  INV_X1 U12958 ( .A(n14832), .ZN(n10335) );
  AOI22_X1 U12959 ( .A1(n10335), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11046), 
        .B2(n14832), .ZN(n10323) );
  NOR2_X1 U12960 ( .A1(n10324), .A2(n10323), .ZN(n10435) );
  AOI21_X1 U12961 ( .B1(n10324), .B2(n10323), .A(n10435), .ZN(n10345) );
  INV_X1 U12962 ( .A(n10325), .ZN(n10327) );
  INV_X1 U12963 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U12964 ( .A1(n10335), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n15626), 
        .B2(n14832), .ZN(n10328) );
  AOI21_X1 U12965 ( .B1(n10329), .B2(n10328), .A(n10420), .ZN(n10333) );
  NOR2_X1 U12966 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10926), .ZN(n10330) );
  AOI21_X1 U12967 ( .B1(n15458), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10330), .ZN(
        n10332) );
  NAND2_X1 U12968 ( .A1(n14926), .A2(n10335), .ZN(n10331) );
  OAI211_X1 U12969 ( .C1(n10333), .C2(n15541), .A(n10332), .B(n10331), .ZN(
        n10334) );
  INV_X1 U12970 ( .A(n10334), .ZN(n10344) );
  MUX2_X1 U12971 ( .A(n11046), .B(n15626), .S(n13279), .Z(n10336) );
  NAND2_X1 U12972 ( .A1(n10336), .A2(n10335), .ZN(n10428) );
  INV_X1 U12973 ( .A(n10336), .ZN(n10337) );
  NAND2_X1 U12974 ( .A1(n10337), .A2(n14832), .ZN(n10338) );
  NAND2_X1 U12975 ( .A1(n10428), .A2(n10338), .ZN(n10339) );
  AND3_X1 U12976 ( .A1(n10341), .A2(n10340), .A3(n10339), .ZN(n10342) );
  OAI21_X1 U12977 ( .B1(n10433), .B2(n10342), .A(n15538), .ZN(n10343) );
  OAI211_X1 U12978 ( .C1(n10345), .C2(n15547), .A(n10344), .B(n10343), .ZN(
        P3_U3190) );
  MUX2_X1 U12979 ( .A(n10347), .B(n10346), .S(n15631), .Z(n10348) );
  OAI21_X1 U12980 ( .B1(n10349), .B2(n13211), .A(n10348), .ZN(P3_U3459) );
  NAND3_X1 U12981 ( .A1(n15547), .A2(n15541), .A3(n14920), .ZN(n10354) );
  NAND2_X1 U12982 ( .A1(n14929), .A2(n9630), .ZN(n10351) );
  AOI22_X1 U12983 ( .A1(n15458), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10350) );
  OAI211_X1 U12984 ( .C1(n10352), .C2(n15547), .A(n10351), .B(n10350), .ZN(
        n10353) );
  AOI21_X1 U12985 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10359) );
  NAND2_X1 U12986 ( .A1(n15538), .A2(n10356), .ZN(n10357) );
  NAND2_X1 U12987 ( .A1(n10359), .A2(n10358), .ZN(P3_U3182) );
  INV_X1 U12988 ( .A(n11110), .ZN(n11033) );
  OAI222_X1 U12989 ( .A1(P2_U3088), .A2(n11033), .B1(n14022), .B2(n10361), 
        .C1(n10360), .C2(n14024), .ZN(P2_U3311) );
  INV_X1 U12990 ( .A(n10362), .ZN(n10363) );
  OAI22_X1 U12991 ( .A1(n14543), .A2(n10364), .B1(n10544), .B2(n14556), .ZN(
        n10365) );
  AOI21_X1 U12992 ( .B1(n14558), .B2(n11961), .A(n10365), .ZN(n10369) );
  MUX2_X1 U12993 ( .A(n10367), .B(n10366), .S(n15098), .Z(n10368) );
  OAI211_X1 U12994 ( .C1(n14601), .C2(n10370), .A(n10369), .B(n10368), .ZN(
        P1_U3289) );
  NAND2_X1 U12995 ( .A1(n14174), .A2(n15135), .ZN(n11930) );
  NAND2_X1 U12996 ( .A1(n15094), .A2(n14538), .ZN(n14389) );
  INV_X1 U12997 ( .A(n14389), .ZN(n10372) );
  OAI21_X1 U12998 ( .B1(n10372), .B2(n14558), .A(n10371), .ZN(n10376) );
  INV_X1 U12999 ( .A(n14556), .ZN(n15085) );
  NAND2_X1 U13000 ( .A1(n6776), .A2(n14570), .ZN(n15132) );
  OAI21_X1 U13001 ( .B1(n15130), .B2(n15178), .A(n15132), .ZN(n10373) );
  AOI21_X1 U13002 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n15085), .A(n10373), .ZN(
        n10374) );
  MUX2_X1 U13003 ( .A(n10374), .B(n9467), .S(n15098), .Z(n10375) );
  OAI211_X1 U13004 ( .C1(n15130), .C2(n14601), .A(n10376), .B(n10375), .ZN(
        P1_U3293) );
  INV_X1 U13005 ( .A(n12022), .ZN(n10386) );
  NAND2_X1 U13006 ( .A1(n10304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10377) );
  XNOR2_X1 U13007 ( .A(n10377), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14296) );
  INV_X1 U13008 ( .A(n14296), .ZN(n14304) );
  OAI222_X1 U13009 ( .A1(n12426), .A2(n10386), .B1(n14304), .B2(P1_U3086), 
        .C1(n6851), .C2(n12296), .ZN(P1_U3338) );
  INV_X1 U13010 ( .A(n15184), .ZN(n15157) );
  OAI21_X1 U13011 ( .B1(n10593), .B2(n15194), .A(n10378), .ZN(n10380) );
  AOI211_X1 U13012 ( .C1(n15157), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        n10383) );
  OR2_X1 U13013 ( .A1(n10383), .A2(n15210), .ZN(n10382) );
  OAI21_X1 U13014 ( .B1(n15213), .B2(n9772), .A(n10382), .ZN(P1_U3533) );
  INV_X1 U13015 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10385) );
  OR2_X1 U13016 ( .A1(n10383), .A2(n15199), .ZN(n10384) );
  OAI21_X1 U13017 ( .B1(n15200), .B2(n10385), .A(n10384), .ZN(P1_U3474) );
  OAI222_X1 U13018 ( .A1(n14024), .A2(n13072), .B1(n14022), .B2(n10386), .C1(
        n13543), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13019 ( .A1(n10388), .A2(n10387), .ZN(n10393) );
  INV_X1 U13020 ( .A(n10389), .ZN(n10390) );
  NAND2_X1 U13021 ( .A1(n10391), .A2(n10390), .ZN(n10392) );
  AND2_X1 U13022 ( .A1(n13513), .A2(n13318), .ZN(n10394) );
  XNOR2_X1 U13023 ( .A(n15224), .B(n13384), .ZN(n10395) );
  NAND2_X1 U13024 ( .A1(n10394), .A2(n10395), .ZN(n10398) );
  INV_X1 U13025 ( .A(n10394), .ZN(n10396) );
  INV_X1 U13026 ( .A(n10395), .ZN(n10403) );
  NAND2_X1 U13027 ( .A1(n10396), .A2(n10403), .ZN(n10397) );
  NAND2_X1 U13028 ( .A1(n10398), .A2(n10397), .ZN(n15219) );
  NAND2_X1 U13029 ( .A1(n13512), .A2(n13318), .ZN(n10557) );
  XNOR2_X1 U13030 ( .A(n15383), .B(n13384), .ZN(n11858) );
  XNOR2_X1 U13031 ( .A(n10557), .B(n11858), .ZN(n10405) );
  INV_X1 U13032 ( .A(n13421), .ZN(n13451) );
  AOI21_X1 U13033 ( .B1(n13451), .B2(n13511), .A(n10399), .ZN(n10401) );
  NAND2_X1 U13034 ( .A1(n13476), .A2(n13854), .ZN(n13409) );
  INV_X1 U13035 ( .A(n13409), .ZN(n13452) );
  NAND2_X1 U13036 ( .A1(n13452), .A2(n13513), .ZN(n10400) );
  OAI211_X1 U13037 ( .C1(n15226), .C2(n10705), .A(n10401), .B(n10400), .ZN(
        n10408) );
  INV_X1 U13038 ( .A(n6621), .ZN(n15218) );
  NOR3_X1 U13039 ( .A1(n10403), .A2(n10402), .A3(n13483), .ZN(n10404) );
  AOI21_X1 U13040 ( .B1(n15218), .B2(n13492), .A(n10404), .ZN(n10406) );
  NOR2_X1 U13041 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  AOI211_X1 U13042 ( .C1(n15383), .C2(n15223), .A(n10408), .B(n10407), .ZN(
        n10409) );
  OAI21_X1 U13043 ( .B1(n11857), .B2(n13480), .A(n10409), .ZN(P2_U3202) );
  OAI21_X1 U13044 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(n10418) );
  AOI22_X1 U13045 ( .A1(n15463), .A2(n10413), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10416) );
  INV_X1 U13046 ( .A(n15467), .ZN(n10414) );
  AOI22_X1 U13047 ( .A1(n10414), .A2(n12599), .B1(n15465), .B2(n15461), .ZN(
        n10415) );
  OAI211_X1 U13048 ( .C1(n12549), .C2(n11148), .A(n10416), .B(n10415), .ZN(
        n10417) );
  AOI21_X1 U13049 ( .B1(n10418), .B2(n15469), .A(n10417), .ZN(n10419) );
  INV_X1 U13050 ( .A(n10419), .ZN(P3_U3170) );
  NAND2_X1 U13051 ( .A1(n10421), .A2(n10441), .ZN(n10765) );
  OAI21_X1 U13052 ( .B1(n10421), .B2(n10441), .A(n10765), .ZN(n10422) );
  INV_X1 U13053 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15629) );
  AOI21_X1 U13054 ( .B1(n10422), .B2(n15629), .A(n10766), .ZN(n10446) );
  MUX2_X1 U13055 ( .A(n10423), .B(n15629), .S(n13279), .Z(n10425) );
  NAND2_X1 U13056 ( .A1(n10425), .A2(n10424), .ZN(n10778) );
  INV_X1 U13057 ( .A(n10425), .ZN(n10426) );
  NAND2_X1 U13058 ( .A1(n10426), .A2(n10441), .ZN(n10427) );
  NAND2_X1 U13059 ( .A1(n10778), .A2(n10427), .ZN(n10429) );
  NAND2_X1 U13060 ( .A1(n10429), .A2(n10428), .ZN(n10432) );
  INV_X1 U13061 ( .A(n10428), .ZN(n10431) );
  INV_X1 U13062 ( .A(n10429), .ZN(n10430) );
  OAI21_X1 U13063 ( .B1(n10433), .B2(n10431), .A(n10430), .ZN(n10779) );
  OAI21_X1 U13064 ( .B1(n10433), .B2(n10432), .A(n10779), .ZN(n10440) );
  AND2_X1 U13065 ( .A1(n14832), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10434) );
  OAI21_X1 U13066 ( .B1(n10436), .B2(n10441), .A(n10758), .ZN(n10437) );
  NOR2_X1 U13067 ( .A1(n10423), .A2(n10437), .ZN(n10759) );
  AOI21_X1 U13068 ( .B1(n10437), .B2(n10423), .A(n10759), .ZN(n10438) );
  NOR2_X1 U13069 ( .A1(n10438), .A2(n15547), .ZN(n10439) );
  AOI21_X1 U13070 ( .B1(n15538), .B2(n10440), .A(n10439), .ZN(n10445) );
  NOR2_X1 U13071 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11082), .ZN(n10443) );
  NOR2_X1 U13072 ( .A1(n15531), .A2(n10441), .ZN(n10442) );
  AOI211_X1 U13073 ( .C1(n15458), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n10443), .B(
        n10442), .ZN(n10444) );
  OAI211_X1 U13074 ( .C1(n10446), .C2(n15541), .A(n10445), .B(n10444), .ZN(
        P3_U3191) );
  NAND2_X1 U13075 ( .A1(n12255), .A2(n14591), .ZN(n10449) );
  OAI21_X1 U13076 ( .B1(n6575), .B2(n15135), .A(n15092), .ZN(n10453) );
  XNOR2_X1 U13077 ( .A(n6776), .B(n10453), .ZN(n10448) );
  MUX2_X1 U13078 ( .A(n10449), .B(n10448), .S(n6817), .Z(n10452) );
  OAI21_X1 U13079 ( .B1(n6817), .B2(n14591), .A(n15178), .ZN(n10451) );
  AOI21_X1 U13080 ( .B1(n10452), .B2(n10451), .A(n10450), .ZN(n15142) );
  OR2_X1 U13081 ( .A1(n10453), .A2(n15091), .ZN(n15141) );
  OAI22_X1 U13082 ( .A1(n14543), .A2(n15141), .B1(n14175), .B2(n14556), .ZN(
        n10456) );
  XOR2_X1 U13083 ( .A(n10454), .B(n12255), .Z(n15140) );
  OAI22_X1 U13084 ( .A1(n6575), .A2(n15088), .B1(n14601), .B2(n15140), .ZN(
        n10455) );
  AOI211_X1 U13085 ( .C1(P1_REG2_REG_1__SCAN_IN), .C2(n15086), .A(n10456), .B(
        n10455), .ZN(n10457) );
  OAI21_X1 U13086 ( .B1(n15098), .B2(n15142), .A(n10457), .ZN(P1_U3292) );
  NAND2_X1 U13087 ( .A1(n10460), .A2(n12234), .ZN(n10462) );
  AOI22_X1 U13088 ( .A1(n12223), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12066), 
        .B2(n14245), .ZN(n10461) );
  NAND2_X1 U13089 ( .A1(n10462), .A2(n10461), .ZN(n11972) );
  XNOR2_X1 U13090 ( .A(n11972), .B(n14168), .ZN(n12259) );
  XNOR2_X1 U13091 ( .A(n10486), .B(n10474), .ZN(n10471) );
  NAND2_X1 U13092 ( .A1(n12147), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10470) );
  INV_X1 U13093 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10463) );
  OR2_X1 U13094 ( .A1(n12149), .A2(n10463), .ZN(n10469) );
  NAND2_X1 U13095 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NAND2_X1 U13096 ( .A1(n10501), .A2(n10466), .ZN(n10897) );
  OR2_X1 U13097 ( .A1(n12202), .A2(n10897), .ZN(n10468) );
  OR2_X1 U13098 ( .A1(n12219), .A2(n9793), .ZN(n10467) );
  NAND4_X1 U13099 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n14167) );
  AOI22_X1 U13100 ( .A1(n14569), .A2(n14169), .B1(n14167), .B2(n14570), .ZN(
        n10753) );
  OAI21_X1 U13101 ( .B1(n10471), .B2(n15178), .A(n10753), .ZN(n15163) );
  INV_X1 U13102 ( .A(n15163), .ZN(n10482) );
  OR2_X1 U13103 ( .A1(n11964), .A2(n14169), .ZN(n10472) );
  NAND2_X1 U13104 ( .A1(n10475), .A2(n10474), .ZN(n10509) );
  OAI21_X1 U13105 ( .B1(n10475), .B2(n10474), .A(n10509), .ZN(n15165) );
  OAI211_X1 U13106 ( .C1(n7091), .C2(n7090), .A(n14538), .B(n10623), .ZN(
        n15162) );
  NAND2_X1 U13107 ( .A1(n14558), .A2(n11972), .ZN(n10479) );
  INV_X1 U13108 ( .A(n10477), .ZN(n10755) );
  AOI22_X1 U13109 ( .A1(n15086), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10755), 
        .B2(n15085), .ZN(n10478) );
  OAI211_X1 U13110 ( .C1(n15162), .C2(n14543), .A(n10479), .B(n10478), .ZN(
        n10480) );
  AOI21_X1 U13111 ( .B1(n15165), .B2(n14562), .A(n10480), .ZN(n10481) );
  OAI21_X1 U13112 ( .B1(n10482), .B2(n15098), .A(n10481), .ZN(P1_U3287) );
  NAND2_X1 U13113 ( .A1(n10483), .A2(n15457), .ZN(n10484) );
  OAI21_X1 U13114 ( .B1(n15457), .B2(n9834), .A(n10484), .ZN(P2_U3502) );
  OR2_X1 U13115 ( .A1(n15098), .A2(n15178), .ZN(n14564) );
  INV_X1 U13116 ( .A(n14168), .ZN(n10487) );
  OR2_X1 U13117 ( .A1(n11972), .A2(n10487), .ZN(n10485) );
  NAND2_X1 U13118 ( .A1(n10486), .A2(n10485), .ZN(n10489) );
  NAND2_X1 U13119 ( .A1(n11972), .A2(n10487), .ZN(n10488) );
  NAND2_X1 U13120 ( .A1(n10490), .A2(n12234), .ZN(n10492) );
  AOI22_X1 U13121 ( .A1(n12223), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12066), 
        .B2(n14258), .ZN(n10491) );
  INV_X1 U13122 ( .A(n14167), .ZN(n10890) );
  AND2_X1 U13123 ( .A1(n15170), .A2(n10890), .ZN(n10493) );
  OR2_X1 U13124 ( .A1(n15170), .A2(n10890), .ZN(n10494) );
  NAND2_X1 U13125 ( .A1(n10495), .A2(n12234), .ZN(n10498) );
  AOI22_X1 U13126 ( .A1(n12223), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12066), 
        .B2(n10496), .ZN(n10497) );
  NAND2_X1 U13127 ( .A1(n10498), .A2(n10497), .ZN(n11983) );
  NAND2_X1 U13128 ( .A1(n12218), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10507) );
  OR2_X1 U13129 ( .A1(n11348), .A2(n10499), .ZN(n10506) );
  NAND2_X1 U13130 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  NAND2_X1 U13131 ( .A1(n10514), .A2(n10502), .ZN(n11142) );
  OR2_X1 U13132 ( .A1(n12202), .A2(n11142), .ZN(n10505) );
  OR2_X1 U13133 ( .A1(n12219), .A2(n10503), .ZN(n10504) );
  NAND4_X1 U13134 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n14166) );
  INV_X1 U13135 ( .A(n14166), .ZN(n10907) );
  XNOR2_X1 U13136 ( .A(n11983), .B(n10907), .ZN(n12263) );
  INV_X1 U13137 ( .A(n12263), .ZN(n10798) );
  XNOR2_X1 U13138 ( .A(n10799), .B(n10798), .ZN(n15179) );
  OR2_X1 U13139 ( .A1(n11972), .A2(n14168), .ZN(n10508) );
  NAND2_X1 U13140 ( .A1(n10509), .A2(n10508), .ZN(n10616) );
  XNOR2_X1 U13141 ( .A(n15170), .B(n14167), .ZN(n12261) );
  OR2_X1 U13142 ( .A1(n15170), .A2(n14167), .ZN(n10510) );
  NAND2_X1 U13143 ( .A1(n10511), .A2(n12263), .ZN(n10817) );
  OAI21_X1 U13144 ( .B1(n10511), .B2(n12263), .A(n10817), .ZN(n15182) );
  INV_X1 U13145 ( .A(n11983), .ZN(n15177) );
  AND2_X2 U13146 ( .A1(n10626), .A2(n15177), .ZN(n10912) );
  INV_X1 U13147 ( .A(n10912), .ZN(n10512) );
  OAI211_X1 U13148 ( .C1(n15177), .C2(n10626), .A(n10512), .B(n14538), .ZN(
        n15176) );
  NAND2_X1 U13149 ( .A1(n14167), .A2(n14569), .ZN(n10522) );
  NAND2_X1 U13150 ( .A1(n12218), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10520) );
  OR2_X1 U13151 ( .A1(n11348), .A2(n15208), .ZN(n10519) );
  INV_X1 U13152 ( .A(n10822), .ZN(n10516) );
  NAND2_X1 U13153 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  NAND2_X1 U13154 ( .A1(n10516), .A2(n10515), .ZN(n11340) );
  OR2_X1 U13155 ( .A1(n12202), .A2(n11340), .ZN(n10518) );
  OR2_X1 U13156 ( .A1(n12219), .A2(n9810), .ZN(n10517) );
  NAND4_X1 U13157 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n14165) );
  NAND2_X1 U13158 ( .A1(n14165), .A2(n14570), .ZN(n10521) );
  NAND2_X1 U13159 ( .A1(n10522), .A2(n10521), .ZN(n11140) );
  INV_X1 U13160 ( .A(n11140), .ZN(n15175) );
  OAI22_X1 U13161 ( .A1(n15086), .A2(n15175), .B1(n11142), .B2(n14556), .ZN(
        n10524) );
  NOR2_X1 U13162 ( .A1(n15088), .A2(n15177), .ZN(n10523) );
  AOI211_X1 U13163 ( .C1(n15086), .C2(P1_REG2_REG_8__SCAN_IN), .A(n10524), .B(
        n10523), .ZN(n10525) );
  OAI21_X1 U13164 ( .B1(n14543), .B2(n15176), .A(n10525), .ZN(n10526) );
  AOI21_X1 U13165 ( .B1(n15182), .B2(n14562), .A(n10526), .ZN(n10527) );
  OAI21_X1 U13166 ( .B1(n14564), .B2(n15179), .A(n10527), .ZN(P1_U3285) );
  INV_X2 U13167 ( .A(n12371), .ZN(n12411) );
  AOI22_X1 U13168 ( .A1(n12329), .A2(n14170), .B1(n12411), .B2(n11961), .ZN(
        n10529) );
  XOR2_X1 U13169 ( .A(n12327), .B(n10529), .Z(n10588) );
  AOI22_X1 U13170 ( .A1(n12412), .A2(n14171), .B1(n12363), .B2(n14046), .ZN(
        n10537) );
  AOI22_X1 U13171 ( .A1(n12411), .A2(n14046), .B1(n12329), .B2(n14171), .ZN(
        n10530) );
  XNOR2_X1 U13172 ( .A(n10530), .B(n12413), .ZN(n10536) );
  INV_X1 U13173 ( .A(n10531), .ZN(n10532) );
  XOR2_X1 U13174 ( .A(n10537), .B(n10536), .Z(n14043) );
  OAI22_X1 U13175 ( .A1(n12369), .A2(n11960), .B1(n11959), .B2(n12370), .ZN(
        n10585) );
  XOR2_X1 U13176 ( .A(n10589), .B(n10588), .Z(n10538) );
  NAND2_X1 U13177 ( .A1(n10538), .A2(n14119), .ZN(n10543) );
  NAND2_X1 U13178 ( .A1(n14152), .A2(n10539), .ZN(n10540) );
  NAND2_X1 U13179 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14222) );
  NAND2_X1 U13180 ( .A1(n10540), .A2(n14222), .ZN(n10541) );
  AOI21_X1 U13181 ( .B1(n14995), .B2(n11961), .A(n10541), .ZN(n10542) );
  OAI211_X1 U13182 ( .C1(n14998), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        P1_U3230) );
  XOR2_X1 U13183 ( .A(n10546), .B(n10545), .Z(n10551) );
  INV_X1 U13184 ( .A(n11120), .ZN(n10549) );
  NAND2_X1 U13185 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15523) );
  OAI21_X1 U13186 ( .B1(n12576), .B2(n15585), .A(n15523), .ZN(n10548) );
  OAI22_X1 U13187 ( .A1(n7247), .A2(n11083), .B1(n15467), .B2(n11125), .ZN(
        n10547) );
  AOI211_X1 U13188 ( .C1(n10549), .C2(n12573), .A(n10548), .B(n10547), .ZN(
        n10550) );
  OAI21_X1 U13189 ( .B1(n10551), .B2(n12552), .A(n10550), .ZN(P3_U3167) );
  INV_X1 U13190 ( .A(n10552), .ZN(n10553) );
  OAI222_X1 U13191 ( .A1(P3_U3151), .A2(n10555), .B1(n13284), .B2(n10554), 
        .C1(n13282), .C2(n10553), .ZN(P3_U3275) );
  INV_X1 U13192 ( .A(n11858), .ZN(n10556) );
  NAND2_X1 U13193 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  NAND2_X1 U13194 ( .A1(n11857), .A2(n10558), .ZN(n10559) );
  XNOR2_X1 U13195 ( .A(n15390), .B(n13384), .ZN(n10560) );
  NAND2_X1 U13196 ( .A1(n13511), .A2(n13318), .ZN(n10561) );
  XNOR2_X1 U13197 ( .A(n10560), .B(n10561), .ZN(n11859) );
  INV_X1 U13198 ( .A(n10560), .ZN(n10562) );
  NAND2_X1 U13199 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  XNOR2_X1 U13200 ( .A(n15396), .B(n13384), .ZN(n10564) );
  AND2_X1 U13201 ( .A1(n13510), .A2(n13318), .ZN(n10565) );
  NAND2_X1 U13202 ( .A1(n10564), .A2(n10565), .ZN(n10575) );
  INV_X1 U13203 ( .A(n10564), .ZN(n10574) );
  INV_X1 U13204 ( .A(n10565), .ZN(n10566) );
  NAND2_X1 U13205 ( .A1(n10574), .A2(n10566), .ZN(n10567) );
  NAND2_X1 U13206 ( .A1(n10575), .A2(n10567), .ZN(n10640) );
  XNOR2_X1 U13207 ( .A(n15404), .B(n13384), .ZN(n10568) );
  AND2_X1 U13208 ( .A1(n13509), .A2(n13318), .ZN(n10569) );
  NAND2_X1 U13209 ( .A1(n10568), .A2(n10569), .ZN(n11213) );
  INV_X1 U13210 ( .A(n10568), .ZN(n11889) );
  INV_X1 U13211 ( .A(n10569), .ZN(n10570) );
  NAND2_X1 U13212 ( .A1(n11889), .A2(n10570), .ZN(n10571) );
  AND2_X1 U13213 ( .A1(n11213), .A2(n10571), .ZN(n10576) );
  INV_X1 U13214 ( .A(n10576), .ZN(n10572) );
  AOI21_X1 U13215 ( .B1(n10637), .B2(n10572), .A(n13480), .ZN(n10579) );
  NOR3_X1 U13216 ( .A1(n10574), .A2(n10573), .A3(n13483), .ZN(n10578) );
  NAND2_X1 U13217 ( .A1(n10637), .A2(n10575), .ZN(n10577) );
  OAI21_X1 U13218 ( .B1(n10579), .B2(n10578), .A(n11888), .ZN(n10584) );
  OAI21_X1 U13219 ( .B1(n11873), .B2(n13421), .A(n10580), .ZN(n10582) );
  NOR2_X1 U13220 ( .A1(n15226), .A2(n10670), .ZN(n10581) );
  AOI211_X1 U13221 ( .C1(n13452), .C2(n13510), .A(n10582), .B(n10581), .ZN(
        n10583) );
  OAI211_X1 U13222 ( .C1(n10671), .C2(n13447), .A(n10584), .B(n10583), .ZN(
        P2_U3185) );
  NAND2_X1 U13223 ( .A1(n12411), .A2(n11964), .ZN(n10591) );
  NAND2_X1 U13224 ( .A1(n12363), .A2(n14169), .ZN(n10590) );
  NAND2_X1 U13225 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  XNOR2_X1 U13226 ( .A(n10592), .B(n12413), .ZN(n10596) );
  OAI22_X1 U13227 ( .A1(n12369), .A2(n10594), .B1(n10593), .B2(n12370), .ZN(
        n10595) );
  NOR2_X1 U13228 ( .A1(n10596), .A2(n10595), .ZN(n10746) );
  INV_X1 U13229 ( .A(n10746), .ZN(n10597) );
  NAND2_X1 U13230 ( .A1(n10596), .A2(n10595), .ZN(n10745) );
  NAND2_X1 U13231 ( .A1(n10597), .A2(n10745), .ZN(n10598) );
  XNOR2_X1 U13232 ( .A(n10747), .B(n10598), .ZN(n10605) );
  OAI21_X1 U13233 ( .B1(n14124), .B2(n10600), .A(n10599), .ZN(n10603) );
  NOR2_X1 U13234 ( .A1(n14998), .A2(n10601), .ZN(n10602) );
  AOI211_X1 U13235 ( .C1(n14995), .C2(n11964), .A(n10603), .B(n10602), .ZN(
        n10604) );
  OAI21_X1 U13236 ( .B1(n10605), .B2(n14989), .A(n10604), .ZN(P1_U3227) );
  OAI211_X1 U13237 ( .C1(n10608), .C2(n10607), .A(n10606), .B(n15469), .ZN(
        n10613) );
  OAI22_X1 U13238 ( .A1(n6737), .A2(n11083), .B1(n15467), .B2(n10928), .ZN(
        n10611) );
  OAI22_X1 U13239 ( .A1(n12576), .A2(n15589), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10609), .ZN(n10610) );
  NOR2_X1 U13240 ( .A1(n10611), .A2(n10610), .ZN(n10612) );
  OAI211_X1 U13241 ( .C1(n10881), .C2(n12549), .A(n10613), .B(n10612), .ZN(
        P3_U3179) );
  XNOR2_X1 U13242 ( .A(n10614), .B(n10615), .ZN(n10621) );
  OR2_X1 U13243 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  NAND2_X1 U13244 ( .A1(n10618), .A2(n10617), .ZN(n15167) );
  NAND2_X1 U13245 ( .A1(n15167), .A2(n15084), .ZN(n10620) );
  AOI22_X1 U13246 ( .A1(n14569), .A2(n14168), .B1(n14166), .B2(n14570), .ZN(
        n10619) );
  OAI211_X1 U13247 ( .C1(n15178), .C2(n10621), .A(n10620), .B(n10619), .ZN(
        n15174) );
  MUX2_X1 U13248 ( .A(n15174), .B(P1_REG2_REG_7__SCAN_IN), .S(n15098), .Z(
        n10622) );
  INV_X1 U13249 ( .A(n10622), .ZN(n10633) );
  INV_X1 U13250 ( .A(n15170), .ZN(n10630) );
  NAND2_X1 U13251 ( .A1(n10623), .A2(n15170), .ZN(n10624) );
  NAND2_X1 U13252 ( .A1(n10624), .A2(n14538), .ZN(n10625) );
  NOR2_X1 U13253 ( .A1(n10626), .A2(n10625), .ZN(n15168) );
  NAND2_X1 U13254 ( .A1(n15168), .A2(n15094), .ZN(n10629) );
  INV_X1 U13255 ( .A(n10897), .ZN(n10627) );
  NAND2_X1 U13256 ( .A1(n15085), .A2(n10627), .ZN(n10628) );
  OAI211_X1 U13257 ( .C1(n10630), .C2(n15088), .A(n10629), .B(n10628), .ZN(
        n10631) );
  AOI21_X1 U13258 ( .B1(n15167), .B2(n15095), .A(n10631), .ZN(n10632) );
  NAND2_X1 U13259 ( .A1(n10633), .A2(n10632), .ZN(P1_U3286) );
  NAND2_X1 U13260 ( .A1(n13509), .A2(n13851), .ZN(n10635) );
  NAND2_X1 U13261 ( .A1(n13511), .A2(n13854), .ZN(n10634) );
  NAND2_X1 U13262 ( .A1(n10635), .A2(n10634), .ZN(n10681) );
  AOI22_X1 U13263 ( .A1(n10681), .A2(n13476), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10636) );
  OAI21_X1 U13264 ( .B1(n15226), .B2(n10690), .A(n10636), .ZN(n10642) );
  INV_X1 U13265 ( .A(n10637), .ZN(n10638) );
  AOI211_X1 U13266 ( .C1(n10640), .C2(n10639), .A(n13480), .B(n10638), .ZN(
        n10641) );
  AOI211_X1 U13267 ( .C1(n15396), .C2(n15223), .A(n10642), .B(n10641), .ZN(
        n10643) );
  INV_X1 U13268 ( .A(n10643), .ZN(P2_U3211) );
  INV_X1 U13269 ( .A(n15366), .ZN(n10644) );
  NAND2_X1 U13270 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  NAND2_X1 U13271 ( .A1(n6587), .A2(n10647), .ZN(n10677) );
  NAND2_X1 U13272 ( .A1(n6801), .A2(n10677), .ZN(n10648) );
  XNOR2_X1 U13273 ( .A(n10649), .B(n10650), .ZN(n15393) );
  XNOR2_X1 U13274 ( .A(n10651), .B(n10650), .ZN(n10654) );
  NAND2_X1 U13275 ( .A1(n13510), .A2(n13851), .ZN(n10653) );
  NAND2_X1 U13276 ( .A1(n13512), .A2(n13854), .ZN(n10652) );
  NAND2_X1 U13277 ( .A1(n10653), .A2(n10652), .ZN(n11854) );
  AOI21_X1 U13278 ( .B1(n10654), .B2(n15313), .A(n11854), .ZN(n15391) );
  MUX2_X1 U13279 ( .A(n10655), .B(n15391), .S(n13883), .Z(n10661) );
  INV_X1 U13280 ( .A(n10686), .ZN(n10656) );
  AOI211_X1 U13281 ( .C1(n15390), .C2(n10702), .A(n13979), .B(n10656), .ZN(
        n15389) );
  INV_X2 U13282 ( .A(n13883), .ZN(n15316) );
  OAI22_X1 U13283 ( .A1(n14957), .A2(n10658), .B1(n13880), .B2(n11856), .ZN(
        n10659) );
  AOI21_X1 U13284 ( .B1(n15389), .B2(n15326), .A(n10659), .ZN(n10660) );
  OAI211_X1 U13285 ( .C1(n14959), .C2(n15393), .A(n10661), .B(n10660), .ZN(
        P2_U3260) );
  XNOR2_X1 U13286 ( .A(n10662), .B(n10663), .ZN(n15408) );
  XNOR2_X1 U13287 ( .A(n10664), .B(n10663), .ZN(n10665) );
  NAND2_X1 U13288 ( .A1(n10665), .A2(n15313), .ZN(n10667) );
  AOI22_X1 U13289 ( .A1(n13854), .A2(n13510), .B1(n13853), .B2(n13851), .ZN(
        n10666) );
  AND2_X1 U13290 ( .A1(n10667), .A2(n10666), .ZN(n15411) );
  MUX2_X1 U13291 ( .A(n10668), .B(n15411), .S(n13883), .Z(n10674) );
  OAI21_X1 U13292 ( .B1(n10689), .B2(n10671), .A(n15323), .ZN(n10669) );
  NOR2_X1 U13293 ( .A1(n10669), .A2(n13885), .ZN(n15406) );
  OAI22_X1 U13294 ( .A1(n14957), .A2(n10671), .B1(n13880), .B2(n10670), .ZN(
        n10672) );
  AOI21_X1 U13295 ( .B1(n15406), .B2(n15326), .A(n10672), .ZN(n10673) );
  OAI211_X1 U13296 ( .C1(n14959), .C2(n15408), .A(n10674), .B(n10673), .ZN(
        P2_U3258) );
  XNOR2_X1 U13297 ( .A(n10676), .B(n10675), .ZN(n15400) );
  INV_X1 U13298 ( .A(n15400), .ZN(n10695) );
  INV_X1 U13299 ( .A(n10677), .ZN(n10678) );
  NAND2_X1 U13300 ( .A1(n13883), .A2(n10678), .ZN(n13892) );
  INV_X1 U13301 ( .A(n6801), .ZN(n10727) );
  NAND2_X1 U13302 ( .A1(n15400), .A2(n10727), .ZN(n10684) );
  XNOR2_X1 U13303 ( .A(n10680), .B(n10679), .ZN(n10682) );
  AOI21_X1 U13304 ( .B1(n10682), .B2(n15313), .A(n10681), .ZN(n10683) );
  AND2_X1 U13305 ( .A1(n10684), .A2(n10683), .ZN(n15402) );
  MUX2_X1 U13306 ( .A(n10685), .B(n15402), .S(n13883), .Z(n10694) );
  NAND2_X1 U13307 ( .A1(n10686), .A2(n15396), .ZN(n10687) );
  NAND2_X1 U13308 ( .A1(n10687), .A2(n15323), .ZN(n10688) );
  NOR2_X1 U13309 ( .A1(n10689), .A2(n10688), .ZN(n15398) );
  OAI22_X1 U13310 ( .A1(n14957), .A2(n10691), .B1(n13880), .B2(n10690), .ZN(
        n10692) );
  AOI21_X1 U13311 ( .B1(n15398), .B2(n15326), .A(n10692), .ZN(n10693) );
  OAI211_X1 U13312 ( .C1(n10695), .C2(n13892), .A(n10694), .B(n10693), .ZN(
        P2_U3259) );
  XNOR2_X1 U13313 ( .A(n10696), .B(n10697), .ZN(n15386) );
  XNOR2_X1 U13314 ( .A(n10698), .B(n10697), .ZN(n10699) );
  AOI222_X1 U13315 ( .A1(n15313), .A2(n10699), .B1(n13511), .B2(n13851), .C1(
        n13513), .C2(n13854), .ZN(n15385) );
  MUX2_X1 U13316 ( .A(n10700), .B(n15385), .S(n13883), .Z(n10709) );
  INV_X1 U13317 ( .A(n10701), .ZN(n10704) );
  INV_X1 U13318 ( .A(n10702), .ZN(n10703) );
  AOI211_X1 U13319 ( .C1(n15383), .C2(n10704), .A(n13979), .B(n10703), .ZN(
        n15382) );
  OAI22_X1 U13320 ( .A1(n14957), .A2(n10706), .B1(n10705), .B2(n13880), .ZN(
        n10707) );
  AOI21_X1 U13321 ( .B1(n15382), .B2(n15326), .A(n10707), .ZN(n10708) );
  OAI211_X1 U13322 ( .C1(n14959), .C2(n15386), .A(n10709), .B(n10708), .ZN(
        P2_U3261) );
  MUX2_X1 U13323 ( .A(n10711), .B(n10710), .S(n13883), .Z(n10716) );
  INV_X1 U13324 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15215) );
  OAI22_X1 U13325 ( .A1(n14957), .A2(n10712), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13880), .ZN(n10713) );
  AOI21_X1 U13326 ( .B1(n10714), .B2(n15326), .A(n10713), .ZN(n10715) );
  OAI211_X1 U13327 ( .C1(n14959), .C2(n10717), .A(n10716), .B(n10715), .ZN(
        P2_U3262) );
  AOI21_X1 U13328 ( .B1(n10718), .B2(n13883), .A(n15326), .ZN(n10733) );
  INV_X1 U13329 ( .A(n10719), .ZN(n10720) );
  OR2_X1 U13330 ( .A1(n10721), .A2(n10720), .ZN(n15368) );
  INV_X1 U13331 ( .A(n13892), .ZN(n10726) );
  INV_X1 U13332 ( .A(n15369), .ZN(n10725) );
  OAI22_X1 U13333 ( .A1(n13883), .A2(n10723), .B1(n10722), .B2(n13880), .ZN(
        n10724) );
  AOI21_X1 U13334 ( .B1(n10726), .B2(n10725), .A(n10724), .ZN(n10732) );
  NOR2_X1 U13335 ( .A1(n10727), .A2(n15313), .ZN(n10728) );
  OR2_X1 U13336 ( .A1(n15369), .A2(n10728), .ZN(n10730) );
  NAND2_X1 U13337 ( .A1(n13515), .A2(n13851), .ZN(n10729) );
  NAND2_X1 U13338 ( .A1(n10730), .A2(n10729), .ZN(n15371) );
  NAND2_X1 U13339 ( .A1(n15371), .A2(n13883), .ZN(n10731) );
  OAI211_X1 U13340 ( .C1(n10733), .C2(n15368), .A(n10732), .B(n10731), .ZN(
        P2_U3265) );
  OR2_X1 U13341 ( .A1(n10734), .A2(n15606), .ZN(n15569) );
  NAND2_X1 U13342 ( .A1(n10736), .A2(n10735), .ZN(n15573) );
  AOI21_X1 U13343 ( .B1(n15556), .B2(n10738), .A(n15560), .ZN(n10739) );
  AOI211_X1 U13344 ( .C1(n11097), .C2(n15573), .A(n10740), .B(n10739), .ZN(
        n15570) );
  OAI21_X1 U13345 ( .B1(n15552), .B2(n15569), .A(n15570), .ZN(n10741) );
  AOI22_X1 U13346 ( .A1(n10741), .A2(n15566), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14938), .ZN(n10743) );
  AND2_X1 U13347 ( .A1(n15552), .A2(n11682), .ZN(n11037) );
  NAND2_X1 U13348 ( .A1(n15566), .A2(n11037), .ZN(n12704) );
  INV_X1 U13349 ( .A(n12704), .ZN(n11156) );
  NAND2_X1 U13350 ( .A1(n11156), .A2(n15573), .ZN(n10742) );
  OAI211_X1 U13351 ( .C1(n10744), .C2(n15566), .A(n10743), .B(n10742), .ZN(
        P3_U3232) );
  NAND2_X1 U13352 ( .A1(n11972), .A2(n12411), .ZN(n10749) );
  NAND2_X1 U13353 ( .A1(n12363), .A2(n14168), .ZN(n10748) );
  NAND2_X1 U13354 ( .A1(n10749), .A2(n10748), .ZN(n10750) );
  XNOR2_X1 U13355 ( .A(n10750), .B(n12413), .ZN(n10885) );
  AOI22_X1 U13356 ( .A1(n12412), .A2(n14168), .B1(n11972), .B2(n12363), .ZN(
        n10886) );
  XNOR2_X1 U13357 ( .A(n10885), .B(n10886), .ZN(n10751) );
  OAI211_X1 U13358 ( .C1(n6584), .C2(n10751), .A(n10889), .B(n14119), .ZN(
        n10757) );
  INV_X1 U13359 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n14243) );
  OAI22_X1 U13360 ( .A1(n14124), .A2(n10753), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14243), .ZN(n10754) );
  AOI21_X1 U13361 ( .B1(n10755), .B2(n14134), .A(n10754), .ZN(n10756) );
  OAI211_X1 U13362 ( .C1(n7090), .C2(n14128), .A(n10757), .B(n10756), .ZN(
        P1_U3239) );
  INV_X1 U13363 ( .A(n10758), .ZN(n10760) );
  NAND2_X1 U13364 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n10945), .ZN(n10761) );
  OAI21_X1 U13365 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n10945), .A(n10761), 
        .ZN(n10762) );
  AOI21_X1 U13366 ( .B1(n10763), .B2(n10762), .A(n10944), .ZN(n10764) );
  INV_X1 U13367 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14793) );
  OAI22_X1 U13368 ( .A1(n10764), .A2(n15547), .B1(n15529), .B2(n14793), .ZN(
        n10784) );
  INV_X1 U13369 ( .A(n10765), .ZN(n10767) );
  NAND2_X1 U13370 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10945), .ZN(n10768) );
  OAI21_X1 U13371 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n10945), .A(n10768), 
        .ZN(n10769) );
  AOI21_X1 U13372 ( .B1(n10770), .B2(n10769), .A(n10933), .ZN(n10771) );
  NOR2_X1 U13373 ( .A1(n10771), .A2(n15541), .ZN(n10783) );
  INV_X1 U13374 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10772) );
  MUX2_X1 U13375 ( .A(n11208), .B(n10772), .S(n13279), .Z(n10774) );
  NAND2_X1 U13376 ( .A1(n10774), .A2(n10773), .ZN(n10936) );
  INV_X1 U13377 ( .A(n10774), .ZN(n10775) );
  NAND2_X1 U13378 ( .A1(n10775), .A2(n10945), .ZN(n10776) );
  NAND2_X1 U13379 ( .A1(n10936), .A2(n10776), .ZN(n10777) );
  AOI21_X1 U13380 ( .B1(n10779), .B2(n10778), .A(n10777), .ZN(n10938) );
  AND3_X1 U13381 ( .A1(n10779), .A2(n10778), .A3(n10777), .ZN(n10780) );
  OAI21_X1 U13382 ( .B1(n10938), .B2(n10780), .A(n15538), .ZN(n10781) );
  NAND2_X1 U13383 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11270)
         );
  OAI211_X1 U13384 ( .C1(n15531), .C2(n10945), .A(n10781), .B(n11270), .ZN(
        n10782) );
  OR3_X1 U13385 ( .A1(n10784), .A2(n10783), .A3(n10782), .ZN(P3_U3192) );
  INV_X1 U13386 ( .A(n12052), .ZN(n10836) );
  NAND2_X1 U13387 ( .A1(n6729), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10785) );
  XNOR2_X1 U13388 ( .A(n10785), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14316) );
  INV_X1 U13389 ( .A(n14316), .ZN(n14310) );
  OAI222_X1 U13390 ( .A1(n12426), .A2(n10836), .B1(n14310), .B2(P1_U3086), 
        .C1(n10786), .C2(n12296), .ZN(P1_U3337) );
  INV_X1 U13391 ( .A(SI_21_), .ZN(n13175) );
  INV_X1 U13392 ( .A(n10787), .ZN(n10788) );
  OAI222_X1 U13393 ( .A1(P3_U3151), .A2(n10789), .B1(n13284), .B2(n13175), 
        .C1(n13282), .C2(n10788), .ZN(P3_U3274) );
  OAI211_X1 U13394 ( .C1(n10792), .C2(n10791), .A(n10790), .B(n15469), .ZN(
        n10796) );
  NOR2_X1 U13395 ( .A1(n12576), .A2(n15594), .ZN(n10794) );
  OAI22_X1 U13396 ( .A1(n11125), .A2(n11083), .B1(n15467), .B2(n11095), .ZN(
        n10793) );
  AOI211_X1 U13397 ( .C1(P3_REG3_REG_7__SCAN_IN), .C2(P3_U3151), .A(n10794), 
        .B(n10793), .ZN(n10795) );
  OAI211_X1 U13398 ( .C1(n10982), .C2(n12549), .A(n10796), .B(n10795), .ZN(
        P3_U3153) );
  NOR2_X1 U13399 ( .A1(n11983), .A2(n10907), .ZN(n10797) );
  NAND2_X1 U13400 ( .A1(n10800), .A2(n12234), .ZN(n10803) );
  AOI22_X1 U13401 ( .A1(n12223), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12066), 
        .B2(n10801), .ZN(n10802) );
  NAND2_X1 U13402 ( .A1(n10803), .A2(n10802), .ZN(n11987) );
  XNOR2_X1 U13403 ( .A(n11987), .B(n14165), .ZN(n12264) );
  INV_X1 U13404 ( .A(n14165), .ZN(n10804) );
  NAND2_X1 U13405 ( .A1(n11987), .A2(n10804), .ZN(n10805) );
  NAND2_X1 U13406 ( .A1(n10806), .A2(n12234), .ZN(n10808) );
  AOI22_X1 U13407 ( .A1(n12223), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12066), 
        .B2(n14273), .ZN(n10807) );
  NAND2_X1 U13408 ( .A1(n12147), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10813) );
  INV_X1 U13409 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10809) );
  OR2_X1 U13410 ( .A1(n12149), .A2(n10809), .ZN(n10812) );
  XNOR2_X1 U13411 ( .A(n10822), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n11401) );
  OR2_X1 U13412 ( .A1(n12202), .A2(n11401), .ZN(n10811) );
  OR2_X1 U13413 ( .A1(n12219), .A2(n13179), .ZN(n10810) );
  NAND4_X1 U13414 ( .A1(n10813), .A2(n10812), .A3(n10811), .A4(n10810), .ZN(
        n14164) );
  XNOR2_X1 U13415 ( .A(n15191), .B(n14164), .ZN(n12265) );
  AOI21_X1 U13416 ( .B1(n10814), .B2(n10819), .A(n15178), .ZN(n10815) );
  AOI22_X1 U13417 ( .A1(n10815), .A2(n10967), .B1(n14569), .B2(n14165), .ZN(
        n15193) );
  OR2_X1 U13418 ( .A1(n11983), .A2(n14166), .ZN(n10816) );
  INV_X1 U13419 ( .A(n12264), .ZN(n10902) );
  NAND2_X1 U13420 ( .A1(n10903), .A2(n10902), .ZN(n10901) );
  OR2_X1 U13421 ( .A1(n11987), .A2(n14165), .ZN(n10818) );
  NAND2_X1 U13422 ( .A1(n10901), .A2(n10818), .ZN(n10820) );
  NAND2_X1 U13423 ( .A1(n10820), .A2(n10819), .ZN(n10952) );
  OAI21_X1 U13424 ( .B1(n10820), .B2(n10819), .A(n10952), .ZN(n15197) );
  INV_X1 U13425 ( .A(n11987), .ZN(n11337) );
  AOI21_X1 U13426 ( .B1(n10821), .B2(n15191), .A(n15091), .ZN(n10830) );
  NAND2_X1 U13427 ( .A1(n12198), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10829) );
  OR2_X1 U13428 ( .A1(n11348), .A2(n15010), .ZN(n10828) );
  NAND2_X1 U13429 ( .A1(n10822), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10824) );
  INV_X1 U13430 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13431 ( .A1(n10824), .A2(n10823), .ZN(n10825) );
  NAND2_X1 U13432 ( .A1(n10825), .A2(n10960), .ZN(n11586) );
  OR2_X1 U13433 ( .A1(n12202), .A2(n11586), .ZN(n10827) );
  INV_X1 U13434 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10970) );
  OR2_X1 U13435 ( .A1(n12219), .A2(n10970), .ZN(n10826) );
  NAND4_X1 U13436 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n14163) );
  AND2_X1 U13437 ( .A1(n14163), .A2(n14570), .ZN(n11398) );
  AOI21_X1 U13438 ( .B1(n10830), .B2(n10969), .A(n11398), .ZN(n15192) );
  OAI22_X1 U13439 ( .A1(n14547), .A2(n13179), .B1(n11401), .B2(n14556), .ZN(
        n10831) );
  AOI21_X1 U13440 ( .B1(n14558), .B2(n15191), .A(n10831), .ZN(n10832) );
  OAI21_X1 U13441 ( .B1(n15192), .B2(n14543), .A(n10832), .ZN(n10833) );
  AOI21_X1 U13442 ( .B1(n15197), .B2(n14562), .A(n10833), .ZN(n10834) );
  OAI21_X1 U13443 ( .B1(n15098), .B2(n15193), .A(n10834), .ZN(P1_U3283) );
  INV_X1 U13444 ( .A(n13555), .ZN(n13539) );
  OAI222_X1 U13445 ( .A1(P2_U3088), .A2(n13539), .B1(n14022), .B2(n10836), 
        .C1(n10835), .C2(n14024), .ZN(P2_U3309) );
  INV_X1 U13446 ( .A(n14289), .ZN(n14279) );
  INV_X1 U13447 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13448 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14077)
         );
  OAI21_X1 U13449 ( .B1(n15075), .B2(n10837), .A(n14077), .ZN(n10848) );
  INV_X1 U13450 ( .A(n11169), .ZN(n10839) );
  AOI21_X1 U13451 ( .B1(n10839), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10838), 
        .ZN(n15049) );
  INV_X1 U13452 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10840) );
  MUX2_X1 U13453 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10840), .S(n15057), .Z(
        n10841) );
  INV_X1 U13454 ( .A(n10841), .ZN(n15048) );
  NOR2_X1 U13455 ( .A1(n15049), .A2(n15048), .ZN(n15047) );
  AOI21_X1 U13456 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n15057), .A(n15047), 
        .ZN(n10843) );
  NAND2_X1 U13457 ( .A1(n10843), .A2(n10842), .ZN(n10844) );
  XNOR2_X1 U13458 ( .A(n10843), .B(n15068), .ZN(n15066) );
  INV_X1 U13459 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15065) );
  NAND2_X1 U13460 ( .A1(n15066), .A2(n15065), .ZN(n15064) );
  NAND2_X1 U13461 ( .A1(n10844), .A2(n15064), .ZN(n10846) );
  XNOR2_X1 U13462 ( .A(n14279), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10845) );
  NOR2_X1 U13463 ( .A1(n10845), .A2(n10846), .ZN(n14278) );
  AOI211_X1 U13464 ( .C1(n10846), .C2(n10845), .A(n14278), .B(n15046), .ZN(
        n10847) );
  AOI211_X1 U13465 ( .C1(n15067), .C2(n14279), .A(n10848), .B(n10847), .ZN(
        n10858) );
  INV_X1 U13466 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U13467 ( .A1(n15057), .A2(n11190), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10852), .ZN(n15052) );
  OR2_X1 U13468 ( .A1(n10850), .A2(n10849), .ZN(n10851) );
  OAI21_X1 U13469 ( .B1(n11169), .B2(n11173), .A(n10851), .ZN(n15051) );
  NOR2_X1 U13470 ( .A1(n15052), .A2(n15051), .ZN(n15050) );
  AOI21_X1 U13471 ( .B1(n10852), .B2(n11190), .A(n15050), .ZN(n10853) );
  NOR2_X1 U13472 ( .A1(n15068), .A2(n10853), .ZN(n10854) );
  XNOR2_X1 U13473 ( .A(n10853), .B(n15068), .ZN(n15062) );
  NOR2_X1 U13474 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15062), .ZN(n15061) );
  NOR2_X1 U13475 ( .A1(n10854), .A2(n15061), .ZN(n10856) );
  XNOR2_X1 U13476 ( .A(n14289), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13477 ( .A1(n10855), .A2(n10856), .ZN(n14287) );
  OAI211_X1 U13478 ( .C1(n10856), .C2(n10855), .A(n15071), .B(n14287), .ZN(
        n10857) );
  NAND2_X1 U13479 ( .A1(n10858), .A2(n10857), .ZN(P1_U3259) );
  INV_X1 U13480 ( .A(n10859), .ZN(n10868) );
  INV_X1 U13481 ( .A(n10860), .ZN(n10861) );
  NAND2_X1 U13482 ( .A1(n15326), .A2(n10861), .ZN(n10863) );
  INV_X1 U13483 ( .A(n13880), .ZN(n15315) );
  AOI22_X1 U13484 ( .A1(n15316), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n15315), 
        .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10862) );
  OAI211_X1 U13485 ( .C1(n14957), .C2(n10864), .A(n10863), .B(n10862), .ZN(
        n10865) );
  AOI21_X1 U13486 ( .B1(n15327), .B2(n10866), .A(n10865), .ZN(n10867) );
  OAI21_X1 U13487 ( .B1(n10868), .B2(n15316), .A(n10867), .ZN(P2_U3264) );
  INV_X1 U13488 ( .A(n10869), .ZN(n10871) );
  OAI22_X1 U13489 ( .A1(n11841), .A2(P3_U3151), .B1(SI_22_), .B2(n13284), .ZN(
        n10870) );
  AOI21_X1 U13490 ( .B1(n10871), .B2(n14835), .A(n10870), .ZN(P3_U3273) );
  OAI222_X1 U13491 ( .A1(n12426), .A2(n12084), .B1(P1_U3086), .B2(n12222), 
        .C1(n10872), .C2(n12296), .ZN(P1_U3335) );
  XNOR2_X1 U13492 ( .A(n10873), .B(n10877), .ZN(n15590) );
  INV_X1 U13493 ( .A(n11097), .ZN(n11153) );
  OR2_X1 U13494 ( .A1(n11123), .A2(n11657), .ZN(n11121) );
  AND2_X1 U13495 ( .A1(n11121), .A2(n10874), .ZN(n10878) );
  NAND2_X1 U13496 ( .A1(n11121), .A2(n10875), .ZN(n10876) );
  OAI211_X1 U13497 ( .C1(n10878), .C2(n10877), .A(n10876), .B(n12861), .ZN(
        n10880) );
  AOI22_X1 U13498 ( .A1(n12849), .A2(n12599), .B1(n12597), .B2(n8165), .ZN(
        n10879) );
  OAI211_X1 U13499 ( .C1(n11153), .C2(n15590), .A(n10880), .B(n10879), .ZN(
        n15592) );
  NAND2_X1 U13500 ( .A1(n15592), .A2(n15566), .ZN(n10884) );
  OAI22_X1 U13501 ( .A1(n12870), .A2(n15589), .B1(n10881), .B2(n15553), .ZN(
        n10882) );
  AOI21_X1 U13502 ( .B1(n14943), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10882), .ZN(
        n10883) );
  OAI211_X1 U13503 ( .C1(n15590), .C2(n12704), .A(n10884), .B(n10883), .ZN(
        P3_U3227) );
  INV_X1 U13504 ( .A(n10886), .ZN(n10887) );
  NOR2_X1 U13505 ( .A1(n12369), .A2(n10890), .ZN(n10891) );
  AOI21_X1 U13506 ( .B1(n15170), .B2(n12329), .A(n10891), .ZN(n11131) );
  AOI22_X1 U13507 ( .A1(n15170), .A2(n12411), .B1(n12363), .B2(n14167), .ZN(
        n10892) );
  XNOR2_X1 U13508 ( .A(n10892), .B(n12413), .ZN(n11130) );
  XOR2_X1 U13509 ( .A(n11131), .B(n11130), .Z(n10893) );
  OAI211_X1 U13510 ( .C1(n10894), .C2(n10893), .A(n11135), .B(n14119), .ZN(
        n10900) );
  AND2_X1 U13511 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14259) );
  AOI21_X1 U13512 ( .B1(n14141), .B2(n14166), .A(n14259), .ZN(n10896) );
  NAND2_X1 U13513 ( .A1(n14140), .A2(n14168), .ZN(n10895) );
  OAI211_X1 U13514 ( .C1(n14998), .C2(n10897), .A(n10896), .B(n10895), .ZN(
        n10898) );
  AOI21_X1 U13515 ( .B1(n14995), .B2(n15170), .A(n10898), .ZN(n10899) );
  NAND2_X1 U13516 ( .A1(n10900), .A2(n10899), .ZN(P1_U3213) );
  OAI21_X1 U13517 ( .B1(n10903), .B2(n10902), .A(n10901), .ZN(n10904) );
  INV_X1 U13518 ( .A(n10904), .ZN(n15185) );
  OAI21_X1 U13519 ( .B1(n10906), .B2(n12264), .A(n10905), .ZN(n10909) );
  INV_X1 U13520 ( .A(n14164), .ZN(n11394) );
  OAI22_X1 U13521 ( .A1(n10907), .A2(n14591), .B1(n11394), .B2(n14593), .ZN(
        n10908) );
  AOI21_X1 U13522 ( .B1(n10909), .B2(n6917), .A(n10908), .ZN(n10910) );
  OAI21_X1 U13523 ( .B1(n15185), .B2(n10911), .A(n10910), .ZN(n15189) );
  NAND2_X1 U13524 ( .A1(n15189), .A2(n14547), .ZN(n10917) );
  XNOR2_X1 U13525 ( .A(n10912), .B(n11337), .ZN(n10913) );
  NOR2_X1 U13526 ( .A1(n10913), .A2(n15091), .ZN(n15186) );
  NOR2_X1 U13527 ( .A1(n15088), .A2(n11337), .ZN(n10915) );
  OAI22_X1 U13528 ( .A1(n14547), .A2(n9810), .B1(n11340), .B2(n14556), .ZN(
        n10914) );
  AOI211_X1 U13529 ( .C1(n15186), .C2(n15094), .A(n10915), .B(n10914), .ZN(
        n10916) );
  OAI211_X1 U13530 ( .C1(n15185), .C2(n10918), .A(n10917), .B(n10916), .ZN(
        P1_U3284) );
  INV_X1 U13531 ( .A(n12065), .ZN(n11898) );
  OAI222_X1 U13532 ( .A1(n14024), .A2(n10919), .B1(n14022), .B2(n11898), .C1(
        P2_U3088), .C2(n13565), .ZN(P2_U3308) );
  OAI222_X1 U13533 ( .A1(n14024), .A2(n10921), .B1(n14022), .B2(n12084), .C1(
        n10920), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI211_X1 U13534 ( .C1(n10924), .C2(n10923), .A(n10922), .B(n15469), .ZN(
        n10932) );
  INV_X1 U13535 ( .A(n10925), .ZN(n11047) );
  OAI22_X1 U13536 ( .A1(n12576), .A2(n15601), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10926), .ZN(n10930) );
  OAI22_X1 U13537 ( .A1(n10928), .A2(n11083), .B1(n15467), .B2(n10927), .ZN(
        n10929) );
  AOI211_X1 U13538 ( .C1(n11047), .C2(n12573), .A(n10930), .B(n10929), .ZN(
        n10931) );
  NAND2_X1 U13539 ( .A1(n10932), .A2(n10931), .ZN(P3_U3161) );
  INV_X1 U13540 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11323) );
  AOI21_X1 U13541 ( .B1(n11323), .B2(n10934), .A(n11059), .ZN(n10950) );
  INV_X1 U13542 ( .A(n14838), .ZN(n11058) );
  INV_X1 U13543 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13544 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11477)
         );
  OAI21_X1 U13545 ( .B1(n15529), .B2(n10935), .A(n11477), .ZN(n10943) );
  INV_X1 U13546 ( .A(n10936), .ZN(n10937) );
  NOR2_X1 U13547 ( .A1(n10938), .A2(n10937), .ZN(n10940) );
  MUX2_X1 U13548 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13279), .Z(n11069) );
  XNOR2_X1 U13549 ( .A(n11069), .B(n14838), .ZN(n10939) );
  AOI21_X1 U13550 ( .B1(n10940), .B2(n10939), .A(n11071), .ZN(n10941) );
  NOR2_X1 U13551 ( .A1(n10941), .A2(n14920), .ZN(n10942) );
  AOI211_X1 U13552 ( .C1(n14926), .C2(n11058), .A(n10943), .B(n10942), .ZN(
        n10949) );
  AOI21_X1 U13553 ( .B1(n11313), .B2(n10946), .A(n11051), .ZN(n10947) );
  OR2_X1 U13554 ( .A1(n10947), .A2(n15547), .ZN(n10948) );
  OAI211_X1 U13555 ( .C1(n10950), .C2(n15541), .A(n10949), .B(n10948), .ZN(
        P3_U3193) );
  OR2_X1 U13556 ( .A1(n15191), .A2(n14164), .ZN(n10951) );
  NAND2_X1 U13557 ( .A1(n10953), .A2(n12234), .ZN(n10955) );
  AOI22_X1 U13558 ( .A1(n12223), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12066), 
        .B2(n15037), .ZN(n10954) );
  XNOR2_X1 U13559 ( .A(n15005), .B(n14163), .ZN(n12267) );
  INV_X1 U13560 ( .A(n12267), .ZN(n10956) );
  OAI21_X1 U13561 ( .B1(n10957), .B2(n10956), .A(n11160), .ZN(n10958) );
  INV_X1 U13562 ( .A(n10958), .ZN(n15007) );
  NAND2_X1 U13563 ( .A1(n12198), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U13564 ( .A1(n10960), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U13565 ( .A1(n11186), .A2(n10961), .ZN(n11610) );
  OR2_X1 U13566 ( .A1(n12202), .A2(n11610), .ZN(n10964) );
  OR2_X1 U13567 ( .A1(n12219), .A2(n10098), .ZN(n10963) );
  OR2_X1 U13568 ( .A1(n11348), .A2(n14857), .ZN(n10962) );
  NAND4_X1 U13569 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n14162) );
  INV_X1 U13570 ( .A(n14162), .ZN(n11601) );
  OR2_X1 U13571 ( .A1(n15191), .A2(n11394), .ZN(n10966) );
  XNOR2_X1 U13572 ( .A(n11180), .B(n12267), .ZN(n10968) );
  OAI222_X1 U13573 ( .A1(n14593), .A2(n11601), .B1(n10968), .B2(n15178), .C1(
        n14591), .C2(n11394), .ZN(n15009) );
  NAND2_X1 U13574 ( .A1(n15009), .A2(n14547), .ZN(n10974) );
  AOI211_X1 U13575 ( .C1(n15005), .C2(n10969), .A(n15091), .B(n11245), .ZN(
        n15004) );
  NOR2_X1 U13576 ( .A1(n7095), .A2(n15088), .ZN(n10972) );
  OAI22_X1 U13577 ( .A1(n14547), .A2(n10970), .B1(n11586), .B2(n14556), .ZN(
        n10971) );
  AOI211_X1 U13578 ( .C1(n15004), .C2(n15094), .A(n10972), .B(n10971), .ZN(
        n10973) );
  OAI211_X1 U13579 ( .C1(n15007), .C2(n14601), .A(n10974), .B(n10973), .ZN(
        P1_U3282) );
  XNOR2_X1 U13580 ( .A(n10976), .B(n10975), .ZN(n15596) );
  XNOR2_X1 U13581 ( .A(n10977), .B(n11708), .ZN(n10980) );
  AOI22_X1 U13582 ( .A1(n12849), .A2(n12598), .B1(n12596), .B2(n8165), .ZN(
        n10978) );
  OAI21_X1 U13583 ( .B1(n15596), .B2(n11153), .A(n10978), .ZN(n10979) );
  AOI21_X1 U13584 ( .B1(n10980), .B2(n12861), .A(n10979), .ZN(n15593) );
  MUX2_X1 U13585 ( .A(n10981), .B(n15593), .S(n15566), .Z(n10986) );
  INV_X1 U13586 ( .A(n10982), .ZN(n10983) );
  AOI22_X1 U13587 ( .A1(n14944), .A2(n10984), .B1(n14938), .B2(n10983), .ZN(
        n10985) );
  OAI211_X1 U13588 ( .C1(n15596), .C2(n12704), .A(n10986), .B(n10985), .ZN(
        P3_U3226) );
  OR2_X1 U13589 ( .A1(n10988), .A2(n11658), .ZN(n10989) );
  NAND2_X1 U13590 ( .A1(n11146), .A2(n10989), .ZN(n10993) );
  INV_X1 U13591 ( .A(n10993), .ZN(n15578) );
  NAND2_X1 U13592 ( .A1(n10990), .A2(n11658), .ZN(n10991) );
  NAND3_X1 U13593 ( .A1(n10992), .A2(n12861), .A3(n10991), .ZN(n10996) );
  NAND2_X1 U13594 ( .A1(n10993), .A2(n11097), .ZN(n10995) );
  AOI22_X1 U13595 ( .A1(n12849), .A2(n6822), .B1(n12600), .B2(n8165), .ZN(
        n10994) );
  NAND3_X1 U13596 ( .A1(n10996), .A2(n10995), .A3(n10994), .ZN(n15579) );
  MUX2_X1 U13597 ( .A(n15579), .B(P3_REG2_REG_3__SCAN_IN), .S(n14943), .Z(
        n10997) );
  INV_X1 U13598 ( .A(n10997), .ZN(n11001) );
  AOI22_X1 U13599 ( .A1(n14944), .A2(n10999), .B1(n14938), .B2(n10998), .ZN(
        n11000) );
  OAI211_X1 U13600 ( .C1(n15578), .C2(n12704), .A(n11001), .B(n11000), .ZN(
        P3_U3230) );
  NOR2_X1 U13601 ( .A1(n15273), .A2(n11002), .ZN(n11003) );
  AOI21_X1 U13602 ( .B1(n11002), .B2(n15273), .A(n11003), .ZN(n15276) );
  AOI21_X1 U13603 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n11005), .A(n11004), 
        .ZN(n13518) );
  MUX2_X1 U13604 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13824), .S(n11019), .Z(
        n13517) );
  AND2_X1 U13605 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  AOI22_X1 U13606 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n11022), .B1(n15268), 
        .B2(n13804), .ZN(n15261) );
  NOR2_X1 U13607 ( .A1(n15262), .A2(n15261), .ZN(n15260) );
  AOI21_X1 U13608 ( .B1(n11022), .B2(n13804), .A(n15260), .ZN(n15277) );
  NAND2_X1 U13609 ( .A1(n15276), .A2(n15277), .ZN(n15275) );
  NAND2_X1 U13610 ( .A1(n11006), .A2(n11007), .ZN(n11008) );
  XNOR2_X1 U13611 ( .A(n15289), .B(n11007), .ZN(n15293) );
  NAND2_X1 U13612 ( .A1(n15299), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U13613 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15303), .ZN(n15301) );
  NAND2_X1 U13614 ( .A1(n11010), .A2(n15301), .ZN(n11014) );
  NAND2_X1 U13615 ( .A1(n11033), .A2(n8682), .ZN(n11012) );
  INV_X1 U13616 ( .A(n11012), .ZN(n11011) );
  AOI21_X1 U13617 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n11110), .A(n11011), 
        .ZN(n11013) );
  NAND2_X1 U13618 ( .A1(n11110), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11107) );
  OAI211_X1 U13619 ( .C1(n11014), .C2(n11013), .A(n11106), .B(n15302), .ZN(
        n11032) );
  NAND2_X1 U13620 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n13420)
         );
  INV_X1 U13621 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11015) );
  XNOR2_X1 U13622 ( .A(n11110), .B(n11015), .ZN(n11111) );
  NOR2_X1 U13623 ( .A1(n15289), .A2(n11016), .ZN(n11017) );
  AOI21_X1 U13624 ( .B1(n11016), .B2(n15289), .A(n11017), .ZN(n15286) );
  INV_X1 U13625 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15256) );
  NOR2_X1 U13626 ( .A1(n11022), .A2(n15256), .ZN(n11021) );
  NOR2_X1 U13627 ( .A1(n11018), .A2(n8578), .ZN(n13526) );
  MUX2_X1 U13628 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11020), .S(n11019), .Z(
        n13525) );
  OAI21_X1 U13629 ( .B1(n13527), .B2(n13526), .A(n13525), .ZN(n13529) );
  OAI21_X1 U13630 ( .B1(n11020), .B2(n13522), .A(n13529), .ZN(n15258) );
  AOI211_X1 U13631 ( .C1(n11022), .C2(n15256), .A(n11021), .B(n15258), .ZN(
        n15257) );
  AOI21_X1 U13632 ( .B1(n15256), .B2(n11022), .A(n15257), .ZN(n15280) );
  NOR2_X1 U13633 ( .A1(n15273), .A2(n11023), .ZN(n11024) );
  AOI21_X1 U13634 ( .B1(n11023), .B2(n15273), .A(n11024), .ZN(n15279) );
  NAND2_X1 U13635 ( .A1(n15280), .A2(n15279), .ZN(n15278) );
  OAI21_X1 U13636 ( .B1(n15273), .B2(n11023), .A(n15278), .ZN(n15285) );
  NAND2_X1 U13637 ( .A1(n15286), .A2(n15285), .ZN(n15284) );
  OAI21_X1 U13638 ( .B1(n15289), .B2(n11016), .A(n15284), .ZN(n11025) );
  NAND2_X1 U13639 ( .A1(n15299), .A2(n11025), .ZN(n11027) );
  XNOR2_X1 U13640 ( .A(n11026), .B(n11025), .ZN(n15306) );
  NAND2_X1 U13641 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15306), .ZN(n15304) );
  NAND2_X1 U13642 ( .A1(n11027), .A2(n15304), .ZN(n11112) );
  XOR2_X1 U13643 ( .A(n11111), .B(n11112), .Z(n11028) );
  NAND2_X1 U13644 ( .A1(n15305), .A2(n11028), .ZN(n11029) );
  NAND2_X1 U13645 ( .A1(n13420), .A2(n11029), .ZN(n11030) );
  AOI21_X1 U13646 ( .B1(n15298), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11030), 
        .ZN(n11031) );
  OAI211_X1 U13647 ( .C1(n15290), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        P2_U3230) );
  OAI222_X1 U13648 ( .A1(n12426), .A2(n12099), .B1(P1_U3086), .B2(n11925), 
        .C1(n11034), .C2(n12296), .ZN(P1_U3334) );
  OAI222_X1 U13649 ( .A1(n14024), .A2(n11036), .B1(n14022), .B2(n12099), .C1(
        n11035), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U13650 ( .A(n11040), .B(n11718), .ZN(n15603) );
  INV_X1 U13651 ( .A(n11718), .ZN(n11041) );
  XNOR2_X1 U13652 ( .A(n11042), .B(n11041), .ZN(n11043) );
  NAND2_X1 U13653 ( .A1(n11043), .A2(n12861), .ZN(n11045) );
  AOI22_X1 U13654 ( .A1(n12849), .A2(n12597), .B1(n12595), .B2(n8165), .ZN(
        n11044) );
  AND2_X1 U13655 ( .A1(n11045), .A2(n11044), .ZN(n15599) );
  MUX2_X1 U13656 ( .A(n15599), .B(n11046), .S(n14943), .Z(n11049) );
  AOI22_X1 U13657 ( .A1(n14944), .A2(n11721), .B1(n11047), .B2(n14938), .ZN(
        n11048) );
  OAI211_X1 U13658 ( .C1(n12857), .C2(n15603), .A(n11049), .B(n11048), .ZN(
        P3_U3225) );
  NOR2_X1 U13659 ( .A1(n11058), .A2(n11050), .ZN(n11052) );
  MUX2_X1 U13660 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n11053), .S(n11068), .Z(
        n11055) );
  INV_X1 U13661 ( .A(n12618), .ZN(n11054) );
  AOI21_X1 U13662 ( .B1(n11056), .B2(n11055), .A(n11054), .ZN(n11078) );
  NOR2_X1 U13663 ( .A1(n11058), .A2(n11057), .ZN(n11060) );
  INV_X1 U13664 ( .A(n11063), .ZN(n11065) );
  INV_X1 U13665 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11061) );
  MUX2_X1 U13666 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n11061), .S(n11068), .Z(
        n11062) );
  INV_X1 U13667 ( .A(n11062), .ZN(n11064) );
  OAI21_X1 U13668 ( .B1(n11065), .B2(n11064), .A(n12603), .ZN(n11076) );
  NAND2_X1 U13669 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n11067)
         );
  NAND2_X1 U13670 ( .A1(n15458), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11066) );
  OAI211_X1 U13671 ( .C1(n15531), .C2(n12616), .A(n11067), .B(n11066), .ZN(
        n11075) );
  MUX2_X1 U13672 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13279), .Z(n12609) );
  XOR2_X1 U13673 ( .A(n11068), .B(n12609), .Z(n11073) );
  NOR2_X1 U13674 ( .A1(n11069), .A2(n14838), .ZN(n11070) );
  OR2_X1 U13675 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  NOR3_X1 U13676 ( .A1(n11071), .A2(n11070), .A3(n11073), .ZN(n12608) );
  AOI211_X1 U13677 ( .C1(n11073), .C2(n11072), .A(n14920), .B(n12608), .ZN(
        n11074) );
  AOI211_X1 U13678 ( .C1(n14929), .C2(n11076), .A(n11075), .B(n11074), .ZN(
        n11077) );
  OAI21_X1 U13679 ( .B1(n11078), .B2(n15547), .A(n11077), .ZN(P3_U3194) );
  AOI21_X1 U13680 ( .B1(n11081), .B2(n11080), .A(n11079), .ZN(n11087) );
  OAI22_X1 U13681 ( .A1(n12576), .A2(n15607), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11082), .ZN(n11085) );
  OAI22_X1 U13682 ( .A1(n11095), .A2(n11083), .B1(n15467), .B2(n11094), .ZN(
        n11084) );
  AOI211_X1 U13683 ( .C1(n11100), .C2(n12573), .A(n11085), .B(n11084), .ZN(
        n11086) );
  OAI21_X1 U13684 ( .B1(n11087), .B2(n12552), .A(n11086), .ZN(P3_U3171) );
  NAND2_X1 U13685 ( .A1(n11088), .A2(n14835), .ZN(n11089) );
  OAI211_X1 U13686 ( .C1(n11090), .C2(n13284), .A(n11089), .B(n11843), .ZN(
        P3_U3272) );
  XNOR2_X1 U13687 ( .A(n11091), .B(n11092), .ZN(n11099) );
  XNOR2_X1 U13688 ( .A(n11093), .B(n11092), .ZN(n15610) );
  OAI22_X1 U13689 ( .A1(n11095), .A2(n15561), .B1(n11094), .B2(n15563), .ZN(
        n11096) );
  AOI21_X1 U13690 ( .B1(n15610), .B2(n11097), .A(n11096), .ZN(n11098) );
  OAI21_X1 U13691 ( .B1(n11099), .B2(n15560), .A(n11098), .ZN(n15608) );
  INV_X1 U13692 ( .A(n15608), .ZN(n11105) );
  AOI22_X1 U13693 ( .A1(n14944), .A2(n11101), .B1(n14938), .B2(n11100), .ZN(
        n11102) );
  OAI21_X1 U13694 ( .B1(n10423), .B2(n15566), .A(n11102), .ZN(n11103) );
  AOI21_X1 U13695 ( .B1(n15610), .B2(n11156), .A(n11103), .ZN(n11104) );
  OAI21_X1 U13696 ( .B1(n11105), .B2(n14943), .A(n11104), .ZN(P3_U3224) );
  AOI22_X1 U13697 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n13533), .B1(n13543), 
        .B2(n8699), .ZN(n11109) );
  NAND2_X1 U13698 ( .A1(n11109), .A2(n11108), .ZN(n13535) );
  OAI21_X1 U13699 ( .B1(n11109), .B2(n11108), .A(n13535), .ZN(n11117) );
  INV_X1 U13700 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U13701 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13433)
         );
  XNOR2_X1 U13702 ( .A(n13543), .B(n13542), .ZN(n13544) );
  AOI22_X1 U13703 ( .A1(n11112), .A2(n11111), .B1(n11110), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n13545) );
  XOR2_X1 U13704 ( .A(n13544), .B(n13545), .Z(n11113) );
  NAND2_X1 U13705 ( .A1(n11113), .A2(n15305), .ZN(n11114) );
  OAI211_X1 U13706 ( .C1(n14818), .C2(n15297), .A(n13433), .B(n11114), .ZN(
        n11115) );
  AOI21_X1 U13707 ( .B1(n15300), .B2(n13533), .A(n11115), .ZN(n11116) );
  OAI21_X1 U13708 ( .B1(n11117), .B2(n15263), .A(n11116), .ZN(P2_U3231) );
  OAI21_X1 U13709 ( .B1(n11119), .B2(n11657), .A(n11118), .ZN(n15588) );
  OAI22_X1 U13710 ( .A1(n12870), .A2(n15585), .B1(n11120), .B2(n15553), .ZN(
        n11127) );
  INV_X1 U13711 ( .A(n11121), .ZN(n11122) );
  AOI21_X1 U13712 ( .B1(n11657), .B2(n11123), .A(n11122), .ZN(n11124) );
  OAI222_X1 U13713 ( .A1(n15563), .A2(n11125), .B1(n15561), .B2(n7247), .C1(
        n15560), .C2(n11124), .ZN(n15586) );
  MUX2_X1 U13714 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15586), .S(n15566), .Z(
        n11126) );
  AOI211_X1 U13715 ( .C1(n12872), .C2(n15588), .A(n11127), .B(n11126), .ZN(
        n11128) );
  INV_X1 U13716 ( .A(n11128), .ZN(P3_U3228) );
  AOI22_X1 U13717 ( .A1(n11983), .A2(n12411), .B1(n12363), .B2(n14166), .ZN(
        n11129) );
  XNOR2_X1 U13718 ( .A(n11129), .B(n12413), .ZN(n11330) );
  AOI22_X1 U13719 ( .A1(n11983), .A2(n12363), .B1(n12412), .B2(n14166), .ZN(
        n11331) );
  XNOR2_X1 U13720 ( .A(n11330), .B(n11331), .ZN(n11139) );
  INV_X1 U13721 ( .A(n11130), .ZN(n11133) );
  INV_X1 U13722 ( .A(n11131), .ZN(n11132) );
  INV_X1 U13723 ( .A(n11333), .ZN(n11137) );
  AOI21_X1 U13724 ( .B1(n11139), .B2(n11138), .A(n11137), .ZN(n11145) );
  AOI22_X1 U13725 ( .A1(n14152), .A2(n11140), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11141) );
  OAI21_X1 U13726 ( .B1(n14998), .B2(n11142), .A(n11141), .ZN(n11143) );
  AOI21_X1 U13727 ( .B1(n14995), .B2(n11983), .A(n11143), .ZN(n11144) );
  OAI21_X1 U13728 ( .B1(n11145), .B2(n14989), .A(n11144), .ZN(P1_U3221) );
  NAND2_X1 U13729 ( .A1(n11146), .A2(n11693), .ZN(n11147) );
  XNOR2_X1 U13730 ( .A(n11147), .B(n11660), .ZN(n15582) );
  INV_X1 U13731 ( .A(n15582), .ZN(n11157) );
  OAI22_X1 U13732 ( .A1(n12870), .A2(n15581), .B1(n11148), .B2(n15553), .ZN(
        n11155) );
  XNOR2_X1 U13733 ( .A(n11149), .B(n11702), .ZN(n11150) );
  NAND2_X1 U13734 ( .A1(n11150), .A2(n12861), .ZN(n11152) );
  AOI22_X1 U13735 ( .A1(n8165), .A2(n12599), .B1(n15461), .B2(n12849), .ZN(
        n11151) );
  OAI211_X1 U13736 ( .C1(n11153), .C2(n15582), .A(n11152), .B(n11151), .ZN(
        n15584) );
  MUX2_X1 U13737 ( .A(n15584), .B(P3_REG2_REG_4__SCAN_IN), .S(n14943), .Z(
        n11154) );
  AOI211_X1 U13738 ( .C1(n11157), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n11158) );
  INV_X1 U13739 ( .A(n11158), .ZN(P3_U3229) );
  OR2_X1 U13740 ( .A1(n15005), .A2(n14163), .ZN(n11159) );
  NAND2_X1 U13741 ( .A1(n11160), .A2(n11159), .ZN(n11250) );
  NAND2_X1 U13742 ( .A1(n11161), .A2(n12234), .ZN(n11164) );
  AOI22_X1 U13743 ( .A1(n12223), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n12066), 
        .B2(n11162), .ZN(n11163) );
  XNOR2_X1 U13744 ( .A(n12002), .B(n11601), .ZN(n12270) );
  OR2_X1 U13745 ( .A1(n12002), .A2(n14162), .ZN(n11165) );
  NAND2_X1 U13746 ( .A1(n11166), .A2(n12234), .ZN(n11172) );
  OAI22_X1 U13747 ( .A1(n11169), .A2(n11922), .B1(n11168), .B2(n11167), .ZN(
        n11170) );
  INV_X1 U13748 ( .A(n11170), .ZN(n11171) );
  NAND2_X1 U13749 ( .A1(n12218), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11178) );
  INV_X1 U13750 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11173) );
  OR2_X1 U13751 ( .A1(n11348), .A2(n11173), .ZN(n11177) );
  INV_X1 U13752 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11174) );
  XNOR2_X1 U13753 ( .A(n11186), .B(n11174), .ZN(n14109) );
  OR2_X1 U13754 ( .A1(n12202), .A2(n14109), .ZN(n11176) );
  OR2_X1 U13755 ( .A1(n12219), .A2(n10260), .ZN(n11175) );
  NAND4_X1 U13756 ( .A1(n11178), .A2(n11177), .A3(n11176), .A4(n11175), .ZN(
        n14161) );
  XNOR2_X1 U13757 ( .A(n12311), .B(n14981), .ZN(n12269) );
  OAI21_X1 U13758 ( .B1(n11179), .B2(n12269), .A(n11363), .ZN(n15003) );
  INV_X1 U13759 ( .A(n15003), .ZN(n11201) );
  AOI22_X1 U13760 ( .A1(n12311), .A2(n14558), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n15098), .ZN(n11200) );
  INV_X1 U13761 ( .A(n14163), .ZN(n11251) );
  OR2_X1 U13762 ( .A1(n15005), .A2(n11251), .ZN(n11181) );
  NAND2_X1 U13763 ( .A1(n11182), .A2(n11181), .ZN(n11248) );
  INV_X1 U13764 ( .A(n12270), .ZN(n11247) );
  NAND2_X1 U13765 ( .A1(n11248), .A2(n11247), .ZN(n11184) );
  OR2_X1 U13766 ( .A1(n12002), .A2(n11601), .ZN(n11183) );
  NAND2_X1 U13767 ( .A1(n11184), .A2(n11183), .ZN(n11355) );
  XNOR2_X1 U13768 ( .A(n11355), .B(n12269), .ZN(n11185) );
  NAND2_X1 U13769 ( .A1(n11185), .A2(n6917), .ZN(n11196) );
  INV_X1 U13770 ( .A(n11186), .ZN(n11187) );
  AOI21_X1 U13771 ( .B1(n11187), .B2(P1_REG3_REG_13__SCAN_IN), .A(
        P1_REG3_REG_14__SCAN_IN), .ZN(n11188) );
  OR2_X1 U13772 ( .A1(n11188), .A2(n11345), .ZN(n14997) );
  OR2_X1 U13773 ( .A1(n14997), .A2(n12202), .ZN(n11194) );
  INV_X1 U13774 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11189) );
  OR2_X1 U13775 ( .A1(n12149), .A2(n11189), .ZN(n11193) );
  OR2_X1 U13776 ( .A1(n12219), .A2(n10840), .ZN(n11192) );
  OR2_X1 U13777 ( .A1(n11348), .A2(n11190), .ZN(n11191) );
  NAND4_X1 U13778 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(
        n14160) );
  AOI22_X1 U13779 ( .A1(n14569), .A2(n14162), .B1(n14160), .B2(n14570), .ZN(
        n11195) );
  NAND2_X1 U13780 ( .A1(n11196), .A2(n11195), .ZN(n15001) );
  INV_X1 U13781 ( .A(n11197), .ZN(n11246) );
  INV_X1 U13782 ( .A(n12311), .ZN(n15000) );
  OR2_X1 U13783 ( .A1(n11197), .A2(n12311), .ZN(n11366) );
  OAI211_X1 U13784 ( .C1(n11246), .C2(n15000), .A(n14538), .B(n11366), .ZN(
        n14999) );
  OAI22_X1 U13785 ( .A1(n14999), .A2(n14445), .B1(n14556), .B2(n14109), .ZN(
        n11198) );
  OAI21_X1 U13786 ( .B1(n15001), .B2(n11198), .A(n14547), .ZN(n11199) );
  OAI211_X1 U13787 ( .C1(n11201), .C2(n14601), .A(n11200), .B(n11199), .ZN(
        P1_U3280) );
  OAI211_X1 U13788 ( .C1(n6726), .C2(n11731), .A(n12861), .B(n11202), .ZN(
        n11205) );
  NAND2_X1 U13789 ( .A1(n12595), .A2(n12849), .ZN(n11204) );
  NAND2_X1 U13790 ( .A1(n12593), .A2(n8165), .ZN(n11203) );
  AND2_X1 U13791 ( .A1(n11204), .A2(n11203), .ZN(n11271) );
  NAND2_X1 U13792 ( .A1(n11205), .A2(n11271), .ZN(n11277) );
  INV_X1 U13793 ( .A(n11277), .ZN(n11212) );
  OAI21_X1 U13794 ( .B1(n11207), .B2(n11664), .A(n11206), .ZN(n11278) );
  NOR2_X1 U13795 ( .A1(n15566), .A2(n11208), .ZN(n11210) );
  OAI22_X1 U13796 ( .A1(n12870), .A2(n11281), .B1(n11276), .B2(n15553), .ZN(
        n11209) );
  AOI211_X1 U13797 ( .C1(n11278), .C2(n12872), .A(n11210), .B(n11209), .ZN(
        n11211) );
  OAI21_X1 U13798 ( .B1(n11212), .B2(n14943), .A(n11211), .ZN(P3_U3223) );
  XNOR2_X1 U13799 ( .A(n13889), .B(n13384), .ZN(n11876) );
  NAND2_X1 U13800 ( .A1(n13853), .A2(n13318), .ZN(n11215) );
  XNOR2_X1 U13801 ( .A(n11876), .B(n11215), .ZN(n11892) );
  INV_X1 U13802 ( .A(n11876), .ZN(n11216) );
  NAND2_X1 U13803 ( .A1(n11216), .A2(n11215), .ZN(n11217) );
  NAND2_X1 U13804 ( .A1(n11897), .A2(n11217), .ZN(n11218) );
  XNOR2_X1 U13805 ( .A(n13865), .B(n13384), .ZN(n11219) );
  NAND2_X1 U13806 ( .A1(n13508), .A2(n13318), .ZN(n11220) );
  XNOR2_X1 U13807 ( .A(n11219), .B(n11220), .ZN(n11877) );
  INV_X1 U13808 ( .A(n11219), .ZN(n11221) );
  NAND2_X1 U13809 ( .A1(n11221), .A2(n11220), .ZN(n11222) );
  XNOR2_X1 U13810 ( .A(n13845), .B(n13384), .ZN(n11223) );
  AND2_X1 U13811 ( .A1(n13852), .A2(n13318), .ZN(n11224) );
  NAND2_X1 U13812 ( .A1(n11223), .A2(n11224), .ZN(n11227) );
  INV_X1 U13813 ( .A(n11223), .ZN(n11285) );
  INV_X1 U13814 ( .A(n11224), .ZN(n11225) );
  NAND2_X1 U13815 ( .A1(n11285), .A2(n11225), .ZN(n11226) );
  NAND2_X1 U13816 ( .A1(n11227), .A2(n11226), .ZN(n11263) );
  XNOR2_X1 U13817 ( .A(n15435), .B(n13384), .ZN(n11229) );
  NAND2_X1 U13818 ( .A1(n13798), .A2(n13318), .ZN(n11230) );
  XNOR2_X1 U13819 ( .A(n11229), .B(n11230), .ZN(n11294) );
  AND2_X1 U13820 ( .A1(n11294), .A2(n11227), .ZN(n11228) );
  INV_X1 U13821 ( .A(n11229), .ZN(n11231) );
  NAND2_X1 U13822 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  XNOR2_X1 U13823 ( .A(n13808), .B(n13336), .ZN(n11233) );
  NAND2_X1 U13824 ( .A1(n13814), .A2(n13318), .ZN(n11234) );
  AND2_X1 U13825 ( .A1(n11233), .A2(n11234), .ZN(n11297) );
  INV_X1 U13826 ( .A(n11297), .ZN(n11237) );
  INV_X1 U13827 ( .A(n11233), .ZN(n11236) );
  INV_X1 U13828 ( .A(n11234), .ZN(n11235) );
  NAND2_X1 U13829 ( .A1(n11236), .A2(n11235), .ZN(n11296) );
  NAND2_X1 U13830 ( .A1(n11237), .A2(n11296), .ZN(n11238) );
  XNOR2_X1 U13831 ( .A(n11298), .B(n11238), .ZN(n11244) );
  NAND2_X1 U13832 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15269)
         );
  OAI21_X1 U13833 ( .B1(n11239), .B2(n13421), .A(n15269), .ZN(n11240) );
  AOI21_X1 U13834 ( .B1(n13452), .B2(n13798), .A(n11240), .ZN(n11241) );
  OAI21_X1 U13835 ( .B1(n13803), .B2(n15226), .A(n11241), .ZN(n11242) );
  AOI21_X1 U13836 ( .B1(n13808), .B2(n15223), .A(n11242), .ZN(n11243) );
  OAI21_X1 U13837 ( .B1(n11244), .B2(n13480), .A(n11243), .ZN(P2_U3196) );
  AOI211_X1 U13838 ( .C1(n12002), .C2(n7097), .A(n15091), .B(n11246), .ZN(
        n14850) );
  XNOR2_X1 U13839 ( .A(n11248), .B(n11247), .ZN(n11254) );
  OAI21_X1 U13840 ( .B1(n11250), .B2(n12270), .A(n11249), .ZN(n14855) );
  OAI22_X1 U13841 ( .A1(n11251), .A2(n14591), .B1(n14981), .B2(n14593), .ZN(
        n11252) );
  AOI21_X1 U13842 ( .B1(n14855), .B2(n15084), .A(n11252), .ZN(n11253) );
  OAI21_X1 U13843 ( .B1(n15178), .B2(n11254), .A(n11253), .ZN(n14853) );
  AOI21_X1 U13844 ( .B1(n14850), .B2(n9547), .A(n14853), .ZN(n11258) );
  NOR2_X1 U13845 ( .A1(n14852), .A2(n15088), .ZN(n11256) );
  OAI22_X1 U13846 ( .A1(n14547), .A2(n10098), .B1(n11610), .B2(n14556), .ZN(
        n11255) );
  AOI211_X1 U13847 ( .C1(n14855), .C2(n15095), .A(n11256), .B(n11255), .ZN(
        n11257) );
  OAI21_X1 U13848 ( .B1(n11258), .B2(n15086), .A(n11257), .ZN(P1_U3281) );
  OAI21_X1 U13849 ( .B1(n13835), .B2(n13421), .A(n11259), .ZN(n11260) );
  AOI21_X1 U13850 ( .B1(n13452), .B2(n13508), .A(n11260), .ZN(n11261) );
  OAI21_X1 U13851 ( .B1(n13839), .B2(n15226), .A(n11261), .ZN(n11265) );
  AOI211_X1 U13852 ( .C1(n11263), .C2(n11262), .A(n13480), .B(n6722), .ZN(
        n11264) );
  AOI211_X1 U13853 ( .C1(n13845), .C2(n15223), .A(n11265), .B(n11264), .ZN(
        n11266) );
  INV_X1 U13854 ( .A(n11266), .ZN(P2_U3189) );
  OAI211_X1 U13855 ( .C1(n11269), .C2(n11268), .A(n11267), .B(n15469), .ZN(
        n11275) );
  OAI21_X1 U13856 ( .B1(n12571), .B2(n11271), .A(n11270), .ZN(n11272) );
  AOI21_X1 U13857 ( .B1(n11273), .B2(n15463), .A(n11272), .ZN(n11274) );
  OAI211_X1 U13858 ( .C1(n11276), .C2(n12549), .A(n11275), .B(n11274), .ZN(
        P3_U3157) );
  AOI21_X1 U13859 ( .B1(n15600), .B2(n11278), .A(n11277), .ZN(n11284) );
  OAI22_X1 U13860 ( .A1(n13211), .A2(n11281), .B1(n15631), .B2(n10772), .ZN(
        n11279) );
  INV_X1 U13861 ( .A(n11279), .ZN(n11280) );
  OAI21_X1 U13862 ( .B1(n11284), .B2(n15628), .A(n11280), .ZN(P3_U3469) );
  OAI22_X1 U13863 ( .A1(n13263), .A2(n11281), .B1(n15613), .B2(n7894), .ZN(
        n11282) );
  INV_X1 U13864 ( .A(n11282), .ZN(n11283) );
  OAI21_X1 U13865 ( .B1(n11284), .B2(n15612), .A(n11283), .ZN(P3_U3420) );
  NOR3_X1 U13866 ( .A1(n11285), .A2(n11287), .A3(n13483), .ZN(n11286) );
  AOI21_X1 U13867 ( .B1(n6722), .B2(n13492), .A(n11286), .ZN(n11295) );
  NAND2_X1 U13868 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n13521)
         );
  OAI21_X1 U13869 ( .B1(n11287), .B2(n13409), .A(n13521), .ZN(n11288) );
  AOI21_X1 U13870 ( .B1(n13451), .B2(n13814), .A(n11288), .ZN(n11289) );
  OAI21_X1 U13871 ( .B1(n13823), .B2(n15226), .A(n11289), .ZN(n11292) );
  NOR2_X1 U13872 ( .A1(n11290), .A2(n13480), .ZN(n11291) );
  AOI211_X1 U13873 ( .C1(n15435), .C2(n15223), .A(n11292), .B(n11291), .ZN(
        n11293) );
  OAI21_X1 U13874 ( .B1(n11295), .B2(n11294), .A(n11293), .ZN(P2_U3208) );
  XNOR2_X1 U13875 ( .A(n11454), .B(n13384), .ZN(n11494) );
  NAND2_X1 U13876 ( .A1(n13797), .A2(n13318), .ZN(n11492) );
  XNOR2_X1 U13877 ( .A(n11494), .B(n11492), .ZN(n11490) );
  XNOR2_X1 U13878 ( .A(n11299), .B(n11490), .ZN(n11305) );
  NAND2_X1 U13879 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15272)
         );
  OAI21_X1 U13880 ( .B1(n11300), .B2(n13421), .A(n15272), .ZN(n11301) );
  AOI21_X1 U13881 ( .B1(n13452), .B2(n13814), .A(n11301), .ZN(n11302) );
  OAI21_X1 U13882 ( .B1(n11377), .B2(n15226), .A(n11302), .ZN(n11303) );
  AOI21_X1 U13883 ( .B1(n11454), .B2(n15223), .A(n11303), .ZN(n11304) );
  OAI21_X1 U13884 ( .B1(n11305), .B2(n13480), .A(n11304), .ZN(P2_U3206) );
  XNOR2_X1 U13885 ( .A(n11306), .B(n11742), .ZN(n11309) );
  OR2_X1 U13886 ( .A1(n11517), .A2(n15563), .ZN(n11308) );
  NAND2_X1 U13887 ( .A1(n12594), .A2(n12849), .ZN(n11307) );
  AND2_X1 U13888 ( .A1(n11308), .A2(n11307), .ZN(n11478) );
  OAI21_X1 U13889 ( .B1(n11309), .B2(n15560), .A(n11478), .ZN(n11321) );
  INV_X1 U13890 ( .A(n11321), .ZN(n11317) );
  OAI21_X1 U13891 ( .B1(n11312), .B2(n11311), .A(n11310), .ZN(n11322) );
  NOR2_X1 U13892 ( .A1(n15566), .A2(n11313), .ZN(n11315) );
  OAI22_X1 U13893 ( .A1(n12870), .A2(n11326), .B1(n11479), .B2(n15553), .ZN(
        n11314) );
  AOI211_X1 U13894 ( .C1(n11322), .C2(n12872), .A(n11315), .B(n11314), .ZN(
        n11316) );
  OAI21_X1 U13895 ( .B1(n11317), .B2(n14943), .A(n11316), .ZN(P3_U3222) );
  OAI222_X1 U13896 ( .A1(n14024), .A2(n11320), .B1(P2_U3088), .B2(n6783), .C1(
        n14022), .C2(n11318), .ZN(P2_U3305) );
  AOI21_X1 U13897 ( .B1(n15600), .B2(n11322), .A(n11321), .ZN(n11329) );
  OAI22_X1 U13898 ( .A1(n13211), .A2(n11326), .B1(n15631), .B2(n11323), .ZN(
        n11324) );
  INV_X1 U13899 ( .A(n11324), .ZN(n11325) );
  OAI21_X1 U13900 ( .B1(n11329), .B2(n15628), .A(n11325), .ZN(P3_U3470) );
  OAI22_X1 U13901 ( .A1(n13263), .A2(n11326), .B1(n15613), .B2(n7907), .ZN(
        n11327) );
  INV_X1 U13902 ( .A(n11327), .ZN(n11328) );
  OAI21_X1 U13903 ( .B1(n11329), .B2(n15612), .A(n11328), .ZN(P3_U3423) );
  NAND2_X1 U13904 ( .A1(n11330), .A2(n11331), .ZN(n11332) );
  NAND2_X1 U13905 ( .A1(n11987), .A2(n12363), .ZN(n11335) );
  NAND2_X1 U13906 ( .A1(n12412), .A2(n14165), .ZN(n11334) );
  NAND2_X1 U13907 ( .A1(n11335), .A2(n11334), .ZN(n11386) );
  AOI22_X1 U13908 ( .A1(n11987), .A2(n12411), .B1(n12363), .B2(n14165), .ZN(
        n11336) );
  XNOR2_X1 U13909 ( .A(n11336), .B(n12413), .ZN(n11389) );
  XOR2_X1 U13910 ( .A(n11390), .B(n11389), .Z(n11344) );
  NOR2_X1 U13911 ( .A1(n11337), .A2(n15194), .ZN(n15187) );
  AOI22_X1 U13912 ( .A1(n14140), .A2(n14166), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11339) );
  NAND2_X1 U13913 ( .A1(n14141), .A2(n14164), .ZN(n11338) );
  OAI211_X1 U13914 ( .C1(n14998), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        n11341) );
  AOI21_X1 U13915 ( .B1(n11342), .B2(n15187), .A(n11341), .ZN(n11343) );
  OAI21_X1 U13916 ( .B1(n11344), .B2(n14989), .A(n11343), .ZN(P1_U3231) );
  NOR2_X1 U13917 ( .A1(n11345), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11346) );
  OR2_X1 U13918 ( .A1(n11437), .A2(n11346), .ZN(n14154) );
  INV_X1 U13919 ( .A(n14154), .ZN(n11347) );
  NAND2_X1 U13920 ( .A1(n12092), .A2(n11347), .ZN(n11353) );
  INV_X1 U13921 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n13146) );
  OR2_X1 U13922 ( .A1(n11348), .A2(n13146), .ZN(n11352) );
  INV_X1 U13923 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11349) );
  OR2_X1 U13924 ( .A1(n12149), .A2(n11349), .ZN(n11351) );
  OR2_X1 U13925 ( .A1(n12219), .A2(n15065), .ZN(n11350) );
  NAND4_X1 U13926 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n14159) );
  INV_X1 U13927 ( .A(n14159), .ZN(n14984) );
  INV_X1 U13928 ( .A(n12269), .ZN(n11354) );
  NAND2_X1 U13929 ( .A1(n11355), .A2(n11354), .ZN(n11357) );
  OR2_X1 U13930 ( .A1(n12311), .A2(n14981), .ZN(n11356) );
  NAND2_X1 U13931 ( .A1(n11357), .A2(n11356), .ZN(n11435) );
  NAND2_X1 U13932 ( .A1(n11358), .A2(n12234), .ZN(n11360) );
  AOI22_X1 U13933 ( .A1(n15057), .A2(n12066), .B1(n12223), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11359) );
  NAND2_X2 U13934 ( .A1(n11360), .A2(n11359), .ZN(n14994) );
  INV_X1 U13935 ( .A(n14160), .ZN(n14111) );
  OR2_X1 U13936 ( .A1(n14994), .A2(n14111), .ZN(n12017) );
  NAND2_X1 U13937 ( .A1(n14994), .A2(n14111), .ZN(n12011) );
  XNOR2_X1 U13938 ( .A(n11435), .B(n12253), .ZN(n11361) );
  OAI222_X1 U13939 ( .A1(n14593), .A2(n14984), .B1(n14591), .B2(n14981), .C1(
        n15178), .C2(n11361), .ZN(n11419) );
  INV_X1 U13940 ( .A(n11419), .ZN(n11373) );
  OR2_X1 U13941 ( .A1(n12311), .A2(n14161), .ZN(n11362) );
  INV_X1 U13942 ( .A(n11431), .ZN(n11364) );
  AOI21_X1 U13943 ( .B1(n12253), .B2(n11365), .A(n11364), .ZN(n11421) );
  AOI21_X1 U13944 ( .B1(n14994), .B2(n11366), .A(n15091), .ZN(n11367) );
  OR2_X1 U13945 ( .A1(n14994), .A2(n11366), .ZN(n11446) );
  NAND2_X1 U13946 ( .A1(n11367), .A2(n11446), .ZN(n11417) );
  NAND2_X1 U13947 ( .A1(n15086), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11368) );
  OAI21_X1 U13948 ( .B1(n14556), .B2(n14997), .A(n11368), .ZN(n11369) );
  AOI21_X1 U13949 ( .B1(n14994), .B2(n14558), .A(n11369), .ZN(n11370) );
  OAI21_X1 U13950 ( .B1(n11417), .B2(n14543), .A(n11370), .ZN(n11371) );
  AOI21_X1 U13951 ( .B1(n11421), .B2(n14562), .A(n11371), .ZN(n11372) );
  OAI21_X1 U13952 ( .B1(n15086), .B2(n11373), .A(n11372), .ZN(P1_U3279) );
  XNOR2_X1 U13953 ( .A(n11374), .B(n11381), .ZN(n11375) );
  AOI222_X1 U13954 ( .A1(n15313), .A2(n11375), .B1(n13506), .B2(n13851), .C1(
        n13814), .C2(n13854), .ZN(n11456) );
  INV_X1 U13955 ( .A(n11376), .ZN(n13805) );
  AOI211_X1 U13956 ( .C1(n11454), .C2(n13805), .A(n13979), .B(n13788), .ZN(
        n11453) );
  INV_X1 U13957 ( .A(n11377), .ZN(n11378) );
  AOI22_X1 U13958 ( .A1(n15316), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n15315), 
        .B2(n11378), .ZN(n11379) );
  OAI21_X1 U13959 ( .B1(n11380), .B2(n14957), .A(n11379), .ZN(n11384) );
  XNOR2_X1 U13960 ( .A(n11382), .B(n11381), .ZN(n11457) );
  NOR2_X1 U13961 ( .A1(n11457), .A2(n14959), .ZN(n11383) );
  AOI211_X1 U13962 ( .C1(n11453), .C2(n15326), .A(n11384), .B(n11383), .ZN(
        n11385) );
  OAI21_X1 U13963 ( .B1(n11456), .B2(n15316), .A(n11385), .ZN(P2_U3252) );
  INV_X1 U13964 ( .A(n11386), .ZN(n11387) );
  NAND2_X1 U13965 ( .A1(n15191), .A2(n12411), .ZN(n11392) );
  NAND2_X1 U13966 ( .A1(n12363), .A2(n14164), .ZN(n11391) );
  NAND2_X1 U13967 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  XNOR2_X1 U13968 ( .A(n11393), .B(n12327), .ZN(n11575) );
  NOR2_X1 U13969 ( .A1(n12369), .A2(n11394), .ZN(n11395) );
  AOI21_X1 U13970 ( .B1(n15191), .B2(n12329), .A(n11395), .ZN(n11576) );
  XNOR2_X1 U13971 ( .A(n11575), .B(n11576), .ZN(n11396) );
  OAI211_X1 U13972 ( .C1(n11397), .C2(n11396), .A(n11578), .B(n14119), .ZN(
        n11404) );
  AND2_X1 U13973 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14268) );
  AOI21_X1 U13974 ( .B1(n14152), .B2(n11398), .A(n14268), .ZN(n11400) );
  NAND2_X1 U13975 ( .A1(n14140), .A2(n14165), .ZN(n11399) );
  OAI211_X1 U13976 ( .C1(n14998), .C2(n11401), .A(n11400), .B(n11399), .ZN(
        n11402) );
  AOI21_X1 U13977 ( .B1(n14995), .B2(n15191), .A(n11402), .ZN(n11403) );
  NAND2_X1 U13978 ( .A1(n11404), .A2(n11403), .ZN(P1_U3217) );
  INV_X1 U13979 ( .A(n11410), .ZN(n11668) );
  XNOR2_X1 U13980 ( .A(n11405), .B(n11668), .ZN(n11408) );
  OR2_X1 U13981 ( .A1(n11899), .A2(n15563), .ZN(n11407) );
  NAND2_X1 U13982 ( .A1(n12593), .A2(n12849), .ZN(n11406) );
  AND2_X1 U13983 ( .A1(n11407), .A2(n11406), .ZN(n11509) );
  OAI21_X1 U13984 ( .B1(n11408), .B2(n15560), .A(n11509), .ZN(n11552) );
  INV_X1 U13985 ( .A(n11552), .ZN(n11416) );
  OAI21_X1 U13986 ( .B1(n11411), .B2(n11410), .A(n11409), .ZN(n11553) );
  INV_X1 U13987 ( .A(n11412), .ZN(n11512) );
  AOI22_X1 U13988 ( .A1(n14943), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n14938), 
        .B2(n11512), .ZN(n11413) );
  OAI21_X1 U13989 ( .B1(n11557), .B2(n12870), .A(n11413), .ZN(n11414) );
  AOI21_X1 U13990 ( .B1(n11553), .B2(n12872), .A(n11414), .ZN(n11415) );
  OAI21_X1 U13991 ( .B1(n11416), .B2(n14943), .A(n11415), .ZN(P3_U3221) );
  INV_X1 U13992 ( .A(n14994), .ZN(n11418) );
  OAI21_X1 U13993 ( .B1(n11418), .B2(n15194), .A(n11417), .ZN(n11420) );
  AOI211_X1 U13994 ( .C1(n11421), .C2(n15198), .A(n11420), .B(n11419), .ZN(
        n11424) );
  NAND2_X1 U13995 ( .A1(n15210), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11422) );
  OAI21_X1 U13996 ( .B1(n11424), .B2(n15210), .A(n11422), .ZN(P1_U3542) );
  NAND2_X1 U13997 ( .A1(n15199), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11423) );
  OAI21_X1 U13998 ( .B1(n11424), .B2(n15199), .A(n11423), .ZN(P1_U3501) );
  INV_X1 U13999 ( .A(n12111), .ZN(n11426) );
  NAND2_X1 U14000 ( .A1(n14717), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11425) );
  OAI211_X1 U14001 ( .C1(n11426), .C2(n12426), .A(n12293), .B(n11425), .ZN(
        P1_U3332) );
  INV_X1 U14002 ( .A(n14022), .ZN(n14008) );
  NAND2_X1 U14003 ( .A1(n12111), .A2(n14008), .ZN(n11428) );
  OAI211_X1 U14004 ( .C1(n11429), .C2(n14024), .A(n11428), .B(n11427), .ZN(
        P2_U3304) );
  NAND2_X1 U14005 ( .A1(n14994), .A2(n14160), .ZN(n11430) );
  NAND2_X1 U14006 ( .A1(n11432), .A2(n12234), .ZN(n11434) );
  AOI22_X1 U14007 ( .A1(n12223), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12066), 
        .B2(n15068), .ZN(n11433) );
  NAND2_X1 U14008 ( .A1(n14156), .A2(n14984), .ZN(n12032) );
  NAND2_X1 U14009 ( .A1(n12031), .A2(n12032), .ZN(n12272) );
  XNOR2_X1 U14010 ( .A(n11533), .B(n11532), .ZN(n11469) );
  INV_X1 U14011 ( .A(n11469), .ZN(n11452) );
  NAND2_X1 U14012 ( .A1(n11435), .A2(n12253), .ZN(n11436) );
  XNOR2_X1 U14013 ( .A(n11529), .B(n12272), .ZN(n11445) );
  OR2_X1 U14014 ( .A1(n11437), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11438) );
  AND2_X1 U14015 ( .A1(n11538), .A2(n11438), .ZN(n14079) );
  NAND2_X1 U14016 ( .A1(n14079), .A2(n12092), .ZN(n11442) );
  NAND2_X1 U14017 ( .A1(n12147), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14018 ( .A1(n12198), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U14019 ( .A1(n12199), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11439) );
  NAND4_X1 U14020 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n14365) );
  NAND2_X1 U14021 ( .A1(n14365), .A2(n14570), .ZN(n11444) );
  NAND2_X1 U14022 ( .A1(n14160), .A2(n14569), .ZN(n11443) );
  NAND2_X1 U14023 ( .A1(n11444), .A2(n11443), .ZN(n14151) );
  AOI21_X1 U14024 ( .B1(n11445), .B2(n6917), .A(n14151), .ZN(n11466) );
  OAI21_X1 U14025 ( .B1(n14154), .B2(n14556), .A(n11466), .ZN(n11450) );
  AOI21_X1 U14026 ( .B1(n14156), .B2(n11446), .A(n15091), .ZN(n11447) );
  NAND2_X1 U14027 ( .A1(n11447), .A2(n11535), .ZN(n11465) );
  NOR2_X1 U14028 ( .A1(n11465), .A2(n14543), .ZN(n11449) );
  INV_X1 U14029 ( .A(n14156), .ZN(n11467) );
  OAI22_X1 U14030 ( .A1(n11467), .A2(n15088), .B1(n15065), .B2(n14547), .ZN(
        n11448) );
  AOI211_X1 U14031 ( .C1(n11450), .C2(n14547), .A(n11449), .B(n11448), .ZN(
        n11451) );
  OAI21_X1 U14032 ( .B1(n14601), .B2(n11452), .A(n11451), .ZN(P1_U3278) );
  INV_X1 U14033 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11459) );
  AOI21_X1 U14034 ( .B1(n15434), .B2(n11454), .A(n11453), .ZN(n11455) );
  OAI211_X1 U14035 ( .C1(n15407), .C2(n11457), .A(n11456), .B(n11455), .ZN(
        n11460) );
  NAND2_X1 U14036 ( .A1(n11460), .A2(n15444), .ZN(n11458) );
  OAI21_X1 U14037 ( .B1(n15444), .B2(n11459), .A(n11458), .ZN(P2_U3469) );
  NAND2_X1 U14038 ( .A1(n11460), .A2(n15457), .ZN(n11461) );
  OAI21_X1 U14039 ( .B1(n15457), .B2(n11023), .A(n11461), .ZN(P2_U3512) );
  NAND2_X1 U14040 ( .A1(n11462), .A2(n14835), .ZN(n11464) );
  AOI22_X1 U14041 ( .A1(n8194), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_24_), .B2(
        n14834), .ZN(n11463) );
  NAND2_X1 U14042 ( .A1(n11464), .A2(n11463), .ZN(P3_U3271) );
  OAI211_X1 U14043 ( .C1(n11467), .C2(n15194), .A(n11466), .B(n11465), .ZN(
        n11468) );
  AOI21_X1 U14044 ( .B1(n11469), .B2(n15198), .A(n11468), .ZN(n11472) );
  NAND2_X1 U14045 ( .A1(n15210), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11470) );
  OAI21_X1 U14046 ( .B1(n11472), .B2(n15210), .A(n11470), .ZN(P1_U3543) );
  NAND2_X1 U14047 ( .A1(n15199), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11471) );
  OAI21_X1 U14048 ( .B1(n11472), .B2(n15199), .A(n11471), .ZN(P1_U3504) );
  INV_X1 U14049 ( .A(n11473), .ZN(n11475) );
  NOR2_X1 U14050 ( .A1(n11475), .A2(n11474), .ZN(n11476) );
  XNOR2_X1 U14051 ( .A(n11476), .B(n12593), .ZN(n11484) );
  OAI21_X1 U14052 ( .B1(n11478), .B2(n12571), .A(n11477), .ZN(n11481) );
  NOR2_X1 U14053 ( .A1(n12549), .A2(n11479), .ZN(n11480) );
  AOI211_X1 U14054 ( .C1(n15463), .C2(n11482), .A(n11481), .B(n11480), .ZN(
        n11483) );
  OAI21_X1 U14055 ( .B1(n11484), .B2(n12552), .A(n11483), .ZN(P3_U3176) );
  XNOR2_X1 U14056 ( .A(n13792), .B(n13336), .ZN(n11485) );
  NAND2_X1 U14057 ( .A1(n13506), .A2(n13318), .ZN(n11486) );
  NAND2_X1 U14058 ( .A1(n11485), .A2(n11486), .ZN(n11590) );
  INV_X1 U14059 ( .A(n11485), .ZN(n11488) );
  INV_X1 U14060 ( .A(n11486), .ZN(n11487) );
  NAND2_X1 U14061 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  NAND2_X1 U14062 ( .A1(n11590), .A2(n11489), .ZN(n11497) );
  INV_X1 U14063 ( .A(n11492), .ZN(n11493) );
  NAND2_X1 U14064 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  AOI21_X1 U14065 ( .B1(n11497), .B2(n11496), .A(n6716), .ZN(n11503) );
  NAND2_X1 U14066 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15288)
         );
  OAI21_X1 U14067 ( .B1(n11498), .B2(n13421), .A(n15288), .ZN(n11499) );
  AOI21_X1 U14068 ( .B1(n13452), .B2(n13797), .A(n11499), .ZN(n11500) );
  OAI21_X1 U14069 ( .B1(n13789), .B2(n15226), .A(n11500), .ZN(n11501) );
  AOI21_X1 U14070 ( .B1(n13792), .B2(n15223), .A(n11501), .ZN(n11502) );
  OAI21_X1 U14071 ( .B1(n11503), .B2(n13480), .A(n11502), .ZN(P2_U3187) );
  NAND2_X1 U14072 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  XNOR2_X1 U14073 ( .A(n11507), .B(n11506), .ZN(n11514) );
  NOR2_X1 U14074 ( .A1(n12576), .A2(n11557), .ZN(n11511) );
  INV_X1 U14075 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11508) );
  OAI22_X1 U14076 ( .A1(n11509), .A2(n12571), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11508), .ZN(n11510) );
  AOI211_X1 U14077 ( .C1(n12573), .C2(n11512), .A(n11511), .B(n11510), .ZN(
        n11513) );
  OAI21_X1 U14078 ( .B1(n11514), .B2(n12552), .A(n11513), .ZN(P3_U3164) );
  OR2_X1 U14079 ( .A1(n11515), .A2(n11748), .ZN(n11561) );
  NAND2_X1 U14080 ( .A1(n11515), .A2(n11748), .ZN(n11516) );
  NAND3_X1 U14081 ( .A1(n11561), .A2(n12861), .A3(n11516), .ZN(n11520) );
  OR2_X1 U14082 ( .A1(n11517), .A2(n15561), .ZN(n11519) );
  OR2_X1 U14083 ( .A1(n12566), .A2(n15563), .ZN(n11518) );
  AND2_X1 U14084 ( .A1(n11519), .A2(n11518), .ZN(n11903) );
  AND2_X1 U14085 ( .A1(n11520), .A2(n11903), .ZN(n13209) );
  OR2_X1 U14086 ( .A1(n11521), .A2(n11748), .ZN(n11522) );
  NAND2_X1 U14087 ( .A1(n11568), .A2(n11522), .ZN(n13207) );
  INV_X1 U14088 ( .A(n11908), .ZN(n13264) );
  NOR2_X1 U14089 ( .A1(n13264), .A2(n12870), .ZN(n11524) );
  OAI22_X1 U14090 ( .A1(n15566), .A2(n7945), .B1(n11906), .B2(n15553), .ZN(
        n11523) );
  AOI211_X1 U14091 ( .C1(n13207), .C2(n12872), .A(n11524), .B(n11523), .ZN(
        n11525) );
  OAI21_X1 U14092 ( .B1(n13209), .B2(n14943), .A(n11525), .ZN(P3_U3220) );
  NAND2_X1 U14093 ( .A1(n11526), .A2(n12234), .ZN(n11528) );
  AOI22_X1 U14094 ( .A1(n12223), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12066), 
        .B2(n14279), .ZN(n11527) );
  INV_X1 U14095 ( .A(n14365), .ZN(n14592) );
  XNOR2_X1 U14096 ( .A(n14686), .B(n14592), .ZN(n14346) );
  XOR2_X1 U14097 ( .A(n14346), .B(n14347), .Z(n14692) );
  OR2_X1 U14098 ( .A1(n14156), .A2(n14159), .ZN(n11531) );
  NAND2_X1 U14099 ( .A1(n11534), .A2(n14346), .ZN(n14367) );
  OAI21_X1 U14100 ( .B1(n11534), .B2(n14346), .A(n14367), .ZN(n14690) );
  AOI21_X1 U14101 ( .B1(n14686), .B2(n11535), .A(n15091), .ZN(n11536) );
  NAND2_X1 U14102 ( .A1(n11536), .A2(n14584), .ZN(n14688) );
  NAND2_X1 U14103 ( .A1(n11538), .A2(n11537), .ZN(n11539) );
  NAND2_X1 U14104 ( .A1(n12069), .A2(n11539), .ZN(n14585) );
  INV_X1 U14105 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n11540) );
  OR2_X1 U14106 ( .A1(n12149), .A2(n11540), .ZN(n11543) );
  INV_X1 U14107 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11541) );
  OR2_X1 U14108 ( .A1(n12219), .A2(n11541), .ZN(n11542) );
  AND2_X1 U14109 ( .A1(n11543), .A2(n11542), .ZN(n11545) );
  INV_X1 U14110 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14305) );
  OR2_X1 U14111 ( .A1(n11348), .A2(n14305), .ZN(n11544) );
  AOI22_X1 U14112 ( .A1(n14568), .A2(n14570), .B1(n14569), .B2(n14159), .ZN(
        n14687) );
  NAND2_X1 U14113 ( .A1(n15086), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14114 ( .A1(n15085), .A2(n14079), .ZN(n11546) );
  OAI211_X1 U14115 ( .C1(n15098), .C2(n14687), .A(n11547), .B(n11546), .ZN(
        n11548) );
  AOI21_X1 U14116 ( .B1(n14686), .B2(n14558), .A(n11548), .ZN(n11549) );
  OAI21_X1 U14117 ( .B1(n14688), .B2(n14543), .A(n11549), .ZN(n11550) );
  AOI21_X1 U14118 ( .B1(n14690), .B2(n14562), .A(n11550), .ZN(n11551) );
  OAI21_X1 U14119 ( .B1(n14564), .B2(n14692), .A(n11551), .ZN(P1_U3277) );
  AOI21_X1 U14120 ( .B1(n15600), .B2(n11553), .A(n11552), .ZN(n11555) );
  MUX2_X1 U14121 ( .A(n11061), .B(n11555), .S(n15631), .Z(n11554) );
  OAI21_X1 U14122 ( .B1(n11557), .B2(n13211), .A(n11554), .ZN(P3_U3471) );
  MUX2_X1 U14123 ( .A(n7924), .B(n11555), .S(n15613), .Z(n11556) );
  OAI21_X1 U14124 ( .B1(n11557), .B2(n13263), .A(n11556), .ZN(P3_U3426) );
  AND2_X1 U14125 ( .A1(n11559), .A2(n11558), .ZN(n12859) );
  NAND3_X1 U14126 ( .A1(n11561), .A2(n11756), .A3(n11560), .ZN(n11562) );
  NAND3_X1 U14127 ( .A1(n12859), .A2(n12861), .A3(n11562), .ZN(n11566) );
  OR2_X1 U14128 ( .A1(n11899), .A2(n15561), .ZN(n11565) );
  OR2_X1 U14129 ( .A1(n11563), .A2(n15563), .ZN(n11564) );
  AND2_X1 U14130 ( .A1(n11565), .A2(n11564), .ZN(n12461) );
  AND2_X1 U14131 ( .A1(n11566), .A2(n12461), .ZN(n13205) );
  INV_X1 U14132 ( .A(n11756), .ZN(n11567) );
  NAND3_X1 U14133 ( .A1(n11568), .A2(n11567), .A3(n11752), .ZN(n11569) );
  NAND2_X1 U14134 ( .A1(n11570), .A2(n11569), .ZN(n13203) );
  AOI22_X1 U14135 ( .A1(n14943), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14938), 
        .B2(n12463), .ZN(n11571) );
  OAI21_X1 U14136 ( .B1(n13260), .B2(n12870), .A(n11571), .ZN(n11572) );
  AOI21_X1 U14137 ( .B1(n13203), .B2(n12872), .A(n11572), .ZN(n11573) );
  OAI21_X1 U14138 ( .B1(n13205), .B2(n14943), .A(n11573), .ZN(P3_U3219) );
  AOI22_X1 U14139 ( .A1(n15005), .A2(n12411), .B1(n12363), .B2(n14163), .ZN(
        n11574) );
  XNOR2_X1 U14140 ( .A(n11574), .B(n12413), .ZN(n11597) );
  AOI22_X1 U14141 ( .A1(n15005), .A2(n12363), .B1(n12412), .B2(n14163), .ZN(
        n11598) );
  XNOR2_X1 U14142 ( .A(n11597), .B(n11598), .ZN(n11583) );
  INV_X1 U14143 ( .A(n11575), .ZN(n11577) );
  INV_X1 U14144 ( .A(n11582), .ZN(n11580) );
  INV_X1 U14145 ( .A(n11583), .ZN(n11579) );
  INV_X1 U14146 ( .A(n11600), .ZN(n11581) );
  AOI21_X1 U14147 ( .B1(n11583), .B2(n11582), .A(n11581), .ZN(n11589) );
  NAND2_X1 U14148 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15043)
         );
  OAI21_X1 U14149 ( .B1(n14983), .B2(n11601), .A(n15043), .ZN(n11584) );
  AOI21_X1 U14150 ( .B1(n14140), .B2(n14164), .A(n11584), .ZN(n11585) );
  OAI21_X1 U14151 ( .B1(n11586), .B2(n14998), .A(n11585), .ZN(n11587) );
  AOI21_X1 U14152 ( .B1(n14995), .B2(n15005), .A(n11587), .ZN(n11588) );
  OAI21_X1 U14153 ( .B1(n11589), .B2(n14989), .A(n11588), .ZN(P1_U3236) );
  INV_X1 U14154 ( .A(n13981), .ZN(n14958) );
  INV_X1 U14155 ( .A(n13483), .ZN(n13462) );
  NAND2_X1 U14156 ( .A1(n13462), .A2(n13784), .ZN(n11592) );
  AND2_X1 U14157 ( .A1(n13784), .A2(n13318), .ZN(n13288) );
  OR2_X1 U14158 ( .A1(n13288), .A2(n13480), .ZN(n11591) );
  XNOR2_X1 U14159 ( .A(n13981), .B(n13384), .ZN(n13290) );
  MUX2_X1 U14160 ( .A(n11592), .B(n11591), .S(n13289), .Z(n11596) );
  INV_X1 U14161 ( .A(n11593), .ZN(n14955) );
  INV_X1 U14162 ( .A(n15226), .ZN(n13488) );
  AOI22_X1 U14163 ( .A1(n13854), .A2(n13506), .B1(n13505), .B2(n13851), .ZN(
        n13975) );
  OAI22_X1 U14164 ( .A1(n13975), .A2(n15216), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13166), .ZN(n11594) );
  AOI21_X1 U14165 ( .B1(n14955), .B2(n13488), .A(n11594), .ZN(n11595) );
  OAI211_X1 U14166 ( .C1(n14958), .C2(n13447), .A(n11596), .B(n11595), .ZN(
        P2_U3213) );
  NOR2_X1 U14167 ( .A1(n12369), .A2(n11601), .ZN(n11602) );
  AOI21_X1 U14168 ( .B1(n12002), .B2(n12329), .A(n11602), .ZN(n12307) );
  NAND2_X1 U14169 ( .A1(n12002), .A2(n12411), .ZN(n11604) );
  NAND2_X1 U14170 ( .A1(n12363), .A2(n14162), .ZN(n11603) );
  NAND2_X1 U14171 ( .A1(n11604), .A2(n11603), .ZN(n11605) );
  XNOR2_X1 U14172 ( .A(n11605), .B(n12327), .ZN(n12306) );
  XOR2_X1 U14173 ( .A(n12307), .B(n12306), .Z(n11607) );
  AOI21_X1 U14174 ( .B1(n11606), .B2(n11607), .A(n14989), .ZN(n11609) );
  NAND2_X1 U14175 ( .A1(n11609), .A2(n12309), .ZN(n11615) );
  NOR2_X1 U14176 ( .A1(n14998), .A2(n11610), .ZN(n11613) );
  OAI21_X1 U14177 ( .B1(n14983), .B2(n14981), .A(n11611), .ZN(n11612) );
  AOI211_X1 U14178 ( .C1(n14140), .C2(n14163), .A(n11613), .B(n11612), .ZN(
        n11614) );
  OAI211_X1 U14179 ( .C1(n14852), .C2(n14128), .A(n11615), .B(n11614), .ZN(
        P1_U3224) );
  OAI222_X1 U14180 ( .A1(n12426), .A2(n12124), .B1(P1_U3086), .B2(n11617), 
        .C1(n11616), .C2(n12296), .ZN(P1_U3331) );
  OAI222_X1 U14181 ( .A1(P2_U3088), .A2(n11619), .B1(n14022), .B2(n12124), 
        .C1(n11618), .C2(n14024), .ZN(P2_U3303) );
  NOR2_X1 U14182 ( .A1(n11645), .A2(n12448), .ZN(n11828) );
  OAI22_X1 U14183 ( .A1(n12438), .A2(n13176), .B1(P2_DATAO_REG_30__SCAN_IN), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14184 ( .A1(n9294), .A2(SI_30_), .ZN(n11623) );
  INV_X1 U14185 ( .A(n14951), .ZN(n11644) );
  AOI22_X1 U14186 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n14004), .B2(n11629), .ZN(n11630) );
  INV_X1 U14187 ( .A(n11630), .ZN(n11631) );
  NAND2_X1 U14188 ( .A1(n13269), .A2(n11633), .ZN(n11635) );
  NAND2_X1 U14189 ( .A1(n9294), .A2(SI_31_), .ZN(n11634) );
  NAND2_X1 U14190 ( .A1(n11636), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11642) );
  INV_X1 U14191 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n14940) );
  OR2_X1 U14192 ( .A1(n11637), .A2(n14940), .ZN(n11641) );
  INV_X1 U14193 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11638) );
  OR2_X1 U14194 ( .A1(n6570), .A2(n11638), .ZN(n11640) );
  NAND4_X1 U14195 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n14936) );
  INV_X1 U14196 ( .A(n14936), .ZN(n11648) );
  OAI22_X1 U14197 ( .A1(n11644), .A2(n12577), .B1(n14947), .B2(n11648), .ZN(
        n11831) );
  AND2_X1 U14198 ( .A1(n11645), .A2(n12448), .ZN(n11826) );
  AOI21_X1 U14199 ( .B1(n14951), .B2(n11648), .A(n11826), .ZN(n11646) );
  INV_X1 U14200 ( .A(n14947), .ZN(n11649) );
  NAND2_X1 U14201 ( .A1(n14947), .A2(n11648), .ZN(n11830) );
  INV_X1 U14202 ( .A(n12441), .ZN(n11824) );
  NAND2_X1 U14203 ( .A1(n11679), .A2(n11678), .ZN(n11680) );
  INV_X1 U14204 ( .A(n11748), .ZN(n11669) );
  NAND4_X1 U14205 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11661) );
  NOR2_X1 U14206 ( .A1(n11661), .A2(n11660), .ZN(n11666) );
  NAND3_X1 U14207 ( .A1(n11708), .A2(n11662), .A3(n15555), .ZN(n11663) );
  NOR2_X1 U14208 ( .A1(n11663), .A2(n11718), .ZN(n11665) );
  NAND4_X1 U14209 ( .A1(n11666), .A2(n11665), .A3(n11725), .A4(n11664), .ZN(
        n11667) );
  NOR4_X1 U14210 ( .A1(n11669), .A2(n11742), .A3(n11668), .A4(n11667), .ZN(
        n11670) );
  NAND4_X1 U14211 ( .A1(n12842), .A2(n12866), .A3(n11670), .A4(n11756), .ZN(
        n11671) );
  NOR4_X1 U14212 ( .A1(n12804), .A2(n11777), .A3(n12828), .A4(n11671), .ZN(
        n11672) );
  NAND3_X1 U14213 ( .A1(n12759), .A2(n12788), .A3(n11672), .ZN(n11673) );
  NOR4_X1 U14214 ( .A1(n12779), .A2(n12719), .A3(n11680), .A4(n11673), .ZN(
        n11674) );
  NAND4_X1 U14215 ( .A1(n11815), .A2(n12708), .A3(n11674), .A4(n12741), .ZN(
        n11675) );
  NOR2_X1 U14216 ( .A1(n11824), .A2(n11675), .ZN(n11676) );
  MUX2_X1 U14217 ( .A(n11679), .B(n11678), .S(n11795), .Z(n11799) );
  INV_X1 U14218 ( .A(n12779), .ZN(n11794) );
  NAND2_X1 U14219 ( .A1(n11685), .A2(n11682), .ZN(n11681) );
  AOI21_X1 U14220 ( .B1(n11681), .B2(n11688), .A(n11795), .ZN(n11684) );
  NOR2_X1 U14221 ( .A1(n9321), .A2(n11682), .ZN(n11683) );
  NAND2_X1 U14222 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U14223 ( .A1(n11687), .A2(n11795), .ZN(n11690) );
  OAI21_X1 U14224 ( .B1(n11688), .B2(n8226), .A(n15555), .ZN(n11689) );
  AOI21_X1 U14225 ( .B1(n11691), .B2(n11690), .A(n11689), .ZN(n11695) );
  AOI21_X1 U14226 ( .B1(n11693), .B2(n11692), .A(n11795), .ZN(n11694) );
  NAND2_X1 U14227 ( .A1(n11699), .A2(n11701), .ZN(n11696) );
  AOI22_X1 U14228 ( .A1(n11696), .A2(n11702), .B1(n12600), .B2(n15581), .ZN(
        n11697) );
  NAND2_X1 U14229 ( .A1(n11707), .A2(n11706), .ZN(n11713) );
  NAND3_X1 U14230 ( .A1(n11713), .A2(n11795), .A3(n11710), .ZN(n11709) );
  OAI211_X1 U14231 ( .C1(n11795), .C2(n11710), .A(n11709), .B(n11708), .ZN(
        n11711) );
  INV_X1 U14232 ( .A(n11711), .ZN(n11712) );
  INV_X1 U14233 ( .A(n11714), .ZN(n11717) );
  INV_X1 U14234 ( .A(n11715), .ZN(n11716) );
  MUX2_X1 U14235 ( .A(n11717), .B(n11716), .S(n11795), .Z(n11719) );
  NOR2_X1 U14236 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  NAND2_X1 U14237 ( .A1(n11721), .A2(n8226), .ZN(n11723) );
  OR2_X1 U14238 ( .A1(n11721), .A2(n8226), .ZN(n11722) );
  MUX2_X1 U14239 ( .A(n11723), .B(n11722), .S(n12596), .Z(n11724) );
  NAND3_X1 U14240 ( .A1(n11726), .A2(n11725), .A3(n11724), .ZN(n11739) );
  INV_X1 U14241 ( .A(n11727), .ZN(n11730) );
  INV_X1 U14242 ( .A(n11728), .ZN(n11729) );
  MUX2_X1 U14243 ( .A(n11730), .B(n11729), .S(n11795), .Z(n11732) );
  NOR2_X1 U14244 ( .A1(n11732), .A2(n11731), .ZN(n11738) );
  INV_X1 U14245 ( .A(n11733), .ZN(n11736) );
  INV_X1 U14246 ( .A(n11734), .ZN(n11735) );
  MUX2_X1 U14247 ( .A(n11736), .B(n11735), .S(n8226), .Z(n11737) );
  AOI21_X1 U14248 ( .B1(n11739), .B2(n11738), .A(n11737), .ZN(n11743) );
  AND2_X1 U14249 ( .A1(n11749), .A2(n11740), .ZN(n11741) );
  AOI21_X1 U14250 ( .B1(n11746), .B2(n11744), .A(n8226), .ZN(n11745) );
  AOI21_X1 U14251 ( .B1(n11747), .B2(n11746), .A(n11745), .ZN(n11751) );
  OAI21_X1 U14252 ( .B1(n8226), .B2(n11749), .A(n11748), .ZN(n11750) );
  AND2_X1 U14253 ( .A1(n11756), .A2(n11752), .ZN(n11753) );
  AOI22_X1 U14254 ( .A1(n11758), .A2(n11753), .B1(n12590), .B2(n13260), .ZN(
        n11754) );
  NAND4_X1 U14255 ( .A1(n11758), .A2(n11795), .A3(n11757), .A4(n11756), .ZN(
        n11759) );
  NAND2_X1 U14256 ( .A1(n11760), .A2(n11759), .ZN(n11766) );
  NAND2_X1 U14257 ( .A1(n11767), .A2(n11761), .ZN(n11764) );
  NAND2_X1 U14258 ( .A1(n11768), .A2(n11762), .ZN(n11763) );
  MUX2_X1 U14259 ( .A(n11764), .B(n11763), .S(n11795), .Z(n11765) );
  AOI21_X1 U14260 ( .B1(n11766), .B2(n12866), .A(n11765), .ZN(n11772) );
  INV_X1 U14261 ( .A(n11767), .ZN(n11770) );
  INV_X1 U14262 ( .A(n11768), .ZN(n11769) );
  MUX2_X1 U14263 ( .A(n11770), .B(n11769), .S(n8226), .Z(n11771) );
  OR2_X1 U14264 ( .A1(n11772), .A2(n11771), .ZN(n11783) );
  NOR2_X1 U14265 ( .A1(n11777), .A2(n12828), .ZN(n11782) );
  NAND2_X1 U14266 ( .A1(n11776), .A2(n11773), .ZN(n11774) );
  NAND3_X1 U14267 ( .A1(n11785), .A2(n11775), .A3(n11774), .ZN(n11780) );
  OAI211_X1 U14268 ( .C1(n11778), .C2(n11777), .A(n11784), .B(n11776), .ZN(
        n11779) );
  MUX2_X1 U14269 ( .A(n11780), .B(n11779), .S(n8226), .Z(n11781) );
  AOI21_X1 U14270 ( .B1(n11783), .B2(n11782), .A(n11781), .ZN(n11789) );
  INV_X1 U14271 ( .A(n11784), .ZN(n11787) );
  INV_X1 U14272 ( .A(n11785), .ZN(n11786) );
  MUX2_X1 U14273 ( .A(n11787), .B(n11786), .S(n8226), .Z(n11788) );
  MUX2_X1 U14274 ( .A(n11791), .B(n11790), .S(n8226), .Z(n11792) );
  NAND2_X1 U14275 ( .A1(n12586), .A2(n11795), .ZN(n11797) );
  OR2_X1 U14276 ( .A1(n12586), .A2(n11795), .ZN(n11796) );
  MUX2_X1 U14277 ( .A(n11797), .B(n11796), .S(n12781), .Z(n11798) );
  NOR2_X1 U14278 ( .A1(n12584), .A2(n8226), .ZN(n11800) );
  NAND2_X1 U14279 ( .A1(n12741), .A2(n11802), .ZN(n11805) );
  XNOR2_X1 U14280 ( .A(n11803), .B(n8226), .ZN(n11804) );
  NAND2_X1 U14281 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  OAI21_X1 U14282 ( .B1(n12735), .B2(n11807), .A(n11806), .ZN(n11811) );
  MUX2_X1 U14283 ( .A(n11809), .B(n11808), .S(n8226), .Z(n11810) );
  MUX2_X1 U14284 ( .A(n11813), .B(n11812), .S(n8226), .Z(n11814) );
  NAND2_X1 U14285 ( .A1(n11816), .A2(n11815), .ZN(n11823) );
  OAI21_X1 U14286 ( .B1(n11817), .B2(n12701), .A(n11823), .ZN(n11822) );
  INV_X1 U14287 ( .A(n11818), .ZN(n11821) );
  NOR2_X1 U14288 ( .A1(n11819), .A2(n8226), .ZN(n11820) );
  NOR3_X1 U14289 ( .A1(n11824), .A2(n11823), .A3(n8226), .ZN(n11825) );
  NOR3_X1 U14290 ( .A1(n11827), .A2(n11826), .A3(n11825), .ZN(n11829) );
  NAND4_X1 U14291 ( .A1(n12849), .A2(n11839), .A3(n7131), .A4(n11838), .ZN(
        n11840) );
  OAI211_X1 U14292 ( .C1(n11841), .C2(n11843), .A(n11840), .B(P3_B_REG_SCAN_IN), .ZN(n11842) );
  OAI21_X1 U14293 ( .B1(n11844), .B2(n11843), .A(n11842), .ZN(P3_U3296) );
  XNOR2_X1 U14294 ( .A(n11845), .B(n11846), .ZN(n11852) );
  OR2_X1 U14295 ( .A1(n12509), .A2(n15561), .ZN(n11848) );
  NAND2_X1 U14296 ( .A1(n12588), .A2(n8165), .ZN(n11847) );
  AND2_X1 U14297 ( .A1(n11848), .A2(n11847), .ZN(n12818) );
  NAND2_X1 U14298 ( .A1(n12573), .A2(n12821), .ZN(n11849) );
  NAND2_X1 U14299 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12633)
         );
  OAI211_X1 U14300 ( .C1(n12818), .C2(n12571), .A(n11849), .B(n12633), .ZN(
        n11850) );
  AOI21_X1 U14301 ( .B1(n12910), .B2(n15463), .A(n11850), .ZN(n11851) );
  OAI21_X1 U14302 ( .B1(n11852), .B2(n12552), .A(n11851), .ZN(P3_U3178) );
  AOI21_X1 U14303 ( .B1(n11854), .B2(n13476), .A(n11853), .ZN(n11855) );
  OAI21_X1 U14304 ( .B1(n15226), .B2(n11856), .A(n11855), .ZN(n11863) );
  INV_X1 U14305 ( .A(n11857), .ZN(n11861) );
  AOI22_X1 U14306 ( .A1(n13462), .A2(n13512), .B1(n13492), .B2(n11858), .ZN(
        n11860) );
  NOR3_X1 U14307 ( .A1(n11861), .A2(n11860), .A3(n11859), .ZN(n11862) );
  AOI211_X1 U14308 ( .C1(n15390), .C2(n15223), .A(n11863), .B(n11862), .ZN(
        n11864) );
  OAI21_X1 U14309 ( .B1(n11865), .B2(n13480), .A(n11864), .ZN(P2_U3199) );
  INV_X1 U14310 ( .A(n14009), .ZN(n11867) );
  OAI222_X1 U14311 ( .A1(n12296), .A2(n11868), .B1(n12426), .B2(n11867), .C1(
        n11866), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U14312 ( .A(n12195), .ZN(n14715) );
  OAI222_X1 U14313 ( .A1(n14024), .A2(n11870), .B1(n14022), .B2(n14715), .C1(
        n11869), .C2(P2_U3088), .ZN(P2_U3298) );
  INV_X1 U14314 ( .A(n12224), .ZN(n12439) );
  OAI222_X1 U14315 ( .A1(n12296), .A2(n13176), .B1(n11871), .B2(P1_U3086), 
        .C1(n12426), .C2(n12439), .ZN(P1_U3325) );
  OAI21_X1 U14316 ( .B1(n11873), .B2(n13409), .A(n11872), .ZN(n11874) );
  AOI21_X1 U14317 ( .B1(n13451), .B2(n13852), .A(n11874), .ZN(n11875) );
  OAI21_X1 U14318 ( .B1(n13860), .B2(n15226), .A(n11875), .ZN(n11881) );
  INV_X1 U14319 ( .A(n11897), .ZN(n11879) );
  AOI22_X1 U14320 ( .A1(n11876), .A2(n13492), .B1(n13462), .B2(n13853), .ZN(
        n11878) );
  NOR3_X1 U14321 ( .A1(n11879), .A2(n11878), .A3(n11877), .ZN(n11880) );
  AOI211_X1 U14322 ( .C1(n13865), .C2(n15223), .A(n11881), .B(n11880), .ZN(
        n11882) );
  OAI21_X1 U14323 ( .B1(n11883), .B2(n13480), .A(n11882), .ZN(P2_U3203) );
  INV_X1 U14324 ( .A(n11884), .ZN(n11885) );
  AOI21_X1 U14325 ( .B1(n13452), .B2(n13509), .A(n11885), .ZN(n11887) );
  NAND2_X1 U14326 ( .A1(n13451), .A2(n13508), .ZN(n11886) );
  OAI211_X1 U14327 ( .C1(n15226), .C2(n13881), .A(n11887), .B(n11886), .ZN(
        n11895) );
  INV_X1 U14328 ( .A(n11888), .ZN(n11891) );
  NOR3_X1 U14329 ( .A1(n11889), .A2(n13875), .A3(n13483), .ZN(n11890) );
  AOI21_X1 U14330 ( .B1(n11891), .B2(n13492), .A(n11890), .ZN(n11893) );
  NOR2_X1 U14331 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  AOI211_X1 U14332 ( .C1(n13889), .C2(n15223), .A(n11895), .B(n11894), .ZN(
        n11896) );
  OAI21_X1 U14333 ( .B1(n11897), .B2(n13480), .A(n11896), .ZN(P2_U3193) );
  OAI222_X1 U14334 ( .A1(n12296), .A2(n7212), .B1(n12426), .B2(n11898), .C1(
        n9547), .C2(P1_U3086), .ZN(P1_U3336) );
  XNOR2_X1 U14335 ( .A(n11900), .B(n11899), .ZN(n11901) );
  XNOR2_X1 U14336 ( .A(n11902), .B(n11901), .ZN(n11910) );
  INV_X1 U14337 ( .A(n11903), .ZN(n11904) );
  INV_X1 U14338 ( .A(n12571), .ZN(n12547) );
  AOI22_X1 U14339 ( .A1(n11904), .A2(n12547), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11905) );
  OAI21_X1 U14340 ( .B1(n12549), .B2(n11906), .A(n11905), .ZN(n11907) );
  AOI21_X1 U14341 ( .B1(n11908), .B2(n15463), .A(n11907), .ZN(n11909) );
  OAI21_X1 U14342 ( .B1(n11910), .B2(n12552), .A(n11909), .ZN(P3_U3174) );
  NAND2_X1 U14343 ( .A1(n12147), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11918) );
  INV_X1 U14344 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11911) );
  OR2_X1 U14345 ( .A1(n12149), .A2(n11911), .ZN(n11917) );
  OAI21_X1 U14346 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11913), .A(n11912), 
        .ZN(n14121) );
  OR2_X1 U14347 ( .A1(n12202), .A2(n14121), .ZN(n11916) );
  INV_X1 U14348 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11914) );
  OR2_X1 U14349 ( .A1(n12219), .A2(n11914), .ZN(n11915) );
  OR2_X1 U14350 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  XNOR2_X1 U14351 ( .A(n11921), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14720) );
  INV_X1 U14352 ( .A(n14651), .ZN(n14512) );
  NAND2_X1 U14353 ( .A1(n11924), .A2(n11923), .ZN(n11926) );
  NAND2_X1 U14354 ( .A1(n11926), .A2(n11925), .ZN(n12226) );
  NAND2_X4 U14355 ( .A1(n12226), .A2(n11927), .ZN(n12241) );
  MUX2_X1 U14356 ( .A(n14525), .B(n14512), .S(n12207), .Z(n12109) );
  INV_X1 U14357 ( .A(n11934), .ZN(n11935) );
  MUX2_X1 U14358 ( .A(n11938), .B(n6575), .S(n12241), .Z(n11940) );
  NOR2_X1 U14359 ( .A1(n11938), .A2(n6575), .ZN(n11939) );
  AOI21_X1 U14360 ( .B1(n11943), .B2(n11942), .A(n11941), .ZN(n11954) );
  INV_X1 U14361 ( .A(n11946), .ZN(n11945) );
  NAND2_X1 U14362 ( .A1(n14172), .A2(n15148), .ZN(n11948) );
  INV_X1 U14363 ( .A(n11948), .ZN(n11944) );
  NAND2_X1 U14364 ( .A1(n11955), .A2(n11946), .ZN(n11947) );
  NAND2_X1 U14365 ( .A1(n11956), .A2(n11948), .ZN(n11949) );
  OAI21_X1 U14366 ( .B1(n11954), .B2(n11953), .A(n11952), .ZN(n11958) );
  MUX2_X1 U14367 ( .A(n11956), .B(n11955), .S(n12178), .Z(n11957) );
  MUX2_X1 U14368 ( .A(n11960), .B(n11959), .S(n12241), .Z(n11963) );
  MUX2_X1 U14369 ( .A(n11961), .B(n14170), .S(n12241), .Z(n11962) );
  MUX2_X1 U14370 ( .A(n14169), .B(n11964), .S(n12178), .Z(n11967) );
  MUX2_X1 U14371 ( .A(n14169), .B(n11964), .S(n12241), .Z(n11965) );
  NAND2_X1 U14372 ( .A1(n11966), .A2(n11965), .ZN(n11971) );
  INV_X1 U14373 ( .A(n11967), .ZN(n11968) );
  NAND2_X1 U14374 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  MUX2_X1 U14375 ( .A(n14168), .B(n11972), .S(n12241), .Z(n11974) );
  MUX2_X1 U14376 ( .A(n14168), .B(n11972), .S(n12178), .Z(n11973) );
  MUX2_X1 U14377 ( .A(n14167), .B(n15170), .S(n12228), .Z(n11978) );
  NAND2_X1 U14378 ( .A1(n11977), .A2(n11978), .ZN(n11976) );
  MUX2_X1 U14379 ( .A(n14167), .B(n15170), .S(n12241), .Z(n11975) );
  NAND2_X1 U14380 ( .A1(n11976), .A2(n11975), .ZN(n11982) );
  INV_X1 U14381 ( .A(n11977), .ZN(n11980) );
  INV_X1 U14382 ( .A(n11978), .ZN(n11979) );
  MUX2_X1 U14383 ( .A(n14166), .B(n11983), .S(n12207), .Z(n11985) );
  MUX2_X1 U14384 ( .A(n14166), .B(n11983), .S(n12228), .Z(n11984) );
  INV_X1 U14385 ( .A(n11985), .ZN(n11986) );
  MUX2_X1 U14386 ( .A(n14165), .B(n11987), .S(n12228), .Z(n11989) );
  MUX2_X1 U14387 ( .A(n14165), .B(n11987), .S(n12207), .Z(n11988) );
  INV_X1 U14388 ( .A(n11989), .ZN(n11990) );
  MUX2_X1 U14389 ( .A(n14164), .B(n15191), .S(n12207), .Z(n11994) );
  NAND2_X1 U14390 ( .A1(n11993), .A2(n11994), .ZN(n11992) );
  MUX2_X1 U14391 ( .A(n14164), .B(n15191), .S(n12228), .Z(n11991) );
  NAND2_X1 U14392 ( .A1(n11992), .A2(n11991), .ZN(n11998) );
  INV_X1 U14393 ( .A(n11994), .ZN(n11995) );
  NAND2_X1 U14394 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  MUX2_X1 U14395 ( .A(n14163), .B(n15005), .S(n12228), .Z(n12000) );
  MUX2_X1 U14396 ( .A(n14163), .B(n15005), .S(n12207), .Z(n11999) );
  INV_X1 U14397 ( .A(n12000), .ZN(n12001) );
  MUX2_X1 U14398 ( .A(n14162), .B(n12002), .S(n12207), .Z(n12005) );
  NAND2_X1 U14399 ( .A1(n12006), .A2(n12005), .ZN(n12004) );
  MUX2_X1 U14400 ( .A(n14162), .B(n12002), .S(n12228), .Z(n12003) );
  NAND2_X1 U14401 ( .A1(n12004), .A2(n12003), .ZN(n12010) );
  OR2_X1 U14402 ( .A1(n12006), .A2(n12005), .ZN(n12009) );
  MUX2_X1 U14403 ( .A(n14161), .B(n12311), .S(n12178), .Z(n12014) );
  NAND2_X1 U14404 ( .A1(n12311), .A2(n12241), .ZN(n12007) );
  OAI211_X1 U14405 ( .C1(n14981), .C2(n12241), .A(n12014), .B(n12007), .ZN(
        n12008) );
  NAND2_X1 U14406 ( .A1(n12032), .A2(n12011), .ZN(n12016) );
  INV_X1 U14407 ( .A(n12241), .ZN(n12228) );
  OR2_X1 U14408 ( .A1(n14161), .A2(n12241), .ZN(n12012) );
  OAI21_X1 U14409 ( .B1(n12311), .B2(n12228), .A(n12012), .ZN(n12013) );
  NOR2_X1 U14410 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  AOI22_X1 U14411 ( .A1(n12016), .A2(n12241), .B1(n12015), .B2(n12253), .ZN(
        n12020) );
  NAND2_X1 U14412 ( .A1(n12031), .A2(n12017), .ZN(n12018) );
  NAND2_X1 U14413 ( .A1(n12018), .A2(n12228), .ZN(n12019) );
  NAND3_X1 U14414 ( .A1(n12021), .A2(n12020), .A3(n12019), .ZN(n12036) );
  MUX2_X1 U14415 ( .A(n14365), .B(n14686), .S(n12207), .Z(n12045) );
  NOR2_X1 U14416 ( .A1(n14365), .A2(n12228), .ZN(n12044) );
  AOI21_X1 U14417 ( .B1(n12045), .B2(n14568), .A(n12044), .ZN(n12030) );
  NAND2_X1 U14418 ( .A1(n12022), .A2(n12234), .ZN(n12024) );
  AOI22_X1 U14419 ( .A1(n12223), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12066), 
        .B2(n14296), .ZN(n12023) );
  INV_X1 U14420 ( .A(n14682), .ZN(n14588) );
  NAND2_X1 U14421 ( .A1(n14568), .A2(n12228), .ZN(n12039) );
  OR2_X1 U14422 ( .A1(n14686), .A2(n12039), .ZN(n12026) );
  NAND2_X1 U14423 ( .A1(n12044), .A2(n14132), .ZN(n12025) );
  AND2_X1 U14424 ( .A1(n12026), .A2(n12025), .ZN(n12041) );
  NAND2_X1 U14425 ( .A1(n12045), .A2(n14132), .ZN(n12027) );
  OR2_X1 U14426 ( .A1(n14686), .A2(n12241), .ZN(n12037) );
  NAND2_X1 U14427 ( .A1(n12027), .A2(n12037), .ZN(n12028) );
  NAND2_X1 U14428 ( .A1(n12028), .A2(n14588), .ZN(n12029) );
  OAI211_X1 U14429 ( .C1(n12030), .C2(n14588), .A(n12041), .B(n12029), .ZN(
        n12034) );
  MUX2_X1 U14430 ( .A(n12032), .B(n12031), .S(n12207), .Z(n12033) );
  NAND2_X1 U14431 ( .A1(n12036), .A2(n12035), .ZN(n12051) );
  INV_X1 U14432 ( .A(n12037), .ZN(n12038) );
  NAND2_X1 U14433 ( .A1(n12045), .A2(n12038), .ZN(n12040) );
  NAND2_X1 U14434 ( .A1(n12040), .A2(n12039), .ZN(n12043) );
  INV_X1 U14435 ( .A(n12041), .ZN(n12042) );
  AOI22_X1 U14436 ( .A1(n12043), .A2(n14588), .B1(n12045), .B2(n12042), .ZN(
        n12049) );
  NAND2_X1 U14437 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  OAI21_X1 U14438 ( .B1(n12228), .B2(n14568), .A(n12046), .ZN(n12047) );
  NAND2_X1 U14439 ( .A1(n12047), .A2(n14682), .ZN(n12048) );
  NAND2_X1 U14440 ( .A1(n12051), .A2(n12050), .ZN(n12061) );
  NAND2_X1 U14441 ( .A1(n12052), .A2(n12234), .ZN(n12054) );
  AOI22_X1 U14442 ( .A1(n12223), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12066), 
        .B2(n14316), .ZN(n12053) );
  XNOR2_X1 U14443 ( .A(n12069), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U14444 ( .A1(n14577), .A2(n12092), .ZN(n12060) );
  INV_X1 U14445 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U14446 ( .A1(n12218), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U14447 ( .A1(n12199), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n12055) );
  OAI211_X1 U14448 ( .C1(n11348), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12058) );
  INV_X1 U14449 ( .A(n12058), .ZN(n12059) );
  NAND2_X1 U14450 ( .A1(n12060), .A2(n12059), .ZN(n14370) );
  NAND2_X1 U14451 ( .A1(n14677), .A2(n12241), .ZN(n12063) );
  OR2_X1 U14452 ( .A1(n14677), .A2(n12241), .ZN(n12062) );
  MUX2_X1 U14453 ( .A(n12063), .B(n12062), .S(n14370), .Z(n12064) );
  NAND2_X1 U14454 ( .A1(n12065), .A2(n12234), .ZN(n12068) );
  AOI22_X1 U14455 ( .A1(n12223), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14445), 
        .B2(n12066), .ZN(n12067) );
  INV_X1 U14456 ( .A(n12069), .ZN(n12070) );
  AOI21_X1 U14457 ( .B1(n12070), .B2(P1_REG3_REG_18__SCAN_IN), .A(
        P1_REG3_REG_19__SCAN_IN), .ZN(n12071) );
  OR2_X1 U14458 ( .A1(n12071), .A2(n12077), .ZN(n14555) );
  AOI22_X1 U14459 ( .A1(n12147), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n12218), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U14460 ( .A1(n12199), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12072) );
  OAI211_X1 U14461 ( .C1(n14555), .C2(n12202), .A(n12073), .B(n12072), .ZN(
        n14571) );
  INV_X1 U14462 ( .A(n14571), .ZN(n12074) );
  OR2_X1 U14463 ( .A1(n14670), .A2(n12074), .ZN(n12075) );
  NAND2_X1 U14464 ( .A1(n14670), .A2(n12074), .ZN(n14352) );
  AND2_X2 U14465 ( .A1(n12075), .A2(n14352), .ZN(n14553) );
  MUX2_X1 U14466 ( .A(n14352), .B(n12075), .S(n12228), .Z(n12076) );
  NOR2_X1 U14467 ( .A1(n12077), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12078) );
  OR2_X1 U14468 ( .A1(n12089), .A2(n12078), .ZN(n14100) );
  INV_X1 U14469 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U14470 ( .A1(n12199), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U14471 ( .A1(n12218), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U14472 ( .C1(n11348), .C2(n12081), .A(n12080), .B(n12079), .ZN(
        n12082) );
  INV_X1 U14473 ( .A(n12082), .ZN(n12083) );
  NAND2_X1 U14474 ( .A1(n12223), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12085) );
  MUX2_X1 U14475 ( .A(n14526), .B(n14540), .S(n12207), .Z(n12088) );
  OR2_X1 U14476 ( .A1(n12089), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12091) );
  AND2_X1 U14477 ( .A1(n12091), .A2(n12090), .ZN(n14521) );
  NAND2_X1 U14478 ( .A1(n14521), .A2(n12092), .ZN(n12098) );
  INV_X1 U14479 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U14480 ( .A1(n12199), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U14481 ( .A1(n12198), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12093) );
  OAI211_X1 U14482 ( .C1(n11348), .C2(n12095), .A(n12094), .B(n12093), .ZN(
        n12096) );
  INV_X1 U14483 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U14484 ( .A1(n12098), .A2(n12097), .ZN(n14374) );
  NAND2_X1 U14485 ( .A1(n12223), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12100) );
  MUX2_X1 U14486 ( .A(n14374), .B(n14657), .S(n12228), .Z(n12104) );
  MUX2_X1 U14487 ( .A(n14374), .B(n14657), .S(n12207), .Z(n12102) );
  INV_X1 U14488 ( .A(n12104), .ZN(n12105) );
  MUX2_X1 U14489 ( .A(n14376), .B(n14651), .S(n12228), .Z(n12106) );
  INV_X1 U14490 ( .A(n12107), .ZN(n12110) );
  NAND2_X1 U14491 ( .A1(n12111), .A2(n12234), .ZN(n12113) );
  NAND2_X1 U14492 ( .A1(n12223), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12112) );
  MUX2_X1 U14493 ( .A(n14378), .B(n14645), .S(n12228), .Z(n12115) );
  MUX2_X1 U14494 ( .A(n14378), .B(n14645), .S(n12207), .Z(n12114) );
  NAND2_X1 U14495 ( .A1(n12147), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12122) );
  INV_X1 U14496 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n12116) );
  OR2_X1 U14497 ( .A1(n12149), .A2(n12116), .ZN(n12121) );
  INV_X1 U14498 ( .A(n12117), .ZN(n12118) );
  NAND2_X1 U14499 ( .A1(n12118), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12132) );
  OAI21_X1 U14500 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n12118), .A(n12132), 
        .ZN(n14479) );
  OR2_X1 U14501 ( .A1(n12202), .A2(n14479), .ZN(n12120) );
  INV_X1 U14502 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14480) );
  OR2_X1 U14503 ( .A1(n12219), .A2(n14480), .ZN(n12119) );
  NAND4_X1 U14504 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n14488) );
  NAND2_X1 U14505 ( .A1(n12223), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12125) );
  MUX2_X1 U14506 ( .A(n12250), .B(n14488), .S(n12207), .Z(n12127) );
  NAND2_X1 U14507 ( .A1(n12147), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12138) );
  INV_X1 U14508 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n12131) );
  OR2_X1 U14509 ( .A1(n12149), .A2(n12131), .ZN(n12137) );
  INV_X1 U14510 ( .A(n12132), .ZN(n12133) );
  NAND2_X1 U14511 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n12133), .ZN(n12152) );
  OAI21_X1 U14512 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n12133), .A(n12152), 
        .ZN(n14458) );
  OR2_X1 U14513 ( .A1(n12202), .A2(n14458), .ZN(n12136) );
  INV_X1 U14514 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n12134) );
  OR2_X1 U14515 ( .A1(n12219), .A2(n12134), .ZN(n12135) );
  NAND4_X1 U14516 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n14381) );
  NAND2_X1 U14517 ( .A1(n12424), .A2(n12234), .ZN(n12140) );
  NAND2_X1 U14518 ( .A1(n12223), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12139) );
  NAND2_X2 U14519 ( .A1(n12140), .A2(n12139), .ZN(n14635) );
  MUX2_X1 U14520 ( .A(n14381), .B(n14635), .S(n12178), .Z(n12143) );
  MUX2_X1 U14521 ( .A(n14381), .B(n14635), .S(n12207), .Z(n12141) );
  NAND2_X1 U14522 ( .A1(n12295), .A2(n12234), .ZN(n12146) );
  NAND2_X1 U14523 ( .A1(n12223), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U14524 ( .A1(n12147), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12158) );
  INV_X1 U14525 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n12148) );
  OR2_X1 U14526 ( .A1(n12149), .A2(n12148), .ZN(n12157) );
  INV_X1 U14527 ( .A(n12152), .ZN(n12150) );
  NAND2_X1 U14528 ( .A1(n12150), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12169) );
  INV_X1 U14529 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U14530 ( .A1(n12152), .A2(n12151), .ZN(n12153) );
  NAND2_X1 U14531 ( .A1(n12169), .A2(n12153), .ZN(n14437) );
  OR2_X1 U14532 ( .A1(n12202), .A2(n14437), .ZN(n12156) );
  INV_X1 U14533 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n12154) );
  OR2_X1 U14534 ( .A1(n12219), .A2(n12154), .ZN(n12155) );
  NAND4_X1 U14535 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n14452) );
  NAND2_X1 U14536 ( .A1(n12160), .A2(n12159), .ZN(n12166) );
  INV_X1 U14537 ( .A(n12161), .ZN(n12164) );
  NAND2_X1 U14538 ( .A1(n12164), .A2(n12163), .ZN(n12165) );
  NAND2_X1 U14539 ( .A1(n12198), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12175) );
  INV_X1 U14540 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14428) );
  OR2_X1 U14541 ( .A1(n12219), .A2(n14428), .ZN(n12174) );
  INV_X1 U14542 ( .A(n12169), .ZN(n12167) );
  NAND2_X1 U14543 ( .A1(n12167), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12200) );
  INV_X1 U14544 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U14545 ( .A1(n12169), .A2(n12168), .ZN(n12170) );
  NAND2_X1 U14546 ( .A1(n12200), .A2(n12170), .ZN(n14427) );
  OR2_X1 U14547 ( .A1(n12202), .A2(n14427), .ZN(n12173) );
  INV_X1 U14548 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n12171) );
  OR2_X1 U14549 ( .A1(n11348), .A2(n12171), .ZN(n12172) );
  NAND4_X1 U14550 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n14404) );
  NAND2_X1 U14551 ( .A1(n14013), .A2(n12234), .ZN(n12177) );
  NAND2_X1 U14552 ( .A1(n12223), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12176) );
  MUX2_X1 U14553 ( .A(n14404), .B(n14430), .S(n12178), .Z(n12180) );
  MUX2_X1 U14554 ( .A(n14404), .B(n14430), .S(n12241), .Z(n12179) );
  INV_X1 U14555 ( .A(n12180), .ZN(n12181) );
  NAND2_X1 U14556 ( .A1(n12198), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12188) );
  INV_X1 U14557 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n12182) );
  OR2_X1 U14558 ( .A1(n11348), .A2(n12182), .ZN(n12187) );
  INV_X1 U14559 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12183) );
  XNOR2_X1 U14560 ( .A(n12200), .B(n12183), .ZN(n14410) );
  OR2_X1 U14561 ( .A1(n12202), .A2(n14410), .ZN(n12186) );
  INV_X1 U14562 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12184) );
  OR2_X1 U14563 ( .A1(n12219), .A2(n12184), .ZN(n12185) );
  NAND4_X1 U14564 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n14394) );
  NAND2_X1 U14565 ( .A1(n14009), .A2(n12234), .ZN(n12190) );
  NAND2_X1 U14566 ( .A1(n12223), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12189) );
  INV_X1 U14567 ( .A(n12193), .ZN(n12194) );
  NAND2_X1 U14568 ( .A1(n12195), .A2(n12234), .ZN(n12197) );
  NAND2_X1 U14569 ( .A1(n12223), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U14570 ( .A1(n12197), .A2(n12196), .ZN(n12279) );
  NAND2_X1 U14571 ( .A1(n12198), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U14572 ( .A1(n12199), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12205) );
  INV_X1 U14573 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n13036) );
  OR2_X1 U14574 ( .A1(n11348), .A2(n13036), .ZN(n12204) );
  INV_X1 U14575 ( .A(n12200), .ZN(n12201) );
  NAND2_X1 U14576 ( .A1(n12201), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14392) );
  OR2_X1 U14577 ( .A1(n9466), .A2(n14392), .ZN(n12203) );
  NAND4_X1 U14578 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n14403) );
  MUX2_X1 U14579 ( .A(n12279), .B(n14403), .S(n12241), .Z(n12211) );
  INV_X1 U14580 ( .A(n14403), .ZN(n12208) );
  MUX2_X1 U14581 ( .A(n12208), .B(n14611), .S(n12207), .Z(n12209) );
  NAND2_X1 U14582 ( .A1(n12213), .A2(n12212), .ZN(n12231) );
  INV_X1 U14583 ( .A(n12231), .ZN(n12233) );
  INV_X1 U14584 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12217) );
  NAND2_X1 U14585 ( .A1(n12218), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12216) );
  INV_X1 U14586 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12214) );
  OR2_X1 U14587 ( .A1(n12219), .A2(n12214), .ZN(n12215) );
  OAI211_X1 U14588 ( .C1(n11348), .C2(n12217), .A(n12216), .B(n12215), .ZN(
        n14335) );
  INV_X1 U14589 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U14590 ( .A1(n12218), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12221) );
  INV_X1 U14591 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13172) );
  OR2_X1 U14592 ( .A1(n12219), .A2(n13172), .ZN(n12220) );
  OAI211_X1 U14593 ( .C1(n11348), .C2(n13071), .A(n12221), .B(n12220), .ZN(
        n14391) );
  OAI21_X1 U14594 ( .B1(n14335), .B2(n12222), .A(n14391), .ZN(n12225) );
  AOI22_X2 U14595 ( .A1(n12224), .A2(n12234), .B1(n12223), .B2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n14606) );
  MUX2_X1 U14596 ( .A(n12225), .B(n14606), .S(n12241), .Z(n12232) );
  INV_X1 U14597 ( .A(n12232), .ZN(n12230) );
  INV_X1 U14598 ( .A(n14606), .ZN(n14331) );
  NAND2_X1 U14599 ( .A1(n14335), .A2(n12241), .ZN(n12242) );
  NAND2_X1 U14600 ( .A1(n12242), .A2(n12226), .ZN(n12227) );
  AOI22_X1 U14601 ( .A1(n14331), .A2(n12228), .B1(n14391), .B2(n12227), .ZN(
        n12229) );
  NAND2_X1 U14602 ( .A1(n14001), .A2(n12234), .ZN(n12236) );
  NAND2_X1 U14603 ( .A1(n12223), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12235) );
  OR2_X1 U14604 ( .A1(n12238), .A2(n12237), .ZN(n12240) );
  NAND2_X1 U14605 ( .A1(n12240), .A2(n12239), .ZN(n12284) );
  NOR3_X1 U14606 ( .A1(n12245), .A2(n12282), .A3(n12284), .ZN(n12289) );
  MUX2_X1 U14607 ( .A(n14335), .B(n12241), .S(n14336), .Z(n12243) );
  INV_X1 U14608 ( .A(n12244), .ZN(n12286) );
  INV_X1 U14609 ( .A(n14394), .ZN(n12246) );
  NAND2_X1 U14610 ( .A1(n14618), .A2(n12246), .ZN(n14364) );
  OR2_X1 U14611 ( .A1(n14618), .A2(n12246), .ZN(n12247) );
  INV_X1 U14612 ( .A(n14404), .ZN(n14438) );
  NAND2_X1 U14613 ( .A1(n14430), .A2(n14438), .ZN(n14363) );
  OR2_X1 U14614 ( .A1(n14430), .A2(n14438), .ZN(n12248) );
  INV_X1 U14615 ( .A(n14381), .ZN(n14469) );
  NAND2_X1 U14616 ( .A1(n14635), .A2(n14469), .ZN(n14360) );
  OR2_X1 U14617 ( .A1(n14635), .A2(n14469), .ZN(n12249) );
  INV_X1 U14618 ( .A(n14488), .ZN(n14379) );
  INV_X1 U14619 ( .A(n14378), .ZN(n14470) );
  XNOR2_X1 U14620 ( .A(n14645), .B(n14470), .ZN(n14491) );
  INV_X1 U14621 ( .A(n14374), .ZN(n14355) );
  XNOR2_X1 U14622 ( .A(n14657), .B(n14355), .ZN(n14522) );
  OR2_X1 U14623 ( .A1(n14651), .A2(n14525), .ZN(n14357) );
  NAND2_X1 U14624 ( .A1(n14651), .A2(n14525), .ZN(n12251) );
  NAND2_X1 U14625 ( .A1(n14357), .A2(n12251), .ZN(n14509) );
  INV_X1 U14626 ( .A(n14526), .ZN(n14353) );
  XNOR2_X1 U14627 ( .A(n14540), .B(n14353), .ZN(n14546) );
  INV_X1 U14628 ( .A(n14566), .ZN(n12275) );
  INV_X1 U14629 ( .A(n14553), .ZN(n14351) );
  OR2_X1 U14630 ( .A1(n14682), .A2(n14132), .ZN(n14348) );
  NAND2_X1 U14631 ( .A1(n14682), .A2(n14132), .ZN(n12252) );
  NAND2_X1 U14632 ( .A1(n14348), .A2(n12252), .ZN(n14589) );
  INV_X1 U14633 ( .A(n12253), .ZN(n12271) );
  NAND4_X1 U14634 ( .A1(n12255), .A2(n12254), .A3(n15130), .A4(n15080), .ZN(
        n12257) );
  NOR2_X1 U14635 ( .A1(n12257), .A2(n12256), .ZN(n12260) );
  NAND4_X1 U14636 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  NOR2_X1 U14637 ( .A1(n12263), .A2(n12262), .ZN(n12266) );
  NAND4_X1 U14638 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12268) );
  OR4_X1 U14639 ( .A1(n14589), .A2(n12273), .A3(n14346), .A4(n12272), .ZN(
        n12274) );
  OR4_X1 U14640 ( .A1(n14546), .A2(n12275), .A3(n14351), .A4(n12274), .ZN(
        n12276) );
  NOR2_X1 U14641 ( .A1(n14474), .A2(n12277), .ZN(n12278) );
  XOR2_X1 U14642 ( .A(n14391), .B(n14606), .Z(n12280) );
  XNOR2_X1 U14643 ( .A(n12279), .B(n14403), .ZN(n14387) );
  XNOR2_X1 U14644 ( .A(n12281), .B(n9547), .ZN(n12287) );
  NAND2_X1 U14645 ( .A1(n12282), .A2(n7655), .ZN(n12283) );
  MUX2_X1 U14646 ( .A(n12284), .B(n12283), .S(n6648), .Z(n12285) );
  OAI21_X1 U14647 ( .B1(n12287), .B2(n12286), .A(n12285), .ZN(n12288) );
  NOR2_X1 U14648 ( .A1(n14187), .A2(P1_U3086), .ZN(n14716) );
  NAND3_X1 U14649 ( .A1(n12290), .A2(n14569), .A3(n14716), .ZN(n12291) );
  OAI211_X1 U14650 ( .C1(n15133), .C2(n12293), .A(n12291), .B(P1_B_REG_SCAN_IN), .ZN(n12292) );
  OAI21_X1 U14651 ( .B1(n12294), .B2(n12293), .A(n12292), .ZN(P1_U3242) );
  INV_X1 U14652 ( .A(n12295), .ZN(n14018) );
  OAI222_X1 U14653 ( .A1(n12426), .A2(n14018), .B1(P1_U3086), .B2(n12298), 
        .C1(n12297), .C2(n12296), .ZN(P1_U3329) );
  INV_X1 U14654 ( .A(n12299), .ZN(n12301) );
  OAI222_X1 U14655 ( .A1(n12302), .A2(P3_U3151), .B1(n13282), .B2(n12301), 
        .C1(n12300), .C2(n13284), .ZN(P3_U3267) );
  AOI22_X1 U14656 ( .A1(n14682), .A2(n12411), .B1(n12363), .B2(n14568), .ZN(
        n12304) );
  XNOR2_X1 U14657 ( .A(n12304), .B(n12327), .ZN(n12338) );
  NOR2_X1 U14658 ( .A1(n12369), .A2(n14132), .ZN(n12305) );
  AOI21_X1 U14659 ( .B1(n14682), .B2(n12363), .A(n12305), .ZN(n12339) );
  INV_X1 U14660 ( .A(n12306), .ZN(n12308) );
  NOR2_X1 U14661 ( .A1(n12369), .A2(n14981), .ZN(n12310) );
  AOI21_X1 U14662 ( .B1(n12311), .B2(n12329), .A(n12310), .ZN(n12318) );
  AOI22_X1 U14663 ( .A1(n12311), .A2(n12411), .B1(n12363), .B2(n14161), .ZN(
        n12312) );
  XNOR2_X1 U14664 ( .A(n12312), .B(n12413), .ZN(n12317) );
  XOR2_X1 U14665 ( .A(n12318), .B(n12317), .Z(n14107) );
  NAND2_X1 U14666 ( .A1(n14994), .A2(n12411), .ZN(n12314) );
  NAND2_X1 U14667 ( .A1(n12329), .A2(n14160), .ZN(n12313) );
  NAND2_X1 U14668 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  XNOR2_X1 U14669 ( .A(n12315), .B(n12413), .ZN(n12322) );
  NOR2_X1 U14670 ( .A1(n12369), .A2(n14111), .ZN(n12316) );
  AOI21_X1 U14671 ( .B1(n14994), .B2(n12329), .A(n12316), .ZN(n12323) );
  XNOR2_X1 U14672 ( .A(n12322), .B(n12323), .ZN(n14985) );
  INV_X1 U14673 ( .A(n12317), .ZN(n12320) );
  INV_X1 U14674 ( .A(n12318), .ZN(n12319) );
  NAND2_X1 U14675 ( .A1(n12320), .A2(n12319), .ZN(n14986) );
  INV_X1 U14676 ( .A(n12322), .ZN(n12324) );
  NAND2_X1 U14677 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  AOI22_X1 U14678 ( .A1(n14156), .A2(n12411), .B1(n12363), .B2(n14159), .ZN(
        n12326) );
  AOI22_X1 U14679 ( .A1(n14156), .A2(n12363), .B1(n12412), .B2(n14159), .ZN(
        n14149) );
  NAND2_X1 U14680 ( .A1(n14148), .A2(n14149), .ZN(n12328) );
  NAND2_X1 U14681 ( .A1(n14686), .A2(n12411), .ZN(n12331) );
  NAND2_X1 U14682 ( .A1(n12329), .A2(n14365), .ZN(n12330) );
  NAND2_X1 U14683 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  XNOR2_X1 U14684 ( .A(n12332), .B(n12327), .ZN(n12335) );
  AOI22_X1 U14685 ( .A1(n14686), .A2(n12363), .B1(n12412), .B2(n14365), .ZN(
        n12333) );
  XNOR2_X1 U14686 ( .A(n12335), .B(n12333), .ZN(n14074) );
  NAND2_X1 U14687 ( .A1(n14075), .A2(n14074), .ZN(n12337) );
  INV_X1 U14688 ( .A(n12333), .ZN(n12334) );
  NAND2_X1 U14689 ( .A1(n12337), .A2(n12336), .ZN(n14083) );
  XOR2_X1 U14690 ( .A(n12339), .B(n12338), .Z(n14084) );
  NAND2_X1 U14691 ( .A1(n14677), .A2(n12411), .ZN(n12342) );
  NAND2_X1 U14692 ( .A1(n12363), .A2(n14370), .ZN(n12341) );
  NAND2_X1 U14693 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  XNOR2_X1 U14694 ( .A(n12343), .B(n12327), .ZN(n12344) );
  AOI22_X1 U14695 ( .A1(n14677), .A2(n12363), .B1(n12412), .B2(n14370), .ZN(
        n12345) );
  XNOR2_X1 U14696 ( .A(n12344), .B(n12345), .ZN(n14129) );
  INV_X1 U14697 ( .A(n12344), .ZN(n12346) );
  NAND2_X1 U14698 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  AND2_X1 U14699 ( .A1(n12412), .A2(n14571), .ZN(n12348) );
  AOI21_X1 U14700 ( .B1(n14670), .B2(n12363), .A(n12348), .ZN(n12352) );
  NAND2_X1 U14701 ( .A1(n14670), .A2(n12411), .ZN(n12350) );
  NAND2_X1 U14702 ( .A1(n14571), .A2(n12363), .ZN(n12349) );
  NAND2_X1 U14703 ( .A1(n12350), .A2(n12349), .ZN(n12351) );
  XNOR2_X1 U14704 ( .A(n12351), .B(n12327), .ZN(n12354) );
  XOR2_X1 U14705 ( .A(n12352), .B(n12354), .Z(n14050) );
  INV_X1 U14706 ( .A(n12352), .ZN(n12353) );
  NAND2_X1 U14707 ( .A1(n12354), .A2(n12353), .ZN(n12355) );
  AND2_X1 U14708 ( .A1(n14526), .A2(n12412), .ZN(n12356) );
  AOI21_X1 U14709 ( .B1(n14540), .B2(n12363), .A(n12356), .ZN(n12359) );
  AOI22_X1 U14710 ( .A1(n14540), .A2(n12411), .B1(n12363), .B2(n14526), .ZN(
        n12357) );
  XNOR2_X1 U14711 ( .A(n12357), .B(n12327), .ZN(n12358) );
  XOR2_X1 U14712 ( .A(n12359), .B(n12358), .Z(n14098) );
  INV_X1 U14713 ( .A(n12358), .ZN(n12361) );
  INV_X1 U14714 ( .A(n12359), .ZN(n12360) );
  NAND2_X1 U14715 ( .A1(n12361), .A2(n12360), .ZN(n12362) );
  AOI22_X1 U14716 ( .A1(n14657), .A2(n12411), .B1(n12363), .B2(n14374), .ZN(
        n12364) );
  XNOR2_X1 U14717 ( .A(n12364), .B(n12327), .ZN(n12367) );
  AOI22_X1 U14718 ( .A1(n14657), .A2(n12363), .B1(n12412), .B2(n14374), .ZN(
        n12366) );
  XNOR2_X1 U14719 ( .A(n12367), .B(n12366), .ZN(n14061) );
  INV_X1 U14720 ( .A(n14061), .ZN(n12365) );
  NAND2_X1 U14721 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  OAI22_X1 U14722 ( .A1(n14651), .A2(n12370), .B1(n14376), .B2(n12369), .ZN(
        n12374) );
  OAI22_X1 U14723 ( .A1(n14651), .A2(n12371), .B1(n14376), .B2(n12370), .ZN(
        n12372) );
  XNOR2_X1 U14724 ( .A(n12372), .B(n12327), .ZN(n12373) );
  XOR2_X1 U14725 ( .A(n12374), .B(n12373), .Z(n14118) );
  INV_X1 U14726 ( .A(n12373), .ZN(n12376) );
  INV_X1 U14727 ( .A(n12374), .ZN(n12375) );
  NAND2_X1 U14728 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  NAND2_X1 U14729 ( .A1(n14645), .A2(n12411), .ZN(n12379) );
  NAND2_X1 U14730 ( .A1(n12363), .A2(n14378), .ZN(n12378) );
  NAND2_X1 U14731 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  XNOR2_X1 U14732 ( .A(n12380), .B(n12327), .ZN(n12381) );
  AOI22_X1 U14733 ( .A1(n14645), .A2(n12363), .B1(n12412), .B2(n14378), .ZN(
        n12382) );
  XNOR2_X1 U14734 ( .A(n12381), .B(n12382), .ZN(n14036) );
  INV_X1 U14735 ( .A(n12381), .ZN(n12383) );
  NAND2_X1 U14736 ( .A1(n12250), .A2(n12411), .ZN(n12385) );
  NAND2_X1 U14737 ( .A1(n12363), .A2(n14488), .ZN(n12384) );
  NAND2_X1 U14738 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  XNOR2_X1 U14739 ( .A(n12386), .B(n12327), .ZN(n12387) );
  AOI22_X1 U14740 ( .A1(n12250), .A2(n12363), .B1(n12412), .B2(n14488), .ZN(
        n12388) );
  XNOR2_X1 U14741 ( .A(n12387), .B(n12388), .ZN(n14091) );
  NAND2_X1 U14742 ( .A1(n14090), .A2(n14091), .ZN(n12391) );
  INV_X1 U14743 ( .A(n12387), .ZN(n12389) );
  NAND2_X1 U14744 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  NAND2_X1 U14745 ( .A1(n14635), .A2(n12411), .ZN(n12393) );
  NAND2_X1 U14746 ( .A1(n12363), .A2(n14381), .ZN(n12392) );
  NAND2_X1 U14747 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  XNOR2_X1 U14748 ( .A(n12394), .B(n12327), .ZN(n12395) );
  AOI22_X1 U14749 ( .A1(n14635), .A2(n12363), .B1(n12412), .B2(n14381), .ZN(
        n12396) );
  XNOR2_X1 U14750 ( .A(n12395), .B(n12396), .ZN(n14068) );
  INV_X1 U14751 ( .A(n12395), .ZN(n12397) );
  NAND2_X1 U14752 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  NAND2_X1 U14753 ( .A1(n14630), .A2(n12411), .ZN(n12400) );
  NAND2_X1 U14754 ( .A1(n12363), .A2(n14452), .ZN(n12399) );
  NAND2_X1 U14755 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  XNOR2_X1 U14756 ( .A(n12401), .B(n12327), .ZN(n12402) );
  AOI22_X1 U14757 ( .A1(n14630), .A2(n12363), .B1(n12412), .B2(n14452), .ZN(
        n12403) );
  XNOR2_X1 U14758 ( .A(n12402), .B(n12403), .ZN(n14139) );
  INV_X1 U14759 ( .A(n12402), .ZN(n12404) );
  NAND2_X1 U14760 ( .A1(n14430), .A2(n12411), .ZN(n12406) );
  NAND2_X1 U14761 ( .A1(n12363), .A2(n14404), .ZN(n12405) );
  NAND2_X1 U14762 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  XNOR2_X1 U14763 ( .A(n12407), .B(n12413), .ZN(n12408) );
  AOI22_X1 U14764 ( .A1(n14430), .A2(n12363), .B1(n12412), .B2(n14404), .ZN(
        n12409) );
  XNOR2_X1 U14765 ( .A(n12408), .B(n12409), .ZN(n14028) );
  INV_X1 U14766 ( .A(n12408), .ZN(n12410) );
  AOI22_X1 U14767 ( .A1(n14618), .A2(n12411), .B1(n12363), .B2(n14394), .ZN(
        n12416) );
  AOI22_X1 U14768 ( .A1(n14618), .A2(n12363), .B1(n12412), .B2(n14394), .ZN(
        n12414) );
  XNOR2_X1 U14769 ( .A(n12414), .B(n12413), .ZN(n12415) );
  XOR2_X1 U14770 ( .A(n12416), .B(n12415), .Z(n12417) );
  XNOR2_X1 U14771 ( .A(n12418), .B(n12417), .ZN(n12423) );
  AOI22_X1 U14772 ( .A1(n14140), .A2(n14404), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12420) );
  NAND2_X1 U14773 ( .A1(n14141), .A2(n14403), .ZN(n12419) );
  OAI211_X1 U14774 ( .C1(n14998), .C2(n14410), .A(n12420), .B(n12419), .ZN(
        n12421) );
  AOI21_X1 U14775 ( .B1(n14618), .B2(n14995), .A(n12421), .ZN(n12422) );
  OAI21_X1 U14776 ( .B1(n12423), .B2(n14989), .A(n12422), .ZN(P1_U3220) );
  INV_X1 U14777 ( .A(n12424), .ZN(n14021) );
  OAI222_X1 U14778 ( .A1(n12296), .A2(n12987), .B1(n12426), .B2(n14021), .C1(
        n12425), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U14779 ( .A1(n7738), .A2(P3_U3151), .B1(n13282), .B2(n12428), .C1(
        n12427), .C2(n13284), .ZN(P3_U3265) );
  INV_X1 U14780 ( .A(n12429), .ZN(n12433) );
  INV_X1 U14781 ( .A(n12430), .ZN(n12431) );
  AOI22_X1 U14782 ( .A1(n12431), .A2(n15315), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15316), .ZN(n12432) );
  OAI21_X1 U14783 ( .B1(n12433), .B2(n14957), .A(n12432), .ZN(n12435) );
  XNOR2_X1 U14784 ( .A(n12441), .B(n12440), .ZN(n12450) );
  INV_X1 U14785 ( .A(n12450), .ZN(n12442) );
  NAND2_X1 U14786 ( .A1(n12442), .A2(n15469), .ZN(n12456) );
  INV_X1 U14787 ( .A(n12443), .ZN(n12444) );
  NAND4_X1 U14788 ( .A1(n12455), .A2(n15469), .A3(n12444), .A4(n12450), .ZN(
        n12454) );
  NAND2_X1 U14789 ( .A1(n12573), .A2(n12445), .ZN(n12447) );
  AOI22_X1 U14790 ( .A1(n15465), .A2(n12580), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12446) );
  OAI211_X1 U14791 ( .C1(n12448), .C2(n15467), .A(n12447), .B(n12446), .ZN(
        n12452) );
  NOR4_X1 U14792 ( .A1(n12450), .A2(n12449), .A3(n12580), .A4(n12552), .ZN(
        n12451) );
  AOI211_X1 U14793 ( .C1(n15463), .C2(n12691), .A(n12452), .B(n12451), .ZN(
        n12453) );
  OAI211_X1 U14794 ( .C1(n12456), .C2(n12455), .A(n12454), .B(n12453), .ZN(
        P3_U3160) );
  AOI21_X1 U14795 ( .B1(n12457), .B2(n12458), .A(n12552), .ZN(n12460) );
  NAND2_X1 U14796 ( .A1(n12460), .A2(n12459), .ZN(n12465) );
  NAND2_X1 U14797 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12607)
         );
  OAI21_X1 U14798 ( .B1(n12461), .B2(n12571), .A(n12607), .ZN(n12462) );
  AOI21_X1 U14799 ( .B1(n12573), .B2(n12463), .A(n12462), .ZN(n12464) );
  OAI211_X1 U14800 ( .C1(n12576), .C2(n13260), .A(n12465), .B(n12464), .ZN(
        P3_U3155) );
  INV_X1 U14801 ( .A(n12529), .ZN(n12467) );
  AOI21_X1 U14802 ( .B1(n12584), .B2(n12468), .A(n12467), .ZN(n12474) );
  OR2_X1 U14803 ( .A1(n12485), .A2(n15561), .ZN(n12470) );
  NAND2_X1 U14804 ( .A1(n12583), .A2(n8165), .ZN(n12469) );
  NAND2_X1 U14805 ( .A1(n12470), .A2(n12469), .ZN(n12751) );
  AOI22_X1 U14806 ( .A1(n12547), .A2(n12751), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12471) );
  OAI21_X1 U14807 ( .B1(n12549), .B2(n12754), .A(n12471), .ZN(n12472) );
  AOI21_X1 U14808 ( .B1(n12757), .B2(n15463), .A(n12472), .ZN(n12473) );
  OAI21_X1 U14809 ( .B1(n12474), .B2(n12552), .A(n12473), .ZN(P3_U3156) );
  XNOR2_X1 U14810 ( .A(n12475), .B(n12476), .ZN(n12480) );
  AOI22_X1 U14811 ( .A1(n12587), .A2(n8165), .B1(n12849), .B2(n12830), .ZN(
        n12806) );
  NAND2_X1 U14812 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12672)
         );
  OAI21_X1 U14813 ( .B1(n12806), .B2(n12571), .A(n12672), .ZN(n12478) );
  NOR2_X1 U14814 ( .A1(n13244), .A2(n12576), .ZN(n12477) );
  AOI211_X1 U14815 ( .C1(n12809), .C2(n12573), .A(n12478), .B(n12477), .ZN(
        n12479) );
  OAI21_X1 U14816 ( .B1(n12480), .B2(n12552), .A(n12479), .ZN(P3_U3159) );
  INV_X1 U14817 ( .A(n12481), .ZN(n12482) );
  AOI21_X1 U14818 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n12491) );
  INV_X1 U14819 ( .A(n12782), .ZN(n12488) );
  OAI22_X1 U14820 ( .A1(n12486), .A2(n15561), .B1(n12485), .B2(n15563), .ZN(
        n12776) );
  AOI22_X1 U14821 ( .A1(n12776), .A2(n12547), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12487) );
  OAI21_X1 U14822 ( .B1(n12549), .B2(n12488), .A(n12487), .ZN(n12489) );
  AOI21_X1 U14823 ( .B1(n12781), .B2(n15463), .A(n12489), .ZN(n12490) );
  OAI21_X1 U14824 ( .B1(n12491), .B2(n12552), .A(n12490), .ZN(P3_U3163) );
  OR2_X1 U14825 ( .A1(n12492), .A2(n15563), .ZN(n12494) );
  NAND2_X1 U14826 ( .A1(n12583), .A2(n12849), .ZN(n12493) );
  NAND2_X1 U14827 ( .A1(n12494), .A2(n12493), .ZN(n12721) );
  AOI22_X1 U14828 ( .A1(n12547), .A2(n12721), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12495) );
  OAI21_X1 U14829 ( .B1(n12549), .B2(n12728), .A(n12495), .ZN(n12503) );
  AND2_X1 U14830 ( .A1(n12498), .A2(n12497), .ZN(n12531) );
  NAND3_X1 U14831 ( .A1(n12531), .A2(n12500), .A3(n7236), .ZN(n12501) );
  AOI21_X1 U14832 ( .B1(n12496), .B2(n12501), .A(n12552), .ZN(n12502) );
  AOI211_X1 U14833 ( .C1(n15463), .C2(n12727), .A(n12503), .B(n12502), .ZN(
        n12504) );
  INV_X1 U14834 ( .A(n12504), .ZN(P3_U3165) );
  INV_X1 U14835 ( .A(n12505), .ZN(n13253) );
  OAI211_X1 U14836 ( .C1(n12508), .C2(n12507), .A(n12506), .B(n15469), .ZN(
        n12513) );
  OAI22_X1 U14837 ( .A1(n15467), .A2(n12509), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14900), .ZN(n12511) );
  NOR2_X1 U14838 ( .A1(n12549), .A2(n12852), .ZN(n12510) );
  AOI211_X1 U14839 ( .C1(n15465), .C2(n12848), .A(n12511), .B(n12510), .ZN(
        n12512) );
  OAI211_X1 U14840 ( .C1(n13253), .C2(n12576), .A(n12513), .B(n12512), .ZN(
        P3_U3166) );
  NOR2_X1 U14841 ( .A1(n12514), .A2(n6724), .ZN(n12515) );
  XNOR2_X1 U14842 ( .A(n12516), .B(n12515), .ZN(n12522) );
  NAND2_X1 U14843 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14917)
         );
  OAI21_X1 U14844 ( .B1(n15467), .B2(n12517), .A(n14917), .ZN(n12518) );
  AOI21_X1 U14845 ( .B1(n15465), .B2(n12831), .A(n12518), .ZN(n12519) );
  OAI21_X1 U14846 ( .B1(n12549), .B2(n12836), .A(n12519), .ZN(n12520) );
  AOI21_X1 U14847 ( .B1(n12835), .B2(n15463), .A(n12520), .ZN(n12521) );
  OAI21_X1 U14848 ( .B1(n12522), .B2(n12552), .A(n12521), .ZN(P3_U3168) );
  OR2_X1 U14849 ( .A1(n12523), .A2(n15563), .ZN(n12525) );
  NAND2_X1 U14850 ( .A1(n12584), .A2(n12849), .ZN(n12524) );
  NAND2_X1 U14851 ( .A1(n12525), .A2(n12524), .ZN(n12737) );
  AOI22_X1 U14852 ( .A1(n12547), .A2(n12737), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12526) );
  OAI21_X1 U14853 ( .B1(n12549), .B2(n12745), .A(n12526), .ZN(n12533) );
  NAND3_X1 U14854 ( .A1(n12529), .A2(n12527), .A3(n12528), .ZN(n12530) );
  AOI21_X1 U14855 ( .B1(n12531), .B2(n12530), .A(n12552), .ZN(n12532) );
  AOI211_X1 U14856 ( .C1(n15463), .C2(n12744), .A(n12533), .B(n12532), .ZN(
        n12534) );
  INV_X1 U14857 ( .A(n12534), .ZN(P3_U3169) );
  XNOR2_X1 U14858 ( .A(n12535), .B(n12536), .ZN(n12541) );
  AOI22_X1 U14859 ( .A1(n12586), .A2(n8165), .B1(n12849), .B2(n12588), .ZN(
        n12791) );
  OAI22_X1 U14860 ( .A1(n12791), .A2(n12571), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12537), .ZN(n12539) );
  NOR2_X1 U14861 ( .A1(n13240), .A2(n12576), .ZN(n12538) );
  AOI211_X1 U14862 ( .C1(n12797), .C2(n12573), .A(n12539), .B(n12538), .ZN(
        n12540) );
  OAI21_X1 U14863 ( .B1(n12541), .B2(n12552), .A(n12540), .ZN(P3_U3173) );
  INV_X1 U14864 ( .A(n12543), .ZN(n12544) );
  AOI21_X1 U14865 ( .B1(n12585), .B2(n12542), .A(n12544), .ZN(n12553) );
  INV_X1 U14866 ( .A(n12584), .ZN(n12545) );
  OAI22_X1 U14867 ( .A1(n12546), .A2(n15561), .B1(n12545), .B2(n15563), .ZN(
        n12763) );
  AOI22_X1 U14868 ( .A1(n12763), .A2(n12547), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12548) );
  OAI21_X1 U14869 ( .B1(n12549), .B2(n12769), .A(n12548), .ZN(n12550) );
  AOI21_X1 U14870 ( .B1(n12768), .B2(n15463), .A(n12550), .ZN(n12551) );
  OAI21_X1 U14871 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(P3_U3175) );
  NAND2_X1 U14872 ( .A1(n12556), .A2(n15469), .ZN(n12561) );
  INV_X1 U14873 ( .A(n12712), .ZN(n12559) );
  AOI22_X1 U14874 ( .A1(n12582), .A2(n12849), .B1(n8165), .B2(n12580), .ZN(
        n12710) );
  INV_X1 U14875 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12557) );
  OAI22_X1 U14876 ( .A1(n12710), .A2(n12571), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12557), .ZN(n12558) );
  AOI21_X1 U14877 ( .B1(n12559), .B2(n12573), .A(n12558), .ZN(n12560) );
  OAI211_X1 U14878 ( .C1(n13219), .C2(n12576), .A(n12561), .B(n12560), .ZN(
        P3_U3180) );
  INV_X1 U14879 ( .A(n12562), .ZN(n13257) );
  OAI211_X1 U14880 ( .C1(n12565), .C2(n12564), .A(n12563), .B(n15469), .ZN(
        n12575) );
  OR2_X1 U14881 ( .A1(n12566), .A2(n15561), .ZN(n12569) );
  OR2_X1 U14882 ( .A1(n12567), .A2(n15563), .ZN(n12568) );
  AND2_X1 U14883 ( .A1(n12569), .A2(n12568), .ZN(n12863) );
  OAI22_X1 U14884 ( .A1(n12863), .A2(n12571), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12570), .ZN(n12572) );
  AOI21_X1 U14885 ( .B1(n12573), .B2(n12868), .A(n12572), .ZN(n12574) );
  OAI211_X1 U14886 ( .C1(n13257), .C2(n12576), .A(n12575), .B(n12574), .ZN(
        P3_U3181) );
  MUX2_X1 U14887 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n14936), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14888 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12577), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12578), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12579), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14891 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12580), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12581), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14893 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12582), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12583), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14895 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12584), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12585), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12586), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14898 ( .A(n12587), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12589), .Z(
        P3_U3511) );
  MUX2_X1 U14899 ( .A(n12588), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12589), .Z(
        P3_U3510) );
  MUX2_X1 U14900 ( .A(n12830), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12589), .Z(
        P3_U3509) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12847), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12831), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12848), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14904 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12590), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14905 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12591), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12592), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14907 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12593), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12594), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14909 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12595), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14910 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12596), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14911 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12597), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14912 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12598), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14913 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12599), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14914 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12600), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14915 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15461), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14916 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n6822), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14917 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n6800), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14918 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n10153), .S(P3_U3897), .Z(
        P3_U3491) );
  NAND2_X1 U14919 ( .A1(n12616), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12602) );
  NOR2_X1 U14920 ( .A1(n12619), .A2(n12604), .ZN(n12605) );
  INV_X1 U14921 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15534) );
  XNOR2_X1 U14922 ( .A(n12648), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12611) );
  AOI21_X1 U14923 ( .B1(n12606), .B2(n12611), .A(n12627), .ZN(n12626) );
  INV_X1 U14924 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14807) );
  OAI21_X1 U14925 ( .B1(n15529), .B2(n14807), .A(n12607), .ZN(n12615) );
  MUX2_X1 U14926 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13279), .Z(n12610) );
  AOI21_X1 U14927 ( .B1(n12609), .B2(n12616), .A(n12608), .ZN(n15537) );
  XNOR2_X1 U14928 ( .A(n12610), .B(n12619), .ZN(n15536) );
  NAND2_X1 U14929 ( .A1(n15537), .A2(n15536), .ZN(n15535) );
  OAI21_X1 U14930 ( .B1(n12610), .B2(n15530), .A(n15535), .ZN(n12613) );
  XNOR2_X1 U14931 ( .A(n12648), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12621) );
  MUX2_X1 U14932 ( .A(n12621), .B(n12611), .S(n13279), .Z(n12612) );
  NOR2_X1 U14933 ( .A1(n12613), .A2(n12612), .ZN(n12635) );
  AOI211_X1 U14934 ( .C1(n12613), .C2(n12612), .A(n14920), .B(n12635), .ZN(
        n12614) );
  AOI211_X1 U14935 ( .C1(n14926), .C2(n7059), .A(n12615), .B(n12614), .ZN(
        n12625) );
  NAND2_X1 U14936 ( .A1(n12616), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12617) );
  NOR2_X1 U14937 ( .A1(n12622), .A2(n12621), .ZN(n12647) );
  AOI21_X1 U14938 ( .B1(n12622), .B2(n12621), .A(n12647), .ZN(n12623) );
  OR2_X1 U14939 ( .A1(n12623), .A2(n15547), .ZN(n12624) );
  OAI211_X1 U14940 ( .C1(n12626), .C2(n15541), .A(n12625), .B(n12624), .ZN(
        P3_U3196) );
  NOR2_X1 U14941 ( .A1(n12649), .A2(n12628), .ZN(n12629) );
  INV_X1 U14942 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14885) );
  INV_X1 U14943 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13198) );
  XNOR2_X1 U14944 ( .A(n12652), .B(n13198), .ZN(n14909) );
  OR2_X1 U14945 ( .A1(n12652), .A2(n13198), .ZN(n12638) );
  NOR2_X1 U14946 ( .A1(n14925), .A2(n6657), .ZN(n12630) );
  INV_X1 U14947 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13194) );
  INV_X1 U14948 ( .A(n14925), .ZN(n12641) );
  NAND2_X1 U14949 ( .A1(n12657), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12664) );
  OAI21_X1 U14950 ( .B1(n12657), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12664), 
        .ZN(n12631) );
  AOI21_X1 U14951 ( .B1(n12632), .B2(n12631), .A(n6656), .ZN(n12663) );
  INV_X1 U14952 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12634) );
  OAI21_X1 U14953 ( .B1(n15529), .B2(n12634), .A(n12633), .ZN(n12646) );
  MUX2_X1 U14954 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13279), .Z(n12644) );
  MUX2_X1 U14955 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13279), .Z(n12642) );
  MUX2_X1 U14956 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13279), .Z(n12636) );
  XNOR2_X1 U14957 ( .A(n12637), .B(n12649), .ZN(n14881) );
  MUX2_X1 U14958 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13279), .Z(n14882) );
  NOR2_X1 U14959 ( .A1(n14881), .A2(n14882), .ZN(n14880) );
  AOI21_X1 U14960 ( .B1(n12637), .B2(n12649), .A(n14880), .ZN(n14899) );
  OR2_X1 U14961 ( .A1(n12652), .A2(n13162), .ZN(n12654) );
  MUX2_X1 U14962 ( .A(n12654), .B(n12638), .S(n13279), .Z(n14896) );
  INV_X1 U14963 ( .A(n14896), .ZN(n12640) );
  MUX2_X1 U14964 ( .A(n13162), .B(n13198), .S(n13279), .Z(n12639) );
  NAND2_X1 U14965 ( .A1(n12639), .A2(n12652), .ZN(n14897) );
  XOR2_X1 U14966 ( .A(n12642), .B(n14925), .Z(n14922) );
  NOR2_X1 U14967 ( .A1(n14921), .A2(n14922), .ZN(n14919) );
  AOI21_X1 U14968 ( .B1(n12642), .B2(n12641), .A(n14919), .ZN(n12667) );
  XNOR2_X1 U14969 ( .A(n12667), .B(n12666), .ZN(n12643) );
  NOR2_X1 U14970 ( .A1(n12643), .A2(n12644), .ZN(n12665) );
  AOI211_X1 U14971 ( .C1(n14926), .C2(n12666), .A(n12646), .B(n12645), .ZN(
        n12662) );
  NOR2_X1 U14972 ( .A1(n12649), .A2(n12650), .ZN(n12651) );
  NAND2_X1 U14973 ( .A1(n12652), .A2(n13162), .ZN(n12653) );
  NAND2_X1 U14974 ( .A1(n12654), .A2(n12653), .ZN(n14894) );
  NOR2_X1 U14975 ( .A1(n14925), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U14976 ( .A1(n12657), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12674) );
  OAI21_X1 U14977 ( .B1(n12657), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12674), 
        .ZN(n12658) );
  AOI21_X1 U14978 ( .B1(n12659), .B2(n12658), .A(n12676), .ZN(n12660) );
  OAI211_X1 U14979 ( .C1(n12663), .C2(n15541), .A(n12662), .B(n12661), .ZN(
        P3_U3200) );
  XNOR2_X1 U14980 ( .A(n12673), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12668) );
  AOI21_X1 U14981 ( .B1(n12667), .B2(n12666), .A(n12665), .ZN(n12670) );
  XNOR2_X1 U14982 ( .A(n12673), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12677) );
  MUX2_X1 U14983 ( .A(n12668), .B(n12677), .S(n7134), .Z(n12669) );
  XNOR2_X1 U14984 ( .A(n12670), .B(n12669), .ZN(n12680) );
  NAND2_X1 U14985 ( .A1(n15458), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12671) );
  OAI211_X1 U14986 ( .C1(n15531), .C2(n12673), .A(n12672), .B(n12671), .ZN(
        n12679) );
  INV_X1 U14987 ( .A(n12674), .ZN(n12675) );
  NOR2_X1 U14988 ( .A1(n12676), .A2(n12675), .ZN(n12678) );
  INV_X1 U14989 ( .A(n12681), .ZN(n12687) );
  AOI22_X1 U14990 ( .A1(n14943), .A2(P3_REG2_REG_29__SCAN_IN), .B1(n14939), 
        .B2(n14938), .ZN(n12682) );
  OAI21_X1 U14991 ( .B1(n12683), .B2(n12870), .A(n12682), .ZN(n12684) );
  AOI21_X1 U14992 ( .B1(n12685), .B2(n12872), .A(n12684), .ZN(n12686) );
  OAI21_X1 U14993 ( .B1(n12687), .B2(n14943), .A(n12686), .ZN(P3_U3204) );
  INV_X1 U14994 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12689) );
  OAI22_X1 U14995 ( .A1(n15566), .A2(n12689), .B1(n12688), .B2(n15553), .ZN(
        n12690) );
  AOI21_X1 U14996 ( .B1(n12691), .B2(n14944), .A(n12690), .ZN(n12694) );
  NAND2_X1 U14997 ( .A1(n12692), .A2(n12872), .ZN(n12693) );
  OAI211_X1 U14998 ( .C1(n12695), .C2(n14943), .A(n12694), .B(n12693), .ZN(
        P3_U3205) );
  INV_X1 U14999 ( .A(n12696), .ZN(n12705) );
  NAND2_X1 U15000 ( .A1(n12697), .A2(n15566), .ZN(n12703) );
  OAI22_X1 U15001 ( .A1(n15566), .A2(n12699), .B1(n12698), .B2(n15553), .ZN(
        n12700) );
  AOI21_X1 U15002 ( .B1(n12701), .B2(n14944), .A(n12700), .ZN(n12702) );
  OAI211_X1 U15003 ( .C1(n12705), .C2(n12704), .A(n12703), .B(n12702), .ZN(
        P3_U3206) );
  OAI21_X1 U15004 ( .B1(n12708), .B2(n12707), .A(n12706), .ZN(n12875) );
  XOR2_X1 U15005 ( .A(n12709), .B(n12708), .Z(n12711) );
  OAI21_X1 U15006 ( .B1(n12711), .B2(n15560), .A(n12710), .ZN(n12876) );
  NAND2_X1 U15007 ( .A1(n12876), .A2(n15566), .ZN(n12717) );
  OAI22_X1 U15008 ( .A1(n15566), .A2(n12713), .B1(n12712), .B2(n15553), .ZN(
        n12714) );
  AOI21_X1 U15009 ( .B1(n12715), .B2(n14944), .A(n12714), .ZN(n12716) );
  OAI211_X1 U15010 ( .C1(n12857), .C2(n12875), .A(n12717), .B(n12716), .ZN(
        P3_U3207) );
  OAI211_X1 U15011 ( .C1(n12720), .C2(n12719), .A(n12718), .B(n12861), .ZN(
        n12723) );
  INV_X1 U15012 ( .A(n12721), .ZN(n12722) );
  NAND2_X1 U15013 ( .A1(n12723), .A2(n12722), .ZN(n12880) );
  INV_X1 U15014 ( .A(n12880), .ZN(n12733) );
  OAI21_X1 U15015 ( .B1(n12726), .B2(n12725), .A(n12724), .ZN(n12881) );
  INV_X1 U15016 ( .A(n12727), .ZN(n13223) );
  NOR2_X1 U15017 ( .A1(n13223), .A2(n12870), .ZN(n12731) );
  OAI22_X1 U15018 ( .A1(n15566), .A2(n12729), .B1(n12728), .B2(n15553), .ZN(
        n12730) );
  AOI211_X1 U15019 ( .C1(n12881), .C2(n12872), .A(n12731), .B(n12730), .ZN(
        n12732) );
  OAI21_X1 U15020 ( .B1(n12733), .B2(n14943), .A(n12732), .ZN(P3_U3208) );
  OAI211_X1 U15021 ( .C1(n12736), .C2(n12735), .A(n12734), .B(n12861), .ZN(
        n12739) );
  INV_X1 U15022 ( .A(n12737), .ZN(n12738) );
  OR2_X1 U15023 ( .A1(n12741), .A2(n12740), .ZN(n12742) );
  NAND2_X1 U15024 ( .A1(n12743), .A2(n12742), .ZN(n12884) );
  NOR2_X1 U15025 ( .A1(n13227), .A2(n12870), .ZN(n12748) );
  OAI22_X1 U15026 ( .A1(n15566), .A2(n12746), .B1(n12745), .B2(n15553), .ZN(
        n12747) );
  AOI211_X1 U15027 ( .C1(n12884), .C2(n12872), .A(n12748), .B(n12747), .ZN(
        n12749) );
  OAI21_X1 U15028 ( .B1(n12886), .B2(n14943), .A(n12749), .ZN(P3_U3209) );
  AOI21_X1 U15029 ( .B1(n12750), .B2(n12759), .A(n15560), .ZN(n12753) );
  AOI21_X1 U15030 ( .B1(n12753), .B2(n12752), .A(n12751), .ZN(n12891) );
  OAI22_X1 U15031 ( .A1(n15566), .A2(n12755), .B1(n12754), .B2(n15553), .ZN(
        n12756) );
  AOI21_X1 U15032 ( .B1(n12757), .B2(n14944), .A(n12756), .ZN(n12761) );
  XOR2_X1 U15033 ( .A(n12759), .B(n12758), .Z(n12889) );
  NAND2_X1 U15034 ( .A1(n12889), .A2(n12872), .ZN(n12760) );
  OAI211_X1 U15035 ( .C1(n12891), .C2(n14943), .A(n12761), .B(n12760), .ZN(
        P3_U3210) );
  XNOR2_X1 U15036 ( .A(n12762), .B(n12766), .ZN(n12765) );
  INV_X1 U15037 ( .A(n12763), .ZN(n12764) );
  OAI21_X1 U15038 ( .B1(n12765), .B2(n15560), .A(n12764), .ZN(n12893) );
  INV_X1 U15039 ( .A(n12893), .ZN(n12774) );
  XNOR2_X1 U15040 ( .A(n6787), .B(n12766), .ZN(n12894) );
  INV_X1 U15041 ( .A(n12768), .ZN(n13232) );
  NOR2_X1 U15042 ( .A1(n13232), .A2(n12870), .ZN(n12772) );
  OAI22_X1 U15043 ( .A1(n15566), .A2(n12770), .B1(n12769), .B2(n15553), .ZN(
        n12771) );
  AOI211_X1 U15044 ( .C1(n12894), .C2(n12872), .A(n12772), .B(n12771), .ZN(
        n12773) );
  OAI21_X1 U15045 ( .B1(n12774), .B2(n14943), .A(n12773), .ZN(P3_U3211) );
  XNOR2_X1 U15046 ( .A(n12775), .B(n12779), .ZN(n12778) );
  INV_X1 U15047 ( .A(n12776), .ZN(n12777) );
  OAI21_X1 U15048 ( .B1(n12778), .B2(n15560), .A(n12777), .ZN(n12897) );
  INV_X1 U15049 ( .A(n12897), .ZN(n12786) );
  XNOR2_X1 U15050 ( .A(n12780), .B(n12779), .ZN(n12898) );
  INV_X1 U15051 ( .A(n12781), .ZN(n13236) );
  AOI22_X1 U15052 ( .A1(n14943), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14938), 
        .B2(n12782), .ZN(n12783) );
  OAI21_X1 U15053 ( .B1(n13236), .B2(n12870), .A(n12783), .ZN(n12784) );
  AOI21_X1 U15054 ( .B1(n12898), .B2(n12872), .A(n12784), .ZN(n12785) );
  OAI21_X1 U15055 ( .B1(n12786), .B2(n14943), .A(n12785), .ZN(P3_U3212) );
  NAND3_X1 U15056 ( .A1(n12803), .A2(n12788), .A3(n12787), .ZN(n12789) );
  NAND3_X1 U15057 ( .A1(n12790), .A2(n12861), .A3(n12789), .ZN(n12792) );
  NAND2_X1 U15058 ( .A1(n12792), .A2(n12791), .ZN(n12901) );
  INV_X1 U15059 ( .A(n12901), .ZN(n12801) );
  INV_X1 U15060 ( .A(n12793), .ZN(n12794) );
  AOI21_X1 U15061 ( .B1(n12796), .B2(n12795), .A(n12794), .ZN(n12902) );
  AOI22_X1 U15062 ( .A1(n14943), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14938), 
        .B2(n12797), .ZN(n12798) );
  OAI21_X1 U15063 ( .B1(n13240), .B2(n12870), .A(n12798), .ZN(n12799) );
  AOI21_X1 U15064 ( .B1(n12902), .B2(n12872), .A(n12799), .ZN(n12800) );
  OAI21_X1 U15065 ( .B1(n12801), .B2(n14943), .A(n12800), .ZN(P3_U3213) );
  XOR2_X1 U15066 ( .A(n12802), .B(n12804), .Z(n12906) );
  INV_X1 U15067 ( .A(n12906), .ZN(n12813) );
  NAND2_X1 U15068 ( .A1(n12803), .A2(n12861), .ZN(n12808) );
  AOI21_X1 U15069 ( .B1(n12816), .B2(n12805), .A(n12804), .ZN(n12807) );
  OAI21_X1 U15070 ( .B1(n12808), .B2(n12807), .A(n12806), .ZN(n12905) );
  AOI22_X1 U15071 ( .A1(n14943), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14938), 
        .B2(n12809), .ZN(n12810) );
  OAI21_X1 U15072 ( .B1(n13244), .B2(n12870), .A(n12810), .ZN(n12811) );
  AOI21_X1 U15073 ( .B1(n12905), .B2(n15566), .A(n12811), .ZN(n12812) );
  OAI21_X1 U15074 ( .B1(n12857), .B2(n12813), .A(n12812), .ZN(P3_U3214) );
  NAND2_X1 U15075 ( .A1(n12814), .A2(n7559), .ZN(n12815) );
  NAND2_X1 U15076 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  NAND2_X1 U15077 ( .A1(n12817), .A2(n12861), .ZN(n12819) );
  NAND2_X1 U15078 ( .A1(n12819), .A2(n12818), .ZN(n12913) );
  INV_X1 U15079 ( .A(n12913), .ZN(n12826) );
  XNOR2_X1 U15080 ( .A(n12820), .B(n7559), .ZN(n12909) );
  INV_X1 U15081 ( .A(n12910), .ZN(n12823) );
  AOI22_X1 U15082 ( .A1(n14943), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14938), 
        .B2(n12821), .ZN(n12822) );
  OAI21_X1 U15083 ( .B1(n12823), .B2(n12870), .A(n12822), .ZN(n12824) );
  AOI21_X1 U15084 ( .B1(n12909), .B2(n12872), .A(n12824), .ZN(n12825) );
  OAI21_X1 U15085 ( .B1(n12826), .B2(n14943), .A(n12825), .ZN(P3_U3215) );
  OAI211_X1 U15086 ( .C1(n12829), .C2(n12828), .A(n12827), .B(n12861), .ZN(
        n12833) );
  AOI22_X1 U15087 ( .A1(n12831), .A2(n12849), .B1(n8165), .B2(n12830), .ZN(
        n12832) );
  NAND2_X1 U15088 ( .A1(n12833), .A2(n12832), .ZN(n13192) );
  INV_X1 U15089 ( .A(n13192), .ZN(n12841) );
  XNOR2_X1 U15090 ( .A(n12834), .B(n7552), .ZN(n13193) );
  INV_X1 U15091 ( .A(n12835), .ZN(n13249) );
  INV_X1 U15092 ( .A(n12836), .ZN(n12837) );
  AOI22_X1 U15093 ( .A1(n14943), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14938), 
        .B2(n12837), .ZN(n12838) );
  OAI21_X1 U15094 ( .B1(n13249), .B2(n12870), .A(n12838), .ZN(n12839) );
  AOI21_X1 U15095 ( .B1(n13193), .B2(n12872), .A(n12839), .ZN(n12840) );
  OAI21_X1 U15096 ( .B1(n12841), .B2(n14943), .A(n12840), .ZN(P3_U3216) );
  XNOR2_X1 U15097 ( .A(n12843), .B(n12842), .ZN(n13197) );
  INV_X1 U15098 ( .A(n13197), .ZN(n12856) );
  OAI211_X1 U15099 ( .C1(n12846), .C2(n12845), .A(n12844), .B(n12861), .ZN(
        n12851) );
  AOI22_X1 U15100 ( .A1(n12849), .A2(n12848), .B1(n12847), .B2(n8165), .ZN(
        n12850) );
  NAND2_X1 U15101 ( .A1(n12851), .A2(n12850), .ZN(n13196) );
  NOR2_X1 U15102 ( .A1(n13253), .A2(n12870), .ZN(n12854) );
  OAI22_X1 U15103 ( .A1(n15566), .A2(n13162), .B1(n12852), .B2(n15553), .ZN(
        n12853) );
  AOI211_X1 U15104 ( .C1(n13196), .C2(n15566), .A(n12854), .B(n12853), .ZN(
        n12855) );
  OAI21_X1 U15105 ( .B1(n12857), .B2(n12856), .A(n12855), .ZN(P3_U3217) );
  NAND3_X1 U15106 ( .A1(n12859), .A2(n12866), .A3(n12858), .ZN(n12860) );
  NAND3_X1 U15107 ( .A1(n12862), .A2(n12861), .A3(n12860), .ZN(n12864) );
  NAND2_X1 U15108 ( .A1(n12864), .A2(n12863), .ZN(n13200) );
  INV_X1 U15109 ( .A(n13200), .ZN(n12874) );
  OAI21_X1 U15110 ( .B1(n6786), .B2(n12866), .A(n12865), .ZN(n13201) );
  AOI22_X1 U15111 ( .A1(n14943), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14938), 
        .B2(n12868), .ZN(n12869) );
  OAI21_X1 U15112 ( .B1(n13257), .B2(n12870), .A(n12869), .ZN(n12871) );
  AOI21_X1 U15113 ( .B1(n13201), .B2(n12872), .A(n12871), .ZN(n12873) );
  OAI21_X1 U15114 ( .B1(n12874), .B2(n14943), .A(n12873), .ZN(P3_U3218) );
  INV_X1 U15115 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12878) );
  INV_X1 U15116 ( .A(n12875), .ZN(n12877) );
  AOI21_X1 U15117 ( .B1(n12877), .B2(n15600), .A(n12876), .ZN(n13216) );
  MUX2_X1 U15118 ( .A(n12878), .B(n13216), .S(n15631), .Z(n12879) );
  OAI21_X1 U15119 ( .B1(n13219), .B2(n13211), .A(n12879), .ZN(P3_U3485) );
  INV_X1 U15120 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12882) );
  AOI21_X1 U15121 ( .B1(n15600), .B2(n12881), .A(n12880), .ZN(n13220) );
  MUX2_X1 U15122 ( .A(n12882), .B(n13220), .S(n15631), .Z(n12883) );
  OAI21_X1 U15123 ( .B1(n13223), .B2(n13211), .A(n12883), .ZN(P3_U3484) );
  INV_X1 U15124 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12887) );
  NAND2_X1 U15125 ( .A1(n12884), .A2(n15600), .ZN(n12885) );
  AND2_X1 U15126 ( .A1(n12886), .A2(n12885), .ZN(n13224) );
  MUX2_X1 U15127 ( .A(n12887), .B(n13224), .S(n15631), .Z(n12888) );
  OAI21_X1 U15128 ( .B1(n13227), .B2(n13211), .A(n12888), .ZN(P3_U3483) );
  NAND2_X1 U15129 ( .A1(n12889), .A2(n15600), .ZN(n12890) );
  OAI211_X1 U15130 ( .C1(n12892), .C2(n15606), .A(n12891), .B(n12890), .ZN(
        n13228) );
  MUX2_X1 U15131 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13228), .S(n15631), .Z(
        P3_U3482) );
  INV_X1 U15132 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12895) );
  AOI21_X1 U15133 ( .B1(n12894), .B2(n15600), .A(n12893), .ZN(n13229) );
  MUX2_X1 U15134 ( .A(n12895), .B(n13229), .S(n15631), .Z(n12896) );
  OAI21_X1 U15135 ( .B1(n13232), .B2(n13211), .A(n12896), .ZN(P3_U3481) );
  INV_X1 U15136 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12899) );
  AOI21_X1 U15137 ( .B1(n12898), .B2(n15600), .A(n12897), .ZN(n13233) );
  MUX2_X1 U15138 ( .A(n12899), .B(n13233), .S(n15631), .Z(n12900) );
  OAI21_X1 U15139 ( .B1(n13236), .B2(n13211), .A(n12900), .ZN(P3_U3480) );
  INV_X1 U15140 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12903) );
  AOI21_X1 U15141 ( .B1(n12902), .B2(n15600), .A(n12901), .ZN(n13237) );
  MUX2_X1 U15142 ( .A(n12903), .B(n13237), .S(n15631), .Z(n12904) );
  OAI21_X1 U15143 ( .B1(n13240), .B2(n13211), .A(n12904), .ZN(P3_U3479) );
  INV_X1 U15144 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12907) );
  AOI21_X1 U15145 ( .B1(n12906), .B2(n15600), .A(n12905), .ZN(n13241) );
  MUX2_X1 U15146 ( .A(n12907), .B(n13241), .S(n15631), .Z(n12908) );
  OAI21_X1 U15147 ( .B1(n13211), .B2(n13244), .A(n12908), .ZN(P3_U3478) );
  AND2_X1 U15148 ( .A1(n12909), .A2(n15600), .ZN(n12912) );
  AND2_X1 U15149 ( .A1(n12910), .A2(n14950), .ZN(n12911) );
  MUX2_X1 U15150 ( .A(n13245), .B(P3_REG1_REG_18__SCAN_IN), .S(n15628), .Z(
        n13191) );
  INV_X1 U15151 ( .A(keyinput15), .ZN(n13150) );
  NAND4_X1 U15152 ( .A1(keyinput70), .A2(keyinput68), .A3(keyinput9), .A4(
        n13150), .ZN(n12960) );
  NOR2_X1 U15153 ( .A1(keyinput34), .A2(keyinput113), .ZN(n12914) );
  NAND3_X1 U15154 ( .A1(keyinput2), .A2(keyinput48), .A3(n12914), .ZN(n12959)
         );
  NOR2_X1 U15155 ( .A1(keyinput29), .A2(keyinput79), .ZN(n12915) );
  NAND3_X1 U15156 ( .A1(keyinput107), .A2(keyinput106), .A3(n12915), .ZN(
        n12916) );
  NOR3_X1 U15157 ( .A1(keyinput95), .A2(keyinput5), .A3(n12916), .ZN(n12924)
         );
  INV_X1 U15158 ( .A(keyinput6), .ZN(n13161) );
  NAND4_X1 U15159 ( .A1(keyinput118), .A2(keyinput81), .A3(keyinput66), .A4(
        n13161), .ZN(n12922) );
  OR4_X1 U15160 ( .A1(keyinput86), .A2(keyinput8), .A3(keyinput109), .A4(
        keyinput64), .ZN(n12921) );
  NOR2_X1 U15161 ( .A1(keyinput71), .A2(keyinput115), .ZN(n12917) );
  NAND3_X1 U15162 ( .A1(keyinput87), .A2(keyinput94), .A3(n12917), .ZN(n12920)
         );
  INV_X1 U15163 ( .A(keyinput77), .ZN(n12918) );
  NAND4_X1 U15164 ( .A1(keyinput13), .A2(keyinput37), .A3(keyinput121), .A4(
        n12918), .ZN(n12919) );
  NOR4_X1 U15165 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12923) );
  NAND4_X1 U15166 ( .A1(keyinput16), .A2(keyinput75), .A3(n12924), .A4(n12923), 
        .ZN(n12958) );
  NAND2_X1 U15167 ( .A1(keyinput32), .A2(keyinput31), .ZN(n12925) );
  NOR3_X1 U15168 ( .A1(keyinput28), .A2(keyinput21), .A3(n12925), .ZN(n12926)
         );
  NAND3_X1 U15169 ( .A1(keyinput127), .A2(keyinput49), .A3(n12926), .ZN(n12940) );
  INV_X1 U15170 ( .A(keyinput56), .ZN(n12927) );
  NAND4_X1 U15171 ( .A1(keyinput26), .A2(keyinput125), .A3(keyinput91), .A4(
        n12927), .ZN(n12928) );
  NOR3_X1 U15172 ( .A1(keyinput54), .A2(keyinput97), .A3(n12928), .ZN(n12938)
         );
  INV_X1 U15173 ( .A(keyinput40), .ZN(n12929) );
  NAND4_X1 U15174 ( .A1(keyinput100), .A2(keyinput108), .A3(keyinput7), .A4(
        n12929), .ZN(n12936) );
  NOR2_X1 U15175 ( .A1(keyinput119), .A2(keyinput3), .ZN(n12930) );
  NAND3_X1 U15176 ( .A1(keyinput58), .A2(keyinput23), .A3(n12930), .ZN(n12935)
         );
  NOR2_X1 U15177 ( .A1(keyinput89), .A2(keyinput55), .ZN(n12931) );
  NAND3_X1 U15178 ( .A1(keyinput96), .A2(keyinput10), .A3(n12931), .ZN(n12934)
         );
  NOR2_X1 U15179 ( .A1(keyinput41), .A2(keyinput69), .ZN(n12932) );
  NAND3_X1 U15180 ( .A1(keyinput62), .A2(keyinput110), .A3(n12932), .ZN(n12933) );
  NOR4_X1 U15181 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12937) );
  NAND4_X1 U15182 ( .A1(keyinput65), .A2(keyinput24), .A3(n12938), .A4(n12937), 
        .ZN(n12939) );
  NOR4_X1 U15183 ( .A1(keyinput111), .A2(keyinput53), .A3(n12940), .A4(n12939), 
        .ZN(n12956) );
  NAND2_X1 U15184 ( .A1(keyinput46), .A2(keyinput33), .ZN(n12941) );
  NOR3_X1 U15185 ( .A1(keyinput112), .A2(keyinput92), .A3(n12941), .ZN(n12955)
         );
  INV_X1 U15186 ( .A(keyinput30), .ZN(n12942) );
  NOR4_X1 U15187 ( .A1(keyinput82), .A2(keyinput18), .A3(keyinput124), .A4(
        n12942), .ZN(n12954) );
  NAND2_X1 U15188 ( .A1(keyinput73), .A2(keyinput22), .ZN(n12943) );
  NOR3_X1 U15189 ( .A1(keyinput103), .A2(keyinput42), .A3(n12943), .ZN(n12944)
         );
  NAND3_X1 U15190 ( .A1(keyinput38), .A2(keyinput84), .A3(n12944), .ZN(n12952)
         );
  NAND4_X1 U15191 ( .A1(keyinput101), .A2(keyinput47), .A3(keyinput35), .A4(
        keyinput17), .ZN(n12950) );
  NOR2_X1 U15192 ( .A1(keyinput99), .A2(keyinput72), .ZN(n12945) );
  NAND3_X1 U15193 ( .A1(keyinput52), .A2(keyinput27), .A3(n12945), .ZN(n12949)
         );
  NOR3_X1 U15194 ( .A1(keyinput78), .A2(keyinput36), .A3(keyinput67), .ZN(
        n12946) );
  NAND2_X1 U15195 ( .A1(keyinput74), .A2(n12946), .ZN(n12948) );
  NAND4_X1 U15196 ( .A1(keyinput114), .A2(keyinput105), .A3(keyinput120), .A4(
        keyinput102), .ZN(n12947) );
  OR4_X1 U15197 ( .A1(n12950), .A2(n12949), .A3(n12948), .A4(n12947), .ZN(
        n12951) );
  NOR4_X1 U15198 ( .A1(keyinput93), .A2(keyinput39), .A3(n12952), .A4(n12951), 
        .ZN(n12953) );
  NAND4_X1 U15199 ( .A1(n12956), .A2(n12955), .A3(n12954), .A4(n12953), .ZN(
        n12957) );
  NOR4_X1 U15200 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n13189) );
  NAND2_X1 U15201 ( .A1(keyinput0), .A2(keyinput14), .ZN(n12961) );
  NOR3_X1 U15202 ( .A1(keyinput19), .A2(keyinput43), .A3(n12961), .ZN(n12962)
         );
  NAND3_X1 U15203 ( .A1(keyinput90), .A2(keyinput123), .A3(n12962), .ZN(n12974) );
  NOR2_X1 U15204 ( .A1(keyinput12), .A2(keyinput85), .ZN(n12963) );
  NAND3_X1 U15205 ( .A1(keyinput61), .A2(keyinput11), .A3(n12963), .ZN(n12964)
         );
  NOR3_X1 U15206 ( .A1(keyinput98), .A2(keyinput104), .A3(n12964), .ZN(n12972)
         );
  INV_X1 U15207 ( .A(keyinput88), .ZN(n13062) );
  NAND4_X1 U15208 ( .A1(keyinput1), .A2(keyinput117), .A3(keyinput25), .A4(
        n13062), .ZN(n12970) );
  OR4_X1 U15209 ( .A1(keyinput83), .A2(keyinput126), .A3(keyinput57), .A4(
        keyinput80), .ZN(n12969) );
  INV_X1 U15210 ( .A(keyinput63), .ZN(n12965) );
  NAND4_X1 U15211 ( .A1(keyinput116), .A2(keyinput60), .A3(keyinput20), .A4(
        n12965), .ZN(n12968) );
  NOR2_X1 U15212 ( .A1(keyinput59), .A2(keyinput4), .ZN(n12966) );
  NAND3_X1 U15213 ( .A1(keyinput76), .A2(keyinput122), .A3(n12966), .ZN(n12967) );
  NOR4_X1 U15214 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n12971) );
  NAND4_X1 U15215 ( .A1(keyinput50), .A2(keyinput44), .A3(n12972), .A4(n12971), 
        .ZN(n12973) );
  NOR4_X1 U15216 ( .A1(keyinput45), .A2(keyinput51), .A3(n12974), .A4(n12973), 
        .ZN(n13188) );
  INV_X1 U15217 ( .A(SI_22_), .ZN(n12976) );
  AOI22_X1 U15218 ( .A1(n9526), .A2(keyinput59), .B1(n12976), .B2(keyinput122), 
        .ZN(n12975) );
  OAI221_X1 U15219 ( .B1(n9526), .B2(keyinput59), .C1(n12976), .C2(keyinput122), .A(n12975), .ZN(n12984) );
  INV_X1 U15220 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U15221 ( .A1(n15109), .A2(keyinput12), .B1(n12978), .B2(keyinput61), 
        .ZN(n12977) );
  OAI221_X1 U15222 ( .B1(n15109), .B2(keyinput12), .C1(n12978), .C2(keyinput61), .A(n12977), .ZN(n12983) );
  INV_X1 U15223 ( .A(keyinput105), .ZN(n12979) );
  XNOR2_X1 U15224 ( .A(n12979), .B(P3_ADDR_REG_14__SCAN_IN), .ZN(n12982) );
  INV_X1 U15225 ( .A(keyinput14), .ZN(n12980) );
  XNOR2_X1 U15226 ( .A(n12980), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n12981) );
  NOR4_X1 U15227 ( .A1(n12984), .A2(n12983), .A3(n12982), .A4(n12981), .ZN(
        n13019) );
  INV_X1 U15228 ( .A(keyinput60), .ZN(n12986) );
  OAI22_X1 U15229 ( .A1(n12987), .A2(keyinput116), .B1(n12986), .B2(
        P3_DATAO_REG_26__SCAN_IN), .ZN(n12985) );
  AOI221_X1 U15230 ( .B1(n12987), .B2(keyinput116), .C1(
        P3_DATAO_REG_26__SCAN_IN), .C2(n12986), .A(n12985), .ZN(n13018) );
  INV_X1 U15231 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U15232 ( .A1(n15099), .A2(keyinput54), .B1(keyinput97), .B2(n15065), 
        .ZN(n12988) );
  OAI221_X1 U15233 ( .B1(n15099), .B2(keyinput54), .C1(n15065), .C2(keyinput97), .A(n12988), .ZN(n12995) );
  AOI22_X1 U15234 ( .A1(n12699), .A2(keyinput16), .B1(n12990), .B2(keyinput75), 
        .ZN(n12989) );
  OAI221_X1 U15235 ( .B1(n12699), .B2(keyinput16), .C1(n12990), .C2(keyinput75), .A(n12989), .ZN(n12994) );
  INV_X1 U15236 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U15237 ( .A1(n14856), .A2(keyinput30), .B1(n12992), .B2(keyinput18), 
        .ZN(n12991) );
  OAI221_X1 U15238 ( .B1(n14856), .B2(keyinput30), .C1(n12992), .C2(keyinput18), .A(n12991), .ZN(n12993) );
  OR3_X1 U15239 ( .A1(n12995), .A2(n12994), .A3(n12993), .ZN(n13002) );
  INV_X1 U15240 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U15241 ( .A1(n12997), .A2(keyinput65), .B1(keyinput24), .B2(n11002), 
        .ZN(n12996) );
  OAI221_X1 U15242 ( .B1(n12997), .B2(keyinput65), .C1(n11002), .C2(keyinput24), .A(n12996), .ZN(n13001) );
  INV_X1 U15243 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U15244 ( .A1(n12999), .A2(keyinput113), .B1(keyinput48), .B2(n9493), 
        .ZN(n12998) );
  OAI221_X1 U15245 ( .B1(n12999), .B2(keyinput113), .C1(n9493), .C2(keyinput48), .A(n12998), .ZN(n13000) );
  NOR3_X1 U15246 ( .A1(n13002), .A2(n13001), .A3(n13000), .ZN(n13017) );
  INV_X1 U15247 ( .A(keyinput87), .ZN(n13003) );
  XNOR2_X1 U15248 ( .A(n13003), .B(P1_ADDR_REG_0__SCAN_IN), .ZN(n13015) );
  INV_X1 U15249 ( .A(keyinput121), .ZN(n13004) );
  XNOR2_X1 U15250 ( .A(n13004), .B(P3_DATAO_REG_22__SCAN_IN), .ZN(n13014) );
  XNOR2_X1 U15251 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput120), .ZN(n13008) );
  XNOR2_X1 U15252 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput70), .ZN(n13007) );
  XNOR2_X1 U15253 ( .A(P1_REG2_REG_16__SCAN_IN), .B(keyinput1), .ZN(n13006) );
  XNOR2_X1 U15254 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput77), .ZN(n13005) );
  NAND4_X1 U15255 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13013) );
  XNOR2_X1 U15256 ( .A(SI_6_), .B(keyinput115), .ZN(n13011) );
  XNOR2_X1 U15257 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput99), .ZN(n13010)
         );
  XNOR2_X1 U15258 ( .A(keyinput35), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n13009)
         );
  NAND3_X1 U15259 ( .A1(n13011), .A2(n13010), .A3(n13009), .ZN(n13012) );
  NOR4_X1 U15260 ( .A1(n13015), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13016) );
  NAND4_X1 U15261 ( .A1(n13019), .A2(n13018), .A3(n13017), .A4(n13016), .ZN(
        n13086) );
  INV_X1 U15262 ( .A(keyinput2), .ZN(n13021) );
  AOI22_X1 U15263 ( .A1(n13603), .A2(keyinput34), .B1(P3_RD_REG_SCAN_IN), .B2(
        n13021), .ZN(n13020) );
  OAI221_X1 U15264 ( .B1(n13603), .B2(keyinput34), .C1(n13021), .C2(
        P3_RD_REG_SCAN_IN), .A(n13020), .ZN(n13025) );
  INV_X1 U15265 ( .A(keyinput125), .ZN(n13023) );
  AOI22_X1 U15266 ( .A1(n10700), .A2(keyinput91), .B1(P3_DATAO_REG_23__SCAN_IN), .B2(n13023), .ZN(n13022) );
  OAI221_X1 U15267 ( .B1(n10700), .B2(keyinput91), .C1(n13023), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n13022), .ZN(n13024) );
  NOR2_X1 U15268 ( .A1(n13025), .A2(n13024), .ZN(n13046) );
  INV_X1 U15269 ( .A(keyinput108), .ZN(n13027) );
  AOI22_X1 U15270 ( .A1(n7894), .A2(keyinput7), .B1(P3_DATAO_REG_4__SCAN_IN), 
        .B2(n13027), .ZN(n13026) );
  OAI221_X1 U15271 ( .B1(n7894), .B2(keyinput7), .C1(n13027), .C2(
        P3_DATAO_REG_4__SCAN_IN), .A(n13026), .ZN(n13031) );
  INV_X1 U15272 ( .A(keyinput62), .ZN(n13029) );
  AOI22_X1 U15273 ( .A1(n15620), .A2(keyinput41), .B1(P3_ADDR_REG_8__SCAN_IN), 
        .B2(n13029), .ZN(n13028) );
  OAI221_X1 U15274 ( .B1(n15620), .B2(keyinput41), .C1(n13029), .C2(
        P3_ADDR_REG_8__SCAN_IN), .A(n13028), .ZN(n13030) );
  NOR2_X1 U15275 ( .A1(n13031), .A2(n13030), .ZN(n13045) );
  INV_X1 U15276 ( .A(keyinput98), .ZN(n13033) );
  AOI22_X1 U15277 ( .A1(n13251), .A2(keyinput104), .B1(
        P3_DATAO_REG_21__SCAN_IN), .B2(n13033), .ZN(n13032) );
  OAI221_X1 U15278 ( .B1(n13251), .B2(keyinput104), .C1(n13033), .C2(
        P3_DATAO_REG_21__SCAN_IN), .A(n13032), .ZN(n13038) );
  INV_X1 U15279 ( .A(keyinput90), .ZN(n13035) );
  AOI22_X1 U15280 ( .A1(n13036), .A2(keyinput123), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(n13035), .ZN(n13034) );
  OAI221_X1 U15281 ( .B1(n13036), .B2(keyinput123), .C1(n13035), .C2(
        P3_DATAO_REG_13__SCAN_IN), .A(n13034), .ZN(n13037) );
  NOR2_X1 U15282 ( .A1(n13038), .A2(n13037), .ZN(n13044) );
  INV_X1 U15283 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U15284 ( .A1(n14243), .A2(keyinput89), .B1(n15102), .B2(keyinput96), 
        .ZN(n13039) );
  OAI221_X1 U15285 ( .B1(n14243), .B2(keyinput89), .C1(n15102), .C2(keyinput96), .A(n13039), .ZN(n13042) );
  INV_X1 U15286 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15139) );
  INV_X1 U15287 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U15288 ( .A1(n15139), .A2(keyinput85), .B1(n15116), .B2(keyinput11), 
        .ZN(n13040) );
  OAI221_X1 U15289 ( .B1(n15139), .B2(keyinput85), .C1(n15116), .C2(keyinput11), .A(n13040), .ZN(n13041) );
  NOR2_X1 U15290 ( .A1(n13042), .A2(n13041), .ZN(n13043) );
  NAND4_X1 U15291 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13085) );
  INV_X1 U15292 ( .A(keyinput80), .ZN(n13048) );
  AOI22_X1 U15293 ( .A1(n13049), .A2(keyinput57), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n13048), .ZN(n13047) );
  OAI221_X1 U15294 ( .B1(n13049), .B2(keyinput57), .C1(n13048), .C2(
        P1_ADDR_REG_18__SCAN_IN), .A(n13047), .ZN(n13058) );
  AOI22_X1 U15295 ( .A1(n15355), .A2(keyinput101), .B1(keyinput47), .B2(n12746), .ZN(n13050) );
  OAI221_X1 U15296 ( .B1(n15355), .B2(keyinput101), .C1(n12746), .C2(
        keyinput47), .A(n13050), .ZN(n13057) );
  AOI22_X1 U15297 ( .A1(n10300), .A2(keyinput76), .B1(keyinput4), .B2(n12184), 
        .ZN(n13051) );
  OAI221_X1 U15298 ( .B1(n10300), .B2(keyinput76), .C1(n12184), .C2(keyinput4), 
        .A(n13051), .ZN(n13056) );
  INV_X1 U15299 ( .A(P1_B_REG_SCAN_IN), .ZN(n13054) );
  INV_X1 U15300 ( .A(keyinput83), .ZN(n13053) );
  AOI22_X1 U15301 ( .A1(n13054), .A2(keyinput126), .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n13053), .ZN(n13052) );
  OAI221_X1 U15302 ( .B1(n13054), .B2(keyinput126), .C1(n13053), .C2(
        P3_ADDR_REG_12__SCAN_IN), .A(n13052), .ZN(n13055) );
  OR4_X1 U15303 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n13055), .ZN(
        n13084) );
  INV_X1 U15304 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U15305 ( .A1(n13060), .A2(keyinput27), .B1(keyinput72), .B2(n15101), 
        .ZN(n13059) );
  OAI221_X1 U15306 ( .B1(n13060), .B2(keyinput27), .C1(n15101), .C2(keyinput72), .A(n13059), .ZN(n13065) );
  AOI22_X1 U15307 ( .A1(n13063), .A2(keyinput25), .B1(P1_ADDR_REG_7__SCAN_IN), 
        .B2(n13062), .ZN(n13061) );
  OAI221_X1 U15308 ( .B1(n13063), .B2(keyinput25), .C1(n13062), .C2(
        P1_ADDR_REG_7__SCAN_IN), .A(n13061), .ZN(n13064) );
  NOR2_X1 U15309 ( .A1(n13065), .A2(n13064), .ZN(n13082) );
  XNOR2_X1 U15310 ( .A(keyinput94), .B(n10020), .ZN(n13067) );
  XNOR2_X1 U15311 ( .A(keyinput10), .B(n13790), .ZN(n13066) );
  NOR2_X1 U15312 ( .A1(n13067), .A2(n13066), .ZN(n13081) );
  AOI22_X1 U15313 ( .A1(n13069), .A2(keyinput69), .B1(keyinput110), .B2(n14916), .ZN(n13068) );
  OAI221_X1 U15314 ( .B1(n13069), .B2(keyinput69), .C1(n14916), .C2(
        keyinput110), .A(n13068), .ZN(n13074) );
  AOI22_X1 U15315 ( .A1(n13072), .A2(keyinput29), .B1(keyinput106), .B2(n13071), .ZN(n13070) );
  OAI221_X1 U15316 ( .B1(n13072), .B2(keyinput29), .C1(n13071), .C2(
        keyinput106), .A(n13070), .ZN(n13073) );
  NOR2_X1 U15317 ( .A1(n13074), .A2(n13073), .ZN(n13080) );
  INV_X1 U15318 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U15319 ( .A1(n13077), .A2(keyinput95), .B1(keyinput5), .B2(n13076), 
        .ZN(n13075) );
  OAI221_X1 U15320 ( .B1(n13077), .B2(keyinput95), .C1(n13076), .C2(keyinput5), 
        .A(n13075), .ZN(n13078) );
  INV_X1 U15321 ( .A(n13078), .ZN(n13079) );
  NAND4_X1 U15322 ( .A1(n13082), .A2(n13081), .A3(n13080), .A4(n13079), .ZN(
        n13083) );
  NOR4_X1 U15323 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13158) );
  AOI22_X1 U15324 ( .A1(n10366), .A2(keyinput93), .B1(n12755), .B2(keyinput39), 
        .ZN(n13087) );
  OAI221_X1 U15325 ( .B1(n10366), .B2(keyinput93), .C1(n12755), .C2(keyinput39), .A(n13087), .ZN(n13097) );
  AOI22_X1 U15326 ( .A1(n13538), .A2(keyinput103), .B1(keyinput22), .B2(n13089), .ZN(n13088) );
  OAI221_X1 U15327 ( .B1(n13538), .B2(keyinput103), .C1(n13089), .C2(
        keyinput22), .A(n13088), .ZN(n13096) );
  AOI22_X1 U15328 ( .A1(n8559), .A2(keyinput73), .B1(keyinput42), .B2(n13091), 
        .ZN(n13090) );
  OAI221_X1 U15329 ( .B1(n8559), .B2(keyinput73), .C1(n13091), .C2(keyinput42), 
        .A(n13090), .ZN(n13095) );
  AOI22_X1 U15330 ( .A1(n7723), .A2(keyinput38), .B1(keyinput84), .B2(n13093), 
        .ZN(n13092) );
  OAI221_X1 U15331 ( .B1(n7723), .B2(keyinput38), .C1(n13093), .C2(keyinput84), 
        .A(n13092), .ZN(n13094) );
  NOR4_X1 U15332 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        n13157) );
  INV_X1 U15333 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14814) );
  INV_X1 U15334 ( .A(keyinput20), .ZN(n13099) );
  OAI22_X1 U15335 ( .A1(keyinput63), .A2(n14814), .B1(n13099), .B2(
        P3_DATAO_REG_10__SCAN_IN), .ZN(n13098) );
  AOI221_X1 U15336 ( .B1(n14814), .B2(keyinput63), .C1(n13099), .C2(
        P3_DATAO_REG_10__SCAN_IN), .A(n13098), .ZN(n13156) );
  XNOR2_X1 U15337 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput51), .ZN(n13103)
         );
  XNOR2_X1 U15338 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput68), .ZN(n13102)
         );
  XNOR2_X1 U15339 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput56), .ZN(n13101)
         );
  XNOR2_X1 U15340 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput50), .ZN(n13100) );
  NAND4_X1 U15341 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n13109) );
  XNOR2_X1 U15342 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(keyinput100), .ZN(n13107)
         );
  XNOR2_X1 U15343 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput71), .ZN(n13106) );
  XNOR2_X1 U15344 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput67), .ZN(n13105) );
  XNOR2_X1 U15345 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput52), .ZN(n13104) );
  NAND4_X1 U15346 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13108) );
  NOR2_X1 U15347 ( .A1(n13109), .A2(n13108), .ZN(n13143) );
  XNOR2_X1 U15348 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput114), .ZN(n13113) );
  XNOR2_X1 U15349 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput107), .ZN(n13112) );
  XNOR2_X1 U15350 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput82), .ZN(n13111) );
  XNOR2_X1 U15351 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput9), .ZN(n13110) );
  NAND4_X1 U15352 ( .A1(n13113), .A2(n13112), .A3(n13111), .A4(n13110), .ZN(
        n13119) );
  XNOR2_X1 U15353 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput19), .ZN(n13117) );
  XNOR2_X1 U15354 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput17), .ZN(n13116) );
  XNOR2_X1 U15355 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput23), .ZN(n13115)
         );
  XNOR2_X1 U15356 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput55), .ZN(n13114)
         );
  NAND4_X1 U15357 ( .A1(n13117), .A2(n13116), .A3(n13115), .A4(n13114), .ZN(
        n13118) );
  NOR2_X1 U15358 ( .A1(n13119), .A2(n13118), .ZN(n13142) );
  XNOR2_X1 U15359 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput0), .ZN(n13123) );
  XNOR2_X1 U15360 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput33), .ZN(n13122)
         );
  XNOR2_X1 U15361 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput46), .ZN(n13121) );
  XNOR2_X1 U15362 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput79), .ZN(n13120) );
  NAND4_X1 U15363 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13120), .ZN(
        n13129) );
  XNOR2_X1 U15364 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput119), .ZN(n13127) );
  XNOR2_X1 U15365 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput117), .ZN(n13126) );
  XNOR2_X1 U15366 ( .A(P3_IR_REG_18__SCAN_IN), .B(keyinput36), .ZN(n13125) );
  XNOR2_X1 U15367 ( .A(P3_IR_REG_30__SCAN_IN), .B(keyinput40), .ZN(n13124) );
  NAND4_X1 U15368 ( .A1(n13127), .A2(n13126), .A3(n13125), .A4(n13124), .ZN(
        n13128) );
  NOR2_X1 U15369 ( .A1(n13129), .A2(n13128), .ZN(n13141) );
  XNOR2_X1 U15370 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput26), .ZN(n13133) );
  XNOR2_X1 U15371 ( .A(P3_D_REG_1__SCAN_IN), .B(keyinput45), .ZN(n13132) );
  XNOR2_X1 U15372 ( .A(P3_REG1_REG_29__SCAN_IN), .B(keyinput43), .ZN(n13131)
         );
  XNOR2_X1 U15373 ( .A(P3_REG1_REG_28__SCAN_IN), .B(keyinput44), .ZN(n13130)
         );
  NAND4_X1 U15374 ( .A1(n13133), .A2(n13132), .A3(n13131), .A4(n13130), .ZN(
        n13139) );
  XNOR2_X1 U15375 ( .A(keyinput124), .B(P2_REG2_REG_29__SCAN_IN), .ZN(n13137)
         );
  XNOR2_X1 U15376 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(keyinput3), .ZN(n13136) );
  XNOR2_X1 U15377 ( .A(keyinput102), .B(P1_REG0_REG_6__SCAN_IN), .ZN(n13135)
         );
  XNOR2_X1 U15378 ( .A(keyinput92), .B(P2_REG0_REG_4__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U15379 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13138) );
  NOR2_X1 U15380 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  NAND4_X1 U15381 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13154) );
  INV_X1 U15382 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U15383 ( .A1(n14297), .A2(keyinput78), .B1(n7808), .B2(keyinput74), 
        .ZN(n13144) );
  OAI221_X1 U15384 ( .B1(n14297), .B2(keyinput78), .C1(n7808), .C2(keyinput74), 
        .A(n13144), .ZN(n13149) );
  AOI22_X1 U15385 ( .A1(n15338), .A2(keyinput37), .B1(keyinput13), .B2(n13146), 
        .ZN(n13145) );
  OAI221_X1 U15386 ( .B1(n15338), .B2(keyinput37), .C1(n13146), .C2(keyinput13), .A(n13145), .ZN(n13148) );
  INV_X1 U15387 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15111) );
  XNOR2_X1 U15388 ( .A(n15111), .B(keyinput112), .ZN(n13147) );
  OR3_X1 U15389 ( .A1(n13149), .A2(n13148), .A3(n13147), .ZN(n13153) );
  XNOR2_X1 U15390 ( .A(n15331), .B(keyinput58), .ZN(n13152) );
  XNOR2_X1 U15391 ( .A(n13150), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n13151) );
  NOR4_X1 U15392 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13155) );
  NAND4_X1 U15393 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        n13187) );
  INV_X1 U15394 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U15395 ( .A1(n8776), .A2(keyinput86), .B1(keyinput8), .B2(n15125), 
        .ZN(n13159) );
  OAI221_X1 U15396 ( .B1(n8776), .B2(keyinput86), .C1(n15125), .C2(keyinput8), 
        .A(n13159), .ZN(n13170) );
  AOI22_X1 U15397 ( .A1(n13162), .A2(keyinput118), .B1(P3_ADDR_REG_6__SCAN_IN), 
        .B2(n13161), .ZN(n13160) );
  OAI221_X1 U15398 ( .B1(n13162), .B2(keyinput118), .C1(n13161), .C2(
        P3_ADDR_REG_6__SCAN_IN), .A(n13160), .ZN(n13169) );
  INV_X1 U15399 ( .A(keyinput81), .ZN(n13164) );
  AOI22_X1 U15400 ( .A1(n13882), .A2(keyinput66), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n13164), .ZN(n13163) );
  OAI221_X1 U15401 ( .B1(n13882), .B2(keyinput66), .C1(n13164), .C2(
        P3_ADDR_REG_15__SCAN_IN), .A(n13163), .ZN(n13168) );
  INV_X1 U15402 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U15403 ( .A1(n13166), .A2(keyinput109), .B1(keyinput64), .B2(n15373), .ZN(n13165) );
  OAI221_X1 U15404 ( .B1(n13166), .B2(keyinput109), .C1(n15373), .C2(
        keyinput64), .A(n13165), .ZN(n13167) );
  NOR4_X1 U15405 ( .A1(n13170), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13185) );
  AOI22_X1 U15406 ( .A1(n13173), .A2(keyinput28), .B1(keyinput31), .B2(n13172), 
        .ZN(n13171) );
  OAI221_X1 U15407 ( .B1(n13173), .B2(keyinput28), .C1(n13172), .C2(keyinput31), .A(n13171), .ZN(n13183) );
  AOI22_X1 U15408 ( .A1(n13176), .A2(keyinput111), .B1(n13175), .B2(keyinput53), .ZN(n13174) );
  OAI221_X1 U15409 ( .B1(n13176), .B2(keyinput111), .C1(n13175), .C2(
        keyinput53), .A(n13174), .ZN(n13182) );
  AOI22_X1 U15410 ( .A1(n8578), .A2(keyinput127), .B1(n15334), .B2(keyinput49), 
        .ZN(n13177) );
  OAI221_X1 U15411 ( .B1(n8578), .B2(keyinput127), .C1(n15334), .C2(keyinput49), .A(n13177), .ZN(n13181) );
  AOI22_X1 U15412 ( .A1(n13179), .A2(keyinput32), .B1(n8699), .B2(keyinput21), 
        .ZN(n13178) );
  OAI221_X1 U15413 ( .B1(n13179), .B2(keyinput32), .C1(n8699), .C2(keyinput21), 
        .A(n13178), .ZN(n13180) );
  NOR4_X1 U15414 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13184) );
  NAND2_X1 U15415 ( .A1(n13185), .A2(n13184), .ZN(n13186) );
  AOI211_X1 U15416 ( .C1(n13189), .C2(n13188), .A(n13187), .B(n13186), .ZN(
        n13190) );
  XOR2_X1 U15417 ( .A(n13191), .B(n13190), .Z(P3_U3477) );
  AOI21_X1 U15418 ( .B1(n13193), .B2(n15600), .A(n13192), .ZN(n13246) );
  MUX2_X1 U15419 ( .A(n13194), .B(n13246), .S(n15631), .Z(n13195) );
  OAI21_X1 U15420 ( .B1(n13249), .B2(n13211), .A(n13195), .ZN(P3_U3476) );
  AOI21_X1 U15421 ( .B1(n13197), .B2(n15600), .A(n13196), .ZN(n13250) );
  MUX2_X1 U15422 ( .A(n13198), .B(n13250), .S(n15631), .Z(n13199) );
  OAI21_X1 U15423 ( .B1(n13253), .B2(n13211), .A(n13199), .ZN(P3_U3475) );
  AOI21_X1 U15424 ( .B1(n15600), .B2(n13201), .A(n13200), .ZN(n13254) );
  MUX2_X1 U15425 ( .A(n14885), .B(n13254), .S(n15631), .Z(n13202) );
  OAI21_X1 U15426 ( .B1(n13257), .B2(n13211), .A(n13202), .ZN(P3_U3474) );
  NAND2_X1 U15427 ( .A1(n13203), .A2(n15600), .ZN(n13204) );
  AND2_X1 U15428 ( .A1(n13205), .A2(n13204), .ZN(n13258) );
  MUX2_X1 U15429 ( .A(n7058), .B(n13258), .S(n15631), .Z(n13206) );
  OAI21_X1 U15430 ( .B1(n13211), .B2(n13260), .A(n13206), .ZN(P3_U3473) );
  NAND2_X1 U15431 ( .A1(n13207), .A2(n15600), .ZN(n13208) );
  AND2_X1 U15432 ( .A1(n13209), .A2(n13208), .ZN(n13261) );
  MUX2_X1 U15433 ( .A(n15534), .B(n13261), .S(n15631), .Z(n13210) );
  OAI21_X1 U15434 ( .B1(n13264), .B2(n13211), .A(n13210), .ZN(P3_U3472) );
  OAI21_X1 U15435 ( .B1(n13215), .B2(n13263), .A(n13214), .ZN(P3_U3454) );
  MUX2_X1 U15436 ( .A(n13217), .B(n13216), .S(n15613), .Z(n13218) );
  OAI21_X1 U15437 ( .B1(n13219), .B2(n13263), .A(n13218), .ZN(P3_U3453) );
  MUX2_X1 U15438 ( .A(n13221), .B(n13220), .S(n15613), .Z(n13222) );
  OAI21_X1 U15439 ( .B1(n13223), .B2(n13263), .A(n13222), .ZN(P3_U3452) );
  MUX2_X1 U15440 ( .A(n13225), .B(n13224), .S(n15613), .Z(n13226) );
  OAI21_X1 U15441 ( .B1(n13227), .B2(n13263), .A(n13226), .ZN(P3_U3451) );
  MUX2_X1 U15442 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13228), .S(n15613), .Z(
        P3_U3450) );
  MUX2_X1 U15443 ( .A(n13230), .B(n13229), .S(n15613), .Z(n13231) );
  OAI21_X1 U15444 ( .B1(n13232), .B2(n13263), .A(n13231), .ZN(P3_U3449) );
  INV_X1 U15445 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13234) );
  MUX2_X1 U15446 ( .A(n13234), .B(n13233), .S(n15613), .Z(n13235) );
  OAI21_X1 U15447 ( .B1(n13236), .B2(n13263), .A(n13235), .ZN(P3_U3448) );
  MUX2_X1 U15448 ( .A(n13238), .B(n13237), .S(n15613), .Z(n13239) );
  OAI21_X1 U15449 ( .B1(n13240), .B2(n13263), .A(n13239), .ZN(P3_U3447) );
  MUX2_X1 U15450 ( .A(n13242), .B(n13241), .S(n15613), .Z(n13243) );
  OAI21_X1 U15451 ( .B1(n13263), .B2(n13244), .A(n13243), .ZN(P3_U3446) );
  MUX2_X1 U15452 ( .A(n13245), .B(P3_REG0_REG_18__SCAN_IN), .S(n15612), .Z(
        P3_U3444) );
  MUX2_X1 U15453 ( .A(n13247), .B(n13246), .S(n15613), .Z(n13248) );
  OAI21_X1 U15454 ( .B1(n13249), .B2(n13263), .A(n13248), .ZN(P3_U3441) );
  MUX2_X1 U15455 ( .A(n13251), .B(n13250), .S(n15613), .Z(n13252) );
  OAI21_X1 U15456 ( .B1(n13253), .B2(n13263), .A(n13252), .ZN(P3_U3438) );
  MUX2_X1 U15457 ( .A(n13255), .B(n13254), .S(n15613), .Z(n13256) );
  OAI21_X1 U15458 ( .B1(n13257), .B2(n13263), .A(n13256), .ZN(P3_U3435) );
  MUX2_X1 U15459 ( .A(n13258), .B(n7968), .S(n15612), .Z(n13259) );
  OAI21_X1 U15460 ( .B1(n13263), .B2(n13260), .A(n13259), .ZN(P3_U3432) );
  MUX2_X1 U15461 ( .A(n13261), .B(n7948), .S(n15612), .Z(n13262) );
  OAI21_X1 U15462 ( .B1(n13264), .B2(n13263), .A(n13262), .ZN(P3_U3429) );
  MUX2_X1 U15463 ( .A(n13265), .B(P3_D_REG_1__SCAN_IN), .S(n13266), .Z(
        P3_U3377) );
  MUX2_X1 U15464 ( .A(n9319), .B(P3_D_REG_0__SCAN_IN), .S(n13266), .Z(P3_U3376) );
  NAND3_X1 U15465 ( .A1(n13268), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U15466 ( .A1(n13269), .A2(n14835), .ZN(n13271) );
  NAND2_X1 U15467 ( .A1(n14834), .A2(SI_31_), .ZN(n13270) );
  OAI211_X1 U15468 ( .C1(n13267), .C2(n13272), .A(n13271), .B(n13270), .ZN(
        P3_U3264) );
  AOI222_X1 U15469 ( .A1(n13274), .A2(n14835), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6755), .C1(SI_29_), .C2(n14834), .ZN(n13275) );
  INV_X1 U15470 ( .A(n13275), .ZN(P3_U3266) );
  INV_X1 U15471 ( .A(n13276), .ZN(n13278) );
  OAI222_X1 U15472 ( .A1(n13279), .A2(P3_U3151), .B1(n13282), .B2(n13278), 
        .C1(n13277), .C2(n13284), .ZN(P3_U3268) );
  INV_X1 U15473 ( .A(SI_26_), .ZN(n13283) );
  INV_X1 U15474 ( .A(n13280), .ZN(n13281) );
  OAI222_X1 U15475 ( .A1(n13285), .A2(P3_U3151), .B1(n13284), .B2(n13283), 
        .C1(n13282), .C2(n13281), .ZN(P3_U3269) );
  AOI222_X1 U15476 ( .A1(n13286), .A2(n14835), .B1(n8198), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_25_), .C2(n14834), .ZN(n13287) );
  INV_X1 U15477 ( .A(n13287), .ZN(P3_U3270) );
  NAND2_X1 U15478 ( .A1(n13633), .A2(n13318), .ZN(n13341) );
  XNOR2_X1 U15479 ( .A(n13913), .B(n13384), .ZN(n13344) );
  NAND2_X1 U15480 ( .A1(n13289), .A2(n13288), .ZN(n13294) );
  INV_X1 U15481 ( .A(n13290), .ZN(n13291) );
  OR2_X1 U15482 ( .A1(n13292), .A2(n13291), .ZN(n13293) );
  XNOR2_X1 U15483 ( .A(n13967), .B(n13336), .ZN(n13295) );
  NAND2_X1 U15484 ( .A1(n13505), .A2(n13318), .ZN(n13296) );
  NAND2_X1 U15485 ( .A1(n13295), .A2(n13296), .ZN(n13300) );
  INV_X1 U15486 ( .A(n13295), .ZN(n13298) );
  INV_X1 U15487 ( .A(n13296), .ZN(n13297) );
  NAND2_X1 U15488 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U15489 ( .A1(n13300), .A2(n13299), .ZN(n13419) );
  XNOR2_X1 U15490 ( .A(n13962), .B(n13336), .ZN(n13301) );
  NAND2_X1 U15491 ( .A1(n13770), .A2(n13318), .ZN(n13302) );
  NAND2_X1 U15492 ( .A1(n13301), .A2(n13302), .ZN(n13306) );
  INV_X1 U15493 ( .A(n13301), .ZN(n13304) );
  INV_X1 U15494 ( .A(n13302), .ZN(n13303) );
  NAND2_X1 U15495 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  AND2_X1 U15496 ( .A1(n13306), .A2(n13305), .ZN(n13429) );
  XNOR2_X1 U15497 ( .A(n13957), .B(n13336), .ZN(n13307) );
  NAND2_X1 U15498 ( .A1(n13504), .A2(n13318), .ZN(n13308) );
  XNOR2_X1 U15499 ( .A(n13307), .B(n13308), .ZN(n13473) );
  INV_X1 U15500 ( .A(n13307), .ZN(n13310) );
  INV_X1 U15501 ( .A(n13308), .ZN(n13309) );
  NAND2_X1 U15502 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  XNOR2_X1 U15503 ( .A(n13951), .B(n13384), .ZN(n13371) );
  NAND2_X1 U15504 ( .A1(n13448), .A2(n13371), .ZN(n13312) );
  AND2_X1 U15505 ( .A1(n13503), .A2(n13318), .ZN(n13372) );
  NAND2_X1 U15506 ( .A1(n13371), .A2(n13372), .ZN(n13370) );
  NAND2_X1 U15507 ( .A1(n13448), .A2(n13372), .ZN(n13313) );
  XNOR2_X1 U15508 ( .A(n13948), .B(n13384), .ZN(n13314) );
  NAND2_X1 U15509 ( .A1(n13502), .A2(n13318), .ZN(n13315) );
  XNOR2_X1 U15510 ( .A(n13314), .B(n13315), .ZN(n13459) );
  INV_X1 U15511 ( .A(n13314), .ZN(n13316) );
  NAND2_X1 U15512 ( .A1(n13316), .A2(n13315), .ZN(n13317) );
  XNOR2_X1 U15513 ( .A(n13943), .B(n13384), .ZN(n13321) );
  NAND2_X1 U15514 ( .A1(n13501), .A2(n13318), .ZN(n13319) );
  XNOR2_X1 U15515 ( .A(n13321), .B(n13319), .ZN(n13393) );
  INV_X1 U15516 ( .A(n13319), .ZN(n13320) );
  NAND2_X1 U15517 ( .A1(n13321), .A2(n13320), .ZN(n13322) );
  XNOR2_X1 U15518 ( .A(n13937), .B(n13336), .ZN(n13324) );
  XNOR2_X1 U15519 ( .A(n13326), .B(n13324), .ZN(n13463) );
  AND2_X1 U15520 ( .A1(n13461), .A2(n13318), .ZN(n13323) );
  NAND2_X1 U15521 ( .A1(n13463), .A2(n13323), .ZN(n13464) );
  INV_X1 U15522 ( .A(n13324), .ZN(n13325) );
  NAND2_X1 U15523 ( .A1(n13326), .A2(n13325), .ZN(n13327) );
  XNOR2_X1 U15524 ( .A(n13673), .B(n13336), .ZN(n13328) );
  NAND2_X1 U15525 ( .A1(n13466), .A2(n13331), .ZN(n13359) );
  INV_X1 U15526 ( .A(n13328), .ZN(n13329) );
  OR2_X1 U15527 ( .A1(n13330), .A2(n13329), .ZN(n13399) );
  XNOR2_X1 U15528 ( .A(n13920), .B(n13384), .ZN(n13332) );
  AND2_X1 U15529 ( .A1(n13500), .A2(n13331), .ZN(n13333) );
  NAND2_X1 U15530 ( .A1(n13332), .A2(n13333), .ZN(n13342) );
  INV_X1 U15531 ( .A(n13332), .ZN(n13485) );
  INV_X1 U15532 ( .A(n13333), .ZN(n13334) );
  NAND2_X1 U15533 ( .A1(n13485), .A2(n13334), .ZN(n13335) );
  NAND2_X1 U15534 ( .A1(n13342), .A2(n13335), .ZN(n13404) );
  XNOR2_X1 U15535 ( .A(n13925), .B(n13336), .ZN(n13405) );
  NAND2_X1 U15536 ( .A1(n13632), .A2(n13318), .ZN(n13338) );
  AND2_X1 U15537 ( .A1(n13405), .A2(n13338), .ZN(n13402) );
  NOR2_X1 U15538 ( .A1(n13404), .A2(n13402), .ZN(n13337) );
  INV_X1 U15539 ( .A(n13405), .ZN(n13340) );
  INV_X1 U15540 ( .A(n13338), .ZN(n13339) );
  NAND2_X1 U15541 ( .A1(n13340), .A2(n13339), .ZN(n13401) );
  XNOR2_X1 U15542 ( .A(n13344), .B(n13341), .ZN(n13494) );
  AND2_X1 U15543 ( .A1(n13494), .A2(n13342), .ZN(n13343) );
  XNOR2_X1 U15544 ( .A(n13905), .B(n13384), .ZN(n13346) );
  AND2_X1 U15545 ( .A1(n13499), .A2(n13331), .ZN(n13345) );
  NAND2_X1 U15546 ( .A1(n13346), .A2(n13345), .ZN(n13380) );
  OAI21_X1 U15547 ( .B1(n13346), .B2(n13345), .A(n13380), .ZN(n13347) );
  NOR2_X1 U15548 ( .A1(n13348), .A2(n13347), .ZN(n13382) );
  AND2_X1 U15549 ( .A1(n13633), .A2(n13854), .ZN(n13349) );
  AOI21_X1 U15550 ( .B1(n13498), .B2(n13851), .A(n13349), .ZN(n13601) );
  INV_X1 U15551 ( .A(n13604), .ZN(n13350) );
  AOI22_X1 U15552 ( .A1(n13350), .A2(n13488), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13351) );
  OAI21_X1 U15553 ( .B1(n13601), .B2(n15216), .A(n13351), .ZN(n13352) );
  INV_X1 U15554 ( .A(n13352), .ZN(n13353) );
  INV_X1 U15555 ( .A(n13358), .ZN(P2_U3186) );
  NAND2_X1 U15556 ( .A1(n13466), .A2(n13462), .ZN(n13362) );
  NAND2_X1 U15557 ( .A1(n13359), .A2(n13492), .ZN(n13361) );
  MUX2_X1 U15558 ( .A(n13362), .B(n13361), .S(n13360), .Z(n13369) );
  NAND2_X1 U15559 ( .A1(n13632), .A2(n13851), .ZN(n13364) );
  NAND2_X1 U15560 ( .A1(n13461), .A2(n13854), .ZN(n13363) );
  NAND2_X1 U15561 ( .A1(n13364), .A2(n13363), .ZN(n13663) );
  INV_X1 U15562 ( .A(n13666), .ZN(n13366) );
  OAI22_X1 U15563 ( .A1(n13366), .A2(n15226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13365), .ZN(n13367) );
  AOI21_X1 U15564 ( .B1(n13663), .B2(n13476), .A(n13367), .ZN(n13368) );
  OAI211_X1 U15565 ( .C1(n8920), .C2(n13447), .A(n13369), .B(n13368), .ZN(
        P2_U3188) );
  OAI21_X1 U15566 ( .B1(n13372), .B2(n13371), .A(n13370), .ZN(n13373) );
  XOR2_X1 U15567 ( .A(n13373), .B(n13448), .Z(n13379) );
  OAI22_X1 U15568 ( .A1(n13375), .A2(n13872), .B1(n13374), .B2(n13874), .ZN(
        n13727) );
  NAND2_X1 U15569 ( .A1(n13727), .A2(n13476), .ZN(n13376) );
  NAND2_X1 U15570 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13568)
         );
  OAI211_X1 U15571 ( .C1(n15226), .C2(n13734), .A(n13376), .B(n13568), .ZN(
        n13377) );
  AOI21_X1 U15572 ( .B1(n13951), .B2(n15223), .A(n13377), .ZN(n13378) );
  OAI21_X1 U15573 ( .B1(n13379), .B2(n13480), .A(n13378), .ZN(P2_U3191) );
  INV_X1 U15574 ( .A(n13380), .ZN(n13381) );
  NAND2_X1 U15575 ( .A1(n13498), .A2(n13331), .ZN(n13383) );
  XOR2_X1 U15576 ( .A(n13384), .B(n13383), .Z(n13385) );
  XNOR2_X1 U15577 ( .A(n13899), .B(n13385), .ZN(n13386) );
  XNOR2_X1 U15578 ( .A(n13387), .B(n13386), .ZN(n13391) );
  AOI22_X1 U15579 ( .A1(n13497), .A2(n13851), .B1(n13499), .B2(n13854), .ZN(
        n13586) );
  AOI22_X1 U15580 ( .A1(n13593), .A2(n13488), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13388) );
  OAI21_X1 U15581 ( .B1(n13586), .B2(n15216), .A(n13388), .ZN(n13389) );
  AOI21_X1 U15582 ( .B1(n13899), .B2(n15223), .A(n13389), .ZN(n13390) );
  OAI21_X1 U15583 ( .B1(n13391), .B2(n13480), .A(n13390), .ZN(P2_U3192) );
  OAI211_X1 U15584 ( .C1(n13394), .C2(n13393), .A(n13392), .B(n13492), .ZN(
        n13398) );
  AOI22_X1 U15585 ( .A1(n13461), .A2(n13851), .B1(n13854), .B2(n13502), .ZN(
        n13697) );
  OAI22_X1 U15586 ( .A1(n13697), .A2(n15216), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13395), .ZN(n13396) );
  AOI21_X1 U15587 ( .B1(n13701), .B2(n13488), .A(n13396), .ZN(n13397) );
  OAI211_X1 U15588 ( .C1(n7034), .C2(n13447), .A(n13398), .B(n13397), .ZN(
        P2_U3195) );
  AND2_X1 U15589 ( .A1(n13400), .A2(n13399), .ZN(n13440) );
  INV_X1 U15590 ( .A(n13401), .ZN(n13403) );
  NOR2_X1 U15591 ( .A1(n13403), .A2(n13402), .ZN(n13439) );
  NAND2_X1 U15592 ( .A1(n13440), .A2(n13439), .ZN(n13438) );
  AOI21_X1 U15593 ( .B1(n13438), .B2(n13404), .A(n13480), .ZN(n13407) );
  NOR3_X1 U15594 ( .A1(n13405), .A2(n13410), .A3(n13483), .ZN(n13406) );
  OAI21_X1 U15595 ( .B1(n13407), .B2(n13406), .A(n13482), .ZN(n13415) );
  OAI22_X1 U15596 ( .A1(n13410), .A2(n13409), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13408), .ZN(n13413) );
  NOR2_X1 U15597 ( .A1(n13411), .A2(n13421), .ZN(n13412) );
  AOI211_X1 U15598 ( .C1(n13488), .C2(n13638), .A(n13413), .B(n13412), .ZN(
        n13414) );
  OAI211_X1 U15599 ( .C1(n13641), .C2(n13447), .A(n13415), .B(n13414), .ZN(
        P2_U3197) );
  INV_X1 U15600 ( .A(n13416), .ZN(n13417) );
  AOI21_X1 U15601 ( .B1(n13419), .B2(n6782), .A(n13417), .ZN(n13426) );
  OAI21_X1 U15602 ( .B1(n13475), .B2(n13421), .A(n13420), .ZN(n13422) );
  AOI21_X1 U15603 ( .B1(n13452), .B2(n13784), .A(n13422), .ZN(n13423) );
  OAI21_X1 U15604 ( .B1(n13776), .B2(n15226), .A(n13423), .ZN(n13424) );
  AOI21_X1 U15605 ( .B1(n13967), .B2(n15223), .A(n13424), .ZN(n13425) );
  OAI21_X1 U15606 ( .B1(n13426), .B2(n13480), .A(n13425), .ZN(P2_U3198) );
  OAI21_X1 U15607 ( .B1(n13429), .B2(n13428), .A(n13427), .ZN(n13430) );
  NAND2_X1 U15608 ( .A1(n13430), .A2(n13492), .ZN(n13437) );
  NAND2_X1 U15609 ( .A1(n13504), .A2(n13851), .ZN(n13432) );
  NAND2_X1 U15610 ( .A1(n13505), .A2(n13854), .ZN(n13431) );
  NAND2_X1 U15611 ( .A1(n13432), .A2(n13431), .ZN(n13752) );
  INV_X1 U15612 ( .A(n13433), .ZN(n13435) );
  NOR2_X1 U15613 ( .A1(n15226), .A2(n13756), .ZN(n13434) );
  AOI211_X1 U15614 ( .C1(n13476), .C2(n13752), .A(n13435), .B(n13434), .ZN(
        n13436) );
  OAI211_X1 U15615 ( .C1(n7048), .C2(n13447), .A(n13437), .B(n13436), .ZN(
        P2_U3200) );
  INV_X1 U15616 ( .A(n13925), .ZN(n13654) );
  OAI211_X1 U15617 ( .C1(n13440), .C2(n13439), .A(n13438), .B(n13492), .ZN(
        n13446) );
  NAND2_X1 U15618 ( .A1(n13500), .A2(n13851), .ZN(n13442) );
  NAND2_X1 U15619 ( .A1(n13466), .A2(n13854), .ZN(n13441) );
  NAND2_X1 U15620 ( .A1(n13442), .A2(n13441), .ZN(n13648) );
  OAI22_X1 U15621 ( .A1(n13645), .A2(n15226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13443), .ZN(n13444) );
  AOI21_X1 U15622 ( .B1(n13648), .B2(n13476), .A(n13444), .ZN(n13445) );
  OAI211_X1 U15623 ( .C1(n13654), .C2(n13447), .A(n13446), .B(n13445), .ZN(
        P2_U3201) );
  NOR2_X1 U15624 ( .A1(n13713), .A2(n13483), .ZN(n13449) );
  AOI22_X1 U15625 ( .A1(n13450), .A2(n13492), .B1(n13449), .B2(n13448), .ZN(
        n13460) );
  NAND2_X1 U15626 ( .A1(n13501), .A2(n13451), .ZN(n13454) );
  AOI22_X1 U15627 ( .A1(n13452), .A2(n13503), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13453) );
  OAI211_X1 U15628 ( .C1(n15226), .C2(n13717), .A(n13454), .B(n13453), .ZN(
        n13457) );
  NOR2_X1 U15629 ( .A1(n13455), .A2(n13480), .ZN(n13456) );
  AOI211_X1 U15630 ( .C1(n13948), .C2(n15223), .A(n13457), .B(n13456), .ZN(
        n13458) );
  OAI21_X1 U15631 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(P2_U3205) );
  AOI22_X1 U15632 ( .A1(n13463), .A2(n13492), .B1(n13462), .B2(n13461), .ZN(
        n13472) );
  INV_X1 U15633 ( .A(n13464), .ZN(n13471) );
  AND2_X1 U15634 ( .A1(n13501), .A2(n13854), .ZN(n13465) );
  AOI21_X1 U15635 ( .B1(n13466), .B2(n13851), .A(n13465), .ZN(n13681) );
  INV_X1 U15636 ( .A(n13467), .ZN(n13687) );
  AOI22_X1 U15637 ( .A1(n13488), .A2(n13687), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13468) );
  OAI21_X1 U15638 ( .B1(n13681), .B2(n15216), .A(n13468), .ZN(n13469) );
  AOI21_X1 U15639 ( .B1(n13937), .B2(n15223), .A(n13469), .ZN(n13470) );
  OAI21_X1 U15640 ( .B1(n13472), .B2(n13471), .A(n13470), .ZN(P2_U3207) );
  XNOR2_X1 U15641 ( .A(n13474), .B(n13473), .ZN(n13481) );
  OAI22_X1 U15642 ( .A1(n13713), .A2(n13872), .B1(n13475), .B2(n13874), .ZN(
        n13739) );
  AOI22_X1 U15643 ( .A1(n13739), .A2(n13476), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13477) );
  OAI21_X1 U15644 ( .B1(n13742), .B2(n15226), .A(n13477), .ZN(n13478) );
  AOI21_X1 U15645 ( .B1(n13957), .B2(n15223), .A(n13478), .ZN(n13479) );
  OAI21_X1 U15646 ( .B1(n13481), .B2(n13480), .A(n13479), .ZN(P2_U3210) );
  INV_X1 U15647 ( .A(n13482), .ZN(n13487) );
  NOR3_X1 U15648 ( .A1(n13485), .A2(n13484), .A3(n13483), .ZN(n13486) );
  AOI21_X1 U15649 ( .B1(n13487), .B2(n13492), .A(n13486), .ZN(n13495) );
  AOI22_X1 U15650 ( .A1(n13499), .A2(n13851), .B1(n13854), .B2(n13500), .ZN(
        n13615) );
  NAND2_X1 U15651 ( .A1(n13913), .A2(n15223), .ZN(n13490) );
  AOI22_X1 U15652 ( .A1(n13622), .A2(n13488), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13489) );
  OAI211_X1 U15653 ( .C1(n13615), .C2(n15216), .A(n13490), .B(n13489), .ZN(
        n13491) );
  AOI21_X1 U15654 ( .B1(n6649), .B2(n13492), .A(n13491), .ZN(n13493) );
  OAI21_X1 U15655 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(P2_U3212) );
  CLKBUF_X1 U15656 ( .A(n13507), .Z(n13516) );
  MUX2_X1 U15657 ( .A(n13496), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13516), .Z(
        P2_U3561) );
  MUX2_X1 U15658 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13497), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15659 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13498), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15660 ( .A(n13499), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13507), .Z(
        P2_U3558) );
  MUX2_X1 U15661 ( .A(n13633), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13507), .Z(
        P2_U3557) );
  MUX2_X1 U15662 ( .A(n13500), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13516), .Z(
        P2_U3556) );
  MUX2_X1 U15663 ( .A(n13632), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13516), .Z(
        P2_U3555) );
  MUX2_X1 U15664 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13501), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15665 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13502), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15666 ( .A(n13503), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13507), .Z(
        P2_U3550) );
  MUX2_X1 U15667 ( .A(n13504), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13507), .Z(
        P2_U3549) );
  MUX2_X1 U15668 ( .A(n13770), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13516), .Z(
        P2_U3548) );
  MUX2_X1 U15669 ( .A(n13505), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13516), .Z(
        P2_U3547) );
  MUX2_X1 U15670 ( .A(n13784), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13507), .Z(
        P2_U3546) );
  MUX2_X1 U15671 ( .A(n13506), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13507), .Z(
        P2_U3545) );
  MUX2_X1 U15672 ( .A(n13797), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13516), .Z(
        P2_U3544) );
  MUX2_X1 U15673 ( .A(n13814), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13516), .Z(
        P2_U3543) );
  MUX2_X1 U15674 ( .A(n13798), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13507), .Z(
        P2_U3542) );
  MUX2_X1 U15675 ( .A(n13852), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13507), .Z(
        P2_U3541) );
  MUX2_X1 U15676 ( .A(n13508), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13516), .Z(
        P2_U3540) );
  MUX2_X1 U15677 ( .A(n13853), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13516), .Z(
        P2_U3539) );
  MUX2_X1 U15678 ( .A(n13509), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13516), .Z(
        P2_U3538) );
  MUX2_X1 U15679 ( .A(n13510), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13516), .Z(
        P2_U3537) );
  MUX2_X1 U15680 ( .A(n13511), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13516), .Z(
        P2_U3536) );
  MUX2_X1 U15681 ( .A(n13512), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13516), .Z(
        P2_U3535) );
  MUX2_X1 U15682 ( .A(n13513), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13516), .Z(
        P2_U3534) );
  MUX2_X1 U15683 ( .A(n13514), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13516), .Z(
        P2_U3533) );
  MUX2_X1 U15684 ( .A(n13515), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13516), .Z(
        P2_U3532) );
  MUX2_X1 U15685 ( .A(n8959), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13516), .Z(
        P2_U3531) );
  NOR2_X1 U15686 ( .A1(n13518), .A2(n13517), .ZN(n13520) );
  OAI21_X1 U15687 ( .B1(n13520), .B2(n13519), .A(n15302), .ZN(n13532) );
  INV_X1 U15688 ( .A(n13521), .ZN(n13524) );
  NOR2_X1 U15689 ( .A1(n15290), .A2(n13522), .ZN(n13523) );
  AOI211_X1 U15690 ( .C1(n15298), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n13524), 
        .B(n13523), .ZN(n13531) );
  OR3_X1 U15691 ( .A1(n13527), .A2(n13526), .A3(n13525), .ZN(n13528) );
  NAND3_X1 U15692 ( .A1(n13529), .A2(n15305), .A3(n13528), .ZN(n13530) );
  NAND3_X1 U15693 ( .A1(n13532), .A2(n13531), .A3(n13530), .ZN(P2_U3225) );
  NAND2_X1 U15694 ( .A1(n13533), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13534) );
  NOR2_X1 U15695 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13537), .ZN(n13551) );
  AOI21_X1 U15696 ( .B1(n13537), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13551), 
        .ZN(n13549) );
  NOR2_X1 U15697 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13538), .ZN(n13541) );
  NOR2_X1 U15698 ( .A1(n15290), .A2(n13539), .ZN(n13540) );
  AOI211_X1 U15699 ( .C1(n15298), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13541), 
        .B(n13540), .ZN(n13548) );
  OAI22_X1 U15700 ( .A1(n13545), .A2(n13544), .B1(n13543), .B2(n13542), .ZN(
        n13556) );
  XNOR2_X1 U15701 ( .A(n13556), .B(n13555), .ZN(n13553) );
  XNOR2_X1 U15702 ( .A(n13553), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U15703 ( .A1(n13546), .A2(n15305), .ZN(n13547) );
  OAI211_X1 U15704 ( .C1(n13549), .C2(n15263), .A(n13548), .B(n13547), .ZN(
        P2_U3232) );
  NAND2_X1 U15705 ( .A1(n13564), .A2(n15302), .ZN(n13562) );
  INV_X1 U15706 ( .A(n13553), .ZN(n13554) );
  NAND2_X1 U15707 ( .A1(n13554), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U15708 ( .A1(n13556), .A2(n13555), .ZN(n13557) );
  NAND2_X1 U15709 ( .A1(n13558), .A2(n13557), .ZN(n13560) );
  XOR2_X1 U15710 ( .A(n13560), .B(n13559), .Z(n13563) );
  AOI21_X1 U15711 ( .B1(n13563), .B2(n15305), .A(n15300), .ZN(n13561) );
  NAND2_X1 U15712 ( .A1(n13562), .A2(n13561), .ZN(n13567) );
  OAI22_X1 U15713 ( .A1(n13564), .A2(n15263), .B1(n13563), .B2(n15265), .ZN(
        n13566) );
  OAI21_X1 U15714 ( .B1(n15297), .B2(n7722), .A(n13568), .ZN(n13569) );
  NAND2_X1 U15715 ( .A1(n13897), .A2(n13579), .ZN(n13578) );
  XOR2_X1 U15716 ( .A(n13575), .B(n13578), .Z(n13572) );
  NAND2_X1 U15717 ( .A1(n13572), .A2(n15323), .ZN(n13893) );
  NAND2_X1 U15718 ( .A1(n13574), .A2(n13573), .ZN(n13895) );
  NOR2_X1 U15719 ( .A1(n15316), .A2(n13895), .ZN(n13581) );
  INV_X1 U15720 ( .A(n13575), .ZN(n13894) );
  NOR2_X1 U15721 ( .A1(n13894), .A2(n14957), .ZN(n13576) );
  AOI211_X1 U15722 ( .C1(n15316), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13581), 
        .B(n13576), .ZN(n13577) );
  OAI21_X1 U15723 ( .B1(n13893), .B2(n13886), .A(n13577), .ZN(P2_U3234) );
  OAI211_X1 U15724 ( .C1(n13897), .C2(n13579), .A(n15323), .B(n13578), .ZN(
        n13896) );
  NOR2_X1 U15725 ( .A1(n13897), .A2(n14957), .ZN(n13580) );
  AOI211_X1 U15726 ( .C1(n15316), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13581), 
        .B(n13580), .ZN(n13582) );
  OAI21_X1 U15727 ( .B1(n13886), .B2(n13896), .A(n13582), .ZN(P2_U3235) );
  OAI211_X1 U15728 ( .C1(n13585), .C2(n13584), .A(n13583), .B(n15313), .ZN(
        n13587) );
  AND2_X2 U15729 ( .A1(n13587), .A2(n13586), .ZN(n13901) );
  OAI21_X1 U15730 ( .B1(n13590), .B2(n13589), .A(n13588), .ZN(n13902) );
  INV_X1 U15731 ( .A(n13902), .ZN(n13597) );
  AOI21_X1 U15732 ( .B1(n6640), .B2(n13899), .A(n13979), .ZN(n13592) );
  AND2_X1 U15733 ( .A1(n13592), .A2(n13591), .ZN(n13898) );
  NAND2_X1 U15734 ( .A1(n13898), .A2(n15326), .ZN(n13595) );
  AOI22_X1 U15735 ( .A1(n13593), .A2(n15315), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15316), .ZN(n13594) );
  OAI211_X1 U15736 ( .C1(n6774), .C2(n14957), .A(n13595), .B(n13594), .ZN(
        n13596) );
  AOI21_X1 U15737 ( .B1(n13597), .B2(n15327), .A(n13596), .ZN(n13598) );
  OAI21_X1 U15738 ( .B1(n13901), .B2(n15316), .A(n13598), .ZN(P2_U3237) );
  XNOR2_X1 U15739 ( .A(n13599), .B(n13608), .ZN(n13600) );
  NAND2_X1 U15740 ( .A1(n13600), .A2(n15313), .ZN(n13602) );
  NAND2_X1 U15741 ( .A1(n13602), .A2(n13601), .ZN(n13910) );
  INV_X1 U15742 ( .A(n13910), .ZN(n13612) );
  OAI22_X1 U15743 ( .A1(n13604), .A2(n13880), .B1(n13603), .B2(n13883), .ZN(
        n13607) );
  OAI211_X1 U15744 ( .C1(n13605), .C2(n13621), .A(n15323), .B(n6640), .ZN(
        n13906) );
  NOR2_X1 U15745 ( .A1(n13906), .A2(n13886), .ZN(n13606) );
  AOI211_X1 U15746 ( .C1(n15317), .C2(n13905), .A(n13607), .B(n13606), .ZN(
        n13611) );
  NAND2_X1 U15747 ( .A1(n13609), .A2(n13608), .ZN(n13903) );
  NAND3_X1 U15748 ( .A1(n13904), .A2(n13903), .A3(n15327), .ZN(n13610) );
  OAI211_X1 U15749 ( .C1(n15316), .C2(n13612), .A(n13611), .B(n13610), .ZN(
        P2_U3238) );
  XNOR2_X1 U15750 ( .A(n13613), .B(n13617), .ZN(n13614) );
  NAND2_X1 U15751 ( .A1(n13614), .A2(n15313), .ZN(n13616) );
  NAND2_X1 U15752 ( .A1(n13616), .A2(n13615), .ZN(n13918) );
  INV_X1 U15753 ( .A(n13918), .ZN(n13627) );
  XNOR2_X1 U15754 ( .A(n13618), .B(n13617), .ZN(n13914) );
  NAND2_X1 U15755 ( .A1(n13913), .A2(n13636), .ZN(n13619) );
  NAND2_X1 U15756 ( .A1(n13619), .A2(n15323), .ZN(n13620) );
  OR2_X1 U15757 ( .A1(n13621), .A2(n13620), .ZN(n13915) );
  AOI22_X1 U15758 ( .A1(n13622), .A2(n15315), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15316), .ZN(n13624) );
  NAND2_X1 U15759 ( .A1(n13913), .A2(n15317), .ZN(n13623) );
  OAI211_X1 U15760 ( .C1(n13915), .C2(n13886), .A(n13624), .B(n13623), .ZN(
        n13625) );
  AOI21_X1 U15761 ( .B1(n13914), .B2(n15327), .A(n13625), .ZN(n13626) );
  OAI21_X1 U15762 ( .B1(n13627), .B2(n15316), .A(n13626), .ZN(P2_U3239) );
  XOR2_X1 U15763 ( .A(n13630), .B(n13628), .Z(n13923) );
  OAI21_X1 U15764 ( .B1(n13631), .B2(n13630), .A(n13629), .ZN(n13634) );
  AOI222_X1 U15765 ( .A1(n15313), .A2(n13634), .B1(n13633), .B2(n13851), .C1(
        n13632), .C2(n13854), .ZN(n13922) );
  INV_X1 U15766 ( .A(n13922), .ZN(n13643) );
  INV_X1 U15767 ( .A(n13652), .ZN(n13635) );
  AOI21_X1 U15768 ( .B1(n13635), .B2(n13920), .A(n13979), .ZN(n13637) );
  AND2_X1 U15769 ( .A1(n13637), .A2(n13636), .ZN(n13919) );
  NAND2_X1 U15770 ( .A1(n13919), .A2(n15326), .ZN(n13640) );
  AOI22_X1 U15771 ( .A1(n13638), .A2(n15315), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15316), .ZN(n13639) );
  OAI211_X1 U15772 ( .C1(n13641), .C2(n14957), .A(n13640), .B(n13639), .ZN(
        n13642) );
  AOI21_X1 U15773 ( .B1(n13643), .B2(n13883), .A(n13642), .ZN(n13644) );
  OAI21_X1 U15774 ( .B1(n13923), .B2(n14959), .A(n13644), .ZN(P2_U3240) );
  INV_X1 U15775 ( .A(n13645), .ZN(n13651) );
  XNOR2_X1 U15776 ( .A(n13647), .B(n13646), .ZN(n13649) );
  AOI21_X1 U15777 ( .B1(n13649), .B2(n15313), .A(n13648), .ZN(n13929) );
  INV_X1 U15778 ( .A(n13929), .ZN(n13650) );
  AOI21_X1 U15779 ( .B1(n13651), .B2(n15315), .A(n13650), .ZN(n13660) );
  AOI211_X1 U15780 ( .C1(n13925), .C2(n13671), .A(n13979), .B(n13652), .ZN(
        n13924) );
  OAI22_X1 U15781 ( .A1(n13654), .A2(n14957), .B1(n13883), .B2(n13653), .ZN(
        n13655) );
  AOI21_X1 U15782 ( .B1(n13924), .B2(n15326), .A(n13655), .ZN(n13659) );
  NAND2_X1 U15783 ( .A1(n13657), .A2(n13656), .ZN(n13926) );
  NAND3_X1 U15784 ( .A1(n13926), .A2(n13927), .A3(n15327), .ZN(n13658) );
  OAI211_X1 U15785 ( .C1(n13660), .C2(n15316), .A(n13659), .B(n13658), .ZN(
        P2_U3241) );
  XNOR2_X1 U15786 ( .A(n13661), .B(n13667), .ZN(n13662) );
  NAND2_X1 U15787 ( .A1(n13662), .A2(n15313), .ZN(n13665) );
  INV_X1 U15788 ( .A(n13663), .ZN(n13664) );
  NAND2_X1 U15789 ( .A1(n13665), .A2(n13664), .ZN(n13935) );
  AOI21_X1 U15790 ( .B1(n13666), .B2(n15315), .A(n13935), .ZN(n13677) );
  INV_X1 U15791 ( .A(n13667), .ZN(n13668) );
  XNOR2_X1 U15792 ( .A(n13669), .B(n13668), .ZN(n13931) );
  INV_X1 U15793 ( .A(n13670), .ZN(n13685) );
  AOI21_X1 U15794 ( .B1(n13673), .B2(n13685), .A(n13979), .ZN(n13672) );
  NAND2_X1 U15795 ( .A1(n13672), .A2(n13671), .ZN(n13932) );
  AOI22_X1 U15796 ( .A1(n13673), .A2(n15317), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n15316), .ZN(n13674) );
  OAI21_X1 U15797 ( .B1(n13932), .B2(n13886), .A(n13674), .ZN(n13675) );
  AOI21_X1 U15798 ( .B1(n13931), .B2(n15327), .A(n13675), .ZN(n13676) );
  OAI21_X1 U15799 ( .B1(n13677), .B2(n15316), .A(n13676), .ZN(P2_U3242) );
  XNOR2_X1 U15800 ( .A(n13678), .B(n13679), .ZN(n13940) );
  AOI21_X1 U15801 ( .B1(n13680), .B2(n13679), .A(n13712), .ZN(n13684) );
  INV_X1 U15802 ( .A(n13681), .ZN(n13682) );
  AOI21_X1 U15803 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13939) );
  INV_X1 U15804 ( .A(n13939), .ZN(n13692) );
  INV_X1 U15805 ( .A(n13937), .ZN(n13690) );
  AOI21_X1 U15806 ( .B1(n13937), .B2(n13699), .A(n13979), .ZN(n13686) );
  AND2_X1 U15807 ( .A1(n13686), .A2(n13685), .ZN(n13936) );
  NAND2_X1 U15808 ( .A1(n13936), .A2(n15326), .ZN(n13689) );
  AOI22_X1 U15809 ( .A1(n13687), .A2(n15315), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n15316), .ZN(n13688) );
  OAI211_X1 U15810 ( .C1(n13690), .C2(n14957), .A(n13689), .B(n13688), .ZN(
        n13691) );
  AOI21_X1 U15811 ( .B1(n13692), .B2(n13883), .A(n13691), .ZN(n13693) );
  OAI21_X1 U15812 ( .B1(n14959), .B2(n13940), .A(n13693), .ZN(P2_U3243) );
  XOR2_X1 U15813 ( .A(n13695), .B(n13694), .Z(n13945) );
  XNOR2_X1 U15814 ( .A(n13696), .B(n13695), .ZN(n13698) );
  OAI21_X1 U15815 ( .B1(n13698), .B2(n13712), .A(n13697), .ZN(n13941) );
  AOI21_X1 U15816 ( .B1(n13943), .B2(n13715), .A(n13979), .ZN(n13700) );
  AND2_X1 U15817 ( .A1(n13700), .A2(n13699), .ZN(n13942) );
  NAND2_X1 U15818 ( .A1(n13942), .A2(n15326), .ZN(n13703) );
  AOI22_X1 U15819 ( .A1(n13701), .A2(n15315), .B1(n15316), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13702) );
  OAI211_X1 U15820 ( .C1(n7034), .C2(n14957), .A(n13703), .B(n13702), .ZN(
        n13704) );
  AOI21_X1 U15821 ( .B1(n13941), .B2(n13883), .A(n13704), .ZN(n13705) );
  OAI21_X1 U15822 ( .B1(n14959), .B2(n13945), .A(n13705), .ZN(P2_U3244) );
  XNOR2_X1 U15823 ( .A(n13706), .B(n13710), .ZN(n13950) );
  INV_X1 U15824 ( .A(n13707), .ZN(n13708) );
  AOI21_X1 U15825 ( .B1(n13710), .B2(n13709), .A(n13708), .ZN(n13711) );
  OAI222_X1 U15826 ( .A1(n13872), .A2(n13714), .B1(n13874), .B2(n13713), .C1(
        n13712), .C2(n13711), .ZN(n13946) );
  INV_X1 U15827 ( .A(n13948), .ZN(n13721) );
  AOI21_X1 U15828 ( .B1(n13730), .B2(n13948), .A(n13979), .ZN(n13716) );
  AND2_X1 U15829 ( .A1(n13716), .A2(n13715), .ZN(n13947) );
  NAND2_X1 U15830 ( .A1(n13947), .A2(n15326), .ZN(n13720) );
  INV_X1 U15831 ( .A(n13717), .ZN(n13718) );
  AOI22_X1 U15832 ( .A1(n15316), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n15315), 
        .B2(n13718), .ZN(n13719) );
  OAI211_X1 U15833 ( .C1(n13721), .C2(n14957), .A(n13720), .B(n13719), .ZN(
        n13722) );
  AOI21_X1 U15834 ( .B1(n13946), .B2(n13883), .A(n13722), .ZN(n13723) );
  OAI21_X1 U15835 ( .B1(n14959), .B2(n13950), .A(n13723), .ZN(P2_U3245) );
  XOR2_X1 U15836 ( .A(n13724), .B(n13725), .Z(n13955) );
  XOR2_X1 U15837 ( .A(n13726), .B(n13725), .Z(n13728) );
  AOI21_X1 U15838 ( .B1(n13728), .B2(n15313), .A(n13727), .ZN(n13954) );
  INV_X1 U15839 ( .A(n13730), .ZN(n13731) );
  AOI21_X1 U15840 ( .B1(n13951), .B2(n13741), .A(n13731), .ZN(n13952) );
  NAND2_X1 U15841 ( .A1(n13952), .A2(n13732), .ZN(n13733) );
  OAI211_X1 U15842 ( .C1(n13880), .C2(n13734), .A(n13954), .B(n13733), .ZN(
        n13735) );
  NAND2_X1 U15843 ( .A1(n13735), .A2(n13883), .ZN(n13737) );
  AOI22_X1 U15844 ( .A1(n13951), .A2(n15317), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n15316), .ZN(n13736) );
  OAI211_X1 U15845 ( .C1(n13955), .C2(n14959), .A(n13737), .B(n13736), .ZN(
        P2_U3246) );
  XNOR2_X1 U15846 ( .A(n13738), .B(n13747), .ZN(n13740) );
  AOI21_X1 U15847 ( .B1(n13740), .B2(n15313), .A(n13739), .ZN(n13959) );
  AOI211_X1 U15848 ( .C1(n13957), .C2(n13754), .A(n13979), .B(n13729), .ZN(
        n13956) );
  INV_X1 U15849 ( .A(n13957), .ZN(n13745) );
  INV_X1 U15850 ( .A(n13742), .ZN(n13743) );
  AOI22_X1 U15851 ( .A1(n15316), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n15315), 
        .B2(n13743), .ZN(n13744) );
  OAI21_X1 U15852 ( .B1(n13745), .B2(n14957), .A(n13744), .ZN(n13749) );
  XOR2_X1 U15853 ( .A(n13747), .B(n13746), .Z(n13960) );
  NOR2_X1 U15854 ( .A1(n13960), .A2(n14959), .ZN(n13748) );
  AOI211_X1 U15855 ( .C1(n13956), .C2(n15326), .A(n13749), .B(n13748), .ZN(
        n13750) );
  OAI21_X1 U15856 ( .B1(n15316), .B2(n13959), .A(n13750), .ZN(P2_U3247) );
  XOR2_X1 U15857 ( .A(n13759), .B(n13751), .Z(n13753) );
  AOI21_X1 U15858 ( .B1(n13753), .B2(n15313), .A(n13752), .ZN(n13964) );
  INV_X1 U15859 ( .A(n13754), .ZN(n13755) );
  AOI211_X1 U15860 ( .C1(n13962), .C2(n13774), .A(n13979), .B(n13755), .ZN(
        n13961) );
  INV_X1 U15861 ( .A(n13756), .ZN(n13757) );
  AOI22_X1 U15862 ( .A1(n15316), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n15315), 
        .B2(n13757), .ZN(n13758) );
  OAI21_X1 U15863 ( .B1(n7048), .B2(n14957), .A(n13758), .ZN(n13762) );
  XNOR2_X1 U15864 ( .A(n13760), .B(n13759), .ZN(n13965) );
  NOR2_X1 U15865 ( .A1(n13965), .A2(n14959), .ZN(n13761) );
  AOI211_X1 U15866 ( .C1(n13961), .C2(n15326), .A(n13762), .B(n13761), .ZN(
        n13763) );
  OAI21_X1 U15867 ( .B1(n15316), .B2(n13964), .A(n13763), .ZN(P2_U3248) );
  XNOR2_X1 U15868 ( .A(n13765), .B(n13764), .ZN(n13773) );
  NAND2_X1 U15869 ( .A1(n13767), .A2(n13766), .ZN(n13768) );
  NAND2_X1 U15870 ( .A1(n13769), .A2(n13768), .ZN(n13970) );
  AOI22_X1 U15871 ( .A1(n13854), .A2(n13784), .B1(n13770), .B2(n13851), .ZN(
        n13771) );
  OAI21_X1 U15872 ( .B1(n13970), .B2(n6801), .A(n13771), .ZN(n13772) );
  AOI21_X1 U15873 ( .B1(n13773), .B2(n15313), .A(n13772), .ZN(n13969) );
  INV_X1 U15874 ( .A(n13774), .ZN(n13775) );
  AOI211_X1 U15875 ( .C1(n13967), .C2(n7052), .A(n13979), .B(n13775), .ZN(
        n13966) );
  INV_X1 U15876 ( .A(n13776), .ZN(n13777) );
  AOI22_X1 U15877 ( .A1(n15316), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n15315), 
        .B2(n13777), .ZN(n13778) );
  OAI21_X1 U15878 ( .B1(n13779), .B2(n14957), .A(n13778), .ZN(n13781) );
  NOR2_X1 U15879 ( .A1(n13970), .A2(n13892), .ZN(n13780) );
  AOI211_X1 U15880 ( .C1(n13966), .C2(n15326), .A(n13781), .B(n13780), .ZN(
        n13782) );
  OAI21_X1 U15881 ( .B1(n15316), .B2(n13969), .A(n13782), .ZN(P2_U3249) );
  XNOR2_X1 U15882 ( .A(n13783), .B(n13786), .ZN(n13785) );
  AOI222_X1 U15883 ( .A1(n15313), .A2(n13785), .B1(n13784), .B2(n13851), .C1(
        n13797), .C2(n13854), .ZN(n14968) );
  XNOR2_X1 U15884 ( .A(n13787), .B(n13786), .ZN(n14971) );
  OAI211_X1 U15885 ( .C1(n13788), .C2(n14967), .A(n15323), .B(n13980), .ZN(
        n14966) );
  OAI22_X1 U15886 ( .A1(n13883), .A2(n13790), .B1(n13789), .B2(n13880), .ZN(
        n13791) );
  AOI21_X1 U15887 ( .B1(n13792), .B2(n15317), .A(n13791), .ZN(n13793) );
  OAI21_X1 U15888 ( .B1(n14966), .B2(n13886), .A(n13793), .ZN(n13794) );
  AOI21_X1 U15889 ( .B1(n14971), .B2(n15327), .A(n13794), .ZN(n13795) );
  OAI21_X1 U15890 ( .B1(n14968), .B2(n15316), .A(n13795), .ZN(P2_U3251) );
  XNOR2_X1 U15891 ( .A(n13796), .B(n13799), .ZN(n14972) );
  AOI22_X1 U15892 ( .A1(n13854), .A2(n13798), .B1(n13797), .B2(n13851), .ZN(
        n13802) );
  OAI211_X1 U15893 ( .C1(n6718), .C2(n7505), .A(n15313), .B(n13800), .ZN(
        n13801) );
  OAI211_X1 U15894 ( .C1(n14972), .C2(n6801), .A(n13802), .B(n13801), .ZN(
        n14975) );
  NAND2_X1 U15895 ( .A1(n14975), .A2(n13883), .ZN(n13810) );
  OAI22_X1 U15896 ( .A1(n13883), .A2(n13804), .B1(n13803), .B2(n13880), .ZN(
        n13807) );
  OAI211_X1 U15897 ( .C1(n14974), .C2(n13825), .A(n13805), .B(n15323), .ZN(
        n14973) );
  NOR2_X1 U15898 ( .A1(n14973), .A2(n13886), .ZN(n13806) );
  AOI211_X1 U15899 ( .C1(n15317), .C2(n13808), .A(n13807), .B(n13806), .ZN(
        n13809) );
  OAI211_X1 U15900 ( .C1(n14972), .C2(n13892), .A(n13810), .B(n13809), .ZN(
        P2_U3253) );
  OR2_X1 U15901 ( .A1(n13811), .A2(n13815), .ZN(n13812) );
  NAND2_X1 U15902 ( .A1(n13813), .A2(n13812), .ZN(n15439) );
  OR2_X1 U15903 ( .A1(n15439), .A2(n6801), .ZN(n13822) );
  AOI22_X1 U15904 ( .A1(n13851), .A2(n13814), .B1(n13852), .B2(n13854), .ZN(
        n13821) );
  NAND2_X1 U15905 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  NAND2_X1 U15906 ( .A1(n13818), .A2(n13817), .ZN(n13819) );
  NAND2_X1 U15907 ( .A1(n13819), .A2(n15313), .ZN(n13820) );
  NAND3_X1 U15908 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n15441) );
  NAND2_X1 U15909 ( .A1(n15441), .A2(n13883), .ZN(n13831) );
  OAI22_X1 U15910 ( .A1(n13883), .A2(n13824), .B1(n13823), .B2(n13880), .ZN(
        n13829) );
  INV_X1 U15911 ( .A(n13825), .ZN(n13827) );
  AOI21_X1 U15912 ( .B1(n13842), .B2(n15435), .A(n13979), .ZN(n13826) );
  NAND2_X1 U15913 ( .A1(n13827), .A2(n13826), .ZN(n15437) );
  NOR2_X1 U15914 ( .A1(n15437), .A2(n13886), .ZN(n13828) );
  AOI211_X1 U15915 ( .C1(n15317), .C2(n15435), .A(n13829), .B(n13828), .ZN(
        n13830) );
  OAI211_X1 U15916 ( .C1(n15439), .C2(n13892), .A(n13831), .B(n13830), .ZN(
        P2_U3254) );
  XNOR2_X1 U15917 ( .A(n13832), .B(n13833), .ZN(n15426) );
  XNOR2_X1 U15918 ( .A(n13834), .B(n13833), .ZN(n13837) );
  OAI22_X1 U15919 ( .A1(n13873), .A2(n13874), .B1(n13835), .B2(n13872), .ZN(
        n13836) );
  AOI21_X1 U15920 ( .B1(n13837), .B2(n15313), .A(n13836), .ZN(n13838) );
  OAI21_X1 U15921 ( .B1(n15426), .B2(n6801), .A(n13838), .ZN(n15429) );
  NAND2_X1 U15922 ( .A1(n15429), .A2(n13883), .ZN(n13847) );
  OAI22_X1 U15923 ( .A1(n13883), .A2(n13840), .B1(n13839), .B2(n13880), .ZN(
        n13844) );
  OAI211_X1 U15924 ( .C1(n13841), .C2(n8918), .A(n15323), .B(n13842), .ZN(
        n15427) );
  NOR2_X1 U15925 ( .A1(n15427), .A2(n13886), .ZN(n13843) );
  AOI211_X1 U15926 ( .C1(n15317), .C2(n13845), .A(n13844), .B(n13843), .ZN(
        n13846) );
  OAI211_X1 U15927 ( .C1(n15426), .C2(n13892), .A(n13847), .B(n13846), .ZN(
        P2_U3255) );
  OR2_X1 U15928 ( .A1(n13848), .A2(n13855), .ZN(n13849) );
  NAND2_X1 U15929 ( .A1(n13850), .A2(n13849), .ZN(n15420) );
  AOI22_X1 U15930 ( .A1(n13854), .A2(n13853), .B1(n13852), .B2(n13851), .ZN(
        n13859) );
  XNOR2_X1 U15931 ( .A(n13856), .B(n13855), .ZN(n13857) );
  NAND2_X1 U15932 ( .A1(n13857), .A2(n15313), .ZN(n13858) );
  OAI211_X1 U15933 ( .C1(n15420), .C2(n6801), .A(n13859), .B(n13858), .ZN(
        n15423) );
  NAND2_X1 U15934 ( .A1(n15423), .A2(n13883), .ZN(n13867) );
  OAI22_X1 U15935 ( .A1(n13883), .A2(n13861), .B1(n13860), .B2(n13880), .ZN(
        n13864) );
  INV_X1 U15936 ( .A(n13884), .ZN(n13862) );
  INV_X1 U15937 ( .A(n13865), .ZN(n15422) );
  OAI211_X1 U15938 ( .C1(n13862), .C2(n15422), .A(n15323), .B(n7040), .ZN(
        n15421) );
  NOR2_X1 U15939 ( .A1(n15421), .A2(n13886), .ZN(n13863) );
  AOI211_X1 U15940 ( .C1(n15317), .C2(n13865), .A(n13864), .B(n13863), .ZN(
        n13866) );
  OAI211_X1 U15941 ( .C1(n15420), .C2(n13892), .A(n13867), .B(n13866), .ZN(
        P2_U3256) );
  XNOR2_X1 U15942 ( .A(n13869), .B(n13868), .ZN(n15413) );
  XNOR2_X1 U15943 ( .A(n13871), .B(n13870), .ZN(n13877) );
  OAI22_X1 U15944 ( .A1(n13875), .A2(n13874), .B1(n13873), .B2(n13872), .ZN(
        n13876) );
  AOI21_X1 U15945 ( .B1(n13877), .B2(n15313), .A(n13876), .ZN(n13878) );
  OAI21_X1 U15946 ( .B1(n6801), .B2(n15413), .A(n13878), .ZN(n15416) );
  NAND2_X1 U15947 ( .A1(n15416), .A2(n13883), .ZN(n13891) );
  OAI22_X1 U15948 ( .A1(n13883), .A2(n13882), .B1(n13881), .B2(n13880), .ZN(
        n13888) );
  OAI211_X1 U15949 ( .C1(n13885), .C2(n15415), .A(n15323), .B(n13884), .ZN(
        n15414) );
  NOR2_X1 U15950 ( .A1(n15414), .A2(n13886), .ZN(n13887) );
  AOI211_X1 U15951 ( .C1(n15317), .C2(n13889), .A(n13888), .B(n13887), .ZN(
        n13890) );
  OAI211_X1 U15952 ( .C1(n15413), .C2(n13892), .A(n13891), .B(n13890), .ZN(
        P2_U3257) );
  OAI211_X1 U15953 ( .C1(n13894), .C2(n15428), .A(n13893), .B(n13895), .ZN(
        n13983) );
  MUX2_X1 U15954 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13983), .S(n15457), .Z(
        P2_U3530) );
  OAI211_X1 U15955 ( .C1(n13897), .C2(n15428), .A(n13896), .B(n13895), .ZN(
        n13984) );
  MUX2_X1 U15956 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13984), .S(n15457), .Z(
        P2_U3529) );
  AOI21_X1 U15957 ( .B1(n15434), .B2(n13899), .A(n13898), .ZN(n13900) );
  OAI211_X1 U15958 ( .C1(n15407), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        n13985) );
  MUX2_X1 U15959 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13985), .S(n15457), .Z(
        P2_U3527) );
  INV_X1 U15960 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13911) );
  NAND3_X1 U15961 ( .A1(n13904), .A2(n13903), .A3(n15379), .ZN(n13908) );
  NAND2_X1 U15962 ( .A1(n13905), .A2(n15434), .ZN(n13907) );
  NAND3_X1 U15963 ( .A1(n13908), .A2(n13907), .A3(n13906), .ZN(n13909) );
  NOR2_X1 U15964 ( .A1(n13910), .A2(n13909), .ZN(n13986) );
  MUX2_X1 U15965 ( .A(n13911), .B(n13986), .S(n15457), .Z(n13912) );
  INV_X1 U15966 ( .A(n13912), .ZN(P2_U3526) );
  NAND2_X1 U15967 ( .A1(n13914), .A2(n15379), .ZN(n13916) );
  OAI211_X1 U15968 ( .C1(n7274), .C2(n15428), .A(n13916), .B(n13915), .ZN(
        n13917) );
  MUX2_X1 U15969 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13989), .S(n15457), .Z(
        P2_U3525) );
  AOI21_X1 U15970 ( .B1(n15434), .B2(n13920), .A(n13919), .ZN(n13921) );
  OAI211_X1 U15971 ( .C1(n15407), .C2(n13923), .A(n13922), .B(n13921), .ZN(
        n13990) );
  MUX2_X1 U15972 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13990), .S(n15457), .Z(
        P2_U3524) );
  AOI21_X1 U15973 ( .B1(n15434), .B2(n13925), .A(n13924), .ZN(n13930) );
  NAND3_X1 U15974 ( .A1(n13927), .A2(n15379), .A3(n13926), .ZN(n13928) );
  NAND3_X1 U15975 ( .A1(n13930), .A2(n13929), .A3(n13928), .ZN(n13991) );
  MUX2_X1 U15976 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13991), .S(n15457), .Z(
        P2_U3523) );
  NAND2_X1 U15977 ( .A1(n13931), .A2(n15379), .ZN(n13933) );
  OAI211_X1 U15978 ( .C1(n8920), .C2(n15428), .A(n13933), .B(n13932), .ZN(
        n13934) );
  MUX2_X1 U15979 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13992), .S(n15457), .Z(
        P2_U3522) );
  AOI21_X1 U15980 ( .B1(n15434), .B2(n13937), .A(n13936), .ZN(n13938) );
  OAI211_X1 U15981 ( .C1(n15407), .C2(n13940), .A(n13939), .B(n13938), .ZN(
        n13993) );
  MUX2_X1 U15982 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13993), .S(n15457), .Z(
        P2_U3521) );
  AOI211_X1 U15983 ( .C1(n15434), .C2(n13943), .A(n13942), .B(n13941), .ZN(
        n13944) );
  OAI21_X1 U15984 ( .B1(n15407), .B2(n13945), .A(n13944), .ZN(n13994) );
  MUX2_X1 U15985 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13994), .S(n15457), .Z(
        P2_U3520) );
  AOI211_X1 U15986 ( .C1(n15434), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        n13949) );
  OAI21_X1 U15987 ( .B1(n15407), .B2(n13950), .A(n13949), .ZN(n13995) );
  MUX2_X1 U15988 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13995), .S(n15457), .Z(
        P2_U3519) );
  AOI22_X1 U15989 ( .A1(n13952), .A2(n15323), .B1(n15434), .B2(n13951), .ZN(
        n13953) );
  OAI211_X1 U15990 ( .C1(n15407), .C2(n13955), .A(n13954), .B(n13953), .ZN(
        n13996) );
  MUX2_X1 U15991 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13996), .S(n15457), .Z(
        P2_U3518) );
  AOI21_X1 U15992 ( .B1(n15434), .B2(n13957), .A(n13956), .ZN(n13958) );
  OAI211_X1 U15993 ( .C1(n13960), .C2(n15407), .A(n13959), .B(n13958), .ZN(
        n13997) );
  MUX2_X1 U15994 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13997), .S(n15457), .Z(
        P2_U3517) );
  AOI21_X1 U15995 ( .B1(n15434), .B2(n13962), .A(n13961), .ZN(n13963) );
  OAI211_X1 U15996 ( .C1(n15407), .C2(n13965), .A(n13964), .B(n13963), .ZN(
        n13998) );
  MUX2_X1 U15997 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13998), .S(n15457), .Z(
        P2_U3516) );
  AOI21_X1 U15998 ( .B1(n15434), .B2(n13967), .A(n13966), .ZN(n13968) );
  OAI211_X1 U15999 ( .C1(n15438), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        n13999) );
  MUX2_X1 U16000 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13999), .S(n15457), .Z(
        P2_U3515) );
  XNOR2_X1 U16001 ( .A(n13972), .B(n13971), .ZN(n14960) );
  XNOR2_X1 U16002 ( .A(n13974), .B(n13973), .ZN(n13977) );
  INV_X1 U16003 ( .A(n13975), .ZN(n13976) );
  AOI21_X1 U16004 ( .B1(n13977), .B2(n15313), .A(n13976), .ZN(n14965) );
  AOI211_X1 U16005 ( .C1(n13981), .C2(n13980), .A(n13979), .B(n13978), .ZN(
        n14963) );
  AOI21_X1 U16006 ( .B1(n15434), .B2(n13981), .A(n14963), .ZN(n13982) );
  OAI211_X1 U16007 ( .C1(n15407), .C2(n14960), .A(n14965), .B(n13982), .ZN(
        n14000) );
  MUX2_X1 U16008 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14000), .S(n15457), .Z(
        P2_U3514) );
  MUX2_X1 U16009 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13983), .S(n15444), .Z(
        P2_U3498) );
  MUX2_X1 U16010 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13984), .S(n15444), .Z(
        P2_U3497) );
  MUX2_X1 U16011 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13985), .S(n15444), .Z(
        P2_U3495) );
  INV_X1 U16012 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13987) );
  MUX2_X1 U16013 ( .A(n13987), .B(n13986), .S(n15444), .Z(n13988) );
  INV_X1 U16014 ( .A(n13988), .ZN(P2_U3494) );
  MUX2_X1 U16015 ( .A(n13989), .B(P2_REG0_REG_26__SCAN_IN), .S(n15442), .Z(
        P2_U3493) );
  MUX2_X1 U16016 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13990), .S(n15444), .Z(
        P2_U3492) );
  MUX2_X1 U16017 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13991), .S(n15444), .Z(
        P2_U3491) );
  MUX2_X1 U16018 ( .A(n13992), .B(P2_REG0_REG_23__SCAN_IN), .S(n15442), .Z(
        P2_U3490) );
  MUX2_X1 U16019 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13993), .S(n15444), .Z(
        P2_U3489) );
  MUX2_X1 U16020 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13994), .S(n15444), .Z(
        P2_U3488) );
  MUX2_X1 U16021 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13995), .S(n15444), .Z(
        P2_U3487) );
  MUX2_X1 U16022 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13996), .S(n15444), .Z(
        P2_U3486) );
  MUX2_X1 U16023 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13997), .S(n15444), .Z(
        P2_U3484) );
  MUX2_X1 U16024 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13998), .S(n15444), .Z(
        P2_U3481) );
  MUX2_X1 U16025 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13999), .S(n15444), .Z(
        P2_U3478) );
  MUX2_X1 U16026 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14000), .S(n15444), .Z(
        P2_U3475) );
  INV_X1 U16027 ( .A(n14001), .ZN(n14712) );
  NAND3_X1 U16028 ( .A1(n14003), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14005) );
  OAI22_X1 U16029 ( .A1(n14002), .A2(n14005), .B1(n14004), .B2(n14024), .ZN(
        n14006) );
  INV_X1 U16030 ( .A(n14006), .ZN(n14007) );
  OAI21_X1 U16031 ( .B1(n14712), .B2(n14022), .A(n14007), .ZN(P2_U3296) );
  NAND2_X1 U16032 ( .A1(n14009), .A2(n14008), .ZN(n14011) );
  OAI211_X1 U16033 ( .C1(n14024), .C2(n14012), .A(n14011), .B(n14010), .ZN(
        P2_U3299) );
  INV_X1 U16034 ( .A(n14013), .ZN(n14719) );
  OAI222_X1 U16035 ( .A1(n14024), .A2(n14016), .B1(n14022), .B2(n14719), .C1(
        P2_U3088), .C2(n14014), .ZN(P2_U3300) );
  OAI222_X1 U16036 ( .A1(P2_U3088), .A2(n14019), .B1(n14022), .B2(n14018), 
        .C1(n14017), .C2(n14024), .ZN(P2_U3301) );
  OAI222_X1 U16037 ( .A1(n14024), .A2(n14023), .B1(n14022), .B2(n14021), .C1(
        P2_U3088), .C2(n14020), .ZN(P2_U3302) );
  INV_X1 U16038 ( .A(n14025), .ZN(n14026) );
  MUX2_X1 U16039 ( .A(n14026), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16040 ( .A(n14028), .B(n14027), .Z(n14034) );
  NAND2_X1 U16041 ( .A1(n14452), .A2(n14569), .ZN(n14030) );
  NAND2_X1 U16042 ( .A1(n14394), .A2(n14570), .ZN(n14029) );
  NAND2_X1 U16043 ( .A1(n14030), .A2(n14029), .ZN(n14418) );
  AOI22_X1 U16044 ( .A1(n14152), .A2(n14418), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14031) );
  OAI21_X1 U16045 ( .B1(n14998), .B2(n14427), .A(n14031), .ZN(n14032) );
  AOI21_X1 U16046 ( .B1(n14430), .B2(n14995), .A(n14032), .ZN(n14033) );
  OAI21_X1 U16047 ( .B1(n14034), .B2(n14989), .A(n14033), .ZN(P1_U3214) );
  XOR2_X1 U16048 ( .A(n14036), .B(n14035), .Z(n14041) );
  AOI22_X1 U16049 ( .A1(n14140), .A2(n14525), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14038) );
  NAND2_X1 U16050 ( .A1(n14141), .A2(n14488), .ZN(n14037) );
  OAI211_X1 U16051 ( .C1(n14998), .C2(n14494), .A(n14038), .B(n14037), .ZN(
        n14039) );
  AOI21_X1 U16052 ( .B1(n14645), .B2(n14995), .A(n14039), .ZN(n14040) );
  OAI21_X1 U16053 ( .B1(n14041), .B2(n14989), .A(n14040), .ZN(P1_U3216) );
  OAI211_X1 U16054 ( .C1(n14044), .C2(n14043), .A(n14042), .B(n14119), .ZN(
        n14049) );
  AOI22_X1 U16055 ( .A1(n14995), .A2(n14046), .B1(n14152), .B2(n14045), .ZN(
        n14048) );
  MUX2_X1 U16056 ( .A(n14998), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n14047) );
  NAND3_X1 U16057 ( .A1(n14049), .A2(n14048), .A3(n14047), .ZN(P1_U3218) );
  INV_X1 U16058 ( .A(n14670), .ZN(n14057) );
  AOI21_X1 U16059 ( .B1(n14051), .B2(n14050), .A(n14989), .ZN(n14053) );
  NAND2_X1 U16060 ( .A1(n14053), .A2(n14052), .ZN(n14056) );
  INV_X1 U16061 ( .A(n14370), .ZN(n14594) );
  OAI22_X1 U16062 ( .A1(n14353), .A2(n14593), .B1(n14594), .B2(n14591), .ZN(
        n14669) );
  AND2_X1 U16063 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14327) );
  NOR2_X1 U16064 ( .A1(n14998), .A2(n14555), .ZN(n14054) );
  AOI211_X1 U16065 ( .C1(n14152), .C2(n14669), .A(n14327), .B(n14054), .ZN(
        n14055) );
  OAI211_X1 U16066 ( .C1(n14057), .C2(n14128), .A(n14056), .B(n14055), .ZN(
        P1_U3219) );
  INV_X1 U16067 ( .A(n14058), .ZN(n14059) );
  AOI21_X1 U16068 ( .B1(n14061), .B2(n14060), .A(n14059), .ZN(n14066) );
  INV_X1 U16069 ( .A(n14140), .ZN(n14982) );
  NAND2_X1 U16070 ( .A1(n14134), .A2(n14521), .ZN(n14063) );
  AOI22_X1 U16071 ( .A1(n14141), .A2(n14525), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14062) );
  OAI211_X1 U16072 ( .C1(n14353), .C2(n14982), .A(n14063), .B(n14062), .ZN(
        n14064) );
  AOI21_X1 U16073 ( .B1(n14657), .B2(n14995), .A(n14064), .ZN(n14065) );
  OAI21_X1 U16074 ( .B1(n14066), .B2(n14989), .A(n14065), .ZN(P1_U3223) );
  XOR2_X1 U16075 ( .A(n14068), .B(n14067), .Z(n14073) );
  AOI22_X1 U16076 ( .A1(n14140), .A2(n14488), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14070) );
  NAND2_X1 U16077 ( .A1(n14141), .A2(n14452), .ZN(n14069) );
  OAI211_X1 U16078 ( .C1(n14998), .C2(n14458), .A(n14070), .B(n14069), .ZN(
        n14071) );
  AOI21_X1 U16079 ( .B1(n14635), .B2(n14995), .A(n14071), .ZN(n14072) );
  OAI21_X1 U16080 ( .B1(n14073), .B2(n14989), .A(n14072), .ZN(P1_U3225) );
  XOR2_X1 U16081 ( .A(n14075), .B(n14074), .Z(n14082) );
  NAND2_X1 U16082 ( .A1(n14141), .A2(n14568), .ZN(n14076) );
  OAI211_X1 U16083 ( .C1(n14982), .C2(n14984), .A(n14077), .B(n14076), .ZN(
        n14078) );
  AOI21_X1 U16084 ( .B1(n14079), .B2(n14134), .A(n14078), .ZN(n14081) );
  NAND2_X1 U16085 ( .A1(n14686), .A2(n14995), .ZN(n14080) );
  OAI211_X1 U16086 ( .C1(n14082), .C2(n14989), .A(n14081), .B(n14080), .ZN(
        P1_U3226) );
  XOR2_X1 U16087 ( .A(n14083), .B(n14084), .Z(n14089) );
  NAND2_X1 U16088 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14284)
         );
  OAI21_X1 U16089 ( .B1(n14982), .B2(n14592), .A(n14284), .ZN(n14085) );
  AOI21_X1 U16090 ( .B1(n14141), .B2(n14370), .A(n14085), .ZN(n14086) );
  OAI21_X1 U16091 ( .B1(n14585), .B2(n14998), .A(n14086), .ZN(n14087) );
  AOI21_X1 U16092 ( .B1(n14682), .B2(n14995), .A(n14087), .ZN(n14088) );
  OAI21_X1 U16093 ( .B1(n14089), .B2(n14989), .A(n14088), .ZN(P1_U3228) );
  XOR2_X1 U16094 ( .A(n14091), .B(n14090), .Z(n14096) );
  AOI22_X1 U16095 ( .A1(n14140), .A2(n14378), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14093) );
  NAND2_X1 U16096 ( .A1(n14141), .A2(n14381), .ZN(n14092) );
  OAI211_X1 U16097 ( .C1(n14998), .C2(n14479), .A(n14093), .B(n14092), .ZN(
        n14094) );
  AOI21_X1 U16098 ( .B1(n12250), .B2(n14995), .A(n14094), .ZN(n14095) );
  OAI21_X1 U16099 ( .B1(n14096), .B2(n14989), .A(n14095), .ZN(P1_U3229) );
  OAI211_X1 U16100 ( .C1(n14099), .C2(n14098), .A(n14097), .B(n14119), .ZN(
        n14106) );
  INV_X1 U16101 ( .A(n14100), .ZN(n14539) );
  NAND2_X1 U16102 ( .A1(n14374), .A2(n14570), .ZN(n14102) );
  NAND2_X1 U16103 ( .A1(n14571), .A2(n14569), .ZN(n14101) );
  AND2_X1 U16104 ( .A1(n14102), .A2(n14101), .ZN(n14661) );
  INV_X1 U16105 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14103) );
  OAI22_X1 U16106 ( .A1(n14124), .A2(n14661), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14103), .ZN(n14104) );
  AOI21_X1 U16107 ( .B1(n14539), .B2(n14134), .A(n14104), .ZN(n14105) );
  OAI211_X1 U16108 ( .C1(n14663), .C2(n14128), .A(n14106), .B(n14105), .ZN(
        P1_U3233) );
  OAI211_X1 U16109 ( .C1(n6583), .C2(n14107), .A(n14987), .B(n14119), .ZN(
        n14115) );
  NOR2_X1 U16110 ( .A1(n14998), .A2(n14109), .ZN(n14113) );
  OAI21_X1 U16111 ( .B1(n14983), .B2(n14111), .A(n14110), .ZN(n14112) );
  AOI211_X1 U16112 ( .C1(n14140), .C2(n14162), .A(n14113), .B(n14112), .ZN(
        n14114) );
  OAI211_X1 U16113 ( .C1(n15000), .C2(n14128), .A(n14115), .B(n14114), .ZN(
        P1_U3234) );
  OAI21_X1 U16114 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(n14120) );
  NAND2_X1 U16115 ( .A1(n14120), .A2(n14119), .ZN(n14127) );
  INV_X1 U16116 ( .A(n14121), .ZN(n14507) );
  AND2_X1 U16117 ( .A1(n14378), .A2(n14570), .ZN(n14122) );
  AOI21_X1 U16118 ( .B1(n14374), .B2(n14569), .A(n14122), .ZN(n14649) );
  INV_X1 U16119 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14123) );
  OAI22_X1 U16120 ( .A1(n14124), .A2(n14649), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14123), .ZN(n14125) );
  AOI21_X1 U16121 ( .B1(n14507), .B2(n14134), .A(n14125), .ZN(n14126) );
  OAI211_X1 U16122 ( .C1(n14128), .C2(n14651), .A(n14127), .B(n14126), .ZN(
        P1_U3235) );
  XOR2_X1 U16123 ( .A(n14130), .B(n14129), .Z(n14137) );
  NAND2_X1 U16124 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14300)
         );
  NAND2_X1 U16125 ( .A1(n14141), .A2(n14571), .ZN(n14131) );
  OAI211_X1 U16126 ( .C1(n14982), .C2(n14132), .A(n14300), .B(n14131), .ZN(
        n14133) );
  AOI21_X1 U16127 ( .B1(n14577), .B2(n14134), .A(n14133), .ZN(n14136) );
  NAND2_X1 U16128 ( .A1(n14677), .A2(n14995), .ZN(n14135) );
  OAI211_X1 U16129 ( .C1(n14137), .C2(n14989), .A(n14136), .B(n14135), .ZN(
        P1_U3238) );
  XOR2_X1 U16130 ( .A(n14139), .B(n14138), .Z(n14146) );
  AOI22_X1 U16131 ( .A1(n14140), .A2(n14381), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14143) );
  NAND2_X1 U16132 ( .A1(n14141), .A2(n14404), .ZN(n14142) );
  OAI211_X1 U16133 ( .C1(n14998), .C2(n14437), .A(n14143), .B(n14142), .ZN(
        n14144) );
  AOI21_X1 U16134 ( .B1(n14630), .B2(n14995), .A(n14144), .ZN(n14145) );
  OAI21_X1 U16135 ( .B1(n14146), .B2(n14989), .A(n14145), .ZN(P1_U3240) );
  NAND2_X1 U16136 ( .A1(n14148), .A2(n14147), .ZN(n14150) );
  XNOR2_X1 U16137 ( .A(n14150), .B(n14149), .ZN(n14158) );
  NAND2_X1 U16138 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15073)
         );
  NAND2_X1 U16139 ( .A1(n14152), .A2(n14151), .ZN(n14153) );
  OAI211_X1 U16140 ( .C1(n14998), .C2(n14154), .A(n15073), .B(n14153), .ZN(
        n14155) );
  AOI21_X1 U16141 ( .B1(n14156), .B2(n14995), .A(n14155), .ZN(n14157) );
  OAI21_X1 U16142 ( .B1(n14158), .B2(n14989), .A(n14157), .ZN(P1_U3241) );
  MUX2_X1 U16143 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14335), .S(n6576), .Z(
        P1_U3591) );
  MUX2_X1 U16144 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14391), .S(n6576), .Z(
        P1_U3590) );
  MUX2_X1 U16145 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14403), .S(n6576), .Z(
        P1_U3589) );
  MUX2_X1 U16146 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14394), .S(n6576), .Z(
        P1_U3588) );
  MUX2_X1 U16147 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14404), .S(n6576), .Z(
        P1_U3587) );
  MUX2_X1 U16148 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14452), .S(n6576), .Z(
        P1_U3586) );
  MUX2_X1 U16149 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14381), .S(n6576), .Z(
        P1_U3585) );
  MUX2_X1 U16150 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14488), .S(n6576), .Z(
        P1_U3584) );
  MUX2_X1 U16151 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14525), .S(n6576), .Z(
        P1_U3582) );
  MUX2_X1 U16152 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14374), .S(n6576), .Z(
        P1_U3581) );
  MUX2_X1 U16153 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14526), .S(n6576), .Z(
        P1_U3580) );
  MUX2_X1 U16154 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14571), .S(n6576), .Z(
        P1_U3579) );
  MUX2_X1 U16155 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14370), .S(n6576), .Z(
        P1_U3578) );
  MUX2_X1 U16156 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14568), .S(n6576), .Z(
        P1_U3577) );
  MUX2_X1 U16157 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14365), .S(n6576), .Z(
        P1_U3576) );
  MUX2_X1 U16158 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14159), .S(n6576), .Z(
        P1_U3575) );
  MUX2_X1 U16159 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14160), .S(n6576), .Z(
        P1_U3574) );
  MUX2_X1 U16160 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14161), .S(n6576), .Z(
        P1_U3573) );
  MUX2_X1 U16161 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14162), .S(n6576), .Z(
        P1_U3572) );
  MUX2_X1 U16162 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14163), .S(n6576), .Z(
        P1_U3571) );
  MUX2_X1 U16163 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14164), .S(n6576), .Z(
        P1_U3570) );
  MUX2_X1 U16164 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14165), .S(n6576), .Z(
        P1_U3569) );
  MUX2_X1 U16165 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14166), .S(n6576), .Z(
        P1_U3568) );
  MUX2_X1 U16166 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14167), .S(n6576), .Z(
        P1_U3567) );
  MUX2_X1 U16167 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14168), .S(n6576), .Z(
        P1_U3566) );
  MUX2_X1 U16168 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14169), .S(n6576), .Z(
        P1_U3565) );
  MUX2_X1 U16169 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14170), .S(n6576), .Z(
        P1_U3564) );
  MUX2_X1 U16170 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14171), .S(n6576), .Z(
        P1_U3563) );
  MUX2_X1 U16171 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14172), .S(n6576), .Z(
        P1_U3562) );
  MUX2_X1 U16172 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6776), .S(n6576), .Z(
        P1_U3561) );
  MUX2_X1 U16173 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14174), .S(n6576), .Z(
        P1_U3560) );
  OAI22_X1 U16174 ( .A1(n15075), .A2(n14724), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14175), .ZN(n14176) );
  AOI21_X1 U16175 ( .B1(n14177), .B2(n15067), .A(n14176), .ZN(n14186) );
  OAI211_X1 U16176 ( .C1(n14179), .C2(n14189), .A(n15070), .B(n14178), .ZN(
        n14185) );
  MUX2_X1 U16177 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9760), .S(n14180), .Z(
        n14181) );
  OAI21_X1 U16178 ( .B1(n9468), .B2(n14182), .A(n14181), .ZN(n14183) );
  NAND3_X1 U16179 ( .A1(n15071), .A2(n14200), .A3(n14183), .ZN(n14184) );
  NAND3_X1 U16180 ( .A1(n14186), .A2(n14185), .A3(n14184), .ZN(P1_U3244) );
  MUX2_X1 U16181 ( .A(n14189), .B(n14188), .S(n14187), .Z(n14191) );
  NAND2_X1 U16182 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  OAI211_X1 U16183 ( .C1(n14721), .C2(n14193), .A(n14192), .B(n6576), .ZN(
        n14237) );
  OAI22_X1 U16184 ( .A1(n15075), .A2(n14725), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14194), .ZN(n14195) );
  AOI21_X1 U16185 ( .B1(n14196), .B2(n15067), .A(n14195), .ZN(n14207) );
  MUX2_X1 U16186 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9763), .S(n14197), .Z(
        n14198) );
  NAND3_X1 U16187 ( .A1(n14200), .A2(n14199), .A3(n14198), .ZN(n14201) );
  NAND3_X1 U16188 ( .A1(n15071), .A2(n14216), .A3(n14201), .ZN(n14206) );
  OAI211_X1 U16189 ( .C1(n14204), .C2(n14203), .A(n15070), .B(n14202), .ZN(
        n14205) );
  NAND4_X1 U16190 ( .A1(n14237), .A2(n14207), .A3(n14206), .A4(n14205), .ZN(
        P1_U3245) );
  INV_X1 U16191 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14209) );
  INV_X1 U16192 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14208) );
  OAI22_X1 U16193 ( .A1(n15075), .A2(n14209), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14208), .ZN(n14210) );
  AOI21_X1 U16194 ( .B1(n14214), .B2(n15067), .A(n14210), .ZN(n14221) );
  OAI211_X1 U16195 ( .C1(n14213), .C2(n14212), .A(n15070), .B(n14211), .ZN(
        n14220) );
  MUX2_X1 U16196 ( .A(n9759), .B(P1_REG1_REG_3__SCAN_IN), .S(n14214), .Z(
        n14217) );
  NAND3_X1 U16197 ( .A1(n14217), .A2(n14216), .A3(n14215), .ZN(n14218) );
  NAND3_X1 U16198 ( .A1(n15071), .A2(n14231), .A3(n14218), .ZN(n14219) );
  NAND3_X1 U16199 ( .A1(n14221), .A2(n14220), .A3(n14219), .ZN(P1_U3246) );
  INV_X1 U16200 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14223) );
  OAI21_X1 U16201 ( .B1(n15075), .B2(n14223), .A(n14222), .ZN(n14224) );
  AOI21_X1 U16202 ( .B1(n14228), .B2(n15067), .A(n14224), .ZN(n14236) );
  OAI211_X1 U16203 ( .C1(n14227), .C2(n14226), .A(n15070), .B(n14225), .ZN(
        n14235) );
  MUX2_X1 U16204 ( .A(n9768), .B(P1_REG1_REG_4__SCAN_IN), .S(n14228), .Z(
        n14229) );
  NAND3_X1 U16205 ( .A1(n14231), .A2(n14230), .A3(n14229), .ZN(n14232) );
  NAND3_X1 U16206 ( .A1(n15071), .A2(n14233), .A3(n14232), .ZN(n14234) );
  NAND4_X1 U16207 ( .A1(n14237), .A2(n14236), .A3(n14235), .A4(n14234), .ZN(
        P1_U3247) );
  OAI211_X1 U16208 ( .C1(n14239), .C2(n14238), .A(n15071), .B(n14255), .ZN(
        n14249) );
  OAI211_X1 U16209 ( .C1(n14242), .C2(n14241), .A(n15070), .B(n14240), .ZN(
        n14248) );
  NOR2_X1 U16210 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14243), .ZN(n14244) );
  AOI21_X1 U16211 ( .B1(n14269), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14244), .ZN(
        n14247) );
  NAND2_X1 U16212 ( .A1(n15067), .A2(n14245), .ZN(n14246) );
  NAND4_X1 U16213 ( .A1(n14249), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        P1_U3249) );
  OAI211_X1 U16214 ( .C1(n14252), .C2(n14251), .A(n15070), .B(n14250), .ZN(
        n14263) );
  MUX2_X1 U16215 ( .A(n9775), .B(P1_REG1_REG_7__SCAN_IN), .S(n14258), .Z(
        n14253) );
  NAND3_X1 U16216 ( .A1(n14255), .A2(n14254), .A3(n14253), .ZN(n14256) );
  NAND3_X1 U16217 ( .A1(n15071), .A2(n14257), .A3(n14256), .ZN(n14262) );
  NAND2_X1 U16218 ( .A1(n15067), .A2(n14258), .ZN(n14261) );
  AOI21_X1 U16219 ( .B1(n14269), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14259), .ZN(
        n14260) );
  NAND4_X1 U16220 ( .A1(n14263), .A2(n14262), .A3(n14261), .A4(n14260), .ZN(
        P1_U3250) );
  AOI21_X1 U16221 ( .B1(n14265), .B2(n14264), .A(n15053), .ZN(n14267) );
  NAND2_X1 U16222 ( .A1(n14267), .A2(n14266), .ZN(n14277) );
  AOI21_X1 U16223 ( .B1(n14269), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14268), 
        .ZN(n14276) );
  OAI211_X1 U16224 ( .C1(n14272), .C2(n14271), .A(n15070), .B(n14270), .ZN(
        n14275) );
  NAND2_X1 U16225 ( .A1(n15067), .A2(n14273), .ZN(n14274) );
  NAND4_X1 U16226 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14274), .ZN(
        P1_U3253) );
  AOI21_X1 U16227 ( .B1(n14279), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14278), 
        .ZN(n14282) );
  NAND2_X1 U16228 ( .A1(n14296), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14280) );
  OAI21_X1 U16229 ( .B1(n14296), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14280), 
        .ZN(n14281) );
  NOR2_X1 U16230 ( .A1(n14282), .A2(n14281), .ZN(n14295) );
  AOI211_X1 U16231 ( .C1(n14282), .C2(n14281), .A(n14295), .B(n15046), .ZN(
        n14283) );
  INV_X1 U16232 ( .A(n14283), .ZN(n14294) );
  INV_X1 U16233 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14285) );
  OAI21_X1 U16234 ( .B1(n15075), .B2(n14285), .A(n14284), .ZN(n14286) );
  AOI21_X1 U16235 ( .B1(n14296), .B2(n15067), .A(n14286), .ZN(n14293) );
  XNOR2_X1 U16236 ( .A(n14304), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14291) );
  INV_X1 U16237 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14288) );
  OAI21_X1 U16238 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n14290) );
  NAND2_X1 U16239 ( .A1(n14291), .A2(n14290), .ZN(n14303) );
  OAI211_X1 U16240 ( .C1(n14291), .C2(n14290), .A(n15071), .B(n14303), .ZN(
        n14292) );
  NAND3_X1 U16241 ( .A1(n14294), .A2(n14293), .A3(n14292), .ZN(P1_U3260) );
  AOI21_X1 U16242 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14296), .A(n14295), 
        .ZN(n14311) );
  XNOR2_X1 U16243 ( .A(n14310), .B(n14311), .ZN(n14298) );
  NOR2_X1 U16244 ( .A1(n14297), .A2(n14298), .ZN(n14312) );
  AOI211_X1 U16245 ( .C1(n14298), .C2(n14297), .A(n14312), .B(n15046), .ZN(
        n14299) );
  INV_X1 U16246 ( .A(n14299), .ZN(n14309) );
  INV_X1 U16247 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U16248 ( .B1(n15075), .B2(n14301), .A(n14300), .ZN(n14302) );
  AOI21_X1 U16249 ( .B1(n14316), .B2(n15067), .A(n14302), .ZN(n14308) );
  OAI21_X1 U16250 ( .B1(n14305), .B2(n14304), .A(n14303), .ZN(n14315) );
  XNOR2_X1 U16251 ( .A(n14310), .B(n14315), .ZN(n14306) );
  NAND2_X1 U16252 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14306), .ZN(n14318) );
  OAI211_X1 U16253 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14306), .A(n15071), 
        .B(n14318), .ZN(n14307) );
  NAND3_X1 U16254 ( .A1(n14309), .A2(n14308), .A3(n14307), .ZN(P1_U3261) );
  NOR2_X1 U16255 ( .A1(n14311), .A2(n14310), .ZN(n14313) );
  NOR2_X1 U16256 ( .A1(n14313), .A2(n14312), .ZN(n14314) );
  XNOR2_X1 U16257 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14314), .ZN(n14324) );
  INV_X1 U16258 ( .A(n14324), .ZN(n14322) );
  NAND2_X1 U16259 ( .A1(n14316), .A2(n14315), .ZN(n14317) );
  NAND2_X1 U16260 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  XOR2_X1 U16261 ( .A(n14319), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14323) );
  OAI21_X1 U16262 ( .B1(n14323), .B2(n15053), .A(n14320), .ZN(n14321) );
  AOI21_X1 U16263 ( .B1(n14322), .B2(n15070), .A(n14321), .ZN(n14326) );
  AOI22_X1 U16264 ( .A1(n14324), .A2(n15070), .B1(n15071), .B2(n14323), .ZN(
        n14325) );
  MUX2_X1 U16265 ( .A(n14326), .B(n14325), .S(n9547), .Z(n14329) );
  INV_X1 U16266 ( .A(n14327), .ZN(n14328) );
  OAI211_X1 U16267 ( .C1(n7723), .C2(n15075), .A(n14329), .B(n14328), .ZN(
        P1_U3262) );
  INV_X1 U16268 ( .A(n14430), .ZN(n14623) );
  INV_X1 U16269 ( .A(n14635), .ZN(n14330) );
  NAND2_X1 U16270 ( .A1(n14554), .A2(n14663), .ZN(n14537) );
  NAND2_X1 U16271 ( .A1(n14330), .A2(n14477), .ZN(n14461) );
  XNOR2_X1 U16272 ( .A(n14339), .B(n14336), .ZN(n14332) );
  NAND2_X1 U16273 ( .A1(n14332), .A2(n14538), .ZN(n14602) );
  NAND2_X1 U16274 ( .A1(n14333), .A2(P1_B_REG_SCAN_IN), .ZN(n14334) );
  AND2_X1 U16275 ( .A1(n14570), .A2(n14334), .ZN(n14390) );
  NAND2_X1 U16276 ( .A1(n14335), .A2(n14390), .ZN(n14604) );
  NOR2_X1 U16277 ( .A1(n15098), .A2(n14604), .ZN(n14343) );
  INV_X1 U16278 ( .A(n14336), .ZN(n14603) );
  NOR2_X1 U16279 ( .A1(n14603), .A2(n15088), .ZN(n14337) );
  AOI211_X1 U16280 ( .C1(n15098), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14343), 
        .B(n14337), .ZN(n14338) );
  OAI21_X1 U16281 ( .B1(n14602), .B2(n14543), .A(n14338), .ZN(P1_U3263) );
  INV_X1 U16282 ( .A(n14388), .ZN(n14341) );
  INV_X1 U16283 ( .A(n14339), .ZN(n14340) );
  OAI211_X1 U16284 ( .C1(n14606), .C2(n14341), .A(n14340), .B(n14538), .ZN(
        n14605) );
  NOR2_X1 U16285 ( .A1(n14606), .A2(n15088), .ZN(n14342) );
  AOI211_X1 U16286 ( .C1(n15086), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14343), 
        .B(n14342), .ZN(n14344) );
  OAI21_X1 U16287 ( .B1(n14605), .B2(n14543), .A(n14344), .ZN(P1_U3264) );
  INV_X1 U16288 ( .A(n14509), .ZN(n14503) );
  NAND2_X1 U16289 ( .A1(n14686), .A2(n14592), .ZN(n14345) );
  OR2_X1 U16290 ( .A1(n14677), .A2(n14594), .ZN(n14349) );
  OR2_X1 U16291 ( .A1(n14540), .A2(n14353), .ZN(n14354) );
  INV_X1 U16292 ( .A(n14522), .ZN(n14520) );
  NOR2_X1 U16293 ( .A1(n14657), .A2(n14355), .ZN(n14356) );
  NAND2_X1 U16294 ( .A1(n14503), .A2(n14502), .ZN(n14501) );
  NAND2_X1 U16295 ( .A1(n14501), .A2(n14357), .ZN(n14487) );
  INV_X1 U16296 ( .A(n14491), .ZN(n14486) );
  NAND2_X1 U16297 ( .A1(n14487), .A2(n14486), .ZN(n14485) );
  NAND2_X1 U16298 ( .A1(n14645), .A2(n14470), .ZN(n14358) );
  INV_X1 U16299 ( .A(n12250), .ZN(n14478) );
  NAND2_X1 U16300 ( .A1(n14478), .A2(n14488), .ZN(n14359) );
  NAND2_X1 U16301 ( .A1(n14441), .A2(n14442), .ZN(n14440) );
  INV_X1 U16302 ( .A(n14452), .ZN(n14361) );
  NAND2_X1 U16303 ( .A1(n14630), .A2(n14361), .ZN(n14362) );
  NAND2_X1 U16304 ( .A1(n14440), .A2(n14362), .ZN(n14417) );
  OR2_X1 U16305 ( .A1(n14686), .A2(n14365), .ZN(n14366) );
  NAND2_X1 U16306 ( .A1(n14682), .A2(n14568), .ZN(n14368) );
  OR2_X1 U16307 ( .A1(n14677), .A2(n14370), .ZN(n14369) );
  NAND2_X1 U16308 ( .A1(n14677), .A2(n14370), .ZN(n14371) );
  OR2_X1 U16309 ( .A1(n14670), .A2(n14571), .ZN(n14373) );
  INV_X1 U16310 ( .A(n14546), .ZN(n14536) );
  OR2_X1 U16311 ( .A1(n14657), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U16312 ( .A1(n14510), .A2(n14509), .ZN(n14508) );
  NAND2_X1 U16313 ( .A1(n14651), .A2(n14376), .ZN(n14377) );
  NAND2_X1 U16314 ( .A1(n14508), .A2(n14377), .ZN(n14490) );
  NAND2_X1 U16315 ( .A1(n14478), .A2(n14379), .ZN(n14380) );
  NAND2_X1 U16316 ( .A1(n14635), .A2(n14381), .ZN(n14382) );
  INV_X1 U16317 ( .A(n14441), .ZN(n14434) );
  NAND2_X1 U16318 ( .A1(n14435), .A2(n14434), .ZN(n14384) );
  NAND2_X1 U16319 ( .A1(n14630), .A2(n14452), .ZN(n14383) );
  OR2_X1 U16320 ( .A1(n14430), .A2(n14404), .ZN(n14386) );
  OAI21_X1 U16321 ( .B1(n14611), .B2(n14409), .A(n14388), .ZN(n14608) );
  NOR2_X1 U16322 ( .A1(n14608), .A2(n14389), .ZN(n14399) );
  NAND2_X1 U16323 ( .A1(n14391), .A2(n14390), .ZN(n14610) );
  OAI22_X1 U16324 ( .A1(n14393), .A2(n14610), .B1(n14392), .B2(n14556), .ZN(
        n14396) );
  NAND2_X1 U16325 ( .A1(n14394), .A2(n14569), .ZN(n14609) );
  NOR2_X1 U16326 ( .A1(n15086), .A2(n14609), .ZN(n14395) );
  AOI211_X1 U16327 ( .C1(n15098), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14396), 
        .B(n14395), .ZN(n14397) );
  OAI21_X1 U16328 ( .B1(n14611), .B2(n15088), .A(n14397), .ZN(n14398) );
  AOI211_X1 U16329 ( .C1(n14607), .C2(n14562), .A(n14399), .B(n14398), .ZN(
        n14400) );
  OAI21_X1 U16330 ( .B1(n14615), .B2(n14564), .A(n14400), .ZN(P1_U3356) );
  NAND2_X1 U16331 ( .A1(n14403), .A2(n14570), .ZN(n14406) );
  AOI211_X1 U16332 ( .C1(n14618), .C2(n14426), .A(n15091), .B(n14409), .ZN(
        n14617) );
  INV_X1 U16333 ( .A(n14410), .ZN(n14411) );
  AOI22_X1 U16334 ( .A1(n15098), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14411), 
        .B2(n15085), .ZN(n14412) );
  OAI21_X1 U16335 ( .B1(n7101), .B2(n15088), .A(n14412), .ZN(n14415) );
  OAI21_X1 U16336 ( .B1(n14420), .B2(n14417), .A(n14416), .ZN(n14419) );
  AOI21_X1 U16337 ( .B1(n14419), .B2(n6917), .A(n14418), .ZN(n14425) );
  NAND2_X1 U16338 ( .A1(n14421), .A2(n14420), .ZN(n14422) );
  NAND2_X1 U16339 ( .A1(n14423), .A2(n14422), .ZN(n14625) );
  NAND2_X1 U16340 ( .A1(n14625), .A2(n15084), .ZN(n14424) );
  OAI211_X1 U16341 ( .C1(n14623), .C2(n14436), .A(n14538), .B(n14426), .ZN(
        n14622) );
  OAI22_X1 U16342 ( .A1(n14547), .A2(n14428), .B1(n14427), .B2(n14556), .ZN(
        n14429) );
  AOI21_X1 U16343 ( .B1(n14430), .B2(n14558), .A(n14429), .ZN(n14431) );
  OAI21_X1 U16344 ( .B1(n14622), .B2(n14543), .A(n14431), .ZN(n14432) );
  AOI21_X1 U16345 ( .B1(n14625), .B2(n15095), .A(n14432), .ZN(n14433) );
  OAI21_X1 U16346 ( .B1(n14627), .B2(n15098), .A(n14433), .ZN(P1_U3266) );
  XNOR2_X1 U16347 ( .A(n14435), .B(n14434), .ZN(n14633) );
  AOI211_X1 U16348 ( .C1(n14630), .C2(n14461), .A(n15091), .B(n14436), .ZN(
        n14628) );
  INV_X1 U16349 ( .A(n14628), .ZN(n14446) );
  INV_X1 U16350 ( .A(n14437), .ZN(n14439) );
  OAI22_X1 U16351 ( .A1(n14469), .A2(n14591), .B1(n14438), .B2(n14593), .ZN(
        n14629) );
  AOI21_X1 U16352 ( .B1(n15085), .B2(n14439), .A(n14629), .ZN(n14444) );
  OAI21_X1 U16353 ( .B1(n14442), .B2(n14441), .A(n14440), .ZN(n14443) );
  NAND2_X1 U16354 ( .A1(n14443), .A2(n6917), .ZN(n14631) );
  OAI211_X1 U16355 ( .C1(n14446), .C2(n14445), .A(n14444), .B(n14631), .ZN(
        n14447) );
  NAND2_X1 U16356 ( .A1(n14447), .A2(n14547), .ZN(n14449) );
  AOI22_X1 U16357 ( .A1(n14630), .A2(n14558), .B1(n15086), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n14448) );
  OAI211_X1 U16358 ( .C1(n14633), .C2(n14601), .A(n14449), .B(n14448), .ZN(
        P1_U3267) );
  OAI21_X1 U16359 ( .B1(n14451), .B2(n6705), .A(n14450), .ZN(n14453) );
  AOI222_X1 U16360 ( .A1(n6917), .A2(n14453), .B1(n14452), .B2(n14570), .C1(
        n14488), .C2(n14569), .ZN(n14637) );
  OAI21_X1 U16361 ( .B1(n14456), .B2(n14455), .A(n14454), .ZN(n14638) );
  NAND2_X1 U16362 ( .A1(n15086), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14457) );
  OAI21_X1 U16363 ( .B1(n14556), .B2(n14458), .A(n14457), .ZN(n14459) );
  AOI21_X1 U16364 ( .B1(n14635), .B2(n14558), .A(n14459), .ZN(n14464) );
  INV_X1 U16365 ( .A(n14477), .ZN(n14460) );
  AOI21_X1 U16366 ( .B1(n14460), .B2(n14635), .A(n15091), .ZN(n14462) );
  AND2_X1 U16367 ( .A1(n14462), .A2(n14461), .ZN(n14634) );
  NAND2_X1 U16368 ( .A1(n14634), .A2(n15094), .ZN(n14463) );
  OAI211_X1 U16369 ( .C1(n14638), .C2(n14601), .A(n14464), .B(n14463), .ZN(
        n14465) );
  INV_X1 U16370 ( .A(n14465), .ZN(n14466) );
  OAI21_X1 U16371 ( .B1(n14637), .B2(n15098), .A(n14466), .ZN(P1_U3268) );
  OAI21_X1 U16372 ( .B1(n14467), .B2(n14474), .A(n14468), .ZN(n14639) );
  OAI22_X1 U16373 ( .A1(n14470), .A2(n14591), .B1(n14469), .B2(n14593), .ZN(
        n14476) );
  INV_X1 U16374 ( .A(n14471), .ZN(n14472) );
  AOI211_X1 U16375 ( .C1(n14474), .C2(n14473), .A(n15178), .B(n14472), .ZN(
        n14475) );
  AOI211_X1 U16376 ( .C1(n15084), .C2(n14639), .A(n14476), .B(n14475), .ZN(
        n14642) );
  AOI211_X1 U16377 ( .C1(n12250), .C2(n6627), .A(n15091), .B(n14477), .ZN(
        n14640) );
  NOR2_X1 U16378 ( .A1(n14478), .A2(n15088), .ZN(n14482) );
  OAI22_X1 U16379 ( .A1(n14547), .A2(n14480), .B1(n14479), .B2(n14556), .ZN(
        n14481) );
  AOI211_X1 U16380 ( .C1(n14640), .C2(n15094), .A(n14482), .B(n14481), .ZN(
        n14484) );
  NAND2_X1 U16381 ( .A1(n14639), .A2(n15095), .ZN(n14483) );
  OAI211_X1 U16382 ( .C1(n14642), .C2(n15086), .A(n14484), .B(n14483), .ZN(
        P1_U3269) );
  OAI21_X1 U16383 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14489) );
  AOI222_X1 U16384 ( .A1(n6917), .A2(n14489), .B1(n14488), .B2(n14570), .C1(
        n14525), .C2(n14569), .ZN(n14647) );
  OAI21_X1 U16385 ( .B1(n14492), .B2(n14491), .A(n7146), .ZN(n14648) );
  NAND2_X1 U16386 ( .A1(n15086), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14493) );
  OAI21_X1 U16387 ( .B1(n14556), .B2(n14494), .A(n14493), .ZN(n14495) );
  AOI21_X1 U16388 ( .B1(n14645), .B2(n14558), .A(n14495), .ZN(n14498) );
  AOI21_X1 U16389 ( .B1(n14645), .B2(n14511), .A(n15091), .ZN(n14496) );
  AND2_X1 U16390 ( .A1(n14496), .A2(n6627), .ZN(n14644) );
  NAND2_X1 U16391 ( .A1(n14644), .A2(n15094), .ZN(n14497) );
  OAI211_X1 U16392 ( .C1(n14648), .C2(n14601), .A(n14498), .B(n14497), .ZN(
        n14499) );
  INV_X1 U16393 ( .A(n14499), .ZN(n14500) );
  OAI21_X1 U16394 ( .B1(n14647), .B2(n15086), .A(n14500), .ZN(P1_U3270) );
  INV_X1 U16395 ( .A(n14649), .ZN(n14506) );
  OAI21_X1 U16396 ( .B1(n14503), .B2(n14502), .A(n14501), .ZN(n14504) );
  NAND2_X1 U16397 ( .A1(n14504), .A2(n6917), .ZN(n14654) );
  INV_X1 U16398 ( .A(n14654), .ZN(n14505) );
  AOI211_X1 U16399 ( .C1(n15085), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14516) );
  OAI21_X1 U16400 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n14653) );
  OAI211_X1 U16401 ( .C1(n14651), .C2(n14529), .A(n14538), .B(n14511), .ZN(
        n14650) );
  AOI22_X1 U16402 ( .A1(n14512), .A2(n14558), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15098), .ZN(n14513) );
  OAI21_X1 U16403 ( .B1(n14650), .B2(n14543), .A(n14513), .ZN(n14514) );
  AOI21_X1 U16404 ( .B1(n14653), .B2(n14562), .A(n14514), .ZN(n14515) );
  OAI21_X1 U16405 ( .B1(n14516), .B2(n15098), .A(n14515), .ZN(P1_U3271) );
  INV_X1 U16406 ( .A(n14517), .ZN(n14518) );
  AOI21_X1 U16407 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14660) );
  INV_X1 U16408 ( .A(n14521), .ZN(n14527) );
  XNOR2_X1 U16409 ( .A(n14523), .B(n14522), .ZN(n14524) );
  AOI222_X1 U16410 ( .A1(n14526), .A2(n14569), .B1(n14525), .B2(n14570), .C1(
        n6917), .C2(n14524), .ZN(n14659) );
  OAI21_X1 U16411 ( .B1(n14527), .B2(n14556), .A(n14659), .ZN(n14528) );
  NAND2_X1 U16412 ( .A1(n14528), .A2(n14547), .ZN(n14534) );
  AOI211_X1 U16413 ( .C1(n14657), .C2(n14537), .A(n15091), .B(n14529), .ZN(
        n14656) );
  INV_X1 U16414 ( .A(n14657), .ZN(n14531) );
  INV_X1 U16415 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14530) );
  OAI22_X1 U16416 ( .A1(n14531), .A2(n15088), .B1(n14530), .B2(n14547), .ZN(
        n14532) );
  AOI21_X1 U16417 ( .B1(n14656), .B2(n15094), .A(n14532), .ZN(n14533) );
  OAI211_X1 U16418 ( .C1(n14660), .C2(n14601), .A(n14534), .B(n14533), .ZN(
        P1_U3272) );
  AOI21_X1 U16419 ( .B1(n14536), .B2(n14535), .A(n6717), .ZN(n14666) );
  OAI211_X1 U16420 ( .C1(n14554), .C2(n14663), .A(n14538), .B(n14537), .ZN(
        n14662) );
  AOI22_X1 U16421 ( .A1(n15086), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14539), 
        .B2(n15085), .ZN(n14542) );
  NAND2_X1 U16422 ( .A1(n14540), .A2(n14558), .ZN(n14541) );
  OAI211_X1 U16423 ( .C1(n14662), .C2(n14543), .A(n14542), .B(n14541), .ZN(
        n14544) );
  AOI21_X1 U16424 ( .B1(n14666), .B2(n14562), .A(n14544), .ZN(n14550) );
  AOI211_X1 U16425 ( .C1(n14546), .C2(n14545), .A(n15178), .B(n6607), .ZN(
        n14664) );
  INV_X1 U16426 ( .A(n14661), .ZN(n14548) );
  OAI21_X1 U16427 ( .B1(n14664), .B2(n14548), .A(n14547), .ZN(n14549) );
  NAND2_X1 U16428 ( .A1(n14550), .A2(n14549), .ZN(P1_U3273) );
  XNOR2_X1 U16429 ( .A(n14551), .B(n14553), .ZN(n14674) );
  XNOR2_X1 U16430 ( .A(n14552), .B(n14553), .ZN(n14671) );
  AOI211_X1 U16431 ( .C1(n14670), .C2(n14575), .A(n15091), .B(n14554), .ZN(
        n14668) );
  NOR2_X1 U16432 ( .A1(n14556), .A2(n14555), .ZN(n14557) );
  AOI211_X1 U16433 ( .C1(n14668), .C2(n9547), .A(n14557), .B(n14669), .ZN(
        n14560) );
  AOI22_X1 U16434 ( .A1(n14670), .A2(n14558), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n15098), .ZN(n14559) );
  OAI21_X1 U16435 ( .B1(n14560), .B2(n15086), .A(n14559), .ZN(n14561) );
  AOI21_X1 U16436 ( .B1(n14562), .B2(n14671), .A(n14561), .ZN(n14563) );
  OAI21_X1 U16437 ( .B1(n14674), .B2(n14564), .A(n14563), .ZN(P1_U3274) );
  XNOR2_X1 U16438 ( .A(n14565), .B(n14566), .ZN(n14675) );
  XNOR2_X1 U16439 ( .A(n14567), .B(n14566), .ZN(n14573) );
  AOI22_X1 U16440 ( .A1(n14571), .A2(n14570), .B1(n14569), .B2(n14568), .ZN(
        n14572) );
  OAI21_X1 U16441 ( .B1(n14573), .B2(n15178), .A(n14572), .ZN(n14574) );
  AOI21_X1 U16442 ( .B1(n14675), .B2(n15084), .A(n14574), .ZN(n14679) );
  INV_X1 U16443 ( .A(n14575), .ZN(n14576) );
  AOI211_X1 U16444 ( .C1(n14677), .C2(n14583), .A(n15091), .B(n14576), .ZN(
        n14676) );
  NAND2_X1 U16445 ( .A1(n14676), .A2(n15094), .ZN(n14579) );
  AOI22_X1 U16446 ( .A1(n15086), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14577), 
        .B2(n15085), .ZN(n14578) );
  OAI211_X1 U16447 ( .C1(n7103), .C2(n15088), .A(n14579), .B(n14578), .ZN(
        n14580) );
  AOI21_X1 U16448 ( .B1(n15095), .B2(n14675), .A(n14580), .ZN(n14581) );
  OAI21_X1 U16449 ( .B1(n14679), .B2(n15086), .A(n14581), .ZN(P1_U3275) );
  XOR2_X1 U16450 ( .A(n14582), .B(n14589), .Z(n14685) );
  AOI211_X1 U16451 ( .C1(n14682), .C2(n14584), .A(n15091), .B(n7104), .ZN(
        n14681) );
  INV_X1 U16452 ( .A(n14585), .ZN(n14586) );
  AOI22_X1 U16453 ( .A1(n15086), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14586), 
        .B2(n15085), .ZN(n14587) );
  OAI21_X1 U16454 ( .B1(n14588), .B2(n15088), .A(n14587), .ZN(n14599) );
  AOI21_X1 U16455 ( .B1(n14590), .B2(n14589), .A(n15178), .ZN(n14597) );
  OAI22_X1 U16456 ( .A1(n14594), .A2(n14593), .B1(n14592), .B2(n14591), .ZN(
        n14595) );
  AOI21_X1 U16457 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n14684) );
  NOR2_X1 U16458 ( .A1(n14684), .A2(n15086), .ZN(n14598) );
  AOI211_X1 U16459 ( .C1(n14681), .C2(n15094), .A(n14599), .B(n14598), .ZN(
        n14600) );
  OAI21_X1 U16460 ( .B1(n14685), .B2(n14601), .A(n14600), .ZN(P1_U3276) );
  OAI211_X1 U16461 ( .C1(n14603), .C2(n15194), .A(n14602), .B(n14604), .ZN(
        n14693) );
  MUX2_X1 U16462 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14693), .S(n15213), .Z(
        P1_U3559) );
  OAI211_X1 U16463 ( .C1(n14606), .C2(n15194), .A(n14605), .B(n14604), .ZN(
        n14694) );
  MUX2_X1 U16464 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14694), .S(n15213), .Z(
        P1_U3558) );
  NAND2_X1 U16465 ( .A1(n14607), .A2(n15198), .ZN(n14616) );
  NOR2_X1 U16466 ( .A1(n14608), .A2(n15091), .ZN(n14613) );
  OAI211_X1 U16467 ( .C1(n14611), .C2(n15194), .A(n14610), .B(n14609), .ZN(
        n14612) );
  MUX2_X1 U16468 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14695), .S(n15213), .Z(
        P1_U3557) );
  AOI21_X1 U16469 ( .B1(n14618), .B2(n15169), .A(n14617), .ZN(n14619) );
  OAI211_X1 U16470 ( .C1(n15131), .C2(n14621), .A(n14620), .B(n14619), .ZN(
        n14696) );
  MUX2_X1 U16471 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14696), .S(n15213), .Z(
        P1_U3556) );
  OAI21_X1 U16472 ( .B1(n14623), .B2(n15194), .A(n14622), .ZN(n14624) );
  AOI21_X1 U16473 ( .B1(n14625), .B2(n15157), .A(n14624), .ZN(n14626) );
  NAND2_X1 U16474 ( .A1(n14627), .A2(n14626), .ZN(n14697) );
  MUX2_X1 U16475 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14697), .S(n15213), .Z(
        P1_U3555) );
  AOI211_X1 U16476 ( .C1(n14630), .C2(n15169), .A(n14629), .B(n14628), .ZN(
        n14632) );
  OAI211_X1 U16477 ( .C1(n15131), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14698) );
  MUX2_X1 U16478 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14698), .S(n15213), .Z(
        P1_U3554) );
  AOI21_X1 U16479 ( .B1(n14635), .B2(n15169), .A(n14634), .ZN(n14636) );
  OAI211_X1 U16480 ( .C1(n15131), .C2(n14638), .A(n14637), .B(n14636), .ZN(
        n14699) );
  MUX2_X1 U16481 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14699), .S(n15213), .Z(
        P1_U3553) );
  INV_X1 U16482 ( .A(n14639), .ZN(n14643) );
  AOI21_X1 U16483 ( .B1(n12250), .B2(n15169), .A(n14640), .ZN(n14641) );
  OAI211_X1 U16484 ( .C1(n14643), .C2(n15184), .A(n14642), .B(n14641), .ZN(
        n14700) );
  MUX2_X1 U16485 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14700), .S(n15213), .Z(
        P1_U3552) );
  AOI21_X1 U16486 ( .B1(n14645), .B2(n15169), .A(n14644), .ZN(n14646) );
  OAI211_X1 U16487 ( .C1(n15131), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        n14701) );
  MUX2_X1 U16488 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14701), .S(n15213), .Z(
        P1_U3551) );
  OAI211_X1 U16489 ( .C1(n15194), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        n14652) );
  AOI21_X1 U16490 ( .B1(n14653), .B2(n15198), .A(n14652), .ZN(n14655) );
  NAND2_X1 U16491 ( .A1(n14655), .A2(n14654), .ZN(n14702) );
  MUX2_X1 U16492 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14702), .S(n15213), .Z(
        P1_U3550) );
  AOI21_X1 U16493 ( .B1(n14657), .B2(n15169), .A(n14656), .ZN(n14658) );
  OAI211_X1 U16494 ( .C1(n14660), .C2(n15131), .A(n14659), .B(n14658), .ZN(
        n14703) );
  MUX2_X1 U16495 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14703), .S(n15213), .Z(
        P1_U3549) );
  OAI211_X1 U16496 ( .C1(n14663), .C2(n15194), .A(n14662), .B(n14661), .ZN(
        n14665) );
  AOI211_X1 U16497 ( .C1(n14666), .C2(n15198), .A(n14665), .B(n14664), .ZN(
        n14667) );
  INV_X1 U16498 ( .A(n14667), .ZN(n14704) );
  MUX2_X1 U16499 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14704), .S(n15213), .Z(
        P1_U3548) );
  AOI211_X1 U16500 ( .C1(n14670), .C2(n15169), .A(n14669), .B(n14668), .ZN(
        n14673) );
  NAND2_X1 U16501 ( .A1(n14671), .A2(n15198), .ZN(n14672) );
  OAI211_X1 U16502 ( .C1(n15178), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        n14705) );
  MUX2_X1 U16503 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14705), .S(n15213), .Z(
        P1_U3547) );
  INV_X1 U16504 ( .A(n14675), .ZN(n14680) );
  AOI21_X1 U16505 ( .B1(n14677), .B2(n15169), .A(n14676), .ZN(n14678) );
  OAI211_X1 U16506 ( .C1(n14680), .C2(n15184), .A(n14679), .B(n14678), .ZN(
        n14706) );
  MUX2_X1 U16507 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14706), .S(n15213), .Z(
        P1_U3546) );
  AOI21_X1 U16508 ( .B1(n14682), .B2(n15169), .A(n14681), .ZN(n14683) );
  OAI211_X1 U16509 ( .C1(n14685), .C2(n15131), .A(n14684), .B(n14683), .ZN(
        n14707) );
  MUX2_X1 U16510 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14707), .S(n15213), .Z(
        P1_U3545) );
  OAI211_X1 U16511 ( .C1(n7105), .C2(n15194), .A(n14688), .B(n14687), .ZN(
        n14689) );
  AOI21_X1 U16512 ( .B1(n14690), .B2(n15198), .A(n14689), .ZN(n14691) );
  OAI21_X1 U16513 ( .B1(n15178), .B2(n14692), .A(n14691), .ZN(n14708) );
  MUX2_X1 U16514 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14708), .S(n15213), .Z(
        P1_U3544) );
  MUX2_X1 U16515 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14693), .S(n15200), .Z(
        P1_U3527) );
  MUX2_X1 U16516 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14694), .S(n15200), .Z(
        P1_U3526) );
  MUX2_X1 U16517 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14696), .S(n15200), .Z(
        P1_U3524) );
  MUX2_X1 U16518 ( .A(n14697), .B(P1_REG0_REG_27__SCAN_IN), .S(n15199), .Z(
        P1_U3523) );
  MUX2_X1 U16519 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14698), .S(n15200), .Z(
        P1_U3522) );
  MUX2_X1 U16520 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14699), .S(n15200), .Z(
        P1_U3521) );
  MUX2_X1 U16521 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14700), .S(n15200), .Z(
        P1_U3520) );
  MUX2_X1 U16522 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14701), .S(n15200), .Z(
        P1_U3519) );
  MUX2_X1 U16523 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14702), .S(n15200), .Z(
        P1_U3518) );
  MUX2_X1 U16524 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14703), .S(n15200), .Z(
        P1_U3517) );
  MUX2_X1 U16525 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14704), .S(n15200), .Z(
        P1_U3516) );
  MUX2_X1 U16526 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14705), .S(n15200), .Z(
        P1_U3515) );
  MUX2_X1 U16527 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14706), .S(n15200), .Z(
        P1_U3513) );
  MUX2_X1 U16528 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14707), .S(n15200), .Z(
        P1_U3510) );
  MUX2_X1 U16529 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14708), .S(n15200), .Z(
        P1_U3507) );
  NOR4_X1 U16530 ( .A1(n14709), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n9447), .ZN(n14710) );
  AOI21_X1 U16531 ( .B1(n14717), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14710), 
        .ZN(n14711) );
  OAI21_X1 U16532 ( .B1(n14712), .B2(n12426), .A(n14711), .ZN(P1_U3324) );
  OAI222_X1 U16533 ( .A1(n12426), .A2(n14715), .B1(n14714), .B2(P1_U3086), 
        .C1(n14713), .C2(n12296), .ZN(P1_U3326) );
  AOI21_X1 U16534 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n14717), .A(n14716), 
        .ZN(n14718) );
  OAI21_X1 U16535 ( .B1(n14719), .B2(n12426), .A(n14718), .ZN(P1_U3328) );
  MUX2_X1 U16536 ( .A(n15133), .B(n14720), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16537 ( .A(n14722), .B(n14721), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  XOR2_X1 U16538 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(P3_ADDR_REG_18__SCAN_IN), 
        .Z(n14867) );
  NOR2_X1 U16539 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14814), .ZN(n14749) );
  INV_X1 U16540 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14879) );
  INV_X1 U16541 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U16542 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15076), .ZN(n14748) );
  NOR2_X1 U16543 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14807), .ZN(n14747) );
  INV_X1 U16544 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14745) );
  INV_X1 U16545 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14739) );
  INV_X1 U16546 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14738) );
  XNOR2_X1 U16547 ( .A(n14725), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14759) );
  NOR2_X1 U16548 ( .A1(n14726), .A2(n15489), .ZN(n14728) );
  NOR2_X1 U16549 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n14769), .ZN(n14727) );
  NOR2_X1 U16550 ( .A1(n14730), .A2(n15525), .ZN(n14732) );
  NOR2_X1 U16551 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14772), .ZN(n14731) );
  XNOR2_X1 U16552 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(n14734), .ZN(n14778) );
  NOR2_X1 U16553 ( .A1(n14779), .A2(n14778), .ZN(n14733) );
  INV_X1 U16554 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14735) );
  XOR2_X1 U16555 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14786) );
  XOR2_X1 U16556 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14756) );
  NOR2_X1 U16557 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14740), .ZN(n14742) );
  XOR2_X1 U16558 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n14796) );
  NOR2_X1 U16559 ( .A1(n14795), .A2(n14796), .ZN(n14743) );
  XOR2_X1 U16560 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14802) );
  NOR2_X1 U16561 ( .A1(n14801), .A2(n14802), .ZN(n14744) );
  AND2_X1 U16562 ( .A1(n15528), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14746) );
  INV_X1 U16563 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15060) );
  OAI22_X1 U16564 ( .A1(n14747), .A2(n14809), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n15060), .ZN(n14810) );
  OAI22_X1 U16565 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14879), .B1(n14748), 
        .B2(n14810), .ZN(n14816) );
  NAND2_X1 U16566 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14814), .ZN(n14813) );
  OAI21_X1 U16567 ( .B1(n14749), .B2(n14816), .A(n14813), .ZN(n14750) );
  NOR2_X1 U16568 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14750), .ZN(n14752) );
  XOR2_X1 U16569 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14750), .Z(n14817) );
  AND2_X1 U16570 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14817), .ZN(n14751) );
  XNOR2_X1 U16571 ( .A(n14867), .B(n14868), .ZN(n14863) );
  INV_X1 U16572 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15296) );
  XOR2_X1 U16573 ( .A(n15528), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14754) );
  XOR2_X1 U16574 ( .A(n14754), .B(n14753), .Z(n14806) );
  INV_X1 U16575 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14794) );
  XNOR2_X1 U16576 ( .A(n14756), .B(n14755), .ZN(n14790) );
  NAND2_X1 U16577 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14758), .ZN(n14771) );
  XNOR2_X1 U16578 ( .A(n14760), .B(n14759), .ZN(n14768) );
  XOR2_X1 U16579 ( .A(n14762), .B(n14761), .Z(n14764) );
  NAND2_X1 U16580 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14764), .ZN(n14766) );
  AOI21_X1 U16581 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14763), .A(n14762), .ZN(
        n15635) );
  NOR2_X1 U16582 ( .A1(n15635), .A2(n10024), .ZN(n15644) );
  NAND2_X1 U16583 ( .A1(n14766), .A2(n14765), .ZN(n14767) );
  NAND2_X1 U16584 ( .A1(n14768), .A2(n14767), .ZN(n14821) );
  NOR2_X1 U16585 ( .A1(n14768), .A2(n14767), .ZN(n14822) );
  XNOR2_X1 U16586 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14769), .ZN(n15640) );
  NOR2_X1 U16587 ( .A1(n15639), .A2(n15640), .ZN(n14770) );
  INV_X1 U16588 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U16589 ( .A1(n15639), .A2(n15640), .ZN(n15638) );
  OAI21_X1 U16590 ( .B1(n14770), .B2(n15641), .A(n15638), .ZN(n15632) );
  XNOR2_X1 U16591 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14772), .ZN(n14773) );
  NOR2_X1 U16592 ( .A1(n14774), .A2(n14773), .ZN(n14776) );
  XNOR2_X1 U16593 ( .A(n14774), .B(n14773), .ZN(n15634) );
  NOR2_X1 U16594 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15634), .ZN(n14775) );
  NAND2_X1 U16595 ( .A1(n14777), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14780) );
  XNOR2_X1 U16596 ( .A(n14779), .B(n14778), .ZN(n14839) );
  NOR2_X1 U16597 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14781), .ZN(n14784) );
  XNOR2_X1 U16598 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n14781), .ZN(n15637) );
  XNOR2_X1 U16599 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14782), .ZN(n15636) );
  NOR2_X1 U16600 ( .A1(n15637), .A2(n15636), .ZN(n14783) );
  XNOR2_X1 U16601 ( .A(n14786), .B(n14785), .ZN(n14788) );
  NAND2_X1 U16602 ( .A1(n14787), .A2(n14788), .ZN(n14789) );
  XOR2_X1 U16603 ( .A(n14793), .B(n14792), .Z(n14847) );
  XNOR2_X1 U16604 ( .A(n14796), .B(n14795), .ZN(n14798) );
  NOR2_X1 U16605 ( .A1(n14797), .A2(n14798), .ZN(n14800) );
  XNOR2_X1 U16606 ( .A(n14798), .B(n14797), .ZN(n15015) );
  NOR2_X1 U16607 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n15015), .ZN(n14799) );
  XNOR2_X1 U16608 ( .A(n14802), .B(n14801), .ZN(n14803) );
  XNOR2_X1 U16609 ( .A(n14807), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14808) );
  XOR2_X1 U16610 ( .A(n14809), .B(n14808), .Z(n15022) );
  XOR2_X1 U16611 ( .A(n14879), .B(P1_ADDR_REG_15__SCAN_IN), .Z(n14811) );
  OAI21_X1 U16612 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14814), .A(n14813), 
        .ZN(n14815) );
  XOR2_X1 U16613 ( .A(n14816), .B(n14815), .Z(n15029) );
  XNOR2_X1 U16614 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14817), .ZN(n14859) );
  XNOR2_X1 U16615 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14862), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16616 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14819) );
  OAI21_X1 U16617 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14819), 
        .ZN(U28) );
  AOI21_X1 U16618 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14820) );
  OAI21_X1 U16619 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14820), 
        .ZN(U29) );
  INV_X1 U16620 ( .A(n14821), .ZN(n14823) );
  AOI222_X1 U16621 ( .A1(n9881), .A2(n14823), .B1(n9881), .B2(n14822), .C1(
        n15639), .C2(n14821), .ZN(SUB_1596_U61) );
  INV_X1 U16622 ( .A(n14824), .ZN(n14825) );
  AOI22_X1 U16623 ( .A1(n14825), .A2(n14835), .B1(SI_4_), .B2(n14834), .ZN(
        n14826) );
  OAI21_X1 U16624 ( .B1(P3_U3151), .B2(n15504), .A(n14826), .ZN(P3_U3291) );
  INV_X1 U16625 ( .A(n14827), .ZN(n14828) );
  AOI22_X1 U16626 ( .A1(n14828), .A2(n14835), .B1(SI_5_), .B2(n14834), .ZN(
        n14829) );
  OAI21_X1 U16627 ( .B1(P3_U3151), .B2(n15512), .A(n14829), .ZN(P3_U3290) );
  AOI22_X1 U16628 ( .A1(n14830), .A2(n14835), .B1(SI_8_), .B2(n14834), .ZN(
        n14831) );
  OAI21_X1 U16629 ( .B1(P3_U3151), .B2(n14832), .A(n14831), .ZN(P3_U3287) );
  INV_X1 U16630 ( .A(n14833), .ZN(n14836) );
  AOI22_X1 U16631 ( .A1(n14836), .A2(n14835), .B1(SI_11_), .B2(n14834), .ZN(
        n14837) );
  OAI21_X1 U16632 ( .B1(P3_U3151), .B2(n14838), .A(n14837), .ZN(P3_U3284) );
  XOR2_X1 U16633 ( .A(n14840), .B(n14839), .Z(SUB_1596_U57) );
  XOR2_X1 U16634 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14841), .Z(SUB_1596_U55) );
  NOR2_X1 U16635 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  XNOR2_X1 U16636 ( .A(n14845), .B(n14844), .ZN(SUB_1596_U54) );
  AOI21_X1 U16637 ( .B1(n14848), .B2(n14847), .A(n14846), .ZN(n14849) );
  XOR2_X1 U16638 ( .A(n14849), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  INV_X1 U16639 ( .A(n14850), .ZN(n14851) );
  OAI21_X1 U16640 ( .B1(n14852), .B2(n15194), .A(n14851), .ZN(n14854) );
  AOI211_X1 U16641 ( .C1(n15157), .C2(n14855), .A(n14854), .B(n14853), .ZN(
        n14858) );
  AOI22_X1 U16642 ( .A1(n15200), .A2(n14858), .B1(n14856), .B2(n15199), .ZN(
        P1_U3495) );
  AOI22_X1 U16643 ( .A1(n15213), .A2(n14858), .B1(n14857), .B2(n15210), .ZN(
        P1_U3540) );
  AOI21_X1 U16644 ( .B1(n14860), .B2(n14859), .A(n6701), .ZN(n14861) );
  XOR2_X1 U16645 ( .A(n14861), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16646 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14862), .ZN(n14866) );
  NOR2_X1 U16647 ( .A1(n14864), .A2(n14863), .ZN(n14865) );
  NOR2_X2 U16648 ( .A1(n14866), .A2(n14865), .ZN(n14875) );
  NOR2_X1 U16649 ( .A1(n14868), .A2(n14867), .ZN(n14869) );
  AOI21_X1 U16650 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14301), .A(n14869), 
        .ZN(n14873) );
  XNOR2_X1 U16651 ( .A(n14870), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14871) );
  XNOR2_X1 U16652 ( .A(n14871), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14872) );
  XNOR2_X1 U16653 ( .A(n14873), .B(n14872), .ZN(n14874) );
  XNOR2_X1 U16654 ( .A(n14875), .B(n14874), .ZN(SUB_1596_U4) );
  AOI21_X1 U16655 ( .B1(n14878), .B2(n14877), .A(n14876), .ZN(n14891) );
  OAI22_X1 U16656 ( .A1(n15531), .A2(n7055), .B1(n15529), .B2(n14879), .ZN(
        n14889) );
  AOI21_X1 U16657 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14887) );
  AOI21_X1 U16658 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14886) );
  OAI22_X1 U16659 ( .A1(n14887), .A2(n14920), .B1(n14886), .B2(n15541), .ZN(
        n14888) );
  AOI211_X1 U16660 ( .C1(P3_REG3_REG_15__SCAN_IN), .C2(P3_U3151), .A(n14889), 
        .B(n14888), .ZN(n14890) );
  OAI21_X1 U16661 ( .B1(n14891), .B2(n15547), .A(n14890), .ZN(P3_U3197) );
  INV_X1 U16662 ( .A(n14892), .ZN(n14893) );
  AOI21_X1 U16663 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14913) );
  NAND2_X1 U16664 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  XNOR2_X1 U16665 ( .A(n14899), .B(n14898), .ZN(n14905) );
  NOR2_X1 U16666 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14900), .ZN(n14901) );
  AOI21_X1 U16667 ( .B1(n15458), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14901), 
        .ZN(n14902) );
  OAI21_X1 U16668 ( .B1(n15531), .B2(n14903), .A(n14902), .ZN(n14904) );
  AOI21_X1 U16669 ( .B1(n14905), .B2(n15538), .A(n14904), .ZN(n14912) );
  INV_X1 U16670 ( .A(n14906), .ZN(n14907) );
  AOI21_X1 U16671 ( .B1(n14909), .B2(n14908), .A(n14907), .ZN(n14910) );
  OR2_X1 U16672 ( .A1(n14910), .A2(n15541), .ZN(n14911) );
  OAI211_X1 U16673 ( .C1(n14913), .C2(n15547), .A(n14912), .B(n14911), .ZN(
        P3_U3198) );
  AOI21_X1 U16674 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14934) );
  INV_X1 U16675 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14918) );
  OAI21_X1 U16676 ( .B1(n15529), .B2(n14918), .A(n14917), .ZN(n14924) );
  AOI211_X1 U16677 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14923) );
  AOI211_X1 U16678 ( .C1(n14926), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        n14933) );
  INV_X1 U16679 ( .A(n14927), .ZN(n14928) );
  NOR2_X1 U16680 ( .A1(n14928), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14931) );
  OAI21_X1 U16681 ( .B1(n14931), .B2(n14930), .A(n14929), .ZN(n14932) );
  OAI211_X1 U16682 ( .C1(n14934), .C2(n15547), .A(n14933), .B(n14932), .ZN(
        P3_U3199) );
  INV_X1 U16683 ( .A(n14935), .ZN(n14937) );
  AOI22_X1 U16684 ( .A1(n14939), .A2(n14938), .B1(n14949), .B2(n15566), .ZN(
        n14946) );
  NOR2_X1 U16685 ( .A1(n15566), .A2(n14940), .ZN(n14941) );
  AOI21_X1 U16686 ( .B1(n14947), .B2(n14944), .A(n14941), .ZN(n14942) );
  NAND2_X1 U16687 ( .A1(n14946), .A2(n14942), .ZN(P3_U3202) );
  AOI22_X1 U16688 ( .A1(n14951), .A2(n14944), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14943), .ZN(n14945) );
  NAND2_X1 U16689 ( .A1(n14946), .A2(n14945), .ZN(P3_U3203) );
  AOI21_X1 U16690 ( .B1(n14947), .B2(n14950), .A(n14949), .ZN(n14953) );
  INV_X1 U16691 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U16692 ( .A1(n15631), .A2(n14953), .B1(n14948), .B2(n15628), .ZN(
        P3_U3490) );
  AOI21_X1 U16693 ( .B1(n14951), .B2(n14950), .A(n14949), .ZN(n14954) );
  INV_X1 U16694 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U16695 ( .A1(n15631), .A2(n14954), .B1(n14952), .B2(n15628), .ZN(
        P3_U3489) );
  AOI22_X1 U16696 ( .A1(n15613), .A2(n14953), .B1(n11638), .B2(n15612), .ZN(
        P3_U3458) );
  AOI22_X1 U16697 ( .A1(n15613), .A2(n14954), .B1(n9300), .B2(n15612), .ZN(
        P3_U3457) );
  AOI22_X1 U16698 ( .A1(n15316), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n15315), 
        .B2(n14955), .ZN(n14956) );
  OAI21_X1 U16699 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14962) );
  NOR2_X1 U16700 ( .A1(n14960), .A2(n14959), .ZN(n14961) );
  AOI211_X1 U16701 ( .C1(n14963), .C2(n15326), .A(n14962), .B(n14961), .ZN(
        n14964) );
  OAI21_X1 U16702 ( .B1(n15316), .B2(n14965), .A(n14964), .ZN(P2_U3250) );
  OAI21_X1 U16703 ( .B1(n14967), .B2(n15428), .A(n14966), .ZN(n14970) );
  INV_X1 U16704 ( .A(n14968), .ZN(n14969) );
  AOI211_X1 U16705 ( .C1(n14971), .C2(n15379), .A(n14970), .B(n14969), .ZN(
        n14979) );
  AOI22_X1 U16706 ( .A1(n15457), .A2(n14979), .B1(n11016), .B2(n15455), .ZN(
        P2_U3513) );
  INV_X1 U16707 ( .A(n15438), .ZN(n15432) );
  INV_X1 U16708 ( .A(n14972), .ZN(n14977) );
  OAI21_X1 U16709 ( .B1(n14974), .B2(n15428), .A(n14973), .ZN(n14976) );
  AOI211_X1 U16710 ( .C1(n15432), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n14980) );
  AOI22_X1 U16711 ( .A1(n15457), .A2(n14980), .B1(n15256), .B2(n15455), .ZN(
        P2_U3511) );
  INV_X1 U16712 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16713 ( .A1(n15444), .A2(n14979), .B1(n14978), .B2(n15442), .ZN(
        P2_U3472) );
  AOI22_X1 U16714 ( .A1(n15444), .A2(n14980), .B1(n8609), .B2(n15442), .ZN(
        P2_U3466) );
  OAI22_X1 U16715 ( .A1(n14984), .A2(n14983), .B1(n14982), .B2(n14981), .ZN(
        n14993) );
  AOI21_X1 U16716 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14988) );
  INV_X1 U16717 ( .A(n14988), .ZN(n14991) );
  AOI21_X1 U16718 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(n14992) );
  AOI211_X1 U16719 ( .C1(n14995), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14996) );
  NAND2_X1 U16720 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15058)
         );
  OAI211_X1 U16721 ( .C1(n14998), .C2(n14997), .A(n14996), .B(n15058), .ZN(
        P1_U3215) );
  OAI21_X1 U16722 ( .B1(n15000), .B2(n15194), .A(n14999), .ZN(n15002) );
  AOI211_X1 U16723 ( .C1(n15198), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        n15012) );
  AOI22_X1 U16724 ( .A1(n15213), .A2(n15012), .B1(n11173), .B2(n15210), .ZN(
        P1_U3541) );
  AOI21_X1 U16725 ( .B1(n15005), .B2(n15169), .A(n15004), .ZN(n15006) );
  OAI21_X1 U16726 ( .B1(n15007), .B2(n15131), .A(n15006), .ZN(n15008) );
  NOR2_X1 U16727 ( .A1(n15009), .A2(n15008), .ZN(n15014) );
  AOI22_X1 U16728 ( .A1(n15213), .A2(n15014), .B1(n15010), .B2(n15210), .ZN(
        P1_U3539) );
  INV_X1 U16729 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U16730 ( .A1(n15200), .A2(n15012), .B1(n15011), .B2(n15199), .ZN(
        P1_U3498) );
  INV_X1 U16731 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16732 ( .A1(n15200), .A2(n15014), .B1(n15013), .B2(n15199), .ZN(
        P1_U3492) );
  XNOR2_X1 U16733 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15015), .ZN(SUB_1596_U69)
         );
  INV_X1 U16734 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15271) );
  XOR2_X1 U16735 ( .A(n15271), .B(n15016), .Z(SUB_1596_U68) );
  NOR2_X1 U16736 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  XOR2_X1 U16737 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n15019), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16738 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15023) );
  XOR2_X1 U16739 ( .A(n15023), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16740 ( .A1(n15025), .A2(n15024), .ZN(n15026) );
  XOR2_X1 U16741 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15026), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16742 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15030) );
  XOR2_X1 U16743 ( .A(n15030), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16744 ( .B1(n15032), .B2(n15031), .A(n15070), .ZN(n15040) );
  AND2_X1 U16745 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  OAI21_X1 U16746 ( .B1(n15036), .B2(n15035), .A(n15071), .ZN(n15039) );
  NAND2_X1 U16747 ( .A1(n15067), .A2(n15037), .ZN(n15038) );
  OAI211_X1 U16748 ( .C1(n15041), .C2(n15040), .A(n15039), .B(n15038), .ZN(
        n15042) );
  INV_X1 U16749 ( .A(n15042), .ZN(n15044) );
  OAI211_X1 U16750 ( .C1(n15045), .C2(n15075), .A(n15044), .B(n15043), .ZN(
        P1_U3254) );
  AOI211_X1 U16751 ( .C1(n15049), .C2(n15048), .A(n15047), .B(n15046), .ZN(
        n15056) );
  AOI21_X1 U16752 ( .B1(n15052), .B2(n15051), .A(n15050), .ZN(n15054) );
  NOR2_X1 U16753 ( .A1(n15054), .A2(n15053), .ZN(n15055) );
  AOI211_X1 U16754 ( .C1(n15067), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15059) );
  OAI211_X1 U16755 ( .C1(n15060), .C2(n15075), .A(n15059), .B(n15058), .ZN(
        P1_U3257) );
  AOI21_X1 U16756 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n15062), .A(n15061), 
        .ZN(n15063) );
  INV_X1 U16757 ( .A(n15063), .ZN(n15072) );
  OAI21_X1 U16758 ( .B1(n15066), .B2(n15065), .A(n15064), .ZN(n15069) );
  AOI222_X1 U16759 ( .A1(n15072), .A2(n15071), .B1(n15070), .B2(n15069), .C1(
        n15068), .C2(n15067), .ZN(n15074) );
  OAI211_X1 U16760 ( .C1(n15076), .C2(n15075), .A(n15074), .B(n15073), .ZN(
        P1_U3258) );
  XNOR2_X1 U16761 ( .A(n15078), .B(n15077), .ZN(n15152) );
  XNOR2_X1 U16762 ( .A(n15080), .B(n15079), .ZN(n15082) );
  OAI21_X1 U16763 ( .B1(n15082), .B2(n15178), .A(n15081), .ZN(n15083) );
  AOI21_X1 U16764 ( .B1(n15152), .B2(n15084), .A(n15083), .ZN(n15149) );
  AOI22_X1 U16765 ( .A1(n15086), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15085), .ZN(n15087) );
  OAI21_X1 U16766 ( .B1(n15088), .B2(n15148), .A(n15087), .ZN(n15089) );
  INV_X1 U16767 ( .A(n15089), .ZN(n15097) );
  AOI211_X1 U16768 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15146) );
  AOI22_X1 U16769 ( .A1(n15095), .A2(n15152), .B1(n15094), .B2(n15146), .ZN(
        n15096) );
  OAI211_X1 U16770 ( .C1(n15098), .C2(n15149), .A(n15097), .B(n15096), .ZN(
        P1_U3291) );
  NOR2_X1 U16771 ( .A1(n15129), .A2(n15099), .ZN(P1_U3294) );
  INV_X1 U16772 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15100) );
  NOR2_X1 U16773 ( .A1(n15129), .A2(n15100), .ZN(P1_U3295) );
  NOR2_X1 U16774 ( .A1(n15129), .A2(n15101), .ZN(P1_U3296) );
  NOR2_X1 U16775 ( .A1(n15129), .A2(n15102), .ZN(P1_U3297) );
  INV_X1 U16776 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15103) );
  NOR2_X1 U16777 ( .A1(n15129), .A2(n15103), .ZN(P1_U3298) );
  INV_X1 U16778 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15104) );
  NOR2_X1 U16779 ( .A1(n15129), .A2(n15104), .ZN(P1_U3299) );
  INV_X1 U16780 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15105) );
  NOR2_X1 U16781 ( .A1(n15129), .A2(n15105), .ZN(P1_U3300) );
  INV_X1 U16782 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15106) );
  NOR2_X1 U16783 ( .A1(n15129), .A2(n15106), .ZN(P1_U3301) );
  INV_X1 U16784 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U16785 ( .A1(n15129), .A2(n15107), .ZN(P1_U3302) );
  INV_X1 U16786 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U16787 ( .A1(n15129), .A2(n15108), .ZN(P1_U3303) );
  NOR2_X1 U16788 ( .A1(n15129), .A2(n15109), .ZN(P1_U3304) );
  INV_X1 U16789 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15110) );
  NOR2_X1 U16790 ( .A1(n15129), .A2(n15110), .ZN(P1_U3305) );
  NOR2_X1 U16791 ( .A1(n15129), .A2(n15111), .ZN(P1_U3306) );
  INV_X1 U16792 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15112) );
  NOR2_X1 U16793 ( .A1(n15129), .A2(n15112), .ZN(P1_U3307) );
  INV_X1 U16794 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U16795 ( .A1(n15129), .A2(n15113), .ZN(P1_U3308) );
  INV_X1 U16796 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15114) );
  NOR2_X1 U16797 ( .A1(n15129), .A2(n15114), .ZN(P1_U3309) );
  INV_X1 U16798 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16799 ( .A1(n15129), .A2(n15115), .ZN(P1_U3310) );
  NOR2_X1 U16800 ( .A1(n15129), .A2(n15116), .ZN(P1_U3311) );
  INV_X1 U16801 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U16802 ( .A1(n15129), .A2(n15117), .ZN(P1_U3312) );
  INV_X1 U16803 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U16804 ( .A1(n15129), .A2(n15118), .ZN(P1_U3313) );
  INV_X1 U16805 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15119) );
  NOR2_X1 U16806 ( .A1(n15129), .A2(n15119), .ZN(P1_U3314) );
  INV_X1 U16807 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U16808 ( .A1(n15129), .A2(n15120), .ZN(P1_U3315) );
  INV_X1 U16809 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16810 ( .A1(n15129), .A2(n15121), .ZN(P1_U3316) );
  INV_X1 U16811 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U16812 ( .A1(n15129), .A2(n15122), .ZN(P1_U3317) );
  INV_X1 U16813 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U16814 ( .A1(n15129), .A2(n15123), .ZN(P1_U3318) );
  INV_X1 U16815 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16816 ( .A1(n15129), .A2(n15124), .ZN(P1_U3319) );
  NOR2_X1 U16817 ( .A1(n15129), .A2(n15125), .ZN(P1_U3320) );
  INV_X1 U16818 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15126) );
  NOR2_X1 U16819 ( .A1(n15129), .A2(n15126), .ZN(P1_U3321) );
  INV_X1 U16820 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16821 ( .A1(n15129), .A2(n15127), .ZN(P1_U3322) );
  INV_X1 U16822 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15128) );
  NOR2_X1 U16823 ( .A1(n15129), .A2(n15128), .ZN(P1_U3323) );
  AOI21_X1 U16824 ( .B1(n15178), .B2(n15131), .A(n15130), .ZN(n15138) );
  INV_X1 U16825 ( .A(n15132), .ZN(n15137) );
  NOR3_X1 U16826 ( .A1(n15135), .A2(n15134), .A3(n15133), .ZN(n15136) );
  NOR3_X1 U16827 ( .A1(n15138), .A2(n15137), .A3(n15136), .ZN(n15201) );
  AOI22_X1 U16828 ( .A1(n15200), .A2(n15201), .B1(n15139), .B2(n15199), .ZN(
        P1_U3459) );
  INV_X1 U16829 ( .A(n15140), .ZN(n15145) );
  OAI21_X1 U16830 ( .B1(n6575), .B2(n15194), .A(n15141), .ZN(n15144) );
  INV_X1 U16831 ( .A(n15142), .ZN(n15143) );
  AOI211_X1 U16832 ( .C1(n15198), .C2(n15145), .A(n15144), .B(n15143), .ZN(
        n15202) );
  AOI22_X1 U16833 ( .A1(n15200), .A2(n15202), .B1(n9453), .B2(n15199), .ZN(
        P1_U3462) );
  INV_X1 U16834 ( .A(n15146), .ZN(n15147) );
  OAI21_X1 U16835 ( .B1(n15148), .B2(n15194), .A(n15147), .ZN(n15151) );
  INV_X1 U16836 ( .A(n15149), .ZN(n15150) );
  AOI211_X1 U16837 ( .C1(n15157), .C2(n15152), .A(n15151), .B(n15150), .ZN(
        n15203) );
  INV_X1 U16838 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16839 ( .A1(n15200), .A2(n15203), .B1(n15153), .B2(n15199), .ZN(
        P1_U3465) );
  OAI21_X1 U16840 ( .B1(n15155), .B2(n15194), .A(n15154), .ZN(n15156) );
  AOI21_X1 U16841 ( .B1(n15158), .B2(n15157), .A(n15156), .ZN(n15159) );
  AND2_X1 U16842 ( .A1(n15160), .A2(n15159), .ZN(n15204) );
  INV_X1 U16843 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16844 ( .A1(n15200), .A2(n15204), .B1(n15161), .B2(n15199), .ZN(
        P1_U3468) );
  OAI21_X1 U16845 ( .B1(n7090), .B2(n15194), .A(n15162), .ZN(n15164) );
  AOI211_X1 U16846 ( .C1(n15198), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        n15205) );
  INV_X1 U16847 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U16848 ( .A1(n15200), .A2(n15205), .B1(n15166), .B2(n15199), .ZN(
        P1_U3477) );
  INV_X1 U16849 ( .A(n15167), .ZN(n15172) );
  AOI21_X1 U16850 ( .B1(n15170), .B2(n15169), .A(n15168), .ZN(n15171) );
  OAI21_X1 U16851 ( .B1(n15172), .B2(n15184), .A(n15171), .ZN(n15173) );
  NOR2_X1 U16852 ( .A1(n15174), .A2(n15173), .ZN(n15206) );
  AOI22_X1 U16853 ( .A1(n15200), .A2(n15206), .B1(n10463), .B2(n15199), .ZN(
        P1_U3480) );
  OAI211_X1 U16854 ( .C1(n15177), .C2(n15194), .A(n15176), .B(n15175), .ZN(
        n15181) );
  NOR2_X1 U16855 ( .A1(n15179), .A2(n15178), .ZN(n15180) );
  AOI211_X1 U16856 ( .C1(n15198), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15207) );
  INV_X1 U16857 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16858 ( .A1(n15200), .A2(n15207), .B1(n15183), .B2(n15199), .ZN(
        P1_U3483) );
  NOR2_X1 U16859 ( .A1(n15185), .A2(n15184), .ZN(n15188) );
  NOR4_X1 U16860 ( .A1(n15189), .A2(n15188), .A3(n15187), .A4(n15186), .ZN(
        n15209) );
  INV_X1 U16861 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U16862 ( .A1(n15200), .A2(n15209), .B1(n15190), .B2(n15199), .ZN(
        P1_U3486) );
  INV_X1 U16863 ( .A(n15191), .ZN(n15195) );
  OAI211_X1 U16864 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15196) );
  AOI21_X1 U16865 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15212) );
  AOI22_X1 U16866 ( .A1(n15200), .A2(n15212), .B1(n10809), .B2(n15199), .ZN(
        P1_U3489) );
  AOI22_X1 U16867 ( .A1(n15213), .A2(n15201), .B1(n9468), .B2(n15210), .ZN(
        P1_U3528) );
  AOI22_X1 U16868 ( .A1(n15213), .A2(n15202), .B1(n9760), .B2(n15210), .ZN(
        P1_U3529) );
  AOI22_X1 U16869 ( .A1(n15213), .A2(n15203), .B1(n9763), .B2(n15210), .ZN(
        P1_U3530) );
  AOI22_X1 U16870 ( .A1(n15213), .A2(n15204), .B1(n9759), .B2(n15210), .ZN(
        P1_U3531) );
  AOI22_X1 U16871 ( .A1(n15213), .A2(n15205), .B1(n9774), .B2(n15210), .ZN(
        P1_U3534) );
  AOI22_X1 U16872 ( .A1(n15213), .A2(n15206), .B1(n9775), .B2(n15210), .ZN(
        P1_U3535) );
  AOI22_X1 U16873 ( .A1(n15213), .A2(n15207), .B1(n10499), .B2(n15210), .ZN(
        P1_U3536) );
  AOI22_X1 U16874 ( .A1(n15213), .A2(n15209), .B1(n15208), .B2(n15210), .ZN(
        P1_U3537) );
  AOI22_X1 U16875 ( .A1(n15213), .A2(n15212), .B1(n15211), .B2(n15210), .ZN(
        P1_U3538) );
  NOR2_X1 U16876 ( .A1(n15298), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16877 ( .A(n15214), .ZN(n15217) );
  OAI22_X1 U16878 ( .A1(n15217), .A2(n15216), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15215), .ZN(n15222) );
  AOI211_X1 U16879 ( .C1(n15220), .C2(n15219), .A(n13480), .B(n15218), .ZN(
        n15221) );
  AOI211_X1 U16880 ( .C1(n15224), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15225) );
  OAI21_X1 U16881 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n15226), .A(n15225), .ZN(
        P2_U3190) );
  INV_X1 U16882 ( .A(n15227), .ZN(n15242) );
  OAI21_X1 U16883 ( .B1(n15242), .B2(n15228), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15229) );
  OAI21_X1 U16884 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15229), .ZN(n15240) );
  INV_X1 U16885 ( .A(n15230), .ZN(n15233) );
  OAI21_X1 U16886 ( .B1(n10020), .B2(n7308), .A(n15231), .ZN(n15232) );
  NAND3_X1 U16887 ( .A1(n15305), .A2(n15233), .A3(n15232), .ZN(n15239) );
  NAND2_X1 U16888 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15298), .ZN(n15238) );
  AND2_X1 U16889 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15235) );
  OAI211_X1 U16890 ( .C1(n15236), .C2(n15235), .A(n15302), .B(n15234), .ZN(
        n15237) );
  NAND4_X1 U16891 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        P2_U3215) );
  OAI21_X1 U16892 ( .B1(n15242), .B2(n15241), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15243) );
  OAI21_X1 U16893 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15243), .ZN(n15254) );
  OAI211_X1 U16894 ( .C1(n15246), .C2(n15245), .A(n15244), .B(n15305), .ZN(
        n15253) );
  AOI211_X1 U16895 ( .C1(n15249), .C2(n15248), .A(n15263), .B(n15247), .ZN(
        n15250) );
  INV_X1 U16896 ( .A(n15250), .ZN(n15252) );
  NAND2_X1 U16897 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n15298), .ZN(n15251) );
  NAND4_X1 U16898 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        P2_U3220) );
  NOR2_X1 U16899 ( .A1(n15268), .A2(n15256), .ZN(n15255) );
  AOI21_X1 U16900 ( .B1(n15256), .B2(n15268), .A(n15255), .ZN(n15259) );
  AOI21_X1 U16901 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n15266) );
  AOI21_X1 U16902 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15264) );
  OAI22_X1 U16903 ( .A1(n15266), .A2(n15265), .B1(n15264), .B2(n15263), .ZN(
        n15267) );
  AOI21_X1 U16904 ( .B1(n15268), .B2(n15300), .A(n15267), .ZN(n15270) );
  OAI211_X1 U16905 ( .C1(n15271), .C2(n15297), .A(n15270), .B(n15269), .ZN(
        P2_U3226) );
  OAI21_X1 U16906 ( .B1(n15290), .B2(n15273), .A(n15272), .ZN(n15274) );
  AOI21_X1 U16907 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n15298), .A(n15274), 
        .ZN(n15283) );
  OAI211_X1 U16908 ( .C1(n15277), .C2(n15276), .A(n15302), .B(n15275), .ZN(
        n15282) );
  OAI211_X1 U16909 ( .C1(n15280), .C2(n15279), .A(n15305), .B(n15278), .ZN(
        n15281) );
  NAND3_X1 U16910 ( .A1(n15283), .A2(n15282), .A3(n15281), .ZN(P2_U3227) );
  OAI211_X1 U16911 ( .C1(n15286), .C2(n15285), .A(n15305), .B(n15284), .ZN(
        n15287) );
  OAI211_X1 U16912 ( .C1(n15290), .C2(n15289), .A(n15288), .B(n15287), .ZN(
        n15291) );
  INV_X1 U16913 ( .A(n15291), .ZN(n15295) );
  OAI211_X1 U16914 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n15293), .A(n15302), 
        .B(n15292), .ZN(n15294) );
  OAI211_X1 U16915 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        P2_U3228) );
  AOI22_X1 U16916 ( .A1(n15298), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15310) );
  NAND2_X1 U16917 ( .A1(n15300), .A2(n15299), .ZN(n15309) );
  OAI211_X1 U16918 ( .C1(n15303), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15302), 
        .B(n15301), .ZN(n15308) );
  OAI211_X1 U16919 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15306), .A(n15305), 
        .B(n15304), .ZN(n15307) );
  NAND4_X1 U16920 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        P2_U3229) );
  AOI21_X1 U16921 ( .B1(n15314), .B2(n15313), .A(n15312), .ZN(n15376) );
  AOI222_X1 U16922 ( .A1(n15318), .A2(n15317), .B1(P2_REG2_REG_2__SCAN_IN), 
        .B2(n15316), .C1(n15315), .C2(P2_REG3_REG_2__SCAN_IN), .ZN(n15329) );
  XNOR2_X1 U16923 ( .A(n15320), .B(n15319), .ZN(n15380) );
  INV_X1 U16924 ( .A(n15321), .ZN(n15324) );
  OAI211_X1 U16925 ( .C1(n15324), .C2(n7258), .A(n15323), .B(n15322), .ZN(
        n15375) );
  INV_X1 U16926 ( .A(n15375), .ZN(n15325) );
  AOI22_X1 U16927 ( .A1(n15380), .A2(n15327), .B1(n15326), .B2(n15325), .ZN(
        n15328) );
  OAI211_X1 U16928 ( .C1(n15316), .C2(n15376), .A(n15329), .B(n15328), .ZN(
        P2_U3263) );
  NOR2_X4 U16929 ( .A1(n15330), .A2(n15364), .ZN(n15358) );
  NOR2_X1 U16930 ( .A1(n15358), .A2(n15331), .ZN(P2_U3266) );
  INV_X1 U16931 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U16932 ( .A1(n15358), .A2(n15332), .ZN(P2_U3267) );
  INV_X1 U16933 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16934 ( .A1(n15358), .A2(n15333), .ZN(P2_U3268) );
  NOR2_X1 U16935 ( .A1(n15358), .A2(n15334), .ZN(P2_U3269) );
  INV_X1 U16936 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16937 ( .A1(n15358), .A2(n15335), .ZN(P2_U3270) );
  INV_X1 U16938 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U16939 ( .A1(n15358), .A2(n15336), .ZN(P2_U3271) );
  INV_X1 U16940 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16941 ( .A1(n15358), .A2(n15337), .ZN(P2_U3272) );
  NOR2_X1 U16942 ( .A1(n15358), .A2(n15338), .ZN(P2_U3273) );
  INV_X1 U16943 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16944 ( .A1(n15358), .A2(n15339), .ZN(P2_U3274) );
  INV_X1 U16945 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U16946 ( .A1(n15358), .A2(n15340), .ZN(P2_U3275) );
  INV_X1 U16947 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U16948 ( .A1(n15358), .A2(n15341), .ZN(P2_U3276) );
  INV_X1 U16949 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U16950 ( .A1(n15358), .A2(n15342), .ZN(P2_U3277) );
  INV_X1 U16951 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16952 ( .A1(n15358), .A2(n15343), .ZN(P2_U3278) );
  INV_X1 U16953 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15344) );
  NOR2_X1 U16954 ( .A1(n15358), .A2(n15344), .ZN(P2_U3279) );
  INV_X1 U16955 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15345) );
  NOR2_X1 U16956 ( .A1(n15358), .A2(n15345), .ZN(P2_U3280) );
  INV_X1 U16957 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15346) );
  NOR2_X1 U16958 ( .A1(n15358), .A2(n15346), .ZN(P2_U3281) );
  INV_X1 U16959 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16960 ( .A1(n15358), .A2(n15347), .ZN(P2_U3282) );
  INV_X1 U16961 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U16962 ( .A1(n15358), .A2(n15348), .ZN(P2_U3283) );
  INV_X1 U16963 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16964 ( .A1(n15358), .A2(n15349), .ZN(P2_U3284) );
  INV_X1 U16965 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U16966 ( .A1(n15358), .A2(n15350), .ZN(P2_U3285) );
  INV_X1 U16967 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U16968 ( .A1(n15358), .A2(n15351), .ZN(P2_U3286) );
  INV_X1 U16969 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16970 ( .A1(n15358), .A2(n15352), .ZN(P2_U3287) );
  INV_X1 U16971 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15353) );
  NOR2_X1 U16972 ( .A1(n15358), .A2(n15353), .ZN(P2_U3288) );
  INV_X1 U16973 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U16974 ( .A1(n15358), .A2(n15354), .ZN(P2_U3289) );
  NOR2_X1 U16975 ( .A1(n15358), .A2(n15355), .ZN(P2_U3290) );
  INV_X1 U16976 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15356) );
  NOR2_X1 U16977 ( .A1(n15358), .A2(n15356), .ZN(P2_U3291) );
  INV_X1 U16978 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U16979 ( .A1(n15358), .A2(n15357), .ZN(P2_U3292) );
  INV_X1 U16980 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15359) );
  NOR2_X1 U16981 ( .A1(n15358), .A2(n15359), .ZN(P2_U3293) );
  INV_X1 U16982 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15360) );
  NOR2_X1 U16983 ( .A1(n15358), .A2(n15360), .ZN(P2_U3294) );
  INV_X1 U16984 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15361) );
  NOR2_X1 U16985 ( .A1(n15358), .A2(n15361), .ZN(P2_U3295) );
  AOI22_X1 U16986 ( .A1(n15367), .A2(n15363), .B1(n15362), .B2(n15364), .ZN(
        P2_U3416) );
  AOI22_X1 U16987 ( .A1(n15367), .A2(n15366), .B1(n15365), .B2(n15364), .ZN(
        P2_U3417) );
  OAI21_X1 U16988 ( .B1(n15369), .B2(n15438), .A(n15368), .ZN(n15370) );
  NOR2_X1 U16989 ( .A1(n15371), .A2(n15370), .ZN(n15445) );
  INV_X1 U16990 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U16991 ( .A1(n15444), .A2(n15445), .B1(n15372), .B2(n15442), .ZN(
        P2_U3430) );
  AOI22_X1 U16992 ( .A1(n15444), .A2(n15374), .B1(n15373), .B2(n15442), .ZN(
        P2_U3433) );
  OAI21_X1 U16993 ( .B1(n7258), .B2(n15428), .A(n15375), .ZN(n15378) );
  INV_X1 U16994 ( .A(n15376), .ZN(n15377) );
  AOI211_X1 U16995 ( .C1(n15380), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15446) );
  INV_X1 U16996 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15381) );
  AOI22_X1 U16997 ( .A1(n15444), .A2(n15446), .B1(n15381), .B2(n15442), .ZN(
        P2_U3436) );
  AOI21_X1 U16998 ( .B1(n15434), .B2(n15383), .A(n15382), .ZN(n15384) );
  OAI211_X1 U16999 ( .C1(n15407), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15387) );
  INV_X1 U17000 ( .A(n15387), .ZN(n15447) );
  INV_X1 U17001 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U17002 ( .A1(n15444), .A2(n15447), .B1(n15388), .B2(n15442), .ZN(
        P2_U3442) );
  AOI21_X1 U17003 ( .B1(n15434), .B2(n15390), .A(n15389), .ZN(n15392) );
  OAI211_X1 U17004 ( .C1(n15393), .C2(n15407), .A(n15392), .B(n15391), .ZN(
        n15394) );
  INV_X1 U17005 ( .A(n15394), .ZN(n15448) );
  INV_X1 U17006 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U17007 ( .A1(n15444), .A2(n15448), .B1(n15395), .B2(n15442), .ZN(
        P2_U3445) );
  AND2_X1 U17008 ( .A1(n15396), .A2(n15434), .ZN(n15397) );
  OR2_X1 U17009 ( .A1(n15398), .A2(n15397), .ZN(n15399) );
  AOI21_X1 U17010 ( .B1(n15400), .B2(n15432), .A(n15399), .ZN(n15401) );
  AND2_X1 U17011 ( .A1(n15402), .A2(n15401), .ZN(n15449) );
  INV_X1 U17012 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U17013 ( .A1(n15444), .A2(n15449), .B1(n15403), .B2(n15442), .ZN(
        P2_U3448) );
  AND2_X1 U17014 ( .A1(n15404), .A2(n15434), .ZN(n15405) );
  NOR2_X1 U17015 ( .A1(n15406), .A2(n15405), .ZN(n15410) );
  OR2_X1 U17016 ( .A1(n15408), .A2(n15407), .ZN(n15409) );
  INV_X1 U17017 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U17018 ( .A1(n15444), .A2(n15450), .B1(n15412), .B2(n15442), .ZN(
        P2_U3451) );
  INV_X1 U17019 ( .A(n15413), .ZN(n15418) );
  OAI21_X1 U17020 ( .B1(n15415), .B2(n15428), .A(n15414), .ZN(n15417) );
  AOI211_X1 U17021 ( .C1(n15432), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15451) );
  INV_X1 U17022 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U17023 ( .A1(n15444), .A2(n15451), .B1(n15419), .B2(n15442), .ZN(
        P2_U3454) );
  INV_X1 U17024 ( .A(n15420), .ZN(n15425) );
  OAI21_X1 U17025 ( .B1(n15422), .B2(n15428), .A(n15421), .ZN(n15424) );
  AOI211_X1 U17026 ( .C1(n15432), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15453) );
  AOI22_X1 U17027 ( .A1(n15444), .A2(n15453), .B1(n8559), .B2(n15442), .ZN(
        P2_U3457) );
  INV_X1 U17028 ( .A(n15426), .ZN(n15431) );
  OAI21_X1 U17029 ( .B1(n8918), .B2(n15428), .A(n15427), .ZN(n15430) );
  AOI211_X1 U17030 ( .C1(n15432), .C2(n15431), .A(n15430), .B(n15429), .ZN(
        n15454) );
  INV_X1 U17031 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U17032 ( .A1(n15444), .A2(n15454), .B1(n15433), .B2(n15442), .ZN(
        P2_U3460) );
  NAND2_X1 U17033 ( .A1(n15435), .A2(n15434), .ZN(n15436) );
  OAI211_X1 U17034 ( .C1(n15439), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        n15440) );
  NOR2_X1 U17035 ( .A1(n15441), .A2(n15440), .ZN(n15456) );
  INV_X1 U17036 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15443) );
  AOI22_X1 U17037 ( .A1(n15444), .A2(n15456), .B1(n15443), .B2(n15442), .ZN(
        P2_U3463) );
  AOI22_X1 U17038 ( .A1(n15457), .A2(n15445), .B1(n10020), .B2(n15455), .ZN(
        P2_U3499) );
  AOI22_X1 U17039 ( .A1(n15457), .A2(n15446), .B1(n9833), .B2(n15455), .ZN(
        P2_U3501) );
  AOI22_X1 U17040 ( .A1(n15457), .A2(n15447), .B1(n9837), .B2(n15455), .ZN(
        P2_U3503) );
  AOI22_X1 U17041 ( .A1(n15457), .A2(n15448), .B1(n9838), .B2(n15455), .ZN(
        P2_U3504) );
  AOI22_X1 U17042 ( .A1(n15457), .A2(n15449), .B1(n9839), .B2(n15455), .ZN(
        P2_U3505) );
  AOI22_X1 U17043 ( .A1(n15457), .A2(n15450), .B1(n8527), .B2(n15455), .ZN(
        P2_U3506) );
  AOI22_X1 U17044 ( .A1(n15457), .A2(n15451), .B1(n8545), .B2(n15455), .ZN(
        P2_U3507) );
  AOI22_X1 U17045 ( .A1(n15457), .A2(n15453), .B1(n15452), .B2(n15455), .ZN(
        P2_U3508) );
  AOI22_X1 U17046 ( .A1(n15457), .A2(n15454), .B1(n8578), .B2(n15455), .ZN(
        P2_U3509) );
  AOI22_X1 U17047 ( .A1(n15457), .A2(n15456), .B1(n11020), .B2(n15455), .ZN(
        P2_U3510) );
  NOR2_X1 U17048 ( .A1(P3_U3897), .A2(n15458), .ZN(P3_U3150) );
  XNOR2_X1 U17049 ( .A(n15460), .B(n15459), .ZN(n15470) );
  INV_X1 U17050 ( .A(n15461), .ZN(n15562) );
  AOI22_X1 U17051 ( .A1(n15465), .A2(n6800), .B1(n15463), .B2(n15462), .ZN(
        n15466) );
  OAI21_X1 U17052 ( .B1(n15562), .B2(n15467), .A(n15466), .ZN(n15468) );
  AOI21_X1 U17053 ( .B1(n15470), .B2(n15469), .A(n15468), .ZN(n15471) );
  OAI21_X1 U17054 ( .B1(n15472), .B2(n10136), .A(n15471), .ZN(P3_U3177) );
  AOI21_X1 U17055 ( .B1(n15474), .B2(n7780), .A(n15473), .ZN(n15478) );
  AOI21_X1 U17056 ( .B1(n15476), .B2(n15618), .A(n15475), .ZN(n15477) );
  OAI22_X1 U17057 ( .A1(n15478), .A2(n15547), .B1(n15541), .B2(n15477), .ZN(
        n15479) );
  INV_X1 U17058 ( .A(n15479), .ZN(n15484) );
  XNOR2_X1 U17059 ( .A(n15481), .B(n15480), .ZN(n15482) );
  NAND2_X1 U17060 ( .A1(n15482), .A2(n15538), .ZN(n15483) );
  OAI211_X1 U17061 ( .C1(n15531), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15486) );
  INV_X1 U17062 ( .A(n15486), .ZN(n15488) );
  NAND2_X1 U17063 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n15487) );
  OAI211_X1 U17064 ( .C1(n15489), .C2(n15529), .A(n15488), .B(n15487), .ZN(
        P3_U3185) );
  XNOR2_X1 U17065 ( .A(n15491), .B(n15490), .ZN(n15492) );
  NAND2_X1 U17066 ( .A1(n15492), .A2(n15538), .ZN(n15503) );
  AOI21_X1 U17067 ( .B1(n15495), .B2(n15494), .A(n15493), .ZN(n15500) );
  AOI21_X1 U17068 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15499) );
  OAI22_X1 U17069 ( .A1(n15500), .A2(n15547), .B1(n15541), .B2(n15499), .ZN(
        n15501) );
  INV_X1 U17070 ( .A(n15501), .ZN(n15502) );
  OAI211_X1 U17071 ( .C1(n15531), .C2(n15504), .A(n15503), .B(n15502), .ZN(
        n15505) );
  INV_X1 U17072 ( .A(n15505), .ZN(n15507) );
  NAND2_X1 U17073 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15506) );
  OAI211_X1 U17074 ( .C1(n7413), .C2(n15529), .A(n15507), .B(n15506), .ZN(
        P3_U3186) );
  NAND2_X1 U17075 ( .A1(n15509), .A2(n15508), .ZN(n15511) );
  XOR2_X1 U17076 ( .A(n15511), .B(n15510), .Z(n15522) );
  NOR2_X1 U17077 ( .A1(n15531), .A2(n15512), .ZN(n15521) );
  AOI21_X1 U17078 ( .B1(n15515), .B2(n15514), .A(n15513), .ZN(n15519) );
  AOI21_X1 U17079 ( .B1(n15622), .B2(n15517), .A(n15516), .ZN(n15518) );
  OAI22_X1 U17080 ( .A1(n15519), .A2(n15547), .B1(n15541), .B2(n15518), .ZN(
        n15520) );
  AOI211_X1 U17081 ( .C1(n15522), .C2(n15538), .A(n15521), .B(n15520), .ZN(
        n15524) );
  OAI211_X1 U17082 ( .C1(n15525), .C2(n15529), .A(n15524), .B(n15523), .ZN(
        P3_U3187) );
  AOI21_X1 U17083 ( .B1(n7945), .B2(n15527), .A(n15526), .ZN(n15548) );
  OAI22_X1 U17084 ( .A1(n15531), .A2(n15530), .B1(n15529), .B2(n15528), .ZN(
        n15544) );
  AOI21_X1 U17085 ( .B1(n15534), .B2(n15533), .A(n15532), .ZN(n15542) );
  OAI21_X1 U17086 ( .B1(n15537), .B2(n15536), .A(n15535), .ZN(n15539) );
  NAND2_X1 U17087 ( .A1(n15539), .A2(n15538), .ZN(n15540) );
  OAI21_X1 U17088 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15543) );
  AOI211_X1 U17089 ( .C1(P3_REG3_REG_13__SCAN_IN), .C2(P3_U3151), .A(n15544), 
        .B(n15543), .ZN(n15546) );
  OAI21_X1 U17090 ( .B1(n15548), .B2(n15547), .A(n15546), .ZN(P3_U3195) );
  XNOR2_X1 U17091 ( .A(n15549), .B(n15555), .ZN(n15576) );
  NOR2_X1 U17092 ( .A1(n15550), .A2(n15606), .ZN(n15575) );
  INV_X1 U17093 ( .A(n15575), .ZN(n15551) );
  OAI22_X1 U17094 ( .A1(n15553), .A2(n10136), .B1(n15552), .B2(n15551), .ZN(
        n15564) );
  NAND3_X1 U17095 ( .A1(n15556), .A2(n15555), .A3(n15554), .ZN(n15557) );
  AND2_X1 U17096 ( .A1(n15558), .A2(n15557), .ZN(n15559) );
  OAI222_X1 U17097 ( .A1(n15563), .A2(n15562), .B1(n15561), .B2(n8123), .C1(
        n15560), .C2(n15559), .ZN(n15574) );
  AOI211_X1 U17098 ( .C1(n15576), .C2(n15565), .A(n15564), .B(n15574), .ZN(
        n15567) );
  AOI22_X1 U17099 ( .A1(n14943), .A2(n15568), .B1(n15567), .B2(n15566), .ZN(
        P3_U3231) );
  INV_X1 U17100 ( .A(n15569), .ZN(n15572) );
  INV_X1 U17101 ( .A(n15570), .ZN(n15571) );
  AOI211_X1 U17102 ( .C1(n15611), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        n15615) );
  AOI22_X1 U17103 ( .A1(n15613), .A2(n15615), .B1(n7754), .B2(n15612), .ZN(
        P3_U3393) );
  AOI211_X1 U17104 ( .C1(n15576), .C2(n15600), .A(n15575), .B(n15574), .ZN(
        n15617) );
  AOI22_X1 U17105 ( .A1(n15613), .A2(n15617), .B1(n7768), .B2(n15612), .ZN(
        P3_U3396) );
  INV_X1 U17106 ( .A(n15611), .ZN(n15595) );
  OAI22_X1 U17107 ( .A1(n15578), .A2(n15595), .B1(n15606), .B2(n15577), .ZN(
        n15580) );
  NOR2_X1 U17108 ( .A1(n15580), .A2(n15579), .ZN(n15619) );
  AOI22_X1 U17109 ( .A1(n15613), .A2(n15619), .B1(n7779), .B2(n15612), .ZN(
        P3_U3399) );
  OAI22_X1 U17110 ( .A1(n15582), .A2(n15595), .B1(n15606), .B2(n15581), .ZN(
        n15583) );
  NOR2_X1 U17111 ( .A1(n15584), .A2(n15583), .ZN(n15621) );
  AOI22_X1 U17112 ( .A1(n15613), .A2(n15621), .B1(n7791), .B2(n15612), .ZN(
        P3_U3402) );
  NOR2_X1 U17113 ( .A1(n15585), .A2(n15606), .ZN(n15587) );
  AOI211_X1 U17114 ( .C1(n15600), .C2(n15588), .A(n15587), .B(n15586), .ZN(
        n15623) );
  AOI22_X1 U17115 ( .A1(n15613), .A2(n15623), .B1(n7810), .B2(n15612), .ZN(
        P3_U3405) );
  OAI22_X1 U17116 ( .A1(n15590), .A2(n15595), .B1(n15589), .B2(n15606), .ZN(
        n15591) );
  NOR2_X1 U17117 ( .A1(n15592), .A2(n15591), .ZN(n15624) );
  AOI22_X1 U17118 ( .A1(n15613), .A2(n15624), .B1(n7828), .B2(n15612), .ZN(
        P3_U3408) );
  INV_X1 U17119 ( .A(n15593), .ZN(n15598) );
  OAI22_X1 U17120 ( .A1(n15596), .A2(n15595), .B1(n15606), .B2(n15594), .ZN(
        n15597) );
  NOR2_X1 U17121 ( .A1(n15598), .A2(n15597), .ZN(n15625) );
  AOI22_X1 U17122 ( .A1(n15613), .A2(n15625), .B1(n7843), .B2(n15612), .ZN(
        P3_U3411) );
  INV_X1 U17123 ( .A(n15599), .ZN(n15605) );
  INV_X1 U17124 ( .A(n15600), .ZN(n15602) );
  OAI22_X1 U17125 ( .A1(n15603), .A2(n15602), .B1(n15601), .B2(n15606), .ZN(
        n15604) );
  NOR2_X1 U17126 ( .A1(n15605), .A2(n15604), .ZN(n15627) );
  AOI22_X1 U17127 ( .A1(n15613), .A2(n15627), .B1(n7859), .B2(n15612), .ZN(
        P3_U3414) );
  NOR2_X1 U17128 ( .A1(n15607), .A2(n15606), .ZN(n15609) );
  AOI211_X1 U17129 ( .C1(n15611), .C2(n15610), .A(n15609), .B(n15608), .ZN(
        n15630) );
  AOI22_X1 U17130 ( .A1(n15613), .A2(n15630), .B1(n7878), .B2(n15612), .ZN(
        P3_U3417) );
  INV_X1 U17131 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U17132 ( .A1(n15631), .A2(n15615), .B1(n15614), .B2(n15628), .ZN(
        P3_U3460) );
  AOI22_X1 U17133 ( .A1(n15631), .A2(n15617), .B1(n15616), .B2(n15628), .ZN(
        P3_U3461) );
  AOI22_X1 U17134 ( .A1(n15631), .A2(n15619), .B1(n15618), .B2(n15628), .ZN(
        P3_U3462) );
  AOI22_X1 U17135 ( .A1(n15631), .A2(n15621), .B1(n15620), .B2(n15628), .ZN(
        P3_U3463) );
  AOI22_X1 U17136 ( .A1(n15631), .A2(n15623), .B1(n15622), .B2(n15628), .ZN(
        P3_U3464) );
  AOI22_X1 U17137 ( .A1(n15631), .A2(n15624), .B1(n10206), .B2(n15628), .ZN(
        P3_U3465) );
  AOI22_X1 U17138 ( .A1(n15631), .A2(n15625), .B1(n10196), .B2(n15628), .ZN(
        P3_U3466) );
  AOI22_X1 U17139 ( .A1(n15631), .A2(n15627), .B1(n15626), .B2(n15628), .ZN(
        P3_U3467) );
  AOI22_X1 U17140 ( .A1(n15631), .A2(n15630), .B1(n15629), .B2(n15628), .ZN(
        P3_U3468) );
  XOR2_X1 U17141 ( .A(n15633), .B(n15632), .Z(SUB_1596_U59) );
  XNOR2_X1 U17142 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15634), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17143 ( .B1(n15635), .B2(n10024), .A(n15644), .ZN(SUB_1596_U53) );
  XNOR2_X1 U17144 ( .A(n15637), .B(n15636), .ZN(SUB_1596_U56) );
  OAI21_X1 U17145 ( .B1(n15640), .B2(n15639), .A(n15638), .ZN(n15642) );
  XOR2_X1 U17146 ( .A(n15642), .B(n15641), .Z(SUB_1596_U60) );
  XOR2_X1 U17147 ( .A(n15644), .B(n15643), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7321 ( .A(n8429), .Z(n6593) );
  BUF_X1 U7387 ( .A(n10250), .Z(n6573) );
  CLKBUF_X2 U7426 ( .A(n12303), .Z(n12413) );
  CLKBUF_X1 U7427 ( .A(n7654), .Z(n12149) );
  CLKBUF_X1 U7540 ( .A(n13273), .Z(n6755) );
  AND4_X1 U7646 ( .A1(n9416), .A2(n9415), .A3(n9501), .A4(n9692), .ZN(n15648)
         );
endmodule

