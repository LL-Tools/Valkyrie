

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646;

  MUX2_X1 U4907 ( .A(n6630), .B(n6629), .S(n10189), .Z(n6631) );
  MUX2_X1 U4908 ( .A(n10506), .B(n6629), .S(n10194), .Z(n6626) );
  NAND2_X1 U4909 ( .A1(n8391), .A2(n9992), .ZN(n9762) );
  OAI21_X1 U4910 ( .B1(n8032), .B2(n6482), .A(n5083), .ZN(n8158) );
  NAND2_X2 U4911 ( .A1(n6204), .A2(n6203), .ZN(n8188) );
  INV_X1 U4912 ( .A(n8870), .ZN(n8056) );
  BUF_X2 U4913 ( .A(n5321), .Z(n5905) );
  CLKBUF_X2 U4914 ( .A(n5321), .Z(n8736) );
  NAND4_X1 U4915 ( .A1(n6076), .A2(n5111), .A3(n6075), .A4(n6074), .ZN(n10200)
         );
  NAND2_X1 U4916 ( .A1(n5304), .A2(n10112), .ZN(n7217) );
  CLKBUF_X2 U4917 ( .A(n6125), .Z(n6681) );
  BUF_X1 U4918 ( .A(n6072), .Z(n6444) );
  XNOR2_X2 U4919 ( .A(n6086), .B(n6101), .ZN(n7297) );
  CLKBUF_X1 U4920 ( .A(n9484), .Z(n4405) );
  OAI21_X1 U4921 ( .B1(n5950), .B2(n5949), .A(n9913), .ZN(n9484) );
  AND2_X1 U4922 ( .A1(n8897), .A2(n8896), .ZN(n8898) );
  NOR2_X1 U4923 ( .A1(n5328), .A2(n5223), .ZN(n5225) );
  AND2_X1 U4924 ( .A1(n8898), .A2(n8928), .ZN(n8899) );
  CLKBUF_X3 U4925 ( .A(n6087), .Z(n6678) );
  INV_X2 U4926 ( .A(n8738), .ZN(n5876) );
  INV_X1 U4927 ( .A(n7946), .ZN(n6482) );
  NAND2_X1 U4928 ( .A1(n4992), .A2(n4991), .ZN(n7969) );
  AND2_X1 U4929 ( .A1(n5143), .A2(n5180), .ZN(n4526) );
  BUF_X1 U4930 ( .A(n5160), .Z(n5161) );
  INV_X2 U4931 ( .A(n6063), .ZN(n8711) );
  NAND2_X1 U4932 ( .A1(n7091), .A2(n7859), .ZN(n7094) );
  AOI21_X1 U4933 ( .B1(n7085), .B2(n4811), .A(n4520), .ZN(n4810) );
  NAND2_X1 U4934 ( .A1(n6041), .A2(n7168), .ZN(n6657) );
  AND2_X2 U4935 ( .A1(n6952), .A2(n4797), .ZN(n9053) );
  AND3_X1 U4936 ( .A1(n6107), .A2(n6106), .A3(n6105), .ZN(n10231) );
  NOR2_X1 U4937 ( .A1(n8562), .A2(n8647), .ZN(n8652) );
  INV_X1 U4938 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5217) );
  AND4_X1 U4939 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n7579)
         );
  AOI21_X1 U4940 ( .B1(n7544), .B2(n6637), .A(n6636), .ZN(n7744) );
  AOI222_X1 U4941 ( .A1(n10202), .A2(n9070), .B1(n9069), .B2(n10199), .C1(
        n9095), .C2(n9236), .ZN(n9368) );
  OR2_X1 U4942 ( .A1(n4929), .A2(n4719), .ZN(n4717) );
  OAI211_X1 U4943 ( .C1(n7217), .C2(n7250), .A(n4438), .B(n5284), .ZN(n10156)
         );
  AND4_X1 U4944 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n8423)
         );
  INV_X1 U4945 ( .A(n8243), .ZN(n8142) );
  INV_X1 U4946 ( .A(n6034), .ZN(n9443) );
  NAND2_X1 U4947 ( .A1(n6006), .A2(n6427), .ZN(n7912) );
  NAND2_X1 U4949 ( .A1(n5846), .A2(n5845), .ZN(n9611) );
  INV_X1 U4950 ( .A(n5150), .ZN(n10109) );
  AND2_X1 U4951 ( .A1(n4774), .A2(n4472), .ZN(n4406) );
  INV_X2 U4952 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5293) );
  INV_X2 U4953 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5255) );
  NOR2_X2 U4954 ( .A1(n5606), .A2(n5605), .ZN(n4569) );
  AOI21_X2 U4955 ( .B1(n8975), .B2(n8974), .A(n8973), .ZN(n9004) );
  NAND2_X2 U4956 ( .A1(n4930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6012) );
  OR2_X2 U4957 ( .A1(n6157), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6100) );
  NAND2_X2 U4958 ( .A1(n8764), .A2(n4807), .ZN(n7007) );
  NOR4_X2 U4959 ( .A1(n8541), .A2(n8540), .A3(n7797), .A4(n8539), .ZN(n8543)
         );
  NAND2_X2 U4960 ( .A1(n4688), .A2(n5958), .ZN(n5974) );
  AND2_X2 U4961 ( .A1(n5957), .A2(n6154), .ZN(n4688) );
  NOR2_X2 U4962 ( .A1(n9212), .A2(n6915), .ZN(n4803) );
  INV_X4 U4963 ( .A(n4410), .ZN(n7072) );
  NAND3_X2 U4964 ( .A1(n5311), .A2(n4467), .A3(n5312), .ZN(n6537) );
  INV_X1 U4965 ( .A(n8871), .ZN(n8096) );
  NOR4_X2 U4966 ( .A1(n6818), .A2(n9210), .A3(n9201), .A4(n6706), .ZN(n6707)
         );
  NAND2_X1 U4967 ( .A1(n4965), .A2(n4963), .ZN(n4407) );
  NOR2_X2 U4968 ( .A1(n8944), .A2(n5110), .ZN(n8945) );
  AOI21_X2 U4969 ( .B1(n8923), .B2(n8921), .A(n8922), .ZN(n8944) );
  NAND2_X2 U4970 ( .A1(n6728), .A2(n6727), .ZN(n7574) );
  AND2_X2 U4971 ( .A1(n9132), .A2(n4477), .ZN(n4419) );
  XNOR2_X2 U4972 ( .A(n5572), .B(n5571), .ZN(n7360) );
  NAND2_X2 U4973 ( .A1(n5710), .A2(n5709), .ZN(n10014) );
  AOI21_X2 U4974 ( .B1(n8984), .B2(n8983), .A(n8982), .ZN(n8985) );
  AOI21_X1 U4975 ( .B1(n6536), .B2(n9964), .A(n6535), .ZN(n8698) );
  NAND2_X1 U4976 ( .A1(n9774), .A2(n8630), .ZN(n6970) );
  NAND2_X1 U4977 ( .A1(n9520), .A2(n5828), .ZN(n9487) );
  INV_X1 U4978 ( .A(n9760), .ZN(n6608) );
  NAND2_X1 U4979 ( .A1(n6509), .A2(n6508), .ZN(n9767) );
  CLKBUF_X1 U4980 ( .A(n9470), .Z(n4535) );
  NAND2_X1 U4981 ( .A1(n5893), .A2(n5892), .ZN(n9782) );
  NAND2_X1 U4982 ( .A1(n6380), .A2(n6379), .ZN(n9364) );
  NAND2_X1 U4983 ( .A1(n8069), .A2(n4671), .ZN(n8325) );
  AOI21_X1 U4984 ( .B1(n9783), .B2(n5899), .A(n5898), .ZN(n9594) );
  OR2_X1 U4985 ( .A1(n6797), .A2(n6696), .ZN(n9223) );
  AND2_X1 U4986 ( .A1(n8079), .A2(n6198), .ZN(n8208) );
  NAND2_X1 U4987 ( .A1(n5690), .A2(n5689), .ZN(n10018) );
  NAND2_X1 U4988 ( .A1(n5497), .A2(n5496), .ZN(n5520) );
  INV_X1 U4989 ( .A(n8367), .ZN(n4408) );
  NAND2_X1 U4990 ( .A1(n8419), .A2(n9629), .ZN(n8433) );
  NAND2_X1 U4991 ( .A1(n8593), .A2(n8600), .ZN(n8536) );
  INV_X1 U4992 ( .A(n7811), .ZN(n4409) );
  INV_X2 U4993 ( .A(n10156), .ZN(n7768) );
  INV_X2 U4994 ( .A(n5228), .ZN(n8425) );
  NAND4_X1 U4995 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n8874)
         );
  NAND2_X1 U4996 ( .A1(n5227), .A2(n5849), .ZN(n4731) );
  INV_X2 U4997 ( .A(n5849), .ZN(n8734) );
  INV_X1 U4998 ( .A(n8518), .ZN(n8521) );
  INV_X2 U5000 ( .A(n6678), .ZN(n6300) );
  BUF_X1 U5001 ( .A(n7116), .Z(n4562) );
  INV_X2 U5002 ( .A(n7912), .ZN(n4797) );
  INV_X4 U5003 ( .A(n6518), .ZN(n6615) );
  INV_X1 U5004 ( .A(n7780), .ZN(n7448) );
  NAND2_X2 U5005 ( .A1(n4410), .A2(n6449), .ZN(n6041) );
  INV_X2 U5006 ( .A(n5362), .ZN(n7168) );
  OR2_X1 U5007 ( .A1(n8565), .A2(n8564), .ZN(n8682) );
  NOR3_X1 U5008 ( .A1(n6854), .A2(n6714), .A3(n6713), .ZN(n6715) );
  NAND2_X1 U5009 ( .A1(n4929), .A2(n4435), .ZN(n9592) );
  OR2_X1 U5010 ( .A1(n6970), .A2(n8561), .ZN(n6972) );
  NAND2_X1 U5011 ( .A1(n6437), .A2(n6436), .ZN(n8729) );
  AND2_X1 U5012 ( .A1(n8686), .A2(n6969), .ZN(n9763) );
  OR2_X1 U5013 ( .A1(n9012), .A2(n8989), .ZN(n8990) );
  OR2_X1 U5014 ( .A1(n8519), .A2(n8664), .ZN(n8667) );
  AOI21_X1 U5015 ( .B1(n9043), .B2(n10202), .A(n9042), .ZN(n9350) );
  NAND2_X1 U5016 ( .A1(n6968), .A2(n4670), .ZN(n8686) );
  AOI21_X1 U5017 ( .B1(n4695), .B2(n4697), .A(n4464), .ZN(n4693) );
  NAND2_X1 U5018 ( .A1(n6618), .A2(n6617), .ZN(n8519) );
  OAI21_X1 U5019 ( .B1(n5068), .B2(n4588), .A(n4587), .ZN(n6968) );
  NAND2_X1 U5020 ( .A1(n6607), .A2(n6606), .ZN(n9760) );
  OR2_X1 U5021 ( .A1(n8692), .A2(n6528), .ZN(n8574) );
  NAND2_X1 U5022 ( .A1(n6520), .A2(n6519), .ZN(n8692) );
  NAND2_X1 U5023 ( .A1(n5772), .A2(n5771), .ZN(n9554) );
  NAND2_X1 U5024 ( .A1(n5060), .A2(n6574), .ZN(n4587) );
  AOI21_X1 U5025 ( .B1(n9767), .B2(n9781), .A(n9949), .ZN(n6977) );
  OR2_X1 U5026 ( .A1(n5063), .A2(n4589), .ZN(n4588) );
  OAI21_X1 U5027 ( .B1(n10110), .B2(n6657), .A(n6658), .ZN(n6964) );
  AOI21_X1 U5028 ( .B1(n8939), .B2(n4430), .A(n8938), .ZN(n8957) );
  OAI22_X2 U5029 ( .A1(n9094), .A2(n6918), .B1(n9109), .B2(n9380), .ZN(n9081)
         );
  NAND2_X1 U5030 ( .A1(n6394), .A2(n6393), .ZN(n9358) );
  XNOR2_X1 U5031 ( .A(n6511), .B(n6510), .ZN(n6654) );
  NAND2_X1 U5032 ( .A1(n6503), .A2(n6502), .ZN(n6511) );
  NAND2_X1 U5033 ( .A1(n5865), .A2(n5864), .ZN(n9981) );
  XNOR2_X1 U5034 ( .A(n6501), .B(n6500), .ZN(n8703) );
  AOI21_X1 U5035 ( .B1(n4923), .B2(n9468), .A(n4922), .ZN(n4921) );
  NAND3_X1 U5036 ( .A1(n7092), .A2(n7094), .A3(P2_REG2_REG_11__SCAN_IN), .ZN(
        n7857) );
  NAND2_X1 U5037 ( .A1(n5887), .A2(n5886), .ZN(n6501) );
  NAND2_X1 U5038 ( .A1(n6371), .A2(n6370), .ZN(n9370) );
  AND2_X1 U5039 ( .A1(n5941), .A2(n5940), .ZN(n8739) );
  NAND2_X1 U5040 ( .A1(n8325), .A2(n5563), .ZN(n5591) );
  NAND2_X2 U5041 ( .A1(n5808), .A2(n5807), .ZN(n9991) );
  NAND2_X1 U5042 ( .A1(n6346), .A2(n6345), .ZN(n9375) );
  AND2_X1 U5043 ( .A1(n7084), .A2(n7085), .ZN(n7864) );
  NAND2_X1 U5044 ( .A1(n5730), .A2(n5729), .ZN(n9876) );
  NAND2_X1 U5045 ( .A1(n6324), .A2(n6323), .ZN(n9392) );
  NAND2_X1 U5046 ( .A1(n6335), .A2(n6334), .ZN(n9386) );
  NAND2_X1 U5047 ( .A1(n5025), .A2(n5023), .ZN(n9235) );
  AND2_X1 U5048 ( .A1(n5024), .A2(n4427), .ZN(n5023) );
  INV_X1 U5049 ( .A(n5013), .ZN(n5012) );
  AND2_X1 U5050 ( .A1(n6908), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U5051 ( .A1(n5661), .A2(n5660), .ZN(n10023) );
  AND2_X1 U5052 ( .A1(n10039), .A2(n8411), .ZN(n9929) );
  NAND2_X2 U5053 ( .A1(n5547), .A2(n5546), .ZN(n10042) );
  NAND2_X1 U5054 ( .A1(n6244), .A2(n6243), .ZN(n9417) );
  NAND2_X1 U5055 ( .A1(n5683), .A2(n5682), .ZN(n5707) );
  NAND2_X1 U5056 ( .A1(n7464), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U5057 ( .A1(n4976), .A2(n4476), .ZN(n5683) );
  NAND2_X1 U5058 ( .A1(n6222), .A2(n6221), .ZN(n9428) );
  AOI21_X1 U5059 ( .B1(n7482), .B2(n4961), .A(n4958), .ZN(n7759) );
  NAND2_X1 U5060 ( .A1(n5500), .A2(n5499), .ZN(n10053) );
  AND2_X1 U5061 ( .A1(n7155), .A2(n4538), .ZN(n7464) );
  NAND2_X1 U5062 ( .A1(n5449), .A2(n5448), .ZN(n10062) );
  NAND2_X1 U5063 ( .A1(n7017), .A2(n7460), .ZN(n7159) );
  OAI21_X1 U5064 ( .B1(n5520), .B2(n4776), .A(n4406), .ZN(n4770) );
  XNOR2_X1 U5065 ( .A(n4684), .B(n8734), .ZN(n8232) );
  XNOR2_X1 U5066 ( .A(n5520), .B(n5515), .ZN(n7338) );
  NAND2_X1 U5067 ( .A1(n6196), .A2(n6195), .ZN(n8091) );
  NAND2_X1 U5068 ( .A1(n5468), .A2(n5467), .ZN(n8205) );
  NAND2_X1 U5069 ( .A1(n7370), .A2(n7016), .ZN(n7017) );
  OR2_X1 U5070 ( .A1(n8871), .A2(n8109), .ZN(n6902) );
  XNOR2_X1 U5071 ( .A(n5495), .B(n5494), .ZN(n7230) );
  AOI21_X1 U5072 ( .B1(n8731), .B2(n8142), .A(n4685), .ZN(n4684) );
  NAND2_X1 U5073 ( .A1(n4612), .A2(n5381), .ZN(n8367) );
  XNOR2_X1 U5074 ( .A(n5463), .B(n5464), .ZN(n7224) );
  AND2_X1 U5075 ( .A1(n5402), .A2(n5401), .ZN(n8243) );
  NAND2_X1 U5076 ( .A1(n5431), .A2(n5116), .ZN(n4754) );
  INV_X1 U5077 ( .A(n10145), .ZN(n8419) );
  NAND2_X1 U5078 ( .A1(n5251), .A2(n5250), .ZN(n10145) );
  AND2_X1 U5079 ( .A1(n6121), .A2(n6120), .ZN(n10240) );
  AND2_X1 U5080 ( .A1(n5421), .A2(n5420), .ZN(n6478) );
  NAND2_X1 U5081 ( .A1(n7616), .A2(n6747), .ZN(n6890) );
  NAND2_X1 U5082 ( .A1(n8414), .A2(n8592), .ZN(n7811) );
  NAND2_X1 U5083 ( .A1(n4465), .A2(n6051), .ZN(n8878) );
  NAND2_X1 U5084 ( .A1(n6632), .A2(n4461), .ZN(n6728) );
  OR2_X1 U5085 ( .A1(n6089), .A2(n6088), .ZN(n7624) );
  INV_X1 U5086 ( .A(n10200), .ZN(n7387) );
  OR2_X1 U5087 ( .A1(n6160), .A2(n6192), .ZN(n7202) );
  INV_X1 U5088 ( .A(n10221), .ZN(n7548) );
  AND3_X1 U5089 ( .A1(n4788), .A2(n6079), .A3(n6078), .ZN(n10221) );
  AND4_X1 U5090 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n8417)
         );
  AND2_X1 U5091 ( .A1(n5109), .A2(n5496), .ZN(n4765) );
  NAND2_X1 U5092 ( .A1(n5123), .A2(n4605), .ZN(n7640) );
  NAND4_X1 U5093 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n6538)
         );
  NAND2_X1 U5094 ( .A1(n6091), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6046) );
  INV_X1 U5095 ( .A(n6072), .ZN(n6125) );
  AND2_X1 U5096 ( .A1(n6529), .A2(n7823), .ZN(n5223) );
  AND2_X1 U5097 ( .A1(n4903), .A2(n7305), .ZN(n4902) );
  INV_X2 U5098 ( .A(n6657), .ZN(n6675) );
  NAND2_X1 U5099 ( .A1(n5568), .A2(n5515), .ZN(n4776) );
  OR2_X1 U5100 ( .A1(n5626), .A2(n5625), .ZN(n5109) );
  INV_X1 U5101 ( .A(n7116), .ZN(n5328) );
  INV_X2 U5102 ( .A(n6041), .ZN(n6301) );
  NAND2_X1 U5103 ( .A1(n6041), .A2(n7193), .ZN(n6087) );
  MUX2_X1 U5104 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10116), .S(n4414), .Z(n7780)
         );
  OR2_X1 U5105 ( .A1(n7286), .A2(n4443), .ZN(n4903) );
  NAND3_X1 U5106 ( .A1(n5221), .A2(n5220), .A3(n5219), .ZN(n8526) );
  AND2_X1 U5107 ( .A1(n5167), .A2(n5222), .ZN(n6529) );
  AND2_X2 U5108 ( .A1(n5150), .A2(n5154), .ZN(n5899) );
  NAND2_X1 U5109 ( .A1(n5171), .A2(n5170), .ZN(n7823) );
  MUX2_X1 U5110 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6003), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6006) );
  XNOR2_X1 U5111 ( .A(n5174), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U5112 ( .A(n6104), .B(n6103), .ZN(n7305) );
  XNOR2_X1 U5113 ( .A(n6016), .B(n6015), .ZN(n8271) );
  OR2_X1 U5114 ( .A1(n6118), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U5115 ( .A(n5992), .B(n6000), .ZN(n7827) );
  NAND2_X1 U5116 ( .A1(n4525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5003) );
  INV_X2 U5117 ( .A(n6448), .ZN(n4410) );
  NAND2_X1 U5118 ( .A1(n6014), .A2(n6013), .ZN(n8223) );
  NAND2_X1 U5119 ( .A1(n4887), .A2(n6060), .ZN(n6157) );
  INV_X1 U5120 ( .A(n7007), .ZN(n4887) );
  AND2_X1 U5121 ( .A1(n4747), .A2(n6060), .ZN(n5957) );
  AND2_X1 U5122 ( .A1(n6152), .A2(n5954), .ZN(n5958) );
  AND3_X1 U5123 ( .A1(n5993), .A2(n5975), .A3(n5977), .ZN(n5962) );
  AND2_X1 U5124 ( .A1(n5172), .A2(n5145), .ZN(n5180) );
  NOR2_X1 U5125 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5956) );
  INV_X1 U5126 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4964) );
  NOR2_X1 U5127 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5955) );
  INV_X1 U5128 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4746) );
  NOR2_X2 U5129 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4715) );
  INV_X1 U5130 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U5131 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5959) );
  NOR2_X1 U5132 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4747) );
  NOR2_X1 U5133 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5960) );
  NOR2_X1 U5134 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5961) );
  INV_X1 U5135 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5993) );
  INV_X1 U5136 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6000) );
  INV_X1 U5137 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n10625) );
  INV_X1 U5138 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4807) );
  INV_X4 U5139 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5140 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5213) );
  INV_X1 U5141 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6060) );
  INV_X1 U5142 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5182) );
  INV_X1 U5143 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U5144 ( .A1(n6034), .A2(n9446), .ZN(n6072) );
  AND2_X1 U5145 ( .A1(n6025), .A2(n6034), .ZN(n6073) );
  OAI22_X2 U5146 ( .A1(n9235), .A2(n6909), .B1(n9428), .B2(n9225), .ZN(n9224)
         );
  AOI21_X2 U5147 ( .B1(n8967), .B2(n8969), .A(n8968), .ZN(n8999) );
  INV_X2 U5148 ( .A(n8526), .ZN(n5687) );
  NAND2_X1 U5149 ( .A1(n4965), .A2(n4963), .ZN(n4411) );
  NOR2_X2 U5150 ( .A1(n7573), .A2(n6725), .ZN(n7351) );
  NAND2_X1 U5151 ( .A1(n4415), .A2(n7193), .ZN(n4413) );
  NAND2_X1 U5152 ( .A1(n4414), .A2(n7193), .ZN(n6518) );
  INV_X1 U5153 ( .A(n10180), .ZN(n7818) );
  NAND2_X1 U5154 ( .A1(n7651), .A2(n10180), .ZN(n8592) );
  NAND4_X4 U5155 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n10198)
         );
  NAND2_X1 U5156 ( .A1(n6923), .A2(n4447), .ZN(n9038) );
  OAI21_X2 U5157 ( .B1(n7014), .B2(n4443), .A(n4902), .ZN(n7366) );
  NOR2_X2 U5158 ( .A1(n5732), .A2(n5731), .ZN(n4570) );
  OR2_X2 U5159 ( .A1(n5711), .A2(n9548), .ZN(n5732) );
  NAND2_X2 U5160 ( .A1(n9443), .A2(n6025), .ZN(n6090) );
  AOI21_X2 U5161 ( .B1(n4419), .B2(n9104), .A(n4545), .ZN(n9094) );
  NOR4_X1 U5162 ( .A1(n9255), .A2(n8178), .A3(n8094), .A4(n6704), .ZN(n6705)
         );
  NAND2_X1 U5163 ( .A1(n5304), .A2(n10112), .ZN(n4414) );
  NAND2_X2 U5164 ( .A1(n5304), .A2(n10112), .ZN(n4415) );
  NOR4_X1 U5165 ( .A1(n9104), .A2(n9121), .A3(n9139), .A4(n6709), .ZN(n6710)
         );
  AND2_X2 U5166 ( .A1(n9948), .A2(n10097), .ZN(n9922) );
  AND2_X2 U5167 ( .A1(n7816), .A2(n7768), .ZN(n7653) );
  INV_X2 U5168 ( .A(n7803), .ZN(n4992) );
  AND2_X1 U5169 ( .A1(n9811), .A2(n4996), .ZN(n6976) );
  NOR2_X2 U5170 ( .A1(n7948), .A2(n4997), .ZN(n8124) );
  NOR2_X2 U5171 ( .A1(n7969), .A2(n8142), .ZN(n7968) );
  NAND2_X1 U5172 ( .A1(n4415), .A2(n7168), .ZN(n4417) );
  AND2_X1 U5173 ( .A1(n6255), .A2(n5989), .ZN(n6258) );
  INV_X1 U5174 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5989) );
  NOR2_X1 U5175 ( .A1(n5745), .A2(n4987), .ZN(n4986) );
  INV_X1 U5176 ( .A(n4989), .ZN(n4987) );
  OR2_X1 U5177 ( .A1(n7528), .A2(n7526), .ZN(n6951) );
  NAND2_X1 U5178 ( .A1(n4437), .A2(n5962), .ZN(n5963) );
  OR2_X1 U5179 ( .A1(n5073), .A2(n4599), .ZN(n4598) );
  INV_X1 U5180 ( .A(n4600), .ZN(n4599) );
  AND2_X1 U5181 ( .A1(n6514), .A2(n6507), .ZN(n6510) );
  NAND4_X2 U5182 ( .A1(n5186), .A2(n5184), .A3(n4715), .A4(n5142), .ZN(n5246)
         );
  INV_X2 U5184 ( .A(n6670), .ZN(n6122) );
  AOI21_X1 U5185 ( .B1(n9150), .B2(n9149), .A(n6916), .ZN(n9132) );
  OR2_X1 U5186 ( .A1(n9358), .A2(n9062), .ZN(n6922) );
  INV_X1 U5187 ( .A(n6840), .ZN(n4699) );
  NOR2_X1 U5188 ( .A1(n6733), .A2(n4789), .ZN(n6740) );
  AOI21_X1 U5189 ( .B1(n8435), .B2(n8592), .A(n8434), .ZN(n8439) );
  OAI21_X1 U5190 ( .B1(n4841), .B2(n4840), .A(n8444), .ZN(n4839) );
  INV_X1 U5191 ( .A(n8440), .ZN(n4834) );
  INV_X1 U5192 ( .A(n6835), .ZN(n4762) );
  NAND2_X1 U5193 ( .A1(n6903), .A2(n6902), .ZN(n5032) );
  NAND2_X1 U5194 ( .A1(n8513), .A2(n8687), .ZN(n4625) );
  AND2_X1 U5195 ( .A1(n5108), .A2(n4546), .ZN(n6712) );
  NOR2_X1 U5196 ( .A1(n6929), .A2(n4547), .ZN(n4546) );
  NOR2_X1 U5197 ( .A1(n6711), .A2(n4577), .ZN(n5108) );
  INV_X1 U5198 ( .A(n6861), .ZN(n4547) );
  AND2_X1 U5199 ( .A1(n6862), .A2(n6855), .ZN(n6860) );
  NAND2_X1 U5200 ( .A1(n5978), .A2(n5977), .ZN(n5988) );
  INV_X1 U5201 ( .A(n6201), .ZN(n5978) );
  AND2_X1 U5202 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  OR2_X1 U5203 ( .A1(n6964), .A2(n8719), .ZN(n6866) );
  INV_X1 U5204 ( .A(n6358), .ZN(n6347) );
  INV_X1 U5205 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6028) );
  OR2_X1 U5206 ( .A1(n8794), .A2(n9214), .ZN(n6808) );
  NAND2_X1 U5207 ( .A1(n6012), .A2(n5966), .ZN(n6008) );
  OAI211_X1 U5208 ( .C1(n8571), .C2(n5224), .A(n7730), .B(n4562), .ZN(n5227)
         );
  AND2_X1 U5209 ( .A1(n8196), .A2(n8192), .ZN(n4549) );
  XNOR2_X1 U5210 ( .A(n5391), .B(n8734), .ZN(n5482) );
  AOI21_X1 U5211 ( .B1(n4924), .B2(n4921), .A(n4682), .ZN(n4681) );
  INV_X1 U5212 ( .A(n5769), .ZN(n4682) );
  INV_X1 U5213 ( .A(n4921), .ZN(n4683) );
  INV_X1 U5214 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5215 ( .B1(n5619), .B2(n4727), .A(n9514), .ZN(n4726) );
  INV_X1 U5216 ( .A(n9512), .ZN(n4727) );
  INV_X1 U5217 ( .A(n5900), .ZN(n5321) );
  OR2_X1 U5218 ( .A1(n8517), .A2(n4844), .ZN(n4629) );
  NOR2_X1 U5220 ( .A1(n9795), .A2(n5007), .ZN(n5006) );
  INV_X1 U5221 ( .A(n4567), .ZN(n5894) );
  NOR2_X1 U5222 ( .A1(n8553), .A2(n5095), .ZN(n5094) );
  INV_X1 U5223 ( .A(n5097), .ZN(n5095) );
  OAI21_X1 U5224 ( .B1(n4657), .B2(n4655), .A(n9906), .ZN(n4652) );
  NOR2_X1 U5225 ( .A1(n6564), .A2(n4601), .ZN(n4600) );
  INV_X1 U5226 ( .A(n6563), .ZN(n4601) );
  NAND2_X1 U5227 ( .A1(n5071), .A2(n4456), .ZN(n4604) );
  NAND2_X1 U5228 ( .A1(n8547), .A2(n8454), .ZN(n5013) );
  INV_X1 U5229 ( .A(n6552), .ZN(n5084) );
  NAND2_X1 U5230 ( .A1(n4408), .A2(n4609), .ZN(n8444) );
  NAND2_X1 U5231 ( .A1(n6475), .A2(n10156), .ZN(n8600) );
  NAND2_X1 U5232 ( .A1(n7640), .A2(n6469), .ZN(n8412) );
  NAND2_X1 U5233 ( .A1(n6501), .A2(n6500), .ZN(n6503) );
  INV_X1 U5234 ( .A(SI_22_), .ZN(n5747) );
  INV_X1 U5235 ( .A(n4986), .ZN(n4985) );
  AOI21_X1 U5236 ( .B1(n4984), .B2(n4986), .A(n4470), .ZN(n4983) );
  INV_X1 U5237 ( .A(n4990), .ZN(n4984) );
  INV_X1 U5238 ( .A(n5246), .ZN(n4919) );
  OR2_X1 U5239 ( .A1(n6294), .A2(n9187), .ZN(n6295) );
  NAND2_X1 U5240 ( .A1(n8826), .A2(n4952), .ZN(n4951) );
  INV_X1 U5241 ( .A(n6312), .ZN(n4952) );
  AND2_X1 U5242 ( .A1(n7515), .A2(n6084), .ZN(n4962) );
  NOR2_X1 U5243 ( .A1(n8277), .A2(n4955), .ZN(n4954) );
  INV_X1 U5244 ( .A(n6238), .ZN(n4955) );
  BUF_X1 U5245 ( .A(n6090), .Z(n6670) );
  INV_X1 U5246 ( .A(n6915), .ZN(n4804) );
  INV_X1 U5247 ( .A(n9159), .ZN(n4802) );
  NAND2_X1 U5248 ( .A1(n9160), .A2(n6914), .ZN(n4805) );
  AND2_X1 U5249 ( .A1(n5999), .A2(n5998), .ZN(n7540) );
  AND2_X1 U5250 ( .A1(n7827), .A2(n5103), .ZN(n5998) );
  NAND2_X1 U5251 ( .A1(n7533), .A2(n7532), .ZN(n7542) );
  AND2_X1 U5252 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  AOI21_X1 U5253 ( .B1(n6654), .B2(n6675), .A(n4509), .ZN(n8714) );
  AND2_X1 U5254 ( .A1(n4492), .A2(n4696), .ZN(n4695) );
  NOR2_X1 U5255 ( .A1(n9074), .A2(n4785), .ZN(n4782) );
  AOI21_X1 U5256 ( .B1(n4468), .B2(n6823), .A(n4703), .ZN(n4702) );
  INV_X1 U5257 ( .A(n6823), .ZN(n4704) );
  INV_X1 U5258 ( .A(n9261), .ZN(n10199) );
  XNOR2_X1 U5259 ( .A(n6425), .B(n6424), .ZN(n7068) );
  NAND2_X1 U5260 ( .A1(n6407), .A2(n6406), .ZN(n7187) );
  NAND2_X1 U5261 ( .A1(n4806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U5262 ( .A(n6194), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7088) );
  NAND3_X1 U5263 ( .A1(n4728), .A2(n5910), .A3(n5906), .ZN(n7116) );
  INV_X1 U5264 ( .A(n9610), .ZN(n6499) );
  NAND2_X1 U5265 ( .A1(n8526), .A2(n7823), .ZN(n8571) );
  INV_X1 U5266 ( .A(n5936), .ZN(n6524) );
  INV_X2 U5267 ( .A(n6524), .ZN(n6620) );
  OR2_X1 U5268 ( .A1(n7431), .A2(n4504), .ZN(n4871) );
  OR2_X1 U5269 ( .A1(n9765), .A2(n6521), .ZN(n5941) );
  INV_X1 U5270 ( .A(n9595), .ZN(n8398) );
  AOI21_X1 U5271 ( .B1(n5094), .B2(n5092), .A(n4446), .ZN(n5091) );
  INV_X1 U5272 ( .A(n5098), .ZN(n5092) );
  NAND2_X1 U5273 ( .A1(n4602), .A2(n4600), .ZN(n6566) );
  INV_X1 U5274 ( .A(n7217), .ZN(n5688) );
  OR2_X1 U5275 ( .A1(n10110), .A2(n6518), .ZN(n6520) );
  XNOR2_X1 U5276 ( .A(n5148), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U5277 ( .A1(n10104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U5278 ( .A(n5149), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U5279 ( .A1(n4860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5149) );
  OAI21_X1 U5280 ( .B1(n5601), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5633) );
  INV_X1 U5281 ( .A(n8875), .ZN(n7517) );
  AOI21_X1 U5282 ( .B1(n6688), .B2(n5046), .A(n5045), .ZN(n6717) );
  NAND2_X1 U5283 ( .A1(n6403), .A2(n6402), .ZN(n9062) );
  NAND2_X1 U5284 ( .A1(n9065), .A2(n6659), .ZN(n4733) );
  NAND2_X1 U5285 ( .A1(n6353), .A2(n6352), .ZN(n9095) );
  NAND2_X1 U5286 ( .A1(n9350), .A2(n10257), .ZN(n9275) );
  INV_X1 U5287 ( .A(n6728), .ZN(n4794) );
  NAND2_X1 U5288 ( .A1(n4441), .A2(n4792), .ZN(n4791) );
  INV_X1 U5289 ( .A(n6727), .ZN(n4792) );
  NAND2_X1 U5290 ( .A1(n6726), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U5291 ( .A1(n4859), .A2(n4857), .ZN(n8432) );
  AOI21_X1 U5292 ( .B1(n8415), .B2(n8518), .A(n8536), .ZN(n4859) );
  NAND2_X1 U5293 ( .A1(n4519), .A2(n4858), .ZN(n4857) );
  AND2_X1 U5294 ( .A1(n8416), .A2(n8599), .ZN(n4856) );
  NOR2_X1 U5295 ( .A1(n6760), .A2(n6759), .ZN(n6770) );
  NOR2_X1 U5296 ( .A1(n6744), .A2(n9053), .ZN(n4801) );
  AND2_X1 U5297 ( .A1(n6770), .A2(n7742), .ZN(n4799) );
  AND2_X1 U5298 ( .A1(n8453), .A2(n8605), .ZN(n4843) );
  NAND2_X1 U5299 ( .A1(n4839), .A2(n8450), .ZN(n4635) );
  OAI21_X1 U5300 ( .B1(n4466), .B2(n8440), .A(n4841), .ZN(n8448) );
  NAND2_X1 U5301 ( .A1(n4848), .A2(n4847), .ZN(n8471) );
  INV_X1 U5302 ( .A(n9919), .ZN(n4847) );
  AND2_X1 U5303 ( .A1(n4757), .A2(n4489), .ZN(n4755) );
  NOR2_X1 U5304 ( .A1(n4759), .A2(n4758), .ZN(n4757) );
  NOR2_X1 U5305 ( .A1(n4762), .A2(n6834), .ZN(n4761) );
  MUX2_X1 U5306 ( .A(n8644), .B(n8574), .S(n8518), .Z(n8513) );
  NOR2_X1 U5307 ( .A1(n5866), .A2(n9598), .ZN(n4567) );
  INV_X1 U5308 ( .A(n5775), .ZN(n4982) );
  OAI21_X1 U5309 ( .B1(n7193), .B2(n4552), .A(n4551), .ZN(n5570) );
  NAND2_X1 U5310 ( .A1(n7193), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U5311 ( .A1(n7832), .A2(n6144), .ZN(n6145) );
  NOR2_X1 U5312 ( .A1(n6184), .A2(n4936), .ZN(n4933) );
  INV_X1 U5313 ( .A(n4434), .ZN(n4937) );
  NAND3_X1 U5314 ( .A1(n4809), .A2(n4808), .A3(n7126), .ZN(n7128) );
  NOR2_X1 U5315 ( .A1(n8898), .A2(n8928), .ZN(n8919) );
  NOR2_X1 U5316 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n4735) );
  OR2_X1 U5317 ( .A1(n6696), .A2(n6803), .ZN(n4711) );
  NOR2_X1 U5318 ( .A1(n4711), .A2(n4707), .ZN(n4706) );
  INV_X1 U5319 ( .A(n6645), .ZN(n4707) );
  INV_X1 U5320 ( .A(n6214), .ZN(n6032) );
  OR2_X1 U5321 ( .A1(n6205), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6214) );
  AND2_X1 U5322 ( .A1(n6751), .A2(n7703), .ZN(n6741) );
  INV_X1 U5323 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U5324 ( .A1(n8876), .A2(n10227), .ZN(n6700) );
  INV_X1 U5325 ( .A(n6921), .ZN(n4780) );
  OR2_X1 U5326 ( .A1(n9392), .A2(n9136), .ZN(n6828) );
  NAND2_X1 U5327 ( .A1(n9179), .A2(n5053), .ZN(n9116) );
  NOR2_X1 U5328 ( .A1(n6814), .A2(n5054), .ZN(n5053) );
  INV_X1 U5329 ( .A(n6695), .ZN(n5054) );
  NAND2_X1 U5330 ( .A1(n6901), .A2(n6900), .ZN(n8112) );
  INV_X1 U5331 ( .A(n6902), .ZN(n5029) );
  OR2_X1 U5332 ( .A1(n6928), .A2(n7827), .ZN(n6433) );
  INV_X1 U5333 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6021) );
  NOR2_X1 U5334 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5971) );
  INV_X1 U5335 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U5336 ( .A1(n5988), .A2(n5987), .ZN(n6255) );
  NOR2_X1 U5337 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5954) );
  INV_X1 U5338 ( .A(n8232), .ZN(n5429) );
  INV_X1 U5339 ( .A(n7931), .ZN(n4874) );
  NAND2_X1 U5340 ( .A1(n4661), .A2(n4660), .ZN(n4665) );
  NAND2_X1 U5341 ( .A1(n8561), .A2(n8632), .ZN(n4661) );
  NAND2_X1 U5342 ( .A1(n4567), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5934) );
  AOI21_X1 U5343 ( .B1(n4643), .B2(n8576), .A(n4642), .ZN(n4646) );
  INV_X1 U5344 ( .A(n5004), .ZN(n4643) );
  INV_X1 U5345 ( .A(n9809), .ZN(n4642) );
  AND2_X1 U5346 ( .A1(n6497), .A2(n8635), .ZN(n5004) );
  OR2_X1 U5347 ( .A1(n9857), .A2(n6493), .ZN(n8490) );
  NOR2_X1 U5348 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  INV_X1 U5349 ( .A(n8410), .ZN(n4656) );
  INV_X1 U5350 ( .A(n8470), .ZN(n4655) );
  INV_X1 U5351 ( .A(n9933), .ZN(n5076) );
  AND2_X1 U5352 ( .A1(n7915), .A2(n7916), .ZN(n4584) );
  NOR2_X1 U5353 ( .A1(n6477), .A2(n5018), .ZN(n5017) );
  INV_X1 U5354 ( .A(n8598), .ZN(n5018) );
  INV_X1 U5355 ( .A(n9627), .ZN(n8030) );
  NAND2_X1 U5356 ( .A1(n9628), .A2(n6478), .ZN(n8437) );
  NAND2_X1 U5357 ( .A1(n4581), .A2(n6546), .ZN(n7657) );
  NAND2_X1 U5358 ( .A1(n6544), .A2(n7768), .ZN(n8593) );
  OR2_X1 U5359 ( .A1(n6537), .A2(n10173), .ZN(n4861) );
  AND2_X1 U5360 ( .A1(n5944), .A2(n5943), .ZN(n6595) );
  INV_X1 U5361 ( .A(n6574), .ZN(n4589) );
  NAND2_X1 U5362 ( .A1(n5062), .A2(n5064), .ZN(n5061) );
  INV_X1 U5363 ( .A(n5065), .ZN(n5062) );
  NAND2_X1 U5364 ( .A1(n6513), .A2(n5127), .ZN(n6605) );
  INV_X1 U5365 ( .A(n6502), .ZN(n4970) );
  AND2_X1 U5366 ( .A1(n6502), .A2(n5891), .ZN(n6500) );
  NAND2_X1 U5367 ( .A1(n5832), .A2(n5831), .ZN(n5857) );
  AND2_X1 U5368 ( .A1(n5144), .A2(n5143), .ZN(n5181) );
  AND2_X1 U5369 ( .A1(n4983), .A2(n4982), .ZN(n4977) );
  AND2_X1 U5370 ( .A1(n4985), .A2(n4982), .ZN(n4980) );
  NAND2_X1 U5371 ( .A1(n5726), .A2(n10386), .ZN(n4989) );
  OR2_X1 U5372 ( .A1(n5726), .A2(n10386), .ZN(n4990) );
  NOR2_X1 U5373 ( .A1(n5161), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n4678) );
  INV_X1 U5374 ( .A(SI_20_), .ZN(n10386) );
  NAND2_X1 U5375 ( .A1(n4768), .A2(n5518), .ZN(n5569) );
  NOR2_X1 U5376 ( .A1(n5519), .A2(n4767), .ZN(n4769) );
  INV_X1 U5377 ( .A(n5022), .ZN(n5021) );
  OR2_X1 U5378 ( .A1(n6012), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U5379 ( .A1(n6012), .A2(n4425), .ZN(n5019) );
  INV_X1 U5380 ( .A(n6344), .ZN(n4945) );
  OR2_X1 U5381 ( .A1(n6369), .A2(n4943), .ZN(n4942) );
  OR2_X1 U5382 ( .A1(n8372), .A2(n4945), .ZN(n4943) );
  XNOR2_X1 U5383 ( .A(n6917), .B(n8711), .ZN(n8812) );
  NAND2_X1 U5384 ( .A1(n7482), .A2(n4962), .ZN(n7513) );
  AND2_X1 U5385 ( .A1(n6311), .A2(n9164), .ZN(n6312) );
  NOR2_X1 U5386 ( .A1(n8771), .A2(n8772), .ZN(n8770) );
  XNOR2_X1 U5387 ( .A(n10204), .B(n6063), .ZN(n6068) );
  NAND2_X1 U5388 ( .A1(n8786), .A2(n8787), .ZN(n8841) );
  NAND2_X1 U5389 ( .A1(n6240), .A2(n9213), .ZN(n4956) );
  INV_X1 U5390 ( .A(n6862), .ZN(n6854) );
  NOR2_X1 U5391 ( .A1(n5048), .A2(n7912), .ZN(n5045) );
  NAND2_X1 U5392 ( .A1(n4475), .A2(n9346), .ZN(n5048) );
  INV_X1 U5393 ( .A(n7827), .ZN(n6953) );
  NAND2_X1 U5394 ( .A1(n6864), .A2(n6867), .ZN(n4574) );
  INV_X1 U5395 ( .A(n6073), .ZN(n6226) );
  NOR2_X1 U5396 ( .A1(n4443), .A2(n7305), .ZN(n4901) );
  NAND2_X1 U5397 ( .A1(n4573), .A2(n7046), .ZN(n7018) );
  INV_X1 U5398 ( .A(n7017), .ZN(n4573) );
  NAND2_X1 U5399 ( .A1(n4889), .A2(n7603), .ZN(n4893) );
  OR2_X1 U5400 ( .A1(n4421), .A2(n7589), .ZN(n4829) );
  OR2_X1 U5401 ( .A1(n7001), .A2(n7603), .ZN(n4828) );
  OR2_X1 U5402 ( .A1(n4892), .A2(n4891), .ZN(n7600) );
  INV_X1 U5403 ( .A(n7022), .ZN(n4891) );
  NAND2_X1 U5404 ( .A1(n7083), .A2(n7859), .ZN(n7085) );
  NAND2_X1 U5405 ( .A1(n7864), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7863) );
  OR2_X1 U5406 ( .A1(n7128), .A2(n7348), .ZN(n4433) );
  NAND2_X1 U5407 ( .A1(n7128), .A2(n7348), .ZN(n7130) );
  INV_X1 U5408 ( .A(n4410), .ZN(n9009) );
  NAND2_X1 U5409 ( .A1(n6396), .A2(n6395), .ZN(n6440) );
  OR2_X1 U5410 ( .A1(n6336), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5411 ( .A1(n6326), .A2(n6325), .ZN(n6336) );
  NAND2_X1 U5412 ( .A1(n6276), .A2(n4429), .ZN(n6316) );
  INV_X1 U5413 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5414 ( .A1(n6276), .A2(n6275), .ZN(n6287) );
  AND2_X1 U5415 ( .A1(n4439), .A2(n6030), .ZN(n4736) );
  INV_X1 U5416 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6030) );
  INV_X1 U5417 ( .A(n6762), .ZN(n6698) );
  NAND2_X1 U5418 ( .A1(n6029), .A2(n4439), .ZN(n6170) );
  INV_X1 U5419 ( .A(n6042), .ZN(n5040) );
  OAI22_X1 U5420 ( .A1(n6087), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n7320), .B2(
        n6041), .ZN(n6042) );
  NOR2_X1 U5421 ( .A1(n6454), .A2(n10239), .ZN(n6955) );
  NAND2_X1 U5422 ( .A1(n8709), .A2(n10235), .ZN(n6936) );
  AND2_X1 U5423 ( .A1(n9364), .A2(n6920), .ZN(n6843) );
  AND2_X1 U5424 ( .A1(n4778), .A2(n4501), .ZN(n4781) );
  NOR2_X1 U5425 ( .A1(n6834), .A2(n6720), .ZN(n5044) );
  INV_X1 U5426 ( .A(n5033), .ZN(n4545) );
  AOI21_X1 U5427 ( .B1(n9104), .B2(n9105), .A(n5034), .ZN(n5033) );
  NOR2_X1 U5428 ( .A1(n9386), .A2(n9126), .ZN(n5034) );
  NAND2_X1 U5429 ( .A1(n9101), .A2(n6722), .ZN(n6651) );
  AND3_X1 U5430 ( .A1(n6267), .A2(n6266), .A3(n6265), .ZN(n9214) );
  NOR2_X1 U5431 ( .A1(n6797), .A2(n4713), .ZN(n4712) );
  INV_X1 U5432 ( .A(n6646), .ZN(n4713) );
  INV_X1 U5433 ( .A(n10239), .ZN(n9329) );
  AND2_X1 U5434 ( .A1(n6426), .A2(n6950), .ZN(n6939) );
  NOR2_X1 U5435 ( .A1(n6461), .A2(n7181), .ZN(n6941) );
  NAND2_X1 U5436 ( .A1(n8024), .A2(n7912), .ZN(n10239) );
  AND2_X1 U5437 ( .A1(n7070), .A2(n7342), .ZN(n7188) );
  AND2_X1 U5438 ( .A1(n6010), .A2(n6009), .ZN(n6406) );
  NAND2_X1 U5439 ( .A1(n6007), .A2(n5967), .ZN(n6010) );
  INV_X1 U5440 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6015) );
  AND2_X1 U5441 ( .A1(n5981), .A2(n6241), .ZN(n8910) );
  AND2_X1 U5442 ( .A1(n6159), .A2(n6158), .ZN(n6192) );
  NAND2_X1 U5443 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4528) );
  NAND2_X1 U5444 ( .A1(n5222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5924) );
  INV_X1 U5445 ( .A(n4435), .ZN(n4722) );
  AOI21_X1 U5446 ( .B1(n4723), .B2(n4722), .A(n4721), .ZN(n4720) );
  NOR2_X1 U5447 ( .A1(n4432), .A2(n5883), .ZN(n4721) );
  AND2_X1 U5448 ( .A1(n5325), .A2(n4730), .ZN(n5331) );
  INV_X1 U5449 ( .A(n8339), .ZN(n4913) );
  AND2_X1 U5450 ( .A1(n9496), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U5451 ( .A1(n5590), .A2(n8339), .ZN(n4912) );
  NAND2_X1 U5452 ( .A1(n7628), .A2(n7627), .ZN(n9528) );
  NAND2_X1 U5453 ( .A1(n5330), .A2(n5329), .ZN(n7444) );
  OR2_X1 U5454 ( .A1(n5327), .A2(n8738), .ZN(n5330) );
  NAND2_X1 U5455 ( .A1(n4570), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5812) );
  AOI21_X1 U5456 ( .B1(n4681), .B2(n4683), .A(n4471), .ZN(n4680) );
  NAND2_X1 U5457 ( .A1(n8381), .A2(n8383), .ZN(n8380) );
  INV_X1 U5458 ( .A(n9567), .ZN(n9593) );
  NAND2_X1 U5459 ( .A1(n5587), .A2(n5586), .ZN(n8338) );
  AOI21_X1 U5460 ( .B1(n8517), .B2(n9760), .A(n4627), .ZN(n4626) );
  AND4_X1 U5461 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(n8341)
         );
  AND4_X1 U5462 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n8161)
         );
  AND4_X1 U5463 ( .A1(n5275), .A2(n5272), .A3(n5273), .A4(n5274), .ZN(n6475)
         );
  OR2_X1 U5464 ( .A1(n7682), .A2(n4876), .ZN(n4875) );
  AND2_X1 U5465 ( .A1(n7673), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4876) );
  AOI21_X1 U5466 ( .B1(n9684), .B2(P1_REG1_REG_15__SCAN_IN), .A(n4445), .ZN(
        n9687) );
  NOR2_X1 U5467 ( .A1(n5121), .A2(n6573), .ZN(n5065) );
  OAI21_X1 U5468 ( .B1(n5005), .B2(n4647), .A(n4646), .ZN(n9805) );
  AND2_X1 U5469 ( .A1(n8580), .A2(n8637), .ZN(n9809) );
  NAND2_X1 U5470 ( .A1(n5005), .A2(n5004), .ZN(n9829) );
  AND2_X1 U5471 ( .A1(n8494), .A2(n8635), .ZN(n9837) );
  NOR2_X1 U5472 ( .A1(n9857), .A2(n5001), .ZN(n5000) );
  INV_X1 U5473 ( .A(n5002), .ZN(n5001) );
  NAND2_X1 U5474 ( .A1(n5088), .A2(n5085), .ZN(n9855) );
  AND2_X1 U5475 ( .A1(n5086), .A2(n8528), .ZN(n5085) );
  INV_X1 U5476 ( .A(n5094), .ZN(n5093) );
  OR2_X1 U5477 ( .A1(n8530), .A2(n8529), .ZN(n9871) );
  OR2_X1 U5478 ( .A1(n10018), .A2(n9617), .ZN(n5097) );
  NOR2_X1 U5479 ( .A1(n6567), .A2(n5099), .ZN(n5098) );
  INV_X1 U5480 ( .A(n6565), .ZN(n5099) );
  AND2_X1 U5481 ( .A1(n8479), .A2(n8625), .ZN(n8555) );
  INV_X1 U5482 ( .A(n8475), .ZN(n4658) );
  AOI21_X1 U5483 ( .B1(n4657), .B2(n4656), .A(n4655), .ZN(n4649) );
  NAND2_X1 U5484 ( .A1(n5073), .A2(n4603), .ZN(n4602) );
  NOR2_X1 U5485 ( .A1(n4459), .A2(n5079), .ZN(n5078) );
  NOR2_X1 U5486 ( .A1(n6561), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U5487 ( .A1(n6560), .A2(n6559), .ZN(n5080) );
  NOR2_X1 U5488 ( .A1(n6561), .A2(n5082), .ZN(n5081) );
  INV_X1 U5489 ( .A(n6559), .ZN(n5082) );
  NAND2_X1 U5490 ( .A1(n4572), .A2(n4571), .ZN(n9950) );
  INV_X1 U5491 ( .A(n10042), .ZN(n4571) );
  OR2_X1 U5492 ( .A1(n8532), .A2(n9929), .ZN(n9955) );
  NAND2_X1 U5493 ( .A1(n9962), .A2(n9968), .ZN(n5014) );
  NAND2_X1 U5494 ( .A1(n8158), .A2(n6553), .ZN(n4592) );
  AND2_X1 U5495 ( .A1(n8419), .A2(n6478), .ZN(n4991) );
  NAND2_X1 U5496 ( .A1(n4992), .A2(n8419), .ZN(n7922) );
  NAND2_X1 U5497 ( .A1(n9992), .A2(n5687), .ZN(n6597) );
  NAND2_X1 U5498 ( .A1(n6977), .A2(n6590), .ZN(n4580) );
  AND2_X1 U5499 ( .A1(n7823), .A2(n7777), .ZN(n9992) );
  INV_X1 U5500 ( .A(n4606), .ZN(n4605) );
  AND2_X1 U5501 ( .A1(n7777), .A2(n8571), .ZN(n10181) );
  OR2_X1 U5502 ( .A1(n8518), .A2(n8675), .ZN(n10170) );
  AND2_X1 U5503 ( .A1(n8026), .A2(n8584), .ZN(n7777) );
  NOR2_X1 U5504 ( .A1(n4637), .A2(n5176), .ZN(n4636) );
  INV_X1 U5505 ( .A(n5146), .ZN(n4637) );
  NOR2_X2 U5506 ( .A1(n5141), .A2(n5176), .ZN(n5144) );
  NAND2_X1 U5507 ( .A1(n4678), .A2(n4919), .ZN(n5212) );
  OAI21_X1 U5508 ( .B1(n5727), .B2(n4985), .A(n4983), .ZN(n5776) );
  NAND2_X1 U5509 ( .A1(n4919), .A2(n4448), .ZN(n4677) );
  NAND2_X1 U5510 ( .A1(n4976), .A2(n5656), .ZN(n5678) );
  XNOR2_X1 U5511 ( .A(n5208), .B(n4967), .ZN(n5205) );
  INV_X1 U5512 ( .A(SI_4_), .ZN(n4967) );
  AND2_X1 U5513 ( .A1(n6363), .A2(n6362), .ZN(n8817) );
  AOI21_X1 U5514 ( .B1(n9141), .B2(n6659), .A(n6320), .ZN(n9153) );
  INV_X1 U5515 ( .A(n4948), .ZN(n4947) );
  OAI21_X1 U5516 ( .B1(n4951), .B2(n4949), .A(n6322), .ZN(n4948) );
  INV_X1 U5517 ( .A(n9095), .ZN(n8790) );
  NAND2_X1 U5518 ( .A1(n8797), .A2(n8796), .ZN(n8795) );
  AND2_X1 U5519 ( .A1(n8314), .A2(n6234), .ZN(n6235) );
  NAND2_X1 U5520 ( .A1(n4959), .A2(n4458), .ZN(n4958) );
  AND2_X1 U5521 ( .A1(n6378), .A2(n6377), .ZN(n8849) );
  AND2_X1 U5522 ( .A1(n6430), .A2(n6429), .ZN(n6952) );
  INV_X1 U5523 ( .A(n8849), .ZN(n9083) );
  INV_X1 U5524 ( .A(n8817), .ZN(n9109) );
  NAND2_X1 U5525 ( .A1(n6293), .A2(n6292), .ZN(n9187) );
  INV_X1 U5526 ( .A(n9214), .ZN(n6269) );
  AND2_X1 U5527 ( .A1(n7073), .A2(n9450), .ZN(n8761) );
  INV_X1 U5528 ( .A(n9020), .ZN(n8978) );
  NAND2_X1 U5529 ( .A1(n6996), .A2(n7374), .ZN(n4814) );
  NAND2_X1 U5530 ( .A1(n7000), .A2(n7154), .ZN(n7158) );
  AOI21_X1 U5531 ( .B1(n8978), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8977), .ZN(
        n4820) );
  OR2_X1 U5532 ( .A1(n9004), .A2(n4823), .ZN(n4822) );
  NAND2_X1 U5533 ( .A1(n8974), .A2(n8973), .ZN(n4824) );
  NAND2_X1 U5534 ( .A1(n5037), .A2(n4420), .ZN(n4764) );
  OAI22_X1 U5535 ( .A1(n6087), .A2(n7174), .B1(n6041), .B2(n7297), .ZN(n6088)
         );
  NOR2_X1 U5536 ( .A1(n7542), .A2(n7541), .ZN(n10209) );
  NAND2_X1 U5537 ( .A1(n7188), .A2(n6955), .ZN(n9240) );
  INV_X1 U5538 ( .A(n8714), .ZN(n9352) );
  NAND2_X1 U5539 ( .A1(n9041), .A2(n9040), .ZN(n9042) );
  XNOR2_X1 U5540 ( .A(n9038), .B(n9037), .ZN(n9043) );
  NAND2_X1 U5541 ( .A1(n9062), .A2(n9236), .ZN(n9040) );
  NAND2_X1 U5542 ( .A1(n9073), .A2(n4698), .ZN(n4692) );
  NAND2_X1 U5543 ( .A1(n4783), .A2(n4782), .ZN(n9068) );
  XNOR2_X1 U5544 ( .A(n5993), .B(n6299), .ZN(n9017) );
  NAND2_X1 U5545 ( .A1(n5783), .A2(n5782), .ZN(n9844) );
  NAND2_X1 U5546 ( .A1(n7192), .A2(n6615), .ZN(n4612) );
  NAND2_X1 U5547 ( .A1(n5872), .A2(n5871), .ZN(n9610) );
  OR2_X1 U5548 ( .A1(n9813), .A2(n6521), .ZN(n5846) );
  NAND2_X1 U5549 ( .A1(n4884), .A2(n7237), .ZN(n9678) );
  OR2_X1 U5550 ( .A1(n10127), .A2(n9662), .ZN(n4884) );
  AND2_X1 U5551 ( .A1(n4872), .A2(n4482), .ZN(n7431) );
  AOI21_X1 U5552 ( .B1(n9747), .B2(n10135), .A(n10139), .ZN(n4864) );
  OR2_X1 U5553 ( .A1(n9746), .A2(n10128), .ZN(n4865) );
  INV_X1 U5554 ( .A(n9729), .ZN(n10135) );
  INV_X1 U5555 ( .A(n10128), .ZN(n9744) );
  NOR2_X1 U5556 ( .A1(n9749), .A2(n9750), .ZN(n4867) );
  NAND2_X1 U5557 ( .A1(n8561), .A2(n8687), .ZN(n4669) );
  OR2_X1 U5558 ( .A1(n6597), .A2(n8567), .ZN(n9913) );
  NAND2_X1 U5559 ( .A1(n10194), .A2(n10181), .ZN(n10036) );
  INV_X1 U5560 ( .A(n8519), .ZN(n9755) );
  NAND2_X1 U5561 ( .A1(n6513), .A2(n6512), .ZN(n6517) );
  NAND2_X1 U5562 ( .A1(n5658), .A2(n5218), .ZN(n5219) );
  NOR2_X2 U5563 ( .A1(n7070), .A2(n6983), .ZN(P2_U3893) );
  NAND2_X1 U5564 ( .A1(n4794), .A2(n9053), .ZN(n4793) );
  NOR2_X1 U5565 ( .A1(n8590), .A2(n8518), .ZN(n4858) );
  NAND2_X1 U5566 ( .A1(n6763), .A2(n6762), .ZN(n6757) );
  NOR2_X1 U5567 ( .A1(n8439), .A2(n4835), .ZN(n4837) );
  NAND2_X1 U5568 ( .A1(n4838), .A2(n8443), .ZN(n4835) );
  NOR2_X1 U5569 ( .A1(n8445), .A2(n4840), .ZN(n4838) );
  INV_X1 U5570 ( .A(n8443), .ZN(n4608) );
  NAND2_X1 U5571 ( .A1(n8443), .A2(n4842), .ZN(n4841) );
  INV_X1 U5572 ( .A(n8438), .ZN(n4842) );
  OAI21_X1 U5573 ( .B1(n8432), .B2(n8590), .A(n4856), .ZN(n8431) );
  MUX2_X1 U5574 ( .A(n6772), .B(n6771), .S(n6984), .Z(n6773) );
  MUX2_X1 U5575 ( .A(n8457), .B(n8456), .S(n8518), .Z(n8466) );
  NAND2_X1 U5576 ( .A1(n8466), .A2(n8612), .ZN(n4616) );
  NAND2_X1 U5577 ( .A1(n8466), .A2(n8617), .ZN(n4621) );
  NAND2_X1 U5578 ( .A1(n8469), .A2(n8468), .ZN(n4850) );
  NAND2_X1 U5579 ( .A1(n8467), .A2(n8521), .ZN(n4849) );
  NAND2_X1 U5580 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  NOR2_X1 U5581 ( .A1(n4851), .A2(n8616), .ZN(n4614) );
  NAND2_X1 U5582 ( .A1(n4616), .A2(n8617), .ZN(n4615) );
  OR2_X1 U5583 ( .A1(n8461), .A2(n8518), .ZN(n4851) );
  NAND2_X1 U5584 ( .A1(n4619), .A2(n4618), .ZN(n4617) );
  NOR2_X1 U5585 ( .A1(n8620), .A2(n8521), .ZN(n4618) );
  NAND2_X1 U5586 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5587 ( .A1(n8464), .A2(n8465), .ZN(n4620) );
  NAND2_X1 U5588 ( .A1(n6821), .A2(n6984), .ZN(n4748) );
  NAND2_X1 U5589 ( .A1(n4750), .A2(n9053), .ZN(n4749) );
  OAI21_X1 U5590 ( .B1(n6819), .B2(n6818), .A(n4752), .ZN(n4751) );
  AND2_X1 U5591 ( .A1(n6816), .A2(n6817), .ZN(n4752) );
  NOR2_X1 U5592 ( .A1(n6833), .A2(n4422), .ZN(n4759) );
  INV_X1 U5593 ( .A(n8471), .ZN(n8478) );
  AND2_X1 U5594 ( .A1(n4422), .A2(n4491), .ZN(n4756) );
  INV_X1 U5595 ( .A(n5518), .ZN(n4775) );
  OR2_X1 U5596 ( .A1(n7187), .A2(n6422), .ZN(n6453) );
  INV_X1 U5597 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5985) );
  INV_X1 U5598 ( .A(n9501), .ZN(n4908) );
  AND2_X1 U5599 ( .A1(n8519), .A2(n4845), .ZN(n4844) );
  INV_X1 U5600 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U5601 ( .B1(n9760), .B2(n8518), .A(n9606), .ZN(n4846) );
  AOI21_X1 U5602 ( .B1(n6554), .B2(n4595), .A(n4594), .ZN(n4593) );
  INV_X1 U5603 ( .A(n6553), .ZN(n4595) );
  INV_X1 U5604 ( .A(n6556), .ZN(n4594) );
  NOR2_X1 U5605 ( .A1(n4409), .A2(n7649), .ZN(n4582) );
  NAND2_X1 U5606 ( .A1(n9630), .A2(n8425), .ZN(n8597) );
  INV_X1 U5607 ( .A(n5743), .ZN(n5744) );
  INV_X1 U5608 ( .A(n4776), .ZN(n4773) );
  NAND2_X1 U5609 ( .A1(n4975), .A2(n4973), .ZN(n5497) );
  NOR2_X1 U5610 ( .A1(n5494), .A2(n4974), .ZN(n4973) );
  INV_X1 U5611 ( .A(n5435), .ZN(n4974) );
  OAI21_X1 U5612 ( .B1(n7193), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n5366), .ZN(
        n5368) );
  NAND2_X1 U5613 ( .A1(n7193), .A2(n7214), .ZN(n5366) );
  INV_X1 U5614 ( .A(n5348), .ZN(n5351) );
  INV_X1 U5615 ( .A(n5349), .ZN(n5350) );
  OAI21_X1 U5616 ( .B1(n5966), .B2(P2_IR_REG_27__SCAN_IN), .A(n5969), .ZN(
        n5022) );
  NAND2_X1 U5617 ( .A1(n9346), .A2(n9030), .ZN(n6862) );
  INV_X1 U5618 ( .A(n6863), .ZN(n6690) );
  OR2_X1 U5619 ( .A1(n6858), .A2(n6856), .ZN(n6853) );
  AND2_X1 U5620 ( .A1(n7013), .A2(n7287), .ZN(n7328) );
  NAND2_X1 U5621 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  AOI21_X1 U5622 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8958), .A(n8957), .ZN(
        n8959) );
  NOR2_X1 U5623 ( .A1(n8945), .A2(n8980), .ZN(n8965) );
  INV_X1 U5624 ( .A(n4695), .ZN(n4694) );
  AND2_X1 U5625 ( .A1(n6315), .A2(n10380), .ZN(n6326) );
  INV_X1 U5626 ( .A(n6316), .ZN(n6315) );
  AND2_X1 U5627 ( .A1(n6275), .A2(n4744), .ZN(n4743) );
  INV_X1 U5628 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4744) );
  AND2_X1 U5629 ( .A1(n6262), .A2(n10383), .ZN(n6276) );
  INV_X1 U5630 ( .A(n6263), .ZN(n6262) );
  NOR2_X1 U5631 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4740) );
  INV_X1 U5632 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5633 ( .A1(n8007), .A2(n8013), .ZN(n6762) );
  OR2_X1 U5634 ( .A1(n9358), .A2(n8723), .ZN(n6848) );
  OR2_X1 U5635 ( .A1(n9375), .A2(n8790), .ZN(n6835) );
  INV_X1 U5636 ( .A(n6828), .ZN(n4703) );
  CLKBUF_X1 U5637 ( .A(n8112), .Z(n4544) );
  INV_X1 U5638 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5990) );
  INV_X1 U5639 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5984) );
  OAI22_X1 U5640 ( .A1(n5382), .A2(n7818), .B1(n5900), .B2(n7651), .ZN(n4905)
         );
  OR2_X1 U5641 ( .A1(n8738), .A2(n7651), .ZN(n4904) );
  OR2_X1 U5642 ( .A1(n5488), .A2(n8199), .ZN(n5489) );
  NOR2_X1 U5643 ( .A1(n8514), .A2(n4557), .ZN(n4556) );
  INV_X1 U5644 ( .A(n4625), .ZN(n4557) );
  INV_X1 U5645 ( .A(n8513), .ZN(n4624) );
  AND2_X1 U5646 ( .A1(n8667), .A2(n8516), .ZN(n8517) );
  NAND2_X1 U5647 ( .A1(n4628), .A2(n8670), .ZN(n4627) );
  NAND2_X1 U5648 ( .A1(n4844), .A2(n6608), .ZN(n4628) );
  NOR2_X1 U5649 ( .A1(n9767), .A2(n4995), .ZN(n4994) );
  INV_X1 U5650 ( .A(n4996), .ZN(n4995) );
  NOR2_X1 U5651 ( .A1(n9782), .A2(n9981), .ZN(n4996) );
  NOR2_X1 U5652 ( .A1(n9876), .A2(n10014), .ZN(n5002) );
  INV_X1 U5653 ( .A(n8529), .ZN(n5087) );
  NOR2_X1 U5654 ( .A1(n8529), .A2(n5090), .ZN(n5089) );
  INV_X1 U5655 ( .A(n5091), .ZN(n5090) );
  NAND2_X1 U5656 ( .A1(n4604), .A2(n4600), .ZN(n4597) );
  AOI21_X1 U5657 ( .B1(n9968), .B2(n6556), .A(n4463), .ZN(n5100) );
  NAND2_X1 U5658 ( .A1(n4593), .A2(n4596), .ZN(n4591) );
  INV_X1 U5659 ( .A(n6554), .ZN(n4596) );
  NAND2_X1 U5660 ( .A1(n5012), .A2(n6555), .ZN(n5011) );
  INV_X1 U5661 ( .A(n8035), .ZN(n4999) );
  OR2_X1 U5662 ( .A1(n5409), .A2(n5383), .ZN(n5470) );
  CLKBUF_X1 U5663 ( .A(n7948), .Z(n8035) );
  AND2_X1 U5664 ( .A1(n5886), .A2(n5863), .ZN(n5884) );
  AND2_X1 U5665 ( .A1(n5858), .A2(n5836), .ZN(n5856) );
  AND2_X1 U5666 ( .A1(n5831), .A2(n5806), .ZN(n5829) );
  INV_X1 U5667 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5138) );
  INV_X1 U5668 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10408) );
  INV_X1 U5669 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4916) );
  INV_X1 U5670 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5671 ( .A1(n7193), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U5672 ( .A1(n4754), .A2(n4753), .ZN(n4975) );
  AND2_X1 U5673 ( .A1(n5464), .A2(n5432), .ZN(n4753) );
  INV_X1 U5674 ( .A(SI_19_), .ZN(n10379) );
  NAND2_X1 U5675 ( .A1(n7757), .A2(n6145), .ZN(n7829) );
  NAND2_X1 U5677 ( .A1(n4936), .A2(n4434), .ZN(n4935) );
  NOR2_X1 U5678 ( .A1(n6184), .A2(n8870), .ZN(n4550) );
  NAND2_X1 U5679 ( .A1(n4938), .A2(n4937), .ZN(n4931) );
  INV_X1 U5680 ( .A(n8772), .ZN(n4949) );
  OR2_X1 U5681 ( .A1(n6321), .A2(n9125), .ZN(n6322) );
  INV_X1 U5682 ( .A(n4951), .ZN(n4950) );
  NAND2_X1 U5683 ( .A1(n8795), .A2(n4939), .ZN(n8802) );
  NOR2_X1 U5684 ( .A1(n8805), .A2(n4940), .ZN(n4939) );
  INV_X1 U5685 ( .A(n6270), .ZN(n4940) );
  AND2_X1 U5686 ( .A1(n6231), .A2(n8210), .ZN(n4565) );
  XNOR2_X1 U5687 ( .A(n9338), .B(n6063), .ZN(n6056) );
  NAND2_X1 U5688 ( .A1(n7607), .A2(n4960), .ZN(n4959) );
  INV_X1 U5689 ( .A(n6099), .ZN(n4960) );
  NOR2_X1 U5690 ( .A1(n5049), .A2(n5047), .ZN(n5046) );
  NAND2_X1 U5691 ( .A1(n6867), .A2(n4797), .ZN(n5047) );
  NOR2_X1 U5692 ( .A1(n6690), .A2(n9346), .ZN(n5049) );
  AND2_X1 U5693 ( .A1(n6687), .A2(n6686), .ZN(n6689) );
  AND2_X1 U5694 ( .A1(n6687), .A2(n6664), .ZN(n8719) );
  AND2_X1 U5695 ( .A1(n6447), .A2(n6446), .ZN(n8712) );
  NAND2_X1 U5696 ( .A1(n6122), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U5697 ( .A(n7169), .B(n10213), .ZN(n8884) );
  AND2_X1 U5698 ( .A1(n7282), .A2(n4819), .ZN(n7331) );
  NAND2_X1 U5699 ( .A1(n4539), .A2(n7046), .ZN(n4538) );
  INV_X1 U5700 ( .A(n6999), .ZN(n4539) );
  NAND2_X1 U5701 ( .A1(n4517), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U5702 ( .A1(n7158), .A2(n4421), .ZN(n4833) );
  NAND2_X1 U5703 ( .A1(n7158), .A2(n7001), .ZN(n4826) );
  OR2_X1 U5704 ( .A1(n4832), .A2(n4831), .ZN(n7586) );
  NAND2_X1 U5705 ( .A1(n4833), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4832) );
  INV_X1 U5706 ( .A(n7004), .ZN(n4831) );
  INV_X1 U5707 ( .A(n7085), .ZN(n4812) );
  OR2_X1 U5708 ( .A1(n7083), .A2(n7859), .ZN(n7084) );
  NAND2_X1 U5709 ( .A1(n4564), .A2(n8155), .ZN(n7121) );
  INV_X1 U5710 ( .A(n7120), .ZN(n4564) );
  NAND2_X1 U5711 ( .A1(n4502), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7122) );
  NOR2_X1 U5712 ( .A1(n8899), .A2(n8919), .ZN(n8900) );
  XNOR2_X1 U5713 ( .A(n8913), .B(n4815), .ZN(n8914) );
  INV_X1 U5714 ( .A(n8928), .ZN(n4815) );
  NAND2_X1 U5715 ( .A1(n8914), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8939) );
  INV_X1 U5716 ( .A(n9017), .ZN(n9000) );
  OR2_X1 U5717 ( .A1(n6440), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U5718 ( .A1(n6347), .A2(n4506), .ZN(n6397) );
  INV_X1 U5719 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5720 ( .A1(n6347), .A2(n4735), .ZN(n6381) );
  NAND2_X1 U5721 ( .A1(n6347), .A2(n10416), .ZN(n6372) );
  OR2_X1 U5722 ( .A1(n6356), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6358) );
  AOI21_X1 U5723 ( .B1(n9129), .B2(n6659), .A(n6331), .ZN(n9136) );
  NAND2_X1 U5724 ( .A1(n6276), .A2(n4743), .ZN(n6304) );
  NAND2_X1 U5725 ( .A1(n9179), .A2(n6695), .ZN(n9173) );
  AND2_X1 U5726 ( .A1(n9181), .A2(n9183), .ZN(n4541) );
  INV_X1 U5727 ( .A(n4710), .ZN(n4709) );
  OAI21_X1 U5728 ( .B1(n4712), .B2(n4711), .A(n6647), .ZN(n4710) );
  NAND2_X1 U5729 ( .A1(n6246), .A2(n6245), .ZN(n6263) );
  INV_X1 U5730 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6245) );
  INV_X1 U5731 ( .A(n6247), .ZN(n6246) );
  NAND2_X1 U5732 ( .A1(n6032), .A2(n4738), .ZN(n6247) );
  AND2_X1 U5733 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5734 ( .A1(n6032), .A2(n4740), .ZN(n6225) );
  NAND2_X1 U5735 ( .A1(n6032), .A2(n6031), .ZN(n6223) );
  OR2_X1 U5736 ( .A1(n8109), .A2(n8096), .ZN(n8092) );
  OR2_X1 U5737 ( .A1(n6186), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6205) );
  INV_X1 U5738 ( .A(n8869), .ZN(n9258) );
  AND2_X1 U5739 ( .A1(n8092), .A2(n6763), .ZN(n8111) );
  NAND2_X1 U5740 ( .A1(n6029), .A2(n6028), .ZN(n6168) );
  INV_X1 U5741 ( .A(n10202), .ZN(n9256) );
  INV_X1 U5742 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4745) );
  AND2_X1 U5743 ( .A1(n6754), .A2(n7747), .ZN(n7885) );
  NAND2_X1 U5744 ( .A1(n7547), .A2(n6026), .ZN(n6109) );
  OR2_X1 U5745 ( .A1(n6701), .A2(n6700), .ZN(n7618) );
  OR2_X1 U5746 ( .A1(n10198), .A2(n4461), .ZN(n6886) );
  OR2_X1 U5747 ( .A1(n6072), .A2(n10213), .ZN(n6065) );
  AND2_X1 U5748 ( .A1(n7522), .A2(n6932), .ZN(n8098) );
  AND2_X1 U5749 ( .A1(n6954), .A2(n6984), .ZN(n7529) );
  AND3_X1 U5750 ( .A1(n6951), .A2(n6950), .A3(n6949), .ZN(n7533) );
  AND2_X1 U5751 ( .A1(n9030), .A2(n9029), .ZN(n9344) );
  NAND2_X1 U5752 ( .A1(n9039), .A2(n10199), .ZN(n9041) );
  OAI21_X1 U5753 ( .B1(n4781), .B2(n4780), .A(n4462), .ZN(n4777) );
  NAND2_X1 U5754 ( .A1(n6450), .A2(n6041), .ZN(n9050) );
  INV_X1 U5755 ( .A(n9364), .ZN(n4732) );
  NAND2_X1 U5756 ( .A1(n4700), .A2(n6840), .ZN(n9059) );
  NAND2_X1 U5757 ( .A1(n4701), .A2(n6839), .ZN(n4700) );
  INV_X1 U5758 ( .A(n9073), .ZN(n4701) );
  OR2_X1 U5759 ( .A1(n9081), .A2(n6919), .ZN(n4783) );
  AND2_X1 U5760 ( .A1(n6835), .A2(n6838), .ZN(n9082) );
  AND2_X1 U5761 ( .A1(n6355), .A2(n6354), .ZN(n6917) );
  NAND2_X1 U5762 ( .A1(n6314), .A2(n6313), .ZN(n8823) );
  AND2_X1 U5763 ( .A1(n9309), .A2(n9187), .ZN(n9147) );
  OAI21_X2 U5764 ( .B1(n9224), .B2(n6911), .A(n6910), .ZN(n9212) );
  NAND2_X1 U5765 ( .A1(n9050), .A2(n9053), .ZN(n9261) );
  NAND2_X1 U5766 ( .A1(n5052), .A2(n5050), .ZN(n9249) );
  NOR2_X1 U5767 ( .A1(n9255), .A2(n5051), .ZN(n5050) );
  INV_X1 U5768 ( .A(n6775), .ZN(n5051) );
  NAND2_X1 U5769 ( .A1(n5026), .A2(n5030), .ZN(n9252) );
  NAND2_X1 U5770 ( .A1(n4544), .A2(n6902), .ZN(n5026) );
  NAND2_X1 U5771 ( .A1(n6301), .A2(n4537), .ZN(n4788) );
  NOR2_X1 U5772 ( .A1(n4423), .A2(n5055), .ZN(n5056) );
  INV_X1 U5773 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6011) );
  AND2_X1 U5774 ( .A1(n5962), .A2(n6424), .ZN(n4686) );
  AND2_X1 U5775 ( .A1(n6259), .A2(n6271), .ZN(n8937) );
  INV_X1 U5776 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U5777 ( .A1(n4533), .A2(n4531), .ZN(n6077) );
  NAND2_X1 U5778 ( .A1(n4532), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U5779 ( .A1(n4534), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4533) );
  INV_X1 U5780 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4532) );
  INV_X1 U5781 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5406) );
  AND2_X1 U5782 ( .A1(n5558), .A2(n5540), .ZN(n4671) );
  XNOR2_X1 U5783 ( .A(n5267), .B(n4426), .ZN(n5268) );
  AND2_X1 U5784 ( .A1(n5404), .A2(n5403), .ZN(n8235) );
  INV_X1 U5785 ( .A(n9543), .ZN(n4922) );
  OR2_X1 U5786 ( .A1(n5812), .A2(n5811), .ZN(n5840) );
  INV_X1 U5787 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5605) );
  INV_X1 U5788 ( .A(n4569), .ZN(n5639) );
  NAND2_X1 U5789 ( .A1(n9494), .A2(n5619), .ZN(n9511) );
  NAND3_X1 U5790 ( .A1(n9554), .A2(n5773), .A3(n4431), .ZN(n9458) );
  NAND2_X1 U5791 ( .A1(n5342), .A2(n9528), .ZN(n9533) );
  NAND2_X1 U5792 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5270) );
  OR2_X1 U5793 ( .A1(n5692), .A2(n5691), .ZN(n5711) );
  INV_X1 U5794 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9548) );
  INV_X1 U5795 ( .A(n5527), .ZN(n5525) );
  INV_X1 U5796 ( .A(n5488), .ZN(n8301) );
  NAND2_X1 U5797 ( .A1(n4569), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U5798 ( .A1(n5676), .A2(n5675), .ZN(n9564) );
  INV_X1 U5799 ( .A(n5673), .ZN(n5676) );
  OR2_X1 U5800 ( .A1(n5942), .A2(n8567), .ZN(n5950) );
  INV_X1 U5801 ( .A(n7823), .ZN(n8675) );
  AND2_X1 U5802 ( .A1(n5224), .A2(n6529), .ZN(n8671) );
  AND4_X1 U5803 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n8160)
         );
  NAND2_X1 U5804 ( .A1(n5410), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U5805 ( .A1(n6620), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5806 ( .A1(n4853), .A2(n10109), .ZN(n4854) );
  AND2_X1 U5807 ( .A1(n8755), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4853) );
  OR2_X1 U5808 ( .A1(n7474), .A2(n7475), .ZN(n4872) );
  INV_X1 U5809 ( .A(n4872), .ZN(n7473) );
  OR2_X1 U5810 ( .A1(n7436), .A2(n7437), .ZN(n7434) );
  OR2_X1 U5811 ( .A1(n7567), .A2(n7568), .ZN(n7672) );
  OR2_X1 U5812 ( .A1(n7687), .A2(n7688), .ZN(n7685) );
  INV_X1 U5813 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U5814 ( .A1(n4873), .A2(n4518), .ZN(n9685) );
  NOR2_X1 U5815 ( .A1(n4665), .A2(n8687), .ZN(n4659) );
  NAND2_X1 U5816 ( .A1(n4670), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U5817 ( .A1(n9811), .A2(n9801), .ZN(n9796) );
  AND2_X1 U5818 ( .A1(n5934), .A2(n5895), .ZN(n9783) );
  AND2_X1 U5819 ( .A1(n5894), .A2(n5867), .ZN(n9798) );
  INV_X1 U5820 ( .A(n9825), .ZN(n6497) );
  NAND2_X1 U5821 ( .A1(n9887), .A2(n5002), .ZN(n9874) );
  INV_X1 U5822 ( .A(n4570), .ZN(n5753) );
  NAND2_X1 U5823 ( .A1(n4653), .A2(n4651), .ZN(n6488) );
  INV_X1 U5824 ( .A(n4652), .ZN(n4651) );
  INV_X1 U5825 ( .A(n5072), .ZN(n5071) );
  OAI21_X1 U5826 ( .B1(n5076), .B2(n5078), .A(n6562), .ZN(n5072) );
  NOR2_X1 U5827 ( .A1(n5076), .A2(n5077), .ZN(n5074) );
  INV_X1 U5828 ( .A(n5081), .ZN(n5077) );
  INV_X1 U5829 ( .A(n5576), .ZN(n5577) );
  NAND2_X1 U5830 ( .A1(n5576), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5606) );
  NOR2_X2 U5831 ( .A1(n9950), .A2(n10039), .ZN(n9948) );
  NAND2_X1 U5832 ( .A1(n4568), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5527) );
  INV_X1 U5833 ( .A(n5501), .ZN(n4568) );
  NAND2_X1 U5834 ( .A1(n4999), .A2(n6588), .ZN(n8170) );
  NAND2_X1 U5835 ( .A1(n4424), .A2(n4451), .ZN(n5016) );
  NAND2_X1 U5836 ( .A1(n9627), .A2(n8243), .ZN(n8436) );
  NAND2_X1 U5837 ( .A1(n4583), .A2(n6550), .ZN(n7965) );
  INV_X1 U5838 ( .A(n6478), .ZN(n7978) );
  NAND2_X1 U5839 ( .A1(n7659), .A2(n5017), .ZN(n7918) );
  NAND2_X1 U5840 ( .A1(n6476), .A2(n8600), .ZN(n7660) );
  NAND2_X1 U5841 ( .A1(n7660), .A2(n7661), .ZN(n7659) );
  INV_X1 U5842 ( .A(n8536), .ZN(n7649) );
  NOR2_X2 U5843 ( .A1(n7817), .A2(n10180), .ZN(n7816) );
  NOR2_X1 U5844 ( .A1(n7811), .A2(n4648), .ZN(n5008) );
  NAND2_X1 U5845 ( .A1(n7724), .A2(n4861), .ZN(n7641) );
  NAND2_X1 U5846 ( .A1(n10173), .A2(n7448), .ZN(n7735) );
  NAND2_X1 U5847 ( .A1(n6538), .A2(n7780), .ZN(n7726) );
  AOI21_X1 U5848 ( .B1(n5063), .B2(n5059), .A(n4589), .ZN(n4585) );
  NAND2_X1 U5849 ( .A1(n5068), .A2(n5059), .ZN(n4586) );
  OAI21_X1 U5850 ( .B1(n8251), .B2(n6560), .A(n6559), .ZN(n9956) );
  NAND2_X1 U5851 ( .A1(n8159), .A2(n10170), .ZN(n10055) );
  INV_X1 U5852 ( .A(n7718), .ZN(n6627) );
  OR2_X1 U5853 ( .A1(n7721), .A2(n6598), .ZN(n6628) );
  INV_X1 U5854 ( .A(n10055), .ZN(n10185) );
  OAI21_X1 U5855 ( .B1(n6503), .B2(n4971), .A(n4968), .ZN(n4972) );
  INV_X1 U5856 ( .A(n6510), .ZN(n4971) );
  AOI21_X1 U5857 ( .B1(n6510), .B2(n4970), .A(n4969), .ZN(n4968) );
  INV_X1 U5858 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U5859 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5174) );
  AOI21_X1 U5860 ( .B1(n4980), .B2(n4983), .A(n4979), .ZN(n4978) );
  INV_X1 U5861 ( .A(n5774), .ZN(n4979) );
  AND2_X1 U5862 ( .A1(n5801), .A2(n5780), .ZN(n5799) );
  NAND2_X1 U5863 ( .A1(n4988), .A2(n4989), .ZN(n5746) );
  NAND2_X1 U5864 ( .A1(n4676), .A2(n4675), .ZN(n5170) );
  NAND2_X1 U5865 ( .A1(n10426), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U5866 ( .A1(n5633), .A2(n10408), .ZN(n5658) );
  AOI21_X1 U5867 ( .B1(n4919), .B2(n4918), .A(n4917), .ZN(n5601) );
  AND2_X1 U5868 ( .A1(n5217), .A2(n4916), .ZN(n4917) );
  NOR2_X1 U5869 ( .A1(n5161), .A2(n4915), .ZN(n4918) );
  NAND2_X1 U5870 ( .A1(n4916), .A2(n4674), .ZN(n4915) );
  NAND2_X1 U5871 ( .A1(n5212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5573) );
  XNOR2_X1 U5872 ( .A(n5544), .B(n5564), .ZN(n7354) );
  OR2_X1 U5873 ( .A1(n5465), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5874 ( .A1(n4754), .A2(n5432), .ZN(n5463) );
  CLKBUF_X1 U5875 ( .A(n5246), .Z(n5247) );
  OR2_X1 U5876 ( .A1(n5276), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5877 ( .A1(n8313), .A2(n6238), .ZN(n8276) );
  XNOR2_X1 U5878 ( .A(n8811), .B(n8812), .ZN(n8813) );
  AND2_X1 U5879 ( .A1(n8717), .A2(n5105), .ZN(n8718) );
  AND2_X1 U5880 ( .A1(n6342), .A2(n6341), .ZN(n8782) );
  OR2_X1 U5881 ( .A1(n6369), .A2(n4945), .ZN(n4944) );
  AND2_X1 U5882 ( .A1(n4942), .A2(n6368), .ZN(n4941) );
  INV_X1 U5883 ( .A(n8874), .ZN(n7610) );
  NAND2_X1 U5884 ( .A1(n7513), .A2(n6099), .ZN(n7608) );
  NAND2_X1 U5885 ( .A1(n8795), .A2(n6270), .ZN(n8804) );
  AND2_X1 U5886 ( .A1(n7482), .A2(n6084), .ZN(n7514) );
  AND2_X1 U5887 ( .A1(n6310), .A2(n6309), .ZN(n9135) );
  NOR2_X1 U5888 ( .A1(n8770), .A2(n6312), .ZN(n8825) );
  OR2_X1 U5889 ( .A1(n8770), .A2(n4951), .ZN(n8824) );
  INV_X1 U5890 ( .A(n8848), .ZN(n8859) );
  INV_X1 U5891 ( .A(n9237), .ZN(n8284) );
  INV_X1 U5892 ( .A(n8208), .ZN(n6199) );
  AND3_X1 U5893 ( .A1(n6281), .A2(n6280), .A3(n6279), .ZN(n9199) );
  INV_X1 U5894 ( .A(n8863), .ZN(n8317) );
  AND2_X1 U5895 ( .A1(n6435), .A2(n6434), .ZN(n8853) );
  NAND2_X1 U5896 ( .A1(n6439), .A2(n9240), .ZN(n8851) );
  AND2_X1 U5897 ( .A1(n8857), .A2(n4956), .ZN(n4953) );
  AND2_X1 U5898 ( .A1(n4957), .A2(n4956), .ZN(n8858) );
  INV_X1 U5899 ( .A(n8853), .ZN(n8855) );
  NAND2_X1 U5900 ( .A1(n7343), .A2(n8063), .ZN(n8863) );
  INV_X1 U5901 ( .A(n6689), .ZN(n9030) );
  INV_X1 U5902 ( .A(n8719), .ZN(n9039) );
  INV_X1 U5903 ( .A(n8712), .ZN(n9051) );
  INV_X1 U5904 ( .A(n8782), .ZN(n9126) );
  INV_X1 U5905 ( .A(n9153), .ZN(n9125) );
  INV_X1 U5906 ( .A(n9135), .ZN(n9164) );
  INV_X1 U5907 ( .A(n9199), .ZN(n9163) );
  OR2_X1 U5908 ( .A1(n6670), .A2(n7589), .ZN(n6165) );
  NAND4_X2 U5909 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n8872)
         );
  NOR2_X1 U5910 ( .A1(n4450), .A2(n6113), .ZN(n6114) );
  NOR2_X1 U5911 ( .A1(n6095), .A2(n5119), .ZN(n6096) );
  INV_X1 U5912 ( .A(n7579), .ZN(n7397) );
  INV_X1 U5913 ( .A(P2_U3893), .ZN(n8877) );
  OR2_X1 U5914 ( .A1(n7325), .A2(n7326), .ZN(n7323) );
  OR2_X1 U5915 ( .A1(n7364), .A2(n7363), .ZN(n7456) );
  NAND2_X1 U5916 ( .A1(n7055), .A2(n7150), .ZN(n7590) );
  NAND2_X1 U5917 ( .A1(n4895), .A2(n4896), .ZN(n7161) );
  AOI21_X1 U5918 ( .B1(n7159), .B2(n4897), .A(n4514), .ZN(n4896) );
  NAND2_X1 U5919 ( .A1(n4893), .A2(n7022), .ZN(n7598) );
  NAND2_X1 U5920 ( .A1(n7004), .A2(n4833), .ZN(n7588) );
  NOR2_X1 U5921 ( .A1(n7202), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4830) );
  AND2_X1 U5922 ( .A1(n4829), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U5923 ( .A1(n7063), .A2(n7064), .ZN(n7855) );
  AOI21_X1 U5924 ( .B1(n7130), .B2(n9324), .A(n4516), .ZN(n4816) );
  NOR2_X1 U5925 ( .A1(n8999), .A2(n8998), .ZN(n9001) );
  NAND2_X1 U5926 ( .A1(n6286), .A2(n6285), .ZN(n9170) );
  NAND2_X1 U5927 ( .A1(n6301), .A2(n6993), .ZN(n6106) );
  INV_X1 U5928 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U5929 ( .A1(n6301), .A2(n4787), .ZN(n4786) );
  INV_X1 U5930 ( .A(n9204), .ZN(n9265) );
  INV_X1 U5931 ( .A(n7344), .ZN(n7537) );
  NAND2_X1 U5932 ( .A1(n6666), .A2(n6665), .ZN(n9347) );
  NAND2_X1 U5933 ( .A1(n4779), .A2(n4781), .ZN(n9061) );
  NAND2_X1 U5934 ( .A1(n9081), .A2(n4782), .ZN(n4779) );
  INV_X1 U5935 ( .A(n6917), .ZN(n9380) );
  NAND2_X1 U5936 ( .A1(n6274), .A2(n6273), .ZN(n9406) );
  AND2_X1 U5937 ( .A1(n9189), .A2(n9188), .ZN(n9405) );
  AOI21_X1 U5938 ( .B1(n4714), .B2(n4712), .A(n6696), .ZN(n4708) );
  NAND2_X1 U5939 ( .A1(n4714), .A2(n6646), .ZN(n9222) );
  NAND2_X1 U5940 ( .A1(n6410), .A2(n6409), .ZN(n7528) );
  INV_X1 U5941 ( .A(n7188), .ZN(n7181) );
  AND2_X1 U5942 ( .A1(n7068), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7342) );
  NAND2_X1 U5943 ( .A1(n7188), .A2(n7187), .ZN(n7215) );
  INV_X1 U5944 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8333) );
  INV_X1 U5945 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8270) );
  INV_X1 U5946 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8221) );
  INV_X1 U5947 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8025) );
  INV_X1 U5948 ( .A(n6952), .ZN(n8024) );
  INV_X1 U5949 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7910) );
  INV_X1 U5950 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7635) );
  INV_X1 U5951 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7551) );
  INV_X1 U5952 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7409) );
  INV_X1 U5953 ( .A(n8937), .ZN(n8958) );
  AND2_X1 U5954 ( .A1(n4411), .A2(P2_U3151), .ZN(n9453) );
  INV_X1 U5955 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7339) );
  INV_X1 U5956 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U5957 ( .A1(n4529), .A2(n4527), .ZN(n6040) );
  NAND2_X1 U5958 ( .A1(n4807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U5959 ( .A1(n4528), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4527) );
  XNOR2_X1 U5960 ( .A(n5927), .B(n5926), .ZN(n7219) );
  NAND2_X1 U5961 ( .A1(n5925), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U5962 ( .A1(n4720), .A2(n4724), .ZN(n4719) );
  AND2_X1 U5963 ( .A1(n4720), .A2(n4495), .ZN(n4718) );
  NAND2_X1 U5964 ( .A1(n8069), .A2(n5540), .ZN(n8327) );
  NAND2_X1 U5965 ( .A1(n9554), .A2(n5773), .ZN(n9460) );
  AND2_X1 U5966 ( .A1(n8744), .A2(n5931), .ZN(n4561) );
  NAND2_X1 U5967 ( .A1(n5337), .A2(n5336), .ZN(n8382) );
  AND2_X1 U5968 ( .A1(n5333), .A2(n5332), .ZN(n8381) );
  NAND2_X1 U5969 ( .A1(n4920), .A2(n4921), .ZN(n9480) );
  AND2_X1 U5970 ( .A1(n4914), .A2(n8337), .ZN(n9495) );
  NAND2_X1 U5971 ( .A1(n8338), .A2(n8339), .ZN(n4914) );
  NAND2_X1 U5972 ( .A1(n4926), .A2(n9467), .ZN(n9546) );
  NAND2_X1 U5973 ( .A1(n4928), .A2(n4927), .ZN(n4926) );
  INV_X1 U5974 ( .A(n4535), .ZN(n4928) );
  NAND2_X1 U5975 ( .A1(n5752), .A2(n5751), .ZN(n9857) );
  NAND2_X1 U5976 ( .A1(n8380), .A2(n8382), .ZN(n7628) );
  NAND2_X1 U5977 ( .A1(n9591), .A2(n9590), .ZN(n4536) );
  INV_X1 U5978 ( .A(n9602), .ZN(n9558) );
  INV_X1 U5979 ( .A(n8527), .ZN(n8520) );
  OR2_X1 U5980 ( .A1(n8652), .A2(n8563), .ZN(n8564) );
  NAND2_X1 U5981 ( .A1(n5759), .A2(n5758), .ZN(n9614) );
  NAND2_X1 U5982 ( .A1(n5124), .A2(n5414), .ZN(n9628) );
  NAND2_X1 U5983 ( .A1(n5936), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5414) );
  AOI21_X1 U5984 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(n10127) );
  AND2_X1 U5985 ( .A1(n4883), .A2(n4882), .ZN(n9675) );
  INV_X1 U5986 ( .A(n9676), .ZN(n4882) );
  INV_X1 U5987 ( .A(n4880), .ZN(n7276) );
  OAI21_X1 U5988 ( .B1(n9675), .B2(n7263), .A(n4881), .ZN(n4880) );
  AOI21_X1 U5989 ( .B1(n7267), .B2(n10454), .A(n7238), .ZN(n4881) );
  INV_X1 U5990 ( .A(n4871), .ZN(n7556) );
  NAND2_X1 U5991 ( .A1(n4869), .A2(n4868), .ZN(n7557) );
  NAND2_X1 U5992 ( .A1(n7563), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4868) );
  INV_X1 U5993 ( .A(n7555), .ZN(n4870) );
  INV_X1 U5994 ( .A(n4875), .ZN(n7932) );
  XNOR2_X1 U5995 ( .A(n9685), .B(n7938), .ZN(n9684) );
  OR2_X1 U5996 ( .A1(n9706), .A2(n9707), .ZN(n9727) );
  OR2_X1 U5997 ( .A1(n10120), .A2(n8566), .ZN(n9729) );
  OR2_X1 U5998 ( .A1(n9731), .A2(n9730), .ZN(n9741) );
  AND2_X1 U5999 ( .A1(n7220), .A2(n7239), .ZN(n10122) );
  NAND2_X1 U6000 ( .A1(n6975), .A2(n8747), .ZN(n9768) );
  NAND2_X1 U6001 ( .A1(n6970), .A2(n8561), .ZN(n6971) );
  INV_X1 U6002 ( .A(n4580), .ZN(n9769) );
  INV_X1 U6003 ( .A(n5058), .ZN(n9787) );
  AOI21_X1 U6004 ( .B1(n5068), .B2(n5065), .A(n5063), .ZN(n5058) );
  INV_X1 U6005 ( .A(n9777), .ZN(n9778) );
  NAND2_X1 U6006 ( .A1(n9776), .A2(n9964), .ZN(n9779) );
  NAND2_X1 U6007 ( .A1(n5066), .A2(n5070), .ZN(n9794) );
  NAND2_X1 U6008 ( .A1(n5068), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U6009 ( .A1(n8580), .A2(n9805), .ZN(n9791) );
  NAND2_X1 U6010 ( .A1(n9829), .A2(n8576), .ZN(n9806) );
  NAND2_X1 U6011 ( .A1(n5005), .A2(n8635), .ZN(n9826) );
  OAI21_X1 U6012 ( .B1(n6566), .B2(n5093), .A(n5091), .ZN(n9872) );
  NAND2_X1 U6013 ( .A1(n5096), .A2(n5097), .ZN(n9882) );
  NAND2_X1 U6014 ( .A1(n6566), .A2(n5098), .ZN(n5096) );
  NAND2_X1 U6015 ( .A1(n6566), .A2(n6565), .ZN(n8396) );
  INV_X1 U6016 ( .A(n4657), .ZN(n4650) );
  NAND2_X1 U6017 ( .A1(n5635), .A2(n5634), .ZN(n9917) );
  NAND2_X1 U6018 ( .A1(n5075), .A2(n5078), .ZN(n9934) );
  NAND2_X1 U6019 ( .A1(n8251), .A2(n5081), .ZN(n5075) );
  NAND2_X1 U6020 ( .A1(n10056), .A2(n6556), .ZN(n8130) );
  AND2_X1 U6021 ( .A1(n5014), .A2(n8454), .ZN(n8121) );
  OR2_X1 U6022 ( .A1(n9967), .A2(n9968), .ZN(n10056) );
  NAND2_X1 U6023 ( .A1(n7947), .A2(n7946), .ZN(n7945) );
  NAND2_X1 U6024 ( .A1(n8032), .A2(n6552), .ZN(n7947) );
  INV_X1 U6025 ( .A(n7922), .ZN(n6587) );
  AND2_X1 U6026 ( .A1(n9951), .A2(n7785), .ZN(n10163) );
  INV_X1 U6027 ( .A(n10157), .ZN(n9953) );
  NAND2_X1 U6028 ( .A1(n7722), .A2(n9913), .ZN(n9951) );
  OR2_X1 U6029 ( .A1(n7721), .A2(n7720), .ZN(n7722) );
  AND2_X1 U6030 ( .A1(n9951), .A2(n7732), .ZN(n10157) );
  INV_X1 U6031 ( .A(n9913), .ZN(n10154) );
  INV_X1 U6032 ( .A(n9844), .ZN(n10078) );
  INV_X1 U6033 ( .A(n9936), .ZN(n10097) );
  OR2_X1 U6034 ( .A1(n10047), .A2(n10046), .ZN(n10099) );
  INV_X1 U6035 ( .A(n8205), .ZN(n6588) );
  NAND2_X1 U6036 ( .A1(n7219), .A2(n5928), .ZN(n8567) );
  AND2_X1 U6037 ( .A1(n4562), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5928) );
  NAND4_X1 U6038 ( .A1(n5144), .A2(n5143), .A3(n4440), .A4(n5147), .ZN(n10104)
         );
  INV_X1 U6039 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U6040 ( .A1(n4640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4639) );
  INV_X1 U6041 ( .A(n5141), .ZN(n4638) );
  INV_X1 U6042 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8334) );
  INV_X1 U6043 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U6044 ( .A1(n5179), .A2(n5178), .ZN(n8220) );
  MUX2_X1 U6045 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5177), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5179) );
  INV_X1 U6046 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8219) );
  INV_X1 U6047 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8068) );
  INV_X1 U6048 ( .A(n5224), .ZN(n8026) );
  INV_X1 U6049 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7909) );
  INV_X1 U6050 ( .A(n6529), .ZN(n8584) );
  INV_X1 U6051 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8370) );
  INV_X1 U6052 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10607) );
  NOR2_X1 U6053 ( .A1(n7193), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10106) );
  INV_X1 U6054 ( .A(n5205), .ZN(n4966) );
  INV_X1 U6055 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6056 ( .A1(n7073), .A2(n6041), .ZN(n6986) );
  AND3_X1 U6057 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(n6880) );
  NAND2_X1 U6058 ( .A1(n7300), .A2(n4813), .ZN(n7307) );
  NAND2_X1 U6059 ( .A1(n4822), .A2(n9006), .ZN(n4821) );
  NAND2_X1 U6060 ( .A1(n4763), .A2(n8710), .ZN(P2_U3204) );
  NAND2_X1 U6061 ( .A1(n4764), .A2(n10212), .ZN(n4763) );
  NAND2_X1 U6062 ( .A1(n6964), .A2(n6963), .ZN(n6965) );
  NAND2_X1 U6063 ( .A1(n9275), .A2(n9274), .ZN(n9277) );
  NAND2_X1 U6064 ( .A1(n9285), .A2(n4542), .ZN(P2_U3484) );
  INV_X1 U6065 ( .A(n4543), .ZN(n4542) );
  OAI21_X1 U6066 ( .B1(n9373), .B2(n9332), .A(n9284), .ZN(n4543) );
  NAND2_X1 U6067 ( .A1(n6964), .A2(n6946), .ZN(n6947) );
  NOR2_X1 U6068 ( .A1(n4867), .A2(n4523), .ZN(n4866) );
  OR2_X1 U6069 ( .A1(n9755), .A2(n10036), .ZN(n5101) );
  OAI21_X1 U6070 ( .B1(n4993), .B2(n10036), .A(n6599), .ZN(n6600) );
  OR2_X1 U6071 ( .A1(n9755), .A2(n10096), .ZN(n5102) );
  OR2_X1 U6072 ( .A1(n9370), .A2(n8849), .ZN(n6839) );
  OR2_X1 U6073 ( .A1(n9542), .A2(n4925), .ZN(n4924) );
  AND2_X1 U6074 ( .A1(n6848), .A2(n6849), .ZN(n4418) );
  AND2_X1 U6075 ( .A1(n6935), .A2(n6934), .ZN(n4420) );
  AND2_X1 U6076 ( .A1(n7001), .A2(n7603), .ZN(n4421) );
  OR2_X1 U6077 ( .A1(n4762), .A2(n6984), .ZN(n4422) );
  NAND2_X1 U6078 ( .A1(n5972), .A2(n5971), .ZN(n4423) );
  AND2_X1 U6079 ( .A1(n8596), .A2(n8602), .ZN(n4424) );
  AND2_X1 U6080 ( .A1(n5966), .A2(n4455), .ZN(n4425) );
  AND2_X1 U6081 ( .A1(n5266), .A2(n4904), .ZN(n4426) );
  INV_X1 U6082 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9439) );
  AND3_X1 U6083 ( .A1(n4498), .A2(n4611), .A3(n4610), .ZN(n7959) );
  INV_X1 U6084 ( .A(n7959), .ZN(n4609) );
  INV_X1 U6085 ( .A(n4924), .ZN(n4923) );
  INV_X1 U6086 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4674) );
  INV_X1 U6087 ( .A(n5121), .ZN(n5069) );
  NOR2_X1 U6088 ( .A1(n5118), .A2(n4485), .ZN(n4427) );
  NAND2_X1 U6089 ( .A1(n9233), .A2(n6645), .ZN(n4714) );
  AND2_X1 U6090 ( .A1(n4433), .A2(n7130), .ZN(n4428) );
  AND2_X1 U6091 ( .A1(n4743), .A2(n4742), .ZN(n4429) );
  INV_X1 U6092 ( .A(n5410), .ZN(n5816) );
  XNOR2_X1 U6093 ( .A(n5283), .B(n4966), .ZN(n6085) );
  NAND2_X1 U6094 ( .A1(n9811), .A2(n4994), .ZN(n6590) );
  OR2_X1 U6095 ( .A1(n8913), .A2(n8928), .ZN(n4430) );
  NAND2_X1 U6096 ( .A1(n5795), .A2(n5796), .ZN(n4431) );
  XOR2_X1 U6097 ( .A(n8743), .B(n8742), .Z(n4432) );
  NAND2_X1 U6098 ( .A1(n9887), .A2(n9894), .ZN(n9873) );
  XNOR2_X1 U6099 ( .A(n6537), .B(n7733), .ZN(n7723) );
  AND2_X1 U6100 ( .A1(n6185), .A2(n6147), .ZN(n4434) );
  AND2_X1 U6101 ( .A1(n5878), .A2(n5855), .ZN(n4435) );
  AND2_X1 U6102 ( .A1(n5009), .A2(n8465), .ZN(n4436) );
  AND3_X1 U6103 ( .A1(n5959), .A2(n5960), .A3(n5961), .ZN(n4437) );
  INV_X1 U6104 ( .A(n8576), .ZN(n4647) );
  OR2_X1 U6105 ( .A1(n6085), .A2(n6518), .ZN(n4438) );
  INV_X1 U6106 ( .A(n6475), .ZN(n6544) );
  OAI21_X1 U6107 ( .B1(n8373), .B2(n4944), .A(n4941), .ZN(n8786) );
  OR2_X1 U6108 ( .A1(n10053), .A2(n8161), .ZN(n8454) );
  AND2_X1 U6109 ( .A1(n6028), .A2(n4737), .ZN(n4439) );
  OAI21_X1 U6110 ( .B1(n9116), .B2(n4704), .A(n4702), .ZN(n9101) );
  OAI21_X1 U6111 ( .B1(n9928), .B2(n8620), .A(n8410), .ZN(n9918) );
  OAI21_X1 U6112 ( .B1(n9928), .B2(n4650), .A(n4649), .ZN(n9905) );
  AND2_X1 U6113 ( .A1(n5146), .A2(n5183), .ZN(n4440) );
  NAND2_X1 U6114 ( .A1(n4602), .A2(n6563), .ZN(n9897) );
  NAND2_X1 U6115 ( .A1(n6651), .A2(n6719), .ZN(n9092) );
  NAND2_X1 U6116 ( .A1(n4692), .A2(n4695), .ZN(n9036) );
  NAND2_X1 U6117 ( .A1(n5073), .A2(n5071), .ZN(n9912) );
  AND2_X1 U6118 ( .A1(n6728), .A2(n6984), .ZN(n4441) );
  INV_X1 U6119 ( .A(n8687), .ZN(n4668) );
  INV_X1 U6120 ( .A(n7046), .ZN(n7460) );
  AND2_X1 U6121 ( .A1(n6936), .A2(n10245), .ZN(n4442) );
  XNOR2_X1 U6122 ( .A(n6024), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6025) );
  AND2_X1 U6123 ( .A1(n7297), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4443) );
  NOR4_X1 U6124 ( .A1(n9854), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n4444)
         );
  AND2_X1 U6125 ( .A1(n9685), .A2(n9692), .ZN(n4445) );
  NAND2_X1 U6126 ( .A1(n5040), .A2(n5039), .ZN(n9338) );
  NAND2_X1 U6127 ( .A1(n4428), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7129) );
  AND2_X1 U6128 ( .A1(n10014), .A2(n9616), .ZN(n4446) );
  OR2_X1 U6129 ( .A1(n9782), .A2(n9594), .ZN(n8630) );
  OR2_X1 U6130 ( .A1(n9812), .A2(n6498), .ZN(n8580) );
  INV_X1 U6131 ( .A(n8580), .ZN(n5007) );
  INV_X1 U6132 ( .A(n7574), .ZN(n6699) );
  INV_X1 U6133 ( .A(n7169), .ZN(n4787) );
  INV_X1 U6134 ( .A(n8692), .ZN(n4993) );
  NOR2_X1 U6135 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6152) );
  OR2_X1 U6136 ( .A1(n9767), .A2(n8739), .ZN(n8573) );
  NAND3_X2 U6137 ( .A1(n6019), .A2(n6020), .A3(n6411), .ZN(n6063) );
  OR2_X1 U6138 ( .A1(n6924), .A2(n8723), .ZN(n4447) );
  NOR2_X1 U6139 ( .A1(n5162), .A2(n5163), .ZN(n4448) );
  OR2_X1 U6140 ( .A1(n6254), .A2(n6804), .ZN(n4449) );
  NOR2_X1 U6141 ( .A1(n6670), .A2(n10254), .ZN(n4450) );
  INV_X1 U6142 ( .A(n9069), .ZN(n6920) );
  NAND2_X1 U6143 ( .A1(n4733), .A2(n6386), .ZN(n9069) );
  AND2_X1 U6144 ( .A1(n8454), .A2(n8613), .ZN(n9968) );
  INV_X1 U6145 ( .A(n9968), .ZN(n6555) );
  OR2_X1 U6146 ( .A1(n9386), .A2(n8782), .ZN(n6719) );
  AND2_X1 U6147 ( .A1(n8540), .A2(n5017), .ZN(n4451) );
  AND2_X1 U6148 ( .A1(n6511), .A2(n6510), .ZN(n4452) );
  INV_X1 U6149 ( .A(n9468), .ZN(n4927) );
  INV_X1 U6150 ( .A(n9981), .ZN(n9801) );
  AND2_X1 U6151 ( .A1(n5011), .A2(n8463), .ZN(n4453) );
  AND2_X1 U6152 ( .A1(n4783), .A2(n4784), .ZN(n4454) );
  INV_X1 U6153 ( .A(n4698), .ZN(n4697) );
  NOR2_X1 U6154 ( .A1(n5042), .A2(n4699), .ZN(n4698) );
  AND2_X1 U6155 ( .A1(n5967), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U6156 ( .A1(n9917), .A2(n9619), .ZN(n4456) );
  AND2_X1 U6157 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4457) );
  NAND2_X1 U6158 ( .A1(n6117), .A2(n7517), .ZN(n4458) );
  NOR2_X1 U6159 ( .A1(n9954), .A2(n8411), .ZN(n4459) );
  AND2_X1 U6160 ( .A1(n4773), .A2(n4765), .ZN(n4460) );
  AND2_X1 U6161 ( .A1(n5040), .A2(n5039), .ZN(n4461) );
  INV_X1 U6162 ( .A(n4785), .ZN(n4784) );
  AND2_X1 U6163 ( .A1(n5956), .A2(n5955), .ZN(n6154) );
  INV_X1 U6164 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5183) );
  OR2_X1 U6165 ( .A1(n9364), .A2(n9069), .ZN(n4462) );
  INV_X1 U6166 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U6167 ( .A1(n4432), .A2(n5883), .ZN(n4724) );
  NOR2_X1 U6168 ( .A1(n10049), .A2(n9623), .ZN(n4463) );
  AND2_X1 U6169 ( .A1(n6839), .A2(n6840), .ZN(n9074) );
  INV_X1 U6170 ( .A(n9074), .ZN(n4758) );
  AND2_X1 U6171 ( .A1(n9352), .A2(n8712), .ZN(n4464) );
  INV_X1 U6172 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7559) );
  AND3_X1 U6173 ( .A1(n6050), .A2(n6049), .A3(n6048), .ZN(n4465) );
  OR2_X1 U6174 ( .A1(n8439), .A2(n4608), .ZN(n4466) );
  AND2_X1 U6175 ( .A1(n6917), .A2(n9109), .ZN(n6834) );
  AND2_X1 U6176 ( .A1(n4854), .A2(n4855), .ZN(n4467) );
  INV_X1 U6177 ( .A(n6573), .ZN(n5067) );
  NAND2_X1 U6178 ( .A1(n9117), .A2(n9115), .ZN(n4468) );
  OR2_X1 U6179 ( .A1(n9981), .A2(n9610), .ZN(n4469) );
  AND2_X1 U6180 ( .A1(n5744), .A2(SI_21_), .ZN(n4470) );
  INV_X1 U6181 ( .A(n8561), .ZN(n4670) );
  NAND2_X1 U6182 ( .A1(n5768), .A2(n5767), .ZN(n4471) );
  OR2_X1 U6183 ( .A1(n5564), .A2(n5567), .ZN(n4472) );
  NAND2_X1 U6184 ( .A1(n6077), .A2(n6100), .ZN(n7171) );
  INV_X1 U6185 ( .A(n7171), .ZN(n4537) );
  AND2_X1 U6186 ( .A1(n4921), .A2(n5767), .ZN(n4473) );
  INV_X1 U6187 ( .A(n5060), .ZN(n5059) );
  NAND2_X1 U6188 ( .A1(n9786), .A2(n5061), .ZN(n5060) );
  NAND2_X1 U6189 ( .A1(n9069), .A2(n4732), .ZN(n6845) );
  INV_X1 U6190 ( .A(n6845), .ZN(n5041) );
  NAND2_X1 U6191 ( .A1(n4469), .A2(n5070), .ZN(n4474) );
  OR2_X1 U6192 ( .A1(n9347), .A2(n9030), .ZN(n4475) );
  AND2_X1 U6193 ( .A1(n5679), .A2(n5656), .ZN(n4476) );
  NOR2_X1 U6194 ( .A1(n4689), .A2(n5974), .ZN(n6423) );
  AND2_X1 U6195 ( .A1(n9121), .A2(n9139), .ZN(n4477) );
  OR2_X1 U6196 ( .A1(n5041), .A2(n6843), .ZN(n9060) );
  INV_X1 U6197 ( .A(n9060), .ZN(n4578) );
  AND3_X1 U6198 ( .A1(n6077), .A2(n6990), .A3(n6100), .ZN(n4478) );
  AND2_X1 U6199 ( .A1(n4994), .A2(n4993), .ZN(n4479) );
  NOR2_X1 U6200 ( .A1(n8205), .A2(n9626), .ZN(n4480) );
  AND2_X1 U6201 ( .A1(n4782), .A2(n6921), .ZN(n4481) );
  NOR2_X1 U6202 ( .A1(n7430), .A2(n7433), .ZN(n4482) );
  INV_X1 U6203 ( .A(n5496), .ZN(n4767) );
  AND2_X1 U6204 ( .A1(n5100), .A2(n4591), .ZN(n4483) );
  INV_X1 U6205 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5975) );
  AND2_X1 U6206 ( .A1(n4566), .A2(n4820), .ZN(n4484) );
  AND2_X1 U6207 ( .A1(n9328), .A2(n9237), .ZN(n4485) );
  NAND2_X1 U6208 ( .A1(n9252), .A2(n9251), .ZN(n4486) );
  AND2_X1 U6209 ( .A1(n6719), .A2(n6722), .ZN(n9103) );
  OR2_X1 U6210 ( .A1(n5623), .A2(SI_16_), .ZN(n4487) );
  AND2_X1 U6211 ( .A1(n4424), .A2(n5017), .ZN(n4488) );
  OR2_X1 U6212 ( .A1(n4761), .A2(n4760), .ZN(n4489) );
  AND2_X1 U6213 ( .A1(n5311), .A2(n4854), .ZN(n4490) );
  OR2_X1 U6214 ( .A1(n4760), .A2(n6836), .ZN(n4491) );
  NOR2_X1 U6215 ( .A1(n8205), .A2(n10062), .ZN(n4998) );
  AND2_X1 U6216 ( .A1(n4741), .A2(n6848), .ZN(n4492) );
  AND2_X1 U6217 ( .A1(n9201), .A2(n4541), .ZN(n4493) );
  AND2_X1 U6218 ( .A1(n5128), .A2(n6899), .ZN(n4494) );
  OR2_X1 U6219 ( .A1(n4432), .A2(n4722), .ZN(n4495) );
  AND2_X1 U6220 ( .A1(n6800), .A2(n9211), .ZN(n4496) );
  AND2_X1 U6221 ( .A1(n5395), .A2(n5396), .ZN(n4497) );
  AND2_X1 U6222 ( .A1(n5387), .A2(n5388), .ZN(n4498) );
  AND2_X1 U6223 ( .A1(n4850), .A2(n4849), .ZN(n4499) );
  AND2_X1 U6224 ( .A1(n4791), .A2(n4793), .ZN(n4500) );
  INV_X1 U6225 ( .A(n5031), .ZN(n5030) );
  NAND2_X1 U6226 ( .A1(n5032), .A2(n6904), .ZN(n5031) );
  OR2_X1 U6227 ( .A1(n9370), .A2(n9083), .ZN(n4501) );
  INV_X1 U6228 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6424) );
  INV_X1 U6229 ( .A(n5064), .ZN(n5063) );
  NAND2_X1 U6230 ( .A1(n4474), .A2(n5069), .ZN(n5064) );
  INV_X2 U6231 ( .A(n9951), .ZN(n10167) );
  NAND2_X1 U6232 ( .A1(n4826), .A2(n7202), .ZN(n7004) );
  AND2_X1 U6233 ( .A1(n7121), .A2(n7123), .ZN(n4502) );
  NAND2_X1 U6234 ( .A1(n5014), .A2(n5012), .ZN(n8120) );
  AND2_X1 U6235 ( .A1(n4999), .A2(n4998), .ZN(n4503) );
  NAND2_X1 U6236 ( .A1(n6889), .A2(n6888), .ZN(n7545) );
  NAND2_X1 U6237 ( .A1(n5035), .A2(n6899), .ZN(n7872) );
  INV_X1 U6238 ( .A(n4708), .ZN(n9209) );
  NAND2_X1 U6239 ( .A1(n7659), .A2(n8598), .ZN(n7799) );
  INV_X1 U6240 ( .A(n8602), .ZN(n4840) );
  INV_X1 U6241 ( .A(n8155), .ZN(n7348) );
  INV_X1 U6242 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U6243 ( .A1(n6474), .A2(n4416), .ZN(n8589) );
  INV_X1 U6244 ( .A(n8589), .ZN(n4648) );
  AND2_X1 U6245 ( .A1(n7422), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4504) );
  INV_X1 U6246 ( .A(n9467), .ZN(n4925) );
  OR2_X1 U6247 ( .A1(n10069), .A2(n10096), .ZN(n4505) );
  INV_X1 U6248 ( .A(n6406), .ZN(n6408) );
  NAND2_X1 U6249 ( .A1(n4592), .A2(n6554), .ZN(n9967) );
  AND2_X1 U6250 ( .A1(n4735), .A2(n4734), .ZN(n4506) );
  AND2_X1 U6251 ( .A1(n5052), .A2(n6775), .ZN(n4507) );
  AND2_X1 U6252 ( .A1(n9511), .A2(n9512), .ZN(n4508) );
  NOR2_X1 U6253 ( .A1(n6678), .A2(n6655), .ZN(n4509) );
  OR2_X1 U6254 ( .A1(n5246), .A2(n5161), .ZN(n4510) );
  INV_X1 U6255 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6031) );
  OR2_X1 U6256 ( .A1(n10069), .A2(n10036), .ZN(n4511) );
  AND2_X1 U6257 ( .A1(n7829), .A2(n6147), .ZN(n4512) );
  INV_X1 U6258 ( .A(n9964), .ZN(n9945) );
  NAND2_X1 U6259 ( .A1(n6530), .A2(n8523), .ZN(n9964) );
  NAND2_X1 U6260 ( .A1(n5223), .A2(n5687), .ZN(n7730) );
  AND2_X1 U6261 ( .A1(n7810), .A2(n7811), .ZN(n4513) );
  XOR2_X1 U6262 ( .A(n7162), .B(P2_REG2_REG_8__SCAN_IN), .Z(n4514) );
  XNOR2_X1 U6263 ( .A(n6056), .B(n10198), .ZN(n7395) );
  NAND2_X1 U6264 ( .A1(n6887), .A2(n6886), .ZN(n10196) );
  XOR2_X1 U6265 ( .A(n8910), .B(P2_REG2_REG_14__SCAN_IN), .Z(n4515) );
  XOR2_X1 U6266 ( .A(n8910), .B(P2_REG1_REG_14__SCAN_IN), .Z(n4516) );
  AND2_X1 U6267 ( .A1(n8761), .A2(n4410), .ZN(n9006) );
  AND2_X1 U6268 ( .A1(n7018), .A2(n7159), .ZN(n4517) );
  INV_X1 U6269 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n4811) );
  NAND2_X1 U6270 ( .A1(n8761), .A2(n9009), .ZN(n9027) );
  INV_X1 U6271 ( .A(n6514), .ZN(n4969) );
  OR2_X1 U6272 ( .A1(n7929), .A2(n7930), .ZN(n4518) );
  AOI21_X1 U6273 ( .B1(n7797), .B2(n7795), .A(n6547), .ZN(n7913) );
  INV_X1 U6274 ( .A(n6633), .ZN(n7573) );
  OR2_X1 U6275 ( .A1(n8878), .A2(n7537), .ZN(n6633) );
  AND2_X1 U6276 ( .A1(n8586), .A2(n8589), .ZN(n4519) );
  INV_X1 U6277 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4739) );
  INV_X1 U6278 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6153) );
  XOR2_X1 U6279 ( .A(n7125), .B(P2_REG1_REG_12__SCAN_IN), .Z(n4520) );
  NAND2_X1 U6280 ( .A1(n4818), .A2(n7171), .ZN(n7282) );
  INV_X1 U6281 ( .A(n5154), .ZN(n8755) );
  AND2_X1 U6282 ( .A1(n5687), .A2(n8675), .ZN(n4521) );
  AND2_X1 U6283 ( .A1(n6041), .A2(P2_B_REG_SCAN_IN), .ZN(n4522) );
  AND2_X1 U6284 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n4523) );
  INV_X1 U6285 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4879) );
  INV_X1 U6286 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U6287 ( .A1(n5677), .A2(n9564), .ZN(n9470) );
  NAND2_X1 U6288 ( .A1(n7997), .A2(n7998), .ZN(n7996) );
  XNOR2_X1 U6289 ( .A(n4905), .B(n8734), .ZN(n5267) );
  OR2_X1 U6290 ( .A1(n5168), .A2(n5217), .ZN(n5169) );
  INV_X1 U6291 ( .A(n9530), .ZN(n4910) );
  NAND2_X1 U6292 ( .A1(n4524), .A2(n4580), .ZN(n4579) );
  NAND2_X1 U6293 ( .A1(n9763), .A2(n10055), .ZN(n4524) );
  NAND2_X1 U6294 ( .A1(n4772), .A2(n5109), .ZN(n4771) );
  NAND2_X1 U6295 ( .A1(n5568), .A2(n4775), .ZN(n4774) );
  NAND3_X1 U6296 ( .A1(n4598), .A2(n4597), .A3(n5089), .ZN(n5088) );
  NAND2_X1 U6297 ( .A1(n9470), .A2(n4923), .ZN(n4920) );
  NAND2_X1 U6298 ( .A1(n4729), .A2(n5493), .ZN(n7997) );
  OAI21_X4 U6299 ( .B1(n5707), .B2(n5706), .A(n5705), .ZN(n5727) );
  INV_X1 U6300 ( .A(n8125), .ZN(n4572) );
  AND2_X2 U6301 ( .A1(n9811), .A2(n4479), .ZN(n8390) );
  NAND2_X1 U6302 ( .A1(n5144), .A2(n4526), .ZN(n4525) );
  OAI22_X1 U6303 ( .A1(n7206), .A2(n4413), .B1(n4417), .B2(n7207), .ZN(n4606)
         );
  NAND2_X1 U6304 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  NAND2_X1 U6305 ( .A1(n8832), .A2(n6295), .ZN(n8771) );
  NAND2_X1 U6306 ( .A1(n7396), .A2(n7395), .ZN(n6059) );
  NAND2_X1 U6307 ( .A1(n5120), .A2(n6633), .ZN(n7396) );
  NAND2_X1 U6308 ( .A1(n4875), .A2(n4874), .ZN(n4873) );
  OR2_X2 U6309 ( .A1(n6197), .A2(n8056), .ZN(n8079) );
  NAND2_X1 U6310 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  NOR2_X1 U6311 ( .A1(n7276), .A2(n7238), .ZN(n7415) );
  NOR2_X1 U6312 ( .A1(n7557), .A2(n7558), .ZN(n7681) );
  AOI21_X2 U6313 ( .B1(n8778), .B2(n8779), .A(n5106), .ZN(n8373) );
  NAND2_X1 U6314 ( .A1(n4957), .A2(n4953), .ZN(n8856) );
  NAND2_X1 U6315 ( .A1(n4863), .A2(n5687), .ZN(n4862) );
  NOR2_X1 U6316 ( .A1(n9713), .A2(n9712), .ZN(n9721) );
  AOI21_X1 U6317 ( .B1(n9636), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9632), .ZN(
        n7498) );
  NOR2_X2 U6318 ( .A1(n5974), .A2(n5963), .ZN(n6001) );
  NAND2_X1 U6319 ( .A1(n4530), .A2(n4537), .ZN(n7013) );
  INV_X1 U6320 ( .A(n7012), .ZN(n4530) );
  NAND2_X1 U6321 ( .A1(n8882), .A2(n7011), .ZN(n7012) );
  NAND2_X1 U6322 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4534) );
  NAND3_X1 U6323 ( .A1(n4536), .A2(n9592), .A3(n5931), .ZN(n9604) );
  NAND2_X1 U6324 ( .A1(n7014), .A2(n7286), .ZN(n7290) );
  NAND2_X1 U6325 ( .A1(n4554), .A2(n7097), .ZN(n7092) );
  AOI21_X1 U6326 ( .B1(n7123), .B2(n7132), .A(n4515), .ZN(n4900) );
  NAND2_X1 U6327 ( .A1(n9980), .A2(n4511), .ZN(P1_U3549) );
  NAND2_X1 U6328 ( .A1(n10068), .A2(n4505), .ZN(P1_U3517) );
  NAND2_X4 U6329 ( .A1(n5838), .A2(n5837), .ZN(n9812) );
  NAND2_X1 U6330 ( .A1(n6040), .A2(n7007), .ZN(n7186) );
  XNOR2_X2 U6331 ( .A(n5857), .B(n5856), .ZN(n8269) );
  NAND2_X1 U6332 ( .A1(n5655), .A2(n5654), .ZN(n4976) );
  NAND2_X1 U6333 ( .A1(n4766), .A2(n4771), .ZN(n5652) );
  NAND2_X1 U6334 ( .A1(n4646), .A2(n4647), .ZN(n4644) );
  NAND2_X1 U6335 ( .A1(n5005), .A2(n4646), .ZN(n4645) );
  OAI21_X1 U6336 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9977) );
  NOR2_X2 U6337 ( .A1(n8549), .A2(n6485), .ZN(n8463) );
  NOR2_X1 U6338 ( .A1(n8959), .A2(n8980), .ZN(n8971) );
  OAI21_X1 U6339 ( .B1(n4817), .B2(n4433), .A(n4816), .ZN(n8912) );
  NAND2_X1 U6340 ( .A1(n4629), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U6341 ( .A1(n6517), .A2(n6516), .ZN(n10110) );
  NAND2_X1 U6342 ( .A1(n5193), .A2(n5192), .ZN(n6054) );
  NAND2_X1 U6343 ( .A1(n4693), .A2(n4694), .ZN(n4690) );
  NAND2_X1 U6344 ( .A1(n4698), .A2(n6653), .ZN(n4696) );
  NAND2_X1 U6345 ( .A1(n6849), .A2(n5043), .ZN(n5042) );
  OAI21_X2 U6346 ( .B1(n4575), .B2(n4574), .A(n6871), .ZN(n6874) );
  NAND2_X1 U6347 ( .A1(n6853), .A2(n6852), .ZN(n6870) );
  NAND2_X1 U6348 ( .A1(n4749), .A2(n4748), .ZN(n6825) );
  NAND2_X1 U6349 ( .A1(n6812), .A2(n6813), .ZN(n6819) );
  NAND2_X1 U6350 ( .A1(n4751), .A2(n6820), .ZN(n4750) );
  OAI21_X1 U6351 ( .B1(n6837), .B2(n4756), .A(n4755), .ZN(n6842) );
  NAND2_X1 U6352 ( .A1(n6755), .A2(n4801), .ZN(n4800) );
  OAI211_X1 U6353 ( .C1(n6756), .C2(n6984), .A(n4800), .B(n4799), .ZN(n4798)
         );
  NAND2_X1 U6354 ( .A1(n4540), .A2(n8655), .ZN(n9775) );
  NAND3_X1 U6355 ( .A1(n4645), .A2(n4644), .A3(n5006), .ZN(n4540) );
  OR3_X1 U6356 ( .A1(n8583), .A2(n9933), .A3(n8550), .ZN(n8552) );
  NOR2_X1 U6357 ( .A1(n8552), .A2(n8622), .ZN(n8554) );
  NAND3_X1 U6358 ( .A1(n8546), .A2(n8547), .A3(n9968), .ZN(n8548) );
  NAND2_X1 U6359 ( .A1(n5802), .A2(n5801), .ZN(n5830) );
  NAND2_X1 U6360 ( .A1(n4981), .A2(n4978), .ZN(n5800) );
  OR3_X2 U6361 ( .A1(n8537), .A2(n8536), .A3(n8535), .ZN(n8541) );
  NAND4_X1 U6362 ( .A1(n8557), .A2(n9809), .A3(n6497), .A4(n9837), .ZN(n8558)
         );
  NAND2_X1 U6363 ( .A1(n4865), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U6364 ( .A1(n9678), .A2(n9677), .ZN(n4883) );
  NOR2_X1 U6365 ( .A1(n5217), .A2(n4879), .ZN(n4878) );
  OAI211_X1 U6366 ( .C1(n9748), .C2(n5687), .A(n4866), .B(n4862), .ZN(P1_U3262) );
  AOI22_X2 U6367 ( .A1(n4805), .A2(n4804), .B1(n4802), .B2(n4803), .ZN(n9150)
         );
  NAND2_X1 U6368 ( .A1(n5036), .A2(n10202), .ZN(n5037) );
  XNOR2_X2 U6369 ( .A(n5600), .B(n5599), .ZN(n7391) );
  INV_X1 U6370 ( .A(n4770), .ZN(n5628) );
  AOI21_X1 U6371 ( .B1(n4481), .B2(n9081), .A(n4777), .ZN(n9049) );
  OAI22_X1 U6372 ( .A1(n9038), .A2(n6925), .B1(n9352), .B2(n9051), .ZN(n6926)
         );
  NAND2_X1 U6373 ( .A1(n7743), .A2(n7749), .ZN(n5035) );
  NAND2_X1 U6374 ( .A1(n5027), .A2(n5031), .ZN(n5024) );
  NAND2_X1 U6375 ( .A1(n5030), .A2(n5029), .ZN(n5028) );
  OAI21_X2 U6376 ( .B1(n7619), .B2(n6892), .A(n6893), .ZN(n7708) );
  INV_X2 U6377 ( .A(n4731), .ZN(n5382) );
  NAND2_X1 U6378 ( .A1(n8754), .A2(n4561), .ZN(n4560) );
  INV_X1 U6379 ( .A(n4678), .ZN(n4672) );
  NAND2_X1 U6380 ( .A1(n6801), .A2(n4496), .ZN(n6807) );
  NAND2_X2 U6381 ( .A1(n7301), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7368) );
  INV_X1 U6382 ( .A(n7091), .ZN(n4554) );
  NAND2_X1 U6383 ( .A1(n4607), .A2(n5365), .ZN(n5399) );
  NAND2_X1 U6384 ( .A1(n5361), .A2(n5360), .ZN(n5415) );
  NAND2_X1 U6385 ( .A1(n4910), .A2(n4909), .ZN(n9534) );
  NAND2_X1 U6386 ( .A1(n4929), .A2(n5855), .ZN(n9591) );
  NAND2_X1 U6387 ( .A1(n5126), .A2(n4548), .ZN(n4729) );
  NAND2_X1 U6388 ( .A1(n7899), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U6389 ( .A1(n9458), .A2(n9461), .ZN(n9519) );
  NOR2_X1 U6390 ( .A1(n9768), .A2(n4579), .ZN(n6979) );
  NAND2_X1 U6391 ( .A1(n7540), .A2(n7912), .ZN(n6020) );
  AND2_X1 U6392 ( .A1(n4935), .A2(n4550), .ZN(n4934) );
  NAND2_X1 U6393 ( .A1(n4406), .A2(n5627), .ZN(n4772) );
  NAND2_X1 U6394 ( .A1(n8208), .A2(n4565), .ZN(n6236) );
  NAND2_X1 U6395 ( .A1(n5038), .A2(n6891), .ZN(n7619) );
  NAND2_X1 U6396 ( .A1(n6423), .A2(n5057), .ZN(n4806) );
  NAND2_X1 U6397 ( .A1(n8900), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8923) );
  AOI21_X1 U6398 ( .B1(n8945), .B2(n8980), .A(n8965), .ZN(n8946) );
  NAND2_X1 U6399 ( .A1(n8946), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8967) );
  NAND3_X1 U6400 ( .A1(n4622), .A2(n4626), .A3(n4555), .ZN(n8527) );
  OAI21_X1 U6401 ( .B1(n7193), .B2(n4559), .A(n4558), .ZN(n5592) );
  INV_X1 U6402 ( .A(n4972), .ZN(n6513) );
  OAI211_X2 U6403 ( .C1(n5587), .C2(n4913), .A(n4911), .B(n8337), .ZN(n9494)
         );
  NAND2_X2 U6404 ( .A1(n5591), .A2(n5590), .ZN(n8337) );
  NOR2_X2 U6405 ( .A1(n6023), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U6406 ( .A1(n6001), .A2(n5056), .ZN(n6023) );
  OAI211_X1 U6407 ( .C1(n8754), .C2(n8753), .A(n4560), .B(n8752), .ZN(P1_U3220) );
  INV_X1 U6408 ( .A(n9531), .ZN(n4909) );
  NAND3_X1 U6409 ( .A1(n5037), .A2(n4442), .A3(n4420), .ZN(n6945) );
  NAND2_X1 U6410 ( .A1(n7545), .A2(n6890), .ZN(n5038) );
  OAI22_X1 U6411 ( .A1(n5382), .A2(n7768), .B1(n6475), .B2(n5900), .ZN(n5285)
         );
  NAND2_X1 U6412 ( .A1(n4893), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4892) );
  AND2_X2 U6413 ( .A1(n4563), .A2(n7366), .ZN(n7301) );
  NAND2_X1 U6414 ( .A1(n7290), .A2(n4901), .ZN(n4563) );
  NAND2_X1 U6415 ( .A1(n7312), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U6416 ( .A1(n4888), .A2(n7093), .ZN(n7119) );
  NAND2_X1 U6417 ( .A1(n4899), .A2(n4900), .ZN(n8897) );
  OR2_X1 U6418 ( .A1(n7007), .A2(n7025), .ZN(n7010) );
  NAND2_X1 U6419 ( .A1(n4890), .A2(n7021), .ZN(n7090) );
  INV_X1 U6420 ( .A(n7020), .ZN(n4889) );
  NAND2_X1 U6421 ( .A1(n7857), .A2(n7094), .ZN(n4888) );
  NAND2_X1 U6422 ( .A1(n4932), .A2(n4931), .ZN(n6197) );
  NAND4_X1 U6423 ( .A1(n4687), .A2(n4686), .A3(n4437), .A4(n4688), .ZN(n4930)
         );
  OAI21_X1 U6424 ( .B1(n8970), .B2(n8999), .A(n8886), .ZN(n4566) );
  NAND2_X1 U6425 ( .A1(n8371), .A2(n6344), .ZN(n8811) );
  OAI21_X1 U6426 ( .B1(n7757), .B2(n4937), .A(n4934), .ZN(n8080) );
  INV_X1 U6427 ( .A(n6145), .ZN(n4936) );
  AND2_X1 U6428 ( .A1(n6001), .A2(n6000), .ZN(n6005) );
  NAND2_X1 U6429 ( .A1(n5662), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6430 ( .A1(n4586), .A2(n4585), .ZN(n6967) );
  NOR2_X2 U6431 ( .A1(n5548), .A2(n7667), .ZN(n5576) );
  NAND2_X1 U6432 ( .A1(n9969), .A2(n4998), .ZN(n4997) );
  NOR2_X4 U6433 ( .A1(n9821), .A2(n9812), .ZN(n9811) );
  NAND3_X1 U6434 ( .A1(n4484), .A2(n4821), .A3(n8996), .ZN(P2_U3200) );
  INV_X1 U6435 ( .A(n6865), .ZN(n4575) );
  NAND2_X1 U6436 ( .A1(n4798), .A2(n6773), .ZN(n6782) );
  XNOR2_X1 U6437 ( .A(n4576), .B(n9017), .ZN(n6718) );
  NAND2_X1 U6438 ( .A1(n6716), .A2(n6717), .ZN(n4576) );
  NOR4_X2 U6439 ( .A1(n7749), .A2(n7706), .A3(n6702), .A4(n7618), .ZN(n6703)
         );
  NAND2_X1 U6440 ( .A1(n6690), .A2(n6712), .ZN(n6714) );
  NAND3_X1 U6441 ( .A1(n4418), .A2(n9037), .A3(n4578), .ZN(n4577) );
  NAND2_X1 U6442 ( .A1(n7810), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U6443 ( .A1(n7657), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U6444 ( .A1(n4590), .A2(n4483), .ZN(n6558) );
  NAND2_X1 U6445 ( .A1(n8158), .A2(n4593), .ZN(n4590) );
  INV_X1 U6446 ( .A(n4604), .ZN(n4603) );
  INV_X1 U6447 ( .A(n7640), .ZN(n7788) );
  NAND2_X2 U6448 ( .A1(n4415), .A2(n7168), .ZN(n5781) );
  OAI21_X2 U6449 ( .B1(n5399), .B2(n5398), .A(n5371), .ZN(n5431) );
  NAND2_X1 U6450 ( .A1(n5415), .A2(n5363), .ZN(n4607) );
  AND2_X1 U6451 ( .A1(n8444), .A2(n8436), .ZN(n8441) );
  NAND3_X1 U6452 ( .A1(n5394), .A2(n5397), .A3(n4497), .ZN(n9627) );
  NAND3_X1 U6453 ( .A1(n4617), .A2(n4613), .A3(n4499), .ZN(n4848) );
  NAND2_X1 U6454 ( .A1(n4629), .A2(n4623), .ZN(n4622) );
  AND2_X1 U6455 ( .A1(n4625), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U6456 ( .A1(n4630), .A2(n8495), .ZN(n8498) );
  NAND2_X1 U6457 ( .A1(n4631), .A2(n8493), .ZN(n4630) );
  NAND2_X1 U6458 ( .A1(n4634), .A2(n4632), .ZN(n4631) );
  INV_X1 U6459 ( .A(n4633), .ZN(n4632) );
  OAI21_X1 U6460 ( .B1(n8474), .B2(n8473), .A(n4444), .ZN(n4633) );
  NAND2_X1 U6461 ( .A1(n8482), .A2(n8481), .ZN(n4634) );
  NAND3_X1 U6462 ( .A1(n4836), .A2(n4843), .A3(n4635), .ZN(n8446) );
  NAND3_X1 U6463 ( .A1(n5143), .A2(n4638), .A3(n4636), .ZN(n4640) );
  XNOR2_X2 U6464 ( .A(n4639), .B(n5183), .ZN(n10112) );
  INV_X1 U6465 ( .A(n7943), .ZN(n6483) );
  NAND2_X1 U6466 ( .A1(n5015), .A2(n4641), .ZN(n7943) );
  NAND3_X1 U6467 ( .A1(n4488), .A2(n8600), .A3(n6476), .ZN(n4641) );
  NAND2_X1 U6468 ( .A1(n9928), .A2(n4654), .ZN(n4653) );
  AOI21_X2 U6469 ( .B1(n8410), .B2(n8620), .A(n4658), .ZN(n4657) );
  NAND2_X1 U6470 ( .A1(n9774), .A2(n4659), .ZN(n4666) );
  NAND2_X1 U6471 ( .A1(n4665), .A2(n8687), .ZN(n4664) );
  INV_X1 U6472 ( .A(n8508), .ZN(n4660) );
  OAI211_X1 U6473 ( .C1(n9774), .C2(n4669), .A(n4666), .B(n4662), .ZN(n6536)
         );
  INV_X1 U6474 ( .A(n4663), .ZN(n4662) );
  OAI21_X1 U6475 ( .B1(n4665), .B2(n4667), .A(n4664), .ZN(n4663) );
  AND2_X2 U6476 ( .A1(n9592), .A2(n4723), .ZN(n8754) );
  NAND2_X2 U6477 ( .A1(n9487), .A2(n9488), .ZN(n4929) );
  NAND2_X2 U6478 ( .A1(n8070), .A2(n8071), .ZN(n8069) );
  INV_X1 U6479 ( .A(n4677), .ZN(n4676) );
  NOR2_X1 U6480 ( .A1(n4677), .A2(n4672), .ZN(n5168) );
  NOR2_X1 U6481 ( .A1(n5161), .A2(n4673), .ZN(n4675) );
  NAND2_X1 U6482 ( .A1(n9470), .A2(n4681), .ZN(n4679) );
  NAND2_X1 U6483 ( .A1(n4679), .A2(n4680), .ZN(n9553) );
  NOR2_X1 U6484 ( .A1(n8030), .A2(n5900), .ZN(n4685) );
  AND2_X1 U6485 ( .A1(n5958), .A2(n5965), .ZN(n4687) );
  NAND3_X1 U6486 ( .A1(n4437), .A2(n5962), .A3(n5965), .ZN(n4689) );
  NAND2_X1 U6487 ( .A1(n9073), .A2(n4693), .ZN(n4691) );
  NAND3_X1 U6488 ( .A1(n4691), .A2(n6656), .A3(n4690), .ZN(n6930) );
  NAND2_X1 U6489 ( .A1(n9233), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U6490 ( .A1(n4705), .A2(n4709), .ZN(n9200) );
  NAND2_X1 U6491 ( .A1(n10221), .A2(n10200), .ZN(n6747) );
  NOR2_X4 U6492 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5184) );
  AND2_X2 U6493 ( .A1(n5293), .A2(n5255), .ZN(n5186) );
  NAND3_X1 U6494 ( .A1(n4715), .A2(n5186), .A3(n5184), .ZN(n5244) );
  NAND3_X1 U6495 ( .A1(n4717), .A2(n4716), .A3(n5931), .ZN(n5953) );
  NAND2_X1 U6496 ( .A1(n4929), .A2(n4718), .ZN(n4716) );
  OAI21_X2 U6497 ( .B1(n9494), .B2(n4727), .A(n4725), .ZN(n5673) );
  INV_X1 U6498 ( .A(n8220), .ZN(n4728) );
  NAND2_X1 U6499 ( .A1(n7996), .A2(n5514), .ZN(n8070) );
  NAND2_X1 U6500 ( .A1(n4731), .A2(n7780), .ZN(n4730) );
  NAND4_X1 U6501 ( .A1(n4420), .A2(n5037), .A3(n6936), .A4(n10257), .ZN(n6962)
         );
  NAND2_X1 U6502 ( .A1(n6029), .A2(n4736), .ZN(n6186) );
  NAND3_X1 U6503 ( .A1(n5043), .A2(n5041), .A3(n6849), .ZN(n4741) );
  NAND3_X1 U6504 ( .A1(n7547), .A2(n6026), .A3(n6027), .ZN(n6123) );
  NAND4_X1 U6505 ( .A1(n7547), .A2(n6026), .A3(n6027), .A4(n4745), .ZN(n6136)
         );
  NAND3_X2 U6506 ( .A1(n10625), .A2(n4746), .A3(n9750), .ZN(n4965) );
  INV_X2 U6507 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U6508 ( .A1(n6838), .A2(n6984), .ZN(n4760) );
  NAND2_X1 U6509 ( .A1(n5497), .A2(n4460), .ZN(n4766) );
  NAND2_X1 U6510 ( .A1(n5497), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U6511 ( .A1(n4782), .A2(n6919), .ZN(n4778) );
  NOR2_X1 U6512 ( .A1(n8790), .A2(n9087), .ZN(n4785) );
  MUX2_X1 U6513 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9457), .S(n6041), .Z(n7344) );
  NAND3_X1 U6514 ( .A1(n6061), .A2(n6062), .A3(n4786), .ZN(n10204) );
  NAND2_X1 U6515 ( .A1(n7573), .A2(n7912), .ZN(n4795) );
  NAND3_X1 U6516 ( .A1(n4796), .A2(n4441), .A3(n4795), .ZN(n4790) );
  NAND2_X1 U6517 ( .A1(n4796), .A2(n4795), .ZN(n6732) );
  NAND2_X1 U6518 ( .A1(n4790), .A2(n4500), .ZN(n4789) );
  OR2_X1 U6519 ( .A1(n7007), .A2(n7026), .ZN(n6989) );
  NAND2_X1 U6520 ( .A1(n4812), .A2(n4810), .ZN(n4808) );
  OAI21_X1 U6521 ( .B1(n7864), .B2(n4812), .A(n4810), .ZN(n7127) );
  NAND2_X1 U6522 ( .A1(n7864), .A2(n4810), .ZN(n4809) );
  NAND3_X1 U6523 ( .A1(n6996), .A2(n7374), .A3(P2_REG1_REG_5__SCAN_IN), .ZN(
        n7300) );
  NAND2_X1 U6524 ( .A1(n4814), .A2(n10254), .ZN(n4813) );
  INV_X1 U6525 ( .A(n7130), .ZN(n4817) );
  NAND2_X1 U6526 ( .A1(n8887), .A2(n6990), .ZN(n4818) );
  NAND3_X1 U6527 ( .A1(n7282), .A2(n4819), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n7330) );
  NAND2_X1 U6528 ( .A1(n8887), .A2(n4478), .ZN(n4819) );
  NOR2_X1 U6529 ( .A1(n4825), .A2(n4824), .ZN(n4823) );
  INV_X1 U6530 ( .A(n8975), .ZN(n4825) );
  OAI21_X1 U6531 ( .B1(n7158), .B2(n4830), .A(n4827), .ZN(n7002) );
  NAND2_X1 U6532 ( .A1(n4837), .A2(n4834), .ZN(n4836) );
  AND2_X1 U6533 ( .A1(n5312), .A2(n4855), .ZN(n6540) );
  NAND3_X1 U6534 ( .A1(n5150), .A2(n5155), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4855) );
  INV_X4 U6535 ( .A(n4852), .ZN(n6621) );
  NAND2_X2 U6536 ( .A1(n10109), .A2(n8755), .ZN(n4852) );
  NAND3_X1 U6537 ( .A1(n4440), .A2(n5143), .A3(n5144), .ZN(n4860) );
  INV_X2 U6538 ( .A(n5246), .ZN(n5143) );
  NAND3_X1 U6539 ( .A1(n7724), .A2(n4861), .A3(n8412), .ZN(n8586) );
  NAND2_X1 U6540 ( .A1(n7723), .A2(n7725), .ZN(n7724) );
  AOI211_X1 U6541 ( .C1(n8498), .C2(n6497), .A(n8499), .B(n8497), .ZN(n8505)
         );
  NAND2_X2 U6542 ( .A1(n6157), .A2(n4885), .ZN(n7169) );
  NAND2_X1 U6543 ( .A1(n6991), .A2(n7281), .ZN(n7285) );
  NAND2_X1 U6544 ( .A1(n6994), .A2(n6993), .ZN(n6996) );
  MUX2_X1 U6545 ( .A(n10190), .B(P1_REG1_REG_1__SCAN_IN), .S(n9636), .Z(n9633)
         );
  XNOR2_X2 U6546 ( .A(n4878), .B(n4877), .ZN(n9636) );
  AOI21_X1 U6547 ( .B1(n7007), .B2(n4457), .A(n4886), .ZN(n4885) );
  NOR2_X1 U6548 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4886) );
  AND2_X1 U6549 ( .A1(n7092), .A2(n7094), .ZN(n7858) );
  NAND2_X1 U6550 ( .A1(n4892), .A2(n7022), .ZN(n4890) );
  INV_X1 U6551 ( .A(n7018), .ZN(n4894) );
  NAND2_X1 U6552 ( .A1(n4894), .A2(n7159), .ZN(n4895) );
  INV_X1 U6553 ( .A(n7121), .ZN(n4898) );
  NAND2_X1 U6554 ( .A1(n4898), .A2(n7123), .ZN(n4899) );
  INV_X1 U6555 ( .A(n5268), .ZN(n7694) );
  AOI21_X2 U6556 ( .B1(n4906), .B2(n9533), .A(n5125), .ZN(n7899) );
  AND2_X1 U6557 ( .A1(n9534), .A2(n4907), .ZN(n4906) );
  NOR2_X1 U6558 ( .A1(n5290), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U6559 ( .A1(n4920), .A2(n4473), .ZN(n5772) );
  NAND2_X1 U6560 ( .A1(n7757), .A2(n4933), .ZN(n4932) );
  INV_X1 U6561 ( .A(n6184), .ZN(n4938) );
  NAND2_X1 U6562 ( .A1(n8373), .A2(n8372), .ZN(n8371) );
  NAND2_X1 U6563 ( .A1(n8771), .A2(n4950), .ZN(n4946) );
  NAND2_X1 U6564 ( .A1(n4946), .A2(n4947), .ZN(n8778) );
  NAND2_X1 U6565 ( .A1(n8313), .A2(n4954), .ZN(n4957) );
  INV_X1 U6566 ( .A(n4957), .ZN(n8275) );
  AND2_X1 U6567 ( .A1(n4962), .A2(n7607), .ZN(n4961) );
  NAND2_X4 U6568 ( .A1(n4965), .A2(n4963), .ZN(n5362) );
  NAND3_X1 U6569 ( .A1(n4964), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6570 ( .A1(n4975), .A2(n5435), .ZN(n5495) );
  NAND2_X1 U6571 ( .A1(n5727), .A2(n4977), .ZN(n4981) );
  NAND2_X1 U6572 ( .A1(n5727), .A2(n4990), .ZN(n4988) );
  NAND3_X1 U6573 ( .A1(n10173), .A2(n7788), .A3(n7448), .ZN(n7817) );
  AND2_X2 U6574 ( .A1(n9887), .A2(n5000), .ZN(n9856) );
  XNOR2_X2 U6575 ( .A(n5003), .B(n5182), .ZN(n5304) );
  NAND2_X2 U6576 ( .A1(n9836), .A2(n9837), .ZN(n5005) );
  NAND2_X1 U6577 ( .A1(n5008), .A2(n8586), .ZN(n7813) );
  NAND2_X1 U6578 ( .A1(n9962), .A2(n4453), .ZN(n5010) );
  NAND2_X1 U6579 ( .A1(n8463), .A2(n5013), .ZN(n5009) );
  NAND2_X2 U6580 ( .A1(n5010), .A2(n4436), .ZN(n9928) );
  AND2_X1 U6581 ( .A1(n8610), .A2(n5016), .ZN(n5015) );
  NAND3_X1 U6582 ( .A1(n5020), .A2(n5019), .A3(n5021), .ZN(n6448) );
  NAND2_X1 U6583 ( .A1(n8112), .A2(n5027), .ZN(n5025) );
  OAI21_X1 U6584 ( .B1(n4544), .B2(n6903), .A(n6902), .ZN(n8095) );
  NAND2_X1 U6585 ( .A1(n5035), .A2(n4494), .ZN(n6901) );
  XNOR2_X1 U6586 ( .A(n6926), .B(n6929), .ZN(n5036) );
  OR2_X1 U6587 ( .A1(n6657), .A2(n6039), .ZN(n5039) );
  NAND2_X1 U6588 ( .A1(n6073), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6066) );
  XNOR2_X2 U6589 ( .A(n6022), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U6590 ( .B1(n9059), .B2(n6843), .A(n6845), .ZN(n9048) );
  NAND2_X1 U6591 ( .A1(n6843), .A2(n6845), .ZN(n5043) );
  NAND2_X1 U6592 ( .A1(n6651), .A2(n5044), .ZN(n9078) );
  NAND2_X1 U6593 ( .A1(n9078), .A2(n6833), .ZN(n6652) );
  NAND2_X1 U6594 ( .A1(n6644), .A2(n6774), .ZN(n8176) );
  NAND2_X1 U6595 ( .A1(n8176), .A2(n6697), .ZN(n5052) );
  NAND3_X1 U6596 ( .A1(n5965), .A2(n6021), .A3(n6424), .ZN(n5055) );
  NOR2_X1 U6597 ( .A1(n4423), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n5057) );
  INV_X1 U6598 ( .A(n9810), .ZN(n5068) );
  OR2_X1 U6599 ( .A1(n9812), .A2(n9611), .ZN(n5070) );
  NAND2_X1 U6600 ( .A1(n5074), .A2(n8251), .ZN(n5073) );
  AOI21_X1 U6601 ( .B1(n7946), .B2(n5084), .A(n4480), .ZN(n5083) );
  NAND3_X1 U6602 ( .A1(n5087), .A2(n5091), .A3(n5093), .ZN(n5086) );
  AOI211_X1 U6603 ( .C1(n9979), .C2(n10055), .A(n9978), .B(n9977), .ZN(n10066)
         );
  NAND2_X1 U6604 ( .A1(n9856), .A2(n10078), .ZN(n9841) );
  OAI21_X1 U6605 ( .B1(n10173), .B2(n5382), .A(n5313), .ZN(n5314) );
  OAI21_X1 U6606 ( .B1(n4407), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5202), .ZN(
        n5208) );
  INV_X1 U6607 ( .A(n5362), .ZN(n5193) );
  NAND2_X1 U6608 ( .A1(n5362), .A2(n7207), .ZN(n5191) );
  AND2_X1 U6609 ( .A1(n6608), .A2(n8390), .ZN(n6619) );
  NAND2_X1 U6610 ( .A1(n9951), .A2(n8526), .ZN(n10160) );
  NAND2_X1 U6611 ( .A1(n5224), .A2(n8526), .ZN(n6578) );
  INV_X1 U6612 ( .A(n5304), .ZN(n7241) );
  AND2_X2 U6613 ( .A1(n9443), .A2(n9446), .ZN(n6091) );
  AOI21_X1 U6614 ( .B1(n8696), .B2(n10163), .A(n8695), .ZN(n8697) );
  AND2_X1 U6615 ( .A1(n9179), .A2(n9178), .ZN(n9409) );
  OAI21_X1 U6616 ( .B1(n6883), .B2(n10187), .A(n6882), .ZN(n6884) );
  INV_X1 U6617 ( .A(n6025), .ZN(n9446) );
  NAND2_X1 U6618 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  NAND2_X1 U6619 ( .A1(n6023), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6024) );
  INV_X1 U6620 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6621 ( .A1(n6125), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6045) );
  INV_X1 U6622 ( .A(n6814), .ZN(n6649) );
  OR2_X1 U6623 ( .A1(n6628), .A2(n7718), .ZN(n10192) );
  INV_X2 U6624 ( .A(n10192), .ZN(n10194) );
  INV_X2 U6625 ( .A(n10187), .ZN(n10189) );
  NAND2_X1 U6626 ( .A1(n5930), .A2(n5929), .ZN(n9589) );
  INV_X1 U6627 ( .A(n9589), .ZN(n5931) );
  AND2_X1 U6628 ( .A1(n5997), .A2(n5996), .ZN(n5103) );
  OR2_X1 U6629 ( .A1(n6981), .A2(n10036), .ZN(n5104) );
  AND2_X1 U6630 ( .A1(n8724), .A2(n8855), .ZN(n5105) );
  AND2_X1 U6631 ( .A1(n6333), .A2(n9136), .ZN(n5106) );
  OR2_X1 U6632 ( .A1(n6981), .A2(n10096), .ZN(n5107) );
  AND2_X1 U6633 ( .A1(n8958), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6634 ( .A1(n6073), .A2(n7547), .ZN(n5111) );
  AND2_X1 U6635 ( .A1(n5213), .A2(n5214), .ZN(n5112) );
  OR2_X1 U6636 ( .A1(n7217), .A2(n9669), .ZN(n5113) );
  INV_X1 U6637 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U6638 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  INV_X1 U6639 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6325) );
  INV_X1 U6640 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5923) );
  OR2_X1 U6641 ( .A1(n7219), .A2(P1_U3086), .ZN(n8570) );
  INV_X1 U6642 ( .A(n9413), .ZN(n6946) );
  NAND2_X1 U6643 ( .A1(n5217), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5115) );
  INV_X1 U6644 ( .A(n9455), .ZN(n8062) );
  AND2_X1 U6645 ( .A1(n5432), .A2(n5376), .ZN(n5116) );
  AND2_X1 U6646 ( .A1(n6953), .A2(n6873), .ZN(n5117) );
  NOR2_X1 U6647 ( .A1(n6907), .A2(n9253), .ZN(n5118) );
  NOR2_X1 U6648 ( .A1(n6226), .A2(n7622), .ZN(n5119) );
  INV_X1 U6649 ( .A(n8685), .ZN(n6575) );
  INV_X1 U6650 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6296) );
  OR2_X1 U6651 ( .A1(n8711), .A2(n7344), .ZN(n5120) );
  AND2_X1 U6652 ( .A1(n9981), .A2(n9610), .ZN(n5121) );
  OR2_X1 U6653 ( .A1(n7217), .A2(n7267), .ZN(n5122) );
  OR2_X1 U6654 ( .A1(n7217), .A2(n7245), .ZN(n5123) );
  AND3_X1 U6655 ( .A1(n5413), .A2(n5412), .A3(n5411), .ZN(n5124) );
  AND4_X1 U6656 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6469)
         );
  NAND2_X1 U6657 ( .A1(n5347), .A2(n9574), .ZN(n5125) );
  INV_X1 U6658 ( .A(n6976), .ZN(n9781) );
  AND3_X1 U6659 ( .A1(n5486), .A2(n8297), .A3(n5487), .ZN(n5126) );
  OR2_X1 U6660 ( .A1(n6603), .A2(SI_29_), .ZN(n5127) );
  INV_X1 U6661 ( .A(n6964), .ZN(n8707) );
  OR2_X1 U6662 ( .A1(n8013), .A2(n8872), .ZN(n5128) );
  NAND2_X2 U6663 ( .A1(n7542), .A2(n9240), .ZN(n10212) );
  INV_X1 U6664 ( .A(n10257), .ZN(n9273) );
  INV_X2 U6665 ( .A(n10247), .ZN(n10245) );
  AND2_X1 U6666 ( .A1(n6943), .A2(n6942), .ZN(n10247) );
  INV_X1 U6667 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5129) );
  NOR2_X1 U6668 ( .A1(n8664), .A2(n8559), .ZN(n8515) );
  AND3_X1 U6669 ( .A1(n6000), .A2(n6004), .A3(n5964), .ZN(n5965) );
  AOI21_X1 U6670 ( .B1(n9760), .B2(n8518), .A(n8515), .ZN(n8516) );
  NAND2_X1 U6671 ( .A1(n5362), .A2(n7212), .ZN(n5202) );
  OAI21_X1 U6672 ( .B1(n8842), .B2(n9069), .A(n8840), .ZN(n6388) );
  INV_X1 U6673 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10380) );
  INV_X1 U6674 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10383) );
  AND2_X1 U6675 ( .A1(n6748), .A2(n7616), .ZN(n7701) );
  INV_X1 U6676 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5977) );
  INV_X1 U6677 ( .A(n8328), .ZN(n5558) );
  INV_X1 U6678 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5691) );
  INV_X1 U6679 ( .A(SI_26_), .ZN(n5860) );
  INV_X1 U6680 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5214) );
  INV_X1 U6681 ( .A(SI_17_), .ZN(n5629) );
  INV_X1 U6682 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10416) );
  INV_X1 U6683 ( .A(n7485), .ZN(n6080) );
  OR2_X1 U6684 ( .A1(n6282), .A2(n9163), .ZN(n6283) );
  INV_X1 U6685 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6275) );
  INV_X1 U6686 ( .A(n7540), .ZN(n6454) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U6688 ( .A1(n10227), .A2(n8876), .ZN(n7703) );
  OR2_X1 U6689 ( .A1(n6458), .A2(n6984), .ZN(n7522) );
  INV_X1 U6690 ( .A(n9590), .ZN(n5878) );
  INV_X1 U6691 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5731) );
  INV_X1 U6692 ( .A(n9628), .ZN(n7960) );
  AND2_X1 U6693 ( .A1(n8671), .A2(n7492), .ZN(n9595) );
  INV_X1 U6694 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5147) );
  AND2_X1 U6695 ( .A1(n5182), .A2(n5180), .ZN(n5146) );
  NAND2_X1 U6696 ( .A1(n6237), .A2(n9225), .ZN(n6238) );
  INV_X1 U6697 ( .A(n9062), .ZN(n8723) );
  NAND2_X1 U6698 ( .A1(n6268), .A2(n6269), .ZN(n6270) );
  INV_X1 U6699 ( .A(n6181), .ZN(n8050) );
  INV_X1 U6700 ( .A(n9225), .ZN(n9260) );
  OR2_X1 U6701 ( .A1(n9147), .A2(n9146), .ZN(n9172) );
  INV_X1 U6702 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6960) );
  AND2_X1 U6703 ( .A1(n6453), .A2(n7188), .ZN(n6950) );
  INV_X1 U6704 ( .A(n9226), .ZN(n6804) );
  AND2_X1 U6705 ( .A1(n6762), .A2(n6766), .ZN(n7873) );
  INV_X1 U6706 ( .A(n7624), .ZN(n10227) );
  INV_X1 U6707 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6004) );
  AND2_X1 U6708 ( .A1(n5419), .A2(n5122), .ZN(n5420) );
  AND2_X1 U6709 ( .A1(n5230), .A2(n5229), .ZN(n9504) );
  INV_X1 U6710 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9598) );
  INV_X1 U6711 ( .A(n8549), .ZN(n8252) );
  AND2_X1 U6712 ( .A1(n8671), .A2(n10112), .ZN(n9567) );
  AND2_X1 U6713 ( .A1(n8458), .A2(n8612), .ZN(n8547) );
  INV_X1 U6714 ( .A(n9992), .ZN(n9949) );
  AND2_X1 U6715 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5218) );
  OAI21_X1 U6716 ( .B1(n5362), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5191), .ZN(
        n5200) );
  OAI21_X1 U6717 ( .B1(n6924), .B2(n8866), .A(n6465), .ZN(n6466) );
  NAND2_X1 U6718 ( .A1(n6941), .A2(n6451), .ZN(n8861) );
  INV_X1 U6719 ( .A(n8872), .ZN(n8007) );
  INV_X1 U6720 ( .A(n8861), .ZN(n8845) );
  OR2_X1 U6721 ( .A1(n6444), .A2(n7025), .ZN(n6051) );
  OR2_X1 U6722 ( .A1(P2_U3150), .A2(n7071), .ZN(n9020) );
  INV_X1 U6723 ( .A(n9018), .ZN(n8991) );
  AND2_X1 U6724 ( .A1(P2_U3893), .A2(n6449), .ZN(n9023) );
  AND2_X1 U6725 ( .A1(n6933), .A2(n9053), .ZN(n9236) );
  INV_X1 U6726 ( .A(n10240), .ZN(n7891) );
  INV_X1 U6727 ( .A(n9240), .ZN(n10205) );
  INV_X1 U6728 ( .A(n9317), .ZN(n6963) );
  AND2_X1 U6729 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  INV_X1 U6730 ( .A(n9334), .ZN(n10235) );
  OR2_X1 U6731 ( .A1(n8098), .A2(n10235), .ZN(n10238) );
  OR2_X1 U6732 ( .A1(n7187), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U6733 ( .A1(n7445), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9599) );
  INV_X1 U6734 ( .A(n9599), .ZN(n9538) );
  AND3_X1 U6735 ( .A1(n6533), .A2(n6532), .A3(n6531), .ZN(n8559) );
  INV_X1 U6736 ( .A(n5899), .ZN(n6521) );
  OR2_X1 U6737 ( .A1(n10120), .A2(n7492), .ZN(n9745) );
  INV_X1 U6738 ( .A(n9745), .ZN(n10139) );
  OR2_X1 U6739 ( .A1(n8553), .A2(n4446), .ZN(n9883) );
  AND2_X1 U6740 ( .A1(n8476), .A2(n8477), .ZN(n9906) );
  INV_X1 U6741 ( .A(n10160), .ZN(n9971) );
  NAND2_X1 U6742 ( .A1(n5911), .A2(n10103), .ZN(n7718) );
  OR2_X1 U6743 ( .A1(n9970), .A2(n8124), .ZN(n10057) );
  AND2_X1 U6744 ( .A1(n5908), .A2(n5910), .ZN(n7195) );
  INV_X8 U6745 ( .A(n7168), .ZN(n7193) );
  INV_X1 U6746 ( .A(n10114), .ZN(n8065) );
  INV_X1 U6747 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10594) );
  INV_X1 U6748 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10281) );
  INV_X1 U6749 ( .A(n7342), .ZN(n6983) );
  OR3_X1 U6750 ( .A1(n6408), .A2(n8271), .A3(n8223), .ZN(n7070) );
  NAND2_X1 U6751 ( .A1(n8729), .A2(n8718), .ZN(n8728) );
  INV_X1 U6752 ( .A(n9170), .ZN(n9309) );
  INV_X1 U6753 ( .A(n8851), .ZN(n8866) );
  INV_X1 U6754 ( .A(n9006), .ZN(n8976) );
  INV_X1 U6755 ( .A(n9023), .ZN(n8150) );
  NAND2_X1 U6756 ( .A1(n7535), .A2(n10203), .ZN(n9204) );
  INV_X1 U6757 ( .A(n10212), .ZN(n9246) );
  NAND2_X1 U6758 ( .A1(n7543), .A2(n10212), .ZN(n9268) );
  NAND2_X1 U6759 ( .A1(n10257), .A2(n10238), .ZN(n9332) );
  NAND2_X1 U6760 ( .A1(n10257), .A2(n9329), .ZN(n9317) );
  AND2_X2 U6761 ( .A1(n7533), .A2(n6959), .ZN(n10257) );
  INV_X1 U6762 ( .A(n8823), .ZN(n9399) );
  NAND2_X1 U6763 ( .A1(n10245), .A2(n10238), .ZN(n9435) );
  NAND2_X1 U6764 ( .A1(n10245), .A2(n9329), .ZN(n9413) );
  INV_X1 U6765 ( .A(n7215), .ZN(n7216) );
  INV_X1 U6766 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7191) );
  INV_X1 U6767 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10523) );
  INV_X1 U6768 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7406) );
  INV_X2 U6769 ( .A(n9453), .ZN(n9449) );
  INV_X1 U6770 ( .A(n4405), .ZN(n9605) );
  INV_X1 U6771 ( .A(n8739), .ZN(n9608) );
  OR2_X1 U6772 ( .A1(n10120), .A2(n7241), .ZN(n10128) );
  INV_X1 U6773 ( .A(n10122), .ZN(n9749) );
  AND2_X1 U6774 ( .A1(n7963), .A2(n8237), .ZN(n8137) );
  INV_X1 U6775 ( .A(n10163), .ZN(n9957) );
  INV_X1 U6776 ( .A(n9917), .ZN(n10092) );
  NAND2_X1 U6777 ( .A1(n10189), .A2(n10181), .ZN(n10096) );
  OR2_X1 U6778 ( .A1(n6628), .A2(n6627), .ZN(n10187) );
  INV_X1 U6779 ( .A(n10169), .ZN(n10168) );
  OR2_X1 U6780 ( .A1(n8567), .A2(n7195), .ZN(n10169) );
  INV_X1 U6781 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8704) );
  INV_X1 U6782 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10405) );
  INV_X1 U6783 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10592) );
  INV_X1 U6784 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7233) );
  INV_X2 U6785 ( .A(n10106), .ZN(n10115) );
  OR4_X1 U6786 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(P2_U3192)
         );
  AND2_X2 U6787 ( .A1(n7219), .A2(n7117), .ZN(P1_U3973) );
  NAND2_X1 U6788 ( .A1(n6602), .A2(n6601), .ZN(P1_U3551) );
  NOR2_X1 U6789 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5132) );
  NOR2_X2 U6790 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5131) );
  NOR2_X2 U6791 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5130) );
  NAND4_X1 U6792 ( .A1(n5132), .A2(n5131), .A3(n5130), .A4(n5129), .ZN(n5160)
         );
  INV_X1 U6793 ( .A(n5160), .ZN(n5134) );
  NOR2_X1 U6794 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5133) );
  NAND2_X1 U6795 ( .A1(n5134), .A2(n5133), .ZN(n5141) );
  NOR2_X1 U6796 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5137) );
  NOR2_X1 U6797 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5136) );
  NOR2_X1 U6798 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5135) );
  AND3_X1 U6799 ( .A1(n5137), .A2(n5136), .A3(n5135), .ZN(n5140) );
  NAND3_X1 U6800 ( .A1(n5213), .A2(n5138), .A3(n4916), .ZN(n5162) );
  INV_X1 U6801 ( .A(n5162), .ZN(n5139) );
  NAND2_X1 U6802 ( .A1(n5140), .A2(n5139), .ZN(n5176) );
  NAND2_X1 U6803 ( .A1(n6621), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5159) );
  AND2_X2 U6804 ( .A1(n8755), .A2(n5150), .ZN(n5936) );
  NAND2_X1 U6805 ( .A1(n5936), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5158) );
  INV_X1 U6806 ( .A(n5270), .ZN(n5151) );
  NAND2_X1 U6807 ( .A1(n5151), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5233) );
  INV_X1 U6808 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6809 ( .A1(n5270), .A2(n5152), .ZN(n5153) );
  AND2_X1 U6810 ( .A1(n5233), .A2(n5153), .ZN(n9506) );
  NAND2_X1 U6811 ( .A1(n5899), .A2(n9506), .ZN(n5157) );
  AND2_X4 U6812 ( .A1(n5155), .A2(n10109), .ZN(n5410) );
  NAND2_X1 U6813 ( .A1(n5410), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6814 ( .A1(n10408), .A2(n5214), .ZN(n5163) );
  NAND2_X1 U6815 ( .A1(n5170), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5164) );
  MUX2_X1 U6816 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5164), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n5167) );
  INV_X1 U6817 ( .A(n5170), .ZN(n5166) );
  INV_X1 U6818 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6819 ( .A1(n5166), .A2(n5165), .ZN(n5222) );
  MUX2_X1 U6820 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5169), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5171) );
  NAND2_X1 U6821 ( .A1(n5181), .A2(n5172), .ZN(n5173) );
  INV_X1 U6822 ( .A(n5181), .ZN(n5178) );
  NAND2_X1 U6823 ( .A1(n5178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5175) );
  XNOR2_X1 U6824 ( .A(n5175), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5906) );
  OAI21_X1 U6825 ( .B1(n5212), .B2(n5176), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5177) );
  NAND2_X2 U6826 ( .A1(n5223), .A2(n4562), .ZN(n5900) );
  INV_X1 U6827 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6828 ( .A1(n5185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5294) );
  INV_X1 U6829 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6830 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6831 ( .A1(n5294), .A2(n5188), .ZN(n5276) );
  NAND2_X1 U6832 ( .A1(n5278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  INV_X1 U6833 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6834 ( .A(n5190), .B(n5189), .ZN(n9661) );
  INV_X1 U6835 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7170) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7207) );
  XNOR2_X1 U6837 ( .A(n5200), .B(SI_2_), .ZN(n5292) );
  AND2_X1 U6838 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5192) );
  AND2_X1 U6839 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6840 ( .A1(n5362), .A2(n5194), .ZN(n5323) );
  NAND2_X1 U6841 ( .A1(n6054), .A2(n5323), .ZN(n5301) );
  INV_X1 U6842 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U6843 ( .A1(n5362), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5195) );
  INV_X1 U6844 ( .A(SI_1_), .ZN(n5300) );
  OAI211_X1 U6845 ( .C1(n4407), .C2(n7185), .A(n5195), .B(n5300), .ZN(n5196)
         );
  NAND2_X1 U6846 ( .A1(n5301), .A2(n5196), .ZN(n5199) );
  INV_X1 U6847 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U6848 ( .A1(n5362), .A2(n7221), .ZN(n5197) );
  OAI211_X1 U6849 ( .C1(n4407), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5197), .B(
        SI_1_), .ZN(n5198) );
  NAND2_X1 U6850 ( .A1(n5199), .A2(n5198), .ZN(n5291) );
  NAND2_X1 U6851 ( .A1(n5292), .A2(n5291), .ZN(n5258) );
  INV_X1 U6852 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6853 ( .A1(n5201), .A2(SI_2_), .ZN(n5257) );
  INV_X1 U6854 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7172) );
  INV_X1 U6855 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7204) );
  MUX2_X1 U6856 ( .A(n7172), .B(n7204), .S(n5362), .Z(n5259) );
  INV_X1 U6857 ( .A(n5259), .ZN(n5203) );
  NAND2_X1 U6858 ( .A1(n5203), .A2(SI_3_), .ZN(n5281) );
  NAND3_X1 U6859 ( .A1(n5258), .A2(n5257), .A3(n5281), .ZN(n5207) );
  INV_X1 U6860 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7174) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7212) );
  NOR2_X1 U6862 ( .A1(n5203), .A2(SI_3_), .ZN(n5204) );
  NOR2_X1 U6863 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  NAND2_X1 U6864 ( .A1(n5207), .A2(n5206), .ZN(n5353) );
  INV_X1 U6865 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6866 ( .A1(n5209), .A2(SI_4_), .ZN(n5349) );
  NAND2_X1 U6867 ( .A1(n5353), .A2(n5349), .ZN(n5240) );
  INV_X1 U6868 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7173) );
  INV_X1 U6869 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7211) );
  MUX2_X1 U6870 ( .A(n7173), .B(n7211), .S(n4407), .Z(n5241) );
  XNOR2_X1 U6871 ( .A(n5241), .B(SI_5_), .ZN(n5239) );
  XNOR2_X1 U6872 ( .A(n5240), .B(n5239), .ZN(n7210) );
  OR2_X1 U6873 ( .A1(n7210), .A2(n6518), .ZN(n5211) );
  OR2_X1 U6874 ( .A1(n5781), .A2(n7211), .ZN(n5210) );
  OAI211_X1 U6875 ( .C1(n7217), .C2(n9661), .A(n5211), .B(n5210), .ZN(n5228)
         );
  INV_X1 U6876 ( .A(n5658), .ZN(n5215) );
  NAND2_X1 U6877 ( .A1(n5215), .A2(n5112), .ZN(n5221) );
  NAND2_X1 U6878 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5216) );
  NAND2_X1 U6879 ( .A1(n5114), .A2(n5115), .ZN(n5220) );
  XNOR2_X2 U6880 ( .A(n5924), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5224) );
  NAND2_X4 U6881 ( .A1(n5225), .A2(n6578), .ZN(n5849) );
  OAI22_X1 U6882 ( .A1(n8417), .A2(n5900), .B1(n8425), .B2(n5382), .ZN(n5226)
         );
  XNOR2_X1 U6883 ( .A(n5226), .B(n8734), .ZN(n9576) );
  BUF_X2 U6884 ( .A(n5227), .Z(n8738) );
  OR2_X1 U6885 ( .A1(n8417), .A2(n8738), .ZN(n5230) );
  NAND2_X1 U6886 ( .A1(n5228), .A2(n8736), .ZN(n5229) );
  NAND2_X1 U6887 ( .A1(n6621), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6888 ( .A1(n5936), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5237) );
  INV_X1 U6889 ( .A(n5233), .ZN(n5231) );
  NAND2_X1 U6890 ( .A1(n5231), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5407) );
  INV_X1 U6891 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6892 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  AND2_X1 U6893 ( .A1(n5407), .A2(n5234), .ZN(n10144) );
  NAND2_X1 U6894 ( .A1(n5899), .A2(n10144), .ZN(n5236) );
  NAND2_X1 U6895 ( .A1(n5410), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6896 ( .A1(n5240), .A2(n5239), .ZN(n5242) );
  INV_X1 U6897 ( .A(n5241), .ZN(n5354) );
  NAND2_X1 U6898 ( .A1(n5354), .A2(SI_5_), .ZN(n5348) );
  NAND2_X1 U6899 ( .A1(n5242), .A2(n5348), .ZN(n5243) );
  MUX2_X1 U6900 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4407), .Z(n5359) );
  XNOR2_X1 U6901 ( .A(n5359), .B(SI_6_), .ZN(n5356) );
  XNOR2_X1 U6902 ( .A(n5243), .B(n5356), .ZN(n7177) );
  NAND2_X1 U6903 ( .A1(n7177), .A2(n6615), .ZN(n5251) );
  INV_X1 U6904 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7209) );
  OR2_X1 U6905 ( .A1(n5781), .A2(n7209), .ZN(n5249) );
  NAND2_X1 U6906 ( .A1(n5244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5245) );
  MUX2_X1 U6907 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5245), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5248) );
  NAND2_X1 U6908 ( .A1(n5248), .A2(n5247), .ZN(n9669) );
  AND2_X1 U6909 ( .A1(n5249), .A2(n5113), .ZN(n5250) );
  OAI22_X1 U6910 ( .A1(n8423), .A2(n5900), .B1(n8419), .B2(n5382), .ZN(n5252)
         );
  XNOR2_X1 U6911 ( .A(n5252), .B(n5849), .ZN(n5343) );
  OR2_X1 U6912 ( .A1(n8423), .A2(n8738), .ZN(n5254) );
  NAND2_X1 U6913 ( .A1(n10145), .A2(n5905), .ZN(n5253) );
  NAND2_X1 U6914 ( .A1(n5254), .A2(n5253), .ZN(n5344) );
  NAND2_X1 U6915 ( .A1(n5343), .A2(n5344), .ZN(n9575) );
  OAI21_X1 U6916 ( .B1(n9576), .B2(n9504), .A(n9575), .ZN(n5290) );
  NAND2_X1 U6917 ( .A1(n5294), .A2(n5293), .ZN(n5296) );
  NAND2_X1 U6918 ( .A1(n5296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  XNOR2_X1 U6919 ( .A(n5256), .B(n5255), .ZN(n9644) );
  NAND2_X1 U6920 ( .A1(n5258), .A2(n5257), .ZN(n5280) );
  XNOR2_X1 U6921 ( .A(n5259), .B(SI_3_), .ZN(n5279) );
  XNOR2_X1 U6922 ( .A(n5280), .B(n5279), .ZN(n7203) );
  OR2_X1 U6923 ( .A1(n6518), .A2(n7203), .ZN(n5261) );
  OR2_X1 U6924 ( .A1(n5781), .A2(n7204), .ZN(n5260) );
  OAI211_X2 U6925 ( .C1(n7217), .C2(n9644), .A(n5261), .B(n5260), .ZN(n10180)
         );
  NAND2_X1 U6926 ( .A1(n5936), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6927 ( .A1(n6621), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5264) );
  INV_X1 U6928 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U6929 ( .A1(n5899), .A2(n7697), .ZN(n5263) );
  NAND2_X1 U6930 ( .A1(n5410), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5262) );
  AND4_X2 U6931 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n7651)
         );
  NAND2_X1 U6932 ( .A1(n10180), .A2(n8736), .ZN(n5266) );
  NAND2_X1 U6933 ( .A1(n5267), .A2(n4426), .ZN(n5341) );
  NAND2_X1 U6934 ( .A1(n5268), .A2(n5341), .ZN(n9530) );
  NAND2_X1 U6935 ( .A1(n6621), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5275) );
  INV_X1 U6936 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6937 ( .A1(n5269), .A2(n7697), .ZN(n5271) );
  AND2_X1 U6938 ( .A1(n5271), .A2(n5270), .ZN(n10155) );
  NAND2_X1 U6939 ( .A1(n5899), .A2(n10155), .ZN(n5274) );
  NAND2_X1 U6940 ( .A1(n5410), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6941 ( .A1(n5936), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6942 ( .A1(n5276), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6943 ( .A1(n5278), .A2(n5277), .ZN(n7250) );
  OR2_X1 U6944 ( .A1(n5781), .A2(n7212), .ZN(n5284) );
  NAND2_X1 U6945 ( .A1(n5280), .A2(n5279), .ZN(n5282) );
  NAND2_X1 U6946 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  XNOR2_X1 U6947 ( .A(n5285), .B(n5849), .ZN(n5289) );
  OR2_X1 U6948 ( .A1(n6475), .A2(n8738), .ZN(n5287) );
  NAND2_X1 U6949 ( .A1(n10156), .A2(n8736), .ZN(n5286) );
  NAND2_X1 U6950 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  XNOR2_X1 U6951 ( .A(n5289), .B(n5288), .ZN(n9531) );
  NAND2_X1 U6952 ( .A1(n5289), .A2(n5288), .ZN(n9501) );
  NAND2_X1 U6953 ( .A1(n6621), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U6954 ( .A1(n5936), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U6955 ( .A1(n5899), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U6956 ( .A1(n5410), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6470) );
  XNOR2_X1 U6957 ( .A(n5291), .B(n5292), .ZN(n7206) );
  OR2_X1 U6958 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  NAND2_X1 U6959 ( .A1(n5296), .A2(n5295), .ZN(n7245) );
  OAI22_X1 U6960 ( .A1(n6469), .A2(n5900), .B1(n4416), .B2(n5382), .ZN(n5297)
         );
  XNOR2_X1 U6961 ( .A(n5297), .B(n8734), .ZN(n5340) );
  OR2_X1 U6962 ( .A1(n6469), .A2(n8738), .ZN(n5299) );
  NAND2_X1 U6963 ( .A1(n7640), .A2(n8736), .ZN(n5298) );
  NAND2_X1 U6964 ( .A1(n5299), .A2(n5298), .ZN(n5338) );
  XNOR2_X1 U6965 ( .A(n5340), .B(n5338), .ZN(n7627) );
  XNOR2_X1 U6966 ( .A(n5301), .B(n5300), .ZN(n5303) );
  MUX2_X1 U6967 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5362), .Z(n5302) );
  XNOR2_X1 U6968 ( .A(n5303), .B(n5302), .ZN(n7222) );
  AND2_X1 U6969 ( .A1(n7222), .A2(n7193), .ZN(n5310) );
  OAI21_X1 U6970 ( .B1(n7193), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7241), .ZN(
        n5309) );
  CLKBUF_X1 U6971 ( .A(n5304), .Z(n7493) );
  NAND3_X1 U6972 ( .A1(n10112), .A2(n9636), .A3(n7493), .ZN(n5308) );
  INV_X1 U6973 ( .A(n10112), .ZN(n7492) );
  NAND2_X1 U6974 ( .A1(n7168), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5305) );
  OAI21_X1 U6975 ( .B1(n7222), .B2(n7168), .A(n5305), .ZN(n5306) );
  NAND2_X1 U6976 ( .A1(n7492), .A2(n5306), .ZN(n5307) );
  OAI211_X2 U6977 ( .C1(n5310), .C2(n5309), .A(n5308), .B(n5307), .ZN(n7733)
         );
  NAND2_X1 U6978 ( .A1(n5936), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6979 ( .A1(n5410), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6980 ( .A1(n6537), .A2(n8736), .ZN(n5313) );
  XNOR2_X1 U6981 ( .A(n5314), .B(n5849), .ZN(n5334) );
  NAND2_X1 U6982 ( .A1(n6537), .A2(n5876), .ZN(n5316) );
  NAND2_X1 U6983 ( .A1(n5905), .A2(n7733), .ZN(n5315) );
  NAND2_X1 U6984 ( .A1(n5316), .A2(n5315), .ZN(n5335) );
  NAND2_X1 U6985 ( .A1(n5334), .A2(n5335), .ZN(n8383) );
  NAND2_X1 U6986 ( .A1(n6621), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6987 ( .A1(n5936), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6988 ( .A1(n5899), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6989 ( .A1(n5410), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6990 ( .A1(n6538), .A2(n8736), .ZN(n5325) );
  INV_X1 U6991 ( .A(SI_0_), .ZN(n6053) );
  INV_X1 U6992 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5322) );
  OAI21_X1 U6993 ( .B1(n7168), .B2(n6053), .A(n5322), .ZN(n5324) );
  AND2_X1 U6994 ( .A1(n5324), .A2(n5323), .ZN(n10116) );
  NAND2_X1 U6995 ( .A1(n5328), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6996 ( .A1(n5331), .A2(n5326), .ZN(n7443) );
  INV_X1 U6997 ( .A(n6538), .ZN(n5327) );
  AOI22_X1 U6998 ( .A1(n7780), .A2(n8736), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5328), .ZN(n5329) );
  NAND2_X1 U6999 ( .A1(n7443), .A2(n7444), .ZN(n5333) );
  NAND2_X1 U7000 ( .A1(n5331), .A2(n8734), .ZN(n5332) );
  INV_X1 U7001 ( .A(n5334), .ZN(n5337) );
  INV_X1 U7002 ( .A(n5335), .ZN(n5336) );
  INV_X1 U7003 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U7004 ( .A1(n5340), .A2(n5339), .ZN(n7695) );
  AND2_X1 U7005 ( .A1(n7695), .A2(n5341), .ZN(n9527) );
  AND2_X1 U7006 ( .A1(n9527), .A2(n4909), .ZN(n5342) );
  NAND3_X1 U7007 ( .A1(n9575), .A2(n9504), .A3(n9576), .ZN(n5347) );
  INV_X1 U7008 ( .A(n5343), .ZN(n5346) );
  INV_X1 U7009 ( .A(n5344), .ZN(n5345) );
  NAND2_X1 U7010 ( .A1(n5346), .A2(n5345), .ZN(n9574) );
  NOR2_X1 U7011 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  NAND2_X1 U7012 ( .A1(n5353), .A2(n5352), .ZN(n5358) );
  NOR2_X1 U7013 ( .A1(n5354), .A2(SI_5_), .ZN(n5355) );
  NOR2_X1 U7014 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U7015 ( .A1(n5358), .A2(n5357), .ZN(n5361) );
  NAND2_X1 U7016 ( .A1(n5359), .A2(SI_6_), .ZN(n5360) );
  MUX2_X1 U7017 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4407), .Z(n5364) );
  XNOR2_X1 U7018 ( .A(n5364), .B(SI_7_), .ZN(n5416) );
  INV_X1 U7019 ( .A(n5416), .ZN(n5363) );
  NAND2_X1 U7020 ( .A1(n5364), .A2(SI_7_), .ZN(n5365) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7184) );
  INV_X1 U7022 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7214) );
  INV_X1 U7023 ( .A(SI_8_), .ZN(n5367) );
  NAND2_X1 U7024 ( .A1(n5368), .A2(n5367), .ZN(n5371) );
  INV_X1 U7025 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U7026 ( .A1(n5369), .A2(SI_8_), .ZN(n5370) );
  NAND2_X1 U7027 ( .A1(n5371), .A2(n5370), .ZN(n5398) );
  INV_X1 U7028 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7200) );
  INV_X1 U7029 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5372) );
  MUX2_X1 U7030 ( .A(n7200), .B(n5372), .S(n7193), .Z(n5374) );
  INV_X1 U7031 ( .A(SI_9_), .ZN(n5373) );
  NAND2_X1 U7032 ( .A1(n5374), .A2(n5373), .ZN(n5432) );
  INV_X1 U7033 ( .A(n5374), .ZN(n5375) );
  NAND2_X1 U7034 ( .A1(n5375), .A2(SI_9_), .ZN(n5376) );
  XNOR2_X1 U7035 ( .A(n5431), .B(n5116), .ZN(n7192) );
  INV_X1 U7036 ( .A(n5781), .ZN(n5377) );
  NAND2_X1 U7037 ( .A1(n5143), .A2(n5417), .ZN(n5440) );
  NAND2_X1 U7038 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5400) );
  INV_X1 U7039 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U7040 ( .A1(n5400), .A2(n5378), .ZN(n5379) );
  NAND2_X1 U7041 ( .A1(n5379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U7042 ( .A(n5380), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7479) );
  AOI22_X1 U7043 ( .A1(n5377), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5688), .B2(
        n7479), .ZN(n5381) );
  INV_X4 U7044 ( .A(n5382), .ZN(n8731) );
  NAND2_X1 U7045 ( .A1(n8367), .A2(n8731), .ZN(n5390) );
  NAND2_X1 U7046 ( .A1(n6621), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5388) );
  OR2_X2 U7047 ( .A1(n5407), .A2(n5406), .ZN(n5409) );
  NAND2_X1 U7048 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .ZN(n5383) );
  INV_X1 U7049 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5385) );
  INV_X1 U7050 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U7051 ( .B1(n5409), .B2(n5385), .A(n5384), .ZN(n5386) );
  AND2_X1 U7052 ( .A1(n5470), .A2(n5386), .ZN(n8349) );
  NAND2_X1 U7053 ( .A1(n5899), .A2(n8349), .ZN(n5387) );
  OR2_X1 U7054 ( .A1(n7959), .A2(n5900), .ZN(n5389) );
  NAND2_X1 U7055 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  NAND2_X1 U7056 ( .A1(n8367), .A2(n5905), .ZN(n5393) );
  OR2_X1 U7057 ( .A1(n7959), .A2(n8738), .ZN(n5392) );
  AND2_X1 U7058 ( .A1(n5393), .A2(n5392), .ZN(n5483) );
  NAND2_X1 U7059 ( .A1(n5482), .A2(n5483), .ZN(n8360) );
  NAND2_X1 U7060 ( .A1(n6620), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U7061 ( .A1(n6621), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5396) );
  XNOR2_X1 U7062 ( .A(n5409), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U7063 ( .A1(n5899), .A2(n8240), .ZN(n5395) );
  NAND2_X1 U7064 ( .A1(n5410), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U7065 ( .A(n5399), .B(n5398), .ZN(n7182) );
  NAND2_X1 U7066 ( .A1(n7182), .A2(n6615), .ZN(n5402) );
  XNOR2_X1 U7067 ( .A(n5400), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U7068 ( .A1(n5377), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5688), .B2(
        n7418), .ZN(n5401) );
  OR2_X1 U7069 ( .A1(n8030), .A2(n8738), .ZN(n5404) );
  NAND2_X1 U7070 ( .A1(n8142), .A2(n8736), .ZN(n5403) );
  NAND2_X1 U7071 ( .A1(n5429), .A2(n8235), .ZN(n5405) );
  AND2_X1 U7072 ( .A1(n8360), .A2(n5405), .ZN(n8196) );
  NAND2_X1 U7073 ( .A1(n6621), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7074 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  AND2_X1 U7075 ( .A1(n5409), .A2(n5408), .ZN(n7977) );
  NAND2_X1 U7076 ( .A1(n5899), .A2(n7977), .ZN(n5412) );
  NAND2_X1 U7077 ( .A1(n5410), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U7078 ( .A(n5415), .B(n5416), .ZN(n7175) );
  NAND2_X1 U7079 ( .A1(n7175), .A2(n6615), .ZN(n5421) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10321) );
  OR2_X1 U7081 ( .A1(n5781), .A2(n10321), .ZN(n5419) );
  NAND2_X1 U7082 ( .A1(n5247), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U7083 ( .A(n5418), .B(n5417), .ZN(n7267) );
  OAI22_X1 U7084 ( .A1(n7960), .A2(n5900), .B1(n6478), .B2(n5382), .ZN(n5422)
         );
  XNOR2_X1 U7085 ( .A(n5422), .B(n8734), .ZN(n5425) );
  OR2_X1 U7086 ( .A1(n7960), .A2(n8738), .ZN(n5424) );
  NAND2_X1 U7087 ( .A1(n7978), .A2(n8736), .ZN(n5423) );
  AND2_X1 U7088 ( .A1(n5424), .A2(n5423), .ZN(n5426) );
  NAND2_X1 U7089 ( .A1(n5425), .A2(n5426), .ZN(n8192) );
  INV_X1 U7090 ( .A(n5425), .ZN(n5428) );
  INV_X1 U7091 ( .A(n5426), .ZN(n5427) );
  AND2_X1 U7092 ( .A1(n5428), .A2(n5427), .ZN(n7897) );
  INV_X1 U7093 ( .A(n8235), .ZN(n5430) );
  AND2_X1 U7094 ( .A1(n8232), .A2(n5430), .ZN(n8194) );
  OAI21_X1 U7095 ( .B1(n7897), .B2(n8194), .A(n8196), .ZN(n5487) );
  INV_X1 U7096 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7225) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7227) );
  MUX2_X1 U7098 ( .A(n7225), .B(n7227), .S(n7193), .Z(n5433) );
  XNOR2_X1 U7099 ( .A(n5433), .B(SI_10_), .ZN(n5464) );
  INV_X1 U7100 ( .A(n5433), .ZN(n5434) );
  NAND2_X1 U7101 ( .A1(n5434), .A2(SI_10_), .ZN(n5435) );
  MUX2_X1 U7102 ( .A(n7231), .B(n7233), .S(n7193), .Z(n5437) );
  INV_X1 U7103 ( .A(SI_11_), .ZN(n5436) );
  NAND2_X1 U7104 ( .A1(n5437), .A2(n5436), .ZN(n5496) );
  INV_X1 U7105 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U7106 ( .A1(n5438), .A2(SI_11_), .ZN(n5439) );
  NAND2_X1 U7107 ( .A1(n5496), .A2(n5439), .ZN(n5494) );
  NAND2_X1 U7108 ( .A1(n7230), .A2(n6615), .ZN(n5449) );
  INV_X1 U7109 ( .A(n5440), .ZN(n5442) );
  NOR2_X1 U7110 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5441) );
  NAND2_X1 U7111 ( .A1(n5442), .A2(n5441), .ZN(n5465) );
  NAND2_X1 U7112 ( .A1(n5444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5443) );
  MUX2_X1 U7113 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5443), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n5447) );
  INV_X1 U7114 ( .A(n5444), .ZN(n5446) );
  INV_X1 U7115 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7116 ( .A1(n5446), .A2(n5445), .ZN(n5521) );
  NAND2_X1 U7117 ( .A1(n5447), .A2(n5521), .ZN(n7554) );
  INV_X1 U7118 ( .A(n7554), .ZN(n7563) );
  AOI22_X1 U7119 ( .A1(n5377), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5688), .B2(
        n7563), .ZN(n5448) );
  NAND2_X1 U7120 ( .A1(n10062), .A2(n8731), .ZN(n5459) );
  NAND2_X1 U7121 ( .A1(n6620), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7122 ( .A1(n6621), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5456) );
  INV_X1 U7123 ( .A(n5470), .ZN(n5450) );
  NAND2_X1 U7124 ( .A1(n5450), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5472) );
  INV_X1 U7125 ( .A(n5472), .ZN(n5451) );
  NAND2_X1 U7126 ( .A1(n5451), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5501) );
  INV_X1 U7127 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7128 ( .A1(n5472), .A2(n5452), .ZN(n5453) );
  AND2_X1 U7129 ( .A1(n5501), .A2(n5453), .ZN(n8171) );
  NAND2_X1 U7130 ( .A1(n5899), .A2(n8171), .ZN(n5455) );
  NAND2_X1 U7131 ( .A1(n5410), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5454) );
  NAND4_X1 U7132 ( .A1(n5457), .A2(n5456), .A3(n5455), .A4(n5454), .ZN(n9625)
         );
  NAND2_X1 U7133 ( .A1(n9625), .A2(n8736), .ZN(n5458) );
  NAND2_X1 U7134 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  XNOR2_X1 U7135 ( .A(n5460), .B(n5849), .ZN(n8299) );
  NAND2_X1 U7136 ( .A1(n10062), .A2(n8736), .ZN(n5462) );
  NAND2_X1 U7137 ( .A1(n9625), .A2(n5876), .ZN(n5461) );
  NAND2_X1 U7138 ( .A1(n5462), .A2(n5461), .ZN(n8298) );
  NAND2_X1 U7139 ( .A1(n8299), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U7140 ( .A1(n7224), .A2(n6615), .ZN(n5468) );
  NAND2_X1 U7141 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5466) );
  XNOR2_X1 U7142 ( .A(n5466), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7422) );
  AOI22_X1 U7143 ( .A1(n5377), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5688), .B2(
        n7422), .ZN(n5467) );
  NAND2_X1 U7144 ( .A1(n8205), .A2(n8736), .ZN(n5478) );
  NAND2_X1 U7145 ( .A1(n6621), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7146 ( .A1(n5410), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5475) );
  INV_X1 U7147 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7148 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  AND2_X1 U7149 ( .A1(n5472), .A2(n5471), .ZN(n8200) );
  NAND2_X1 U7150 ( .A1(n5899), .A2(n8200), .ZN(n5474) );
  NAND2_X1 U7151 ( .A1(n6620), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5473) );
  OR2_X1 U7152 ( .A1(n8160), .A2(n8738), .ZN(n5477) );
  NAND2_X1 U7153 ( .A1(n5478), .A2(n5477), .ZN(n8199) );
  NAND2_X1 U7154 ( .A1(n8205), .A2(n8731), .ZN(n5480) );
  OR2_X1 U7155 ( .A1(n8160), .A2(n5900), .ZN(n5479) );
  NAND2_X1 U7156 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  XNOR2_X1 U7157 ( .A(n5481), .B(n5849), .ZN(n5488) );
  INV_X1 U7158 ( .A(n5482), .ZN(n5485) );
  INV_X1 U7159 ( .A(n5483), .ZN(n5484) );
  AND2_X1 U7160 ( .A1(n5485), .A2(n5484), .ZN(n8359) );
  AOI21_X1 U7161 ( .B1(n8199), .B2(n5488), .A(n8359), .ZN(n5486) );
  INV_X1 U7162 ( .A(n8299), .ZN(n5492) );
  NAND2_X1 U7163 ( .A1(n5489), .A2(n8298), .ZN(n5491) );
  NOR2_X1 U7164 ( .A1(n8298), .A2(n8199), .ZN(n5490) );
  AOI22_X1 U7165 ( .A1(n5492), .A2(n5491), .B1(n5490), .B2(n8301), .ZN(n5493)
         );
  MUX2_X1 U7166 ( .A(n7339), .B(n10607), .S(n7193), .Z(n5516) );
  XNOR2_X1 U7167 ( .A(n5516), .B(SI_12_), .ZN(n5515) );
  NAND2_X1 U7168 ( .A1(n7338), .A2(n6615), .ZN(n5500) );
  NAND2_X1 U7169 ( .A1(n5521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U7170 ( .A(n5498), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7670) );
  AOI22_X1 U7171 ( .A1(n5377), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5688), .B2(
        n7670), .ZN(n5499) );
  NAND2_X1 U7172 ( .A1(n10053), .A2(n8731), .ZN(n5508) );
  NAND2_X1 U7173 ( .A1(n6620), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7174 ( .A1(n6621), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7175 ( .A1(n5501), .A2(n7559), .ZN(n5502) );
  AND2_X1 U7176 ( .A1(n5527), .A2(n5502), .ZN(n9966) );
  NAND2_X1 U7177 ( .A1(n5899), .A2(n9966), .ZN(n5504) );
  NAND2_X1 U7178 ( .A1(n5410), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5503) );
  OR2_X1 U7179 ( .A1(n8161), .A2(n5900), .ZN(n5507) );
  NAND2_X1 U7180 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  XNOR2_X1 U7181 ( .A(n5509), .B(n8734), .ZN(n5512) );
  NOR2_X1 U7182 ( .A1(n8161), .A2(n8738), .ZN(n5510) );
  AOI21_X1 U7183 ( .B1(n10053), .B2(n5905), .A(n5510), .ZN(n5511) );
  NAND2_X1 U7184 ( .A1(n5512), .A2(n5511), .ZN(n5514) );
  OR2_X1 U7185 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  AND2_X1 U7186 ( .A1(n5514), .A2(n5513), .ZN(n7998) );
  INV_X1 U7187 ( .A(n5515), .ZN(n5519) );
  INV_X1 U7188 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U7189 ( .A1(n5517), .A2(SI_12_), .ZN(n5518) );
  MUX2_X1 U7190 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7193), .Z(n5542) );
  XNOR2_X1 U7191 ( .A(n5542), .B(SI_13_), .ZN(n5541) );
  XNOR2_X1 U7192 ( .A(n5541), .B(n5569), .ZN(n7347) );
  NAND2_X1 U7193 ( .A1(n7347), .A2(n6615), .ZN(n5524) );
  OAI21_X1 U7194 ( .B1(n5521), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5522) );
  XNOR2_X1 U7195 ( .A(n5522), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7673) );
  AOI22_X1 U7196 ( .A1(n5377), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5688), .B2(
        n7673), .ZN(n5523) );
  NAND2_X2 U7197 ( .A1(n5524), .A2(n5523), .ZN(n10049) );
  NAND2_X1 U7198 ( .A1(n10049), .A2(n8731), .ZN(n5534) );
  NAND2_X1 U7199 ( .A1(n6620), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7200 ( .A1(n6621), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7201 ( .A1(n5525), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5548) );
  INV_X1 U7202 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7203 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  AND2_X1 U7204 ( .A1(n5548), .A2(n5528), .ZN(n8127) );
  NAND2_X1 U7205 ( .A1(n5899), .A2(n8127), .ZN(n5530) );
  NAND2_X1 U7206 ( .A1(n5410), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5529) );
  NAND4_X1 U7207 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n9623)
         );
  NAND2_X1 U7208 ( .A1(n9623), .A2(n5905), .ZN(n5533) );
  NAND2_X1 U7209 ( .A1(n5534), .A2(n5533), .ZN(n5535) );
  XNOR2_X1 U7210 ( .A(n5535), .B(n5849), .ZN(n5537) );
  AND2_X1 U7211 ( .A1(n9623), .A2(n5876), .ZN(n5536) );
  AOI21_X1 U7212 ( .B1(n10049), .B2(n8736), .A(n5536), .ZN(n5538) );
  XNOR2_X1 U7213 ( .A(n5537), .B(n5538), .ZN(n8071) );
  INV_X1 U7214 ( .A(n5537), .ZN(n5539) );
  NAND2_X1 U7215 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  INV_X1 U7216 ( .A(n5541), .ZN(n5565) );
  NAND2_X1 U7217 ( .A1(n5569), .A2(n5565), .ZN(n5543) );
  NAND2_X1 U7218 ( .A1(n5542), .A2(SI_13_), .ZN(n5567) );
  NAND2_X1 U7219 ( .A1(n5543), .A2(n5567), .ZN(n5544) );
  XNOR2_X1 U7220 ( .A(n5570), .B(SI_14_), .ZN(n5564) );
  NAND2_X1 U7221 ( .A1(n7354), .A2(n6615), .ZN(n5547) );
  NAND2_X1 U7222 ( .A1(n4510), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5545) );
  XNOR2_X1 U7223 ( .A(n5545), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7935) );
  AOI22_X1 U7224 ( .A1(n5377), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5688), .B2(
        n7935), .ZN(n5546) );
  NAND2_X1 U7225 ( .A1(n10042), .A2(n8731), .ZN(n5555) );
  NAND2_X1 U7226 ( .A1(n6621), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7227 ( .A1(n5410), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7228 ( .A1(n5548), .A2(n7667), .ZN(n5549) );
  AND2_X1 U7229 ( .A1(n5577), .A2(n5549), .ZN(n8261) );
  NAND2_X1 U7230 ( .A1(n5899), .A2(n8261), .ZN(n5551) );
  NAND2_X1 U7231 ( .A1(n6620), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5550) );
  NAND4_X1 U7232 ( .A1(n5553), .A2(n5552), .A3(n5551), .A4(n5550), .ZN(n9622)
         );
  NAND2_X1 U7233 ( .A1(n9622), .A2(n5905), .ZN(n5554) );
  NAND2_X1 U7234 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  XNOR2_X1 U7235 ( .A(n5556), .B(n8734), .ZN(n5559) );
  AND2_X1 U7236 ( .A1(n9622), .A2(n5876), .ZN(n5557) );
  AOI21_X1 U7237 ( .B1(n10042), .B2(n5905), .A(n5557), .ZN(n5560) );
  XNOR2_X1 U7238 ( .A(n5559), .B(n5560), .ZN(n8328) );
  INV_X1 U7239 ( .A(n5559), .ZN(n5562) );
  INV_X1 U7240 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7241 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  INV_X1 U7242 ( .A(n5591), .ZN(n5587) );
  INV_X1 U7243 ( .A(n5564), .ZN(n5566) );
  AND2_X1 U7244 ( .A1(n5566), .A2(n5565), .ZN(n5568) );
  NAND2_X1 U7245 ( .A1(n5570), .A2(SI_14_), .ZN(n5594) );
  NAND2_X1 U7246 ( .A1(n5628), .A2(n5594), .ZN(n5572) );
  XNOR2_X1 U7247 ( .A(n5592), .B(SI_15_), .ZN(n5571) );
  NAND2_X1 U7248 ( .A1(n7360), .A2(n6615), .ZN(n5575) );
  XNOR2_X1 U7249 ( .A(n5573), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9692) );
  AOI22_X1 U7250 ( .A1(n5377), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5688), .B2(
        n9692), .ZN(n5574) );
  NAND2_X2 U7251 ( .A1(n5575), .A2(n5574), .ZN(n10039) );
  NAND2_X1 U7252 ( .A1(n10039), .A2(n8731), .ZN(n5584) );
  NAND2_X1 U7253 ( .A1(n6620), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7254 ( .A1(n6621), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5581) );
  INV_X1 U7255 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U7256 ( .A1(n5577), .A2(n8344), .ZN(n5578) );
  AND2_X1 U7257 ( .A1(n5606), .A2(n5578), .ZN(n9947) );
  NAND2_X1 U7258 ( .A1(n5899), .A2(n9947), .ZN(n5580) );
  NAND2_X1 U7259 ( .A1(n5410), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5579) );
  NAND4_X1 U7260 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .ZN(n9621)
         );
  NAND2_X1 U7261 ( .A1(n9621), .A2(n5905), .ZN(n5583) );
  NAND2_X1 U7262 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  XNOR2_X1 U7263 ( .A(n5585), .B(n5849), .ZN(n5590) );
  INV_X1 U7264 ( .A(n5590), .ZN(n5586) );
  NAND2_X1 U7265 ( .A1(n10039), .A2(n5905), .ZN(n5589) );
  NAND2_X1 U7266 ( .A1(n9621), .A2(n5876), .ZN(n5588) );
  NAND2_X1 U7267 ( .A1(n5589), .A2(n5588), .ZN(n8339) );
  INV_X1 U7268 ( .A(n5592), .ZN(n5596) );
  INV_X1 U7269 ( .A(SI_15_), .ZN(n5595) );
  OR2_X1 U7270 ( .A1(n5596), .A2(n5595), .ZN(n5593) );
  AND2_X1 U7271 ( .A1(n5594), .A2(n5593), .ZN(n5621) );
  NAND2_X1 U7272 ( .A1(n5628), .A2(n5621), .ZN(n5597) );
  NAND2_X1 U7273 ( .A1(n5596), .A2(n5595), .ZN(n5624) );
  NAND2_X1 U7274 ( .A1(n5597), .A2(n5624), .ZN(n5600) );
  INV_X1 U7275 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5598) );
  MUX2_X1 U7276 ( .A(n7406), .B(n5598), .S(n4407), .Z(n5620) );
  XNOR2_X1 U7277 ( .A(n5620), .B(SI_16_), .ZN(n5599) );
  NAND2_X1 U7278 ( .A1(n7391), .A2(n6615), .ZN(n5604) );
  NAND2_X1 U7279 ( .A1(n5601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5602) );
  XNOR2_X1 U7280 ( .A(n5602), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U7281 ( .A1(n5377), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5688), .B2(
        n9702), .ZN(n5603) );
  NAND2_X2 U7282 ( .A1(n5604), .A2(n5603), .ZN(n9936) );
  NAND2_X1 U7283 ( .A1(n9936), .A2(n8731), .ZN(n5613) );
  NAND2_X1 U7284 ( .A1(n6620), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7285 ( .A1(n6621), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7286 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  AND2_X1 U7287 ( .A1(n5639), .A2(n5607), .ZN(n9937) );
  NAND2_X1 U7288 ( .A1(n5899), .A2(n9937), .ZN(n5609) );
  NAND2_X1 U7289 ( .A1(n5410), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5608) );
  OR2_X1 U7290 ( .A1(n8341), .A2(n5900), .ZN(n5612) );
  NAND2_X1 U7291 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  XNOR2_X1 U7292 ( .A(n5614), .B(n8734), .ZN(n5617) );
  NOR2_X1 U7293 ( .A1(n8341), .A2(n8738), .ZN(n5615) );
  AOI21_X1 U7294 ( .B1(n9936), .B2(n5905), .A(n5615), .ZN(n5616) );
  NAND2_X1 U7295 ( .A1(n5617), .A2(n5616), .ZN(n5619) );
  OR2_X1 U7296 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  AND2_X1 U7297 ( .A1(n5619), .A2(n5618), .ZN(n9496) );
  INV_X1 U7298 ( .A(n5620), .ZN(n5623) );
  NAND2_X1 U7299 ( .A1(n5623), .A2(SI_16_), .ZN(n5622) );
  AND2_X1 U7300 ( .A1(n5621), .A2(n5622), .ZN(n5627) );
  INV_X1 U7301 ( .A(n5622), .ZN(n5626) );
  AND2_X1 U7302 ( .A1(n5624), .A2(n4487), .ZN(n5625) );
  MUX2_X1 U7303 ( .A(n7409), .B(n10592), .S(n7193), .Z(n5630) );
  NAND2_X1 U7304 ( .A1(n5630), .A2(n5629), .ZN(n5656) );
  INV_X1 U7305 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7306 ( .A1(n5631), .A2(SI_17_), .ZN(n5632) );
  NAND2_X1 U7307 ( .A1(n5656), .A2(n5632), .ZN(n5653) );
  XNOR2_X1 U7308 ( .A(n5652), .B(n5653), .ZN(n7408) );
  NAND2_X1 U7309 ( .A1(n7408), .A2(n6615), .ZN(n5635) );
  XNOR2_X1 U7310 ( .A(n5633), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U7311 ( .A1(n5377), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5688), .B2(
        n9725), .ZN(n5634) );
  NAND2_X1 U7312 ( .A1(n9917), .A2(n8731), .ZN(n5644) );
  INV_X1 U7313 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U7314 ( .A1(n6620), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7315 ( .A1(n6621), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5636) );
  AND2_X1 U7316 ( .A1(n5637), .A2(n5636), .ZN(n5642) );
  INV_X1 U7317 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7318 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  NAND2_X1 U7319 ( .A1(n5664), .A2(n5640), .ZN(n9914) );
  OR2_X1 U7320 ( .A1(n9914), .A2(n6521), .ZN(n5641) );
  OAI211_X1 U7321 ( .C1(n5816), .C2(n9915), .A(n5642), .B(n5641), .ZN(n9619)
         );
  NAND2_X1 U7322 ( .A1(n9619), .A2(n5905), .ZN(n5643) );
  NAND2_X1 U7323 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  XNOR2_X1 U7324 ( .A(n5645), .B(n5849), .ZN(n5648) );
  NAND2_X1 U7325 ( .A1(n9917), .A2(n5905), .ZN(n5647) );
  NAND2_X1 U7326 ( .A1(n9619), .A2(n5876), .ZN(n5646) );
  NAND2_X1 U7327 ( .A1(n5647), .A2(n5646), .ZN(n5649) );
  NAND2_X1 U7328 ( .A1(n5648), .A2(n5649), .ZN(n9512) );
  INV_X1 U7329 ( .A(n5648), .ZN(n5651) );
  INV_X1 U7330 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7331 ( .A1(n5651), .A2(n5650), .ZN(n9514) );
  INV_X1 U7332 ( .A(n5652), .ZN(n5655) );
  INV_X1 U7333 ( .A(n5653), .ZN(n5654) );
  INV_X1 U7334 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5657) );
  MUX2_X1 U7335 ( .A(n7551), .B(n5657), .S(n7193), .Z(n5680) );
  XNOR2_X1 U7336 ( .A(n5680), .B(SI_18_), .ZN(n5679) );
  XNOR2_X1 U7337 ( .A(n5678), .B(n5679), .ZN(n7511) );
  NAND2_X1 U7338 ( .A1(n7511), .A2(n6615), .ZN(n5661) );
  NAND2_X1 U7339 ( .A1(n5658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U7340 ( .A(n5659), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U7341 ( .A1(n5377), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5688), .B2(
        n9739), .ZN(n5660) );
  NAND2_X1 U7342 ( .A1(n10023), .A2(n8731), .ZN(n5669) );
  INV_X1 U7343 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9728) );
  INV_X1 U7344 ( .A(n5664), .ZN(n5662) );
  INV_X1 U7345 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7346 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  NAND2_X1 U7347 ( .A1(n5692), .A2(n5665), .ZN(n9901) );
  OR2_X1 U7348 ( .A1(n9901), .A2(n6521), .ZN(n5667) );
  AOI22_X1 U7349 ( .A1(n6620), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6621), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5666) );
  OAI211_X1 U7350 ( .C1(n5816), .C2(n9728), .A(n5667), .B(n5666), .ZN(n9618)
         );
  NAND2_X1 U7351 ( .A1(n9618), .A2(n5905), .ZN(n5668) );
  NAND2_X1 U7352 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U7353 ( .A(n5670), .B(n8734), .ZN(n5674) );
  NAND2_X1 U7354 ( .A1(n5673), .A2(n5674), .ZN(n9563) );
  NAND2_X1 U7355 ( .A1(n10023), .A2(n5905), .ZN(n5672) );
  NAND2_X1 U7356 ( .A1(n9618), .A2(n5876), .ZN(n5671) );
  NAND2_X1 U7357 ( .A1(n5672), .A2(n5671), .ZN(n9566) );
  NAND2_X1 U7358 ( .A1(n9563), .A2(n9566), .ZN(n5677) );
  INV_X1 U7359 ( .A(n5674), .ZN(n5675) );
  INV_X1 U7360 ( .A(n5680), .ZN(n5681) );
  NAND2_X1 U7361 ( .A1(n5681), .A2(SI_18_), .ZN(n5682) );
  MUX2_X1 U7362 ( .A(n7635), .B(n8370), .S(n7193), .Z(n5684) );
  NAND2_X1 U7363 ( .A1(n5684), .A2(n10379), .ZN(n5705) );
  INV_X1 U7364 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U7365 ( .A1(n5685), .A2(SI_19_), .ZN(n5686) );
  NAND2_X1 U7366 ( .A1(n5705), .A2(n5686), .ZN(n5706) );
  XNOR2_X1 U7367 ( .A(n5707), .B(n5706), .ZN(n7634) );
  NAND2_X1 U7368 ( .A1(n7634), .A2(n6615), .ZN(n5690) );
  AOI22_X1 U7369 ( .A1(n5377), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5687), .B2(
        n5688), .ZN(n5689) );
  NAND2_X1 U7370 ( .A1(n10018), .A2(n8731), .ZN(n5697) );
  INV_X1 U7371 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U7372 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U7373 ( .A1(n5711), .A2(n5693), .ZN(n9473) );
  OR2_X1 U7374 ( .A1(n9473), .A2(n6521), .ZN(n5695) );
  AOI22_X1 U7375 ( .A1(n6620), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6621), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5694) );
  OAI211_X1 U7376 ( .C1(n5816), .C2(n8402), .A(n5695), .B(n5694), .ZN(n9617)
         );
  NAND2_X1 U7377 ( .A1(n9617), .A2(n5905), .ZN(n5696) );
  NAND2_X1 U7378 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  XNOR2_X1 U7379 ( .A(n5698), .B(n5849), .ZN(n5701) );
  NAND2_X1 U7380 ( .A1(n10018), .A2(n5905), .ZN(n5700) );
  NAND2_X1 U7381 ( .A1(n9617), .A2(n5876), .ZN(n5699) );
  NAND2_X1 U7382 ( .A1(n5700), .A2(n5699), .ZN(n5702) );
  AND2_X1 U7383 ( .A1(n5701), .A2(n5702), .ZN(n9468) );
  INV_X1 U7384 ( .A(n5701), .ZN(n5704) );
  INV_X1 U7385 ( .A(n5702), .ZN(n5703) );
  NAND2_X1 U7386 ( .A1(n5704), .A2(n5703), .ZN(n9467) );
  MUX2_X1 U7387 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7193), .Z(n5725) );
  XNOR2_X1 U7388 ( .A(n5725), .B(n10386), .ZN(n5708) );
  XNOR2_X1 U7389 ( .A(n5727), .B(n5708), .ZN(n7822) );
  NAND2_X1 U7390 ( .A1(n7822), .A2(n6615), .ZN(n5710) );
  INV_X1 U7391 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7824) );
  OR2_X1 U7392 ( .A1(n5781), .A2(n7824), .ZN(n5709) );
  NAND2_X1 U7393 ( .A1(n10014), .A2(n8731), .ZN(n5718) );
  NAND2_X1 U7394 ( .A1(n5711), .A2(n9548), .ZN(n5712) );
  NAND2_X1 U7395 ( .A1(n5732), .A2(n5712), .ZN(n9890) );
  INV_X1 U7396 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U7397 ( .A1(n6620), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7398 ( .A1(n5410), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5713) );
  OAI211_X1 U7399 ( .C1(n4852), .C2(n10395), .A(n5714), .B(n5713), .ZN(n5715)
         );
  INV_X1 U7400 ( .A(n5715), .ZN(n5716) );
  OAI21_X1 U7401 ( .B1(n9890), .B2(n6521), .A(n5716), .ZN(n9616) );
  NAND2_X1 U7402 ( .A1(n9616), .A2(n5905), .ZN(n5717) );
  NAND2_X1 U7403 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  XNOR2_X1 U7404 ( .A(n5719), .B(n8734), .ZN(n5721) );
  AND2_X1 U7405 ( .A1(n9616), .A2(n5876), .ZN(n5720) );
  AOI21_X1 U7406 ( .B1(n10014), .B2(n5905), .A(n5720), .ZN(n5722) );
  AND2_X1 U7407 ( .A1(n5721), .A2(n5722), .ZN(n9542) );
  INV_X1 U7408 ( .A(n5721), .ZN(n5724) );
  INV_X1 U7409 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U7410 ( .A1(n5724), .A2(n5723), .ZN(n9543) );
  INV_X1 U7411 ( .A(n5725), .ZN(n5726) );
  MUX2_X1 U7412 ( .A(n7910), .B(n7909), .S(n7193), .Z(n5743) );
  XNOR2_X1 U7413 ( .A(n5743), .B(SI_21_), .ZN(n5728) );
  XNOR2_X1 U7414 ( .A(n5746), .B(n5728), .ZN(n7908) );
  NAND2_X1 U7415 ( .A1(n7908), .A2(n6615), .ZN(n5730) );
  OR2_X1 U7416 ( .A1(n5781), .A2(n7909), .ZN(n5729) );
  NAND2_X1 U7417 ( .A1(n9876), .A2(n8731), .ZN(n5740) );
  NAND2_X1 U7418 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  AND2_X1 U7419 ( .A1(n5753), .A2(n5733), .ZN(n9870) );
  NAND2_X1 U7420 ( .A1(n9870), .A2(n5899), .ZN(n5738) );
  INV_X1 U7421 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U7422 ( .A1(n6620), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7423 ( .A1(n5410), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7424 ( .C1(n4852), .C2(n10537), .A(n5735), .B(n5734), .ZN(n5736)
         );
  INV_X1 U7425 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7426 ( .A1(n5738), .A2(n5737), .ZN(n9615) );
  NAND2_X1 U7427 ( .A1(n9615), .A2(n5905), .ZN(n5739) );
  NAND2_X1 U7428 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  XNOR2_X1 U7429 ( .A(n5741), .B(n8734), .ZN(n9478) );
  AND2_X1 U7430 ( .A1(n9615), .A2(n5876), .ZN(n5742) );
  AOI21_X1 U7431 ( .B1(n9876), .B2(n5905), .A(n5742), .ZN(n5763) );
  NAND2_X1 U7432 ( .A1(n9478), .A2(n5763), .ZN(n5769) );
  NOR2_X1 U7433 ( .A1(n5744), .A2(SI_21_), .ZN(n5745) );
  MUX2_X1 U7434 ( .A(n8025), .B(n10405), .S(n7193), .Z(n5748) );
  NAND2_X1 U7435 ( .A1(n5748), .A2(n5747), .ZN(n5774) );
  INV_X1 U7436 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7437 ( .A1(n5749), .A2(SI_22_), .ZN(n5750) );
  NAND2_X1 U7438 ( .A1(n5774), .A2(n5750), .ZN(n5775) );
  XNOR2_X1 U7439 ( .A(n5776), .B(n5775), .ZN(n8023) );
  NAND2_X1 U7440 ( .A1(n8023), .A2(n6615), .ZN(n5752) );
  OR2_X1 U7441 ( .A1(n5781), .A2(n10405), .ZN(n5751) );
  NAND2_X1 U7442 ( .A1(n9857), .A2(n8731), .ZN(n5761) );
  INV_X1 U7443 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U7444 ( .A1(n5753), .A2(n10505), .ZN(n5754) );
  NAND2_X1 U7445 ( .A1(n5812), .A2(n5754), .ZN(n9859) );
  OR2_X1 U7446 ( .A1(n9859), .A2(n6521), .ZN(n5759) );
  INV_X1 U7447 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U7448 ( .A1(n6621), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7449 ( .A1(n6620), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5755) );
  OAI211_X1 U7450 ( .C1(n9858), .C2(n5816), .A(n5756), .B(n5755), .ZN(n5757)
         );
  INV_X1 U7451 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7452 ( .A1(n9614), .A2(n5905), .ZN(n5760) );
  NAND2_X1 U7453 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  XNOR2_X1 U7454 ( .A(n5762), .B(n8734), .ZN(n5768) );
  INV_X1 U7455 ( .A(n9478), .ZN(n5764) );
  INV_X1 U7456 ( .A(n5763), .ZN(n9477) );
  NAND2_X1 U7457 ( .A1(n5764), .A2(n9477), .ZN(n5767) );
  NAND2_X1 U7458 ( .A1(n9857), .A2(n5905), .ZN(n5766) );
  NAND2_X1 U7459 ( .A1(n9614), .A2(n5876), .ZN(n5765) );
  NAND2_X1 U7460 ( .A1(n5766), .A2(n5765), .ZN(n9556) );
  NAND2_X1 U7461 ( .A1(n9553), .A2(n9556), .ZN(n5773) );
  INV_X1 U7462 ( .A(n5768), .ZN(n5770) );
  AND2_X1 U7463 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  MUX2_X1 U7464 ( .A(n10523), .B(n8068), .S(n7193), .Z(n5778) );
  INV_X1 U7465 ( .A(SI_23_), .ZN(n5777) );
  NAND2_X1 U7466 ( .A1(n5778), .A2(n5777), .ZN(n5801) );
  INV_X1 U7467 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U7468 ( .A1(n5779), .A2(SI_23_), .ZN(n5780) );
  XNOR2_X1 U7469 ( .A(n5800), .B(n5799), .ZN(n8066) );
  NAND2_X1 U7470 ( .A1(n8066), .A2(n6615), .ZN(n5783) );
  OR2_X1 U7471 ( .A1(n5781), .A2(n8068), .ZN(n5782) );
  NAND2_X1 U7472 ( .A1(n9844), .A2(n8731), .ZN(n5791) );
  XNOR2_X1 U7473 ( .A(n5812), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U7474 ( .A1(n9845), .A2(n5899), .ZN(n5789) );
  INV_X1 U7475 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7476 ( .A1(n6620), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7477 ( .A1(n6621), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5784) );
  OAI211_X1 U7478 ( .C1(n5786), .C2(n5816), .A(n5785), .B(n5784), .ZN(n5787)
         );
  INV_X1 U7479 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7480 ( .A1(n5789), .A2(n5788), .ZN(n9613) );
  NAND2_X1 U7481 ( .A1(n9613), .A2(n5905), .ZN(n5790) );
  NAND2_X1 U7482 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  XNOR2_X1 U7483 ( .A(n5792), .B(n5849), .ZN(n5795) );
  NAND2_X1 U7484 ( .A1(n9844), .A2(n5905), .ZN(n5794) );
  NAND2_X1 U7485 ( .A1(n9613), .A2(n5876), .ZN(n5793) );
  NAND2_X1 U7486 ( .A1(n5794), .A2(n5793), .ZN(n5796) );
  INV_X1 U7487 ( .A(n5795), .ZN(n5798) );
  INV_X1 U7488 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U7489 ( .A1(n5798), .A2(n5797), .ZN(n9461) );
  NAND2_X1 U7490 ( .A1(n5800), .A2(n5799), .ZN(n5802) );
  MUX2_X1 U7491 ( .A(n8221), .B(n8219), .S(n7193), .Z(n5804) );
  INV_X1 U7492 ( .A(SI_24_), .ZN(n5803) );
  NAND2_X1 U7493 ( .A1(n5804), .A2(n5803), .ZN(n5831) );
  INV_X1 U7494 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U7495 ( .A1(n5805), .A2(SI_24_), .ZN(n5806) );
  XNOR2_X1 U7496 ( .A(n5830), .B(n5829), .ZN(n8218) );
  NAND2_X1 U7497 ( .A1(n8218), .A2(n6615), .ZN(n5808) );
  OR2_X1 U7498 ( .A1(n5781), .A2(n8219), .ZN(n5807) );
  NAND2_X1 U7499 ( .A1(n9991), .A2(n8731), .ZN(n5822) );
  INV_X1 U7500 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5810) );
  INV_X1 U7501 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5809) );
  OAI21_X1 U7502 ( .B1(n5812), .B2(n5810), .A(n5809), .ZN(n5813) );
  NAND2_X1 U7503 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5811) );
  AND2_X1 U7504 ( .A1(n5813), .A2(n5840), .ZN(n9822) );
  NAND2_X1 U7505 ( .A1(n9822), .A2(n5899), .ZN(n5820) );
  INV_X1 U7506 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7507 ( .A1(n6620), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7508 ( .A1(n6621), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5814) );
  OAI211_X1 U7509 ( .C1(n5817), .C2(n5816), .A(n5815), .B(n5814), .ZN(n5818)
         );
  INV_X1 U7510 ( .A(n5818), .ZN(n5819) );
  NAND2_X1 U7511 ( .A1(n5820), .A2(n5819), .ZN(n9612) );
  NAND2_X1 U7512 ( .A1(n9612), .A2(n5905), .ZN(n5821) );
  NAND2_X1 U7513 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U7514 ( .A(n5823), .B(n5849), .ZN(n5825) );
  AND2_X1 U7515 ( .A1(n9612), .A2(n5876), .ZN(n5824) );
  AOI21_X1 U7516 ( .B1(n9991), .B2(n5905), .A(n5824), .ZN(n5826) );
  XNOR2_X1 U7517 ( .A(n5825), .B(n5826), .ZN(n9521) );
  NAND2_X1 U7518 ( .A1(n9519), .A2(n9521), .ZN(n9520) );
  INV_X1 U7519 ( .A(n5825), .ZN(n5827) );
  NAND2_X1 U7520 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND2_X1 U7521 ( .A1(n5830), .A2(n5829), .ZN(n5832) );
  MUX2_X1 U7522 ( .A(n8270), .B(n8272), .S(n7193), .Z(n5834) );
  INV_X1 U7523 ( .A(SI_25_), .ZN(n5833) );
  NAND2_X1 U7524 ( .A1(n5834), .A2(n5833), .ZN(n5858) );
  INV_X1 U7525 ( .A(n5834), .ZN(n5835) );
  NAND2_X1 U7526 ( .A1(n5835), .A2(SI_25_), .ZN(n5836) );
  NAND2_X1 U7527 ( .A1(n8269), .A2(n6615), .ZN(n5838) );
  OR2_X1 U7528 ( .A1(n5781), .A2(n8272), .ZN(n5837) );
  NAND2_X1 U7529 ( .A1(n9812), .A2(n8731), .ZN(n5848) );
  INV_X1 U7530 ( .A(n5840), .ZN(n5839) );
  NAND2_X1 U7531 ( .A1(n5839), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5866) );
  INV_X1 U7532 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10509) );
  NAND2_X1 U7533 ( .A1(n5840), .A2(n10509), .ZN(n5841) );
  NAND2_X1 U7534 ( .A1(n5866), .A2(n5841), .ZN(n9813) );
  INV_X1 U7535 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U7536 ( .A1(n6620), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7537 ( .A1(n5410), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5842) );
  OAI211_X1 U7538 ( .C1(n4852), .C2(n10406), .A(n5843), .B(n5842), .ZN(n5844)
         );
  INV_X1 U7539 ( .A(n5844), .ZN(n5845) );
  NAND2_X1 U7540 ( .A1(n9611), .A2(n5905), .ZN(n5847) );
  NAND2_X1 U7541 ( .A1(n5848), .A2(n5847), .ZN(n5850) );
  XNOR2_X1 U7542 ( .A(n5850), .B(n5849), .ZN(n5852) );
  AND2_X1 U7543 ( .A1(n9611), .A2(n5876), .ZN(n5851) );
  AOI21_X1 U7544 ( .B1(n9812), .B2(n5905), .A(n5851), .ZN(n5853) );
  XNOR2_X1 U7545 ( .A(n5852), .B(n5853), .ZN(n9488) );
  INV_X1 U7546 ( .A(n5852), .ZN(n5854) );
  NAND2_X1 U7547 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U7548 ( .A1(n5857), .A2(n5856), .ZN(n5859) );
  NAND2_X1 U7549 ( .A1(n5859), .A2(n5858), .ZN(n5885) );
  MUX2_X1 U7550 ( .A(n8333), .B(n8334), .S(n7193), .Z(n5861) );
  NAND2_X1 U7551 ( .A1(n5861), .A2(n5860), .ZN(n5886) );
  INV_X1 U7552 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U7553 ( .A1(n5862), .A2(SI_26_), .ZN(n5863) );
  XNOR2_X1 U7554 ( .A(n5885), .B(n5884), .ZN(n8332) );
  NAND2_X1 U7555 ( .A1(n8332), .A2(n6615), .ZN(n5865) );
  OR2_X1 U7556 ( .A1(n5781), .A2(n8334), .ZN(n5864) );
  NAND2_X1 U7557 ( .A1(n9981), .A2(n8731), .ZN(n5874) );
  NAND2_X1 U7558 ( .A1(n5866), .A2(n9598), .ZN(n5867) );
  NAND2_X1 U7559 ( .A1(n9798), .A2(n5899), .ZN(n5872) );
  INV_X1 U7560 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U7561 ( .A1(n5410), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7562 ( .A1(n6621), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5868) );
  OAI211_X1 U7563 ( .C1(n6524), .C2(n10443), .A(n5869), .B(n5868), .ZN(n5870)
         );
  INV_X1 U7564 ( .A(n5870), .ZN(n5871) );
  NAND2_X1 U7565 ( .A1(n9610), .A2(n5905), .ZN(n5873) );
  NAND2_X1 U7566 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  XNOR2_X1 U7567 ( .A(n5875), .B(n8734), .ZN(n5879) );
  AND2_X1 U7568 ( .A1(n9610), .A2(n5876), .ZN(n5877) );
  AOI21_X1 U7569 ( .B1(n9981), .B2(n5905), .A(n5877), .ZN(n5880) );
  XNOR2_X1 U7570 ( .A(n5879), .B(n5880), .ZN(n9590) );
  INV_X1 U7571 ( .A(n5879), .ZN(n5882) );
  INV_X1 U7572 ( .A(n5880), .ZN(n5881) );
  NAND2_X1 U7573 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  NAND2_X1 U7574 ( .A1(n5885), .A2(n5884), .ZN(n5887) );
  MUX2_X1 U7575 ( .A(n6392), .B(n8704), .S(n7193), .Z(n5889) );
  INV_X1 U7576 ( .A(SI_27_), .ZN(n5888) );
  NAND2_X1 U7577 ( .A1(n5889), .A2(n5888), .ZN(n6502) );
  INV_X1 U7578 ( .A(n5889), .ZN(n5890) );
  NAND2_X1 U7579 ( .A1(n5890), .A2(SI_27_), .ZN(n5891) );
  NAND2_X1 U7580 ( .A1(n8703), .A2(n6615), .ZN(n5893) );
  OR2_X1 U7581 ( .A1(n5781), .A2(n8704), .ZN(n5892) );
  NAND2_X1 U7582 ( .A1(n9782), .A2(n8731), .ZN(n5902) );
  INV_X1 U7583 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7584 ( .A1(n5894), .A2(n5946), .ZN(n5895) );
  INV_X1 U7585 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U7586 ( .A1(n5410), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7587 ( .A1(n6621), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5896) );
  OAI211_X1 U7588 ( .C1(n6524), .C2(n10456), .A(n5897), .B(n5896), .ZN(n5898)
         );
  OR2_X1 U7589 ( .A1(n9594), .A2(n5900), .ZN(n5901) );
  NAND2_X1 U7590 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  XNOR2_X1 U7591 ( .A(n5903), .B(n8734), .ZN(n8743) );
  NOR2_X1 U7592 ( .A1(n9594), .A2(n8738), .ZN(n5904) );
  AOI21_X1 U7593 ( .B1(n9782), .B2(n5905), .A(n5904), .ZN(n8742) );
  INV_X1 U7594 ( .A(n5906), .ZN(n8274) );
  NAND2_X1 U7595 ( .A1(n8274), .A2(P1_B_REG_SCAN_IN), .ZN(n5907) );
  MUX2_X1 U7596 ( .A(P1_B_REG_SCAN_IN), .B(n5907), .S(n8220), .Z(n5908) );
  INV_X1 U7597 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7598 ( .A1(n7195), .A2(n5909), .ZN(n5911) );
  INV_X1 U7599 ( .A(n5910), .ZN(n8336) );
  NAND2_X1 U7600 ( .A1(n8220), .A2(n8336), .ZN(n10103) );
  INV_X1 U7601 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7199) );
  NAND2_X1 U7602 ( .A1(n7195), .A2(n7199), .ZN(n5912) );
  NAND2_X1 U7603 ( .A1(n8336), .A2(n8274), .ZN(n7196) );
  NAND2_X1 U7604 ( .A1(n5912), .A2(n7196), .ZN(n6596) );
  INV_X1 U7605 ( .A(n6596), .ZN(n7719) );
  INV_X1 U7606 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10546) );
  INV_X1 U7607 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10414) );
  INV_X1 U7608 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10470) );
  INV_X1 U7609 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10474) );
  NAND4_X1 U7610 ( .A1(n10546), .A2(n10414), .A3(n10470), .A4(n10474), .ZN(
        n5913) );
  NOR4_X1 U7611 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(n5913), .ZN(n10334) );
  NOR4_X1 U7612 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5914) );
  INV_X1 U7613 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10533) );
  INV_X1 U7614 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10407) );
  NAND3_X1 U7615 ( .A1(n5914), .A2(n10533), .A3(n10407), .ZN(n5920) );
  NOR4_X1 U7616 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5918) );
  NOR4_X1 U7617 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5917) );
  NOR4_X1 U7618 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5916) );
  NOR4_X1 U7619 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U7620 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n5919)
         );
  NOR3_X1 U7621 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n5920), .A3(n5919), .ZN(n5921) );
  NAND2_X1 U7622 ( .A1(n10334), .A2(n5921), .ZN(n5922) );
  NAND2_X1 U7623 ( .A1(n7195), .A2(n5922), .ZN(n6594) );
  NAND3_X1 U7624 ( .A1(n6627), .A2(n7719), .A3(n6594), .ZN(n5942) );
  NAND2_X1 U7625 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  INV_X1 U7626 ( .A(n5950), .ZN(n5930) );
  NOR2_X1 U7627 ( .A1(n10181), .A2(n8671), .ZN(n5929) );
  INV_X1 U7628 ( .A(n5934), .ZN(n5932) );
  NAND2_X1 U7629 ( .A1(n5932), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8690) );
  INV_X1 U7630 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7631 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  NAND2_X1 U7632 ( .A1(n8690), .A2(n5935), .ZN(n9765) );
  INV_X1 U7633 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U7634 ( .A1(n5936), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7635 ( .A1(n5410), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5937) );
  OAI211_X1 U7636 ( .C1(n4852), .C2(n10473), .A(n5938), .B(n5937), .ZN(n5939)
         );
  INV_X1 U7637 ( .A(n5939), .ZN(n5940) );
  OAI22_X1 U7638 ( .A1(n8739), .A2(n9593), .B1(n6499), .B2(n8398), .ZN(n9777)
         );
  NOR2_X2 U7639 ( .A1(n5950), .A2(n8571), .ZN(n9602) );
  INV_X1 U7640 ( .A(n9783), .ZN(n5947) );
  NAND2_X1 U7641 ( .A1(n5942), .A2(n6597), .ZN(n5945) );
  AND2_X1 U7642 ( .A1(n7219), .A2(n4562), .ZN(n5944) );
  NAND2_X1 U7643 ( .A1(n8671), .A2(n8571), .ZN(n5943) );
  NAND2_X1 U7644 ( .A1(n5945), .A2(n6595), .ZN(n7445) );
  OAI22_X1 U7645 ( .A1(n5947), .A2(n9599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5946), .ZN(n5948) );
  AOI21_X1 U7646 ( .B1(n9777), .B2(n9602), .A(n5948), .ZN(n5952) );
  AND2_X1 U7647 ( .A1(n7777), .A2(n8675), .ZN(n7732) );
  INV_X1 U7648 ( .A(n7732), .ZN(n5949) );
  NAND2_X1 U7649 ( .A1(n9782), .A2(n4405), .ZN(n5951) );
  NAND3_X1 U7650 ( .A1(n5953), .A2(n5952), .A3(n5951), .ZN(P1_U3214) );
  NAND2_X1 U7651 ( .A1(n6011), .A2(n6015), .ZN(n5970) );
  NAND2_X1 U7652 ( .A1(n5970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5966) );
  INV_X1 U7653 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U7654 ( .B1(n5967), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U7655 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_27__SCAN_IN), .A(
        n5968), .ZN(n5969) );
  INV_X1 U7656 ( .A(n5970), .ZN(n5972) );
  XNOR2_X2 U7657 ( .A(n5973), .B(n6021), .ZN(n6449) );
  NAND2_X1 U7658 ( .A1(n7354), .A2(n6675), .ZN(n5983) );
  INV_X1 U7659 ( .A(n5974), .ZN(n5976) );
  NAND2_X1 U7660 ( .A1(n5976), .A2(n5975), .ZN(n6201) );
  NAND2_X1 U7661 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  AOI21_X1 U7662 ( .B1(n6220), .B2(n5985), .A(n9439), .ZN(n5979) );
  NAND2_X1 U7663 ( .A1(n5979), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5981) );
  INV_X1 U7664 ( .A(n5979), .ZN(n5980) );
  NAND2_X1 U7665 ( .A1(n5980), .A2(n5984), .ZN(n6241) );
  AOI22_X1 U7666 ( .A1(n6300), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6301), .B2(
        n8910), .ZN(n5982) );
  NAND2_X2 U7667 ( .A1(n5983), .A2(n5982), .ZN(n9423) );
  INV_X1 U7668 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5986) );
  NAND3_X1 U7669 ( .A1(n5986), .A2(n5985), .A3(n5984), .ZN(n5987) );
  NAND2_X1 U7670 ( .A1(n6258), .A2(n5990), .ZN(n6284) );
  AND2_X1 U7671 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5991) );
  NAND2_X1 U7672 ( .A1(n6284), .A2(n5991), .ZN(n5999) );
  INV_X1 U7673 ( .A(n6001), .ZN(n5997) );
  NAND2_X1 U7674 ( .A1(n5997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7675 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n5994) );
  NAND2_X1 U7676 ( .A1(n5994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5995) );
  OAI21_X1 U7677 ( .B1(n5993), .B2(P2_IR_REG_31__SCAN_IN), .A(n5995), .ZN(
        n5996) );
  INV_X1 U7678 ( .A(n6005), .ZN(n6002) );
  NAND2_X1 U7679 ( .A1(n6002), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7680 ( .A1(n6005), .A2(n6004), .ZN(n6427) );
  INV_X1 U7681 ( .A(n6008), .ZN(n6007) );
  NAND2_X1 U7682 ( .A1(n6008), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7683 ( .A1(n6012), .A2(n6011), .ZN(n6014) );
  OR2_X1 U7684 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7685 ( .A1(n6408), .A2(n8223), .ZN(n7189) );
  NAND2_X1 U7686 ( .A1(n4797), .A2(n6953), .ZN(n6927) );
  AND2_X1 U7687 ( .A1(n7189), .A2(n6927), .ZN(n6019) );
  NAND2_X1 U7688 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7689 ( .A(n8223), .B(P2_B_REG_SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7690 ( .A1(n8271), .A2(n6017), .ZN(n6407) );
  AND2_X1 U7691 ( .A1(n6406), .A2(n7191), .ZN(n6018) );
  NAND2_X1 U7692 ( .A1(n6407), .A2(n6018), .ZN(n6411) );
  XNOR2_X1 U7693 ( .A(n9423), .B(n4553), .ZN(n6239) );
  INV_X1 U7694 ( .A(n6239), .ZN(n6240) );
  OR2_X2 U7695 ( .A1(n9438), .A2(n9439), .ZN(n6022) );
  BUF_X4 U7696 ( .A(n6091), .Z(n6682) );
  NAND2_X1 U7697 ( .A1(n6682), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7698 ( .A1(n6122), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6037) );
  INV_X1 U7699 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6026) );
  INV_X1 U7700 ( .A(n6136), .ZN(n6029) );
  NAND2_X1 U7701 ( .A1(n6225), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7702 ( .A1(n6247), .A2(n6033), .ZN(n9230) );
  NAND2_X1 U7703 ( .A1(n6659), .A2(n9230), .ZN(n6036) );
  NAND2_X1 U7704 ( .A1(n6681), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6035) );
  NAND4_X1 U7705 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n9238)
         );
  INV_X1 U7706 ( .A(n9238), .ZN(n9213) );
  INV_X1 U7707 ( .A(n7222), .ZN(n6039) );
  INV_X1 U7708 ( .A(n7186), .ZN(n7320) );
  NAND2_X1 U7709 ( .A1(n6073), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6047) );
  INV_X1 U7710 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7711 ( .A1(n6090), .A2(n6043), .ZN(n6044) );
  NAND2_X1 U7712 ( .A1(n6073), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7713 ( .A1(n6091), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6049) );
  INV_X1 U7714 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7026) );
  OR2_X1 U7715 ( .A1(n6090), .A2(n7026), .ZN(n6048) );
  INV_X1 U7716 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7025) );
  INV_X1 U7717 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U7718 ( .B1(n7193), .B2(n6053), .A(n6052), .ZN(n6055) );
  AND2_X1 U7719 ( .A1(n6054), .A2(n6055), .ZN(n9457) );
  INV_X1 U7720 ( .A(n6056), .ZN(n6057) );
  OR2_X1 U7721 ( .A1(n6057), .A2(n10198), .ZN(n6058) );
  NAND2_X1 U7722 ( .A1(n6059), .A2(n6058), .ZN(n7384) );
  OR2_X1 U7723 ( .A1(n6087), .A2(n7170), .ZN(n6062) );
  OR2_X1 U7724 ( .A1(n6657), .A2(n7206), .ZN(n6061) );
  NAND2_X1 U7725 ( .A1(n6091), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6067) );
  INV_X1 U7726 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10213) );
  INV_X1 U7727 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10248) );
  OR2_X1 U7728 ( .A1(n6090), .A2(n10248), .ZN(n6064) );
  XNOR2_X1 U7729 ( .A(n6068), .B(n7579), .ZN(n7385) );
  NAND2_X1 U7730 ( .A1(n7384), .A2(n7385), .ZN(n6071) );
  INV_X1 U7731 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7732 ( .A1(n7579), .A2(n6069), .ZN(n6070) );
  NAND2_X1 U7733 ( .A1(n6071), .A2(n6070), .ZN(n7484) );
  INV_X1 U7734 ( .A(n7484), .ZN(n6081) );
  INV_X1 U7735 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10467) );
  OR2_X1 U7736 ( .A1(n6072), .A2(n10467), .ZN(n6076) );
  NAND2_X1 U7737 ( .A1(n6091), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6075) );
  INV_X1 U7738 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10250) );
  OR2_X1 U7739 ( .A1(n6090), .A2(n10250), .ZN(n6074) );
  OR2_X1 U7740 ( .A1(n7203), .A2(n6657), .ZN(n6079) );
  OR2_X1 U7741 ( .A1(n6087), .A2(n7172), .ZN(n6078) );
  XNOR2_X1 U7742 ( .A(n7548), .B(n8711), .ZN(n6082) );
  XNOR2_X1 U7743 ( .A(n7387), .B(n6082), .ZN(n7485) );
  NAND2_X1 U7744 ( .A1(n6081), .A2(n6080), .ZN(n7482) );
  INV_X1 U7745 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7746 ( .A1(n10200), .A2(n6083), .ZN(n6084) );
  NOR2_X1 U7747 ( .A1(n6085), .A2(n6657), .ZN(n6089) );
  NAND2_X1 U7748 ( .A1(n6100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7749 ( .A(n7624), .B(n8711), .ZN(n6098) );
  NAND2_X1 U7750 ( .A1(n6681), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6097) );
  INV_X1 U7751 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10252) );
  OR2_X1 U7752 ( .A1(n6090), .A2(n10252), .ZN(n6093) );
  NAND2_X1 U7753 ( .A1(n6091), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7754 ( .A1(n6093), .A2(n6092), .ZN(n6095) );
  NAND2_X1 U7755 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6094) );
  AND2_X1 U7756 ( .A1(n6109), .A2(n6094), .ZN(n7622) );
  NAND2_X2 U7757 ( .A1(n6097), .A2(n6096), .ZN(n8876) );
  XNOR2_X1 U7758 ( .A(n6098), .B(n8876), .ZN(n7515) );
  INV_X1 U7759 ( .A(n8876), .ZN(n7488) );
  NAND2_X1 U7760 ( .A1(n7488), .A2(n6098), .ZN(n6099) );
  OR2_X1 U7761 ( .A1(n7210), .A2(n6657), .ZN(n6107) );
  INV_X1 U7762 ( .A(n6100), .ZN(n6102) );
  NAND2_X1 U7763 ( .A1(n6102), .A2(n6101), .ZN(n6118) );
  NAND2_X1 U7764 ( .A1(n6118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6104) );
  INV_X1 U7765 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7766 ( .A1(n6678), .A2(n7173), .ZN(n6105) );
  XNOR2_X1 U7767 ( .A(n10231), .B(n8711), .ZN(n6116) );
  INV_X1 U7768 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7769 ( .A1(n6444), .A2(n6108), .ZN(n6115) );
  INV_X1 U7770 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U7771 ( .A1(n6109), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6110) );
  AND2_X1 U7772 ( .A1(n6123), .A2(n6110), .ZN(n7714) );
  OR2_X1 U7773 ( .A1(n6226), .A2(n7714), .ZN(n6112) );
  NAND2_X1 U7774 ( .A1(n6682), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6111) );
  NAND2_X2 U7775 ( .A1(n6115), .A2(n6114), .ZN(n8875) );
  XNOR2_X1 U7776 ( .A(n6116), .B(n7517), .ZN(n7607) );
  INV_X1 U7777 ( .A(n6116), .ZN(n6117) );
  NAND2_X1 U7778 ( .A1(n7177), .A2(n6675), .ZN(n6121) );
  NAND2_X1 U7779 ( .A1(n6130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6119) );
  XNOR2_X1 U7780 ( .A(n6119), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7373) );
  AOI22_X1 U7781 ( .A1(n6300), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6301), .B2(
        n7373), .ZN(n6120) );
  XNOR2_X1 U7782 ( .A(n10240), .B(n6063), .ZN(n6142) );
  NAND2_X1 U7783 ( .A1(n6123), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6124) );
  AND2_X1 U7784 ( .A1(n6136), .A2(n6124), .ZN(n7889) );
  OR2_X1 U7785 ( .A1(n6226), .A2(n7889), .ZN(n6128) );
  NAND2_X1 U7786 ( .A1(n6682), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7787 ( .A1(n6681), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6126) );
  XNOR2_X1 U7788 ( .A(n6142), .B(n8874), .ZN(n7758) );
  NAND2_X1 U7789 ( .A1(n7759), .A2(n7758), .ZN(n7757) );
  NAND2_X1 U7790 ( .A1(n7175), .A2(n6675), .ZN(n6134) );
  INV_X1 U7791 ( .A(n6130), .ZN(n6132) );
  INV_X1 U7792 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7793 ( .A1(n6132), .A2(n6131), .ZN(n6148) );
  NAND2_X1 U7794 ( .A1(n6148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U7795 ( .A(n6176), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U7796 ( .A1(n6300), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6301), .B2(
        n7046), .ZN(n6133) );
  NAND2_X1 U7797 ( .A1(n6134), .A2(n6133), .ZN(n7838) );
  XNOR2_X1 U7798 ( .A(n7838), .B(n8711), .ZN(n6146) );
  NAND2_X1 U7799 ( .A1(n6122), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6141) );
  INV_X2 U7800 ( .A(n6682), .ZN(n6667) );
  INV_X1 U7801 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7802 ( .A1(n6667), .A2(n6135), .ZN(n6140) );
  NAND2_X1 U7803 ( .A1(n6136), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6137) );
  AND2_X1 U7804 ( .A1(n6168), .A2(n6137), .ZN(n7844) );
  OR2_X1 U7805 ( .A1(n6226), .A2(n7844), .ZN(n6139) );
  OR2_X1 U7806 ( .A1(n6444), .A2(n4897), .ZN(n6138) );
  AND4_X2 U7807 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n8009)
         );
  XNOR2_X1 U7808 ( .A(n6146), .B(n8009), .ZN(n7832) );
  INV_X1 U7809 ( .A(n6142), .ZN(n6143) );
  NAND2_X1 U7810 ( .A1(n6143), .A2(n8874), .ZN(n7828) );
  INV_X1 U7811 ( .A(n7828), .ZN(n6144) );
  NAND2_X1 U7812 ( .A1(n6146), .A2(n8009), .ZN(n6147) );
  NAND2_X1 U7813 ( .A1(n7192), .A2(n6675), .ZN(n6162) );
  INV_X1 U7814 ( .A(n6148), .ZN(n6150) );
  NOR2_X1 U7815 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6149) );
  AOI21_X1 U7816 ( .B1(n6150), .B2(n6149), .A(n9439), .ZN(n6151) );
  MUX2_X1 U7817 ( .A(n9439), .B(n6151), .S(P2_IR_REG_9__SCAN_IN), .Z(n6160) );
  NAND2_X1 U7818 ( .A1(n6152), .A2(n6153), .ZN(n6156) );
  INV_X1 U7819 ( .A(n6154), .ZN(n6155) );
  NOR2_X1 U7820 ( .A1(n6156), .A2(n6155), .ZN(n6159) );
  INV_X1 U7821 ( .A(n6157), .ZN(n6158) );
  INV_X1 U7822 ( .A(n7202), .ZN(n7603) );
  AOI22_X1 U7823 ( .A1(n6300), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6301), .B2(
        n7603), .ZN(n6161) );
  NAND2_X1 U7824 ( .A1(n6162), .A2(n6161), .ZN(n8109) );
  XNOR2_X1 U7825 ( .A(n8109), .B(n8711), .ZN(n8052) );
  NAND2_X1 U7826 ( .A1(n6170), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6163) );
  AND2_X1 U7827 ( .A1(n6186), .A2(n6163), .ZN(n8110) );
  OR2_X1 U7828 ( .A1(n6226), .A2(n8110), .ZN(n6167) );
  INV_X1 U7829 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10468) );
  OR2_X1 U7830 ( .A1(n6444), .A2(n10468), .ZN(n6166) );
  NAND2_X1 U7831 ( .A1(n6682), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7832 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n8871)
         );
  INV_X1 U7833 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10376) );
  OR2_X1 U7834 ( .A1(n6670), .A2(n10376), .ZN(n6174) );
  NAND2_X1 U7835 ( .A1(n6168), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6169) );
  AND2_X1 U7836 ( .A1(n6170), .A2(n6169), .ZN(n8016) );
  OR2_X1 U7837 ( .A1(n6226), .A2(n8016), .ZN(n6173) );
  NAND2_X1 U7838 ( .A1(n6682), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7839 ( .A1(n6125), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7840 ( .A1(n7182), .A2(n6675), .ZN(n6180) );
  INV_X1 U7841 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7842 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  NAND2_X1 U7843 ( .A1(n6177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7844 ( .A(n6178), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7162) );
  AOI22_X1 U7845 ( .A1(n6300), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6301), .B2(
        n7162), .ZN(n6179) );
  NAND2_X1 U7846 ( .A1(n6180), .A2(n6179), .ZN(n8013) );
  XNOR2_X1 U7847 ( .A(n8013), .B(n8711), .ZN(n6181) );
  AOI22_X1 U7848 ( .A1(n8052), .A2(n8096), .B1(n8007), .B2(n6181), .ZN(n6185)
         );
  AOI21_X1 U7849 ( .B1(n8050), .B2(n8872), .A(n8871), .ZN(n6183) );
  NAND3_X1 U7850 ( .A1(n8050), .A2(n8871), .A3(n8872), .ZN(n6182) );
  OAI21_X1 U7851 ( .B1(n8052), .B2(n6183), .A(n6182), .ZN(n6184) );
  NAND2_X1 U7852 ( .A1(n6122), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7853 ( .A1(n6186), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6187) );
  AND2_X1 U7854 ( .A1(n6205), .A2(n6187), .ZN(n8244) );
  OR2_X1 U7855 ( .A1(n6226), .A2(n8244), .ZN(n6190) );
  NAND2_X1 U7856 ( .A1(n6682), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7857 ( .A1(n6681), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6188) );
  NAND4_X1 U7858 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n8870)
         );
  NAND2_X1 U7859 ( .A1(n7224), .A2(n6675), .ZN(n6196) );
  INV_X1 U7860 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7861 ( .A1(n6193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  AOI22_X1 U7862 ( .A1(n6300), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6301), .B2(
        n7088), .ZN(n6195) );
  XNOR2_X1 U7863 ( .A(n8091), .B(n4553), .ZN(n8083) );
  NAND2_X1 U7864 ( .A1(n8080), .A2(n8083), .ZN(n6198) );
  NAND2_X1 U7865 ( .A1(n7230), .A2(n6675), .ZN(n6204) );
  NAND2_X1 U7866 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7867 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6200), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n6202) );
  NAND2_X1 U7868 ( .A1(n6202), .A2(n6201), .ZN(n7859) );
  INV_X1 U7869 ( .A(n7859), .ZN(n7097) );
  AOI22_X1 U7870 ( .A1(n6300), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6301), .B2(
        n7097), .ZN(n6203) );
  INV_X1 U7871 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10564) );
  OR2_X1 U7872 ( .A1(n6667), .A2(n10564), .ZN(n6210) );
  NAND2_X1 U7873 ( .A1(n6205), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6206) );
  AND2_X1 U7874 ( .A1(n6214), .A2(n6206), .ZN(n8187) );
  OR2_X1 U7875 ( .A1(n6226), .A2(n8187), .ZN(n6209) );
  NAND2_X1 U7876 ( .A1(n6122), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7877 ( .A1(n6681), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6207) );
  NAND4_X1 U7878 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n8869)
         );
  XNOR2_X1 U7879 ( .A(n8188), .B(n8869), .ZN(n6697) );
  XNOR2_X1 U7880 ( .A(n6697), .B(n8711), .ZN(n8210) );
  NAND2_X1 U7881 ( .A1(n7338), .A2(n6675), .ZN(n6213) );
  NAND2_X1 U7882 ( .A1(n6201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6211) );
  XNOR2_X1 U7883 ( .A(n6211), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7125) );
  AOI22_X1 U7884 ( .A1(n6300), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6301), .B2(
        n7125), .ZN(n6212) );
  NAND2_X2 U7885 ( .A1(n6213), .A2(n6212), .ZN(n9328) );
  XNOR2_X1 U7886 ( .A(n9328), .B(n4553), .ZN(n8285) );
  NAND2_X1 U7887 ( .A1(n6122), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7888 ( .A1(n6214), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6215) );
  AND2_X1 U7889 ( .A1(n6223), .A2(n6215), .ZN(n8291) );
  OR2_X1 U7890 ( .A1(n6226), .A2(n8291), .ZN(n6218) );
  NAND2_X1 U7891 ( .A1(n6682), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7892 ( .A1(n6681), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6216) );
  NAND4_X1 U7893 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n9237)
         );
  NAND2_X1 U7894 ( .A1(n8285), .A2(n9237), .ZN(n6231) );
  NAND2_X1 U7895 ( .A1(n7347), .A2(n6675), .ZN(n6222) );
  XNOR2_X1 U7896 ( .A(n6220), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8155) );
  AOI22_X1 U7897 ( .A1(n6300), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6301), .B2(
        n8155), .ZN(n6221) );
  XNOR2_X1 U7898 ( .A(n9428), .B(n4553), .ZN(n6237) );
  INV_X1 U7899 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10355) );
  OR2_X1 U7900 ( .A1(n6667), .A2(n10355), .ZN(n6230) );
  NAND2_X1 U7901 ( .A1(n6223), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6224) );
  AND2_X1 U7902 ( .A1(n6225), .A2(n6224), .ZN(n9241) );
  OR2_X1 U7903 ( .A1(n6226), .A2(n9241), .ZN(n6229) );
  NAND2_X1 U7904 ( .A1(n6122), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7905 ( .A1(n6681), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6227) );
  NAND4_X1 U7906 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n9225)
         );
  XNOR2_X1 U7907 ( .A(n6237), .B(n9260), .ZN(n8314) );
  INV_X1 U7908 ( .A(n8210), .ZN(n8287) );
  NAND3_X1 U7909 ( .A1(n6231), .A2(n8287), .A3(n9258), .ZN(n6233) );
  INV_X1 U7910 ( .A(n8285), .ZN(n6232) );
  NAND2_X1 U7911 ( .A1(n6232), .A2(n8284), .ZN(n8311) );
  AND2_X1 U7912 ( .A1(n6233), .A2(n8311), .ZN(n6234) );
  NAND2_X1 U7913 ( .A1(n6236), .A2(n6235), .ZN(n8313) );
  XNOR2_X1 U7914 ( .A(n6239), .B(n9238), .ZN(n8277) );
  NAND2_X1 U7915 ( .A1(n7360), .A2(n6675), .ZN(n6244) );
  NAND2_X1 U7916 ( .A1(n6241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7917 ( .A(n6242), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8928) );
  AOI22_X1 U7918 ( .A1(n6300), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6301), .B2(
        n8928), .ZN(n6243) );
  XNOR2_X1 U7919 ( .A(n9417), .B(n4553), .ZN(n6253) );
  NAND2_X1 U7920 ( .A1(n6247), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7921 ( .A1(n6263), .A2(n6248), .ZN(n9218) );
  NAND2_X1 U7922 ( .A1(n9218), .A2(n6659), .ZN(n6252) );
  NAND2_X1 U7923 ( .A1(n6122), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7924 ( .A1(n6682), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7925 ( .A1(n6681), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6249) );
  NAND4_X1 U7926 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n9226)
         );
  XNOR2_X1 U7927 ( .A(n6253), .B(n6804), .ZN(n8857) );
  INV_X1 U7928 ( .A(n6253), .ZN(n6254) );
  NAND2_X1 U7929 ( .A1(n8856), .A2(n4449), .ZN(n8797) );
  NAND2_X1 U7930 ( .A1(n7391), .A2(n6675), .ZN(n6261) );
  INV_X1 U7931 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7932 ( .A1(n6256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6257) );
  MUX2_X1 U7933 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6257), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6259) );
  INV_X1 U7934 ( .A(n6258), .ZN(n6271) );
  AOI22_X1 U7935 ( .A1(n6300), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6301), .B2(
        n8937), .ZN(n6260) );
  NAND2_X1 U7936 ( .A1(n6261), .A2(n6260), .ZN(n8794) );
  XNOR2_X1 U7937 ( .A(n8794), .B(n4553), .ZN(n6268) );
  INV_X1 U7938 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7939 ( .A1(n6263), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7940 ( .A1(n6277), .A2(n6264), .ZN(n9202) );
  NAND2_X1 U7941 ( .A1(n9202), .A2(n6659), .ZN(n6267) );
  AOI22_X1 U7942 ( .A1(n6681), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6682), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7943 ( .A1(n6122), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6265) );
  XNOR2_X1 U7944 ( .A(n6268), .B(n9214), .ZN(n8796) );
  NAND2_X1 U7945 ( .A1(n7408), .A2(n6675), .ZN(n6274) );
  NAND2_X1 U7946 ( .A1(n6271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U7947 ( .A(n6272), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8980) );
  AOI22_X1 U7948 ( .A1(n6300), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6301), .B2(
        n8980), .ZN(n6273) );
  XNOR2_X1 U7949 ( .A(n9406), .B(n4553), .ZN(n6282) );
  NAND2_X1 U7950 ( .A1(n6277), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7951 ( .A1(n6287), .A2(n6278), .ZN(n9191) );
  NAND2_X1 U7952 ( .A1(n9191), .A2(n6659), .ZN(n6281) );
  AOI22_X1 U7953 ( .A1(n6681), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6682), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7954 ( .A1(n6122), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6279) );
  XNOR2_X1 U7955 ( .A(n6282), .B(n9163), .ZN(n8805) );
  NAND2_X1 U7956 ( .A1(n8802), .A2(n6283), .ZN(n8833) );
  NAND2_X1 U7957 ( .A1(n7511), .A2(n6675), .ZN(n6286) );
  NAND2_X1 U7958 ( .A1(n6284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U7959 ( .A(n6297), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8993) );
  AOI22_X1 U7960 ( .A1(n6300), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8993), .B2(
        n6301), .ZN(n6285) );
  XNOR2_X1 U7961 ( .A(n9170), .B(n4553), .ZN(n6294) );
  NAND2_X1 U7962 ( .A1(n6287), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7963 ( .A1(n6304), .A2(n6288), .ZN(n9166) );
  NAND2_X1 U7964 ( .A1(n9166), .A2(n6659), .ZN(n6293) );
  INV_X1 U7965 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U7966 ( .A1(n6122), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7967 ( .A1(n6681), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6289) );
  OAI211_X1 U7968 ( .C1(n6667), .C2(n10445), .A(n6290), .B(n6289), .ZN(n6291)
         );
  INV_X1 U7969 ( .A(n6291), .ZN(n6292) );
  INV_X1 U7970 ( .A(n9187), .ZN(n9152) );
  XNOR2_X1 U7971 ( .A(n6294), .B(n9152), .ZN(n8834) );
  NAND2_X1 U7972 ( .A1(n8833), .A2(n8834), .ZN(n8832) );
  NAND2_X1 U7973 ( .A1(n7634), .A2(n6675), .ZN(n6303) );
  NAND2_X1 U7974 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  NAND2_X1 U7975 ( .A1(n6298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  AOI22_X1 U7976 ( .A1(n9000), .A2(n6301), .B1(n6300), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7977 ( .A1(n6303), .A2(n6302), .ZN(n9302) );
  XNOR2_X1 U7978 ( .A(n9302), .B(n4553), .ZN(n6311) );
  NAND2_X1 U7979 ( .A1(n6304), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7980 ( .A1(n6316), .A2(n6305), .ZN(n9154) );
  NAND2_X1 U7981 ( .A1(n9154), .A2(n6659), .ZN(n6310) );
  INV_X1 U7982 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U7983 ( .A1(n6122), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6307) );
  INV_X1 U7984 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10486) );
  OR2_X1 U7985 ( .A1(n6667), .A2(n10486), .ZN(n6306) );
  OAI211_X1 U7986 ( .C1(n10476), .C2(n6444), .A(n6307), .B(n6306), .ZN(n6308)
         );
  INV_X1 U7987 ( .A(n6308), .ZN(n6309) );
  XNOR2_X1 U7988 ( .A(n6311), .B(n9164), .ZN(n8772) );
  NAND2_X1 U7989 ( .A1(n7822), .A2(n6675), .ZN(n6314) );
  INV_X1 U7990 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7825) );
  OR2_X1 U7991 ( .A1(n6678), .A2(n7825), .ZN(n6313) );
  XNOR2_X1 U7992 ( .A(n8823), .B(n4553), .ZN(n6321) );
  INV_X1 U7993 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U7994 ( .A1(n6316), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7995 ( .A1(n6327), .A2(n6317), .ZN(n9141) );
  INV_X1 U7996 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U7997 ( .A1(n6681), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7998 ( .A1(n6682), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6318) );
  OAI211_X1 U7999 ( .C1(n6670), .C2(n10489), .A(n6319), .B(n6318), .ZN(n6320)
         );
  XNOR2_X1 U8000 ( .A(n6321), .B(n9153), .ZN(n8826) );
  NAND2_X1 U8001 ( .A1(n7908), .A2(n6675), .ZN(n6324) );
  OR2_X1 U8002 ( .A1(n6678), .A2(n7910), .ZN(n6323) );
  XNOR2_X1 U8003 ( .A(n9392), .B(n4553), .ZN(n6332) );
  NAND2_X1 U8004 ( .A1(n6327), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U8005 ( .A1(n6336), .A2(n6328), .ZN(n9129) );
  INV_X1 U8006 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U8007 ( .A1(n6122), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8008 ( .A1(n6682), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6329) );
  OAI211_X1 U8009 ( .C1(n9128), .C2(n6444), .A(n6330), .B(n6329), .ZN(n6331)
         );
  XNOR2_X1 U8010 ( .A(n6332), .B(n9136), .ZN(n8779) );
  INV_X1 U8011 ( .A(n6332), .ZN(n6333) );
  NAND2_X1 U8012 ( .A1(n8023), .A2(n6675), .ZN(n6335) );
  OR2_X1 U8013 ( .A1(n6678), .A2(n8025), .ZN(n6334) );
  XNOR2_X1 U8014 ( .A(n9386), .B(n4553), .ZN(n6343) );
  NAND2_X1 U8015 ( .A1(n6336), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U8016 ( .A1(n6356), .A2(n6337), .ZN(n9112) );
  NAND2_X1 U8017 ( .A1(n9112), .A2(n6659), .ZN(n6342) );
  INV_X1 U8018 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U8019 ( .A1(n6681), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U8020 ( .A1(n6682), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6338) );
  OAI211_X1 U8021 ( .C1(n6670), .C2(n10565), .A(n6339), .B(n6338), .ZN(n6340)
         );
  INV_X1 U8022 ( .A(n6340), .ZN(n6341) );
  XNOR2_X1 U8023 ( .A(n6343), .B(n8782), .ZN(n8372) );
  NAND2_X1 U8024 ( .A1(n6343), .A2(n9126), .ZN(n6344) );
  NAND2_X1 U8025 ( .A1(n8218), .A2(n6675), .ZN(n6346) );
  OR2_X1 U8026 ( .A1(n6678), .A2(n8221), .ZN(n6345) );
  XNOR2_X1 U8027 ( .A(n9375), .B(n4553), .ZN(n8814) );
  INV_X1 U8028 ( .A(n8814), .ZN(n6367) );
  NAND2_X1 U8029 ( .A1(n6358), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8030 ( .A1(n6372), .A2(n6348), .ZN(n9085) );
  NAND2_X1 U8031 ( .A1(n9085), .A2(n6659), .ZN(n6353) );
  INV_X1 U8032 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U8033 ( .A1(n6122), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U8034 ( .A1(n6681), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6349) );
  OAI211_X1 U8035 ( .C1(n6667), .C2(n10508), .A(n6350), .B(n6349), .ZN(n6351)
         );
  INV_X1 U8036 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U8037 ( .A1(n8066), .A2(n6675), .ZN(n6355) );
  OR2_X1 U8038 ( .A1(n6678), .A2(n10523), .ZN(n6354) );
  INV_X1 U8039 ( .A(n8812), .ZN(n6364) );
  NAND2_X1 U8040 ( .A1(n6356), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U8041 ( .A1(n6358), .A2(n6357), .ZN(n9098) );
  NAND2_X1 U8042 ( .A1(n9098), .A2(n6659), .ZN(n6363) );
  INV_X1 U8043 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U8044 ( .A1(n6681), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8045 ( .A1(n6122), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6359) );
  OAI211_X1 U8046 ( .C1(n6667), .C2(n10548), .A(n6360), .B(n6359), .ZN(n6361)
         );
  INV_X1 U8047 ( .A(n6361), .ZN(n6362) );
  OAI22_X1 U8048 ( .A1(n6367), .A2(n8790), .B1(n6364), .B2(n8817), .ZN(n6369)
         );
  OAI21_X1 U8049 ( .B1(n8812), .B2(n9109), .A(n9095), .ZN(n6366) );
  NOR3_X1 U8050 ( .A1(n8812), .A2(n9095), .A3(n9109), .ZN(n6365) );
  AOI21_X1 U8051 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6368) );
  NAND2_X1 U8052 ( .A1(n8269), .A2(n6675), .ZN(n6371) );
  OR2_X1 U8053 ( .A1(n6678), .A2(n8270), .ZN(n6370) );
  XNOR2_X1 U8054 ( .A(n9370), .B(n8711), .ZN(n6387) );
  NAND2_X1 U8055 ( .A1(n6372), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8056 ( .A1(n6381), .A2(n6373), .ZN(n9071) );
  NAND2_X1 U8057 ( .A1(n9071), .A2(n6659), .ZN(n6378) );
  INV_X1 U8058 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U8059 ( .A1(n6122), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8060 ( .A1(n6682), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6374) );
  OAI211_X1 U8061 ( .C1(n9075), .C2(n6444), .A(n6375), .B(n6374), .ZN(n6376)
         );
  INV_X1 U8062 ( .A(n6376), .ZN(n6377) );
  XNOR2_X1 U8063 ( .A(n6387), .B(n9083), .ZN(n8787) );
  NAND2_X1 U8064 ( .A1(n8332), .A2(n6675), .ZN(n6380) );
  OR2_X1 U8065 ( .A1(n6678), .A2(n8333), .ZN(n6379) );
  XNOR2_X1 U8066 ( .A(n9364), .B(n4553), .ZN(n8842) );
  NAND2_X1 U8067 ( .A1(n6381), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8068 ( .A1(n6397), .A2(n6382), .ZN(n9065) );
  INV_X1 U8069 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U8070 ( .A1(n6122), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8071 ( .A1(n6682), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6383) );
  OAI211_X1 U8072 ( .C1(n9064), .C2(n6444), .A(n6384), .B(n6383), .ZN(n6385)
         );
  INV_X1 U8073 ( .A(n6385), .ZN(n6386) );
  NAND2_X1 U8074 ( .A1(n6387), .A2(n8849), .ZN(n8840) );
  INV_X1 U8075 ( .A(n6388), .ZN(n6389) );
  NAND2_X1 U8076 ( .A1(n8841), .A2(n6389), .ZN(n6391) );
  NAND2_X1 U8077 ( .A1(n8842), .A2(n9069), .ZN(n6390) );
  NAND2_X1 U8078 ( .A1(n6391), .A2(n6390), .ZN(n6437) );
  INV_X1 U8079 ( .A(n6437), .ZN(n6405) );
  NAND2_X1 U8080 ( .A1(n8703), .A2(n6675), .ZN(n6394) );
  OR2_X1 U8081 ( .A1(n6678), .A2(n6392), .ZN(n6393) );
  XNOR2_X1 U8082 ( .A(n9358), .B(n8711), .ZN(n8722) );
  INV_X1 U8083 ( .A(n6397), .ZN(n6396) );
  INV_X1 U8084 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8085 ( .A1(n6397), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8086 ( .A1(n6440), .A2(n6398), .ZN(n9056) );
  NAND2_X1 U8087 ( .A1(n9056), .A2(n6659), .ZN(n6403) );
  INV_X1 U8088 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U8089 ( .A1(n6682), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8090 ( .A1(n6122), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6399) );
  OAI211_X1 U8091 ( .C1(n9055), .C2(n6444), .A(n6400), .B(n6399), .ZN(n6401)
         );
  INV_X1 U8092 ( .A(n6401), .ZN(n6402) );
  NOR2_X1 U8093 ( .A1(n8722), .A2(n8723), .ZN(n8716) );
  AOI21_X1 U8094 ( .B1(n8722), .B2(n8723), .A(n8716), .ZN(n6436) );
  INV_X1 U8095 ( .A(n6436), .ZN(n6404) );
  NAND2_X1 U8096 ( .A1(n6405), .A2(n6404), .ZN(n6438) );
  NAND2_X1 U8097 ( .A1(n8271), .A2(n6408), .ZN(n6409) );
  NAND2_X1 U8098 ( .A1(n6411), .A2(n7189), .ZN(n7526) );
  INV_X1 U8099 ( .A(n6951), .ZN(n6426) );
  NOR2_X1 U8100 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .ZN(
        n6415) );
  NOR4_X1 U8101 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6414) );
  NOR4_X1 U8102 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6413) );
  NOR4_X1 U8103 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6412) );
  NAND4_X1 U8104 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n6421)
         );
  NOR4_X1 U8105 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6419) );
  NOR4_X1 U8106 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6418) );
  NOR4_X1 U8107 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6417) );
  NOR4_X1 U8108 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6416) );
  NAND4_X1 U8109 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n6420)
         );
  NOR2_X1 U8110 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  INV_X1 U8111 ( .A(n6423), .ZN(n6429) );
  NAND2_X1 U8112 ( .A1(n6429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8113 ( .A1(n6427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6428) );
  MUX2_X1 U8114 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6428), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n6430) );
  NAND2_X1 U8115 ( .A1(n9000), .A2(n6952), .ZN(n6928) );
  NOR2_X1 U8116 ( .A1(n9053), .A2(n9329), .ZN(n6431) );
  NAND2_X1 U8117 ( .A1(n6433), .A2(n6431), .ZN(n6455) );
  INV_X1 U8118 ( .A(n6455), .ZN(n6432) );
  NAND2_X1 U8119 ( .A1(n6939), .A2(n6432), .ZN(n6435) );
  NAND3_X1 U8120 ( .A1(n7528), .A2(n7526), .A3(n6453), .ZN(n6461) );
  OR2_X1 U8121 ( .A1(n6433), .A2(n4797), .ZN(n6937) );
  INV_X1 U8122 ( .A(n6937), .ZN(n6457) );
  NAND2_X1 U8123 ( .A1(n6941), .A2(n6457), .ZN(n6434) );
  NAND3_X1 U8124 ( .A1(n6438), .A2(n8855), .A3(n8729), .ZN(n6468) );
  INV_X1 U8125 ( .A(n9358), .ZN(n6924) );
  NAND2_X1 U8126 ( .A1(n6939), .A2(n9329), .ZN(n6439) );
  NAND2_X1 U8127 ( .A1(n6440), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8128 ( .A1(n8705), .A2(n6441), .ZN(n9045) );
  NAND2_X1 U8129 ( .A1(n9045), .A2(n6659), .ZN(n6447) );
  INV_X1 U8130 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U8131 ( .A1(n6122), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8132 ( .A1(n6682), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6442) );
  OAI211_X1 U8133 ( .C1(n9044), .C2(n6444), .A(n6443), .B(n6442), .ZN(n6445)
         );
  INV_X1 U8134 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8135 ( .A1(n9017), .A2(n7827), .ZN(n6458) );
  INV_X1 U8136 ( .A(n6449), .ZN(n7074) );
  NAND2_X1 U8137 ( .A1(n9009), .A2(n7074), .ZN(n6450) );
  INV_X1 U8138 ( .A(n9050), .ZN(n6933) );
  NOR2_X1 U8139 ( .A1(n7522), .A2(n6933), .ZN(n6451) );
  NOR2_X1 U8140 ( .A1(n7522), .A2(n9050), .ZN(n6452) );
  NAND2_X1 U8141 ( .A1(n6941), .A2(n6452), .ZN(n8848) );
  INV_X1 U8142 ( .A(n6453), .ZN(n6456) );
  NAND2_X1 U8143 ( .A1(n9329), .A2(n6454), .ZN(n9242) );
  NAND2_X1 U8144 ( .A1(n6455), .A2(n9242), .ZN(n6940) );
  OAI21_X1 U8145 ( .B1(n6456), .B2(n6951), .A(n6940), .ZN(n6460) );
  NAND2_X1 U8146 ( .A1(n6457), .A2(n6461), .ZN(n6459) );
  NAND2_X1 U8147 ( .A1(n6458), .A2(n9053), .ZN(n6949) );
  NAND4_X1 U8148 ( .A1(n6460), .A2(n6459), .A3(n7070), .A4(n6949), .ZN(n6462)
         );
  NOR2_X1 U8149 ( .A1(n7522), .A2(n7181), .ZN(n6875) );
  AOI22_X1 U8150 ( .A1(n6462), .A2(P2_STATE_REG_SCAN_IN), .B1(n6875), .B2(
        n6461), .ZN(n7343) );
  NOR2_X1 U8151 ( .A1(n7068), .A2(P2_U3151), .ZN(n6873) );
  INV_X1 U8152 ( .A(n6873), .ZN(n8063) );
  AOI22_X1 U8153 ( .A1(n9056), .A2(n8863), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6463) );
  OAI21_X1 U8154 ( .B1(n6920), .B2(n8848), .A(n6463), .ZN(n6464) );
  AOI21_X1 U8155 ( .B1(n9051), .B2(n8845), .A(n6464), .ZN(n6465) );
  INV_X1 U8156 ( .A(n6466), .ZN(n6467) );
  NAND2_X1 U8157 ( .A1(n6468), .A2(n6467), .ZN(P2_U3154) );
  NOR2_X1 U8158 ( .A1(n6538), .A2(n7448), .ZN(n7725) );
  NAND4_X1 U8159 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6474)
         );
  INV_X1 U8160 ( .A(n7651), .ZN(n9631) );
  NAND2_X1 U8161 ( .A1(n9631), .A2(n7818), .ZN(n8414) );
  NAND2_X1 U8162 ( .A1(n7813), .A2(n8592), .ZN(n7650) );
  NAND2_X1 U8163 ( .A1(n7650), .A2(n8593), .ZN(n6476) );
  NAND2_X1 U8164 ( .A1(n8417), .A2(n5228), .ZN(n8598) );
  INV_X1 U8165 ( .A(n8417), .ZN(n9630) );
  NAND2_X1 U8166 ( .A1(n8598), .A2(n8597), .ZN(n8540) );
  INV_X1 U8167 ( .A(n8540), .ZN(n7661) );
  NAND2_X1 U8168 ( .A1(n8423), .A2(n10145), .ZN(n8599) );
  INV_X1 U8169 ( .A(n8599), .ZN(n6477) );
  NAND2_X1 U8170 ( .A1(n7960), .A2(n7978), .ZN(n7955) );
  NAND2_X1 U8171 ( .A1(n8030), .A2(n8142), .ZN(n8442) );
  AND2_X1 U8172 ( .A1(n7955), .A2(n8442), .ZN(n8596) );
  NAND2_X1 U8173 ( .A1(n8367), .A2(n7959), .ZN(n8602) );
  INV_X1 U8174 ( .A(n8423), .ZN(n9629) );
  NAND2_X1 U8175 ( .A1(n8433), .A2(n8437), .ZN(n6479) );
  NAND2_X1 U8176 ( .A1(n8596), .A2(n6479), .ZN(n6480) );
  NAND2_X1 U8177 ( .A1(n8441), .A2(n6480), .ZN(n6481) );
  NAND2_X1 U8178 ( .A1(n6481), .A2(n8602), .ZN(n8610) );
  OR2_X1 U8179 ( .A1(n8205), .A2(n8160), .ZN(n8605) );
  NAND2_X1 U8180 ( .A1(n8205), .A2(n8160), .ZN(n8450) );
  NAND2_X1 U8181 ( .A1(n8605), .A2(n8450), .ZN(n7946) );
  NAND2_X1 U8182 ( .A1(n6483), .A2(n6482), .ZN(n8164) );
  INV_X1 U8183 ( .A(n9625), .ZN(n8000) );
  OR2_X1 U8184 ( .A1(n10062), .A2(n8000), .ZN(n8453) );
  NAND2_X1 U8185 ( .A1(n10062), .A2(n8000), .ZN(n8451) );
  NAND2_X1 U8186 ( .A1(n8453), .A2(n8451), .ZN(n8544) );
  INV_X1 U8187 ( .A(n8450), .ZN(n8445) );
  NOR2_X1 U8188 ( .A1(n8544), .A2(n8445), .ZN(n6484) );
  NAND2_X1 U8189 ( .A1(n8164), .A2(n6484), .ZN(n8165) );
  NAND2_X1 U8190 ( .A1(n8165), .A2(n8453), .ZN(n9962) );
  NAND2_X1 U8191 ( .A1(n10053), .A2(n8161), .ZN(n8613) );
  INV_X1 U8192 ( .A(n9623), .ZN(n8001) );
  OR2_X1 U8193 ( .A1(n10049), .A2(n8001), .ZN(n8458) );
  NAND2_X1 U8194 ( .A1(n10049), .A2(n8001), .ZN(n8612) );
  INV_X1 U8195 ( .A(n9622), .ZN(n8073) );
  OR2_X1 U8196 ( .A1(n10042), .A2(n8073), .ZN(n8465) );
  NAND2_X1 U8197 ( .A1(n10042), .A2(n8073), .ZN(n8459) );
  NAND2_X1 U8198 ( .A1(n8465), .A2(n8459), .ZN(n8549) );
  INV_X1 U8199 ( .A(n8612), .ZN(n6485) );
  OR2_X1 U8200 ( .A1(n9936), .A2(n8341), .ZN(n8462) );
  INV_X1 U8201 ( .A(n9621), .ZN(n8411) );
  OR2_X1 U8202 ( .A1(n10039), .A2(n8411), .ZN(n8531) );
  NAND2_X1 U8203 ( .A1(n8462), .A2(n8531), .ZN(n8620) );
  NAND2_X1 U8204 ( .A1(n8462), .A2(n9929), .ZN(n6486) );
  NAND2_X1 U8205 ( .A1(n9936), .A2(n8341), .ZN(n8619) );
  AND2_X1 U8206 ( .A1(n6486), .A2(n8619), .ZN(n8410) );
  INV_X1 U8207 ( .A(n9619), .ZN(n6487) );
  OR2_X1 U8208 ( .A1(n9917), .A2(n6487), .ZN(n8475) );
  NAND2_X1 U8209 ( .A1(n9917), .A2(n6487), .ZN(n8470) );
  INV_X1 U8210 ( .A(n9618), .ZN(n8399) );
  OR2_X1 U8211 ( .A1(n10023), .A2(n8399), .ZN(n8476) );
  NAND2_X1 U8212 ( .A1(n10023), .A2(n8399), .ZN(n8477) );
  NAND2_X1 U8213 ( .A1(n6488), .A2(n8477), .ZN(n8397) );
  INV_X1 U8214 ( .A(n9617), .ZN(n6489) );
  OR2_X1 U8215 ( .A1(n10018), .A2(n6489), .ZN(n8479) );
  NAND2_X1 U8216 ( .A1(n10018), .A2(n6489), .ZN(n8625) );
  NAND2_X1 U8217 ( .A1(n8397), .A2(n8555), .ZN(n6490) );
  NAND2_X1 U8218 ( .A1(n6490), .A2(n8625), .ZN(n8654) );
  INV_X1 U8219 ( .A(n9615), .ZN(n8483) );
  OR2_X1 U8220 ( .A1(n9876), .A2(n8483), .ZN(n8480) );
  INV_X1 U8221 ( .A(n9616), .ZN(n8400) );
  OR2_X1 U8222 ( .A1(n10014), .A2(n8400), .ZN(n8486) );
  AND2_X1 U8223 ( .A1(n8480), .A2(n8486), .ZN(n8581) );
  NAND2_X1 U8224 ( .A1(n8654), .A2(n8581), .ZN(n6492) );
  NAND2_X1 U8225 ( .A1(n9876), .A2(n8483), .ZN(n8472) );
  NAND2_X1 U8226 ( .A1(n10014), .A2(n8400), .ZN(n9865) );
  NAND2_X1 U8227 ( .A1(n8472), .A2(n9865), .ZN(n6491) );
  NAND2_X1 U8228 ( .A1(n6491), .A2(n8480), .ZN(n8633) );
  NAND2_X1 U8229 ( .A1(n6492), .A2(n8633), .ZN(n9851) );
  INV_X1 U8230 ( .A(n9614), .ZN(n6493) );
  NAND2_X1 U8231 ( .A1(n9851), .A2(n8490), .ZN(n6494) );
  NAND2_X1 U8232 ( .A1(n9857), .A2(n6493), .ZN(n8634) );
  NAND2_X1 U8233 ( .A1(n6494), .A2(n8634), .ZN(n9836) );
  INV_X1 U8234 ( .A(n9613), .ZN(n6495) );
  OR2_X1 U8235 ( .A1(n9844), .A2(n6495), .ZN(n8494) );
  NAND2_X1 U8236 ( .A1(n9844), .A2(n6495), .ZN(n8635) );
  INV_X1 U8237 ( .A(n9612), .ZN(n6496) );
  OR2_X2 U8238 ( .A1(n9991), .A2(n6496), .ZN(n8576) );
  NAND2_X1 U8239 ( .A1(n9991), .A2(n6496), .ZN(n8636) );
  NAND2_X1 U8240 ( .A1(n8576), .A2(n8636), .ZN(n9825) );
  INV_X1 U8241 ( .A(n9611), .ZN(n6498) );
  NAND2_X1 U8242 ( .A1(n9812), .A2(n6498), .ZN(n8637) );
  XNOR2_X1 U8243 ( .A(n9981), .B(n6499), .ZN(n9795) );
  NAND2_X1 U8244 ( .A1(n9981), .A2(n6499), .ZN(n8655) );
  NAND2_X1 U8245 ( .A1(n9782), .A2(n9594), .ZN(n8502) );
  NAND2_X1 U8246 ( .A1(n8630), .A2(n8502), .ZN(n9786) );
  OR2_X2 U8247 ( .A1(n9775), .A2(n9786), .ZN(n9774) );
  INV_X1 U8248 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6655) );
  MUX2_X1 U8249 ( .A(n6655), .B(n10588), .S(n7193), .Z(n6505) );
  INV_X1 U8250 ( .A(SI_28_), .ZN(n6504) );
  NAND2_X1 U8251 ( .A1(n6505), .A2(n6504), .ZN(n6514) );
  INV_X1 U8252 ( .A(n6505), .ZN(n6506) );
  NAND2_X1 U8253 ( .A1(n6506), .A2(SI_28_), .ZN(n6507) );
  NAND2_X1 U8254 ( .A1(n6654), .A2(n6615), .ZN(n6509) );
  OR2_X1 U8255 ( .A1(n5781), .A2(n10588), .ZN(n6508) );
  NAND2_X1 U8256 ( .A1(n9767), .A2(n8739), .ZN(n8503) );
  AND2_X2 U8257 ( .A1(n8573), .A2(n8503), .ZN(n8561) );
  MUX2_X1 U8258 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7193), .Z(n6603) );
  XNOR2_X1 U8259 ( .A(n6603), .B(SI_29_), .ZN(n6515) );
  INV_X1 U8260 ( .A(n6515), .ZN(n6512) );
  OAI21_X1 U8261 ( .B1(n4452), .B2(n4969), .A(n6515), .ZN(n6516) );
  INV_X1 U8262 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10111) );
  OR2_X1 U8263 ( .A1(n5781), .A2(n10111), .ZN(n6519) );
  OR2_X1 U8264 ( .A1(n8690), .A2(n6521), .ZN(n6527) );
  INV_X1 U8265 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10519) );
  NAND2_X1 U8266 ( .A1(n5410), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8267 ( .A1(n6621), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8268 ( .C1(n10519), .C2(n6524), .A(n6523), .B(n6522), .ZN(n6525)
         );
  INV_X1 U8269 ( .A(n6525), .ZN(n6526) );
  NAND2_X1 U8270 ( .A1(n6527), .A2(n6526), .ZN(n9607) );
  INV_X1 U8271 ( .A(n9607), .ZN(n6528) );
  NAND2_X1 U8272 ( .A1(n8692), .A2(n6528), .ZN(n8644) );
  NAND2_X2 U8273 ( .A1(n8574), .A2(n8644), .ZN(n8687) );
  NAND2_X1 U8274 ( .A1(n5687), .A2(n5224), .ZN(n6530) );
  NAND2_X1 U8275 ( .A1(n6529), .A2(n8675), .ZN(n8523) );
  NAND2_X1 U8276 ( .A1(n6620), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8277 ( .A1(n5410), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8278 ( .A1(n6621), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8279 ( .A1(n7241), .A2(P1_B_REG_SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8280 ( .A1(n9567), .A2(n6534), .ZN(n6625) );
  OAI22_X1 U8281 ( .A1(n8739), .A2(n8398), .B1(n8559), .B2(n6625), .ZN(n6535)
         );
  NAND2_X1 U8282 ( .A1(n6537), .A2(n7733), .ZN(n6539) );
  NAND2_X1 U8283 ( .A1(n6539), .A2(n7726), .ZN(n6542) );
  INV_X2 U8284 ( .A(n7733), .ZN(n10173) );
  NAND3_X1 U8285 ( .A1(n4490), .A2(n6540), .A3(n10173), .ZN(n6541) );
  NAND2_X1 U8286 ( .A1(n6542), .A2(n6541), .ZN(n7638) );
  NAND2_X1 U8287 ( .A1(n8412), .A2(n8589), .ZN(n7636) );
  NAND2_X1 U8288 ( .A1(n7638), .A2(n7636), .ZN(n7637) );
  NAND2_X1 U8289 ( .A1(n6469), .A2(n4416), .ZN(n6543) );
  NAND2_X1 U8290 ( .A1(n7637), .A2(n6543), .ZN(n7810) );
  NOR2_X1 U8291 ( .A1(n9631), .A2(n10180), .ZN(n7647) );
  NOR2_X1 U8292 ( .A1(n6544), .A2(n10156), .ZN(n6545) );
  AOI21_X1 U8293 ( .B1(n8536), .B2(n7647), .A(n6545), .ZN(n6546) );
  NAND2_X1 U8294 ( .A1(n8433), .A2(n8599), .ZN(n7797) );
  AND2_X1 U8295 ( .A1(n8540), .A2(n7797), .ZN(n7915) );
  NAND2_X1 U8296 ( .A1(n7955), .A2(n8437), .ZN(n7916) );
  NOR2_X1 U8297 ( .A1(n9630), .A2(n5228), .ZN(n7795) );
  NOR2_X1 U8298 ( .A1(n9629), .A2(n10145), .ZN(n6547) );
  INV_X1 U8299 ( .A(n7916), .ZN(n8430) );
  NAND2_X1 U8300 ( .A1(n7960), .A2(n6478), .ZN(n6548) );
  OAI21_X1 U8301 ( .B1(n7913), .B2(n8430), .A(n6548), .ZN(n6549) );
  INV_X1 U8302 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8303 ( .A1(n8442), .A2(n8436), .ZN(n7964) );
  NAND2_X1 U8304 ( .A1(n7965), .A2(n7964), .ZN(n7967) );
  NAND2_X1 U8305 ( .A1(n8030), .A2(n8243), .ZN(n6551) );
  NAND2_X1 U8306 ( .A1(n7967), .A2(n6551), .ZN(n8034) );
  NAND2_X1 U8307 ( .A1(n8444), .A2(n8602), .ZN(n8033) );
  NAND2_X1 U8308 ( .A1(n8034), .A2(n8033), .ZN(n8032) );
  OR2_X1 U8309 ( .A1(n8367), .A2(n4609), .ZN(n6552) );
  INV_X1 U8310 ( .A(n8160), .ZN(n9626) );
  NAND2_X1 U8311 ( .A1(n10062), .A2(n9625), .ZN(n6553) );
  OR2_X1 U8312 ( .A1(n10062), .A2(n9625), .ZN(n6554) );
  INV_X1 U8313 ( .A(n8161), .ZN(n9624) );
  NAND2_X1 U8314 ( .A1(n10053), .A2(n9624), .ZN(n6556) );
  NAND2_X1 U8315 ( .A1(n10049), .A2(n9623), .ZN(n6557) );
  NAND2_X1 U8316 ( .A1(n6558), .A2(n6557), .ZN(n8251) );
  AND2_X1 U8317 ( .A1(n10042), .A2(n9622), .ZN(n6560) );
  OR2_X1 U8318 ( .A1(n10042), .A2(n9622), .ZN(n6559) );
  NOR2_X1 U8319 ( .A1(n10039), .A2(n9621), .ZN(n6561) );
  INV_X1 U8320 ( .A(n10039), .ZN(n9954) );
  NAND2_X1 U8321 ( .A1(n8462), .A2(n8619), .ZN(n9933) );
  INV_X1 U8322 ( .A(n8341), .ZN(n9620) );
  NAND2_X1 U8323 ( .A1(n9936), .A2(n9620), .ZN(n6562) );
  OR2_X1 U8324 ( .A1(n9917), .A2(n9619), .ZN(n6563) );
  NOR2_X1 U8325 ( .A1(n10023), .A2(n9618), .ZN(n6564) );
  NAND2_X1 U8326 ( .A1(n10023), .A2(n9618), .ZN(n6565) );
  AND2_X1 U8327 ( .A1(n10018), .A2(n9617), .ZN(n6567) );
  NOR2_X1 U8328 ( .A1(n10014), .A2(n9616), .ZN(n8553) );
  AND2_X1 U8329 ( .A1(n9876), .A2(n9615), .ZN(n8529) );
  OR2_X1 U8330 ( .A1(n9876), .A2(n9615), .ZN(n8528) );
  NOR2_X1 U8331 ( .A1(n9857), .A2(n9614), .ZN(n6569) );
  NAND2_X1 U8332 ( .A1(n9857), .A2(n9614), .ZN(n6568) );
  OAI21_X1 U8333 ( .B1(n9855), .B2(n6569), .A(n6568), .ZN(n9835) );
  AND2_X1 U8334 ( .A1(n9844), .A2(n9613), .ZN(n6570) );
  OAI22_X1 U8335 ( .A1(n9835), .A2(n6570), .B1(n9844), .B2(n9613), .ZN(n9820)
         );
  NOR2_X1 U8336 ( .A1(n9991), .A2(n9612), .ZN(n6572) );
  NAND2_X1 U8337 ( .A1(n9991), .A2(n9612), .ZN(n6571) );
  OAI21_X1 U8338 ( .B1(n9820), .B2(n6572), .A(n6571), .ZN(n9810) );
  AND2_X1 U8339 ( .A1(n9812), .A2(n9611), .ZN(n6573) );
  INV_X1 U8340 ( .A(n9594), .ZN(n9609) );
  OR2_X1 U8341 ( .A1(n9782), .A2(n9609), .ZN(n6574) );
  NAND2_X1 U8342 ( .A1(n8687), .A2(n4670), .ZN(n6586) );
  AND2_X1 U8343 ( .A1(n9767), .A2(n9608), .ZN(n8685) );
  NAND2_X1 U8344 ( .A1(n4668), .A2(n6575), .ZN(n6582) );
  INV_X1 U8345 ( .A(n6582), .ZN(n6576) );
  NAND2_X1 U8346 ( .A1(n6967), .A2(n6576), .ZN(n6585) );
  INV_X1 U8347 ( .A(n8671), .ZN(n6577) );
  OR2_X1 U8348 ( .A1(n6577), .A2(n8571), .ZN(n8568) );
  INV_X1 U8349 ( .A(n7777), .ZN(n6580) );
  NAND2_X1 U8350 ( .A1(n6578), .A2(n8571), .ZN(n6579) );
  NAND3_X1 U8351 ( .A1(n8568), .A2(n6580), .A3(n6579), .ZN(n8159) );
  NAND2_X2 U8352 ( .A1(n5687), .A2(n8026), .ZN(n8518) );
  AOI21_X1 U8353 ( .B1(n8687), .B2(n8685), .A(n10185), .ZN(n6581) );
  OAI21_X1 U8354 ( .B1(n6582), .B2(n4670), .A(n6581), .ZN(n6583) );
  INV_X1 U8355 ( .A(n6583), .ZN(n6584) );
  OAI211_X1 U8356 ( .C1(n6967), .C2(n6586), .A(n6585), .B(n6584), .ZN(n6593)
         );
  NAND2_X1 U8357 ( .A1(n7653), .A2(n8425), .ZN(n7803) );
  NAND2_X1 U8358 ( .A1(n7968), .A2(n4408), .ZN(n7948) );
  INV_X1 U8359 ( .A(n10053), .ZN(n9969) );
  INV_X1 U8360 ( .A(n10049), .ZN(n8129) );
  NAND2_X1 U8361 ( .A1(n8124), .A2(n8129), .ZN(n8125) );
  NAND2_X1 U8362 ( .A1(n9922), .A2(n10092), .ZN(n9898) );
  OR2_X2 U8363 ( .A1(n9898), .A2(n10023), .ZN(n9899) );
  NOR2_X4 U8364 ( .A1(n9899), .A2(n10018), .ZN(n9887) );
  INV_X1 U8365 ( .A(n10014), .ZN(n9894) );
  NOR2_X2 U8366 ( .A1(n9841), .A2(n9991), .ZN(n6589) );
  INV_X1 U8367 ( .A(n6589), .ZN(n9821) );
  AOI21_X1 U8368 ( .B1(n8692), .B2(n6590), .A(n9949), .ZN(n6592) );
  INV_X1 U8369 ( .A(n8390), .ZN(n6591) );
  NAND2_X1 U8370 ( .A1(n6592), .A2(n6591), .ZN(n8694) );
  NAND3_X1 U8371 ( .A1(n8698), .A2(n6593), .A3(n8694), .ZN(n6883) );
  NAND3_X1 U8372 ( .A1(n6595), .A2(P1_STATE_REG_SCAN_IN), .A3(n6594), .ZN(
        n7721) );
  NAND2_X1 U8373 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  NAND2_X1 U8374 ( .A1(n6883), .A2(n10194), .ZN(n6602) );
  OR2_X1 U8375 ( .A1(n10194), .A2(n10519), .ZN(n6599) );
  INV_X1 U8376 ( .A(n6600), .ZN(n6601) );
  INV_X1 U8377 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U8378 ( .A1(n6603), .A2(SI_29_), .ZN(n6604) );
  NAND2_X1 U8379 ( .A1(n6605), .A2(n6604), .ZN(n6611) );
  MUX2_X1 U8380 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7193), .Z(n6609) );
  XNOR2_X1 U8381 ( .A(n6609), .B(SI_30_), .ZN(n6610) );
  XNOR2_X1 U8382 ( .A(n6611), .B(n6610), .ZN(n8756) );
  NAND2_X1 U8383 ( .A1(n8756), .A2(n6615), .ZN(n6607) );
  INV_X1 U8384 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8757) );
  OR2_X1 U8385 ( .A1(n5781), .A2(n8757), .ZN(n6606) );
  OAI22_X1 U8386 ( .A1(n6611), .A2(n6610), .B1(SI_30_), .B2(n6609), .ZN(n6614)
         );
  INV_X1 U8387 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6677) );
  INV_X1 U8388 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6616) );
  MUX2_X1 U8389 ( .A(n6677), .B(n6616), .S(n7193), .Z(n6612) );
  XNOR2_X1 U8390 ( .A(n6612), .B(SI_31_), .ZN(n6613) );
  XNOR2_X1 U8391 ( .A(n6614), .B(n6613), .ZN(n6676) );
  NAND2_X1 U8392 ( .A1(n6676), .A2(n6615), .ZN(n6618) );
  OR2_X1 U8393 ( .A1(n5781), .A2(n6616), .ZN(n6617) );
  XNOR2_X1 U8394 ( .A(n6619), .B(n8519), .ZN(n9751) );
  NAND2_X1 U8395 ( .A1(n6620), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U8396 ( .A1(n6621), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8397 ( .A1(n5410), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6622) );
  AND3_X1 U8398 ( .A1(n6624), .A2(n6623), .A3(n6622), .ZN(n8664) );
  NOR2_X1 U8399 ( .A1(n8664), .A2(n6625), .ZN(n9752) );
  AOI21_X1 U8400 ( .B1(n9751), .B2(n9992), .A(n9752), .ZN(n6629) );
  NAND2_X1 U8401 ( .A1(n6626), .A2(n5101), .ZN(P1_U3553) );
  INV_X1 U8402 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U8403 ( .A1(n6631), .A2(n5102), .ZN(P1_U3521) );
  INV_X1 U8404 ( .A(n10198), .ZN(n6632) );
  NAND2_X1 U8405 ( .A1(n10198), .A2(n9338), .ZN(n6727) );
  NAND2_X1 U8406 ( .A1(n6699), .A2(n7573), .ZN(n7575) );
  NAND2_X1 U8407 ( .A1(n7575), .A2(n6728), .ZN(n10195) );
  INV_X1 U8408 ( .A(n10204), .ZN(n10216) );
  NAND2_X1 U8409 ( .A1(n7397), .A2(n10216), .ZN(n6734) );
  NAND2_X1 U8410 ( .A1(n7579), .A2(n10204), .ZN(n6735) );
  NAND2_X1 U8411 ( .A1(n6734), .A2(n6735), .ZN(n10197) );
  INV_X1 U8412 ( .A(n10197), .ZN(n6730) );
  NAND2_X1 U8413 ( .A1(n10195), .A2(n6730), .ZN(n6634) );
  NAND2_X1 U8414 ( .A1(n6634), .A2(n6735), .ZN(n7544) );
  NAND2_X2 U8415 ( .A1(n7387), .A2(n7548), .ZN(n7616) );
  INV_X1 U8416 ( .A(n6890), .ZN(n7615) );
  NAND2_X1 U8417 ( .A1(n8875), .A2(n10231), .ZN(n6751) );
  AND2_X1 U8418 ( .A1(n7615), .A2(n6741), .ZN(n6637) );
  INV_X1 U8419 ( .A(n6741), .ZN(n6635) );
  INV_X1 U8420 ( .A(n6700), .ZN(n6748) );
  NOR2_X1 U8421 ( .A1(n6635), .A2(n7701), .ZN(n6636) );
  NAND2_X1 U8422 ( .A1(n7610), .A2(n7891), .ZN(n7747) );
  INV_X1 U8423 ( .A(n10231), .ZN(n6638) );
  NAND2_X1 U8424 ( .A1(n7517), .A2(n6638), .ZN(n7878) );
  NAND2_X1 U8425 ( .A1(n7747), .A2(n7878), .ZN(n6743) );
  NAND2_X1 U8426 ( .A1(n8009), .A2(n7838), .ZN(n6761) );
  INV_X1 U8427 ( .A(n6761), .ZN(n6639) );
  NOR2_X1 U8428 ( .A1(n6743), .A2(n6639), .ZN(n6640) );
  NAND2_X1 U8429 ( .A1(n7744), .A2(n6640), .ZN(n6643) );
  INV_X1 U8430 ( .A(n8013), .ZN(n8017) );
  NAND2_X1 U8431 ( .A1(n8017), .A2(n8872), .ZN(n6766) );
  AND2_X1 U8432 ( .A1(n8874), .A2(n10240), .ZN(n6744) );
  NAND2_X1 U8433 ( .A1(n6761), .A2(n6744), .ZN(n6641) );
  INV_X1 U8434 ( .A(n8009), .ZN(n8873) );
  INV_X1 U8435 ( .A(n7838), .ZN(n7845) );
  NAND2_X1 U8436 ( .A1(n8873), .A2(n7845), .ZN(n7869) );
  AND3_X1 U8437 ( .A1(n6766), .A2(n6641), .A3(n7869), .ZN(n6642) );
  AOI21_X1 U8438 ( .B1(n6643), .B2(n6642), .A(n6698), .ZN(n8106) );
  NAND2_X1 U8439 ( .A1(n8109), .A2(n8096), .ZN(n6763) );
  NAND2_X1 U8440 ( .A1(n8106), .A2(n8111), .ZN(n8108) );
  OR2_X1 U8441 ( .A1(n8091), .A2(n8056), .ZN(n6776) );
  AND2_X1 U8442 ( .A1(n6776), .A2(n8092), .ZN(n6767) );
  NAND2_X1 U8443 ( .A1(n8108), .A2(n6767), .ZN(n6644) );
  NAND2_X1 U8444 ( .A1(n8091), .A2(n8056), .ZN(n6774) );
  NAND2_X1 U8445 ( .A1(n8188), .A2(n9258), .ZN(n6775) );
  XNOR2_X1 U8446 ( .A(n9328), .B(n8284), .ZN(n9255) );
  OR2_X1 U8447 ( .A1(n9328), .A2(n8284), .ZN(n6786) );
  NAND2_X1 U8448 ( .A1(n9249), .A2(n6786), .ZN(n9233) );
  NAND2_X1 U8449 ( .A1(n9428), .A2(n9260), .ZN(n6645) );
  OR2_X1 U8450 ( .A1(n9428), .A2(n9260), .ZN(n6646) );
  INV_X1 U8451 ( .A(n9423), .ZN(n9228) );
  AND2_X1 U8452 ( .A1(n9228), .A2(n9238), .ZN(n6797) );
  NAND2_X1 U8453 ( .A1(n9423), .A2(n9213), .ZN(n6799) );
  AND2_X1 U8454 ( .A1(n9417), .A2(n6804), .ZN(n6803) );
  OR2_X1 U8455 ( .A1(n9417), .A2(n6804), .ZN(n6647) );
  NAND2_X1 U8456 ( .A1(n8794), .A2(n9214), .ZN(n6809) );
  INV_X1 U8457 ( .A(n6808), .ZN(n6648) );
  AOI21_X1 U8458 ( .B1(n9200), .B2(n6809), .A(n6648), .ZN(n9177) );
  OR2_X1 U8459 ( .A1(n9406), .A2(n9199), .ZN(n6693) );
  NAND2_X1 U8460 ( .A1(n9406), .A2(n9199), .ZN(n6695) );
  NAND2_X1 U8461 ( .A1(n6693), .A2(n6695), .ZN(n9183) );
  INV_X1 U8462 ( .A(n9183), .ZN(n9176) );
  NAND2_X1 U8463 ( .A1(n9177), .A2(n9176), .ZN(n9179) );
  NAND2_X1 U8464 ( .A1(n9302), .A2(n9135), .ZN(n6820) );
  NAND2_X1 U8465 ( .A1(n9170), .A2(n9152), .ZN(n9145) );
  NAND2_X1 U8466 ( .A1(n6820), .A2(n9145), .ZN(n6814) );
  OR2_X1 U8467 ( .A1(n8823), .A2(n9153), .ZN(n9117) );
  NAND2_X1 U8468 ( .A1(n6820), .A2(n9147), .ZN(n6650) );
  OR2_X1 U8469 ( .A1(n9302), .A2(n9135), .ZN(n6817) );
  AND2_X1 U8470 ( .A1(n6650), .A2(n6817), .ZN(n9115) );
  NAND2_X1 U8471 ( .A1(n9392), .A2(n9136), .ZN(n6827) );
  NAND2_X1 U8472 ( .A1(n8823), .A2(n9153), .ZN(n9118) );
  AND2_X1 U8473 ( .A1(n6827), .A2(n9118), .ZN(n6823) );
  NAND2_X1 U8474 ( .A1(n9386), .A2(n8782), .ZN(n6722) );
  NAND2_X1 U8475 ( .A1(n9375), .A2(n8790), .ZN(n6838) );
  NAND2_X1 U8476 ( .A1(n9380), .A2(n8817), .ZN(n9079) );
  AND2_X1 U8477 ( .A1(n6838), .A2(n9079), .ZN(n6833) );
  NAND2_X1 U8478 ( .A1(n6652), .A2(n6835), .ZN(n9073) );
  INV_X1 U8479 ( .A(n6839), .ZN(n6653) );
  NAND2_X1 U8480 ( .A1(n9370), .A2(n8849), .ZN(n6840) );
  NAND2_X1 U8481 ( .A1(n9358), .A2(n8723), .ZN(n6849) );
  OR2_X1 U8482 ( .A1(n8712), .A2(n9352), .ZN(n6656) );
  INV_X1 U8483 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9448) );
  OR2_X1 U8484 ( .A1(n6678), .A2(n9448), .ZN(n6658) );
  INV_X1 U8485 ( .A(n8705), .ZN(n6660) );
  NAND2_X1 U8486 ( .A1(n6660), .A2(n6659), .ZN(n6687) );
  INV_X1 U8487 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10453) );
  NAND2_X1 U8488 ( .A1(n6122), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U8489 ( .A1(n6681), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6661) );
  OAI211_X1 U8490 ( .C1(n6667), .C2(n10453), .A(n6662), .B(n6661), .ZN(n6663)
         );
  INV_X1 U8491 ( .A(n6663), .ZN(n6664) );
  INV_X1 U8492 ( .A(n6866), .ZN(n6674) );
  NAND2_X1 U8493 ( .A1(n8756), .A2(n6675), .ZN(n6666) );
  INV_X1 U8494 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9445) );
  OR2_X1 U8495 ( .A1(n6678), .A2(n9445), .ZN(n6665) );
  INV_X1 U8496 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U8497 ( .A1(n6681), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6669) );
  INV_X1 U8498 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10392) );
  OR2_X1 U8499 ( .A1(n6667), .A2(n10392), .ZN(n6668) );
  OAI211_X1 U8500 ( .C1(n6670), .C2(n10458), .A(n6669), .B(n6668), .ZN(n6671)
         );
  INV_X1 U8501 ( .A(n6671), .ZN(n6672) );
  NAND2_X1 U8502 ( .A1(n6687), .A2(n6672), .ZN(n8868) );
  INV_X1 U8503 ( .A(n8868), .ZN(n6673) );
  NAND2_X1 U8504 ( .A1(n9347), .A2(n6673), .ZN(n6861) );
  NAND2_X1 U8505 ( .A1(n6964), .A2(n8719), .ZN(n6692) );
  AND2_X1 U8506 ( .A1(n6861), .A2(n6692), .ZN(n6855) );
  OAI21_X1 U8507 ( .B1(n6930), .B2(n6674), .A(n6855), .ZN(n6688) );
  NAND2_X1 U8508 ( .A1(n6676), .A2(n6675), .ZN(n6680) );
  OR2_X1 U8509 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  NAND2_X1 U8510 ( .A1(n6680), .A2(n6679), .ZN(n6691) );
  NAND2_X1 U8511 ( .A1(n6681), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U8512 ( .A1(n6122), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8513 ( .A1(n6682), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6683) );
  AND3_X1 U8514 ( .A1(n6685), .A2(n6684), .A3(n6683), .ZN(n6686) );
  NAND2_X1 U8515 ( .A1(n6691), .A2(n6689), .ZN(n6867) );
  INV_X1 U8516 ( .A(n9347), .ZN(n9035) );
  AND2_X1 U8517 ( .A1(n9035), .A2(n8868), .ZN(n6863) );
  INV_X1 U8518 ( .A(n6691), .ZN(n9346) );
  NAND2_X1 U8519 ( .A1(n6866), .A2(n6692), .ZN(n6929) );
  XNOR2_X1 U8520 ( .A(n8714), .B(n8712), .ZN(n9037) );
  INV_X1 U8521 ( .A(n9079), .ZN(n6836) );
  NOR2_X1 U8522 ( .A1(n6834), .A2(n6836), .ZN(n9093) );
  INV_X1 U8523 ( .A(n9103), .ZN(n9104) );
  NAND2_X1 U8524 ( .A1(n6828), .A2(n6827), .ZN(n9121) );
  NAND2_X1 U8525 ( .A1(n9117), .A2(n9118), .ZN(n9139) );
  NAND2_X1 U8526 ( .A1(n6817), .A2(n6820), .ZN(n9149) );
  INV_X1 U8527 ( .A(n9149), .ZN(n6708) );
  INV_X1 U8528 ( .A(n6693), .ZN(n6694) );
  NOR2_X1 U8529 ( .A1(n9147), .A2(n6694), .ZN(n6723) );
  NAND2_X1 U8530 ( .A1(n9145), .A2(n6695), .ZN(n6818) );
  XNOR2_X1 U8531 ( .A(n9417), .B(n6804), .ZN(n9210) );
  NAND2_X1 U8532 ( .A1(n6808), .A2(n6809), .ZN(n9201) );
  INV_X1 U8533 ( .A(n6799), .ZN(n6696) );
  INV_X2 U8534 ( .A(n9223), .ZN(n9221) );
  INV_X1 U8535 ( .A(n6697), .ZN(n8178) );
  XNOR2_X1 U8536 ( .A(n8091), .B(n8056), .ZN(n8094) );
  INV_X1 U8537 ( .A(n6744), .ZN(n6754) );
  NAND2_X1 U8538 ( .A1(n6761), .A2(n7869), .ZN(n7749) );
  NAND2_X1 U8539 ( .A1(n7878), .A2(n6751), .ZN(n7706) );
  AND2_X1 U8540 ( .A1(n8878), .A2(n7537), .ZN(n6725) );
  NAND4_X1 U8541 ( .A1(n6699), .A2(n7615), .A3(n6730), .A4(n7351), .ZN(n6702)
         );
  INV_X1 U8542 ( .A(n7703), .ZN(n6701) );
  NAND4_X1 U8543 ( .A1(n8111), .A2(n7873), .A3(n7885), .A4(n6703), .ZN(n6704)
         );
  XNOR2_X1 U8544 ( .A(n9428), .B(n9225), .ZN(n9234) );
  NAND3_X1 U8545 ( .A1(n9221), .A2(n6705), .A3(n9234), .ZN(n6706) );
  NAND3_X1 U8546 ( .A1(n6708), .A2(n6723), .A3(n6707), .ZN(n6709) );
  NAND4_X1 U8547 ( .A1(n9074), .A2(n9082), .A3(n9093), .A4(n6710), .ZN(n6711)
         );
  INV_X1 U8548 ( .A(n6867), .ZN(n6713) );
  NAND2_X1 U8549 ( .A1(n6715), .A2(n7912), .ZN(n6716) );
  NAND2_X1 U8550 ( .A1(n6718), .A2(n5117), .ZN(n6881) );
  INV_X1 U8551 ( .A(n6719), .ZN(n6720) );
  NOR2_X1 U8552 ( .A1(n6834), .A2(n6720), .ZN(n6721) );
  MUX2_X1 U8553 ( .A(n6722), .B(n6721), .S(n9053), .Z(n6832) );
  INV_X1 U8554 ( .A(n9118), .ZN(n6826) );
  INV_X1 U8555 ( .A(n6723), .ZN(n6724) );
  NAND2_X1 U8556 ( .A1(n6724), .A2(n6984), .ZN(n6813) );
  INV_X1 U8557 ( .A(n6725), .ZN(n6729) );
  AND2_X1 U8558 ( .A1(n6729), .A2(n8024), .ZN(n6726) );
  NAND2_X1 U8559 ( .A1(n6699), .A2(n6729), .ZN(n6731) );
  OAI21_X1 U8560 ( .B1(n6732), .B2(n6731), .A(n6730), .ZN(n6733) );
  NAND2_X1 U8561 ( .A1(n6747), .A2(n6734), .ZN(n6737) );
  NAND2_X1 U8562 ( .A1(n7616), .A2(n6735), .ZN(n6736) );
  MUX2_X1 U8563 ( .A(n6737), .B(n6736), .S(n6984), .Z(n6739) );
  INV_X1 U8564 ( .A(n7618), .ZN(n6738) );
  OAI21_X1 U8565 ( .B1(n6740), .B2(n6739), .A(n6738), .ZN(n6750) );
  INV_X1 U8566 ( .A(n7616), .ZN(n6742) );
  OAI21_X1 U8567 ( .B1(n6750), .B2(n6742), .A(n6741), .ZN(n6746) );
  INV_X1 U8568 ( .A(n6743), .ZN(n6745) );
  AOI21_X1 U8569 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(n6756) );
  INV_X1 U8570 ( .A(n6747), .ZN(n6749) );
  OAI211_X1 U8571 ( .C1(n6750), .C2(n6749), .A(n7878), .B(n6748), .ZN(n6752)
         );
  NAND2_X1 U8572 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  NAND2_X1 U8573 ( .A1(n6753), .A2(n7747), .ZN(n6755) );
  INV_X1 U8574 ( .A(n6766), .ZN(n6758) );
  MUX2_X1 U8575 ( .A(n6758), .B(n6757), .S(n6984), .Z(n6760) );
  INV_X1 U8576 ( .A(n8092), .ZN(n6759) );
  INV_X1 U8577 ( .A(n7749), .ZN(n7742) );
  NAND2_X1 U8578 ( .A1(n6762), .A2(n6761), .ZN(n6765) );
  NAND2_X1 U8579 ( .A1(n6774), .A2(n6763), .ZN(n6764) );
  AOI21_X1 U8580 ( .B1(n6770), .B2(n6765), .A(n6764), .ZN(n6772) );
  NAND2_X1 U8581 ( .A1(n6766), .A2(n7869), .ZN(n6769) );
  INV_X1 U8582 ( .A(n6767), .ZN(n6768) );
  AOI21_X1 U8583 ( .B1(n6770), .B2(n6769), .A(n6768), .ZN(n6771) );
  NAND2_X1 U8584 ( .A1(n9328), .A2(n8284), .ZN(n6787) );
  NAND4_X1 U8585 ( .A1(n6787), .A2(n6775), .A3(n6774), .A4(n6984), .ZN(n6780)
         );
  OAI211_X1 U8586 ( .C1(n8188), .C2(n9258), .A(n9053), .B(n6776), .ZN(n6777)
         );
  INV_X1 U8587 ( .A(n6777), .ZN(n6778) );
  NAND2_X1 U8588 ( .A1(n6786), .A2(n6778), .ZN(n6779) );
  NAND2_X1 U8589 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  NAND3_X1 U8590 ( .A1(n6782), .A2(n9234), .A3(n6781), .ZN(n6796) );
  NAND2_X1 U8591 ( .A1(n6786), .A2(n9053), .ZN(n6784) );
  NAND2_X1 U8592 ( .A1(n6787), .A2(n6984), .ZN(n6783) );
  NAND2_X1 U8593 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  NAND2_X1 U8594 ( .A1(n6785), .A2(n9255), .ZN(n6790) );
  NAND4_X1 U8595 ( .A1(n6786), .A2(n9258), .A3(n9053), .A4(n8188), .ZN(n6789)
         );
  INV_X1 U8596 ( .A(n8188), .ZN(n8217) );
  NAND4_X1 U8597 ( .A1(n6787), .A2(n8217), .A3(n6984), .A4(n8869), .ZN(n6788)
         );
  NAND3_X1 U8598 ( .A1(n6790), .A2(n6789), .A3(n6788), .ZN(n6791) );
  NAND2_X1 U8599 ( .A1(n9234), .A2(n6791), .ZN(n6795) );
  NAND2_X1 U8600 ( .A1(n9428), .A2(n9053), .ZN(n6793) );
  OR2_X1 U8601 ( .A1(n9428), .A2(n9053), .ZN(n6792) );
  MUX2_X1 U8602 ( .A(n6793), .B(n6792), .S(n9225), .Z(n6794) );
  NAND4_X1 U8603 ( .A1(n6796), .A2(n9221), .A3(n6795), .A4(n6794), .ZN(n6801)
         );
  INV_X1 U8604 ( .A(n9210), .ZN(n9211) );
  INV_X1 U8605 ( .A(n6797), .ZN(n6798) );
  MUX2_X1 U8606 ( .A(n6799), .B(n6798), .S(n9053), .Z(n6800) );
  NAND2_X1 U8607 ( .A1(n6808), .A2(n6984), .ZN(n6802) );
  OAI21_X1 U8608 ( .B1(n9201), .B2(n6803), .A(n6802), .ZN(n6806) );
  OR3_X1 U8609 ( .A1(n9417), .A2(n6804), .A3(n9053), .ZN(n6805) );
  NAND3_X1 U8610 ( .A1(n6807), .A2(n6806), .A3(n6805), .ZN(n6811) );
  MUX2_X1 U8611 ( .A(n6809), .B(n6808), .S(n9053), .Z(n6810) );
  NAND3_X1 U8612 ( .A1(n6811), .A2(n9176), .A3(n6810), .ZN(n6812) );
  NAND2_X1 U8613 ( .A1(n6819), .A2(n6649), .ZN(n6815) );
  NAND3_X1 U8614 ( .A1(n6815), .A2(n9117), .A3(n6817), .ZN(n6821) );
  INV_X1 U8615 ( .A(n9147), .ZN(n6816) );
  AND2_X1 U8616 ( .A1(n6828), .A2(n9117), .ZN(n6822) );
  MUX2_X1 U8617 ( .A(n6823), .B(n6822), .S(n9053), .Z(n6824) );
  OAI21_X1 U8618 ( .B1(n6826), .B2(n6825), .A(n6824), .ZN(n6830) );
  MUX2_X1 U8619 ( .A(n6828), .B(n6827), .S(n9053), .Z(n6829) );
  NAND3_X1 U8620 ( .A1(n6830), .A2(n9103), .A3(n6829), .ZN(n6831) );
  NAND2_X1 U8621 ( .A1(n6832), .A2(n6831), .ZN(n6837) );
  MUX2_X1 U8622 ( .A(n6840), .B(n6839), .S(n9053), .Z(n6841) );
  NAND3_X1 U8623 ( .A1(n6842), .A2(n4578), .A3(n6841), .ZN(n6847) );
  INV_X1 U8624 ( .A(n6843), .ZN(n6844) );
  MUX2_X1 U8625 ( .A(n6845), .B(n6844), .S(n9053), .Z(n6846) );
  NAND3_X1 U8626 ( .A1(n6847), .A2(n4418), .A3(n6846), .ZN(n6851) );
  MUX2_X1 U8627 ( .A(n6849), .B(n6848), .S(n9053), .Z(n6850) );
  NAND2_X1 U8628 ( .A1(n6851), .A2(n6850), .ZN(n6858) );
  MUX2_X1 U8629 ( .A(n9051), .B(n9352), .S(n6984), .Z(n6856) );
  INV_X1 U8630 ( .A(n6929), .ZN(n6852) );
  INV_X1 U8631 ( .A(n6856), .ZN(n6857) );
  NOR2_X1 U8632 ( .A1(n6929), .A2(n6857), .ZN(n6859) );
  NAND2_X1 U8633 ( .A1(n6859), .A2(n6858), .ZN(n6868) );
  OAI211_X1 U8634 ( .C1(n6870), .C2(n9051), .A(n6860), .B(n6868), .ZN(n6865)
         );
  OAI211_X1 U8635 ( .C1(n6863), .C2(n9053), .A(n6862), .B(n6861), .ZN(n6864)
         );
  AND4_X1 U8636 ( .A1(n6867), .A2(n9053), .A3(n6866), .A4(n6690), .ZN(n6869)
         );
  OAI211_X1 U8637 ( .C1(n6870), .C2(n9352), .A(n6869), .B(n6868), .ZN(n6871)
         );
  INV_X1 U8638 ( .A(n6874), .ZN(n6872) );
  NAND3_X1 U8639 ( .A1(n6872), .A2(n6873), .A3(n7540), .ZN(n6879) );
  NAND4_X1 U8640 ( .A1(n6874), .A2(n6873), .A3(n9017), .A4(n7827), .ZN(n6878)
         );
  NAND3_X1 U8641 ( .A1(n6875), .A2(n7074), .A3(n4410), .ZN(n6876) );
  OAI211_X1 U8642 ( .C1(n6952), .C2(n8063), .A(n6876), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6877) );
  NAND2_X1 U8643 ( .A1(n6881), .A2(n6880), .ZN(P2_U3296) );
  OR2_X1 U8644 ( .A1(n10189), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6882) );
  OAI21_X1 U8645 ( .B1(n10096), .B2(n4993), .A(n6884), .ZN(P1_U3519) );
  NOR2_X1 U8646 ( .A1(n8823), .A2(n9125), .ZN(n9122) );
  NAND2_X1 U8647 ( .A1(n9121), .A2(n9122), .ZN(n6885) );
  INV_X1 U8648 ( .A(n9136), .ZN(n9108) );
  OR2_X1 U8649 ( .A1(n9392), .A2(n9108), .ZN(n9102) );
  NAND2_X1 U8650 ( .A1(n6885), .A2(n9102), .ZN(n9105) );
  NAND2_X1 U8651 ( .A1(n8878), .A2(n7344), .ZN(n7577) );
  NAND2_X1 U8652 ( .A1(n7574), .A2(n7577), .ZN(n6887) );
  NAND2_X1 U8653 ( .A1(n10196), .A2(n10197), .ZN(n6889) );
  NAND2_X1 U8654 ( .A1(n7579), .A2(n10216), .ZN(n6888) );
  NAND2_X1 U8655 ( .A1(n7387), .A2(n10221), .ZN(n6891) );
  NOR2_X1 U8656 ( .A1(n8876), .A2(n7624), .ZN(n6892) );
  NAND2_X1 U8657 ( .A1(n8876), .A2(n7624), .ZN(n6893) );
  NAND2_X1 U8658 ( .A1(n8874), .A2(n7891), .ZN(n6894) );
  NAND2_X1 U8659 ( .A1(n7706), .A2(n6894), .ZN(n6898) );
  NAND2_X1 U8660 ( .A1(n7517), .A2(n10231), .ZN(n6895) );
  NAND2_X1 U8661 ( .A1(n6895), .A2(n8874), .ZN(n6896) );
  INV_X1 U8662 ( .A(n6895), .ZN(n7883) );
  AOI22_X1 U8663 ( .A1(n10240), .A2(n6896), .B1(n7883), .B2(n7610), .ZN(n6897)
         );
  OAI21_X2 U8664 ( .B1(n7708), .B2(n6898), .A(n6897), .ZN(n7743) );
  NAND2_X1 U8665 ( .A1(n8009), .A2(n7845), .ZN(n6899) );
  NAND2_X1 U8666 ( .A1(n8013), .A2(n8872), .ZN(n6900) );
  AND2_X1 U8667 ( .A1(n8109), .A2(n8871), .ZN(n6903) );
  NAND2_X1 U8668 ( .A1(n8091), .A2(n8870), .ZN(n6904) );
  OR2_X1 U8669 ( .A1(n8091), .A2(n8870), .ZN(n8177) );
  OR2_X1 U8670 ( .A1(n8188), .A2(n8869), .ZN(n6905) );
  AND2_X1 U8671 ( .A1(n6905), .A2(n8177), .ZN(n9251) );
  NOR2_X1 U8672 ( .A1(n9328), .A2(n9237), .ZN(n6907) );
  INV_X1 U8673 ( .A(n6907), .ZN(n6906) );
  AND2_X1 U8674 ( .A1(n6906), .A2(n9251), .ZN(n6908) );
  NAND2_X1 U8675 ( .A1(n8188), .A2(n8869), .ZN(n9253) );
  AND2_X1 U8676 ( .A1(n9428), .A2(n9225), .ZN(n6909) );
  NOR2_X1 U8677 ( .A1(n9423), .A2(n9238), .ZN(n6911) );
  NAND2_X1 U8678 ( .A1(n9423), .A2(n9238), .ZN(n6910) );
  AND2_X1 U8679 ( .A1(n9417), .A2(n9226), .ZN(n9180) );
  AND2_X1 U8680 ( .A1(n8794), .A2(n6269), .ZN(n9184) );
  AOI22_X1 U8681 ( .A1(n9183), .A2(n9184), .B1(n9406), .B2(n9163), .ZN(n6912)
         );
  INV_X1 U8682 ( .A(n6912), .ZN(n6913) );
  OR2_X1 U8683 ( .A1(n9180), .A2(n6913), .ZN(n9159) );
  AND2_X1 U8684 ( .A1(n9170), .A2(n9187), .ZN(n6915) );
  OR2_X1 U8685 ( .A1(n9170), .A2(n9187), .ZN(n6914) );
  OR2_X1 U8686 ( .A1(n9417), .A2(n9226), .ZN(n9181) );
  OR2_X1 U8687 ( .A1(n6913), .A2(n4493), .ZN(n9160) );
  AND2_X1 U8688 ( .A1(n9302), .A2(n9164), .ZN(n6916) );
  NOR2_X1 U8689 ( .A1(n6917), .A2(n8817), .ZN(n6918) );
  NOR2_X1 U8690 ( .A1(n9375), .A2(n9095), .ZN(n6919) );
  INV_X1 U8691 ( .A(n9375), .ZN(n9087) );
  NAND2_X1 U8692 ( .A1(n9364), .A2(n9069), .ZN(n6921) );
  NAND2_X1 U8693 ( .A1(n9049), .A2(n6922), .ZN(n6923) );
  NOR2_X1 U8694 ( .A1(n8714), .A2(n8712), .ZN(n6925) );
  NAND2_X2 U8695 ( .A1(n6928), .A2(n6927), .ZN(n10202) );
  XNOR2_X1 U8696 ( .A(n6930), .B(n6929), .ZN(n8709) );
  NAND2_X1 U8697 ( .A1(n8024), .A2(n6953), .ZN(n6931) );
  AND3_X1 U8698 ( .A1(n9017), .A2(n6931), .A3(n10239), .ZN(n6932) );
  NAND2_X1 U8699 ( .A1(n8709), .A2(n8098), .ZN(n6935) );
  NOR2_X1 U8700 ( .A1(n9261), .A2(n4522), .ZN(n9029) );
  AOI22_X1 U8701 ( .A1(n9236), .A2(n9051), .B1(n8868), .B2(n9029), .ZN(n6934)
         );
  NAND2_X1 U8702 ( .A1(n7540), .A2(n8024), .ZN(n9334) );
  NAND2_X1 U8703 ( .A1(n6937), .A2(n7522), .ZN(n6938) );
  NAND2_X1 U8704 ( .A1(n6939), .A2(n6938), .ZN(n6943) );
  NAND2_X1 U8705 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  NAND2_X1 U8706 ( .A1(n10247), .A2(n10453), .ZN(n6944) );
  NAND2_X1 U8707 ( .A1(n6945), .A2(n6944), .ZN(n6948) );
  NAND2_X1 U8708 ( .A1(n6948), .A2(n6947), .ZN(P2_U3456) );
  NAND3_X1 U8709 ( .A1(n9017), .A2(n6953), .A3(n6952), .ZN(n6954) );
  OAI21_X1 U8710 ( .B1(n7526), .B2(n6955), .A(n7529), .ZN(n6958) );
  INV_X1 U8711 ( .A(n7529), .ZN(n6956) );
  NAND2_X1 U8712 ( .A1(n6956), .A2(n7528), .ZN(n6957) );
  NAND2_X1 U8713 ( .A1(n9273), .A2(n6960), .ZN(n6961) );
  NAND2_X1 U8714 ( .A1(n6962), .A2(n6961), .ZN(n6966) );
  NAND2_X1 U8715 ( .A1(n6966), .A2(n6965), .ZN(P2_U3488) );
  NAND2_X1 U8716 ( .A1(n6967), .A2(n8561), .ZN(n6969) );
  NAND3_X1 U8717 ( .A1(n6972), .A2(n6971), .A3(n9964), .ZN(n6975) );
  NAND2_X1 U8718 ( .A1(n9607), .A2(n9567), .ZN(n6974) );
  NAND2_X1 U8719 ( .A1(n9609), .A2(n9595), .ZN(n6973) );
  AND2_X1 U8720 ( .A1(n6974), .A2(n6973), .ZN(n8747) );
  MUX2_X1 U8721 ( .A(n10473), .B(n6979), .S(n10189), .Z(n6978) );
  INV_X1 U8722 ( .A(n9767), .ZN(n6981) );
  NAND2_X1 U8723 ( .A1(n6978), .A2(n5107), .ZN(P1_U3518) );
  INV_X1 U8724 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8725 ( .A(n6980), .B(n6979), .S(n10194), .Z(n6982) );
  NAND2_X1 U8726 ( .A1(n6982), .A2(n5104), .ZN(P1_U3550) );
  NAND2_X1 U8727 ( .A1(n6984), .A2(n7070), .ZN(n6985) );
  NAND2_X1 U8728 ( .A1(n6985), .A2(n7068), .ZN(n7073) );
  NAND2_X1 U8729 ( .A1(n6986), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U8730 ( .A1(n8764), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6987) );
  OAI21_X1 U8731 ( .B1(n7186), .B2(n6987), .A(n6989), .ZN(n6988) );
  INV_X1 U8732 ( .A(n6988), .ZN(n7315) );
  NAND2_X1 U8733 ( .A1(n7315), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U8734 ( .A1(n7314), .A2(n6989), .ZN(n8888) );
  XNOR2_X1 U8735 ( .A(n7169), .B(n10248), .ZN(n8889) );
  NAND2_X1 U8736 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  NAND2_X1 U8737 ( .A1(n7169), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8738 ( .A1(n7330), .A2(n7282), .ZN(n6991) );
  XNOR2_X1 U8739 ( .A(n7297), .B(n10252), .ZN(n7281) );
  NAND2_X1 U8740 ( .A1(n7297), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U8741 ( .A1(n7285), .A2(n6992), .ZN(n6995) );
  INV_X1 U8742 ( .A(n6995), .ZN(n6994) );
  INV_X1 U8743 ( .A(n7305), .ZN(n6993) );
  NAND2_X1 U8744 ( .A1(n6995), .A2(n7305), .ZN(n7374) );
  NAND2_X1 U8745 ( .A1(n7300), .A2(n7374), .ZN(n6997) );
  XNOR2_X1 U8746 ( .A(n7373), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U8747 ( .A1(n6997), .A2(n7375), .ZN(n7378) );
  INV_X1 U8748 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7042) );
  OR2_X1 U8749 ( .A1(n7373), .A2(n7042), .ZN(n6998) );
  NAND2_X1 U8750 ( .A1(n7378), .A2(n6998), .ZN(n6999) );
  NAND2_X1 U8751 ( .A1(n6999), .A2(n7460), .ZN(n7155) );
  NAND2_X1 U8752 ( .A1(n7463), .A2(n7155), .ZN(n7000) );
  XNOR2_X1 U8753 ( .A(n7162), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7154) );
  OR2_X1 U8754 ( .A1(n7162), .A2(n10376), .ZN(n7001) );
  INV_X1 U8755 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7589) );
  XNOR2_X1 U8756 ( .A(n7088), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8757 ( .A1(n7002), .A2(n7003), .ZN(n7082) );
  INV_X1 U8758 ( .A(n7003), .ZN(n7005) );
  NAND3_X1 U8759 ( .A1(n7586), .A2(n7005), .A3(n7004), .ZN(n7006) );
  NOR2_X1 U8760 ( .A1(n6449), .A2(P2_U3151), .ZN(n9450) );
  AOI21_X1 U8761 ( .B1(n7082), .B2(n7006), .A(n8976), .ZN(n7080) );
  AND2_X1 U8762 ( .A1(n8764), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7008) );
  OAI21_X1 U8763 ( .B1(n7186), .B2(n7008), .A(n7010), .ZN(n7009) );
  INV_X1 U8764 ( .A(n7009), .ZN(n7312) );
  NAND2_X1 U8765 ( .A1(n7311), .A2(n7010), .ZN(n8883) );
  NAND2_X1 U8766 ( .A1(n8883), .A2(n8884), .ZN(n8882) );
  NAND2_X1 U8767 ( .A1(n7169), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U8768 ( .A1(n7012), .A2(n7171), .ZN(n7287) );
  NAND2_X1 U8769 ( .A1(n7328), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U8770 ( .A1(n7327), .A2(n7287), .ZN(n7014) );
  INV_X1 U8771 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7621) );
  XNOR2_X1 U8772 ( .A(n7297), .B(n7621), .ZN(n7286) );
  NAND2_X1 U8773 ( .A1(n7368), .A2(n7366), .ZN(n7015) );
  XNOR2_X1 U8774 ( .A(n7373), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7365) );
  NAND2_X1 U8775 ( .A1(n7015), .A2(n7365), .ZN(n7370) );
  INV_X1 U8776 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7888) );
  OR2_X1 U8777 ( .A1(n7373), .A2(n7888), .ZN(n7016) );
  INV_X1 U8778 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7051) );
  OR2_X1 U8779 ( .A1(n7162), .A2(n7051), .ZN(n7019) );
  NAND2_X1 U8780 ( .A1(n7161), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U8781 ( .A1(n7020), .A2(n7202), .ZN(n7022) );
  XNOR2_X1 U8782 ( .A(n7088), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7021) );
  INV_X1 U8783 ( .A(n7021), .ZN(n7023) );
  NAND3_X1 U8784 ( .A1(n7600), .A2(n7023), .A3(n7022), .ZN(n7024) );
  AOI21_X1 U8785 ( .B1(n7090), .B2(n7024), .A(n9027), .ZN(n7079) );
  MUX2_X1 U8786 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n6448), .Z(n7027) );
  XNOR2_X1 U8787 ( .A(n7027), .B(n7320), .ZN(n7310) );
  MUX2_X1 U8788 ( .A(n7026), .B(n7025), .S(n7072), .Z(n8759) );
  NAND2_X1 U8789 ( .A1(n8759), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U8790 ( .A1(n7310), .A2(n8758), .ZN(n7029) );
  NAND2_X1 U8791 ( .A1(n7027), .A2(n7186), .ZN(n7028) );
  NAND2_X1 U8792 ( .A1(n7029), .A2(n7028), .ZN(n8879) );
  MUX2_X1 U8793 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n7072), .Z(n7030) );
  XNOR2_X1 U8794 ( .A(n7030), .B(n4787), .ZN(n8880) );
  NAND2_X1 U8795 ( .A1(n8879), .A2(n8880), .ZN(n7032) );
  NAND2_X1 U8796 ( .A1(n7030), .A2(n7169), .ZN(n7031) );
  NAND2_X1 U8797 ( .A1(n7032), .A2(n7031), .ZN(n7325) );
  MUX2_X1 U8798 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n7072), .Z(n7034) );
  XNOR2_X1 U8799 ( .A(n7034), .B(n7171), .ZN(n7326) );
  MUX2_X1 U8800 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n7072), .Z(n7037) );
  INV_X1 U8801 ( .A(n7297), .ZN(n7033) );
  XNOR2_X1 U8802 ( .A(n7037), .B(n7033), .ZN(n7279) );
  INV_X1 U8803 ( .A(n7034), .ZN(n7035) );
  NAND2_X1 U8804 ( .A1(n7035), .A2(n4537), .ZN(n7277) );
  AND2_X1 U8805 ( .A1(n7279), .A2(n7277), .ZN(n7036) );
  NAND2_X1 U8806 ( .A1(n7323), .A2(n7036), .ZN(n7278) );
  NAND2_X1 U8807 ( .A1(n7037), .A2(n7297), .ZN(n7038) );
  NAND2_X1 U8808 ( .A1(n7278), .A2(n7038), .ZN(n7299) );
  MUX2_X1 U8809 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n7072), .Z(n7039) );
  XNOR2_X1 U8810 ( .A(n7039), .B(n6993), .ZN(n7298) );
  NAND2_X1 U8811 ( .A1(n7299), .A2(n7298), .ZN(n7041) );
  NAND2_X1 U8812 ( .A1(n7039), .A2(n7305), .ZN(n7040) );
  NAND2_X1 U8813 ( .A1(n7041), .A2(n7040), .ZN(n7364) );
  MUX2_X1 U8814 ( .A(n7042), .B(n7888), .S(n7072), .Z(n7043) );
  NAND2_X1 U8815 ( .A1(n7043), .A2(n7373), .ZN(n7451) );
  INV_X1 U8816 ( .A(n7043), .ZN(n7044) );
  INV_X1 U8817 ( .A(n7373), .ZN(n7178) );
  NAND2_X1 U8818 ( .A1(n7044), .A2(n7178), .ZN(n7045) );
  NAND2_X1 U8819 ( .A1(n7451), .A2(n7045), .ZN(n7363) );
  NAND2_X1 U8820 ( .A1(n7456), .A2(n7451), .ZN(n7050) );
  INV_X1 U8821 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7895) );
  MUX2_X1 U8822 ( .A(n7895), .B(n4897), .S(n7072), .Z(n7047) );
  NAND2_X1 U8823 ( .A1(n7047), .A2(n7046), .ZN(n7152) );
  INV_X1 U8824 ( .A(n7047), .ZN(n7048) );
  NAND2_X1 U8825 ( .A1(n7048), .A2(n7460), .ZN(n7049) );
  AND2_X1 U8826 ( .A1(n7152), .A2(n7049), .ZN(n7453) );
  NAND2_X1 U8827 ( .A1(n7050), .A2(n7453), .ZN(n7454) );
  NAND2_X1 U8828 ( .A1(n7454), .A2(n7152), .ZN(n7055) );
  MUX2_X1 U8829 ( .A(n10376), .B(n7051), .S(n7072), .Z(n7052) );
  NAND2_X1 U8830 ( .A1(n7052), .A2(n7162), .ZN(n7591) );
  INV_X1 U8831 ( .A(n7052), .ZN(n7053) );
  INV_X1 U8832 ( .A(n7162), .ZN(n7183) );
  NAND2_X1 U8833 ( .A1(n7053), .A2(n7183), .ZN(n7054) );
  AND2_X1 U8834 ( .A1(n7591), .A2(n7054), .ZN(n7150) );
  NAND2_X1 U8835 ( .A1(n7590), .A2(n7591), .ZN(n7059) );
  MUX2_X1 U8836 ( .A(n7589), .B(n10468), .S(n9009), .Z(n7056) );
  NAND2_X1 U8837 ( .A1(n7056), .A2(n7603), .ZN(n7066) );
  INV_X1 U8838 ( .A(n7056), .ZN(n7057) );
  NAND2_X1 U8839 ( .A1(n7057), .A2(n7202), .ZN(n7058) );
  AND2_X1 U8840 ( .A1(n7066), .A2(n7058), .ZN(n7592) );
  NAND2_X1 U8841 ( .A1(n7059), .A2(n7592), .ZN(n7595) );
  NAND2_X1 U8842 ( .A1(n7595), .A2(n7066), .ZN(n7063) );
  INV_X1 U8843 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8104) );
  INV_X1 U8844 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7087) );
  MUX2_X1 U8845 ( .A(n8104), .B(n7087), .S(n9009), .Z(n7060) );
  NAND2_X1 U8846 ( .A1(n7060), .A2(n7088), .ZN(n7850) );
  INV_X1 U8847 ( .A(n7060), .ZN(n7061) );
  INV_X1 U8848 ( .A(n7088), .ZN(n7226) );
  NAND2_X1 U8849 ( .A1(n7061), .A2(n7226), .ZN(n7062) );
  AND2_X1 U8850 ( .A1(n7850), .A2(n7062), .ZN(n7064) );
  INV_X1 U8851 ( .A(n7064), .ZN(n7065) );
  NAND3_X1 U8852 ( .A1(n7595), .A2(n7066), .A3(n7065), .ZN(n7067) );
  AOI21_X1 U8853 ( .B1(n7855), .B2(n7067), .A(n8150), .ZN(n7078) );
  INV_X1 U8854 ( .A(n7068), .ZN(n7069) );
  NOR2_X1 U8855 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  AND2_X1 U8856 ( .A1(n7072), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9452) );
  NAND2_X1 U8857 ( .A1(n7073), .A2(n9452), .ZN(n7075) );
  MUX2_X1 U8858 ( .A(n7075), .B(n8877), .S(n7074), .Z(n9018) );
  NAND2_X1 U8859 ( .A1(n8991), .A2(n7088), .ZN(n7076) );
  NAND2_X1 U8860 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8085) );
  OAI211_X1 U8861 ( .C1(n10281), .C2(n9020), .A(n7076), .B(n8085), .ZN(n7077)
         );
  OR2_X1 U8862 ( .A1(n7088), .A2(n8104), .ZN(n7081) );
  NAND2_X1 U8863 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  NAND3_X1 U8864 ( .A1(n7863), .A2(n4520), .A3(n7085), .ZN(n7086) );
  AOI21_X1 U8865 ( .B1(n7127), .B2(n7086), .A(n8976), .ZN(n7115) );
  OR2_X1 U8866 ( .A1(n7088), .A2(n7087), .ZN(n7089) );
  XNOR2_X1 U8867 ( .A(n7125), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7093) );
  INV_X1 U8868 ( .A(n7093), .ZN(n7095) );
  NAND3_X1 U8869 ( .A1(n7857), .A2(n7095), .A3(n7094), .ZN(n7096) );
  AOI21_X1 U8870 ( .B1(n7119), .B2(n7096), .A(n9027), .ZN(n7114) );
  NAND2_X1 U8871 ( .A1(n7855), .A2(n7850), .ZN(n7101) );
  INV_X1 U8872 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8186) );
  MUX2_X1 U8873 ( .A(n4811), .B(n8186), .S(n9009), .Z(n7098) );
  NAND2_X1 U8874 ( .A1(n7098), .A2(n7097), .ZN(n7108) );
  INV_X1 U8875 ( .A(n7098), .ZN(n7099) );
  NAND2_X1 U8876 ( .A1(n7099), .A2(n7859), .ZN(n7100) );
  AND2_X1 U8877 ( .A1(n7108), .A2(n7100), .ZN(n7852) );
  NAND2_X1 U8878 ( .A1(n7101), .A2(n7852), .ZN(n7853) );
  NAND2_X1 U8879 ( .A1(n7853), .A2(n7108), .ZN(n7105) );
  INV_X1 U8880 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9330) );
  INV_X1 U8881 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9263) );
  MUX2_X1 U8882 ( .A(n9330), .B(n9263), .S(n9009), .Z(n7102) );
  NAND2_X1 U8883 ( .A1(n7102), .A2(n7125), .ZN(n8148) );
  INV_X1 U8884 ( .A(n7102), .ZN(n7103) );
  INV_X1 U8885 ( .A(n7125), .ZN(n7341) );
  NAND2_X1 U8886 ( .A1(n7103), .A2(n7341), .ZN(n7104) );
  AND2_X1 U8887 ( .A1(n8148), .A2(n7104), .ZN(n7106) );
  NAND2_X1 U8888 ( .A1(n7105), .A2(n7106), .ZN(n8149) );
  INV_X1 U8889 ( .A(n7106), .ZN(n7107) );
  NAND3_X1 U8890 ( .A1(n7853), .A2(n7108), .A3(n7107), .ZN(n7109) );
  AOI21_X1 U8891 ( .B1(n8149), .B2(n7109), .A(n8150), .ZN(n7113) );
  NAND2_X1 U8892 ( .A1(n8978), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U8893 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n7110) );
  OAI211_X1 U8894 ( .C1(n9018), .C2(n7341), .A(n7111), .B(n7110), .ZN(n7112)
         );
  OR4_X1 U8895 ( .A1(n7115), .A2(n7114), .A3(n7113), .A4(n7112), .ZN(P2_U3194)
         );
  INV_X4 U8896 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U8897 ( .A1(n4562), .A2(P1_U3086), .ZN(n7117) );
  OR2_X1 U8898 ( .A1(n7125), .A2(n9263), .ZN(n7118) );
  NAND2_X1 U8899 ( .A1(n7120), .A2(n7348), .ZN(n7123) );
  NAND3_X1 U8900 ( .A1(n7122), .A2(n4515), .A3(n7123), .ZN(n7124) );
  AOI21_X1 U8901 ( .B1(n8897), .B2(n7124), .A(n9027), .ZN(n7149) );
  OR2_X1 U8902 ( .A1(n7125), .A2(n9330), .ZN(n7126) );
  NAND3_X1 U8903 ( .A1(n7129), .A2(n4516), .A3(n7130), .ZN(n7131) );
  AOI21_X1 U8904 ( .B1(n8912), .B2(n7131), .A(n8976), .ZN(n7148) );
  NAND2_X1 U8905 ( .A1(n8149), .A2(n8148), .ZN(n7136) );
  INV_X1 U8906 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9324) );
  INV_X1 U8907 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7132) );
  MUX2_X1 U8908 ( .A(n9324), .B(n7132), .S(n9009), .Z(n7133) );
  NAND2_X1 U8909 ( .A1(n7133), .A2(n8155), .ZN(n7143) );
  INV_X1 U8910 ( .A(n7133), .ZN(n7134) );
  NAND2_X1 U8911 ( .A1(n7134), .A2(n7348), .ZN(n7135) );
  AND2_X1 U8912 ( .A1(n7143), .A2(n7135), .ZN(n8146) );
  NAND2_X1 U8913 ( .A1(n7136), .A2(n8146), .ZN(n8152) );
  NAND2_X1 U8914 ( .A1(n8152), .A2(n7143), .ZN(n7140) );
  INV_X1 U8915 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9321) );
  INV_X1 U8916 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U8917 ( .A(n9321), .B(n8895), .S(n9009), .Z(n7137) );
  NAND2_X1 U8918 ( .A1(n7137), .A2(n8910), .ZN(n8902) );
  INV_X1 U8919 ( .A(n7137), .ZN(n7138) );
  INV_X1 U8920 ( .A(n8910), .ZN(n7355) );
  NAND2_X1 U8921 ( .A1(n7138), .A2(n7355), .ZN(n7139) );
  AND2_X1 U8922 ( .A1(n8902), .A2(n7139), .ZN(n7141) );
  NAND2_X1 U8923 ( .A1(n7140), .A2(n7141), .ZN(n8903) );
  INV_X1 U8924 ( .A(n7141), .ZN(n7142) );
  NAND3_X1 U8925 ( .A1(n8152), .A2(n7143), .A3(n7142), .ZN(n7144) );
  AOI21_X1 U8926 ( .B1(n8903), .B2(n7144), .A(n8150), .ZN(n7147) );
  NOR2_X1 U8927 ( .A1(n4739), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8278) );
  AOI21_X1 U8928 ( .B1(n8978), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n8278), .ZN(
        n7145) );
  OAI21_X1 U8929 ( .B1(n7355), .B2(n9018), .A(n7145), .ZN(n7146) );
  OR4_X1 U8930 ( .A1(n7149), .A2(n7148), .A3(n7147), .A4(n7146), .ZN(P2_U3196)
         );
  INV_X1 U8931 ( .A(n7150), .ZN(n7151) );
  NAND3_X1 U8932 ( .A1(n7454), .A2(n7152), .A3(n7151), .ZN(n7153) );
  AOI21_X1 U8933 ( .B1(n7590), .B2(n7153), .A(n8150), .ZN(n7167) );
  INV_X1 U8934 ( .A(n7154), .ZN(n7156) );
  NAND3_X1 U8935 ( .A1(n7463), .A2(n7156), .A3(n7155), .ZN(n7157) );
  AOI21_X1 U8936 ( .B1(n7158), .B2(n7157), .A(n8976), .ZN(n7166) );
  NAND3_X1 U8937 ( .A1(n7458), .A2(n4514), .A3(n7159), .ZN(n7160) );
  AOI21_X1 U8938 ( .B1(n7161), .B2(n7160), .A(n9027), .ZN(n7165) );
  INV_X1 U8939 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U8940 ( .A1(n8991), .A2(n7162), .ZN(n7163) );
  NAND2_X1 U8941 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8008) );
  OAI211_X1 U8942 ( .C1(n10274), .C2(n9020), .A(n7163), .B(n8008), .ZN(n7164)
         );
  OR4_X1 U8943 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(P2_U3190)
         );
  NAND2_X2 U8944 ( .A1(n7168), .A2(P2_U3151), .ZN(n9455) );
  OAI222_X1 U8945 ( .A1(n9449), .A2(n7170), .B1(n9455), .B2(n7206), .C1(
        P2_U3151), .C2(n7169), .ZN(P2_U3293) );
  OAI222_X1 U8946 ( .A1(n9449), .A2(n7172), .B1(n9455), .B2(n7203), .C1(
        P2_U3151), .C2(n7171), .ZN(P2_U3292) );
  OAI222_X1 U8947 ( .A1(n9449), .A2(n7173), .B1(n9455), .B2(n7210), .C1(
        P2_U3151), .C2(n7305), .ZN(P2_U3290) );
  OAI222_X1 U8948 ( .A1(n9449), .A2(n7174), .B1(n9455), .B2(n6085), .C1(
        P2_U3151), .C2(n7297), .ZN(P2_U3291) );
  INV_X1 U8949 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7176) );
  INV_X1 U8950 ( .A(n7175), .ZN(n7205) );
  OAI222_X1 U8951 ( .A1(n9449), .A2(n7176), .B1(n9455), .B2(n7205), .C1(
        P2_U3151), .C2(n7460), .ZN(P2_U3288) );
  INV_X1 U8952 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7179) );
  INV_X1 U8953 ( .A(n7177), .ZN(n7208) );
  OAI222_X1 U8954 ( .A1(n9449), .A2(n7179), .B1(n9455), .B2(n7208), .C1(
        P2_U3151), .C2(n7178), .ZN(P2_U3289) );
  NAND2_X1 U8955 ( .A1(n7181), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7180) );
  OAI21_X1 U8956 ( .B1(n7528), .B2(n7181), .A(n7180), .ZN(P2_U3377) );
  INV_X1 U8957 ( .A(n7182), .ZN(n7213) );
  OAI222_X1 U8958 ( .A1(n9449), .A2(n7184), .B1(n9455), .B2(n7213), .C1(
        P2_U3151), .C2(n7183), .ZN(P2_U3287) );
  OAI222_X1 U8959 ( .A1(n7186), .A2(P2_U3151), .B1(n9455), .B2(n7222), .C1(
        n7185), .C2(n9449), .ZN(P2_U3294) );
  INV_X1 U8960 ( .A(n7189), .ZN(n7190) );
  AOI22_X1 U8961 ( .A1(n7215), .A2(n7191), .B1(n7342), .B2(n7190), .ZN(
        P2_U3376) );
  INV_X1 U8962 ( .A(n7192), .ZN(n7201) );
  NAND2_X2 U8963 ( .A1(n4411), .A2(P1_U3086), .ZN(n10114) );
  AOI22_X1 U8964 ( .A1(n7479), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10106), .ZN(n7194) );
  OAI21_X1 U8965 ( .B1(n7201), .B2(n10114), .A(n7194), .ZN(P1_U3346) );
  INV_X1 U8966 ( .A(n8567), .ZN(n7198) );
  INV_X1 U8967 ( .A(n7196), .ZN(n7197) );
  AOI22_X1 U8968 ( .A1(n10169), .A2(n7199), .B1(n7198), .B2(n7197), .ZN(
        P1_U3440) );
  AND2_X1 U8969 ( .A1(n7215), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8970 ( .A1(n7215), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8971 ( .A1(n7215), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8972 ( .A1(n7215), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8973 ( .A1(n7215), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8974 ( .A1(n7215), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8975 ( .A1(n7215), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8976 ( .A1(n7215), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8977 ( .A1(n7215), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8978 ( .A1(n7215), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8979 ( .A1(n7215), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8980 ( .A1(n7215), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8981 ( .A1(n7215), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8982 ( .A1(n7215), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8983 ( .A1(n7215), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8984 ( .A1(n7215), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8985 ( .A1(n7215), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8986 ( .A1(n7215), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8987 ( .A1(n7215), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8988 ( .A1(n7215), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8989 ( .A1(n7215), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8990 ( .A1(n7215), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8991 ( .A1(n7215), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8992 ( .A1(n7215), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  OAI222_X1 U8993 ( .A1(P2_U3151), .A2(n7202), .B1(n9455), .B2(n7201), .C1(
        n7200), .C2(n9449), .ZN(P2_U3286) );
  OAI222_X1 U8994 ( .A1(n10115), .A2(n7204), .B1(n10114), .B2(n7203), .C1(
        P1_U3086), .C2(n9644), .ZN(P1_U3352) );
  OAI222_X1 U8995 ( .A1(n10115), .A2(n10321), .B1(n10114), .B2(n7205), .C1(
        P1_U3086), .C2(n7267), .ZN(P1_U3348) );
  OAI222_X1 U8996 ( .A1(n10115), .A2(n7207), .B1(n10114), .B2(n7206), .C1(
        P1_U3086), .C2(n7245), .ZN(P1_U3353) );
  OAI222_X1 U8997 ( .A1(n10115), .A2(n7209), .B1(n10114), .B2(n7208), .C1(
        P1_U3086), .C2(n9669), .ZN(P1_U3349) );
  OAI222_X1 U8998 ( .A1(n10115), .A2(n7211), .B1(n10114), .B2(n7210), .C1(
        P1_U3086), .C2(n9661), .ZN(P1_U3350) );
  OAI222_X1 U8999 ( .A1(n10115), .A2(n7212), .B1(n10114), .B2(n6085), .C1(
        P1_U3086), .C2(n7250), .ZN(P1_U3351) );
  INV_X1 U9000 ( .A(n7418), .ZN(n7413) );
  OAI222_X1 U9001 ( .A1(n10115), .A2(n7214), .B1(n10114), .B2(n7213), .C1(
        P1_U3086), .C2(n7413), .ZN(P1_U3347) );
  INV_X1 U9002 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U9003 ( .A1(n7216), .A2(n10554), .ZN(P2_U3239) );
  INV_X1 U9004 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10608) );
  NOR2_X1 U9005 ( .A1(n7216), .A2(n10608), .ZN(P2_U3245) );
  INV_X1 U9006 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10447) );
  NOR2_X1 U9007 ( .A1(n7216), .A2(n10447), .ZN(P2_U3240) );
  INV_X1 U9008 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10536) );
  NOR2_X1 U9009 ( .A1(n7216), .A2(n10536), .ZN(P2_U3243) );
  INV_X1 U9010 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10524) );
  NOR2_X1 U9011 ( .A1(n7216), .A2(n10524), .ZN(P2_U3255) );
  INV_X1 U9012 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10423) );
  NOR2_X1 U9013 ( .A1(n7216), .A2(n10423), .ZN(P2_U3247) );
  NAND2_X1 U9014 ( .A1(n8671), .A2(n7219), .ZN(n7218) );
  AND2_X1 U9015 ( .A1(n7218), .A2(n7217), .ZN(n7240) );
  INV_X1 U9016 ( .A(n7240), .ZN(n7220) );
  NAND2_X1 U9017 ( .A1(n8570), .A2(n8567), .ZN(n7239) );
  NOR2_X1 U9018 ( .A1(n10122), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U9019 ( .A(n9636), .ZN(n7223) );
  OAI222_X1 U9020 ( .A1(n7223), .A2(P1_U3086), .B1(n10114), .B2(n7222), .C1(
        n7221), .C2(n10115), .ZN(P1_U3354) );
  INV_X1 U9021 ( .A(n7224), .ZN(n7228) );
  OAI222_X1 U9022 ( .A1(P2_U3151), .A2(n7226), .B1(n9455), .B2(n7228), .C1(
        n7225), .C2(n9449), .ZN(P2_U3285) );
  INV_X1 U9023 ( .A(n7422), .ZN(n7439) );
  OAI222_X1 U9024 ( .A1(P1_U3086), .A2(n7439), .B1(n10114), .B2(n7228), .C1(
        n7227), .C2(n10115), .ZN(P1_U3345) );
  INV_X1 U9025 ( .A(n8664), .ZN(n8669) );
  NAND2_X1 U9026 ( .A1(n8669), .A2(P1_U3973), .ZN(n7229) );
  OAI21_X1 U9027 ( .B1(P1_U3973), .B2(n6677), .A(n7229), .ZN(P1_U3585) );
  INV_X1 U9028 ( .A(n7230), .ZN(n7232) );
  OAI222_X1 U9029 ( .A1(n9449), .A2(n7231), .B1(n9455), .B2(n7232), .C1(
        P2_U3151), .C2(n7859), .ZN(P2_U3284) );
  OAI222_X1 U9030 ( .A1(n10115), .A2(n7233), .B1(n10114), .B2(n7232), .C1(
        P1_U3086), .C2(n7554), .ZN(P1_U3344) );
  INV_X1 U9031 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10454) );
  NOR2_X1 U9032 ( .A1(n7267), .A2(n10454), .ZN(n7238) );
  INV_X1 U9033 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U9034 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9634) );
  NOR2_X1 U9035 ( .A1(n9633), .A2(n9634), .ZN(n9632) );
  INV_X1 U9036 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10534) );
  MUX2_X1 U9037 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10534), .S(n7245), .Z(n7497)
         );
  OAI22_X1 U9038 ( .A1(n7498), .A2(n7497), .B1(n10534), .B2(n7245), .ZN(n9649)
         );
  INV_X1 U9039 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7234) );
  MUX2_X1 U9040 ( .A(n7234), .B(P1_REG1_REG_3__SCAN_IN), .S(n9644), .Z(n9650)
         );
  NAND2_X1 U9041 ( .A1(n9649), .A2(n9650), .ZN(n10125) );
  INV_X1 U9042 ( .A(n9644), .ZN(n7235) );
  NAND2_X1 U9043 ( .A1(n7235), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10124) );
  INV_X1 U9044 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10574) );
  MUX2_X1 U9045 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10574), .S(n7250), .Z(n10123) );
  NOR2_X1 U9046 ( .A1(n7250), .A2(n10574), .ZN(n9662) );
  INV_X1 U9047 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7236) );
  MUX2_X1 U9048 ( .A(n7236), .B(P1_REG1_REG_5__SCAN_IN), .S(n9661), .Z(n7237)
         );
  INV_X1 U9049 ( .A(n9661), .ZN(n9657) );
  NAND2_X1 U9050 ( .A1(n9657), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9677) );
  INV_X1 U9051 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10422) );
  MUX2_X1 U9052 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10422), .S(n9669), .Z(n9676)
         );
  NOR2_X1 U9053 ( .A1(n9669), .A2(n10422), .ZN(n7263) );
  XNOR2_X1 U9054 ( .A(n7418), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7414) );
  XNOR2_X1 U9055 ( .A(n7415), .B(n7414), .ZN(n7262) );
  NAND2_X1 U9056 ( .A1(n7240), .A2(n7239), .ZN(n10120) );
  AND2_X1 U9057 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8239) );
  NOR2_X1 U9058 ( .A1(n9745), .A2(n7413), .ZN(n7242) );
  AOI211_X1 U9059 ( .C1(n10122), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n8239), .B(
        n7242), .ZN(n7261) );
  INV_X1 U9060 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7243) );
  XNOR2_X1 U9061 ( .A(n7418), .B(n7243), .ZN(n7259) );
  INV_X1 U9062 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7736) );
  MUX2_X1 U9063 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7736), .S(n9636), .Z(n9639)
         );
  AND2_X1 U9064 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9638) );
  NAND2_X1 U9065 ( .A1(n9639), .A2(n9638), .ZN(n9637) );
  NAND2_X1 U9066 ( .A1(n9636), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U9067 ( .A1(n9637), .A2(n7244), .ZN(n7500) );
  INV_X1 U9068 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7787) );
  MUX2_X1 U9069 ( .A(n7787), .B(P1_REG2_REG_2__SCAN_IN), .S(n7245), .Z(n7501)
         );
  NAND2_X1 U9070 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  INV_X1 U9071 ( .A(n7245), .ZN(n7506) );
  NAND2_X1 U9072 ( .A1(n7506), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U9073 ( .A1(n7499), .A2(n7246), .ZN(n9647) );
  INV_X1 U9074 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7247) );
  MUX2_X1 U9075 ( .A(n7247), .B(P1_REG2_REG_3__SCAN_IN), .S(n9644), .Z(n9648)
         );
  NAND2_X1 U9076 ( .A1(n9647), .A2(n9648), .ZN(n10132) );
  OR2_X1 U9077 ( .A1(n9644), .A2(n7247), .ZN(n10130) );
  NAND2_X1 U9078 ( .A1(n10132), .A2(n10130), .ZN(n7249) );
  INV_X1 U9079 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7248) );
  MUX2_X1 U9080 ( .A(n7248), .B(P1_REG2_REG_4__SCAN_IN), .S(n7250), .Z(n10129)
         );
  NAND2_X1 U9081 ( .A1(n7249), .A2(n10129), .ZN(n10134) );
  INV_X1 U9082 ( .A(n7250), .ZN(n10138) );
  NAND2_X1 U9083 ( .A1(n10138), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7251) );
  NAND2_X1 U9084 ( .A1(n10134), .A2(n7251), .ZN(n9659) );
  XNOR2_X1 U9085 ( .A(n9661), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U9086 ( .A1(n9659), .A2(n9660), .ZN(n9658) );
  NAND2_X1 U9087 ( .A1(n9657), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U9088 ( .A1(n9658), .A2(n7252), .ZN(n9673) );
  INV_X1 U9089 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7253) );
  MUX2_X1 U9090 ( .A(n7253), .B(P1_REG2_REG_6__SCAN_IN), .S(n9669), .Z(n9674)
         );
  NAND2_X1 U9091 ( .A1(n9673), .A2(n9674), .ZN(n9672) );
  INV_X1 U9092 ( .A(n9669), .ZN(n7254) );
  NAND2_X1 U9093 ( .A1(n7254), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U9094 ( .A1(n9672), .A2(n7255), .ZN(n7271) );
  XNOR2_X1 U9095 ( .A(n7267), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U9096 ( .A1(n7271), .A2(n7272), .ZN(n7270) );
  INV_X1 U9097 ( .A(n7267), .ZN(n7256) );
  NAND2_X1 U9098 ( .A1(n7256), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U9099 ( .A1(n7270), .A2(n7257), .ZN(n7258) );
  OR2_X1 U9100 ( .A1(n10112), .A2(n5304), .ZN(n8566) );
  NAND2_X1 U9101 ( .A1(n7258), .A2(n7259), .ZN(n7420) );
  OAI211_X1 U9102 ( .C1(n7259), .C2(n7258), .A(n10135), .B(n7420), .ZN(n7260)
         );
  OAI211_X1 U9103 ( .C1(n7262), .C2(n10128), .A(n7261), .B(n7260), .ZN(
        P1_U3251) );
  MUX2_X1 U9104 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10454), .S(n7267), .Z(n7265)
         );
  INV_X1 U9105 ( .A(n7263), .ZN(n7264) );
  NAND2_X1 U9106 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  OAI21_X1 U9107 ( .B1(n9675), .B2(n7266), .A(n9744), .ZN(n7275) );
  NAND2_X1 U9108 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7903) );
  INV_X1 U9109 ( .A(n7903), .ZN(n7269) );
  NOR2_X1 U9110 ( .A1(n9745), .A2(n7267), .ZN(n7268) );
  AOI211_X1 U9111 ( .C1(n10122), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7269), .B(
        n7268), .ZN(n7274) );
  OAI211_X1 U9112 ( .C1(n7272), .C2(n7271), .A(n10135), .B(n7270), .ZN(n7273)
         );
  OAI211_X1 U9113 ( .C1(n7276), .C2(n7275), .A(n7274), .B(n7273), .ZN(P1_U3250) );
  AND2_X1 U9114 ( .A1(n7323), .A2(n7277), .ZN(n7280) );
  OAI211_X1 U9115 ( .C1(n7280), .C2(n7279), .A(n9023), .B(n7278), .ZN(n7296)
         );
  INV_X1 U9116 ( .A(n7281), .ZN(n7283) );
  NAND3_X1 U9117 ( .A1(n7330), .A2(n7283), .A3(n7282), .ZN(n7284) );
  AOI21_X1 U9118 ( .B1(n7285), .B2(n7284), .A(n8976), .ZN(n7294) );
  INV_X1 U9119 ( .A(n7286), .ZN(n7288) );
  NAND3_X1 U9120 ( .A1(n7327), .A2(n7288), .A3(n7287), .ZN(n7289) );
  AOI21_X1 U9121 ( .B1(n7290), .B2(n7289), .A(n9027), .ZN(n7293) );
  INV_X1 U9122 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7291) );
  NOR2_X1 U9123 ( .A1(n9020), .A2(n7291), .ZN(n7292) );
  AND2_X1 U9124 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7519) );
  NOR4_X1 U9125 ( .A1(n7294), .A2(n7293), .A3(n7292), .A4(n7519), .ZN(n7295)
         );
  OAI211_X1 U9126 ( .C1(n9018), .C2(n7297), .A(n7296), .B(n7295), .ZN(P2_U3186) );
  XNOR2_X1 U9127 ( .A(n7299), .B(n7298), .ZN(n7309) );
  AND2_X1 U9128 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7612) );
  AOI21_X1 U9129 ( .B1(n8978), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7612), .ZN(
        n7304) );
  OAI21_X1 U9130 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7301), .A(n7368), .ZN(
        n7302) );
  INV_X1 U9131 ( .A(n9027), .ZN(n8886) );
  NAND2_X1 U9132 ( .A1(n7302), .A2(n8886), .ZN(n7303) );
  OAI211_X1 U9133 ( .C1(n9018), .C2(n7305), .A(n7304), .B(n7303), .ZN(n7306)
         );
  AOI21_X1 U9134 ( .B1(n9006), .B2(n7307), .A(n7306), .ZN(n7308) );
  OAI21_X1 U9135 ( .B1(n7309), .B2(n8150), .A(n7308), .ZN(P2_U3187) );
  XNOR2_X1 U9136 ( .A(n7310), .B(n8758), .ZN(n7322) );
  INV_X1 U9137 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10263) );
  OAI21_X1 U9138 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n7312), .A(n7311), .ZN(
        n7313) );
  AOI22_X1 U9139 ( .A1(n8886), .A2(n7313), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n7318) );
  OAI21_X1 U9140 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7315), .A(n7314), .ZN(
        n7316) );
  NAND2_X1 U9141 ( .A1(n9006), .A2(n7316), .ZN(n7317) );
  OAI211_X1 U9142 ( .C1(n10263), .C2(n9020), .A(n7318), .B(n7317), .ZN(n7319)
         );
  AOI21_X1 U9143 ( .B1(n7320), .B2(n8991), .A(n7319), .ZN(n7321) );
  OAI21_X1 U9144 ( .B1(n8150), .B2(n7322), .A(n7321), .ZN(P2_U3183) );
  INV_X1 U9145 ( .A(n7323), .ZN(n7324) );
  AOI21_X1 U9146 ( .B1(n7326), .B2(n7325), .A(n7324), .ZN(n7337) );
  INV_X1 U9147 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10521) );
  OAI21_X1 U9148 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7328), .A(n7327), .ZN(
        n7329) );
  AOI22_X1 U9149 ( .A1(n8886), .A2(n7329), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n7334) );
  OAI21_X1 U9150 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7331), .A(n7330), .ZN(
        n7332) );
  NAND2_X1 U9151 ( .A1(n9006), .A2(n7332), .ZN(n7333) );
  OAI211_X1 U9152 ( .C1(n10521), .C2(n9020), .A(n7334), .B(n7333), .ZN(n7335)
         );
  AOI21_X1 U9153 ( .B1(n4537), .B2(n8991), .A(n7335), .ZN(n7336) );
  OAI21_X1 U9154 ( .B1(n7337), .B2(n8150), .A(n7336), .ZN(P2_U3185) );
  INV_X1 U9155 ( .A(n7670), .ZN(n7560) );
  INV_X1 U9156 ( .A(n7338), .ZN(n7340) );
  OAI222_X1 U9157 ( .A1(P1_U3086), .A2(n7560), .B1(n10114), .B2(n7340), .C1(
        n10607), .C2(n10115), .ZN(P1_U3343) );
  OAI222_X1 U9158 ( .A1(P2_U3151), .A2(n7341), .B1(n9455), .B2(n7340), .C1(
        n7339), .C2(n9449), .ZN(P2_U3283) );
  NAND2_X1 U9159 ( .A1(n7343), .A2(n7342), .ZN(n7399) );
  INV_X1 U9160 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U9161 ( .A1(n7399), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7346) );
  AOI22_X1 U9162 ( .A1(n8845), .A2(n10198), .B1(n8851), .B2(n7344), .ZN(n7345)
         );
  OAI211_X1 U9163 ( .C1(n7351), .C2(n8853), .A(n7346), .B(n7345), .ZN(P2_U3172) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10377) );
  INV_X1 U9165 ( .A(n7347), .ZN(n7349) );
  OAI222_X1 U9166 ( .A1(n9449), .A2(n10377), .B1(n9455), .B2(n7349), .C1(
        P2_U3151), .C2(n7348), .ZN(P2_U3282) );
  INV_X1 U9167 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7350) );
  INV_X1 U9168 ( .A(n7673), .ZN(n7690) );
  OAI222_X1 U9169 ( .A1(n10115), .A2(n7350), .B1(n10114), .B2(n7349), .C1(
        P1_U3086), .C2(n7690), .ZN(P1_U3342) );
  INV_X1 U9170 ( .A(n7351), .ZN(n7523) );
  OAI21_X1 U9171 ( .B1(n10202), .B2(n10238), .A(n7523), .ZN(n7352) );
  NAND2_X1 U9172 ( .A1(n10198), .A2(n10199), .ZN(n7524) );
  OAI211_X1 U9173 ( .C1(n10239), .C2(n7537), .A(n7352), .B(n7524), .ZN(n7358)
         );
  NAND2_X1 U9174 ( .A1(n7358), .A2(n10257), .ZN(n7353) );
  OAI21_X1 U9175 ( .B1(n10257), .B2(n7026), .A(n7353), .ZN(P2_U3459) );
  INV_X1 U9176 ( .A(n7354), .ZN(n7356) );
  OAI222_X1 U9177 ( .A1(n9449), .A2(n4552), .B1(n9455), .B2(n7356), .C1(
        P2_U3151), .C2(n7355), .ZN(P2_U3281) );
  INV_X1 U9178 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7357) );
  INV_X1 U9179 ( .A(n7935), .ZN(n7929) );
  OAI222_X1 U9180 ( .A1(n10115), .A2(n7357), .B1(n10114), .B2(n7356), .C1(
        P1_U3086), .C2(n7929), .ZN(P1_U3341) );
  INV_X1 U9181 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U9182 ( .A1(n7358), .A2(n10245), .ZN(n7359) );
  OAI21_X1 U9183 ( .B1(n10396), .B2(n10245), .A(n7359), .ZN(P2_U3390) );
  INV_X1 U9184 ( .A(n7360), .ZN(n7393) );
  AOI22_X1 U9185 ( .A1(n8928), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9453), .ZN(n7361) );
  OAI21_X1 U9186 ( .B1(n7393), .B2(n9455), .A(n7361), .ZN(P2_U3280) );
  INV_X1 U9187 ( .A(n7456), .ZN(n7362) );
  AOI21_X1 U9188 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(n7383) );
  NAND2_X1 U9189 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7760) );
  OAI21_X1 U9190 ( .B1(n9020), .B2(n10637), .A(n7760), .ZN(n7372) );
  INV_X1 U9191 ( .A(n7365), .ZN(n7367) );
  NAND3_X1 U9192 ( .A1(n7368), .A2(n7367), .A3(n7366), .ZN(n7369) );
  AOI21_X1 U9193 ( .B1(n7370), .B2(n7369), .A(n9027), .ZN(n7371) );
  AOI211_X1 U9194 ( .C1(n8991), .C2(n7373), .A(n7372), .B(n7371), .ZN(n7382)
         );
  INV_X1 U9195 ( .A(n7300), .ZN(n7377) );
  INV_X1 U9196 ( .A(n7374), .ZN(n7376) );
  NOR3_X1 U9197 ( .A1(n7377), .A2(n7376), .A3(n7375), .ZN(n7380) );
  INV_X1 U9198 ( .A(n7378), .ZN(n7379) );
  OAI21_X1 U9199 ( .B1(n7380), .B2(n7379), .A(n9006), .ZN(n7381) );
  OAI211_X1 U9200 ( .C1(n7383), .C2(n8150), .A(n7382), .B(n7381), .ZN(P2_U3188) );
  XOR2_X1 U9201 ( .A(n7384), .B(n7385), .Z(n7390) );
  AOI22_X1 U9202 ( .A1(n8859), .A2(n10198), .B1(n8851), .B2(n10204), .ZN(n7386) );
  OAI21_X1 U9203 ( .B1(n7387), .B2(n8861), .A(n7386), .ZN(n7388) );
  AOI21_X1 U9204 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7399), .A(n7388), .ZN(
        n7389) );
  OAI21_X1 U9205 ( .B1(n8853), .B2(n7390), .A(n7389), .ZN(P2_U3177) );
  INV_X1 U9206 ( .A(n7391), .ZN(n7407) );
  AOI22_X1 U9207 ( .A1(n9702), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10106), .ZN(n7392) );
  OAI21_X1 U9208 ( .B1(n7407), .B2(n10114), .A(n7392), .ZN(P1_U3339) );
  INV_X1 U9209 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7394) );
  INV_X1 U9210 ( .A(n9692), .ZN(n7938) );
  OAI222_X1 U9211 ( .A1(n10115), .A2(n7394), .B1(n10114), .B2(n7393), .C1(
        P1_U3086), .C2(n7938), .ZN(P1_U3340) );
  XOR2_X1 U9212 ( .A(n7396), .B(n7395), .Z(n7405) );
  INV_X1 U9213 ( .A(n8878), .ZN(n7398) );
  OAI22_X1 U9214 ( .A1(n8866), .A2(n9338), .B1(n7398), .B2(n8848), .ZN(n7403)
         );
  INV_X1 U9215 ( .A(n7399), .ZN(n7401) );
  INV_X1 U9216 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7400) );
  NOR2_X1 U9217 ( .A1(n7401), .A2(n7400), .ZN(n7402) );
  AOI211_X1 U9218 ( .C1(n8845), .C2(n7397), .A(n7403), .B(n7402), .ZN(n7404)
         );
  OAI21_X1 U9219 ( .B1(n8853), .B2(n7405), .A(n7404), .ZN(P2_U3162) );
  OAI222_X1 U9220 ( .A1(P2_U3151), .A2(n8958), .B1(n9455), .B2(n7407), .C1(
        n7406), .C2(n9449), .ZN(P2_U3279) );
  INV_X1 U9221 ( .A(n7408), .ZN(n7411) );
  INV_X1 U9222 ( .A(n8980), .ZN(n8954) );
  OAI222_X1 U9223 ( .A1(n9449), .A2(n7409), .B1(n9455), .B2(n7411), .C1(
        P2_U3151), .C2(n8954), .ZN(P2_U3278) );
  INV_X1 U9224 ( .A(n9725), .ZN(n7410) );
  OAI222_X1 U9225 ( .A1(n10115), .A2(n10592), .B1(n10114), .B2(n7411), .C1(
        P1_U3086), .C2(n7410), .ZN(P1_U3338) );
  INV_X1 U9226 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7412) );
  OAI22_X1 U9227 ( .A1(n7415), .A2(n7414), .B1(n7413), .B2(n7412), .ZN(n7474)
         );
  XNOR2_X1 U9228 ( .A(n7479), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7475) );
  NOR2_X1 U9229 ( .A1(n7479), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7430) );
  XNOR2_X1 U9230 ( .A(n7422), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7433) );
  INV_X1 U9231 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7553) );
  XNOR2_X1 U9232 ( .A(n7554), .B(n7553), .ZN(n7555) );
  XNOR2_X1 U9233 ( .A(n7556), .B(n7555), .ZN(n7429) );
  AND2_X1 U9234 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7417) );
  NOR2_X1 U9235 ( .A1(n9745), .A2(n7554), .ZN(n7416) );
  AOI211_X1 U9236 ( .C1(n10122), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7417), .B(
        n7416), .ZN(n7428) );
  NAND2_X1 U9237 ( .A1(n7418), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7419) );
  NAND2_X1 U9238 ( .A1(n7420), .A2(n7419), .ZN(n7471) );
  XNOR2_X1 U9239 ( .A(n7479), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7472) );
  OR2_X1 U9240 ( .A1(n7471), .A2(n7472), .ZN(n7469) );
  OR2_X1 U9241 ( .A1(n7479), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U9242 ( .A1(n7469), .A2(n7421), .ZN(n7436) );
  XNOR2_X1 U9243 ( .A(n7422), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9244 ( .A1(n7422), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9245 ( .A1(n7434), .A2(n7423), .ZN(n7426) );
  INV_X1 U9246 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7424) );
  MUX2_X1 U9247 ( .A(n7424), .B(P1_REG2_REG_11__SCAN_IN), .S(n7554), .Z(n7425)
         );
  NAND2_X1 U9248 ( .A1(n7426), .A2(n7425), .ZN(n7565) );
  OAI211_X1 U9249 ( .C1(n7426), .C2(n7425), .A(n7565), .B(n10135), .ZN(n7427)
         );
  OAI211_X1 U9250 ( .C1(n7429), .C2(n10128), .A(n7428), .B(n7427), .ZN(
        P1_U3254) );
  OR2_X1 U9251 ( .A1(n7473), .A2(n7430), .ZN(n7432) );
  AOI211_X1 U9252 ( .C1(n7433), .C2(n7432), .A(n10128), .B(n7431), .ZN(n7442)
         );
  INV_X1 U9253 ( .A(n7434), .ZN(n7435) );
  AOI211_X1 U9254 ( .C1(n7437), .C2(n7436), .A(n9729), .B(n7435), .ZN(n7441)
         );
  NAND2_X1 U9255 ( .A1(n10122), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U9256 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8202) );
  OAI211_X1 U9257 ( .C1(n9745), .C2(n7439), .A(n7438), .B(n8202), .ZN(n7440)
         );
  OR3_X1 U9258 ( .A1(n7442), .A2(n7441), .A3(n7440), .ZN(P1_U3253) );
  XNOR2_X1 U9259 ( .A(n7444), .B(n7443), .ZN(n7491) );
  AND2_X1 U9260 ( .A1(n6537), .A2(n9567), .ZN(n7779) );
  OR2_X1 U9261 ( .A1(n7445), .A2(P1_U3086), .ZN(n8386) );
  AOI22_X1 U9262 ( .A1(n9602), .A2(n7779), .B1(n8386), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U9263 ( .A1(n4405), .A2(n7780), .ZN(n7446) );
  OAI211_X1 U9264 ( .C1(n7491), .C2(n9589), .A(n7447), .B(n7446), .ZN(P1_U3232) );
  AND2_X1 U9265 ( .A1(n6538), .A2(n7448), .ZN(n8585) );
  NOR2_X1 U9266 ( .A1(n7725), .A2(n8585), .ZN(n8534) );
  AOI21_X1 U9267 ( .B1(n10185), .B2(n9945), .A(n8534), .ZN(n7449) );
  AOI211_X1 U9268 ( .C1(n7777), .C2(n7780), .A(n7779), .B(n7449), .ZN(n7508)
         );
  NAND2_X1 U9269 ( .A1(n10192), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7450) );
  OAI21_X1 U9270 ( .B1(n7508), .B2(n10192), .A(n7450), .ZN(P1_U3522) );
  INV_X1 U9271 ( .A(n7451), .ZN(n7452) );
  NOR2_X1 U9272 ( .A1(n7453), .A2(n7452), .ZN(n7457) );
  INV_X1 U9273 ( .A(n7454), .ZN(n7455) );
  AOI21_X1 U9274 ( .B1(n7457), .B2(n7456), .A(n7455), .ZN(n7468) );
  OAI21_X1 U9275 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n4517), .A(n7458), .ZN(
        n7462) );
  NAND2_X1 U9276 ( .A1(n8978), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7459) );
  NAND2_X1 U9277 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7833) );
  OAI211_X1 U9278 ( .C1(n9018), .C2(n7460), .A(n7459), .B(n7833), .ZN(n7461)
         );
  AOI21_X1 U9279 ( .B1(n7462), .B2(n8886), .A(n7461), .ZN(n7467) );
  OAI21_X1 U9280 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7464), .A(n7463), .ZN(
        n7465) );
  NAND2_X1 U9281 ( .A1(n7465), .A2(n9006), .ZN(n7466) );
  OAI211_X1 U9282 ( .C1(n7468), .C2(n8150), .A(n7467), .B(n7466), .ZN(P2_U3189) );
  INV_X1 U9283 ( .A(n7469), .ZN(n7470) );
  AOI21_X1 U9284 ( .B1(n7472), .B2(n7471), .A(n7470), .ZN(n7481) );
  NAND2_X1 U9285 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8353) );
  OAI21_X1 U9286 ( .B1(n9749), .B2(n10594), .A(n8353), .ZN(n7478) );
  AOI21_X1 U9287 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7476) );
  NOR2_X1 U9288 ( .A1(n7476), .A2(n10128), .ZN(n7477) );
  AOI211_X1 U9289 ( .C1(n10139), .C2(n7479), .A(n7478), .B(n7477), .ZN(n7480)
         );
  OAI21_X1 U9290 ( .B1(n7481), .B2(n9729), .A(n7480), .ZN(P1_U3252) );
  INV_X1 U9291 ( .A(n7482), .ZN(n7483) );
  AOI211_X1 U9292 ( .C1(n7485), .C2(n7484), .A(n8853), .B(n7483), .ZN(n7490)
         );
  MUX2_X1 U9293 ( .A(P2_STATE_REG_SCAN_IN), .B(n8317), .S(n7547), .Z(n7487) );
  AOI22_X1 U9294 ( .A1(n8859), .A2(n7397), .B1(n8851), .B2(n7548), .ZN(n7486)
         );
  OAI211_X1 U9295 ( .C1(n7488), .C2(n8861), .A(n7487), .B(n7486), .ZN(n7489)
         );
  OR2_X1 U9296 ( .A1(n7490), .A2(n7489), .ZN(P2_U3158) );
  NAND3_X1 U9297 ( .A1(n7491), .A2(n7492), .A3(n7493), .ZN(n7496) );
  OAI21_X1 U9298 ( .B1(n7493), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7492), .ZN(
        n10117) );
  INV_X1 U9299 ( .A(n8566), .ZN(n7494) );
  AOI22_X1 U9300 ( .A1(n4879), .A2(n10117), .B1(n7494), .B2(n9638), .ZN(n7495)
         );
  NAND3_X1 U9301 ( .A1(n7496), .A2(P1_U3973), .A3(n7495), .ZN(n10140) );
  INV_X1 U9302 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10575) );
  INV_X1 U9303 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10483) );
  OAI22_X1 U9304 ( .A1(n9749), .A2(n10575), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10483), .ZN(n7505) );
  XNOR2_X1 U9305 ( .A(n7498), .B(n7497), .ZN(n7503) );
  OAI211_X1 U9306 ( .C1(n7501), .C2(n7500), .A(n10135), .B(n7499), .ZN(n7502)
         );
  OAI21_X1 U9307 ( .B1(n10128), .B2(n7503), .A(n7502), .ZN(n7504) );
  AOI211_X1 U9308 ( .C1(n7506), .C2(n10139), .A(n7505), .B(n7504), .ZN(n7507)
         );
  NAND2_X1 U9309 ( .A1(n10140), .A2(n7507), .ZN(P1_U3245) );
  INV_X1 U9310 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7510) );
  OR2_X1 U9311 ( .A1(n7508), .A2(n10187), .ZN(n7509) );
  OAI21_X1 U9312 ( .B1(n10189), .B2(n7510), .A(n7509), .ZN(P1_U3453) );
  INV_X1 U9313 ( .A(n7511), .ZN(n7552) );
  AOI22_X1 U9314 ( .A1(n9739), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10106), .ZN(n7512) );
  OAI21_X1 U9315 ( .B1(n7552), .B2(n10114), .A(n7512), .ZN(P1_U3337) );
  OAI21_X1 U9316 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7516) );
  NAND2_X1 U9317 ( .A1(n7516), .A2(n8855), .ZN(n7521) );
  OAI22_X1 U9318 ( .A1(n8866), .A2(n10227), .B1(n7517), .B2(n8861), .ZN(n7518)
         );
  AOI211_X1 U9319 ( .C1(n8859), .C2(n10200), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI211_X1 U9320 ( .C1(n7622), .C2(n8317), .A(n7521), .B(n7520), .ZN(P2_U3170) );
  NAND3_X1 U9321 ( .A1(n7523), .A2(n7522), .A3(n10239), .ZN(n7525) );
  NAND2_X1 U9322 ( .A1(n7525), .A2(n7524), .ZN(n7534) );
  INV_X1 U9323 ( .A(n7526), .ZN(n7527) );
  OR2_X1 U9324 ( .A1(n7527), .A2(n7529), .ZN(n7531) );
  NAND2_X1 U9325 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  MUX2_X1 U9326 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n7534), .S(n10212), .Z(n7539)
         );
  INV_X1 U9327 ( .A(n7542), .ZN(n7535) );
  INV_X1 U9328 ( .A(n9242), .ZN(n10203) );
  OAI22_X1 U9329 ( .A1(n9204), .A2(n7537), .B1(n7536), .B2(n9240), .ZN(n7538)
         );
  OR2_X1 U9330 ( .A1(n7539), .A2(n7538), .ZN(P2_U3233) );
  NAND2_X1 U9331 ( .A1(n7540), .A2(n4797), .ZN(n7541) );
  OR2_X1 U9332 ( .A1(n10209), .A2(n8098), .ZN(n7543) );
  XNOR2_X1 U9333 ( .A(n6890), .B(n7544), .ZN(n10219) );
  XNOR2_X1 U9334 ( .A(n6890), .B(n7545), .ZN(n7546) );
  AOI222_X1 U9335 ( .A1(n10202), .A2(n7546), .B1(n8876), .B2(n10199), .C1(
        n7397), .C2(n9236), .ZN(n10220) );
  MUX2_X1 U9336 ( .A(n10467), .B(n10220), .S(n10212), .Z(n7550) );
  AOI22_X1 U9337 ( .A1(n9265), .A2(n7548), .B1(n10205), .B2(n7547), .ZN(n7549)
         );
  OAI211_X1 U9338 ( .C1(n9268), .C2(n10219), .A(n7550), .B(n7549), .ZN(
        P2_U3230) );
  INV_X1 U9339 ( .A(n8993), .ZN(n9014) );
  OAI222_X1 U9340 ( .A1(P2_U3151), .A2(n9014), .B1(n9455), .B2(n7552), .C1(
        n7551), .C2(n9449), .ZN(P2_U3277) );
  XNOR2_X1 U9341 ( .A(n7670), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7558) );
  AOI21_X1 U9342 ( .B1(n7558), .B2(n7557), .A(n7681), .ZN(n7572) );
  NOR2_X1 U9343 ( .A1(n7559), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8004) );
  NOR2_X1 U9344 ( .A1(n9745), .A2(n7560), .ZN(n7561) );
  AOI211_X1 U9345 ( .C1(n10122), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n8004), .B(
        n7561), .ZN(n7571) );
  INV_X1 U9346 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7562) );
  MUX2_X1 U9347 ( .A(n7562), .B(P1_REG2_REG_12__SCAN_IN), .S(n7670), .Z(n7568)
         );
  NAND2_X1 U9348 ( .A1(n7563), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9349 ( .A1(n7565), .A2(n7564), .ZN(n7567) );
  INV_X1 U9350 ( .A(n7672), .ZN(n7566) );
  AOI21_X1 U9351 ( .B1(n7568), .B2(n7567), .A(n7566), .ZN(n7569) );
  OR2_X1 U9352 ( .A1(n7569), .A2(n9729), .ZN(n7570) );
  OAI211_X1 U9353 ( .C1(n7572), .C2(n10128), .A(n7571), .B(n7570), .ZN(
        P1_U3255) );
  NAND2_X1 U9354 ( .A1(n6633), .A2(n7574), .ZN(n7576) );
  NAND2_X1 U9355 ( .A1(n7576), .A2(n7575), .ZN(n9340) );
  INV_X1 U9356 ( .A(n9340), .ZN(n7585) );
  XNOR2_X1 U9357 ( .A(n7574), .B(n7577), .ZN(n7581) );
  NAND2_X1 U9358 ( .A1(n8878), .A2(n9236), .ZN(n7578) );
  OAI21_X1 U9359 ( .B1(n7579), .B2(n9261), .A(n7578), .ZN(n7580) );
  AOI21_X1 U9360 ( .B1(n7581), .B2(n10202), .A(n7580), .ZN(n9341) );
  INV_X1 U9361 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7582) );
  MUX2_X1 U9362 ( .A(n9341), .B(n7582), .S(n9246), .Z(n7584) );
  AOI22_X1 U9363 ( .A1(n9265), .A2(n4461), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10205), .ZN(n7583) );
  OAI211_X1 U9364 ( .C1(n7585), .C2(n9268), .A(n7584), .B(n7583), .ZN(P2_U3232) );
  INV_X1 U9365 ( .A(n7586), .ZN(n7587) );
  AOI21_X1 U9366 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7606) );
  INV_X1 U9367 ( .A(n7590), .ZN(n7594) );
  INV_X1 U9368 ( .A(n7591), .ZN(n7593) );
  NOR3_X1 U9369 ( .A1(n7594), .A2(n7593), .A3(n7592), .ZN(n7597) );
  INV_X1 U9370 ( .A(n7595), .ZN(n7596) );
  OAI21_X1 U9371 ( .B1(n7597), .B2(n7596), .A(n9023), .ZN(n7605) );
  INV_X1 U9372 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U9373 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8055) );
  OAI21_X1 U9374 ( .B1(n9020), .B2(n10277), .A(n8055), .ZN(n7602) );
  NAND2_X1 U9375 ( .A1(n7598), .A2(n10468), .ZN(n7599) );
  AOI21_X1 U9376 ( .B1(n7600), .B2(n7599), .A(n9027), .ZN(n7601) );
  AOI211_X1 U9377 ( .C1(n8991), .C2(n7603), .A(n7602), .B(n7601), .ZN(n7604)
         );
  OAI211_X1 U9378 ( .C1(n7606), .C2(n8976), .A(n7605), .B(n7604), .ZN(P2_U3191) );
  XNOR2_X1 U9379 ( .A(n7608), .B(n7607), .ZN(n7609) );
  NAND2_X1 U9380 ( .A1(n7609), .A2(n8855), .ZN(n7614) );
  OAI22_X1 U9381 ( .A1(n8866), .A2(n10231), .B1(n7610), .B2(n8861), .ZN(n7611)
         );
  AOI211_X1 U9382 ( .C1(n8859), .C2(n8876), .A(n7612), .B(n7611), .ZN(n7613)
         );
  OAI211_X1 U9383 ( .C1(n7714), .C2(n8317), .A(n7614), .B(n7613), .ZN(P2_U3167) );
  NAND2_X1 U9384 ( .A1(n7544), .A2(n7615), .ZN(n7702) );
  NAND2_X1 U9385 ( .A1(n7702), .A2(n7616), .ZN(n7617) );
  XNOR2_X1 U9386 ( .A(n7617), .B(n7618), .ZN(n10225) );
  XNOR2_X1 U9387 ( .A(n7619), .B(n7618), .ZN(n7620) );
  AOI222_X1 U9388 ( .A1(n10202), .A2(n7620), .B1(n8875), .B2(n10199), .C1(
        n10200), .C2(n9236), .ZN(n10226) );
  MUX2_X1 U9389 ( .A(n7621), .B(n10226), .S(n10212), .Z(n7626) );
  INV_X1 U9390 ( .A(n7622), .ZN(n7623) );
  AOI22_X1 U9391 ( .A1(n9265), .A2(n7624), .B1(n10205), .B2(n7623), .ZN(n7625)
         );
  OAI211_X1 U9392 ( .C1(n9268), .C2(n10225), .A(n7626), .B(n7625), .ZN(
        P2_U3229) );
  XNOR2_X1 U9393 ( .A(n7628), .B(n7627), .ZN(n7629) );
  NAND2_X1 U9394 ( .A1(n7629), .A2(n5931), .ZN(n7633) );
  OR2_X1 U9395 ( .A1(n7651), .A2(n9593), .ZN(n7631) );
  NAND2_X1 U9396 ( .A1(n6537), .A2(n9595), .ZN(n7630) );
  NAND2_X1 U9397 ( .A1(n7631), .A2(n7630), .ZN(n7642) );
  AOI22_X1 U9398 ( .A1(n7642), .A2(n9602), .B1(n8386), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7632) );
  OAI211_X1 U9399 ( .C1(n4416), .C2(n9605), .A(n7633), .B(n7632), .ZN(P1_U3237) );
  INV_X1 U9400 ( .A(n7634), .ZN(n8369) );
  OAI222_X1 U9401 ( .A1(n9449), .A2(n7635), .B1(n9455), .B2(n8369), .C1(n9017), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI21_X1 U9402 ( .B1(n7638), .B2(n7636), .A(n7637), .ZN(n7784) );
  INV_X1 U9403 ( .A(n7817), .ZN(n7639) );
  AOI211_X1 U9404 ( .C1(n7640), .C2(n7735), .A(n9949), .B(n7639), .ZN(n7791)
         );
  XNOR2_X1 U9405 ( .A(n7641), .B(n7636), .ZN(n7644) );
  INV_X1 U9406 ( .A(n7642), .ZN(n7643) );
  OAI21_X1 U9407 ( .B1(n7644), .B2(n9945), .A(n7643), .ZN(n7786) );
  AOI211_X1 U9408 ( .C1(n10055), .C2(n7784), .A(n7791), .B(n7786), .ZN(n7767)
         );
  OAI22_X1 U9409 ( .A1(n10036), .A2(n4416), .B1(n10194), .B2(n10534), .ZN(
        n7645) );
  INV_X1 U9410 ( .A(n7645), .ZN(n7646) );
  OAI21_X1 U9411 ( .B1(n7767), .B2(n10192), .A(n7646), .ZN(P1_U3524) );
  NOR2_X1 U9412 ( .A1(n4513), .A2(n7647), .ZN(n7648) );
  XNOR2_X1 U9413 ( .A(n7648), .B(n8536), .ZN(n10153) );
  XNOR2_X1 U9414 ( .A(n7650), .B(n7649), .ZN(n7652) );
  OAI22_X1 U9415 ( .A1(n7651), .A2(n8398), .B1(n8417), .B2(n9593), .ZN(n9537)
         );
  AOI21_X1 U9416 ( .B1(n7652), .B2(n9964), .A(n9537), .ZN(n10166) );
  INV_X1 U9417 ( .A(n7653), .ZN(n7654) );
  OAI211_X1 U9418 ( .C1(n7768), .C2(n7816), .A(n7654), .B(n9992), .ZN(n10161)
         );
  OAI211_X1 U9419 ( .C1(n10185), .C2(n10153), .A(n10166), .B(n10161), .ZN(
        n7770) );
  OAI22_X1 U9420 ( .A1(n10036), .A2(n7768), .B1(n10194), .B2(n10574), .ZN(
        n7655) );
  AOI21_X1 U9421 ( .B1(n7770), .B2(n10194), .A(n7655), .ZN(n7656) );
  INV_X1 U9422 ( .A(n7656), .ZN(P1_U3526) );
  INV_X1 U9423 ( .A(n7657), .ZN(n7658) );
  NOR2_X1 U9424 ( .A1(n7658), .A2(n7661), .ZN(n7796) );
  AOI21_X1 U9425 ( .B1(n7658), .B2(n7661), .A(n7796), .ZN(n7986) );
  OAI21_X1 U9426 ( .B1(n7661), .B2(n7660), .A(n7659), .ZN(n7664) );
  OR2_X1 U9427 ( .A1(n6475), .A2(n8398), .ZN(n7663) );
  OR2_X1 U9428 ( .A1(n8423), .A2(n9593), .ZN(n7662) );
  NAND2_X1 U9429 ( .A1(n7663), .A2(n7662), .ZN(n9507) );
  AOI21_X1 U9430 ( .B1(n7664), .B2(n9964), .A(n9507), .ZN(n7993) );
  OAI211_X1 U9431 ( .C1(n7653), .C2(n8425), .A(n9992), .B(n7803), .ZN(n7989)
         );
  OAI211_X1 U9432 ( .C1(n10185), .C2(n7986), .A(n7993), .B(n7989), .ZN(n7774)
         );
  OAI22_X1 U9433 ( .A1(n10036), .A2(n8425), .B1(n10194), .B2(n7236), .ZN(n7665) );
  AOI21_X1 U9434 ( .B1(n7774), .B2(n10194), .A(n7665), .ZN(n7666) );
  INV_X1 U9435 ( .A(n7666), .ZN(P1_U3527) );
  NOR2_X1 U9436 ( .A1(n7670), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7680) );
  XNOR2_X1 U9437 ( .A(n7673), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7684) );
  NOR3_X1 U9438 ( .A1(n7681), .A2(n7680), .A3(n7684), .ZN(n7682) );
  XNOR2_X1 U9439 ( .A(n7935), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7931) );
  XNOR2_X1 U9440 ( .A(n7932), .B(n7931), .ZN(n7679) );
  NOR2_X1 U9441 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7667), .ZN(n7669) );
  NOR2_X1 U9442 ( .A1(n9745), .A2(n7929), .ZN(n7668) );
  AOI211_X1 U9443 ( .C1(n10122), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7669), .B(
        n7668), .ZN(n7678) );
  OR2_X1 U9444 ( .A1(n7670), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9445 ( .A1(n7672), .A2(n7671), .ZN(n7687) );
  XNOR2_X1 U9446 ( .A(n7673), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9447 ( .A1(n7673), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9448 ( .A1(n7685), .A2(n7674), .ZN(n7676) );
  INV_X1 U9449 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8262) );
  XNOR2_X1 U9450 ( .A(n7935), .B(n8262), .ZN(n7675) );
  NAND2_X1 U9451 ( .A1(n7676), .A2(n7675), .ZN(n7937) );
  OAI211_X1 U9452 ( .C1(n7676), .C2(n7675), .A(n7937), .B(n10135), .ZN(n7677)
         );
  OAI211_X1 U9453 ( .C1(n7679), .C2(n10128), .A(n7678), .B(n7677), .ZN(
        P1_U3257) );
  OR2_X1 U9454 ( .A1(n7681), .A2(n7680), .ZN(n7683) );
  AOI211_X1 U9455 ( .C1(n7684), .C2(n7683), .A(n10128), .B(n7682), .ZN(n7693)
         );
  INV_X1 U9456 ( .A(n7685), .ZN(n7686) );
  AOI211_X1 U9457 ( .C1(n7688), .C2(n7687), .A(n9729), .B(n7686), .ZN(n7692)
         );
  NAND2_X1 U9458 ( .A1(n10122), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9459 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8074) );
  OAI211_X1 U9460 ( .C1(n9745), .C2(n7690), .A(n7689), .B(n8074), .ZN(n7691)
         );
  OR3_X1 U9461 ( .A1(n7693), .A2(n7692), .A3(n7691), .ZN(P1_U3256) );
  NAND2_X1 U9462 ( .A1(n9528), .A2(n7695), .ZN(n7696) );
  XOR2_X1 U9463 ( .A(n7694), .B(n7696), .Z(n7700) );
  OAI22_X1 U9464 ( .A1(n6469), .A2(n8398), .B1(n6475), .B2(n9593), .ZN(n7814)
         );
  AOI22_X1 U9465 ( .A1(n7814), .A2(n9602), .B1(n10180), .B2(n4405), .ZN(n7699)
         );
  MUX2_X1 U9466 ( .A(P1_STATE_REG_SCAN_IN), .B(n9599), .S(n7697), .Z(n7698) );
  OAI211_X1 U9467 ( .C1(n7700), .C2(n9589), .A(n7699), .B(n7698), .ZN(P1_U3218) );
  NAND2_X1 U9468 ( .A1(n7702), .A2(n7701), .ZN(n7704) );
  NAND2_X1 U9469 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  XNOR2_X1 U9470 ( .A(n7705), .B(n7706), .ZN(n10234) );
  NAND2_X1 U9471 ( .A1(n10234), .A2(n8098), .ZN(n7712) );
  AOI22_X1 U9472 ( .A1(n9236), .A2(n8876), .B1(n8874), .B2(n10199), .ZN(n7711)
         );
  INV_X1 U9473 ( .A(n7706), .ZN(n7707) );
  NOR2_X1 U9474 ( .A1(n7708), .A2(n7707), .ZN(n7884) );
  AND2_X1 U9475 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  OAI21_X1 U9476 ( .B1(n7884), .B2(n7709), .A(n10202), .ZN(n7710) );
  NAND3_X1 U9477 ( .A1(n7712), .A2(n7711), .A3(n7710), .ZN(n10232) );
  MUX2_X1 U9478 ( .A(n10232), .B(P2_REG2_REG_5__SCAN_IN), .S(n9246), .Z(n7713)
         );
  INV_X1 U9479 ( .A(n7713), .ZN(n7717) );
  OAI22_X1 U9480 ( .A1(n9204), .A2(n10231), .B1(n7714), .B2(n9240), .ZN(n7715)
         );
  AOI21_X1 U9481 ( .B1(n10234), .B2(n10209), .A(n7715), .ZN(n7716) );
  NAND2_X1 U9482 ( .A1(n7717), .A2(n7716), .ZN(P2_U3228) );
  NAND2_X1 U9483 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  OAI21_X1 U9484 ( .B1(n7725), .B2(n7723), .A(n7724), .ZN(n7729) );
  OAI22_X1 U9485 ( .A1(n5327), .A2(n8398), .B1(n6469), .B2(n9593), .ZN(n8387)
         );
  INV_X1 U9486 ( .A(n7723), .ZN(n8535) );
  XNOR2_X1 U9487 ( .A(n8535), .B(n7726), .ZN(n10177) );
  INV_X1 U9488 ( .A(n10177), .ZN(n7727) );
  NOR2_X1 U9489 ( .A1(n7727), .A2(n8159), .ZN(n7728) );
  AOI211_X1 U9490 ( .C1(n9964), .C2(n7729), .A(n8387), .B(n7728), .ZN(n10174)
         );
  INV_X1 U9491 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U9492 ( .A1(n9951), .A2(n7731), .ZN(n8268) );
  INV_X1 U9493 ( .A(n8268), .ZN(n7740) );
  NAND2_X1 U9494 ( .A1(n7780), .A2(n7733), .ZN(n7734) );
  NAND3_X1 U9495 ( .A1(n7735), .A2(n9992), .A3(n7734), .ZN(n10171) );
  OAI22_X1 U9496 ( .A1(n9953), .A2(n10173), .B1(n10171), .B2(n10160), .ZN(
        n7739) );
  INV_X1 U9497 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7737) );
  OAI22_X1 U9498 ( .A1(n9913), .A2(n7737), .B1(n7736), .B2(n9951), .ZN(n7738)
         );
  AOI211_X1 U9499 ( .C1(n10177), .C2(n7740), .A(n7739), .B(n7738), .ZN(n7741)
         );
  OAI21_X1 U9500 ( .B1(n10167), .B2(n10174), .A(n7741), .ZN(P1_U3292) );
  XNOR2_X1 U9501 ( .A(n7743), .B(n7742), .ZN(n7754) );
  NAND2_X1 U9502 ( .A1(n7744), .A2(n7878), .ZN(n7745) );
  NAND2_X1 U9503 ( .A1(n7745), .A2(n7885), .ZN(n7880) );
  NAND2_X1 U9504 ( .A1(n7880), .A2(n7747), .ZN(n7746) );
  NAND2_X1 U9505 ( .A1(n7746), .A2(n7749), .ZN(n7751) );
  INV_X1 U9506 ( .A(n7747), .ZN(n7748) );
  NOR2_X1 U9507 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  NAND2_X1 U9508 ( .A1(n7880), .A2(n7750), .ZN(n7870) );
  NAND2_X1 U9509 ( .A1(n7751), .A2(n7870), .ZN(n7843) );
  INV_X1 U9510 ( .A(n8098), .ZN(n10207) );
  OR2_X1 U9511 ( .A1(n7843), .A2(n10207), .ZN(n7753) );
  AOI22_X1 U9512 ( .A1(n9236), .A2(n8874), .B1(n8872), .B2(n10199), .ZN(n7752)
         );
  OAI211_X1 U9513 ( .C1(n9256), .C2(n7754), .A(n7753), .B(n7752), .ZN(n7841)
         );
  OAI22_X1 U9514 ( .A1(n7843), .A2(n9334), .B1(n7845), .B2(n10239), .ZN(n7755)
         );
  NOR2_X1 U9515 ( .A1(n7841), .A2(n7755), .ZN(n7894) );
  NAND2_X1 U9516 ( .A1(n10247), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7756) );
  OAI21_X1 U9517 ( .B1(n7894), .B2(n10247), .A(n7756), .ZN(P2_U3411) );
  OAI211_X1 U9518 ( .C1(n7759), .C2(n7758), .A(n7757), .B(n8855), .ZN(n7764)
         );
  NAND2_X1 U9519 ( .A1(n8859), .A2(n8875), .ZN(n7761) );
  OAI211_X1 U9520 ( .C1(n8009), .C2(n8861), .A(n7761), .B(n7760), .ZN(n7762)
         );
  AOI21_X1 U9521 ( .B1(n7891), .B2(n8851), .A(n7762), .ZN(n7763) );
  OAI211_X1 U9522 ( .C1(n7889), .C2(n8317), .A(n7764), .B(n7763), .ZN(P2_U3179) );
  INV_X1 U9523 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10527) );
  OAI22_X1 U9524 ( .A1(n10096), .A2(n4416), .B1(n10189), .B2(n10527), .ZN(
        n7765) );
  INV_X1 U9525 ( .A(n7765), .ZN(n7766) );
  OAI21_X1 U9526 ( .B1(n7767), .B2(n10187), .A(n7766), .ZN(P1_U3459) );
  INV_X1 U9527 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10605) );
  OAI22_X1 U9528 ( .A1(n10096), .A2(n7768), .B1(n10189), .B2(n10605), .ZN(
        n7769) );
  AOI21_X1 U9529 ( .B1(n7770), .B2(n10189), .A(n7769), .ZN(n7771) );
  INV_X1 U9530 ( .A(n7771), .ZN(P1_U3465) );
  INV_X1 U9531 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7772) );
  OAI22_X1 U9532 ( .A1(n10096), .A2(n8425), .B1(n10189), .B2(n7772), .ZN(n7773) );
  AOI21_X1 U9533 ( .B1(n7774), .B2(n10189), .A(n7773), .ZN(n7775) );
  INV_X1 U9534 ( .A(n7775), .ZN(P1_U3468) );
  INV_X1 U9535 ( .A(n8568), .ZN(n7776) );
  NOR3_X1 U9536 ( .A1(n8534), .A2(n7777), .A3(n7776), .ZN(n7778) );
  AOI211_X1 U9537 ( .C1(n10154), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7779), .B(
        n7778), .ZN(n7783) );
  NAND2_X1 U9538 ( .A1(n10167), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7782) );
  NOR2_X1 U9539 ( .A1(n10160), .A2(n9949), .ZN(n9833) );
  OAI21_X1 U9540 ( .B1(n9833), .B2(n10157), .A(n7780), .ZN(n7781) );
  OAI211_X1 U9541 ( .C1(n7783), .C2(n10167), .A(n7782), .B(n7781), .ZN(
        P1_U3293) );
  INV_X1 U9542 ( .A(n7784), .ZN(n7794) );
  NAND2_X1 U9543 ( .A1(n8159), .A2(n7730), .ZN(n7785) );
  NAND2_X1 U9544 ( .A1(n7786), .A2(n9951), .ZN(n7793) );
  OAI22_X1 U9545 ( .A1(n9951), .A2(n7787), .B1(n10483), .B2(n9913), .ZN(n7790)
         );
  NOR2_X1 U9546 ( .A1(n9953), .A2(n4416), .ZN(n7789) );
  AOI211_X1 U9547 ( .C1(n7791), .C2(n9971), .A(n7790), .B(n7789), .ZN(n7792)
         );
  OAI211_X1 U9548 ( .C1(n7794), .C2(n9957), .A(n7793), .B(n7792), .ZN(P1_U3291) );
  NOR2_X1 U9549 ( .A1(n7796), .A2(n7795), .ZN(n7798) );
  XNOR2_X1 U9550 ( .A(n7798), .B(n7797), .ZN(n10143) );
  XOR2_X1 U9551 ( .A(n7799), .B(n7797), .Z(n7802) );
  OR2_X1 U9552 ( .A1(n8417), .A2(n8398), .ZN(n7801) );
  OR2_X1 U9553 ( .A1(n7960), .A2(n9593), .ZN(n7800) );
  NAND2_X1 U9554 ( .A1(n7801), .A2(n7800), .ZN(n9583) );
  AOI21_X1 U9555 ( .B1(n7802), .B2(n9964), .A(n9583), .ZN(n10152) );
  OAI211_X1 U9556 ( .C1(n4992), .C2(n8419), .A(n9992), .B(n7922), .ZN(n10148)
         );
  OAI211_X1 U9557 ( .C1(n10185), .C2(n10143), .A(n10152), .B(n10148), .ZN(
        n7808) );
  OAI22_X1 U9558 ( .A1(n10036), .A2(n8419), .B1(n10194), .B2(n10422), .ZN(
        n7804) );
  AOI21_X1 U9559 ( .B1(n7808), .B2(n10194), .A(n7804), .ZN(n7805) );
  INV_X1 U9560 ( .A(n7805), .ZN(P1_U3528) );
  INV_X1 U9561 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7806) );
  OAI22_X1 U9562 ( .A1(n10096), .A2(n8419), .B1(n10189), .B2(n7806), .ZN(n7807) );
  AOI21_X1 U9563 ( .B1(n7808), .B2(n10189), .A(n7807), .ZN(n7809) );
  INV_X1 U9564 ( .A(n7809), .ZN(P1_U3471) );
  INV_X1 U9565 ( .A(n7810), .ZN(n7812) );
  AOI21_X1 U9566 ( .B1(n7812), .B2(n4409), .A(n4513), .ZN(n10184) );
  OAI21_X1 U9567 ( .B1(n4519), .B2(n4409), .A(n7813), .ZN(n7815) );
  AOI21_X1 U9568 ( .B1(n7815), .B2(n9964), .A(n7814), .ZN(n10183) );
  MUX2_X1 U9569 ( .A(n10183), .B(n7247), .S(n10167), .Z(n7821) );
  AOI211_X1 U9570 ( .C1(n10180), .C2(n7817), .A(n9949), .B(n7816), .ZN(n10179)
         );
  OAI22_X1 U9571 ( .A1(n9953), .A2(n7818), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9913), .ZN(n7819) );
  AOI21_X1 U9572 ( .B1(n10179), .B2(n9971), .A(n7819), .ZN(n7820) );
  OAI211_X1 U9573 ( .C1(n10184), .C2(n9957), .A(n7821), .B(n7820), .ZN(
        P1_U3290) );
  INV_X1 U9574 ( .A(n7822), .ZN(n7826) );
  OAI222_X1 U9575 ( .A1(n10115), .A2(n7824), .B1(n10114), .B2(n7826), .C1(
        n7823), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U9576 ( .A1(P2_U3151), .A2(n7827), .B1(n9455), .B2(n7826), .C1(
        n7825), .C2(n9449), .ZN(P2_U3275) );
  NAND2_X1 U9577 ( .A1(n7757), .A2(n7828), .ZN(n7831) );
  INV_X1 U9578 ( .A(n7829), .ZN(n7830) );
  AOI21_X1 U9579 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7840) );
  INV_X1 U9580 ( .A(n7833), .ZN(n7834) );
  AOI21_X1 U9581 ( .B1(n8859), .B2(n8874), .A(n7834), .ZN(n7835) );
  OAI21_X1 U9582 ( .B1(n8007), .B2(n8861), .A(n7835), .ZN(n7837) );
  NOR2_X1 U9583 ( .A1(n8317), .A2(n7844), .ZN(n7836) );
  AOI211_X1 U9584 ( .C1(n7838), .C2(n8851), .A(n7837), .B(n7836), .ZN(n7839)
         );
  OAI21_X1 U9585 ( .B1(n7840), .B2(n8853), .A(n7839), .ZN(P2_U3153) );
  MUX2_X1 U9586 ( .A(n7841), .B(P2_REG2_REG_7__SCAN_IN), .S(n9246), .Z(n7842)
         );
  INV_X1 U9587 ( .A(n7842), .ZN(n7849) );
  INV_X1 U9588 ( .A(n7843), .ZN(n7847) );
  OAI22_X1 U9589 ( .A1(n9204), .A2(n7845), .B1(n7844), .B2(n9240), .ZN(n7846)
         );
  AOI21_X1 U9590 ( .B1(n7847), .B2(n10209), .A(n7846), .ZN(n7848) );
  NAND2_X1 U9591 ( .A1(n7849), .A2(n7848), .ZN(P2_U3226) );
  INV_X1 U9592 ( .A(n7850), .ZN(n7851) );
  NOR2_X1 U9593 ( .A1(n7852), .A2(n7851), .ZN(n7856) );
  INV_X1 U9594 ( .A(n7853), .ZN(n7854) );
  AOI21_X1 U9595 ( .B1(n7856), .B2(n7855), .A(n7854), .ZN(n7868) );
  OAI21_X1 U9596 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7858), .A(n7857), .ZN(
        n7862) );
  NOR2_X1 U9597 ( .A1(n9018), .A2(n7859), .ZN(n7861) );
  INV_X1 U9598 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U9599 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8211) );
  OAI21_X1 U9600 ( .B1(n9020), .B2(n10260), .A(n8211), .ZN(n7860) );
  AOI211_X1 U9601 ( .C1(n7862), .C2(n8886), .A(n7861), .B(n7860), .ZN(n7867)
         );
  OAI21_X1 U9602 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7864), .A(n7863), .ZN(
        n7865) );
  NAND2_X1 U9603 ( .A1(n7865), .A2(n9006), .ZN(n7866) );
  OAI211_X1 U9604 ( .C1(n7868), .C2(n8150), .A(n7867), .B(n7866), .ZN(P2_U3193) );
  NAND2_X1 U9605 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  XOR2_X1 U9606 ( .A(n7873), .B(n7871), .Z(n8021) );
  INV_X1 U9607 ( .A(n9236), .ZN(n9259) );
  XNOR2_X1 U9608 ( .A(n7872), .B(n7873), .ZN(n7874) );
  OAI222_X1 U9609 ( .A1(n9261), .A2(n8096), .B1(n9259), .B2(n8009), .C1(n9256), 
        .C2(n7874), .ZN(n8018) );
  AOI21_X1 U9610 ( .B1(n10238), .B2(n8021), .A(n8018), .ZN(n7994) );
  INV_X1 U9611 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7875) );
  OAI22_X1 U9612 ( .A1(n9413), .A2(n8017), .B1(n7875), .B2(n10245), .ZN(n7876)
         );
  INV_X1 U9613 ( .A(n7876), .ZN(n7877) );
  OAI21_X1 U9614 ( .B1(n7994), .B2(n10247), .A(n7877), .ZN(P2_U3414) );
  INV_X1 U9615 ( .A(n7878), .ZN(n7879) );
  NOR2_X1 U9616 ( .A1(n7885), .A2(n7879), .ZN(n7882) );
  INV_X1 U9617 ( .A(n7880), .ZN(n7881) );
  AOI21_X1 U9618 ( .B1(n7882), .B2(n7744), .A(n7881), .ZN(n10242) );
  NOR2_X1 U9619 ( .A1(n7884), .A2(n7883), .ZN(n7886) );
  XNOR2_X1 U9620 ( .A(n7886), .B(n7885), .ZN(n7887) );
  AOI222_X1 U9621 ( .A1(n10202), .A2(n7887), .B1(n8873), .B2(n10199), .C1(
        n8875), .C2(n9236), .ZN(n10237) );
  MUX2_X1 U9622 ( .A(n7888), .B(n10237), .S(n10212), .Z(n7893) );
  INV_X1 U9623 ( .A(n7889), .ZN(n7890) );
  AOI22_X1 U9624 ( .A1(n9265), .A2(n7891), .B1(n10205), .B2(n7890), .ZN(n7892)
         );
  OAI211_X1 U9625 ( .C1(n10242), .C2(n9268), .A(n7893), .B(n7892), .ZN(
        P2_U3227) );
  MUX2_X1 U9626 ( .A(n7895), .B(n7894), .S(n10257), .Z(n7896) );
  INV_X1 U9627 ( .A(n7896), .ZN(P2_U3466) );
  INV_X1 U9628 ( .A(n7897), .ZN(n7898) );
  AND2_X1 U9629 ( .A1(n7898), .A2(n8192), .ZN(n7901) );
  INV_X1 U9630 ( .A(n7899), .ZN(n7900) );
  NAND2_X1 U9631 ( .A1(n7900), .A2(n7901), .ZN(n8193) );
  OAI21_X1 U9632 ( .B1(n7901), .B2(n7900), .A(n8193), .ZN(n7902) );
  NAND2_X1 U9633 ( .A1(n7902), .A2(n5931), .ZN(n7907) );
  OAI22_X1 U9634 ( .A1(n8030), .A2(n9593), .B1(n8423), .B2(n8398), .ZN(n7920)
         );
  INV_X1 U9635 ( .A(n7920), .ZN(n7904) );
  OAI21_X1 U9636 ( .B1(n7904), .B2(n9558), .A(n7903), .ZN(n7905) );
  AOI21_X1 U9637 ( .B1(n7977), .B2(n9538), .A(n7905), .ZN(n7906) );
  OAI211_X1 U9638 ( .C1(n6478), .C2(n9605), .A(n7907), .B(n7906), .ZN(P1_U3213) );
  INV_X1 U9639 ( .A(n7908), .ZN(n7911) );
  OAI222_X1 U9640 ( .A1(n10115), .A2(n7909), .B1(n10114), .B2(n7911), .C1(
        n8584), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U9641 ( .A1(P2_U3151), .A2(n7912), .B1(n9455), .B2(n7911), .C1(
        n7910), .C2(n9449), .ZN(P2_U3274) );
  INV_X1 U9642 ( .A(n7913), .ZN(n7914) );
  AOI21_X1 U9643 ( .B1(n7657), .B2(n7915), .A(n7914), .ZN(n7917) );
  XNOR2_X1 U9644 ( .A(n7917), .B(n7916), .ZN(n7976) );
  AND2_X1 U9645 ( .A1(n7918), .A2(n8433), .ZN(n7919) );
  NAND2_X1 U9646 ( .A1(n7919), .A2(n8430), .ZN(n7956) );
  OAI21_X1 U9647 ( .B1(n8430), .B2(n7919), .A(n7956), .ZN(n7921) );
  AOI21_X1 U9648 ( .B1(n7921), .B2(n9964), .A(n7920), .ZN(n7985) );
  OAI211_X1 U9649 ( .C1(n6587), .C2(n6478), .A(n9992), .B(n7969), .ZN(n7981)
         );
  OAI211_X1 U9650 ( .C1(n10185), .C2(n7976), .A(n7985), .B(n7981), .ZN(n7927)
         );
  OAI22_X1 U9651 ( .A1(n10036), .A2(n6478), .B1(n10194), .B2(n10454), .ZN(
        n7923) );
  AOI21_X1 U9652 ( .B1(n7927), .B2(n10194), .A(n7923), .ZN(n7924) );
  INV_X1 U9653 ( .A(n7924), .ZN(P1_U3529) );
  INV_X1 U9654 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7925) );
  OAI22_X1 U9655 ( .A1(n10096), .A2(n6478), .B1(n10189), .B2(n7925), .ZN(n7926) );
  AOI21_X1 U9656 ( .B1(n7927), .B2(n10189), .A(n7926), .ZN(n7928) );
  INV_X1 U9657 ( .A(n7928), .ZN(P1_U3474) );
  INV_X1 U9658 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7930) );
  XNOR2_X1 U9659 ( .A(n9684), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7942) );
  NOR2_X1 U9660 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8344), .ZN(n7934) );
  NOR2_X1 U9661 ( .A1(n9745), .A2(n7938), .ZN(n7933) );
  AOI211_X1 U9662 ( .C1(n10122), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7934), .B(
        n7933), .ZN(n7941) );
  NAND2_X1 U9663 ( .A1(n7935), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U9664 ( .A1(n7937), .A2(n7936), .ZN(n9693) );
  XNOR2_X1 U9665 ( .A(n9693), .B(n7938), .ZN(n7939) );
  NAND2_X1 U9666 ( .A1(n7939), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9695) );
  OAI211_X1 U9667 ( .C1(n7939), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9695), .B(
        n10135), .ZN(n7940) );
  OAI211_X1 U9668 ( .C1(n7942), .C2(n10128), .A(n7941), .B(n7940), .ZN(
        P1_U3258) );
  XNOR2_X1 U9669 ( .A(n7943), .B(n6482), .ZN(n7944) );
  AOI22_X1 U9670 ( .A1(n4609), .A2(n9595), .B1(n9567), .B2(n9625), .ZN(n8203)
         );
  OAI21_X1 U9671 ( .B1(n7944), .B2(n9945), .A(n8203), .ZN(n8042) );
  INV_X1 U9672 ( .A(n8042), .ZN(n7954) );
  OAI21_X1 U9673 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n8044) );
  INV_X1 U9674 ( .A(n8170), .ZN(n7949) );
  AOI211_X1 U9675 ( .C1(n8205), .C2(n8035), .A(n9949), .B(n7949), .ZN(n8043)
         );
  NAND2_X1 U9676 ( .A1(n8043), .A2(n9971), .ZN(n7951) );
  AOI22_X1 U9677 ( .A1(n10167), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8200), .B2(
        n10154), .ZN(n7950) );
  OAI211_X1 U9678 ( .C1(n6588), .C2(n9953), .A(n7951), .B(n7950), .ZN(n7952)
         );
  AOI21_X1 U9679 ( .B1(n10163), .B2(n8044), .A(n7952), .ZN(n7953) );
  OAI21_X1 U9680 ( .B1(n7954), .B2(n10167), .A(n7953), .ZN(P1_U3283) );
  AND2_X1 U9681 ( .A1(n7956), .A2(n7955), .ZN(n7958) );
  INV_X1 U9682 ( .A(n7964), .ZN(n7957) );
  NAND2_X1 U9683 ( .A1(n7958), .A2(n7957), .ZN(n8028) );
  OAI211_X1 U9684 ( .C1(n7958), .C2(n7957), .A(n8028), .B(n9964), .ZN(n7963)
         );
  OR2_X1 U9685 ( .A1(n7959), .A2(n9593), .ZN(n7962) );
  OR2_X1 U9686 ( .A1(n7960), .A2(n8398), .ZN(n7961) );
  AND2_X1 U9687 ( .A1(n7962), .A2(n7961), .ZN(n8237) );
  OR2_X1 U9688 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U9689 ( .A1(n7967), .A2(n7966), .ZN(n8135) );
  NAND2_X1 U9690 ( .A1(n7969), .A2(n8142), .ZN(n7970) );
  NAND2_X1 U9691 ( .A1(n7970), .A2(n9992), .ZN(n7971) );
  NOR2_X1 U9692 ( .A1(n7968), .A2(n7971), .ZN(n8134) );
  NAND2_X1 U9693 ( .A1(n8134), .A2(n9971), .ZN(n7973) );
  AOI22_X1 U9694 ( .A1(n10167), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8240), .B2(
        n10154), .ZN(n7972) );
  OAI211_X1 U9695 ( .C1(n8243), .C2(n9953), .A(n7973), .B(n7972), .ZN(n7974)
         );
  AOI21_X1 U9696 ( .B1(n10163), .B2(n8135), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9697 ( .B1(n8137), .B2(n10167), .A(n7975), .ZN(P1_U3285) );
  INV_X1 U9698 ( .A(n7976), .ZN(n7983) );
  AOI22_X1 U9699 ( .A1(n10167), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7977), .B2(
        n10154), .ZN(n7980) );
  NAND2_X1 U9700 ( .A1(n10157), .A2(n7978), .ZN(n7979) );
  OAI211_X1 U9701 ( .C1(n7981), .C2(n10160), .A(n7980), .B(n7979), .ZN(n7982)
         );
  AOI21_X1 U9702 ( .B1(n7983), .B2(n10163), .A(n7982), .ZN(n7984) );
  OAI21_X1 U9703 ( .B1(n7985), .B2(n10167), .A(n7984), .ZN(P1_U3286) );
  INV_X1 U9704 ( .A(n7986), .ZN(n7991) );
  AOI22_X1 U9705 ( .A1(n10167), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9506), .B2(
        n10154), .ZN(n7988) );
  NAND2_X1 U9706 ( .A1(n10157), .A2(n5228), .ZN(n7987) );
  OAI211_X1 U9707 ( .C1(n7989), .C2(n10160), .A(n7988), .B(n7987), .ZN(n7990)
         );
  AOI21_X1 U9708 ( .B1(n7991), .B2(n10163), .A(n7990), .ZN(n7992) );
  OAI21_X1 U9709 ( .B1(n10167), .B2(n7993), .A(n7992), .ZN(P1_U3288) );
  MUX2_X1 U9710 ( .A(n10376), .B(n7994), .S(n10257), .Z(n7995) );
  OAI21_X1 U9711 ( .B1(n8017), .B2(n9317), .A(n7995), .ZN(P2_U3467) );
  OAI21_X1 U9712 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n7999) );
  NAND2_X1 U9713 ( .A1(n7999), .A2(n5931), .ZN(n8006) );
  OAI22_X1 U9714 ( .A1(n8001), .A2(n9593), .B1(n8000), .B2(n8398), .ZN(n9963)
         );
  INV_X1 U9715 ( .A(n9966), .ZN(n8002) );
  NOR2_X1 U9716 ( .A1(n9599), .A2(n8002), .ZN(n8003) );
  AOI211_X1 U9717 ( .C1(n9602), .C2(n9963), .A(n8004), .B(n8003), .ZN(n8005)
         );
  OAI211_X1 U9718 ( .C1(n9969), .C2(n9605), .A(n8006), .B(n8005), .ZN(P1_U3224) );
  XNOR2_X1 U9719 ( .A(n4512), .B(n8050), .ZN(n8051) );
  XNOR2_X1 U9720 ( .A(n8051), .B(n8007), .ZN(n8015) );
  OAI21_X1 U9721 ( .B1(n8848), .B2(n8009), .A(n8008), .ZN(n8010) );
  AOI21_X1 U9722 ( .B1(n8845), .B2(n8871), .A(n8010), .ZN(n8011) );
  OAI21_X1 U9723 ( .B1(n8317), .B2(n8016), .A(n8011), .ZN(n8012) );
  AOI21_X1 U9724 ( .B1(n8013), .B2(n8851), .A(n8012), .ZN(n8014) );
  OAI21_X1 U9725 ( .B1(n8015), .B2(n8853), .A(n8014), .ZN(P2_U3161) );
  INV_X1 U9726 ( .A(n9268), .ZN(n9206) );
  OAI22_X1 U9727 ( .A1(n9204), .A2(n8017), .B1(n8016), .B2(n9240), .ZN(n8020)
         );
  MUX2_X1 U9728 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n8018), .S(n10212), .Z(n8019)
         );
  AOI211_X1 U9729 ( .C1(n9206), .C2(n8021), .A(n8020), .B(n8019), .ZN(n8022)
         );
  INV_X1 U9730 ( .A(n8022), .ZN(P2_U3225) );
  INV_X1 U9731 ( .A(n8023), .ZN(n8027) );
  OAI222_X1 U9732 ( .A1(n9449), .A2(n8025), .B1(n9455), .B2(n8027), .C1(n8024), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9733 ( .A1(n10115), .A2(n10405), .B1(n10114), .B2(n8027), .C1(
        P1_U3086), .C2(n8026), .ZN(P1_U3333) );
  NAND2_X1 U9734 ( .A1(n8028), .A2(n8436), .ZN(n8029) );
  INV_X1 U9735 ( .A(n8033), .ZN(n8542) );
  XNOR2_X1 U9736 ( .A(n8029), .B(n8542), .ZN(n8031) );
  OR2_X1 U9737 ( .A1(n8030), .A2(n8398), .ZN(n8351) );
  OAI21_X1 U9738 ( .B1(n8031), .B2(n9945), .A(n8351), .ZN(n8224) );
  INV_X1 U9739 ( .A(n8224), .ZN(n8041) );
  OAI21_X1 U9740 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8226) );
  OAI211_X1 U9741 ( .C1(n7968), .C2(n4408), .A(n8035), .B(n9992), .ZN(n8036)
         );
  OR2_X1 U9742 ( .A1(n8160), .A2(n9593), .ZN(n8350) );
  NAND2_X1 U9743 ( .A1(n8036), .A2(n8350), .ZN(n8225) );
  NAND2_X1 U9744 ( .A1(n8225), .A2(n9971), .ZN(n8038) );
  AOI22_X1 U9745 ( .A1(n10167), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8349), .B2(
        n10154), .ZN(n8037) );
  OAI211_X1 U9746 ( .C1(n4408), .C2(n9953), .A(n8038), .B(n8037), .ZN(n8039)
         );
  AOI21_X1 U9747 ( .B1(n8226), .B2(n10163), .A(n8039), .ZN(n8040) );
  OAI21_X1 U9748 ( .B1(n8041), .B2(n10167), .A(n8040), .ZN(P1_U3284) );
  INV_X1 U9749 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8045) );
  AOI211_X1 U9750 ( .C1(n10055), .C2(n8044), .A(n8043), .B(n8042), .ZN(n8047)
         );
  MUX2_X1 U9751 ( .A(n8045), .B(n8047), .S(n10189), .Z(n8046) );
  OAI21_X1 U9752 ( .B1(n6588), .B2(n10096), .A(n8046), .ZN(P1_U3483) );
  INV_X1 U9753 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8048) );
  MUX2_X1 U9754 ( .A(n8048), .B(n8047), .S(n10194), .Z(n8049) );
  OAI21_X1 U9755 ( .B1(n6588), .B2(n10036), .A(n8049), .ZN(P1_U3532) );
  OAI22_X1 U9756 ( .A1(n8051), .A2(n8872), .B1(n4512), .B2(n8050), .ZN(n8054)
         );
  XNOR2_X1 U9757 ( .A(n8052), .B(n8096), .ZN(n8053) );
  XNOR2_X1 U9758 ( .A(n8054), .B(n8053), .ZN(n8061) );
  OAI21_X1 U9759 ( .B1(n8861), .B2(n8056), .A(n8055), .ZN(n8057) );
  AOI21_X1 U9760 ( .B1(n8859), .B2(n8872), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9761 ( .B1(n8317), .B2(n8110), .A(n8058), .ZN(n8059) );
  AOI21_X1 U9762 ( .B1(n8109), .B2(n8851), .A(n8059), .ZN(n8060) );
  OAI21_X1 U9763 ( .B1(n8061), .B2(n8853), .A(n8060), .ZN(P2_U3171) );
  NAND2_X1 U9764 ( .A1(n8066), .A2(n8062), .ZN(n8064) );
  OAI211_X1 U9765 ( .C1(n10523), .C2(n9449), .A(n8064), .B(n8063), .ZN(
        P2_U3272) );
  NAND2_X1 U9766 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  OAI211_X1 U9767 ( .C1(n8068), .C2(n10115), .A(n8067), .B(n8570), .ZN(
        P1_U3332) );
  OAI21_X1 U9768 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n8072) );
  NAND2_X1 U9769 ( .A1(n8072), .A2(n5931), .ZN(n8078) );
  OAI22_X1 U9770 ( .A1(n8073), .A2(n9593), .B1(n8161), .B2(n8398), .ZN(n8122)
         );
  INV_X1 U9771 ( .A(n8122), .ZN(n8075) );
  OAI21_X1 U9772 ( .B1(n8075), .B2(n9558), .A(n8074), .ZN(n8076) );
  AOI21_X1 U9773 ( .B1(n8127), .B2(n9538), .A(n8076), .ZN(n8077) );
  OAI211_X1 U9774 ( .C1(n8129), .C2(n9605), .A(n8078), .B(n8077), .ZN(P1_U3234) );
  INV_X1 U9775 ( .A(n8079), .ZN(n8082) );
  INV_X1 U9776 ( .A(n8080), .ZN(n8081) );
  NOR2_X1 U9777 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  XNOR2_X1 U9778 ( .A(n8084), .B(n8083), .ZN(n8090) );
  OAI21_X1 U9779 ( .B1(n8861), .B2(n9258), .A(n8085), .ZN(n8086) );
  AOI21_X1 U9780 ( .B1(n8859), .B2(n8871), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9781 ( .B1(n8317), .B2(n8244), .A(n8087), .ZN(n8088) );
  AOI21_X1 U9782 ( .B1(n8091), .B2(n8851), .A(n8088), .ZN(n8089) );
  OAI21_X1 U9783 ( .B1(n8090), .B2(n8853), .A(n8089), .ZN(P2_U3157) );
  INV_X1 U9784 ( .A(n8091), .ZN(n8245) );
  INV_X1 U9785 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U9786 ( .A1(n8108), .A2(n8092), .ZN(n8093) );
  XNOR2_X1 U9787 ( .A(n8093), .B(n8094), .ZN(n8249) );
  XOR2_X1 U9788 ( .A(n8095), .B(n8094), .Z(n8100) );
  OAI22_X1 U9789 ( .A1(n8096), .A2(n9259), .B1(n9258), .B2(n9261), .ZN(n8097)
         );
  AOI21_X1 U9790 ( .B1(n8249), .B2(n8098), .A(n8097), .ZN(n8099) );
  OAI21_X1 U9791 ( .B1(n8100), .B2(n9256), .A(n8099), .ZN(n8246) );
  AOI21_X1 U9792 ( .B1(n10235), .B2(n8249), .A(n8246), .ZN(n8103) );
  MUX2_X1 U9793 ( .A(n8101), .B(n8103), .S(n10245), .Z(n8102) );
  OAI21_X1 U9794 ( .B1(n8245), .B2(n9413), .A(n8102), .ZN(P2_U3420) );
  MUX2_X1 U9795 ( .A(n8104), .B(n8103), .S(n10257), .Z(n8105) );
  OAI21_X1 U9796 ( .B1(n8245), .B2(n9317), .A(n8105), .ZN(P2_U3469) );
  OR2_X1 U9797 ( .A1(n8106), .A2(n8111), .ZN(n8107) );
  NAND2_X1 U9798 ( .A1(n8108), .A2(n8107), .ZN(n9335) );
  INV_X1 U9799 ( .A(n9335), .ZN(n8118) );
  INV_X1 U9800 ( .A(n8109), .ZN(n9333) );
  OAI22_X1 U9801 ( .A1(n9204), .A2(n9333), .B1(n8110), .B2(n9240), .ZN(n8117)
         );
  XNOR2_X1 U9802 ( .A(n4544), .B(n8111), .ZN(n8113) );
  NAND2_X1 U9803 ( .A1(n8113), .A2(n10202), .ZN(n8115) );
  AOI22_X1 U9804 ( .A1(n9236), .A2(n8872), .B1(n8870), .B2(n10199), .ZN(n8114)
         );
  OAI211_X1 U9805 ( .C1(n10207), .C2(n9335), .A(n8115), .B(n8114), .ZN(n9337)
         );
  MUX2_X1 U9806 ( .A(n9337), .B(P2_REG2_REG_9__SCAN_IN), .S(n9246), .Z(n8116)
         );
  AOI211_X1 U9807 ( .C1(n8118), .C2(n10209), .A(n8117), .B(n8116), .ZN(n8119)
         );
  INV_X1 U9808 ( .A(n8119), .ZN(P2_U3224) );
  OAI21_X1 U9809 ( .B1(n8121), .B2(n8547), .A(n8120), .ZN(n8123) );
  AOI21_X1 U9810 ( .B1(n8123), .B2(n9964), .A(n8122), .ZN(n10051) );
  INV_X1 U9811 ( .A(n8124), .ZN(n8126) );
  AOI211_X1 U9812 ( .C1(n10049), .C2(n8126), .A(n9949), .B(n4572), .ZN(n10048)
         );
  AOI22_X1 U9813 ( .A1(n10167), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8127), .B2(
        n10154), .ZN(n8128) );
  OAI21_X1 U9814 ( .B1(n8129), .B2(n9953), .A(n8128), .ZN(n8132) );
  XOR2_X1 U9815 ( .A(n8130), .B(n8547), .Z(n10052) );
  NOR2_X1 U9816 ( .A1(n10052), .A2(n9957), .ZN(n8131) );
  AOI211_X1 U9817 ( .C1(n10048), .C2(n9971), .A(n8132), .B(n8131), .ZN(n8133)
         );
  OAI21_X1 U9818 ( .B1(n10167), .B2(n10051), .A(n8133), .ZN(P1_U3280) );
  INV_X1 U9819 ( .A(n10096), .ZN(n8701) );
  AOI21_X1 U9820 ( .B1(n8135), .B2(n10055), .A(n8134), .ZN(n8136) );
  NAND2_X1 U9821 ( .A1(n8137), .A2(n8136), .ZN(n8140) );
  MUX2_X1 U9822 ( .A(n8140), .B(P1_REG0_REG_8__SCAN_IN), .S(n10187), .Z(n8138)
         );
  AOI21_X1 U9823 ( .B1(n8701), .B2(n8142), .A(n8138), .ZN(n8139) );
  INV_X1 U9824 ( .A(n8139), .ZN(P1_U3477) );
  INV_X1 U9825 ( .A(n10036), .ZN(n8394) );
  MUX2_X1 U9826 ( .A(n8140), .B(P1_REG1_REG_8__SCAN_IN), .S(n10192), .Z(n8141)
         );
  AOI21_X1 U9827 ( .B1(n8394), .B2(n8142), .A(n8141), .ZN(n8143) );
  INV_X1 U9828 ( .A(n8143), .ZN(P1_U3530) );
  OAI21_X1 U9829 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n4428), .A(n7129), .ZN(
        n8145) );
  OAI21_X1 U9830 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n4502), .A(n7122), .ZN(
        n8144) );
  AOI22_X1 U9831 ( .A1(n9006), .A2(n8145), .B1(n8144), .B2(n8886), .ZN(n8157)
         );
  INV_X1 U9832 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U9833 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8316) );
  OAI21_X1 U9834 ( .B1(n9020), .B2(n10286), .A(n8316), .ZN(n8154) );
  INV_X1 U9835 ( .A(n8146), .ZN(n8147) );
  NAND3_X1 U9836 ( .A1(n8149), .A2(n8148), .A3(n8147), .ZN(n8151) );
  AOI21_X1 U9837 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8153) );
  AOI211_X1 U9838 ( .C1(n8991), .C2(n8155), .A(n8154), .B(n8153), .ZN(n8156)
         );
  NAND2_X1 U9839 ( .A1(n8157), .A2(n8156), .ZN(P2_U3195) );
  XNOR2_X1 U9840 ( .A(n8158), .B(n8544), .ZN(n8169) );
  INV_X1 U9841 ( .A(n8169), .ZN(n10065) );
  INV_X1 U9842 ( .A(n8159), .ZN(n8257) );
  OR2_X1 U9843 ( .A1(n8160), .A2(n8398), .ZN(n8163) );
  OR2_X1 U9844 ( .A1(n8161), .A2(n9593), .ZN(n8162) );
  NAND2_X1 U9845 ( .A1(n8163), .A2(n8162), .ZN(n8305) );
  NAND2_X1 U9846 ( .A1(n8164), .A2(n8450), .ZN(n8167) );
  INV_X1 U9847 ( .A(n8165), .ZN(n8166) );
  AOI211_X1 U9848 ( .C1(n8544), .C2(n8167), .A(n9945), .B(n8166), .ZN(n8168)
         );
  AOI211_X1 U9849 ( .C1(n8257), .C2(n8169), .A(n8305), .B(n8168), .ZN(n10064)
         );
  MUX2_X1 U9850 ( .A(n7424), .B(n10064), .S(n9951), .Z(n8175) );
  AOI211_X1 U9851 ( .C1(n10062), .C2(n8170), .A(n9949), .B(n4503), .ZN(n10061)
         );
  INV_X1 U9852 ( .A(n10062), .ZN(n8172) );
  INV_X1 U9853 ( .A(n8171), .ZN(n8307) );
  OAI22_X1 U9854 ( .A1(n8172), .A2(n9953), .B1(n9913), .B2(n8307), .ZN(n8173)
         );
  AOI21_X1 U9855 ( .B1(n10061), .B2(n9971), .A(n8173), .ZN(n8174) );
  OAI211_X1 U9856 ( .C1(n10065), .C2(n8268), .A(n8175), .B(n8174), .ZN(
        P1_U3282) );
  XNOR2_X1 U9857 ( .A(n8176), .B(n8178), .ZN(n8191) );
  NAND2_X1 U9858 ( .A1(n9252), .A2(n8177), .ZN(n8179) );
  XNOR2_X1 U9859 ( .A(n8179), .B(n8178), .ZN(n8180) );
  AOI222_X1 U9860 ( .A1(n10202), .A2(n8180), .B1(n9237), .B2(n10199), .C1(
        n8870), .C2(n9236), .ZN(n8185) );
  MUX2_X1 U9861 ( .A(n10564), .B(n8185), .S(n10245), .Z(n8182) );
  NAND2_X1 U9862 ( .A1(n6946), .A2(n8188), .ZN(n8181) );
  OAI211_X1 U9863 ( .C1(n8191), .C2(n9435), .A(n8182), .B(n8181), .ZN(P2_U3423) );
  MUX2_X1 U9864 ( .A(n4811), .B(n8185), .S(n10257), .Z(n8184) );
  NAND2_X1 U9865 ( .A1(n8188), .A2(n6963), .ZN(n8183) );
  OAI211_X1 U9866 ( .C1(n8191), .C2(n9332), .A(n8184), .B(n8183), .ZN(P2_U3470) );
  MUX2_X1 U9867 ( .A(n8186), .B(n8185), .S(n10212), .Z(n8190) );
  INV_X1 U9868 ( .A(n8187), .ZN(n8214) );
  AOI22_X1 U9869 ( .A1(n8188), .A2(n9265), .B1(n10205), .B2(n8214), .ZN(n8189)
         );
  OAI211_X1 U9870 ( .C1(n8191), .C2(n9268), .A(n8190), .B(n8189), .ZN(P2_U3222) );
  NAND2_X1 U9871 ( .A1(n8193), .A2(n8192), .ZN(n8231) );
  INV_X1 U9872 ( .A(n8194), .ZN(n8195) );
  NAND2_X1 U9873 ( .A1(n8231), .A2(n8195), .ZN(n8197) );
  AOI21_X1 U9874 ( .B1(n8197), .B2(n8196), .A(n8359), .ZN(n8302) );
  XNOR2_X1 U9875 ( .A(n8302), .B(n8301), .ZN(n8198) );
  NOR2_X1 U9876 ( .A1(n8198), .A2(n8199), .ZN(n8300) );
  AOI21_X1 U9877 ( .B1(n8199), .B2(n8198), .A(n8300), .ZN(n8207) );
  NAND2_X1 U9878 ( .A1(n9538), .A2(n8200), .ZN(n8201) );
  OAI211_X1 U9879 ( .C1(n8203), .C2(n9558), .A(n8202), .B(n8201), .ZN(n8204)
         );
  AOI21_X1 U9880 ( .B1(n8205), .B2(n4405), .A(n8204), .ZN(n8206) );
  OAI21_X1 U9881 ( .B1(n8207), .B2(n9589), .A(n8206), .ZN(P1_U3217) );
  NOR2_X1 U9882 ( .A1(n8208), .A2(n8287), .ZN(n8286) );
  INV_X1 U9883 ( .A(n8286), .ZN(n8209) );
  OAI211_X1 U9884 ( .C1(n8210), .C2(n6199), .A(n8209), .B(n8855), .ZN(n8216)
         );
  NAND2_X1 U9885 ( .A1(n8859), .A2(n8870), .ZN(n8212) );
  OAI211_X1 U9886 ( .C1(n8284), .C2(n8861), .A(n8212), .B(n8211), .ZN(n8213)
         );
  AOI21_X1 U9887 ( .B1(n8863), .B2(n8214), .A(n8213), .ZN(n8215) );
  OAI211_X1 U9888 ( .C1(n8217), .C2(n8866), .A(n8216), .B(n8215), .ZN(P2_U3176) );
  INV_X1 U9889 ( .A(n8218), .ZN(n8222) );
  OAI222_X1 U9890 ( .A1(P1_U3086), .A2(n8220), .B1(n10114), .B2(n8222), .C1(
        n8219), .C2(n10115), .ZN(P1_U3331) );
  OAI222_X1 U9891 ( .A1(n8223), .A2(P2_U3151), .B1(n9455), .B2(n8222), .C1(
        n8221), .C2(n9449), .ZN(P2_U3271) );
  INV_X1 U9892 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10471) );
  AOI211_X1 U9893 ( .C1(n10055), .C2(n8226), .A(n8225), .B(n8224), .ZN(n8228)
         );
  MUX2_X1 U9894 ( .A(n10471), .B(n8228), .S(n10189), .Z(n8227) );
  OAI21_X1 U9895 ( .B1(n4408), .B2(n10096), .A(n8227), .ZN(P1_U3480) );
  INV_X1 U9896 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8229) );
  MUX2_X1 U9897 ( .A(n8229), .B(n8228), .S(n10194), .Z(n8230) );
  OAI21_X1 U9898 ( .B1(n4408), .B2(n10036), .A(n8230), .ZN(P1_U3531) );
  INV_X1 U9899 ( .A(n8231), .ZN(n8233) );
  NOR2_X1 U9900 ( .A1(n8233), .A2(n8232), .ZN(n8356) );
  AOI21_X1 U9901 ( .B1(n8233), .B2(n8232), .A(n8356), .ZN(n8234) );
  NAND2_X1 U9902 ( .A1(n8234), .A2(n8235), .ZN(n8358) );
  OAI21_X1 U9903 ( .B1(n8235), .B2(n8234), .A(n8358), .ZN(n8236) );
  NAND2_X1 U9904 ( .A1(n8236), .A2(n5931), .ZN(n8242) );
  NOR2_X1 U9905 ( .A1(n8237), .A2(n9558), .ZN(n8238) );
  AOI211_X1 U9906 ( .C1(n9538), .C2(n8240), .A(n8239), .B(n8238), .ZN(n8241)
         );
  OAI211_X1 U9907 ( .C1(n8243), .C2(n9605), .A(n8242), .B(n8241), .ZN(P1_U3221) );
  OAI22_X1 U9908 ( .A1(n8245), .A2(n9204), .B1(n8244), .B2(n9240), .ZN(n8248)
         );
  MUX2_X1 U9909 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8246), .S(n10212), .Z(n8247) );
  AOI211_X1 U9910 ( .C1(n8249), .C2(n10209), .A(n8248), .B(n8247), .ZN(n8250)
         );
  INV_X1 U9911 ( .A(n8250), .ZN(P2_U3223) );
  XNOR2_X1 U9912 ( .A(n8251), .B(n8252), .ZN(n8258) );
  INV_X1 U9913 ( .A(n8258), .ZN(n10045) );
  NAND2_X1 U9914 ( .A1(n8120), .A2(n8612), .ZN(n8253) );
  XNOR2_X1 U9915 ( .A(n8253), .B(n8252), .ZN(n8254) );
  NAND2_X1 U9916 ( .A1(n8254), .A2(n9964), .ZN(n8260) );
  NAND2_X1 U9917 ( .A1(n9621), .A2(n9567), .ZN(n8256) );
  NAND2_X1 U9918 ( .A1(n9623), .A2(n9595), .ZN(n8255) );
  NAND2_X1 U9919 ( .A1(n8256), .A2(n8255), .ZN(n8322) );
  AOI21_X1 U9920 ( .B1(n8258), .B2(n8257), .A(n8322), .ZN(n8259) );
  NAND2_X1 U9921 ( .A1(n8260), .A2(n8259), .ZN(n10047) );
  NAND2_X1 U9922 ( .A1(n10047), .A2(n9951), .ZN(n8267) );
  INV_X1 U9923 ( .A(n8261), .ZN(n8324) );
  OAI22_X1 U9924 ( .A1(n9951), .A2(n8262), .B1(n8324), .B2(n9913), .ZN(n8265)
         );
  AOI21_X1 U9925 ( .B1(n8125), .B2(n10042), .A(n9949), .ZN(n8263) );
  NAND2_X1 U9926 ( .A1(n8263), .A2(n9950), .ZN(n10043) );
  NOR2_X1 U9927 ( .A1(n10043), .A2(n10160), .ZN(n8264) );
  AOI211_X1 U9928 ( .C1(n10157), .C2(n10042), .A(n8265), .B(n8264), .ZN(n8266)
         );
  OAI211_X1 U9929 ( .C1(n10045), .C2(n8268), .A(n8267), .B(n8266), .ZN(
        P1_U3279) );
  INV_X1 U9930 ( .A(n8269), .ZN(n8273) );
  OAI222_X1 U9931 ( .A1(n8271), .A2(P2_U3151), .B1(n9455), .B2(n8273), .C1(
        n8270), .C2(n9449), .ZN(P2_U3270) );
  OAI222_X1 U9932 ( .A1(P1_U3086), .A2(n8274), .B1(n10114), .B2(n8273), .C1(
        n8272), .C2(n10115), .ZN(P1_U3330) );
  AOI21_X1 U9933 ( .B1(n8277), .B2(n8276), .A(n8275), .ZN(n8283) );
  NAND2_X1 U9934 ( .A1(n8863), .A2(n9230), .ZN(n8280) );
  AOI21_X1 U9935 ( .B1(n8845), .B2(n9226), .A(n8278), .ZN(n8279) );
  OAI211_X1 U9936 ( .C1(n9260), .C2(n8848), .A(n8280), .B(n8279), .ZN(n8281)
         );
  AOI21_X1 U9937 ( .B1(n9423), .B2(n8851), .A(n8281), .ZN(n8282) );
  OAI21_X1 U9938 ( .B1(n8283), .B2(n8853), .A(n8282), .ZN(P2_U3155) );
  INV_X1 U9939 ( .A(n9328), .ZN(n8296) );
  XNOR2_X1 U9940 ( .A(n8285), .B(n8284), .ZN(n8289) );
  AOI21_X1 U9941 ( .B1(n8869), .B2(n8287), .A(n8286), .ZN(n8288) );
  NAND2_X1 U9942 ( .A1(n8288), .A2(n8289), .ZN(n8312) );
  OAI21_X1 U9943 ( .B1(n8289), .B2(n8288), .A(n8312), .ZN(n8290) );
  NAND2_X1 U9944 ( .A1(n8290), .A2(n8855), .ZN(n8295) );
  INV_X1 U9945 ( .A(n8291), .ZN(n9264) );
  AOI22_X1 U9946 ( .A1(n8845), .A2(n9225), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3151), .ZN(n8292) );
  OAI21_X1 U9947 ( .B1(n9258), .B2(n8848), .A(n8292), .ZN(n8293) );
  AOI21_X1 U9948 ( .B1(n9264), .B2(n8863), .A(n8293), .ZN(n8294) );
  OAI211_X1 U9949 ( .C1(n8296), .C2(n8866), .A(n8295), .B(n8294), .ZN(P2_U3164) );
  OAI21_X1 U9950 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8304) );
  AOI21_X1 U9951 ( .B1(n8302), .B2(n8301), .A(n8300), .ZN(n8303) );
  XOR2_X1 U9952 ( .A(n8304), .B(n8303), .Z(n8310) );
  AOI22_X1 U9953 ( .A1(n8305), .A2(n9602), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8306) );
  OAI21_X1 U9954 ( .B1(n8307), .B2(n9599), .A(n8306), .ZN(n8308) );
  AOI21_X1 U9955 ( .B1(n10062), .B2(n4405), .A(n8308), .ZN(n8309) );
  OAI21_X1 U9956 ( .B1(n8310), .B2(n9589), .A(n8309), .ZN(P1_U3236) );
  INV_X1 U9957 ( .A(n9428), .ZN(n9243) );
  AND2_X1 U9958 ( .A1(n8312), .A2(n8311), .ZN(n8315) );
  OAI211_X1 U9959 ( .C1(n8315), .C2(n8314), .A(n8855), .B(n8313), .ZN(n8321)
         );
  OAI21_X1 U9960 ( .B1(n8861), .B2(n9213), .A(n8316), .ZN(n8319) );
  NOR2_X1 U9961 ( .A1(n8317), .A2(n9241), .ZN(n8318) );
  AOI211_X1 U9962 ( .C1(n8859), .C2(n9237), .A(n8319), .B(n8318), .ZN(n8320)
         );
  OAI211_X1 U9963 ( .C1(n9243), .C2(n8866), .A(n8321), .B(n8320), .ZN(P2_U3174) );
  AOI22_X1 U9964 ( .A1(n9602), .A2(n8322), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8323) );
  OAI21_X1 U9965 ( .B1(n8324), .B2(n9599), .A(n8323), .ZN(n8330) );
  INV_X1 U9966 ( .A(n8325), .ZN(n8326) );
  AOI211_X1 U9967 ( .C1(n8328), .C2(n8327), .A(n9589), .B(n8326), .ZN(n8329)
         );
  AOI211_X1 U9968 ( .C1(n10042), .C2(n4405), .A(n8330), .B(n8329), .ZN(n8331)
         );
  INV_X1 U9969 ( .A(n8331), .ZN(P1_U3215) );
  INV_X1 U9970 ( .A(n8332), .ZN(n8335) );
  OAI222_X1 U9971 ( .A1(n6408), .A2(P2_U3151), .B1(n9455), .B2(n8335), .C1(
        n8333), .C2(n9449), .ZN(P2_U3269) );
  OAI222_X1 U9972 ( .A1(P1_U3086), .A2(n8336), .B1(n10114), .B2(n8335), .C1(
        n8334), .C2(n10115), .ZN(P1_U3329) );
  NAND2_X1 U9973 ( .A1(n8338), .A2(n8337), .ZN(n8340) );
  XOR2_X1 U9974 ( .A(n8340), .B(n8339), .Z(n8348) );
  OR2_X1 U9975 ( .A1(n8341), .A2(n9593), .ZN(n8343) );
  NAND2_X1 U9976 ( .A1(n9622), .A2(n9595), .ZN(n8342) );
  AND2_X1 U9977 ( .A1(n8343), .A2(n8342), .ZN(n9944) );
  OAI22_X1 U9978 ( .A1(n9944), .A2(n9558), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8344), .ZN(n8346) );
  NOR2_X1 U9979 ( .A1(n9954), .A2(n9605), .ZN(n8345) );
  AOI211_X1 U9980 ( .C1(n9538), .C2(n9947), .A(n8346), .B(n8345), .ZN(n8347)
         );
  OAI21_X1 U9981 ( .B1(n8348), .B2(n9589), .A(n8347), .ZN(P1_U3241) );
  INV_X1 U9982 ( .A(n8349), .ZN(n8355) );
  NAND2_X1 U9983 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U9984 ( .A1(n8352), .A2(n9602), .ZN(n8354) );
  OAI211_X1 U9985 ( .C1(n9599), .C2(n8355), .A(n8354), .B(n8353), .ZN(n8366)
         );
  INV_X1 U9986 ( .A(n8356), .ZN(n8357) );
  NAND2_X1 U9987 ( .A1(n8358), .A2(n8357), .ZN(n8363) );
  INV_X1 U9988 ( .A(n8359), .ZN(n8361) );
  NAND2_X1 U9989 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  XNOR2_X1 U9990 ( .A(n8363), .B(n8362), .ZN(n8364) );
  NOR2_X1 U9991 ( .A1(n8364), .A2(n9589), .ZN(n8365) );
  AOI211_X1 U9992 ( .C1(n8367), .C2(n4405), .A(n8366), .B(n8365), .ZN(n8368)
         );
  INV_X1 U9993 ( .A(n8368), .ZN(P1_U3231) );
  OAI222_X1 U9994 ( .A1(n10115), .A2(n8370), .B1(n10114), .B2(n8369), .C1(
        P1_U3086), .C2(n8526), .ZN(P1_U3336) );
  INV_X1 U9995 ( .A(n9386), .ZN(n8378) );
  OAI211_X1 U9996 ( .C1(n8373), .C2(n8372), .A(n8371), .B(n8855), .ZN(n8377)
         );
  AOI22_X1 U9997 ( .A1(n9108), .A2(n8859), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8374) );
  OAI21_X1 U9998 ( .B1(n8817), .B2(n8861), .A(n8374), .ZN(n8375) );
  AOI21_X1 U9999 ( .B1(n9112), .B2(n8863), .A(n8375), .ZN(n8376) );
  OAI211_X1 U10000 ( .C1(n8378), .C2(n8866), .A(n8377), .B(n8376), .ZN(
        P2_U3175) );
  INV_X1 U10001 ( .A(n8382), .ZN(n8379) );
  NOR2_X1 U10002 ( .A1(n8380), .A2(n8379), .ZN(n8385) );
  AOI21_X1 U10003 ( .B1(n8383), .B2(n8382), .A(n8381), .ZN(n8384) );
  OAI21_X1 U10004 ( .B1(n8385), .B2(n8384), .A(n5931), .ZN(n8389) );
  AOI22_X1 U10005 ( .A1(n8387), .A2(n9602), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8386), .ZN(n8388) );
  OAI211_X1 U10006 ( .C1(n10173), .C2(n9605), .A(n8389), .B(n8388), .ZN(
        P1_U3222) );
  XNOR2_X1 U10007 ( .A(n8390), .B(n9760), .ZN(n8391) );
  INV_X1 U10008 ( .A(n9752), .ZN(n8392) );
  NAND2_X1 U10009 ( .A1(n9762), .A2(n8392), .ZN(n8699) );
  MUX2_X1 U10010 ( .A(n8699), .B(P1_REG1_REG_30__SCAN_IN), .S(n10192), .Z(
        n8393) );
  AOI21_X1 U10011 ( .B1(n8394), .B2(n9760), .A(n8393), .ZN(n8395) );
  INV_X1 U10012 ( .A(n8395), .ZN(P1_U3552) );
  XOR2_X1 U10013 ( .A(n8396), .B(n8555), .Z(n10021) );
  XNOR2_X1 U10014 ( .A(n8397), .B(n8555), .ZN(n8401) );
  OAI22_X1 U10015 ( .A1(n8400), .A2(n9593), .B1(n8399), .B2(n8398), .ZN(n9471)
         );
  AOI21_X1 U10016 ( .B1(n8401), .B2(n9964), .A(n9471), .ZN(n10020) );
  OAI22_X1 U10017 ( .A1(n9951), .A2(n8402), .B1(n9473), .B2(n9913), .ZN(n8403)
         );
  AOI21_X1 U10018 ( .B1(n10018), .B2(n10157), .A(n8403), .ZN(n8407) );
  NAND2_X1 U10019 ( .A1(n9899), .A2(n10018), .ZN(n8404) );
  NAND2_X1 U10020 ( .A1(n8404), .A2(n9992), .ZN(n8405) );
  NOR2_X1 U10021 ( .A1(n9887), .A2(n8405), .ZN(n10017) );
  NAND2_X1 U10022 ( .A1(n10017), .A2(n9971), .ZN(n8406) );
  OAI211_X1 U10023 ( .C1(n10020), .C2(n10167), .A(n8407), .B(n8406), .ZN(n8408) );
  INV_X1 U10024 ( .A(n8408), .ZN(n8409) );
  OAI21_X1 U10025 ( .B1(n10021), .B2(n9957), .A(n8409), .ZN(P1_U3274) );
  NAND2_X1 U10026 ( .A1(n8519), .A2(n8664), .ZN(n8670) );
  INV_X1 U10027 ( .A(n8670), .ZN(n8522) );
  OAI21_X1 U10028 ( .B1(n10039), .B2(n8518), .A(n8410), .ZN(n8469) );
  INV_X1 U10029 ( .A(n8619), .ZN(n8461) );
  OAI21_X1 U10030 ( .B1(n8461), .B2(n8411), .A(n8521), .ZN(n8468) );
  NAND2_X1 U10031 ( .A1(n8592), .A2(n8412), .ZN(n8413) );
  AOI21_X1 U10032 ( .B1(n7641), .B2(n8589), .A(n8413), .ZN(n8415) );
  INV_X1 U10033 ( .A(n8414), .ZN(n8590) );
  AND3_X1 U10034 ( .A1(n8598), .A2(n8600), .A3(n8518), .ZN(n8416) );
  NAND2_X1 U10035 ( .A1(n8417), .A2(n8521), .ZN(n8426) );
  OAI21_X1 U10036 ( .B1(n8426), .B2(n9629), .A(n5228), .ZN(n8422) );
  OR2_X1 U10037 ( .A1(n8417), .A2(n8521), .ZN(n8418) );
  OAI21_X1 U10038 ( .B1(n8418), .B2(n8423), .A(n8425), .ZN(n8421) );
  OAI22_X1 U10039 ( .A1(n8418), .A2(n5228), .B1(n8423), .B2(n8521), .ZN(n8420)
         );
  AOI22_X1 U10040 ( .A1(n8422), .A2(n8421), .B1(n8420), .B2(n8419), .ZN(n8429)
         );
  NAND2_X1 U10041 ( .A1(n8423), .A2(n8521), .ZN(n8424) );
  OAI21_X1 U10042 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8427) );
  NAND2_X1 U10043 ( .A1(n8427), .A2(n10145), .ZN(n8428) );
  NAND4_X1 U10044 ( .A1(n8431), .A2(n8430), .A3(n8429), .A4(n8428), .ZN(n8440)
         );
  INV_X1 U10045 ( .A(n8432), .ZN(n8435) );
  NAND4_X1 U10046 ( .A1(n8593), .A2(n8433), .A3(n8597), .A4(n8521), .ZN(n8434)
         );
  AND2_X1 U10047 ( .A1(n8437), .A2(n8436), .ZN(n8538) );
  MUX2_X1 U10048 ( .A(n8538), .B(n8596), .S(n8518), .Z(n8438) );
  MUX2_X1 U10049 ( .A(n8442), .B(n8441), .S(n8518), .Z(n8443) );
  NAND3_X1 U10050 ( .A1(n8446), .A2(n8451), .A3(n8613), .ZN(n8447) );
  NAND2_X1 U10051 ( .A1(n8447), .A2(n8454), .ZN(n8457) );
  INV_X1 U10052 ( .A(n8448), .ZN(n8449) );
  NAND2_X1 U10053 ( .A1(n8449), .A2(n8602), .ZN(n8452) );
  NAND2_X1 U10054 ( .A1(n8451), .A2(n8450), .ZN(n8609) );
  AOI21_X1 U10055 ( .B1(n8452), .B2(n8605), .A(n8609), .ZN(n8455) );
  NAND2_X1 U10056 ( .A1(n8454), .A2(n8453), .ZN(n8614) );
  OAI21_X1 U10057 ( .B1(n8455), .B2(n8614), .A(n8613), .ZN(n8456) );
  AND2_X1 U10058 ( .A1(n8465), .A2(n8458), .ZN(n8617) );
  INV_X1 U10059 ( .A(n8459), .ZN(n8460) );
  OR2_X1 U10060 ( .A1(n9929), .A2(n8460), .ZN(n8616) );
  INV_X1 U10061 ( .A(n8462), .ZN(n8467) );
  INV_X1 U10062 ( .A(n8463), .ZN(n8464) );
  NAND2_X1 U10063 ( .A1(n8475), .A2(n8470), .ZN(n9919) );
  AND2_X1 U10064 ( .A1(n8477), .A2(n8470), .ZN(n8551) );
  NAND2_X1 U10065 ( .A1(n8479), .A2(n8476), .ZN(n8626) );
  AOI21_X1 U10066 ( .B1(n8471), .B2(n8551), .A(n8626), .ZN(n8474) );
  NAND4_X1 U10067 ( .A1(n8472), .A2(n9865), .A3(n8625), .A4(n8518), .ZN(n8473)
         );
  NAND2_X1 U10068 ( .A1(n8476), .A2(n8475), .ZN(n8583) );
  OAI211_X1 U10069 ( .C1(n8478), .C2(n8583), .A(n8625), .B(n8477), .ZN(n8482)
         );
  AND4_X1 U10070 ( .A1(n8480), .A2(n8521), .A3(n8479), .A4(n8486), .ZN(n8481)
         );
  NAND2_X1 U10071 ( .A1(n8490), .A2(n8634), .ZN(n9854) );
  INV_X1 U10072 ( .A(n9876), .ZN(n10085) );
  AOI211_X1 U10073 ( .C1(n9615), .C2(n9865), .A(n8518), .B(n10085), .ZN(n8489)
         );
  AOI211_X1 U10074 ( .C1(n8483), .C2(n8486), .A(n8521), .B(n9876), .ZN(n8488)
         );
  NAND2_X1 U10075 ( .A1(n9615), .A2(n8518), .ZN(n8485) );
  OR2_X1 U10076 ( .A1(n9615), .A2(n8518), .ZN(n8484) );
  OAI22_X1 U10077 ( .A1(n8486), .A2(n8485), .B1(n9865), .B2(n8484), .ZN(n8487)
         );
  NAND2_X1 U10078 ( .A1(n8494), .A2(n8490), .ZN(n8575) );
  NAND2_X1 U10079 ( .A1(n8635), .A2(n8634), .ZN(n8491) );
  MUX2_X1 U10080 ( .A(n8575), .B(n8491), .S(n8518), .Z(n8492) );
  INV_X1 U10081 ( .A(n8492), .ZN(n8493) );
  MUX2_X1 U10082 ( .A(n8635), .B(n8494), .S(n8518), .Z(n8495) );
  NAND2_X1 U10083 ( .A1(n8655), .A2(n8637), .ZN(n8499) );
  NAND2_X1 U10084 ( .A1(n9801), .A2(n9610), .ZN(n8500) );
  MUX2_X1 U10085 ( .A(n8636), .B(n8576), .S(n8518), .Z(n8496) );
  NAND3_X1 U10086 ( .A1(n8500), .A2(n8580), .A3(n8496), .ZN(n8497) );
  INV_X1 U10087 ( .A(n8499), .ZN(n8507) );
  INV_X1 U10088 ( .A(n8500), .ZN(n8631) );
  AOI21_X1 U10089 ( .B1(n8507), .B2(n5007), .A(n8631), .ZN(n8501) );
  OAI21_X1 U10090 ( .B1(n8501), .B2(n8518), .A(n8630), .ZN(n8504) );
  AND2_X1 U10091 ( .A1(n8503), .A2(n8502), .ZN(n8506) );
  OAI21_X1 U10092 ( .B1(n8505), .B2(n8504), .A(n8506), .ZN(n8512) );
  INV_X1 U10093 ( .A(n8506), .ZN(n8640) );
  NOR3_X1 U10094 ( .A1(n8507), .A2(n8631), .A3(n8521), .ZN(n8509) );
  INV_X1 U10095 ( .A(n8573), .ZN(n8508) );
  AOI211_X1 U10096 ( .C1(n8518), .C2(n8640), .A(n8509), .B(n8508), .ZN(n8511)
         );
  OAI21_X1 U10097 ( .B1(n8640), .B2(n8630), .A(n8573), .ZN(n8510) );
  AOI22_X1 U10098 ( .A1(n8512), .A2(n8511), .B1(n8518), .B2(n8510), .ZN(n8514)
         );
  INV_X1 U10099 ( .A(n8559), .ZN(n9606) );
  AOI21_X1 U10100 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8684) );
  INV_X1 U10101 ( .A(n8570), .ZN(n8525) );
  NOR2_X1 U10102 ( .A1(n8523), .A2(n5224), .ZN(n8524) );
  OAI211_X1 U10103 ( .C1(n8667), .C2(n8526), .A(n8525), .B(n8524), .ZN(n8683)
         );
  AOI21_X1 U10104 ( .B1(n8527), .B2(n5224), .A(n8584), .ZN(n8565) );
  INV_X1 U10105 ( .A(n8528), .ZN(n8530) );
  INV_X1 U10106 ( .A(n8531), .ZN(n8532) );
  INV_X1 U10107 ( .A(n7636), .ZN(n8533) );
  NAND4_X1 U10108 ( .A1(n8534), .A2(n4409), .A3(n8533), .A4(n8584), .ZN(n8537)
         );
  INV_X1 U10109 ( .A(n8538), .ZN(n8539) );
  NAND4_X1 U10110 ( .A1(n8543), .A2(n6482), .A3(n8596), .A4(n8542), .ZN(n8545)
         );
  NOR2_X1 U10111 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  OR3_X1 U10112 ( .A1(n9955), .A2(n8549), .A3(n8548), .ZN(n8550) );
  INV_X1 U10113 ( .A(n8551), .ZN(n8622) );
  NAND4_X1 U10114 ( .A1(n9871), .A2(n8555), .A3(n8554), .A4(n9883), .ZN(n8556)
         );
  NOR2_X1 U10115 ( .A1(n8556), .A2(n9854), .ZN(n8557) );
  NOR4_X1 U10116 ( .A1(n8687), .A2(n9795), .A3(n9786), .A4(n8558), .ZN(n8560)
         );
  NAND2_X1 U10117 ( .A1(n9760), .A2(n8559), .ZN(n8645) );
  NAND4_X1 U10118 ( .A1(n8667), .A2(n8561), .A3(n8560), .A4(n8645), .ZN(n8562)
         );
  NAND2_X1 U10119 ( .A1(n6608), .A2(n9606), .ZN(n8663) );
  NAND2_X1 U10120 ( .A1(n8670), .A2(n8663), .ZN(n8647) );
  NAND2_X1 U10121 ( .A1(n8525), .A2(n4521), .ZN(n8563) );
  OR3_X1 U10122 ( .A1(n8568), .A2(n8567), .A3(n8566), .ZN(n8569) );
  OAI211_X1 U10123 ( .C1(n5224), .C2(n8570), .A(n8569), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8673) );
  INV_X1 U10124 ( .A(n8673), .ZN(n8680) );
  NOR2_X1 U10125 ( .A1(n8570), .A2(n4521), .ZN(n8679) );
  INV_X1 U10126 ( .A(n8571), .ZN(n8572) );
  NAND2_X1 U10127 ( .A1(n8673), .A2(n8572), .ZN(n8651) );
  NAND2_X1 U10128 ( .A1(n8673), .A2(n5687), .ZN(n8650) );
  AND2_X1 U10129 ( .A1(n8574), .A2(n8573), .ZN(n8659) );
  NAND2_X1 U10130 ( .A1(n8575), .A2(n8635), .ZN(n8577) );
  NAND2_X1 U10131 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U10132 ( .A1(n8578), .A2(n8636), .ZN(n8579) );
  NAND2_X1 U10133 ( .A1(n8580), .A2(n8579), .ZN(n8639) );
  INV_X1 U10134 ( .A(n8581), .ZN(n8582) );
  NOR2_X1 U10135 ( .A1(n8639), .A2(n8582), .ZN(n8653) );
  INV_X1 U10136 ( .A(n8583), .ZN(n8624) );
  AOI21_X1 U10137 ( .B1(n6537), .B2(n10173), .A(n8584), .ZN(n8588) );
  INV_X1 U10138 ( .A(n8585), .ZN(n8587) );
  AOI21_X1 U10139 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8591) );
  NOR3_X1 U10140 ( .A1(n8591), .A2(n4648), .A3(n8590), .ZN(n8595) );
  INV_X1 U10141 ( .A(n8592), .ZN(n8594) );
  OAI211_X1 U10142 ( .C1(n8595), .C2(n8594), .A(n8597), .B(n8593), .ZN(n8608)
         );
  INV_X1 U10143 ( .A(n8596), .ZN(n8604) );
  INV_X1 U10144 ( .A(n8597), .ZN(n8601) );
  OAI211_X1 U10145 ( .C1(n8601), .C2(n8600), .A(n8599), .B(n8598), .ZN(n8603)
         );
  NOR3_X1 U10146 ( .A1(n8604), .A2(n8603), .A3(n4840), .ZN(n8607) );
  INV_X1 U10147 ( .A(n8605), .ZN(n8606) );
  AOI21_X1 U10148 ( .B1(n8608), .B2(n8607), .A(n8606), .ZN(n8611) );
  AOI21_X1 U10149 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8615) );
  OAI211_X1 U10150 ( .C1(n8615), .C2(n8614), .A(n8613), .B(n8612), .ZN(n8618)
         );
  AOI21_X1 U10151 ( .B1(n8618), .B2(n8617), .A(n8616), .ZN(n8621) );
  OAI21_X1 U10152 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(n8623) );
  AOI21_X1 U10153 ( .B1(n8624), .B2(n8623), .A(n8622), .ZN(n8627) );
  OAI21_X1 U10154 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8629) );
  INV_X1 U10155 ( .A(n8655), .ZN(n8628) );
  AOI21_X1 U10156 ( .B1(n8653), .B2(n8629), .A(n8628), .ZN(n8643) );
  INV_X1 U10157 ( .A(n8630), .ZN(n8632) );
  NOR2_X1 U10158 ( .A1(n8632), .A2(n8631), .ZN(n8658) );
  INV_X1 U10159 ( .A(n8658), .ZN(n8642) );
  AND4_X1 U10160 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(n8638)
         );
  OAI21_X1 U10161 ( .B1(n8639), .B2(n8638), .A(n8637), .ZN(n8641) );
  AOI21_X1 U10162 ( .B1(n8658), .B2(n8641), .A(n8640), .ZN(n8662) );
  OAI21_X1 U10163 ( .B1(n8643), .B2(n8642), .A(n8662), .ZN(n8646) );
  NAND2_X1 U10164 ( .A1(n8645), .A2(n8644), .ZN(n8665) );
  AOI21_X1 U10165 ( .B1(n8659), .B2(n8646), .A(n8665), .ZN(n8648) );
  OAI21_X1 U10166 ( .B1(n8648), .B2(n8647), .A(n8667), .ZN(n8649) );
  MUX2_X1 U10167 ( .A(n8651), .B(n8650), .S(n8649), .Z(n8678) );
  INV_X1 U10168 ( .A(n8652), .ZN(n8676) );
  INV_X1 U10169 ( .A(n8653), .ZN(n8656) );
  INV_X1 U10170 ( .A(n8654), .ZN(n9884) );
  OAI21_X1 U10171 ( .B1(n8656), .B2(n9884), .A(n8655), .ZN(n8657) );
  NAND2_X1 U10172 ( .A1(n8658), .A2(n8657), .ZN(n8661) );
  INV_X1 U10173 ( .A(n8659), .ZN(n8660) );
  AOI21_X1 U10174 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8666) );
  OAI22_X1 U10175 ( .A1(n8666), .A2(n8665), .B1(n8664), .B2(n8663), .ZN(n8668)
         );
  OAI211_X1 U10176 ( .C1(n6608), .C2(n8669), .A(n8668), .B(n8667), .ZN(n8672)
         );
  NAND3_X1 U10177 ( .A1(n8672), .A2(n8671), .A3(n8670), .ZN(n8674) );
  NAND4_X1 U10178 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n8677)
         );
  OAI211_X1 U10179 ( .C1(n8680), .C2(n8679), .A(n8678), .B(n8677), .ZN(n8681)
         );
  OAI211_X1 U10180 ( .C1(n8684), .C2(n8683), .A(n8682), .B(n8681), .ZN(
        P1_U3242) );
  NAND2_X1 U10181 ( .A1(n8686), .A2(n6575), .ZN(n8688) );
  XNOR2_X1 U10182 ( .A(n8688), .B(n4668), .ZN(n8696) );
  INV_X1 U10183 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8689) );
  OAI22_X1 U10184 ( .A1(n8690), .A2(n9913), .B1(n8689), .B2(n9951), .ZN(n8691)
         );
  AOI21_X1 U10185 ( .B1(n8692), .B2(n10157), .A(n8691), .ZN(n8693) );
  OAI21_X1 U10186 ( .B1(n8694), .B2(n10160), .A(n8693), .ZN(n8695) );
  OAI21_X1 U10187 ( .B1(n8698), .B2(n10167), .A(n8697), .ZN(P1_U3356) );
  MUX2_X1 U10188 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n8699), .S(n10189), .Z(
        n8700) );
  AOI21_X1 U10189 ( .B1(n8701), .B2(n9760), .A(n8700), .ZN(n8702) );
  INV_X1 U10190 ( .A(n8702), .ZN(P1_U3520) );
  INV_X1 U10191 ( .A(n8703), .ZN(n9456) );
  OAI222_X1 U10192 ( .A1(n10115), .A2(n8704), .B1(n10114), .B2(n9456), .C1(
        n5304), .C2(P1_U3086), .ZN(P1_U3328) );
  NOR2_X1 U10193 ( .A1(n8705), .A2(n9240), .ZN(n9031) );
  AOI21_X1 U10194 ( .B1(n9246), .B2(P2_REG2_REG_29__SCAN_IN), .A(n9031), .ZN(
        n8706) );
  OAI21_X1 U10195 ( .B1(n8707), .B2(n9204), .A(n8706), .ZN(n8708) );
  AOI21_X1 U10196 ( .B1(n8709), .B2(n10209), .A(n8708), .ZN(n8710) );
  XNOR2_X1 U10197 ( .A(n8712), .B(n8711), .ZN(n8713) );
  XNOR2_X1 U10198 ( .A(n8714), .B(n8713), .ZN(n8724) );
  INV_X1 U10199 ( .A(n8724), .ZN(n8715) );
  NAND2_X1 U10200 ( .A1(n8715), .A2(n8855), .ZN(n8730) );
  INV_X1 U10201 ( .A(n8716), .ZN(n8717) );
  NAND2_X1 U10202 ( .A1(n9039), .A2(n8845), .ZN(n8721) );
  AOI22_X1 U10203 ( .A1(n9045), .A2(n8863), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8720) );
  OAI211_X1 U10204 ( .C1(n8723), .C2(n8848), .A(n8721), .B(n8720), .ZN(n8726)
         );
  NOR4_X1 U10205 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8853), .ZN(n8725)
         );
  AOI211_X1 U10206 ( .C1(n9352), .C2(n8851), .A(n8726), .B(n8725), .ZN(n8727)
         );
  OAI211_X1 U10207 ( .C1(n8730), .C2(n8729), .A(n8728), .B(n8727), .ZN(
        P2_U3160) );
  NAND2_X1 U10208 ( .A1(n9767), .A2(n8731), .ZN(n8733) );
  NAND2_X1 U10209 ( .A1(n9608), .A2(n5905), .ZN(n8732) );
  NAND2_X1 U10210 ( .A1(n8733), .A2(n8732), .ZN(n8735) );
  XNOR2_X1 U10211 ( .A(n8735), .B(n8734), .ZN(n8741) );
  NAND2_X1 U10212 ( .A1(n9767), .A2(n8736), .ZN(n8737) );
  OAI21_X1 U10213 ( .B1(n8739), .B2(n8738), .A(n8737), .ZN(n8740) );
  XNOR2_X1 U10214 ( .A(n8741), .B(n8740), .ZN(n8744) );
  INV_X1 U10215 ( .A(n8744), .ZN(n8749) );
  NAND2_X1 U10216 ( .A1(n8743), .A2(n8742), .ZN(n8748) );
  NAND3_X1 U10217 ( .A1(n8749), .A2(n5931), .A3(n8748), .ZN(n8753) );
  INV_X1 U10218 ( .A(n9765), .ZN(n8745) );
  AOI22_X1 U10219 ( .A1(n8745), .A2(n9538), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8746) );
  OAI21_X1 U10220 ( .B1(n8747), .B2(n9558), .A(n8746), .ZN(n8751) );
  NOR3_X1 U10221 ( .A1(n8749), .A2(n9589), .A3(n8748), .ZN(n8750) );
  AOI211_X1 U10222 ( .C1(n9767), .C2(n4405), .A(n8751), .B(n8750), .ZN(n8752)
         );
  INV_X1 U10223 ( .A(n8756), .ZN(n9444) );
  OAI222_X1 U10224 ( .A1(P1_U3086), .A2(n8755), .B1(n10114), .B2(n9444), .C1(
        n8757), .C2(n10115), .ZN(P1_U3325) );
  AOI22_X1 U10225 ( .A1(n8978), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n8763) );
  OAI21_X1 U10226 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n8759), .A(n8758), .ZN(
        n8760) );
  OAI21_X1 U10227 ( .B1(n8761), .B2(n9023), .A(n8760), .ZN(n8762) );
  OAI211_X1 U10228 ( .C1(n9018), .C2(n8764), .A(n8763), .B(n8762), .ZN(
        P2_U3182) );
  XNOR2_X1 U10229 ( .A(n8813), .B(n8817), .ZN(n8769) );
  AOI22_X1 U10230 ( .A1(n9126), .A2(n8859), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8766) );
  NAND2_X1 U10231 ( .A1(n9098), .A2(n8863), .ZN(n8765) );
  OAI211_X1 U10232 ( .C1(n8790), .C2(n8861), .A(n8766), .B(n8765), .ZN(n8767)
         );
  AOI21_X1 U10233 ( .B1(n9380), .B2(n8851), .A(n8767), .ZN(n8768) );
  OAI21_X1 U10234 ( .B1(n8769), .B2(n8853), .A(n8768), .ZN(P2_U3156) );
  INV_X1 U10235 ( .A(n9302), .ZN(n9156) );
  AOI211_X1 U10236 ( .C1(n8772), .C2(n8771), .A(n8853), .B(n8770), .ZN(n8773)
         );
  INV_X1 U10237 ( .A(n8773), .ZN(n8777) );
  NAND2_X1 U10238 ( .A1(n9187), .A2(n8859), .ZN(n8774) );
  NAND2_X1 U10239 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9019) );
  OAI211_X1 U10240 ( .C1(n9153), .C2(n8861), .A(n8774), .B(n9019), .ZN(n8775)
         );
  AOI21_X1 U10241 ( .B1(n9154), .B2(n8863), .A(n8775), .ZN(n8776) );
  OAI211_X1 U10242 ( .C1(n9156), .C2(n8866), .A(n8777), .B(n8776), .ZN(
        P2_U3159) );
  XOR2_X1 U10243 ( .A(n8779), .B(n8778), .Z(n8785) );
  AOI22_X1 U10244 ( .A1(n9125), .A2(n8859), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8781) );
  NAND2_X1 U10245 ( .A1(n9129), .A2(n8863), .ZN(n8780) );
  OAI211_X1 U10246 ( .C1(n8782), .C2(n8861), .A(n8781), .B(n8780), .ZN(n8783)
         );
  AOI21_X1 U10247 ( .B1(n9392), .B2(n8851), .A(n8783), .ZN(n8784) );
  OAI21_X1 U10248 ( .B1(n8785), .B2(n8853), .A(n8784), .ZN(P2_U3163) );
  XOR2_X1 U10249 ( .A(n8787), .B(n8786), .Z(n8793) );
  NAND2_X1 U10250 ( .A1(n9069), .A2(n8845), .ZN(n8789) );
  AOI22_X1 U10251 ( .A1(n9071), .A2(n8863), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8788) );
  OAI211_X1 U10252 ( .C1(n8790), .C2(n8848), .A(n8789), .B(n8788), .ZN(n8791)
         );
  AOI21_X1 U10253 ( .B1(n9370), .B2(n8851), .A(n8791), .ZN(n8792) );
  OAI21_X1 U10254 ( .B1(n8793), .B2(n8853), .A(n8792), .ZN(P2_U3165) );
  INV_X1 U10255 ( .A(n8794), .ZN(n9414) );
  OAI211_X1 U10256 ( .C1(n8797), .C2(n8796), .A(n8795), .B(n8855), .ZN(n8801)
         );
  NAND2_X1 U10257 ( .A1(n8859), .A2(n9226), .ZN(n8798) );
  NAND2_X1 U10258 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8933) );
  OAI211_X1 U10259 ( .C1(n9199), .C2(n8861), .A(n8798), .B(n8933), .ZN(n8799)
         );
  AOI21_X1 U10260 ( .B1(n8863), .B2(n9202), .A(n8799), .ZN(n8800) );
  OAI211_X1 U10261 ( .C1(n9414), .C2(n8866), .A(n8801), .B(n8800), .ZN(
        P2_U3166) );
  INV_X1 U10262 ( .A(n8802), .ZN(n8803) );
  AOI21_X1 U10263 ( .B1(n8805), .B2(n8804), .A(n8803), .ZN(n8810) );
  NAND2_X1 U10264 ( .A1(n9187), .A2(n8845), .ZN(n8806) );
  NAND2_X1 U10265 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8952) );
  OAI211_X1 U10266 ( .C1(n9214), .C2(n8848), .A(n8806), .B(n8952), .ZN(n8807)
         );
  AOI21_X1 U10267 ( .B1(n8863), .B2(n9191), .A(n8807), .ZN(n8809) );
  NAND2_X1 U10268 ( .A1(n9406), .A2(n8851), .ZN(n8808) );
  OAI211_X1 U10269 ( .C1(n8810), .C2(n8853), .A(n8809), .B(n8808), .ZN(
        P2_U3168) );
  OAI22_X1 U10270 ( .A1(n8813), .A2(n9109), .B1(n8812), .B2(n8811), .ZN(n8816)
         );
  XNOR2_X1 U10271 ( .A(n8814), .B(n9095), .ZN(n8815) );
  XNOR2_X1 U10272 ( .A(n8816), .B(n8815), .ZN(n8822) );
  OAI22_X1 U10273 ( .A1(n8817), .A2(n8848), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10416), .ZN(n8818) );
  AOI21_X1 U10274 ( .B1(n9085), .B2(n8863), .A(n8818), .ZN(n8819) );
  OAI21_X1 U10275 ( .B1(n8849), .B2(n8861), .A(n8819), .ZN(n8820) );
  AOI21_X1 U10276 ( .B1(n9375), .B2(n8851), .A(n8820), .ZN(n8821) );
  OAI21_X1 U10277 ( .B1(n8822), .B2(n8853), .A(n8821), .ZN(P2_U3169) );
  OAI21_X1 U10278 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(n8827) );
  NAND2_X1 U10279 ( .A1(n8827), .A2(n8855), .ZN(n8831) );
  AOI22_X1 U10280 ( .A1(n9108), .A2(n8845), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8828) );
  OAI21_X1 U10281 ( .B1(n9135), .B2(n8848), .A(n8828), .ZN(n8829) );
  AOI21_X1 U10282 ( .B1(n9141), .B2(n8863), .A(n8829), .ZN(n8830) );
  OAI211_X1 U10283 ( .C1(n9399), .C2(n8866), .A(n8831), .B(n8830), .ZN(
        P2_U3173) );
  OAI21_X1 U10284 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8835) );
  NAND2_X1 U10285 ( .A1(n8835), .A2(n8855), .ZN(n8839) );
  AND2_X1 U10286 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8977) );
  AOI21_X1 U10287 ( .B1(n9164), .B2(n8845), .A(n8977), .ZN(n8836) );
  OAI21_X1 U10288 ( .B1(n9199), .B2(n8848), .A(n8836), .ZN(n8837) );
  AOI21_X1 U10289 ( .B1(n9166), .B2(n8863), .A(n8837), .ZN(n8838) );
  OAI211_X1 U10290 ( .C1(n9309), .C2(n8866), .A(n8839), .B(n8838), .ZN(
        P2_U3178) );
  NAND2_X1 U10291 ( .A1(n8841), .A2(n8840), .ZN(n8844) );
  XNOR2_X1 U10292 ( .A(n8842), .B(n9069), .ZN(n8843) );
  XNOR2_X1 U10293 ( .A(n8844), .B(n8843), .ZN(n8854) );
  NAND2_X1 U10294 ( .A1(n9062), .A2(n8845), .ZN(n8847) );
  AOI22_X1 U10295 ( .A1(n9065), .A2(n8863), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8846) );
  OAI211_X1 U10296 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8850)
         );
  AOI21_X1 U10297 ( .B1(n9364), .B2(n8851), .A(n8850), .ZN(n8852) );
  OAI21_X1 U10298 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(P2_U3180) );
  INV_X1 U10299 ( .A(n9417), .ZN(n8867) );
  OAI211_X1 U10300 ( .C1(n8858), .C2(n8857), .A(n8856), .B(n8855), .ZN(n8865)
         );
  NAND2_X1 U10301 ( .A1(n8859), .A2(n9238), .ZN(n8860) );
  NAND2_X1 U10302 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8906) );
  OAI211_X1 U10303 ( .C1(n9214), .C2(n8861), .A(n8860), .B(n8906), .ZN(n8862)
         );
  AOI21_X1 U10304 ( .B1(n8863), .B2(n9218), .A(n8862), .ZN(n8864) );
  OAI211_X1 U10305 ( .C1(n8867), .C2(n8866), .A(n8865), .B(n8864), .ZN(
        P2_U3181) );
  MUX2_X1 U10306 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9030), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10307 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8868), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10308 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9039), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10309 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9051), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10310 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9062), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10311 ( .A(n9069), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8877), .Z(
        P2_U3517) );
  MUX2_X1 U10312 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9083), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10313 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9095), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10314 ( .A(n9109), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8877), .Z(
        P2_U3514) );
  MUX2_X1 U10315 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9126), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10316 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9108), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10317 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9125), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10318 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9164), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9187), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10320 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9163), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10321 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n6269), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10322 ( .A(n9226), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8877), .Z(
        P2_U3506) );
  MUX2_X1 U10323 ( .A(n9238), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8877), .Z(
        P2_U3505) );
  MUX2_X1 U10324 ( .A(n9225), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8877), .Z(
        P2_U3504) );
  MUX2_X1 U10325 ( .A(n9237), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8877), .Z(
        P2_U3503) );
  MUX2_X1 U10326 ( .A(n8869), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8877), .Z(
        P2_U3502) );
  MUX2_X1 U10327 ( .A(n8870), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8877), .Z(
        P2_U3501) );
  MUX2_X1 U10328 ( .A(n8871), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8877), .Z(
        P2_U3500) );
  MUX2_X1 U10329 ( .A(n8872), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8877), .Z(
        P2_U3499) );
  MUX2_X1 U10330 ( .A(n8873), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8877), .Z(
        P2_U3498) );
  MUX2_X1 U10331 ( .A(n8874), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8877), .Z(
        P2_U3497) );
  MUX2_X1 U10332 ( .A(n8875), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8877), .Z(
        P2_U3496) );
  MUX2_X1 U10333 ( .A(n8876), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8877), .Z(
        P2_U3495) );
  MUX2_X1 U10334 ( .A(n10200), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8877), .Z(
        P2_U3494) );
  MUX2_X1 U10335 ( .A(n7397), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8877), .Z(
        P2_U3493) );
  MUX2_X1 U10336 ( .A(n10198), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8877), .Z(
        P2_U3492) );
  MUX2_X1 U10337 ( .A(n8878), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8877), .Z(
        P2_U3491) );
  XOR2_X1 U10338 ( .A(n8879), .B(n8880), .Z(n8881) );
  NAND2_X1 U10339 ( .A1(n8881), .A2(n9023), .ZN(n8894) );
  OAI21_X1 U10340 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n8885) );
  AOI22_X1 U10341 ( .A1(n8886), .A2(n8885), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n8893) );
  OAI21_X1 U10342 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n8890) );
  AOI22_X1 U10343 ( .A1(n8978), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n9006), .B2(
        n8890), .ZN(n8892) );
  NAND2_X1 U10344 ( .A1(n8991), .A2(n4787), .ZN(n8891) );
  NAND4_X1 U10345 ( .A1(n8894), .A2(n8893), .A3(n8892), .A4(n8891), .ZN(
        P2_U3184) );
  OR2_X1 U10346 ( .A1(n8910), .A2(n8895), .ZN(n8896) );
  OAI21_X1 U10347 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8900), .A(n8923), .ZN(
        n8901) );
  INV_X1 U10348 ( .A(n8901), .ZN(n8918) );
  NAND2_X1 U10349 ( .A1(n8903), .A2(n8902), .ZN(n8905) );
  MUX2_X1 U10350 ( .A(P2_REG1_REG_15__SCAN_IN), .B(P2_REG2_REG_15__SCAN_IN), 
        .S(n9009), .Z(n8927) );
  XNOR2_X1 U10351 ( .A(n8927), .B(n8928), .ZN(n8904) );
  NAND2_X1 U10352 ( .A1(n8905), .A2(n8904), .ZN(n8931) );
  OAI21_X1 U10353 ( .B1(n8905), .B2(n8904), .A(n8931), .ZN(n8909) );
  INV_X1 U10354 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U10355 ( .A1(n8991), .A2(n8928), .ZN(n8907) );
  OAI211_X1 U10356 ( .C1(n9020), .C2(n10292), .A(n8907), .B(n8906), .ZN(n8908)
         );
  AOI21_X1 U10357 ( .B1(n8909), .B2(n9023), .A(n8908), .ZN(n8917) );
  OR2_X1 U10358 ( .A1(n8910), .A2(n9321), .ZN(n8911) );
  OAI21_X1 U10359 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8914), .A(n8939), .ZN(
        n8915) );
  NAND2_X1 U10360 ( .A1(n8915), .A2(n9006), .ZN(n8916) );
  OAI211_X1 U10361 ( .C1(n8918), .C2(n9027), .A(n8917), .B(n8916), .ZN(
        P2_U3197) );
  INV_X1 U10362 ( .A(n8919), .ZN(n8921) );
  INV_X1 U10363 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U10364 ( .A(n8937), .B(n8920), .ZN(n8922) );
  AND3_X1 U10365 ( .A1(n8923), .A2(n8922), .A3(n8921), .ZN(n8924) );
  NOR2_X1 U10366 ( .A1(n8944), .A2(n8924), .ZN(n8943) );
  MUX2_X1 U10367 ( .A(P2_REG1_REG_16__SCAN_IN), .B(P2_REG2_REG_16__SCAN_IN), 
        .S(n9009), .Z(n8926) );
  INV_X1 U10368 ( .A(n8926), .ZN(n8925) );
  NAND2_X1 U10369 ( .A1(n8925), .A2(n8937), .ZN(n8950) );
  NAND2_X1 U10370 ( .A1(n8926), .A2(n8958), .ZN(n8948) );
  NAND2_X1 U10371 ( .A1(n8950), .A2(n8948), .ZN(n8932) );
  INV_X1 U10372 ( .A(n8927), .ZN(n8929) );
  NAND2_X1 U10373 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  NAND2_X1 U10374 ( .A1(n8931), .A2(n8930), .ZN(n8949) );
  XOR2_X1 U10375 ( .A(n8932), .B(n8949), .Z(n8936) );
  NAND2_X1 U10376 ( .A1(n8978), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8934) );
  OAI211_X1 U10377 ( .C1(n9018), .C2(n8958), .A(n8934), .B(n8933), .ZN(n8935)
         );
  AOI21_X1 U10378 ( .B1(n8936), .B2(n9023), .A(n8935), .ZN(n8942) );
  INV_X1 U10379 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9315) );
  XNOR2_X1 U10380 ( .A(n8937), .B(n9315), .ZN(n8938) );
  AND3_X1 U10381 ( .A1(n8939), .A2(n8938), .A3(n4430), .ZN(n8940) );
  OAI21_X1 U10382 ( .B1(n8957), .B2(n8940), .A(n9006), .ZN(n8941) );
  OAI211_X1 U10383 ( .C1(n8943), .C2(n9027), .A(n8942), .B(n8941), .ZN(
        P2_U3198) );
  OAI21_X1 U10384 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8946), .A(n8967), .ZN(
        n8947) );
  INV_X1 U10385 ( .A(n8947), .ZN(n8964) );
  NAND2_X1 U10386 ( .A1(n8949), .A2(n8948), .ZN(n8951) );
  NAND2_X1 U10387 ( .A1(n8951), .A2(n8950), .ZN(n8984) );
  MUX2_X1 U10388 ( .A(P2_REG1_REG_17__SCAN_IN), .B(P2_REG2_REG_17__SCAN_IN), 
        .S(n9009), .Z(n8979) );
  XNOR2_X1 U10389 ( .A(n8979), .B(n8980), .ZN(n8983) );
  XNOR2_X1 U10390 ( .A(n8984), .B(n8983), .ZN(n8956) );
  NAND2_X1 U10391 ( .A1(n8978), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U10392 ( .C1(n9018), .C2(n8954), .A(n8953), .B(n8952), .ZN(n8955)
         );
  AOI21_X1 U10393 ( .B1(n8956), .B2(n9023), .A(n8955), .ZN(n8963) );
  AOI21_X1 U10394 ( .B1(n8959), .B2(n8980), .A(n8971), .ZN(n8960) );
  NAND2_X1 U10395 ( .A1(n8960), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8975) );
  OAI21_X1 U10396 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8960), .A(n8975), .ZN(
        n8961) );
  NAND2_X1 U10397 ( .A1(n8961), .A2(n9006), .ZN(n8962) );
  OAI211_X1 U10398 ( .C1(n8964), .C2(n9027), .A(n8963), .B(n8962), .ZN(
        P2_U3199) );
  INV_X1 U10399 ( .A(n8965), .ZN(n8969) );
  INV_X1 U10400 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9168) );
  OR2_X1 U10401 ( .A1(n8993), .A2(n9168), .ZN(n8997) );
  NAND2_X1 U10402 ( .A1(n8993), .A2(n9168), .ZN(n8966) );
  NAND2_X1 U10403 ( .A1(n8997), .A2(n8966), .ZN(n8968) );
  AND3_X1 U10404 ( .A1(n8967), .A2(n8969), .A3(n8968), .ZN(n8970) );
  INV_X1 U10405 ( .A(n8971), .ZN(n8974) );
  INV_X1 U10406 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10582) );
  OR2_X1 U10407 ( .A1(n8993), .A2(n10582), .ZN(n9002) );
  NAND2_X1 U10408 ( .A1(n8993), .A2(n10582), .ZN(n8972) );
  NAND2_X1 U10409 ( .A1(n9002), .A2(n8972), .ZN(n8973) );
  INV_X1 U10410 ( .A(n8979), .ZN(n8981) );
  AND2_X1 U10411 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  MUX2_X1 U10412 ( .A(P2_REG1_REG_18__SCAN_IN), .B(P2_REG2_REG_18__SCAN_IN), 
        .S(n9009), .Z(n8986) );
  AND2_X1 U10413 ( .A1(n8985), .A2(n8986), .ZN(n9012) );
  INV_X1 U10414 ( .A(n8985), .ZN(n8988) );
  INV_X1 U10415 ( .A(n8986), .ZN(n8987) );
  NAND2_X1 U10416 ( .A1(n8988), .A2(n8987), .ZN(n9013) );
  INV_X1 U10417 ( .A(n9013), .ZN(n8989) );
  NAND2_X1 U10418 ( .A1(n8990), .A2(n9023), .ZN(n8995) );
  INV_X1 U10419 ( .A(n8990), .ZN(n8992) );
  AOI21_X1 U10420 ( .B1(n8992), .B2(P2_U3893), .A(n8991), .ZN(n8994) );
  MUX2_X1 U10421 ( .A(n8995), .B(n8994), .S(n8993), .Z(n8996) );
  INV_X1 U10422 ( .A(n8997), .ZN(n8998) );
  XNOR2_X1 U10423 ( .A(n9000), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U10424 ( .A(n9001), .B(n9008), .ZN(n9028) );
  INV_X1 U10425 ( .A(n9002), .ZN(n9003) );
  NOR2_X1 U10426 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  XNOR2_X1 U10427 ( .A(n9017), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U10428 ( .A(n9005), .B(n9011), .ZN(n9007) );
  NAND2_X1 U10429 ( .A1(n9007), .A2(n9006), .ZN(n9026) );
  INV_X1 U10430 ( .A(n9008), .ZN(n9010) );
  MUX2_X1 U10431 ( .A(n9011), .B(n9010), .S(n9009), .Z(n9016) );
  AOI21_X1 U10432 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9015) );
  XOR2_X1 U10433 ( .A(n9016), .B(n9015), .Z(n9024) );
  NOR2_X1 U10434 ( .A1(n9018), .A2(n9017), .ZN(n9022) );
  OAI21_X1 U10435 ( .B1(n9020), .B2(n10625), .A(n9019), .ZN(n9021) );
  AOI211_X1 U10436 ( .C1(n9024), .C2(n9023), .A(n9022), .B(n9021), .ZN(n9025)
         );
  OAI211_X1 U10437 ( .C1(n9028), .C2(n9027), .A(n9026), .B(n9025), .ZN(
        P2_U3201) );
  AOI21_X1 U10438 ( .B1(n9344), .B2(n10212), .A(n9031), .ZN(n9034) );
  NAND2_X1 U10439 ( .A1(n9246), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9032) );
  OAI211_X1 U10440 ( .C1(n9346), .C2(n9204), .A(n9034), .B(n9032), .ZN(
        P2_U3202) );
  NAND2_X1 U10441 ( .A1(n9246), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9033) );
  OAI211_X1 U10442 ( .C1(n9035), .C2(n9204), .A(n9034), .B(n9033), .ZN(
        P2_U3203) );
  XNOR2_X1 U10443 ( .A(n9036), .B(n9037), .ZN(n9355) );
  MUX2_X1 U10444 ( .A(n9044), .B(n9350), .S(n10212), .Z(n9047) );
  AOI22_X1 U10445 ( .A1(n9352), .A2(n9265), .B1(n10205), .B2(n9045), .ZN(n9046) );
  OAI211_X1 U10446 ( .C1(n9355), .C2(n9268), .A(n9047), .B(n9046), .ZN(
        P2_U3205) );
  XNOR2_X1 U10447 ( .A(n9048), .B(n4418), .ZN(n9361) );
  XNOR2_X1 U10448 ( .A(n9049), .B(n4418), .ZN(n9054) );
  MUX2_X1 U10449 ( .A(n9069), .B(n9051), .S(n9050), .Z(n9052) );
  AOI22_X1 U10450 ( .A1(n9054), .A2(n10202), .B1(n9053), .B2(n9052), .ZN(n9356) );
  MUX2_X1 U10451 ( .A(n9055), .B(n9356), .S(n10212), .Z(n9058) );
  AOI22_X1 U10452 ( .A1(n9358), .A2(n9265), .B1(n10205), .B2(n9056), .ZN(n9057) );
  OAI211_X1 U10453 ( .C1(n9361), .C2(n9268), .A(n9058), .B(n9057), .ZN(
        P2_U3206) );
  XNOR2_X1 U10454 ( .A(n9059), .B(n9060), .ZN(n9367) );
  XNOR2_X1 U10455 ( .A(n9061), .B(n9060), .ZN(n9063) );
  AOI222_X1 U10456 ( .A1(n10202), .A2(n9063), .B1(n9062), .B2(n10199), .C1(
        n9083), .C2(n9236), .ZN(n9362) );
  MUX2_X1 U10457 ( .A(n9064), .B(n9362), .S(n10212), .Z(n9067) );
  AOI22_X1 U10458 ( .A1(n9364), .A2(n9265), .B1(n10205), .B2(n9065), .ZN(n9066) );
  OAI211_X1 U10459 ( .C1(n9367), .C2(n9268), .A(n9067), .B(n9066), .ZN(
        P2_U3207) );
  OAI21_X1 U10460 ( .B1(n4454), .B2(n4758), .A(n9068), .ZN(n9070) );
  AOI22_X1 U10461 ( .A1(n9370), .A2(n10203), .B1(n10205), .B2(n9071), .ZN(
        n9072) );
  AOI21_X1 U10462 ( .B1(n9368), .B2(n9072), .A(n9246), .ZN(n9077) );
  XNOR2_X1 U10463 ( .A(n9073), .B(n9074), .ZN(n9373) );
  OAI22_X1 U10464 ( .A1(n9373), .A2(n9268), .B1(n9075), .B2(n10212), .ZN(n9076) );
  OR2_X1 U10465 ( .A1(n9077), .A2(n9076), .ZN(P2_U3208) );
  NAND2_X1 U10466 ( .A1(n9078), .A2(n9079), .ZN(n9080) );
  XOR2_X1 U10467 ( .A(n9082), .B(n9080), .Z(n9378) );
  XOR2_X1 U10468 ( .A(n9082), .B(n9081), .Z(n9084) );
  AOI222_X1 U10469 ( .A1(n10202), .A2(n9084), .B1(n9083), .B2(n10199), .C1(
        n9109), .C2(n9236), .ZN(n9374) );
  INV_X1 U10470 ( .A(n9374), .ZN(n9089) );
  INV_X1 U10471 ( .A(n9085), .ZN(n9086) );
  OAI22_X1 U10472 ( .A1(n9087), .A2(n9242), .B1(n9086), .B2(n9240), .ZN(n9088)
         );
  OAI21_X1 U10473 ( .B1(n9089), .B2(n9088), .A(n10212), .ZN(n9091) );
  NAND2_X1 U10474 ( .A1(n9246), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9090) );
  OAI211_X1 U10475 ( .C1(n9378), .C2(n9268), .A(n9091), .B(n9090), .ZN(
        P2_U3209) );
  XNOR2_X1 U10476 ( .A(n9092), .B(n9093), .ZN(n9383) );
  INV_X1 U10477 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U10478 ( .A(n9094), .B(n9093), .ZN(n9096) );
  AOI222_X1 U10479 ( .A1(n10202), .A2(n9096), .B1(n9095), .B2(n10199), .C1(
        n9126), .C2(n9236), .ZN(n9379) );
  MUX2_X1 U10480 ( .A(n9097), .B(n9379), .S(n10212), .Z(n9100) );
  AOI22_X1 U10481 ( .A1(n9380), .A2(n9265), .B1(n10205), .B2(n9098), .ZN(n9099) );
  OAI211_X1 U10482 ( .C1(n9383), .C2(n9268), .A(n9100), .B(n9099), .ZN(
        P2_U3210) );
  XNOR2_X1 U10483 ( .A(n9101), .B(n9103), .ZN(n9389) );
  INV_X1 U10484 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9111) );
  AND2_X1 U10485 ( .A1(n9132), .A2(n9139), .ZN(n9134) );
  OAI21_X1 U10486 ( .B1(n9134), .B2(n9122), .A(n9121), .ZN(n9124) );
  NAND3_X1 U10487 ( .A1(n9124), .A2(n9103), .A3(n9102), .ZN(n9107) );
  OAI21_X1 U10488 ( .B1(n4419), .B2(n9105), .A(n9104), .ZN(n9106) );
  NAND2_X1 U10489 ( .A1(n9107), .A2(n9106), .ZN(n9110) );
  AOI222_X1 U10490 ( .A1(n10202), .A2(n9110), .B1(n9109), .B2(n10199), .C1(
        n9108), .C2(n9236), .ZN(n9384) );
  MUX2_X1 U10491 ( .A(n9111), .B(n9384), .S(n10212), .Z(n9114) );
  AOI22_X1 U10492 ( .A1(n9386), .A2(n9265), .B1(n10205), .B2(n9112), .ZN(n9113) );
  OAI211_X1 U10493 ( .C1(n9389), .C2(n9268), .A(n9114), .B(n9113), .ZN(
        P2_U3211) );
  NAND2_X1 U10494 ( .A1(n9116), .A2(n9115), .ZN(n9140) );
  INV_X1 U10495 ( .A(n9117), .ZN(n9119) );
  OAI21_X1 U10496 ( .B1(n9140), .B2(n9119), .A(n9118), .ZN(n9120) );
  XNOR2_X1 U10497 ( .A(n9120), .B(n9121), .ZN(n9395) );
  OR3_X1 U10498 ( .A1(n9134), .A2(n9122), .A3(n9121), .ZN(n9123) );
  NAND2_X1 U10499 ( .A1(n9124), .A2(n9123), .ZN(n9127) );
  AOI222_X1 U10500 ( .A1(n10202), .A2(n9127), .B1(n9126), .B2(n10199), .C1(
        n9125), .C2(n9236), .ZN(n9390) );
  MUX2_X1 U10501 ( .A(n9128), .B(n9390), .S(n10212), .Z(n9131) );
  AOI22_X1 U10502 ( .A1(n9392), .A2(n9265), .B1(n10205), .B2(n9129), .ZN(n9130) );
  OAI211_X1 U10503 ( .C1(n9395), .C2(n9268), .A(n9131), .B(n9130), .ZN(
        P2_U3212) );
  NOR2_X1 U10504 ( .A1(n9132), .A2(n9139), .ZN(n9133) );
  OR2_X1 U10505 ( .A1(n9134), .A2(n9133), .ZN(n9138) );
  OAI22_X1 U10506 ( .A1(n9136), .A2(n9261), .B1(n9135), .B2(n9259), .ZN(n9137)
         );
  AOI21_X1 U10507 ( .B1(n9138), .B2(n10202), .A(n9137), .ZN(n9299) );
  XNOR2_X1 U10508 ( .A(n9140), .B(n9139), .ZN(n9297) );
  AOI22_X1 U10509 ( .A1(n9141), .A2(n10205), .B1(n9246), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n9142) );
  OAI21_X1 U10510 ( .B1(n9399), .B2(n9204), .A(n9142), .ZN(n9143) );
  AOI21_X1 U10511 ( .B1(n9297), .B2(n9206), .A(n9143), .ZN(n9144) );
  OAI21_X1 U10512 ( .B1(n9299), .B2(n9246), .A(n9144), .ZN(P2_U3213) );
  INV_X1 U10513 ( .A(n9145), .ZN(n9146) );
  NOR2_X1 U10514 ( .A1(n9173), .A2(n9172), .ZN(n9171) );
  NOR2_X1 U10515 ( .A1(n9171), .A2(n9147), .ZN(n9148) );
  XNOR2_X1 U10516 ( .A(n9148), .B(n9149), .ZN(n9402) );
  XNOR2_X1 U10517 ( .A(n9150), .B(n9149), .ZN(n9151) );
  OAI222_X1 U10518 ( .A1(n9261), .A2(n9153), .B1(n9259), .B2(n9152), .C1(n9151), .C2(n9256), .ZN(n9301) );
  AOI22_X1 U10519 ( .A1(n9246), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9154), .B2(
        n10205), .ZN(n9155) );
  OAI21_X1 U10520 ( .B1(n9156), .B2(n9204), .A(n9155), .ZN(n9157) );
  AOI21_X1 U10521 ( .B1(n9301), .B2(n10212), .A(n9157), .ZN(n9158) );
  OAI21_X1 U10522 ( .B1(n9402), .B2(n9268), .A(n9158), .ZN(P2_U3214) );
  OR2_X1 U10523 ( .A1(n9212), .A2(n9159), .ZN(n9161) );
  AND2_X1 U10524 ( .A1(n9161), .A2(n9160), .ZN(n9162) );
  XOR2_X1 U10525 ( .A(n9172), .B(n9162), .Z(n9165) );
  AOI222_X1 U10526 ( .A1(n10202), .A2(n9165), .B1(n9164), .B2(n10199), .C1(
        n9163), .C2(n9236), .ZN(n9308) );
  INV_X1 U10527 ( .A(n9166), .ZN(n9167) );
  OAI22_X1 U10528 ( .A1(n10212), .A2(n9168), .B1(n9167), .B2(n9240), .ZN(n9169) );
  AOI21_X1 U10529 ( .B1(n9170), .B2(n9265), .A(n9169), .ZN(n9175) );
  INV_X1 U10530 ( .A(n9171), .ZN(n9306) );
  NAND2_X1 U10531 ( .A1(n9173), .A2(n9172), .ZN(n9305) );
  NAND3_X1 U10532 ( .A1(n9306), .A2(n9206), .A3(n9305), .ZN(n9174) );
  OAI211_X1 U10533 ( .C1(n9308), .C2(n9246), .A(n9175), .B(n9174), .ZN(
        P2_U3215) );
  OR2_X1 U10534 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  OR2_X1 U10535 ( .A1(n9212), .A2(n9180), .ZN(n9182) );
  NAND2_X1 U10536 ( .A1(n9182), .A2(n9181), .ZN(n9195) );
  INV_X1 U10537 ( .A(n9201), .ZN(n9196) );
  NOR2_X1 U10538 ( .A1(n9195), .A2(n9196), .ZN(n9194) );
  OAI21_X1 U10539 ( .B1(n9194), .B2(n9184), .A(n9183), .ZN(n9186) );
  OR3_X1 U10540 ( .A1(n9194), .A2(n9184), .A3(n9183), .ZN(n9185) );
  NAND3_X1 U10541 ( .A1(n9186), .A2(n10202), .A3(n9185), .ZN(n9189) );
  AOI22_X1 U10542 ( .A1(n9187), .A2(n10199), .B1(n6269), .B2(n9236), .ZN(n9188) );
  INV_X1 U10543 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U10544 ( .A(n9405), .B(n9190), .S(n9246), .Z(n9193) );
  AOI22_X1 U10545 ( .A1(n9406), .A2(n9265), .B1(n10205), .B2(n9191), .ZN(n9192) );
  OAI211_X1 U10546 ( .C1(n9409), .C2(n9268), .A(n9193), .B(n9192), .ZN(
        P2_U3216) );
  AOI211_X1 U10547 ( .C1(n9196), .C2(n9195), .A(n9256), .B(n9194), .ZN(n9197)
         );
  AOI21_X1 U10548 ( .B1(n9236), .B2(n9226), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10549 ( .B1(n9199), .B2(n9261), .A(n9198), .ZN(n9313) );
  INV_X1 U10550 ( .A(n9313), .ZN(n9208) );
  XNOR2_X1 U10551 ( .A(n9200), .B(n9201), .ZN(n9314) );
  AOI22_X1 U10552 ( .A1(n9246), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10205), 
        .B2(n9202), .ZN(n9203) );
  OAI21_X1 U10553 ( .B1(n9414), .B2(n9204), .A(n9203), .ZN(n9205) );
  AOI21_X1 U10554 ( .B1(n9314), .B2(n9206), .A(n9205), .ZN(n9207) );
  OAI21_X1 U10555 ( .B1(n9208), .B2(n9246), .A(n9207), .ZN(P2_U3217) );
  XNOR2_X1 U10556 ( .A(n9209), .B(n9210), .ZN(n9420) );
  INV_X1 U10557 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9217) );
  XNOR2_X1 U10558 ( .A(n9212), .B(n9211), .ZN(n9216) );
  OAI22_X1 U10559 ( .A1(n9214), .A2(n9261), .B1(n9213), .B2(n9259), .ZN(n9215)
         );
  AOI21_X1 U10560 ( .B1(n9216), .B2(n10202), .A(n9215), .ZN(n9415) );
  MUX2_X1 U10561 ( .A(n9217), .B(n9415), .S(n10212), .Z(n9220) );
  AOI22_X1 U10562 ( .A1(n9417), .A2(n9265), .B1(n10205), .B2(n9218), .ZN(n9219) );
  OAI211_X1 U10563 ( .C1(n9420), .C2(n9268), .A(n9220), .B(n9219), .ZN(
        P2_U3218) );
  XNOR2_X1 U10564 ( .A(n9222), .B(n9221), .ZN(n9426) );
  XNOR2_X1 U10565 ( .A(n9224), .B(n9223), .ZN(n9227) );
  AOI222_X1 U10566 ( .A1(n10202), .A2(n9227), .B1(n9226), .B2(n10199), .C1(
        n9225), .C2(n9236), .ZN(n9421) );
  OAI21_X1 U10567 ( .B1(n9228), .B2(n9242), .A(n9421), .ZN(n9229) );
  NAND2_X1 U10568 ( .A1(n9229), .A2(n10212), .ZN(n9232) );
  AOI22_X1 U10569 ( .A1(n9246), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10205), 
        .B2(n9230), .ZN(n9231) );
  OAI211_X1 U10570 ( .C1(n9426), .C2(n9268), .A(n9232), .B(n9231), .ZN(
        P2_U3219) );
  XNOR2_X1 U10571 ( .A(n9233), .B(n9234), .ZN(n9431) );
  XNOR2_X1 U10572 ( .A(n9235), .B(n9234), .ZN(n9239) );
  AOI222_X1 U10573 ( .A1(n10202), .A2(n9239), .B1(n9238), .B2(n10199), .C1(
        n9237), .C2(n9236), .ZN(n9427) );
  INV_X1 U10574 ( .A(n9427), .ZN(n9245) );
  OAI22_X1 U10575 ( .A1(n9243), .A2(n9242), .B1(n9241), .B2(n9240), .ZN(n9244)
         );
  OAI21_X1 U10576 ( .B1(n9245), .B2(n9244), .A(n10212), .ZN(n9248) );
  NAND2_X1 U10577 ( .A1(n9246), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9247) );
  OAI211_X1 U10578 ( .C1(n9431), .C2(n9268), .A(n9248), .B(n9247), .ZN(
        P2_U3220) );
  INV_X1 U10579 ( .A(n9255), .ZN(n9250) );
  OAI21_X1 U10580 ( .B1(n4507), .B2(n9250), .A(n9249), .ZN(n9436) );
  AND2_X1 U10581 ( .A1(n4486), .A2(n9253), .ZN(n9254) );
  XOR2_X1 U10582 ( .A(n9255), .B(n9254), .Z(n9257) );
  OAI222_X1 U10583 ( .A1(n9261), .A2(n9260), .B1(n9259), .B2(n9258), .C1(n9257), .C2(n9256), .ZN(n9327) );
  INV_X1 U10584 ( .A(n9327), .ZN(n9262) );
  MUX2_X1 U10585 ( .A(n9263), .B(n9262), .S(n10212), .Z(n9267) );
  AOI22_X1 U10586 ( .A1(n9328), .A2(n9265), .B1(n10205), .B2(n9264), .ZN(n9266) );
  OAI211_X1 U10587 ( .C1(n9436), .C2(n9268), .A(n9267), .B(n9266), .ZN(
        P2_U3221) );
  NAND2_X1 U10588 ( .A1(n9344), .A2(n10257), .ZN(n9270) );
  NAND2_X1 U10589 ( .A1(n9273), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9269) );
  OAI211_X1 U10590 ( .C1(n9346), .C2(n9317), .A(n9270), .B(n9269), .ZN(
        P2_U3490) );
  NAND2_X1 U10591 ( .A1(n9347), .A2(n6963), .ZN(n9271) );
  OAI211_X1 U10592 ( .C1(n10257), .C2(n10458), .A(n9271), .B(n9270), .ZN(
        P2_U3489) );
  INV_X1 U10593 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U10594 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U10595 ( .A1(n9352), .A2(n6963), .ZN(n9276) );
  OAI211_X1 U10596 ( .C1(n9355), .C2(n9332), .A(n9277), .B(n9276), .ZN(
        P2_U3487) );
  INV_X1 U10597 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9278) );
  MUX2_X1 U10598 ( .A(n9278), .B(n9356), .S(n10257), .Z(n9280) );
  NAND2_X1 U10599 ( .A1(n9358), .A2(n6963), .ZN(n9279) );
  OAI211_X1 U10600 ( .C1(n9361), .C2(n9332), .A(n9280), .B(n9279), .ZN(
        P2_U3486) );
  INV_X1 U10601 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9281) );
  MUX2_X1 U10602 ( .A(n9281), .B(n9362), .S(n10257), .Z(n9283) );
  NAND2_X1 U10603 ( .A1(n9364), .A2(n6963), .ZN(n9282) );
  OAI211_X1 U10604 ( .C1(n9332), .C2(n9367), .A(n9283), .B(n9282), .ZN(
        P2_U3485) );
  INV_X1 U10605 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10320) );
  MUX2_X1 U10606 ( .A(n10320), .B(n9368), .S(n10257), .Z(n9285) );
  NAND2_X1 U10607 ( .A1(n9370), .A2(n6963), .ZN(n9284) );
  INV_X1 U10608 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9286) );
  MUX2_X1 U10609 ( .A(n9286), .B(n9374), .S(n10257), .Z(n9288) );
  NAND2_X1 U10610 ( .A1(n9375), .A2(n6963), .ZN(n9287) );
  OAI211_X1 U10611 ( .C1(n9332), .C2(n9378), .A(n9288), .B(n9287), .ZN(
        P2_U3483) );
  INV_X1 U10612 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9289) );
  MUX2_X1 U10613 ( .A(n9289), .B(n9379), .S(n10257), .Z(n9291) );
  NAND2_X1 U10614 ( .A1(n9380), .A2(n6963), .ZN(n9290) );
  OAI211_X1 U10615 ( .C1(n9383), .C2(n9332), .A(n9291), .B(n9290), .ZN(
        P2_U3482) );
  MUX2_X1 U10616 ( .A(n10565), .B(n9384), .S(n10257), .Z(n9293) );
  NAND2_X1 U10617 ( .A1(n9386), .A2(n6963), .ZN(n9292) );
  OAI211_X1 U10618 ( .C1(n9389), .C2(n9332), .A(n9293), .B(n9292), .ZN(
        P2_U3481) );
  INV_X1 U10619 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9294) );
  MUX2_X1 U10620 ( .A(n9294), .B(n9390), .S(n10257), .Z(n9296) );
  NAND2_X1 U10621 ( .A1(n9392), .A2(n6963), .ZN(n9295) );
  OAI211_X1 U10622 ( .C1(n9332), .C2(n9395), .A(n9296), .B(n9295), .ZN(
        P2_U3480) );
  NAND2_X1 U10623 ( .A1(n9297), .A2(n10238), .ZN(n9298) );
  AND2_X1 U10624 ( .A1(n9299), .A2(n9298), .ZN(n9396) );
  MUX2_X1 U10625 ( .A(n10489), .B(n9396), .S(n10257), .Z(n9300) );
  OAI21_X1 U10626 ( .B1(n9399), .B2(n9317), .A(n9300), .ZN(P2_U3479) );
  INV_X1 U10627 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9303) );
  AOI21_X1 U10628 ( .B1(n9329), .B2(n9302), .A(n9301), .ZN(n9400) );
  MUX2_X1 U10629 ( .A(n9303), .B(n9400), .S(n10257), .Z(n9304) );
  OAI21_X1 U10630 ( .B1(n9402), .B2(n9332), .A(n9304), .ZN(P2_U3478) );
  NAND3_X1 U10631 ( .A1(n9306), .A2(n10238), .A3(n9305), .ZN(n9307) );
  OAI211_X1 U10632 ( .C1(n9309), .C2(n10239), .A(n9308), .B(n9307), .ZN(n9403)
         );
  MUX2_X1 U10633 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9403), .S(n10257), .Z(
        P2_U3477) );
  INV_X1 U10634 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9310) );
  MUX2_X1 U10635 ( .A(n9310), .B(n9405), .S(n10257), .Z(n9312) );
  NAND2_X1 U10636 ( .A1(n9406), .A2(n6963), .ZN(n9311) );
  OAI211_X1 U10637 ( .C1(n9409), .C2(n9332), .A(n9312), .B(n9311), .ZN(
        P2_U3476) );
  AOI21_X1 U10638 ( .B1(n10238), .B2(n9314), .A(n9313), .ZN(n9410) );
  MUX2_X1 U10639 ( .A(n9315), .B(n9410), .S(n10257), .Z(n9316) );
  OAI21_X1 U10640 ( .B1(n9414), .B2(n9317), .A(n9316), .ZN(P2_U3475) );
  INV_X1 U10641 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9318) );
  MUX2_X1 U10642 ( .A(n9318), .B(n9415), .S(n10257), .Z(n9320) );
  NAND2_X1 U10643 ( .A1(n9417), .A2(n6963), .ZN(n9319) );
  OAI211_X1 U10644 ( .C1(n9420), .C2(n9332), .A(n9320), .B(n9319), .ZN(
        P2_U3474) );
  MUX2_X1 U10645 ( .A(n9321), .B(n9421), .S(n10257), .Z(n9323) );
  NAND2_X1 U10646 ( .A1(n9423), .A2(n6963), .ZN(n9322) );
  OAI211_X1 U10647 ( .C1(n9426), .C2(n9332), .A(n9323), .B(n9322), .ZN(
        P2_U3473) );
  MUX2_X1 U10648 ( .A(n9324), .B(n9427), .S(n10257), .Z(n9326) );
  NAND2_X1 U10649 ( .A1(n9428), .A2(n6963), .ZN(n9325) );
  OAI211_X1 U10650 ( .C1(n9332), .C2(n9431), .A(n9326), .B(n9325), .ZN(
        P2_U3472) );
  AOI21_X1 U10651 ( .B1(n9329), .B2(n9328), .A(n9327), .ZN(n9432) );
  MUX2_X1 U10652 ( .A(n9330), .B(n9432), .S(n10257), .Z(n9331) );
  OAI21_X1 U10653 ( .B1(n9332), .B2(n9436), .A(n9331), .ZN(P2_U3471) );
  OAI22_X1 U10654 ( .A1(n9335), .A2(n9334), .B1(n9333), .B2(n10239), .ZN(n9336) );
  OR2_X1 U10655 ( .A1(n9337), .A2(n9336), .ZN(n9437) );
  MUX2_X1 U10656 ( .A(n9437), .B(P2_REG1_REG_9__SCAN_IN), .S(n9273), .Z(
        P2_U3468) );
  NOR2_X1 U10657 ( .A1(n9338), .A2(n10239), .ZN(n9339) );
  AOI21_X1 U10658 ( .B1(n9340), .B2(n10238), .A(n9339), .ZN(n9342) );
  AND2_X1 U10659 ( .A1(n9342), .A2(n9341), .ZN(n10214) );
  INV_X1 U10660 ( .A(n10214), .ZN(n9343) );
  MUX2_X1 U10661 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9343), .S(n10257), .Z(
        P2_U3460) );
  NAND2_X1 U10662 ( .A1(n9344), .A2(n10245), .ZN(n9348) );
  NAND2_X1 U10663 ( .A1(n10247), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9345) );
  OAI211_X1 U10664 ( .C1(n9346), .C2(n9413), .A(n9348), .B(n9345), .ZN(
        P2_U3458) );
  NAND2_X1 U10665 ( .A1(n9347), .A2(n6946), .ZN(n9349) );
  OAI211_X1 U10666 ( .C1(n10245), .C2(n10392), .A(n9349), .B(n9348), .ZN(
        P2_U3457) );
  INV_X1 U10667 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9351) );
  MUX2_X1 U10668 ( .A(n9351), .B(n9350), .S(n10245), .Z(n9354) );
  NAND2_X1 U10669 ( .A1(n9352), .A2(n6946), .ZN(n9353) );
  OAI211_X1 U10670 ( .C1(n9355), .C2(n9435), .A(n9354), .B(n9353), .ZN(
        P2_U3455) );
  INV_X1 U10671 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9357) );
  MUX2_X1 U10672 ( .A(n9357), .B(n9356), .S(n10245), .Z(n9360) );
  NAND2_X1 U10673 ( .A1(n9358), .A2(n6946), .ZN(n9359) );
  OAI211_X1 U10674 ( .C1(n9361), .C2(n9435), .A(n9360), .B(n9359), .ZN(
        P2_U3454) );
  INV_X1 U10675 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9363) );
  MUX2_X1 U10676 ( .A(n9363), .B(n9362), .S(n10245), .Z(n9366) );
  NAND2_X1 U10677 ( .A1(n9364), .A2(n6946), .ZN(n9365) );
  OAI211_X1 U10678 ( .C1(n9367), .C2(n9435), .A(n9366), .B(n9365), .ZN(
        P2_U3453) );
  INV_X1 U10679 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9369) );
  MUX2_X1 U10680 ( .A(n9369), .B(n9368), .S(n10245), .Z(n9372) );
  NAND2_X1 U10681 ( .A1(n9370), .A2(n6946), .ZN(n9371) );
  OAI211_X1 U10682 ( .C1(n9373), .C2(n9435), .A(n9372), .B(n9371), .ZN(
        P2_U3452) );
  MUX2_X1 U10683 ( .A(n10508), .B(n9374), .S(n10245), .Z(n9377) );
  NAND2_X1 U10684 ( .A1(n9375), .A2(n6946), .ZN(n9376) );
  OAI211_X1 U10685 ( .C1(n9378), .C2(n9435), .A(n9377), .B(n9376), .ZN(
        P2_U3451) );
  MUX2_X1 U10686 ( .A(n10548), .B(n9379), .S(n10245), .Z(n9382) );
  NAND2_X1 U10687 ( .A1(n9380), .A2(n6946), .ZN(n9381) );
  OAI211_X1 U10688 ( .C1(n9383), .C2(n9435), .A(n9382), .B(n9381), .ZN(
        P2_U3450) );
  INV_X1 U10689 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9385) );
  MUX2_X1 U10690 ( .A(n9385), .B(n9384), .S(n10245), .Z(n9388) );
  NAND2_X1 U10691 ( .A1(n9386), .A2(n6946), .ZN(n9387) );
  OAI211_X1 U10692 ( .C1(n9389), .C2(n9435), .A(n9388), .B(n9387), .ZN(
        P2_U3449) );
  INV_X1 U10693 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9391) );
  MUX2_X1 U10694 ( .A(n9391), .B(n9390), .S(n10245), .Z(n9394) );
  NAND2_X1 U10695 ( .A1(n9392), .A2(n6946), .ZN(n9393) );
  OAI211_X1 U10696 ( .C1(n9395), .C2(n9435), .A(n9394), .B(n9393), .ZN(
        P2_U3448) );
  INV_X1 U10697 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9397) );
  MUX2_X1 U10698 ( .A(n9397), .B(n9396), .S(n10245), .Z(n9398) );
  OAI21_X1 U10699 ( .B1(n9399), .B2(n9413), .A(n9398), .ZN(P2_U3447) );
  MUX2_X1 U10700 ( .A(n10486), .B(n9400), .S(n10245), .Z(n9401) );
  OAI21_X1 U10701 ( .B1(n9402), .B2(n9435), .A(n9401), .ZN(P2_U3446) );
  MUX2_X1 U10702 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9403), .S(n10245), .Z(
        P2_U3444) );
  INV_X1 U10703 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9404) );
  MUX2_X1 U10704 ( .A(n9405), .B(n9404), .S(n10247), .Z(n9408) );
  NAND2_X1 U10705 ( .A1(n9406), .A2(n6946), .ZN(n9407) );
  OAI211_X1 U10706 ( .C1(n9409), .C2(n9435), .A(n9408), .B(n9407), .ZN(
        P2_U3441) );
  INV_X1 U10707 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U10708 ( .A(n9411), .B(n9410), .S(n10245), .Z(n9412) );
  OAI21_X1 U10709 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(P2_U3438) );
  INV_X1 U10710 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9416) );
  MUX2_X1 U10711 ( .A(n9416), .B(n9415), .S(n10245), .Z(n9419) );
  NAND2_X1 U10712 ( .A1(n9417), .A2(n6946), .ZN(n9418) );
  OAI211_X1 U10713 ( .C1(n9420), .C2(n9435), .A(n9419), .B(n9418), .ZN(
        P2_U3435) );
  INV_X1 U10714 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9422) );
  MUX2_X1 U10715 ( .A(n9422), .B(n9421), .S(n10245), .Z(n9425) );
  NAND2_X1 U10716 ( .A1(n9423), .A2(n6946), .ZN(n9424) );
  OAI211_X1 U10717 ( .C1(n9426), .C2(n9435), .A(n9425), .B(n9424), .ZN(
        P2_U3432) );
  MUX2_X1 U10718 ( .A(n10355), .B(n9427), .S(n10245), .Z(n9430) );
  NAND2_X1 U10719 ( .A1(n9428), .A2(n6946), .ZN(n9429) );
  OAI211_X1 U10720 ( .C1(n9431), .C2(n9435), .A(n9430), .B(n9429), .ZN(
        P2_U3429) );
  INV_X1 U10721 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9433) );
  MUX2_X1 U10722 ( .A(n9433), .B(n9432), .S(n10245), .Z(n9434) );
  OAI21_X1 U10723 ( .B1(n9436), .B2(n9435), .A(n9434), .ZN(P2_U3426) );
  MUX2_X1 U10724 ( .A(n9437), .B(P2_REG0_REG_9__SCAN_IN), .S(n10247), .Z(
        P2_U3417) );
  INV_X1 U10725 ( .A(n6676), .ZN(n10108) );
  INV_X1 U10726 ( .A(n9438), .ZN(n9440) );
  NOR4_X1 U10727 ( .A1(n9440), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9439), .A4(
        P2_U3151), .ZN(n9441) );
  AOI21_X1 U10728 ( .B1(n9453), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9441), .ZN(
        n9442) );
  OAI21_X1 U10729 ( .B1(n10108), .B2(n9455), .A(n9442), .ZN(P2_U3264) );
  OAI222_X1 U10730 ( .A1(n9449), .A2(n9445), .B1(n9455), .B2(n9444), .C1(n9443), .C2(P2_U3151), .ZN(P2_U3265) );
  OAI222_X1 U10731 ( .A1(n9449), .A2(n9448), .B1(P2_U3151), .B2(n9446), .C1(
        n9455), .C2(n10110), .ZN(P2_U3266) );
  INV_X1 U10732 ( .A(n6654), .ZN(n10113) );
  AOI21_X1 U10733 ( .B1(n9453), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9450), .ZN(
        n9451) );
  OAI21_X1 U10734 ( .B1(n10113), .B2(n9455), .A(n9451), .ZN(P2_U3267) );
  AOI21_X1 U10735 ( .B1(n9453), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n9452), .ZN(
        n9454) );
  OAI21_X1 U10736 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(P2_U3268) );
  MUX2_X1 U10737 ( .A(n9457), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10738 ( .A(n9458), .ZN(n9462) );
  NAND2_X1 U10739 ( .A1(n4431), .A2(n9461), .ZN(n9459) );
  AOI22_X1 U10740 ( .A1(n9462), .A2(n9461), .B1(n9460), .B2(n9459), .ZN(n9466)
         );
  AOI22_X1 U10741 ( .A1(n9612), .A2(n9567), .B1(n9595), .B2(n9614), .ZN(n9839)
         );
  AOI22_X1 U10742 ( .A1(n9845), .A2(n9538), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9463) );
  OAI21_X1 U10743 ( .B1(n9839), .B2(n9558), .A(n9463), .ZN(n9464) );
  AOI21_X1 U10744 ( .B1(n9844), .B2(n4405), .A(n9464), .ZN(n9465) );
  OAI21_X1 U10745 ( .B1(n9466), .B2(n9589), .A(n9465), .ZN(P1_U3216) );
  NOR2_X1 U10746 ( .A1(n4925), .A2(n9468), .ZN(n9469) );
  XNOR2_X1 U10747 ( .A(n4535), .B(n9469), .ZN(n9476) );
  AOI22_X1 U10748 ( .A1(n9471), .A2(n9602), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9472) );
  OAI21_X1 U10749 ( .B1(n9473), .B2(n9599), .A(n9472), .ZN(n9474) );
  AOI21_X1 U10750 ( .B1(n10018), .B2(n4405), .A(n9474), .ZN(n9475) );
  OAI21_X1 U10751 ( .B1(n9476), .B2(n9589), .A(n9475), .ZN(P1_U3219) );
  XNOR2_X1 U10752 ( .A(n9478), .B(n9477), .ZN(n9479) );
  XNOR2_X1 U10753 ( .A(n9480), .B(n9479), .ZN(n9486) );
  AND2_X1 U10754 ( .A1(n9616), .A2(n9595), .ZN(n9481) );
  AOI21_X1 U10755 ( .B1(n9614), .B2(n9567), .A(n9481), .ZN(n9868) );
  AOI22_X1 U10756 ( .A1(n9870), .A2(n9538), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9482) );
  OAI21_X1 U10757 ( .B1(n9868), .B2(n9558), .A(n9482), .ZN(n9483) );
  AOI21_X1 U10758 ( .B1(n9876), .B2(n4405), .A(n9483), .ZN(n9485) );
  OAI21_X1 U10759 ( .B1(n9486), .B2(n9589), .A(n9485), .ZN(P1_U3223) );
  XOR2_X1 U10760 ( .A(n9488), .B(n9487), .Z(n9493) );
  AND2_X1 U10761 ( .A1(n9612), .A2(n9595), .ZN(n9489) );
  AOI21_X1 U10762 ( .B1(n9610), .B2(n9567), .A(n9489), .ZN(n9807) );
  NOR2_X1 U10763 ( .A1(n9807), .A2(n9558), .ZN(n9491) );
  OAI22_X1 U10764 ( .A1(n9813), .A2(n9599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10509), .ZN(n9490) );
  AOI211_X1 U10765 ( .C1(n9812), .C2(n4405), .A(n9491), .B(n9490), .ZN(n9492)
         );
  OAI21_X1 U10766 ( .B1(n9493), .B2(n9589), .A(n9492), .ZN(P1_U3225) );
  OAI21_X1 U10767 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  NAND2_X1 U10768 ( .A1(n9497), .A2(n5931), .ZN(n9500) );
  AOI22_X1 U10769 ( .A1(n9619), .A2(n9567), .B1(n9621), .B2(n9595), .ZN(n9931)
         );
  NAND2_X1 U10770 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9689) );
  OAI21_X1 U10771 ( .B1(n9931), .B2(n9558), .A(n9689), .ZN(n9498) );
  AOI21_X1 U10772 ( .B1(n9937), .B2(n9538), .A(n9498), .ZN(n9499) );
  OAI211_X1 U10773 ( .C1(n10097), .C2(n9605), .A(n9500), .B(n9499), .ZN(
        P1_U3226) );
  AND2_X1 U10774 ( .A1(n9534), .A2(n9501), .ZN(n9502) );
  NAND2_X1 U10775 ( .A1(n9533), .A2(n9502), .ZN(n9578) );
  XNOR2_X1 U10776 ( .A(n9578), .B(n9576), .ZN(n9503) );
  NAND2_X1 U10777 ( .A1(n9503), .A2(n9504), .ZN(n9577) );
  OAI21_X1 U10778 ( .B1(n9504), .B2(n9503), .A(n9577), .ZN(n9505) );
  NAND2_X1 U10779 ( .A1(n9505), .A2(n5931), .ZN(n9510) );
  AOI22_X1 U10780 ( .A1(n9506), .A2(n9538), .B1(n4405), .B2(n5228), .ZN(n9509)
         );
  NAND2_X1 U10781 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U10782 ( .A1(n9507), .A2(n9602), .ZN(n9508) );
  NAND4_X1 U10783 ( .A1(n9510), .A2(n9509), .A3(n9654), .A4(n9508), .ZN(
        P1_U3227) );
  AOI21_X1 U10784 ( .B1(n9512), .B2(n9514), .A(n9511), .ZN(n9513) );
  AOI21_X1 U10785 ( .B1(n4508), .B2(n9514), .A(n9513), .ZN(n9518) );
  NOR2_X1 U10786 ( .A1(n9599), .A2(n9914), .ZN(n9516) );
  AOI22_X1 U10787 ( .A1(n9595), .A2(n9620), .B1(n9618), .B2(n9567), .ZN(n9920)
         );
  NAND2_X1 U10788 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9708) );
  OAI21_X1 U10789 ( .B1(n9920), .B2(n9558), .A(n9708), .ZN(n9515) );
  AOI211_X1 U10790 ( .C1(n9917), .C2(n4405), .A(n9516), .B(n9515), .ZN(n9517)
         );
  OAI21_X1 U10791 ( .B1(n9518), .B2(n9589), .A(n9517), .ZN(P1_U3228) );
  OAI21_X1 U10792 ( .B1(n9521), .B2(n9519), .A(n9520), .ZN(n9525) );
  AOI22_X1 U10793 ( .A1(n9611), .A2(n9567), .B1(n9595), .B2(n9613), .ZN(n9827)
         );
  NAND2_X1 U10794 ( .A1(n9991), .A2(n4405), .ZN(n9523) );
  AOI22_X1 U10795 ( .A1(n9822), .A2(n9538), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9522) );
  OAI211_X1 U10796 ( .C1(n9827), .C2(n9558), .A(n9523), .B(n9522), .ZN(n9524)
         );
  AOI21_X1 U10797 ( .B1(n9525), .B2(n5931), .A(n9524), .ZN(n9526) );
  INV_X1 U10798 ( .A(n9526), .ZN(P1_U3229) );
  NAND2_X1 U10799 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  AND2_X1 U10800 ( .A1(n9530), .A2(n9529), .ZN(n9532) );
  AOI21_X1 U10801 ( .B1(n9532), .B2(n9531), .A(n9589), .ZN(n9536) );
  AND2_X1 U10802 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  NAND2_X1 U10803 ( .A1(n9536), .A2(n9535), .ZN(n9541) );
  AOI22_X1 U10804 ( .A1(n9537), .A2(n9602), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n9540) );
  AOI22_X1 U10805 ( .A1(n9538), .A2(n10155), .B1(n4405), .B2(n10156), .ZN(
        n9539) );
  NAND3_X1 U10806 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(P1_U3230) );
  INV_X1 U10807 ( .A(n9542), .ZN(n9544) );
  NAND2_X1 U10808 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  XNOR2_X1 U10809 ( .A(n9546), .B(n9545), .ZN(n9552) );
  NOR2_X1 U10810 ( .A1(n9890), .A2(n9599), .ZN(n9550) );
  AND2_X1 U10811 ( .A1(n9617), .A2(n9595), .ZN(n9547) );
  AOI21_X1 U10812 ( .B1(n9615), .B2(n9567), .A(n9547), .ZN(n9885) );
  OAI22_X1 U10813 ( .A1(n9885), .A2(n9558), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9548), .ZN(n9549) );
  AOI211_X1 U10814 ( .C1(n10014), .C2(n4405), .A(n9550), .B(n9549), .ZN(n9551)
         );
  OAI21_X1 U10815 ( .B1(n9552), .B2(n9589), .A(n9551), .ZN(P1_U3233) );
  NAND2_X1 U10816 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  XOR2_X1 U10817 ( .A(n9556), .B(n9555), .Z(n9562) );
  AND2_X1 U10818 ( .A1(n9615), .A2(n9595), .ZN(n9557) );
  AOI21_X1 U10819 ( .B1(n9613), .B2(n9567), .A(n9557), .ZN(n9852) );
  NOR2_X1 U10820 ( .A1(n9852), .A2(n9558), .ZN(n9560) );
  OAI22_X1 U10821 ( .A1(n9859), .A2(n9599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10505), .ZN(n9559) );
  AOI211_X1 U10822 ( .C1(n9857), .C2(n4405), .A(n9560), .B(n9559), .ZN(n9561)
         );
  OAI21_X1 U10823 ( .B1(n9562), .B2(n9589), .A(n9561), .ZN(P1_U3235) );
  NAND2_X1 U10824 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  XOR2_X1 U10825 ( .A(n9566), .B(n9565), .Z(n9573) );
  NAND2_X1 U10826 ( .A1(n9617), .A2(n9567), .ZN(n9569) );
  NAND2_X1 U10827 ( .A1(n9619), .A2(n9595), .ZN(n9568) );
  NAND2_X1 U10828 ( .A1(n9569), .A2(n9568), .ZN(n9907) );
  AOI22_X1 U10829 ( .A1(n9907), .A2(n9602), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9570) );
  OAI21_X1 U10830 ( .B1(n9901), .B2(n9599), .A(n9570), .ZN(n9571) );
  AOI21_X1 U10831 ( .B1(n10023), .B2(n4405), .A(n9571), .ZN(n9572) );
  OAI21_X1 U10832 ( .B1(n9573), .B2(n9589), .A(n9572), .ZN(P1_U3238) );
  NAND2_X1 U10833 ( .A1(n9575), .A2(n9574), .ZN(n9581) );
  INV_X1 U10834 ( .A(n9576), .ZN(n9579) );
  OAI21_X1 U10835 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9580) );
  XOR2_X1 U10836 ( .A(n9581), .B(n9580), .Z(n9582) );
  NAND2_X1 U10837 ( .A1(n9582), .A2(n5931), .ZN(n9588) );
  AOI22_X1 U10838 ( .A1(n9583), .A2(n9602), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n9587) );
  NAND2_X1 U10839 ( .A1(n4405), .A2(n10145), .ZN(n9586) );
  INV_X1 U10840 ( .A(n10144), .ZN(n9584) );
  OR2_X1 U10841 ( .A1(n9599), .A2(n9584), .ZN(n9585) );
  NAND4_X1 U10842 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(
        P1_U3239) );
  OR2_X1 U10843 ( .A1(n9594), .A2(n9593), .ZN(n9597) );
  NAND2_X1 U10844 ( .A1(n9611), .A2(n9595), .ZN(n9596) );
  NAND2_X1 U10845 ( .A1(n9597), .A2(n9596), .ZN(n9792) );
  INV_X1 U10846 ( .A(n9798), .ZN(n9600) );
  OAI22_X1 U10847 ( .A1(n9600), .A2(n9599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9598), .ZN(n9601) );
  AOI21_X1 U10848 ( .B1(n9792), .B2(n9602), .A(n9601), .ZN(n9603) );
  OAI211_X1 U10849 ( .C1(n9801), .C2(n9605), .A(n9604), .B(n9603), .ZN(
        P1_U3240) );
  MUX2_X1 U10850 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9606), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10851 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9607), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10852 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9608), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10853 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9609), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10854 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9610), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10855 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9611), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10856 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9612), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10857 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9613), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10858 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9614), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10859 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9615), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10860 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9616), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10861 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9617), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10862 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9618), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10863 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9619), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10864 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9620), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10865 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9621), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10866 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9622), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10867 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9623), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10868 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9624), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10869 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9625), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10870 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9626), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10871 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n4609), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10872 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9627), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10873 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9628), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10874 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9629), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10875 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9630), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10876 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n6544), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10877 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9631), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10878 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6474), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10879 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6537), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10880 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6538), .S(P1_U3973), .Z(
        P1_U3554) );
  AOI211_X1 U10881 ( .C1(n9634), .C2(n9633), .A(n9632), .B(n10128), .ZN(n9635)
         );
  INV_X1 U10882 ( .A(n9635), .ZN(n9643) );
  AOI22_X1 U10883 ( .A1(n10122), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9642) );
  NAND2_X1 U10884 ( .A1(n10139), .A2(n9636), .ZN(n9641) );
  OAI211_X1 U10885 ( .C1(n9639), .C2(n9638), .A(n10135), .B(n9637), .ZN(n9640)
         );
  NAND4_X1 U10886 ( .A1(n9643), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(
        P1_U3244) );
  AND2_X1 U10887 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9646) );
  NOR2_X1 U10888 ( .A1(n9745), .A2(n9644), .ZN(n9645) );
  AOI211_X1 U10889 ( .C1(n10122), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9646), .B(
        n9645), .ZN(n9653) );
  OAI211_X1 U10890 ( .C1(n9648), .C2(n9647), .A(n10135), .B(n10132), .ZN(n9652) );
  OAI211_X1 U10891 ( .C1(n9650), .C2(n9649), .A(n9744), .B(n10125), .ZN(n9651)
         );
  NAND3_X1 U10892 ( .A1(n9653), .A2(n9652), .A3(n9651), .ZN(P1_U3246) );
  INV_X1 U10893 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9655) );
  OAI21_X1 U10894 ( .B1(n9749), .B2(n9655), .A(n9654), .ZN(n9656) );
  AOI21_X1 U10895 ( .B1(n9657), .B2(n10139), .A(n9656), .ZN(n9668) );
  OAI211_X1 U10896 ( .C1(n9660), .C2(n9659), .A(n10135), .B(n9658), .ZN(n9667)
         );
  MUX2_X1 U10897 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7236), .S(n9661), .Z(n9664)
         );
  INV_X1 U10898 ( .A(n9662), .ZN(n9663) );
  NAND2_X1 U10899 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  OAI211_X1 U10900 ( .C1(n10127), .C2(n9665), .A(n9744), .B(n9678), .ZN(n9666)
         );
  NAND3_X1 U10901 ( .A1(n9668), .A2(n9667), .A3(n9666), .ZN(P1_U3248) );
  AND2_X1 U10902 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U10903 ( .A1(n9745), .A2(n9669), .ZN(n9670) );
  AOI211_X1 U10904 ( .C1(n10122), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9671), .B(
        n9670), .ZN(n9683) );
  OAI211_X1 U10905 ( .C1(n9674), .C2(n9673), .A(n10135), .B(n9672), .ZN(n9682)
         );
  INV_X1 U10906 ( .A(n9675), .ZN(n9680) );
  NAND3_X1 U10907 ( .A1(n9678), .A2(n9677), .A3(n9676), .ZN(n9679) );
  NAND3_X1 U10908 ( .A1(n9744), .A2(n9680), .A3(n9679), .ZN(n9681) );
  NAND3_X1 U10909 ( .A1(n9683), .A2(n9682), .A3(n9681), .ZN(P1_U3249) );
  NOR2_X1 U10910 ( .A1(n9702), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9710) );
  AOI21_X1 U10911 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9702), .A(n9710), .ZN(
        n9686) );
  NOR2_X1 U10912 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  AND2_X1 U10913 ( .A1(n9687), .A2(n9686), .ZN(n9711) );
  OAI21_X1 U10914 ( .B1(n9688), .B2(n9711), .A(n9744), .ZN(n9701) );
  INV_X1 U10915 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9690) );
  OAI21_X1 U10916 ( .B1(n9749), .B2(n9690), .A(n9689), .ZN(n9691) );
  AOI21_X1 U10917 ( .B1(n9702), .B2(n10139), .A(n9691), .ZN(n9700) );
  NAND2_X1 U10918 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  NAND2_X1 U10919 ( .A1(n9695), .A2(n9694), .ZN(n9698) );
  INV_X1 U10920 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9696) );
  MUX2_X1 U10921 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n9696), .S(n9702), .Z(n9697) );
  NAND2_X1 U10922 ( .A1(n9698), .A2(n9697), .ZN(n9704) );
  OAI211_X1 U10923 ( .C1(n9698), .C2(n9697), .A(n9704), .B(n10135), .ZN(n9699)
         );
  NAND3_X1 U10924 ( .A1(n9701), .A2(n9700), .A3(n9699), .ZN(P1_U3259) );
  MUX2_X1 U10925 ( .A(n9915), .B(P1_REG2_REG_17__SCAN_IN), .S(n9725), .Z(n9707) );
  NAND2_X1 U10926 ( .A1(n9702), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U10927 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  INV_X1 U10928 ( .A(n9727), .ZN(n9705) );
  AOI21_X1 U10929 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9718) );
  INV_X1 U10930 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9709) );
  OAI21_X1 U10931 ( .B1(n9749), .B2(n9709), .A(n9708), .ZN(n9716) );
  NOR2_X1 U10932 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  XNOR2_X1 U10933 ( .A(n9725), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9712) );
  AOI21_X1 U10934 ( .B1(n9713), .B2(n9712), .A(n9721), .ZN(n9714) );
  NOR2_X1 U10935 ( .A1(n9714), .A2(n10128), .ZN(n9715) );
  AOI211_X1 U10936 ( .C1(n10139), .C2(n9725), .A(n9716), .B(n9715), .ZN(n9717)
         );
  OAI21_X1 U10937 ( .B1(n9718), .B2(n9729), .A(n9717), .ZN(P1_U3260) );
  NOR2_X1 U10938 ( .A1(n9725), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9720) );
  XNOR2_X1 U10939 ( .A(n9739), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9719) );
  NOR3_X1 U10940 ( .A1(n9721), .A2(n9720), .A3(n9719), .ZN(n9737) );
  INV_X1 U10941 ( .A(n9737), .ZN(n9723) );
  OAI21_X1 U10942 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9722) );
  NAND3_X1 U10943 ( .A1(n9723), .A2(n9744), .A3(n9722), .ZN(n9736) );
  AND2_X1 U10944 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9724) );
  AOI21_X1 U10945 ( .B1(n10122), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9724), .ZN(
        n9735) );
  OR2_X1 U10946 ( .A1(n9725), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U10947 ( .A1(n9727), .A2(n9726), .ZN(n9731) );
  MUX2_X1 U10948 ( .A(n9728), .B(P1_REG2_REG_18__SCAN_IN), .S(n9739), .Z(n9730) );
  AOI21_X1 U10949 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9732) );
  NAND2_X1 U10950 ( .A1(n9732), .A2(n9741), .ZN(n9734) );
  NAND2_X1 U10951 ( .A1(n10139), .A2(n9739), .ZN(n9733) );
  NAND4_X1 U10952 ( .A1(n9736), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(
        P1_U3261) );
  INV_X1 U10953 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9750) );
  AOI21_X1 U10954 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9739), .A(n9737), .ZN(
        n9738) );
  XNOR2_X1 U10955 ( .A(n9738), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U10956 ( .A1(n9739), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U10957 ( .A1(n9741), .A2(n9740), .ZN(n9742) );
  XNOR2_X1 U10958 ( .A(n9742), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9747) );
  INV_X1 U10959 ( .A(n9747), .ZN(n9743) );
  AOI22_X1 U10960 ( .A1(n9746), .A2(n9744), .B1(n10135), .B2(n9743), .ZN(n9748) );
  NAND2_X1 U10961 ( .A1(n9751), .A2(n9833), .ZN(n9754) );
  AND2_X1 U10962 ( .A1(n9752), .A2(n9951), .ZN(n9756) );
  AOI21_X1 U10963 ( .B1(n10167), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9756), .ZN(
        n9753) );
  OAI211_X1 U10964 ( .C1(n9755), .C2(n9953), .A(n9754), .B(n9753), .ZN(
        P1_U3263) );
  INV_X1 U10965 ( .A(n9756), .ZN(n9758) );
  NAND2_X1 U10966 ( .A1(n10167), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U10967 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  AOI21_X1 U10968 ( .B1(n9760), .B2(n10157), .A(n9759), .ZN(n9761) );
  OAI21_X1 U10969 ( .B1(n9762), .B2(n10160), .A(n9761), .ZN(P1_U3264) );
  NAND2_X1 U10970 ( .A1(n9763), .A2(n10163), .ZN(n9773) );
  INV_X1 U10971 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9764) );
  OAI22_X1 U10972 ( .A1(n9765), .A2(n9913), .B1(n9764), .B2(n9951), .ZN(n9766)
         );
  AOI21_X1 U10973 ( .B1(n9767), .B2(n10157), .A(n9766), .ZN(n9772) );
  NAND2_X1 U10974 ( .A1(n9768), .A2(n9951), .ZN(n9771) );
  NAND2_X1 U10975 ( .A1(n9769), .A2(n9971), .ZN(n9770) );
  NAND4_X1 U10976 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(
        P1_U3265) );
  INV_X1 U10977 ( .A(n9774), .ZN(n9780) );
  NAND2_X1 U10978 ( .A1(n9775), .A2(n9786), .ZN(n9776) );
  INV_X1 U10979 ( .A(n9977), .ZN(n9790) );
  AOI211_X1 U10980 ( .C1(n9782), .C2(n9796), .A(n9949), .B(n6976), .ZN(n9978)
         );
  INV_X1 U10981 ( .A(n9782), .ZN(n10069) );
  AOI22_X1 U10982 ( .A1(n9783), .A2(n10154), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10167), .ZN(n9784) );
  OAI21_X1 U10983 ( .B1(n10069), .B2(n9953), .A(n9784), .ZN(n9785) );
  AOI21_X1 U10984 ( .B1(n9978), .B2(n9971), .A(n9785), .ZN(n9789) );
  XNOR2_X1 U10985 ( .A(n9787), .B(n9786), .ZN(n9979) );
  NAND2_X1 U10986 ( .A1(n9979), .A2(n10163), .ZN(n9788) );
  OAI211_X1 U10987 ( .C1(n9790), .C2(n10167), .A(n9789), .B(n9788), .ZN(
        P1_U3266) );
  XNOR2_X1 U10988 ( .A(n9791), .B(n9795), .ZN(n9793) );
  AOI21_X1 U10989 ( .B1(n9793), .B2(n9964), .A(n9792), .ZN(n9984) );
  XOR2_X1 U10990 ( .A(n9795), .B(n9794), .Z(n9985) );
  INV_X1 U10991 ( .A(n9985), .ZN(n9803) );
  OR2_X1 U10992 ( .A1(n9801), .A2(n9811), .ZN(n9797) );
  AND2_X1 U10993 ( .A1(n9797), .A2(n9796), .ZN(n9982) );
  NAND2_X1 U10994 ( .A1(n9982), .A2(n9833), .ZN(n9800) );
  AOI22_X1 U10995 ( .A1(n9798), .A2(n10154), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10167), .ZN(n9799) );
  OAI211_X1 U10996 ( .C1(n9801), .C2(n9953), .A(n9800), .B(n9799), .ZN(n9802)
         );
  AOI21_X1 U10997 ( .B1(n9803), .B2(n10163), .A(n9802), .ZN(n9804) );
  OAI21_X1 U10998 ( .B1(n10167), .B2(n9984), .A(n9804), .ZN(P1_U3267) );
  OAI211_X1 U10999 ( .C1(n9806), .C2(n9809), .A(n9805), .B(n9964), .ZN(n9808)
         );
  NAND2_X1 U11000 ( .A1(n9808), .A2(n9807), .ZN(n9986) );
  INV_X1 U11001 ( .A(n9986), .ZN(n9819) );
  XNOR2_X1 U11002 ( .A(n9809), .B(n9810), .ZN(n9988) );
  NAND2_X1 U11003 ( .A1(n9988), .A2(n10163), .ZN(n9818) );
  AOI211_X1 U11004 ( .C1(n9812), .C2(n9821), .A(n9949), .B(n9811), .ZN(n9987)
         );
  INV_X1 U11005 ( .A(n9812), .ZN(n10073) );
  INV_X1 U11006 ( .A(n9813), .ZN(n9814) );
  AOI22_X1 U11007 ( .A1(n9814), .A2(n10154), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10167), .ZN(n9815) );
  OAI21_X1 U11008 ( .B1(n10073), .B2(n9953), .A(n9815), .ZN(n9816) );
  AOI21_X1 U11009 ( .B1(n9987), .B2(n9971), .A(n9816), .ZN(n9817) );
  OAI211_X1 U11010 ( .C1(n10167), .C2(n9819), .A(n9818), .B(n9817), .ZN(
        P1_U3268) );
  XNOR2_X1 U11011 ( .A(n9820), .B(n6497), .ZN(n9996) );
  AOI21_X1 U11012 ( .B1(n9991), .B2(n9841), .A(n6589), .ZN(n9993) );
  INV_X1 U11013 ( .A(n9991), .ZN(n9824) );
  AOI22_X1 U11014 ( .A1(n9822), .A2(n10154), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10167), .ZN(n9823) );
  OAI21_X1 U11015 ( .B1(n9824), .B2(n9953), .A(n9823), .ZN(n9832) );
  AOI21_X1 U11016 ( .B1(n9826), .B2(n9825), .A(n9945), .ZN(n9830) );
  INV_X1 U11017 ( .A(n9827), .ZN(n9828) );
  AOI21_X1 U11018 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9995) );
  NOR2_X1 U11019 ( .A1(n9995), .A2(n10167), .ZN(n9831) );
  AOI211_X1 U11020 ( .C1(n9993), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9834)
         );
  OAI21_X1 U11021 ( .B1(n9996), .B2(n9957), .A(n9834), .ZN(P1_U3269) );
  XNOR2_X1 U11022 ( .A(n9835), .B(n9837), .ZN(n9999) );
  INV_X1 U11023 ( .A(n9999), .ZN(n9850) );
  XNOR2_X1 U11024 ( .A(n9836), .B(n9837), .ZN(n9838) );
  NAND2_X1 U11025 ( .A1(n9838), .A2(n9964), .ZN(n9840) );
  NAND2_X1 U11026 ( .A1(n9840), .A2(n9839), .ZN(n9997) );
  INV_X1 U11027 ( .A(n9856), .ZN(n9843) );
  INV_X1 U11028 ( .A(n9841), .ZN(n9842) );
  AOI211_X1 U11029 ( .C1(n9844), .C2(n9843), .A(n9949), .B(n9842), .ZN(n9998)
         );
  NAND2_X1 U11030 ( .A1(n9998), .A2(n9971), .ZN(n9847) );
  AOI22_X1 U11031 ( .A1(n9845), .A2(n10154), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10167), .ZN(n9846) );
  OAI211_X1 U11032 ( .C1(n10078), .C2(n9953), .A(n9847), .B(n9846), .ZN(n9848)
         );
  AOI21_X1 U11033 ( .B1(n9951), .B2(n9997), .A(n9848), .ZN(n9849) );
  OAI21_X1 U11034 ( .B1(n9850), .B2(n9957), .A(n9849), .ZN(P1_U3270) );
  XNOR2_X1 U11035 ( .A(n9851), .B(n9854), .ZN(n9853) );
  OAI21_X1 U11036 ( .B1(n9853), .B2(n9945), .A(n9852), .ZN(n10002) );
  INV_X1 U11037 ( .A(n10002), .ZN(n9864) );
  XNOR2_X1 U11038 ( .A(n9855), .B(n9854), .ZN(n10004) );
  NAND2_X1 U11039 ( .A1(n10004), .A2(n10163), .ZN(n9863) );
  AOI211_X1 U11040 ( .C1(n9857), .C2(n9874), .A(n9949), .B(n9856), .ZN(n10003)
         );
  INV_X1 U11041 ( .A(n9857), .ZN(n10082) );
  NOR2_X1 U11042 ( .A1(n10082), .A2(n9953), .ZN(n9861) );
  OAI22_X1 U11043 ( .A1(n9859), .A2(n9913), .B1(n9858), .B2(n9951), .ZN(n9860)
         );
  AOI211_X1 U11044 ( .C1(n10003), .C2(n9971), .A(n9861), .B(n9860), .ZN(n9862)
         );
  OAI211_X1 U11045 ( .C1(n10167), .C2(n9864), .A(n9863), .B(n9862), .ZN(
        P1_U3271) );
  INV_X1 U11046 ( .A(n9865), .ZN(n9866) );
  AOI21_X1 U11047 ( .B1(n8654), .B2(n9883), .A(n9866), .ZN(n9867) );
  XNOR2_X1 U11048 ( .A(n9867), .B(n9871), .ZN(n9869) );
  OAI21_X1 U11049 ( .B1(n9869), .B2(n9945), .A(n9868), .ZN(n10007) );
  AOI21_X1 U11050 ( .B1(n9870), .B2(n10154), .A(n10007), .ZN(n9881) );
  XNOR2_X1 U11051 ( .A(n9872), .B(n9871), .ZN(n10009) );
  INV_X1 U11052 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U11053 ( .C1(n9876), .C2(n9873), .A(n9949), .B(n9875), .ZN(n10008)
         );
  INV_X1 U11054 ( .A(n10008), .ZN(n9878) );
  AOI22_X1 U11055 ( .A1(n9876), .A2(n10157), .B1(n10167), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9877) );
  OAI21_X1 U11056 ( .B1(n9878), .B2(n10160), .A(n9877), .ZN(n9879) );
  AOI21_X1 U11057 ( .B1(n10009), .B2(n10163), .A(n9879), .ZN(n9880) );
  OAI21_X1 U11058 ( .B1(n9881), .B2(n10167), .A(n9880), .ZN(P1_U3272) );
  XNOR2_X1 U11059 ( .A(n9882), .B(n9883), .ZN(n10016) );
  XNOR2_X1 U11060 ( .A(n9884), .B(n9883), .ZN(n9886) );
  OAI21_X1 U11061 ( .B1(n9886), .B2(n9945), .A(n9885), .ZN(n10012) );
  INV_X1 U11062 ( .A(n9887), .ZN(n9889) );
  INV_X1 U11063 ( .A(n9873), .ZN(n9888) );
  AOI211_X1 U11064 ( .C1(n10014), .C2(n9889), .A(n9949), .B(n9888), .ZN(n10013) );
  NAND2_X1 U11065 ( .A1(n10013), .A2(n9971), .ZN(n9893) );
  INV_X1 U11066 ( .A(n9890), .ZN(n9891) );
  AOI22_X1 U11067 ( .A1(n9891), .A2(n10154), .B1(n10167), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9892) );
  OAI211_X1 U11068 ( .C1(n9894), .C2(n9953), .A(n9893), .B(n9892), .ZN(n9895)
         );
  AOI21_X1 U11069 ( .B1(n10012), .B2(n9951), .A(n9895), .ZN(n9896) );
  OAI21_X1 U11070 ( .B1(n9957), .B2(n10016), .A(n9896), .ZN(P1_U3273) );
  XNOR2_X1 U11071 ( .A(n9897), .B(n9906), .ZN(n10026) );
  INV_X1 U11072 ( .A(n9899), .ZN(n9900) );
  AOI211_X1 U11073 ( .C1(n10023), .C2(n9898), .A(n9949), .B(n9900), .ZN(n10022) );
  INV_X1 U11074 ( .A(n10023), .ZN(n9904) );
  INV_X1 U11075 ( .A(n9901), .ZN(n9902) );
  AOI22_X1 U11076 ( .A1(n10167), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9902), 
        .B2(n10154), .ZN(n9903) );
  OAI21_X1 U11077 ( .B1(n9904), .B2(n9953), .A(n9903), .ZN(n9910) );
  XNOR2_X1 U11078 ( .A(n9905), .B(n9906), .ZN(n9908) );
  AOI21_X1 U11079 ( .B1(n9908), .B2(n9964), .A(n9907), .ZN(n10025) );
  NOR2_X1 U11080 ( .A1(n10025), .A2(n10167), .ZN(n9909) );
  AOI211_X1 U11081 ( .C1(n10022), .C2(n9971), .A(n9910), .B(n9909), .ZN(n9911)
         );
  OAI21_X1 U11082 ( .B1(n10026), .B2(n9957), .A(n9911), .ZN(P1_U3275) );
  XOR2_X1 U11083 ( .A(n9912), .B(n9919), .Z(n10029) );
  NAND2_X1 U11084 ( .A1(n10029), .A2(n10163), .ZN(n9927) );
  OAI22_X1 U11085 ( .A1(n9951), .A2(n9915), .B1(n9914), .B2(n9913), .ZN(n9916)
         );
  AOI21_X1 U11086 ( .B1(n9917), .B2(n10157), .A(n9916), .ZN(n9926) );
  XNOR2_X1 U11087 ( .A(n9918), .B(n9919), .ZN(n9921) );
  OAI21_X1 U11088 ( .B1(n9921), .B2(n9945), .A(n9920), .ZN(n10027) );
  NAND2_X1 U11089 ( .A1(n10027), .A2(n9951), .ZN(n9925) );
  OR2_X1 U11090 ( .A1(n9922), .A2(n10092), .ZN(n9923) );
  AND3_X1 U11091 ( .A1(n9898), .A2(n9923), .A3(n9992), .ZN(n10028) );
  NAND2_X1 U11092 ( .A1(n10028), .A2(n9971), .ZN(n9924) );
  NAND4_X1 U11093 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(
        P1_U3276) );
  NOR2_X1 U11094 ( .A1(n9928), .A2(n9955), .ZN(n9943) );
  NOR2_X1 U11095 ( .A1(n9943), .A2(n9929), .ZN(n9930) );
  XOR2_X1 U11096 ( .A(n9933), .B(n9930), .Z(n9932) );
  OAI21_X1 U11097 ( .B1(n9932), .B2(n9945), .A(n9931), .ZN(n10031) );
  INV_X1 U11098 ( .A(n10031), .ZN(n9942) );
  XOR2_X1 U11099 ( .A(n9934), .B(n9933), .Z(n10033) );
  INV_X1 U11100 ( .A(n9948), .ZN(n9935) );
  AOI211_X1 U11101 ( .C1(n9936), .C2(n9935), .A(n9949), .B(n9922), .ZN(n10032)
         );
  NAND2_X1 U11102 ( .A1(n10032), .A2(n9971), .ZN(n9939) );
  AOI22_X1 U11103 ( .A1(n10167), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9937), 
        .B2(n10154), .ZN(n9938) );
  OAI211_X1 U11104 ( .C1(n10097), .C2(n9953), .A(n9939), .B(n9938), .ZN(n9940)
         );
  AOI21_X1 U11105 ( .B1(n10033), .B2(n10163), .A(n9940), .ZN(n9941) );
  OAI21_X1 U11106 ( .B1(n9942), .B2(n10167), .A(n9941), .ZN(P1_U3277) );
  AOI21_X1 U11107 ( .B1(n9928), .B2(n9955), .A(n9943), .ZN(n9946) );
  OAI21_X1 U11108 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n10037) );
  AOI21_X1 U11109 ( .B1(n9947), .B2(n10154), .A(n10037), .ZN(n9961) );
  AOI211_X1 U11110 ( .C1(n10039), .C2(n9950), .A(n9949), .B(n9948), .ZN(n10038) );
  INV_X1 U11111 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9952) );
  OAI22_X1 U11112 ( .A1(n9954), .A2(n9953), .B1(n9952), .B2(n9951), .ZN(n9959)
         );
  XOR2_X1 U11113 ( .A(n9956), .B(n9955), .Z(n10041) );
  NOR2_X1 U11114 ( .A1(n10041), .A2(n9957), .ZN(n9958) );
  AOI211_X1 U11115 ( .C1(n10038), .C2(n9971), .A(n9959), .B(n9958), .ZN(n9960)
         );
  OAI21_X1 U11116 ( .B1(n9961), .B2(n10167), .A(n9960), .ZN(P1_U3278) );
  XOR2_X1 U11117 ( .A(n9962), .B(n9968), .Z(n9965) );
  AOI21_X1 U11118 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n10060) );
  MUX2_X1 U11119 ( .A(n10060), .B(n7562), .S(n10167), .Z(n9976) );
  AOI22_X1 U11120 ( .A1(n10053), .A2(n10157), .B1(n10154), .B2(n9966), .ZN(
        n9975) );
  NAND2_X1 U11121 ( .A1(n9967), .A2(n9968), .ZN(n10054) );
  NAND3_X1 U11122 ( .A1(n10056), .A2(n10054), .A3(n10163), .ZN(n9974) );
  OAI21_X1 U11123 ( .B1(n4503), .B2(n9969), .A(n9992), .ZN(n9970) );
  INV_X1 U11124 ( .A(n10057), .ZN(n9972) );
  NAND2_X1 U11125 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  NAND4_X1 U11126 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(
        P1_U3281) );
  MUX2_X1 U11127 ( .A(n10456), .B(n10066), .S(n10194), .Z(n9980) );
  AOI22_X1 U11128 ( .A1(n9982), .A2(n9992), .B1(n10181), .B2(n9981), .ZN(n9983) );
  OAI211_X1 U11129 ( .C1(n9985), .C2(n10185), .A(n9984), .B(n9983), .ZN(n10070) );
  MUX2_X1 U11130 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10070), .S(n10194), .Z(
        P1_U3548) );
  INV_X1 U11131 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9989) );
  AOI211_X1 U11132 ( .C1(n9988), .C2(n10055), .A(n9987), .B(n9986), .ZN(n10071) );
  MUX2_X1 U11133 ( .A(n9989), .B(n10071), .S(n10194), .Z(n9990) );
  OAI21_X1 U11134 ( .B1(n10073), .B2(n10036), .A(n9990), .ZN(P1_U3547) );
  AOI22_X1 U11135 ( .A1(n9993), .A2(n9992), .B1(n10181), .B2(n9991), .ZN(n9994) );
  OAI211_X1 U11136 ( .C1(n9996), .C2(n10185), .A(n9995), .B(n9994), .ZN(n10074) );
  MUX2_X1 U11137 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10074), .S(n10194), .Z(
        P1_U3546) );
  INV_X1 U11138 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10000) );
  AOI211_X1 U11139 ( .C1(n9999), .C2(n10055), .A(n9998), .B(n9997), .ZN(n10075) );
  MUX2_X1 U11140 ( .A(n10000), .B(n10075), .S(n10194), .Z(n10001) );
  OAI21_X1 U11141 ( .B1(n10078), .B2(n10036), .A(n10001), .ZN(P1_U3545) );
  INV_X1 U11142 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10005) );
  AOI211_X1 U11143 ( .C1(n10004), .C2(n10055), .A(n10003), .B(n10002), .ZN(
        n10079) );
  MUX2_X1 U11144 ( .A(n10005), .B(n10079), .S(n10194), .Z(n10006) );
  OAI21_X1 U11145 ( .B1(n10082), .B2(n10036), .A(n10006), .ZN(P1_U3544) );
  INV_X1 U11146 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10010) );
  AOI211_X1 U11147 ( .C1(n10055), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10083) );
  MUX2_X1 U11148 ( .A(n10010), .B(n10083), .S(n10194), .Z(n10011) );
  OAI21_X1 U11149 ( .B1(n10085), .B2(n10036), .A(n10011), .ZN(P1_U3543) );
  AOI211_X1 U11150 ( .C1(n10181), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        n10015) );
  OAI21_X1 U11151 ( .B1(n10185), .B2(n10016), .A(n10015), .ZN(n10086) );
  MUX2_X1 U11152 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10086), .S(n10194), .Z(
        P1_U3542) );
  AOI21_X1 U11153 ( .B1(n10181), .B2(n10018), .A(n10017), .ZN(n10019) );
  OAI211_X1 U11154 ( .C1(n10021), .C2(n10185), .A(n10020), .B(n10019), .ZN(
        n10087) );
  MUX2_X1 U11155 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10087), .S(n10194), .Z(
        P1_U3541) );
  AOI21_X1 U11156 ( .B1(n10181), .B2(n10023), .A(n10022), .ZN(n10024) );
  OAI211_X1 U11157 ( .C1(n10026), .C2(n10185), .A(n10025), .B(n10024), .ZN(
        n10088) );
  MUX2_X1 U11158 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10088), .S(n10194), .Z(
        P1_U3540) );
  INV_X1 U11159 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10503) );
  AOI211_X1 U11160 ( .C1(n10029), .C2(n10055), .A(n10028), .B(n10027), .ZN(
        n10089) );
  MUX2_X1 U11161 ( .A(n10503), .B(n10089), .S(n10194), .Z(n10030) );
  OAI21_X1 U11162 ( .B1(n10092), .B2(n10036), .A(n10030), .ZN(P1_U3539) );
  INV_X1 U11163 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10034) );
  AOI211_X1 U11164 ( .C1(n10033), .C2(n10055), .A(n10032), .B(n10031), .ZN(
        n10093) );
  MUX2_X1 U11165 ( .A(n10034), .B(n10093), .S(n10194), .Z(n10035) );
  OAI21_X1 U11166 ( .B1(n10097), .B2(n10036), .A(n10035), .ZN(P1_U3538) );
  AOI211_X1 U11167 ( .C1(n10181), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10040) );
  OAI21_X1 U11168 ( .B1(n10185), .B2(n10041), .A(n10040), .ZN(n10098) );
  MUX2_X1 U11169 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10098), .S(n10194), .Z(
        P1_U3537) );
  NAND2_X1 U11170 ( .A1(n10042), .A2(n10181), .ZN(n10044) );
  OAI211_X1 U11171 ( .C1(n10045), .C2(n10170), .A(n10044), .B(n10043), .ZN(
        n10046) );
  MUX2_X1 U11172 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10099), .S(n10194), .Z(
        P1_U3536) );
  AOI21_X1 U11173 ( .B1(n10181), .B2(n10049), .A(n10048), .ZN(n10050) );
  OAI211_X1 U11174 ( .C1(n10185), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        n10100) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10100), .S(n10194), .Z(
        P1_U3535) );
  NAND2_X1 U11176 ( .A1(n10053), .A2(n10181), .ZN(n10059) );
  NAND3_X1 U11177 ( .A1(n10056), .A2(n10055), .A3(n10054), .ZN(n10058) );
  NAND4_X1 U11178 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10101) );
  MUX2_X1 U11179 ( .A(n10101), .B(P1_REG1_REG_12__SCAN_IN), .S(n10192), .Z(
        P1_U3534) );
  AOI21_X1 U11180 ( .B1(n10181), .B2(n10062), .A(n10061), .ZN(n10063) );
  OAI211_X1 U11181 ( .C1(n10065), .C2(n10170), .A(n10064), .B(n10063), .ZN(
        n10102) );
  MUX2_X1 U11182 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10102), .S(n10194), .Z(
        P1_U3533) );
  INV_X1 U11183 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U11184 ( .A(n10067), .B(n10066), .S(n10189), .Z(n10068) );
  MUX2_X1 U11185 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10070), .S(n10189), .Z(
        P1_U3516) );
  MUX2_X1 U11186 ( .A(n10406), .B(n10071), .S(n10189), .Z(n10072) );
  OAI21_X1 U11187 ( .B1(n10073), .B2(n10096), .A(n10072), .ZN(P1_U3515) );
  MUX2_X1 U11188 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10074), .S(n10189), .Z(
        P1_U3514) );
  INV_X1 U11189 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10076) );
  MUX2_X1 U11190 ( .A(n10076), .B(n10075), .S(n10189), .Z(n10077) );
  OAI21_X1 U11191 ( .B1(n10078), .B2(n10096), .A(n10077), .ZN(P1_U3513) );
  INV_X1 U11192 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U11193 ( .A(n10080), .B(n10079), .S(n10189), .Z(n10081) );
  OAI21_X1 U11194 ( .B1(n10082), .B2(n10096), .A(n10081), .ZN(P1_U3512) );
  MUX2_X1 U11195 ( .A(n10537), .B(n10083), .S(n10189), .Z(n10084) );
  OAI21_X1 U11196 ( .B1(n10085), .B2(n10096), .A(n10084), .ZN(P1_U3511) );
  MUX2_X1 U11197 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10086), .S(n10189), .Z(
        P1_U3510) );
  MUX2_X1 U11198 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10087), .S(n10189), .Z(
        P1_U3509) );
  MUX2_X1 U11199 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10088), .S(n10189), .Z(
        P1_U3507) );
  INV_X1 U11200 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U11201 ( .A(n10090), .B(n10089), .S(n10189), .Z(n10091) );
  OAI21_X1 U11202 ( .B1(n10092), .B2(n10096), .A(n10091), .ZN(P1_U3504) );
  INV_X1 U11203 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10094) );
  MUX2_X1 U11204 ( .A(n10094), .B(n10093), .S(n10189), .Z(n10095) );
  OAI21_X1 U11205 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(P1_U3501) );
  MUX2_X1 U11206 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10098), .S(n10189), .Z(
        P1_U3498) );
  MUX2_X1 U11207 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10099), .S(n10189), .Z(
        P1_U3495) );
  MUX2_X1 U11208 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10100), .S(n10189), .Z(
        P1_U3492) );
  MUX2_X1 U11209 ( .A(n10101), .B(P1_REG0_REG_12__SCAN_IN), .S(n10187), .Z(
        P1_U3489) );
  MUX2_X1 U11210 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10102), .S(n10189), .Z(
        P1_U3486) );
  MUX2_X1 U11211 ( .A(n10103), .B(P1_D_REG_0__SCAN_IN), .S(n10169), .Z(
        P1_U3439) );
  NOR4_X1 U11212 ( .A1(n10104), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5217), .A4(
        P1_U3086), .ZN(n10105) );
  AOI21_X1 U11213 ( .B1(n10106), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10105), 
        .ZN(n10107) );
  OAI21_X1 U11214 ( .B1(n10108), .B2(n10114), .A(n10107), .ZN(P1_U3324) );
  OAI222_X1 U11215 ( .A1(n10115), .A2(n10111), .B1(n10114), .B2(n10110), .C1(
        n10109), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U11216 ( .A1(n10115), .A2(n10588), .B1(n10114), .B2(n10113), .C1(
        n10112), .C2(P1_U3086), .ZN(P1_U3327) );
  MUX2_X1 U11217 ( .A(n10116), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11218 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11219 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11220 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10354) );
  AOI21_X1 U11221 ( .B1(n5304), .B2(n10354), .A(n10117), .ZN(n10118) );
  XNOR2_X1 U11222 ( .A(n10118), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11223 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10122), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10119) );
  OAI21_X1 U11224 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(P1_U3243) );
  AOI22_X1 U11225 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n10122), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(P1_U3086), .ZN(n10142) );
  AND3_X1 U11226 ( .A1(n10125), .A2(n10124), .A3(n10123), .ZN(n10126) );
  NOR3_X1 U11227 ( .A1(n10128), .A2(n10127), .A3(n10126), .ZN(n10137) );
  INV_X1 U11228 ( .A(n10129), .ZN(n10131) );
  NAND3_X1 U11229 ( .A1(n10132), .A2(n10131), .A3(n10130), .ZN(n10133) );
  AND3_X1 U11230 ( .A1(n10135), .A2(n10134), .A3(n10133), .ZN(n10136) );
  AOI211_X1 U11231 ( .C1(n10139), .C2(n10138), .A(n10137), .B(n10136), .ZN(
        n10141) );
  NAND3_X1 U11232 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(P1_U3247) );
  INV_X1 U11233 ( .A(n10143), .ZN(n10150) );
  AOI22_X1 U11234 ( .A1(n10167), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10144), 
        .B2(n10154), .ZN(n10147) );
  NAND2_X1 U11235 ( .A1(n10157), .A2(n10145), .ZN(n10146) );
  OAI211_X1 U11236 ( .C1(n10148), .C2(n10160), .A(n10147), .B(n10146), .ZN(
        n10149) );
  AOI21_X1 U11237 ( .B1(n10150), .B2(n10163), .A(n10149), .ZN(n10151) );
  OAI21_X1 U11238 ( .B1(n10167), .B2(n10152), .A(n10151), .ZN(P1_U3287) );
  INV_X1 U11239 ( .A(n10153), .ZN(n10164) );
  AOI22_X1 U11240 ( .A1(n10167), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10155), 
        .B2(n10154), .ZN(n10159) );
  NAND2_X1 U11241 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  OAI211_X1 U11242 ( .C1(n10161), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n10162) );
  AOI21_X1 U11243 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10165) );
  OAI21_X1 U11244 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(P1_U3289) );
  NOR2_X1 U11245 ( .A1(n10168), .A2(n10407), .ZN(P1_U3294) );
  AND2_X1 U11246 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10169), .ZN(P1_U3295) );
  INV_X1 U11247 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10484) );
  NOR2_X1 U11248 ( .A1(n10168), .A2(n10484), .ZN(P1_U3296) );
  AND2_X1 U11249 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10169), .ZN(P1_U3297) );
  AND2_X1 U11250 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10169), .ZN(P1_U3298) );
  AND2_X1 U11251 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10169), .ZN(P1_U3299) );
  AND2_X1 U11252 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10169), .ZN(P1_U3300) );
  AND2_X1 U11253 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10169), .ZN(P1_U3301) );
  AND2_X1 U11254 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10169), .ZN(P1_U3302) );
  INV_X1 U11255 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U11256 ( .A1(n10168), .A2(n10563), .ZN(P1_U3303) );
  NOR2_X1 U11257 ( .A1(n10168), .A2(n10533), .ZN(P1_U3304) );
  AND2_X1 U11258 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10169), .ZN(P1_U3305) );
  NOR2_X1 U11259 ( .A1(n10168), .A2(n10414), .ZN(P1_U3306) );
  AND2_X1 U11260 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10169), .ZN(P1_U3307) );
  AND2_X1 U11261 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10169), .ZN(P1_U3308) );
  NOR2_X1 U11262 ( .A1(n10168), .A2(n10470), .ZN(P1_U3309) );
  AND2_X1 U11263 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10169), .ZN(P1_U3310) );
  AND2_X1 U11264 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10169), .ZN(P1_U3311) );
  AND2_X1 U11265 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10169), .ZN(P1_U3312) );
  INV_X1 U11266 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10459) );
  NOR2_X1 U11267 ( .A1(n10168), .A2(n10459), .ZN(P1_U3313) );
  INV_X1 U11268 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10502) );
  NOR2_X1 U11269 ( .A1(n10168), .A2(n10502), .ZN(P1_U3314) );
  NOR2_X1 U11270 ( .A1(n10168), .A2(n10474), .ZN(P1_U3315) );
  AND2_X1 U11271 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10169), .ZN(P1_U3316) );
  AND2_X1 U11272 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10169), .ZN(P1_U3317) );
  INV_X1 U11273 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10442) );
  NOR2_X1 U11274 ( .A1(n10168), .A2(n10442), .ZN(P1_U3318) );
  AND2_X1 U11275 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10169), .ZN(P1_U3319) );
  NOR2_X1 U11276 ( .A1(n10168), .A2(n10546), .ZN(P1_U3320) );
  AND2_X1 U11277 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10169), .ZN(P1_U3321) );
  INV_X1 U11278 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10425) );
  NOR2_X1 U11279 ( .A1(n10168), .A2(n10425), .ZN(P1_U3322) );
  AND2_X1 U11280 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10169), .ZN(P1_U3323) );
  INV_X1 U11281 ( .A(n10170), .ZN(n10178) );
  INV_X1 U11282 ( .A(n10181), .ZN(n10172) );
  OAI21_X1 U11283 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10176) );
  INV_X1 U11284 ( .A(n10174), .ZN(n10175) );
  AOI211_X1 U11285 ( .C1(n10178), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10191) );
  INV_X1 U11286 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U11287 ( .A1(n10189), .A2(n10191), .B1(n10439), .B2(n10187), .ZN(
        P1_U3456) );
  AOI21_X1 U11288 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(n10182) );
  OAI211_X1 U11289 ( .C1(n10185), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        n10186) );
  INV_X1 U11290 ( .A(n10186), .ZN(n10193) );
  INV_X1 U11291 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U11292 ( .A1(n10189), .A2(n10193), .B1(n10188), .B2(n10187), .ZN(
        P1_U3462) );
  AOI22_X1 U11293 ( .A1(n10194), .A2(n10191), .B1(n10190), .B2(n10192), .ZN(
        P1_U3523) );
  AOI22_X1 U11294 ( .A1(n10194), .A2(n10193), .B1(n7234), .B2(n10192), .ZN(
        P1_U3525) );
  XNOR2_X1 U11295 ( .A(n10195), .B(n10197), .ZN(n10208) );
  XNOR2_X1 U11296 ( .A(n10197), .B(n10196), .ZN(n10201) );
  AOI222_X1 U11297 ( .A1(n10202), .A2(n10201), .B1(n10200), .B2(n10199), .C1(
        n10198), .C2(n9236), .ZN(n10215) );
  AOI22_X1 U11298 ( .A1(n10205), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n10204), 
        .B2(n10203), .ZN(n10206) );
  OAI211_X1 U11299 ( .C1(n10207), .C2(n10208), .A(n10215), .B(n10206), .ZN(
        n10210) );
  INV_X1 U11300 ( .A(n10208), .ZN(n10218) );
  AOI22_X1 U11301 ( .A1(n10210), .A2(n10212), .B1(n10218), .B2(n10209), .ZN(
        n10211) );
  OAI21_X1 U11302 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(P2_U3231) );
  INV_X1 U11303 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U11304 ( .A1(n10247), .A2(n10413), .B1(n10214), .B2(n10245), .ZN(
        P2_U3393) );
  INV_X1 U11305 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10440) );
  OAI21_X1 U11306 ( .B1(n10216), .B2(n10239), .A(n10215), .ZN(n10217) );
  AOI21_X1 U11307 ( .B1(n10218), .B2(n10238), .A(n10217), .ZN(n10249) );
  AOI22_X1 U11308 ( .A1(n10247), .A2(n10440), .B1(n10249), .B2(n10245), .ZN(
        P2_U3396) );
  INV_X1 U11309 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10224) );
  INV_X1 U11310 ( .A(n10219), .ZN(n10223) );
  OAI21_X1 U11311 ( .B1(n10221), .B2(n10239), .A(n10220), .ZN(n10222) );
  AOI21_X1 U11312 ( .B1(n10223), .B2(n10238), .A(n10222), .ZN(n10251) );
  AOI22_X1 U11313 ( .A1(n10247), .A2(n10224), .B1(n10251), .B2(n10245), .ZN(
        P2_U3399) );
  INV_X1 U11314 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10230) );
  INV_X1 U11315 ( .A(n10225), .ZN(n10229) );
  OAI21_X1 U11316 ( .B1(n10227), .B2(n10239), .A(n10226), .ZN(n10228) );
  AOI21_X1 U11317 ( .B1(n10229), .B2(n10238), .A(n10228), .ZN(n10253) );
  AOI22_X1 U11318 ( .A1(n10247), .A2(n10230), .B1(n10253), .B2(n10245), .ZN(
        P2_U3402) );
  INV_X1 U11319 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U11320 ( .A1(n10231), .A2(n10239), .ZN(n10233) );
  AOI211_X1 U11321 ( .C1(n10235), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10255) );
  AOI22_X1 U11322 ( .A1(n10247), .A2(n10236), .B1(n10255), .B2(n10245), .ZN(
        P2_U3405) );
  INV_X1 U11323 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10246) );
  INV_X1 U11324 ( .A(n10237), .ZN(n10244) );
  INV_X1 U11325 ( .A(n10238), .ZN(n10241) );
  OAI22_X1 U11326 ( .A1(n10242), .A2(n10241), .B1(n10240), .B2(n10239), .ZN(
        n10243) );
  NOR2_X1 U11327 ( .A1(n10244), .A2(n10243), .ZN(n10256) );
  AOI22_X1 U11328 ( .A1(n10247), .A2(n10246), .B1(n10256), .B2(n10245), .ZN(
        P2_U3408) );
  AOI22_X1 U11329 ( .A1(n10257), .A2(n10249), .B1(n10248), .B2(n9273), .ZN(
        P2_U3461) );
  AOI22_X1 U11330 ( .A1(n10257), .A2(n10251), .B1(n10250), .B2(n9273), .ZN(
        P2_U3462) );
  AOI22_X1 U11331 ( .A1(n10257), .A2(n10253), .B1(n10252), .B2(n9273), .ZN(
        P2_U3463) );
  AOI22_X1 U11332 ( .A1(n10257), .A2(n10255), .B1(n10254), .B2(n9273), .ZN(
        P2_U3464) );
  AOI22_X1 U11333 ( .A1(n10257), .A2(n10256), .B1(n7042), .B2(n9273), .ZN(
        P2_U3465) );
  NAND3_X1 U11334 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10262) );
  AOI21_X1 U11335 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10264) );
  INV_X1 U11336 ( .A(n10264), .ZN(n10258) );
  NAND2_X1 U11337 ( .A1(n10262), .A2(n10258), .ZN(n10259) );
  XNOR2_X1 U11338 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10259), .ZN(ADD_1068_U5)
         );
  NOR2_X1 U11339 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10300) );
  NOR2_X1 U11340 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10298) );
  NOR2_X1 U11341 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10295) );
  NOR2_X1 U11342 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10291) );
  NOR2_X1 U11343 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10289) );
  NAND2_X1 U11344 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10285) );
  XOR2_X1 U11345 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n10315) );
  NAND2_X1 U11346 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10283) );
  INV_X1 U11347 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11348 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n10261), .B2(n10260), .ZN(n10317) );
  INV_X1 U11349 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U11350 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .B1(n10518), .B2(n10281), .ZN(n10319) );
  INV_X1 U11351 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10641) );
  NOR2_X1 U11352 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10270) );
  XNOR2_X1 U11353 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10646) );
  NAND2_X1 U11354 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10268) );
  NOR2_X1 U11355 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10366) );
  AOI21_X1 U11356 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10366), .ZN(n10644) );
  NAND2_X1 U11357 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10266) );
  XOR2_X1 U11358 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10634) );
  OAI21_X1 U11359 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10633) );
  NAND2_X1 U11360 ( .A1(n10634), .A2(n10633), .ZN(n10265) );
  NAND2_X1 U11361 ( .A1(n10266), .A2(n10265), .ZN(n10643) );
  NAND2_X1 U11362 ( .A1(n10644), .A2(n10643), .ZN(n10267) );
  NAND2_X1 U11363 ( .A1(n10268), .A2(n10267), .ZN(n10645) );
  NOR2_X1 U11364 ( .A1(n10646), .A2(n10645), .ZN(n10269) );
  NOR2_X1 U11365 ( .A1(n10270), .A2(n10269), .ZN(n10640) );
  NAND2_X1 U11366 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10640), .ZN(n10271) );
  NOR2_X1 U11367 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10640), .ZN(n10639) );
  AOI21_X1 U11368 ( .B1(n10641), .B2(n10271), .A(n10639), .ZN(n10272) );
  NOR2_X1 U11369 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10272), .ZN(n10635) );
  AND2_X1 U11370 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10272), .ZN(n10636) );
  OAI22_X1 U11371 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n10636), .ZN(n10275) );
  INV_X1 U11372 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10273) );
  OAI22_X1 U11373 ( .A1(n10635), .A2(n10275), .B1(n10274), .B2(n10273), .ZN(
        n10276) );
  AOI21_X1 U11374 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10276), .ZN(n10279) );
  OAI22_X1 U11375 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10278)
         );
  OAI22_X1 U11376 ( .A1(n10279), .A2(n10278), .B1(n10277), .B2(n10594), .ZN(
        n10318) );
  NAND2_X1 U11377 ( .A1(n10319), .A2(n10318), .ZN(n10280) );
  OAI21_X1 U11378 ( .B1(n10518), .B2(n10281), .A(n10280), .ZN(n10316) );
  NAND2_X1 U11379 ( .A1(n10317), .A2(n10316), .ZN(n10282) );
  NAND2_X1 U11380 ( .A1(n10283), .A2(n10282), .ZN(n10314) );
  NAND2_X1 U11381 ( .A1(n10315), .A2(n10314), .ZN(n10284) );
  NAND2_X1 U11382 ( .A1(n10285), .A2(n10284), .ZN(n10313) );
  INV_X1 U11383 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11384 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10287), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10286), .ZN(n10312) );
  NOR2_X1 U11385 ( .A1(n10313), .A2(n10312), .ZN(n10288) );
  NOR2_X1 U11386 ( .A1(n10289), .A2(n10288), .ZN(n10311) );
  XNOR2_X1 U11387 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10310) );
  NOR2_X1 U11388 ( .A1(n10311), .A2(n10310), .ZN(n10290) );
  NOR2_X1 U11389 ( .A1(n10291), .A2(n10290), .ZN(n10309) );
  INV_X1 U11390 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U11391 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10293), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10292), .ZN(n10308) );
  NOR2_X1 U11392 ( .A1(n10309), .A2(n10308), .ZN(n10294) );
  NOR2_X1 U11393 ( .A1(n10295), .A2(n10294), .ZN(n10307) );
  INV_X1 U11394 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U11395 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9690), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10296), .ZN(n10306) );
  NOR2_X1 U11396 ( .A1(n10307), .A2(n10306), .ZN(n10297) );
  NOR2_X1 U11397 ( .A1(n10298), .A2(n10297), .ZN(n10305) );
  XNOR2_X1 U11398 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10304) );
  NOR2_X1 U11399 ( .A1(n10305), .A2(n10304), .ZN(n10299) );
  NOR2_X1 U11400 ( .A1(n10300), .A2(n10299), .ZN(n10301) );
  AND2_X1 U11401 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10301), .ZN(n10628) );
  NOR2_X1 U11402 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10301), .ZN(n10630) );
  NOR2_X1 U11403 ( .A1(n10628), .A2(n10630), .ZN(n10303) );
  INV_X1 U11404 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10302) );
  XNOR2_X1 U11405 ( .A(n10303), .B(n10302), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11406 ( .A(n10305), .B(n10304), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11407 ( .A(n10307), .B(n10306), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11408 ( .A(n10309), .B(n10308), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11409 ( .A(n10311), .B(n10310), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11410 ( .A(n10313), .B(n10312), .ZN(ADD_1068_U60) );
  XOR2_X1 U11411 ( .A(n10315), .B(n10314), .Z(ADD_1068_U61) );
  XOR2_X1 U11412 ( .A(n10317), .B(n10316), .Z(ADD_1068_U62) );
  XOR2_X1 U11413 ( .A(n10319), .B(n10318), .Z(ADD_1068_U63) );
  NOR4_X1 U11414 ( .A1(n10321), .A2(n10320), .A3(P1_REG2_REG_22__SCAN_IN), 
        .A4(P2_REG0_REG_1__SCAN_IN), .ZN(n10322) );
  NAND3_X1 U11415 ( .A1(n10322), .A2(P2_REG0_REG_0__SCAN_IN), .A3(
        P2_REG0_REG_30__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U11416 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(SI_20_), .A4(SI_19_), .ZN(n10323) );
  NOR3_X1 U11417 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_WR_REG_SCAN_IN), .A3(
        n10323), .ZN(n10331) );
  NAND4_X1 U11418 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_REG2_REG_28__SCAN_IN), 
        .A3(P1_DATAO_REG_13__SCAN_IN), .A4(P2_REG1_REG_8__SCAN_IN), .ZN(n10324) );
  NOR3_X1 U11419 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(n10324), .A3(
        P1_IR_REG_20__SCAN_IN), .ZN(n10326) );
  INV_X1 U11420 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10325) );
  NAND3_X1 U11421 ( .A1(n10326), .A2(P2_IR_REG_20__SCAN_IN), .A3(n10325), .ZN(
        n10329) );
  NAND4_X1 U11422 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), 
        .A3(n10405), .A4(n10406), .ZN(n10328) );
  NAND4_X1 U11423 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), 
        .A3(P1_D_REG_21__SCAN_IN), .A4(n10537), .ZN(n10327) );
  NOR3_X1 U11424 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10330) );
  NAND4_X1 U11425 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(n10331), .A4(n10330), .ZN(n10332) );
  NOR4_X1 U11426 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n10416), .A3(n10333), .A4(
        n10332), .ZN(n10374) );
  INV_X1 U11427 ( .A(n10334), .ZN(n10372) );
  NOR4_X1 U11428 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .A3(n10508), .A4(n10506), .ZN(n10341) );
  INV_X1 U11429 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10510) );
  NOR4_X1 U11430 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), 
        .A3(P2_DATAO_REG_8__SCAN_IN), .A4(n10510), .ZN(n10340) );
  INV_X1 U11431 ( .A(SI_16_), .ZN(n10526) );
  NAND4_X1 U11432 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(P1_REG0_REG_2__SCAN_IN), 
        .A3(n10526), .A4(n10519), .ZN(n10338) );
  INV_X1 U11433 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10593) );
  INV_X1 U11434 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10590) );
  NAND4_X1 U11435 ( .A1(SI_7_), .A2(n10593), .A3(n10592), .A4(n10590), .ZN(
        n10337) );
  NAND4_X1 U11436 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .A3(n10548), .A4(n10534), .ZN(n10336) );
  INV_X1 U11437 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10549) );
  NAND4_X1 U11438 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(n10505), .A3(n10549), 
        .A4(n7234), .ZN(n10335) );
  NOR4_X1 U11439 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  NAND3_X1 U11440 ( .A1(n10341), .A2(n10340), .A3(n10339), .ZN(n10371) );
  INV_X1 U11441 ( .A(SI_10_), .ZN(n10487) );
  NAND4_X1 U11442 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(P2_REG2_REG_19__SCAN_IN), 
        .A3(P1_REG3_REG_2__SCAN_IN), .A4(n10487), .ZN(n10343) );
  NAND4_X1 U11443 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .A3(P1_REG1_REG_7__SCAN_IN), .A4(n10456), .ZN(n10342) );
  NOR4_X1 U11444 ( .A1(n10574), .A2(n10605), .A3(n10343), .A4(n10342), .ZN(
        n10349) );
  NAND4_X1 U11445 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(P1_REG0_REG_9__SCAN_IN), .A4(n10473), .ZN(n10344) );
  NOR2_X1 U11446 ( .A1(n10344), .A2(n9709), .ZN(n10348) );
  INV_X1 U11447 ( .A(SI_30_), .ZN(n10345) );
  NOR4_X1 U11448 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P1_DATAO_REG_0__SCAN_IN), 
        .A3(n10565), .A4(n10345), .ZN(n10347) );
  NOR4_X1 U11449 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .A3(P1_ADDR_REG_10__SCAN_IN), .A4(n10594), .ZN(n10346) );
  NAND4_X1 U11450 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NOR4_X1 U11451 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .A3(P1_IR_REG_23__SCAN_IN), .A4(n10350), .ZN(n10353) );
  NOR2_X1 U11452 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n10352) );
  INV_X1 U11453 ( .A(SI_6_), .ZN(n10351) );
  NAND4_X1 U11454 ( .A1(n10353), .A2(SI_21_), .A3(n10352), .A4(n10351), .ZN(
        n10360) );
  NAND4_X1 U11455 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), 
        .A3(P1_D_REG_3__SCAN_IN), .A4(n10422), .ZN(n10359) );
  NAND4_X1 U11456 ( .A1(n10354), .A2(P2_IR_REG_8__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n10358) );
  INV_X1 U11457 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10356) );
  NAND4_X1 U11458 ( .A1(n10356), .A2(n10355), .A3(n10564), .A4(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10357) );
  NOR4_X1 U11459 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10369) );
  INV_X1 U11460 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10602) );
  NAND4_X1 U11461 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(n5817), .A3(n10588), .A4(
        n10602), .ZN(n10363) );
  NAND4_X1 U11462 ( .A1(n10637), .A2(n10582), .A3(n10489), .A4(
        P2_REG1_REG_30__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U11463 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .A3(P2_D_REG_20__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10361) );
  NOR3_X1 U11464 ( .A1(n10363), .A2(n10362), .A3(n10361), .ZN(n10368) );
  NAND4_X1 U11465 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .A3(n10445), .A4(n9952), .ZN(n10365) );
  NAND4_X1 U11466 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P2_REG0_REG_2__SCAN_IN), 
        .A3(P1_REG1_REG_26__SCAN_IN), .A4(n10439), .ZN(n10364) );
  NOR2_X1 U11467 ( .A1(n10365), .A2(n10364), .ZN(n10367) );
  NAND4_X1 U11468 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10370) );
  NOR3_X1 U11469 ( .A1(n10372), .A2(n10371), .A3(n10370), .ZN(n10373) );
  AOI21_X1 U11470 ( .B1(n10374), .B2(n10373), .A(P2_IR_REG_10__SCAN_IN), .ZN(
        n10624) );
  AOI22_X1 U11471 ( .A1(n10377), .A2(keyinput122), .B1(keyinput78), .B2(n10376), .ZN(n10375) );
  OAI221_X1 U11472 ( .B1(n10377), .B2(keyinput122), .C1(n10376), .C2(
        keyinput78), .A(n10375), .ZN(n10390) );
  AOI22_X1 U11473 ( .A1(n10380), .A2(keyinput75), .B1(keyinput13), .B2(n10379), 
        .ZN(n10378) );
  OAI221_X1 U11474 ( .B1(n10380), .B2(keyinput75), .C1(n10379), .C2(keyinput13), .A(n10378), .ZN(n10389) );
  INV_X1 U11475 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U11476 ( .A1(n10383), .A2(keyinput126), .B1(keyinput37), .B2(n10382), .ZN(n10381) );
  OAI221_X1 U11477 ( .B1(n10383), .B2(keyinput126), .C1(n10382), .C2(
        keyinput37), .A(n10381), .ZN(n10388) );
  INV_X1 U11478 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U11479 ( .A1(n10386), .A2(keyinput41), .B1(n10385), .B2(keyinput94), 
        .ZN(n10384) );
  OAI221_X1 U11480 ( .B1(n10386), .B2(keyinput41), .C1(n10385), .C2(keyinput94), .A(n10384), .ZN(n10387) );
  NOR4_X1 U11481 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10437) );
  AOI22_X1 U11482 ( .A1(n10392), .A2(keyinput116), .B1(keyinput61), .B2(n9858), 
        .ZN(n10391) );
  OAI221_X1 U11483 ( .B1(n10392), .B2(keyinput116), .C1(n9858), .C2(keyinput61), .A(n10391), .ZN(n10403) );
  INV_X1 U11484 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10394) );
  AOI22_X1 U11485 ( .A1(n10395), .A2(keyinput77), .B1(keyinput24), .B2(n10394), 
        .ZN(n10393) );
  OAI221_X1 U11486 ( .B1(n10395), .B2(keyinput77), .C1(n10394), .C2(keyinput24), .A(n10393), .ZN(n10402) );
  XOR2_X1 U11487 ( .A(n10396), .B(keyinput100), .Z(n10400) );
  XNOR2_X1 U11488 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput86), .ZN(n10399) );
  XNOR2_X1 U11489 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput45), .ZN(n10398)
         );
  XNOR2_X1 U11490 ( .A(P2_REG1_REG_25__SCAN_IN), .B(keyinput105), .ZN(n10397)
         );
  NAND4_X1 U11491 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10401) );
  NOR3_X1 U11492 ( .A1(n10403), .A2(n10402), .A3(n10401), .ZN(n10436) );
  AOI22_X1 U11493 ( .A1(n10406), .A2(keyinput56), .B1(n10405), .B2(keyinput97), 
        .ZN(n10404) );
  OAI221_X1 U11494 ( .B1(n10406), .B2(keyinput56), .C1(n10405), .C2(keyinput97), .A(n10404), .ZN(n10411) );
  XNOR2_X1 U11495 ( .A(n10407), .B(keyinput99), .ZN(n10410) );
  XNOR2_X1 U11496 ( .A(n10408), .B(keyinput49), .ZN(n10409) );
  OR3_X1 U11497 ( .A1(n10411), .A2(n10410), .A3(n10409), .ZN(n10420) );
  AOI22_X1 U11498 ( .A1(n10414), .A2(keyinput76), .B1(n10413), .B2(keyinput7), 
        .ZN(n10412) );
  OAI221_X1 U11499 ( .B1(n10414), .B2(keyinput76), .C1(n10413), .C2(keyinput7), 
        .A(n10412), .ZN(n10419) );
  INV_X1 U11500 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U11501 ( .A1(n10417), .A2(keyinput2), .B1(n10416), .B2(keyinput48), 
        .ZN(n10415) );
  OAI221_X1 U11502 ( .B1(n10417), .B2(keyinput2), .C1(n10416), .C2(keyinput48), 
        .A(n10415), .ZN(n10418) );
  NOR3_X1 U11503 ( .A1(n10420), .A2(n10419), .A3(n10418), .ZN(n10435) );
  AOI22_X1 U11504 ( .A1(n10423), .A2(keyinput47), .B1(keyinput93), .B2(n10422), 
        .ZN(n10421) );
  OAI221_X1 U11505 ( .B1(n10423), .B2(keyinput47), .C1(n10422), .C2(keyinput93), .A(n10421), .ZN(n10433) );
  AOI22_X1 U11506 ( .A1(n4739), .A2(keyinput72), .B1(keyinput85), .B2(n10425), 
        .ZN(n10424) );
  OAI221_X1 U11507 ( .B1(n4739), .B2(keyinput72), .C1(n10425), .C2(keyinput85), 
        .A(n10424), .ZN(n10432) );
  INV_X1 U11508 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10426) );
  XOR2_X1 U11509 ( .A(n10426), .B(keyinput1), .Z(n10430) );
  XNOR2_X1 U11510 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput46), .ZN(n10429)
         );
  XNOR2_X1 U11511 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput55), .ZN(n10428) );
  XNOR2_X1 U11512 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput115), .ZN(n10427) );
  NAND4_X1 U11513 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10431) );
  NOR3_X1 U11514 ( .A1(n10433), .A2(n10432), .A3(n10431), .ZN(n10434) );
  NAND4_X1 U11515 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10622) );
  AOI22_X1 U11516 ( .A1(n10440), .A2(keyinput112), .B1(keyinput57), .B2(n10439), .ZN(n10438) );
  OAI221_X1 U11517 ( .B1(n10440), .B2(keyinput112), .C1(n10439), .C2(
        keyinput57), .A(n10438), .ZN(n10451) );
  AOI22_X1 U11518 ( .A1(n10443), .A2(keyinput43), .B1(n10442), .B2(keyinput33), 
        .ZN(n10441) );
  OAI221_X1 U11519 ( .B1(n10443), .B2(keyinput43), .C1(n10442), .C2(keyinput33), .A(n10441), .ZN(n10450) );
  AOI22_X1 U11520 ( .A1(n10445), .A2(keyinput114), .B1(keyinput120), .B2(n9952), .ZN(n10444) );
  OAI221_X1 U11521 ( .B1(n10445), .B2(keyinput114), .C1(n9952), .C2(
        keyinput120), .A(n10444), .ZN(n10449) );
  AOI22_X1 U11522 ( .A1(n5986), .A2(keyinput70), .B1(keyinput31), .B2(n10447), 
        .ZN(n10446) );
  OAI221_X1 U11523 ( .B1(n5986), .B2(keyinput70), .C1(n10447), .C2(keyinput31), 
        .A(n10446), .ZN(n10448) );
  NOR4_X1 U11524 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10500) );
  AOI22_X1 U11525 ( .A1(n10454), .A2(keyinput104), .B1(n10453), .B2(keyinput95), .ZN(n10452) );
  OAI221_X1 U11526 ( .B1(n10454), .B2(keyinput104), .C1(n10453), .C2(
        keyinput95), .A(n10452), .ZN(n10465) );
  AOI22_X1 U11527 ( .A1(n10456), .A2(keyinput92), .B1(n6296), .B2(keyinput8), 
        .ZN(n10455) );
  OAI221_X1 U11528 ( .B1(n10456), .B2(keyinput92), .C1(n6296), .C2(keyinput8), 
        .A(n10455), .ZN(n10464) );
  AOI22_X1 U11529 ( .A1(n6153), .A2(keyinput111), .B1(keyinput68), .B2(n10458), 
        .ZN(n10457) );
  OAI221_X1 U11530 ( .B1(n6153), .B2(keyinput111), .C1(n10458), .C2(keyinput68), .A(n10457), .ZN(n10463) );
  XOR2_X1 U11531 ( .A(n10459), .B(keyinput84), .Z(n10461) );
  XNOR2_X1 U11532 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput14), .ZN(n10460)
         );
  NAND2_X1 U11533 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  NOR4_X1 U11534 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10499) );
  AOI22_X1 U11535 ( .A1(n10468), .A2(keyinput113), .B1(keyinput69), .B2(n10467), .ZN(n10466) );
  OAI221_X1 U11536 ( .B1(n10468), .B2(keyinput113), .C1(n10467), .C2(
        keyinput69), .A(n10466), .ZN(n10481) );
  AOI22_X1 U11537 ( .A1(n10471), .A2(keyinput28), .B1(n10470), .B2(keyinput117), .ZN(n10469) );
  OAI221_X1 U11538 ( .B1(n10471), .B2(keyinput28), .C1(n10470), .C2(
        keyinput117), .A(n10469), .ZN(n10480) );
  AOI22_X1 U11539 ( .A1(n10474), .A2(keyinput60), .B1(keyinput16), .B2(n10473), 
        .ZN(n10472) );
  OAI221_X1 U11540 ( .B1(n10474), .B2(keyinput60), .C1(n10473), .C2(keyinput16), .A(n10472), .ZN(n10479) );
  INV_X1 U11541 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U11542 ( .A1(n10477), .A2(keyinput64), .B1(n10476), .B2(keyinput125), .ZN(n10475) );
  OAI221_X1 U11543 ( .B1(n10477), .B2(keyinput64), .C1(n10476), .C2(
        keyinput125), .A(n10475), .ZN(n10478) );
  NOR4_X1 U11544 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10498) );
  AOI22_X1 U11545 ( .A1(n10484), .A2(keyinput87), .B1(keyinput80), .B2(n10483), 
        .ZN(n10482) );
  OAI221_X1 U11546 ( .B1(n10484), .B2(keyinput87), .C1(n10483), .C2(keyinput80), .A(n10482), .ZN(n10496) );
  AOI22_X1 U11547 ( .A1(n10487), .A2(keyinput3), .B1(keyinput102), .B2(n10486), 
        .ZN(n10485) );
  OAI221_X1 U11548 ( .B1(n10487), .B2(keyinput3), .C1(n10486), .C2(keyinput102), .A(n10485), .ZN(n10495) );
  INV_X1 U11549 ( .A(SI_21_), .ZN(n10490) );
  AOI22_X1 U11550 ( .A1(n10490), .A2(keyinput6), .B1(keyinput74), .B2(n10489), 
        .ZN(n10488) );
  OAI221_X1 U11551 ( .B1(n10490), .B2(keyinput6), .C1(n10489), .C2(keyinput74), 
        .A(n10488), .ZN(n10494) );
  XNOR2_X1 U11552 ( .A(P2_REG0_REG_13__SCAN_IN), .B(keyinput118), .ZN(n10492)
         );
  XNOR2_X1 U11553 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput35), .ZN(n10491) );
  NAND2_X1 U11554 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  NOR4_X1 U11555 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10497) );
  NAND4_X1 U11556 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10621) );
  AOI22_X1 U11557 ( .A1(n10503), .A2(keyinput27), .B1(n10502), .B2(keyinput123), .ZN(n10501) );
  OAI221_X1 U11558 ( .B1(n10503), .B2(keyinput27), .C1(n10502), .C2(
        keyinput123), .A(n10501), .ZN(n10516) );
  AOI22_X1 U11559 ( .A1(n10506), .A2(keyinput58), .B1(n10505), .B2(keyinput90), 
        .ZN(n10504) );
  OAI221_X1 U11560 ( .B1(n10506), .B2(keyinput58), .C1(n10505), .C2(keyinput90), .A(n10504), .ZN(n10515) );
  AOI22_X1 U11561 ( .A1(n10509), .A2(keyinput39), .B1(n10508), .B2(keyinput71), 
        .ZN(n10507) );
  OAI221_X1 U11562 ( .B1(n10509), .B2(keyinput39), .C1(n10508), .C2(keyinput71), .A(n10507), .ZN(n10514) );
  XOR2_X1 U11563 ( .A(n10510), .B(keyinput9), .Z(n10512) );
  XNOR2_X1 U11564 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput108), .ZN(n10511)
         );
  NAND2_X1 U11565 ( .A1(n10512), .A2(n10511), .ZN(n10513) );
  NOR4_X1 U11566 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10561) );
  AOI22_X1 U11567 ( .A1(n10519), .A2(keyinput50), .B1(keyinput91), .B2(n10518), 
        .ZN(n10517) );
  OAI221_X1 U11568 ( .B1(n10519), .B2(keyinput50), .C1(n10518), .C2(keyinput91), .A(n10517), .ZN(n10531) );
  AOI22_X1 U11569 ( .A1(n9064), .A2(keyinput19), .B1(keyinput44), .B2(n10521), 
        .ZN(n10520) );
  OAI221_X1 U11570 ( .B1(n9064), .B2(keyinput19), .C1(n10521), .C2(keyinput44), 
        .A(n10520), .ZN(n10530) );
  AOI22_X1 U11571 ( .A1(n10524), .A2(keyinput12), .B1(keyinput54), .B2(n10523), 
        .ZN(n10522) );
  OAI221_X1 U11572 ( .B1(n10524), .B2(keyinput12), .C1(n10523), .C2(keyinput54), .A(n10522), .ZN(n10529) );
  AOI22_X1 U11573 ( .A1(n10527), .A2(keyinput15), .B1(n10526), .B2(keyinput63), 
        .ZN(n10525) );
  OAI221_X1 U11574 ( .B1(n10527), .B2(keyinput15), .C1(n10526), .C2(keyinput63), .A(n10525), .ZN(n10528) );
  NOR4_X1 U11575 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10560) );
  AOI22_X1 U11576 ( .A1(n10534), .A2(keyinput62), .B1(n10533), .B2(keyinput67), 
        .ZN(n10532) );
  OAI221_X1 U11577 ( .B1(n10534), .B2(keyinput62), .C1(n10533), .C2(keyinput67), .A(n10532), .ZN(n10544) );
  AOI22_X1 U11578 ( .A1(n10537), .A2(keyinput124), .B1(n10536), .B2(keyinput98), .ZN(n10535) );
  OAI221_X1 U11579 ( .B1(n10537), .B2(keyinput124), .C1(n10536), .C2(
        keyinput98), .A(n10535), .ZN(n10543) );
  INV_X1 U11580 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U11581 ( .A1(n10637), .A2(keyinput73), .B1(n6325), .B2(keyinput36), 
        .ZN(n10538) );
  OAI221_X1 U11582 ( .B1(n10637), .B2(keyinput73), .C1(n6325), .C2(keyinput36), 
        .A(n10538), .ZN(n10542) );
  XOR2_X1 U11583 ( .A(n9044), .B(keyinput20), .Z(n10540) );
  XNOR2_X1 U11584 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput25), .ZN(n10539) );
  NAND2_X1 U11585 ( .A1(n10540), .A2(n10539), .ZN(n10541) );
  NOR4_X1 U11586 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10559) );
  AOI22_X1 U11587 ( .A1(n5923), .A2(keyinput107), .B1(keyinput38), .B2(n10546), 
        .ZN(n10545) );
  OAI221_X1 U11588 ( .B1(n5923), .B2(keyinput107), .C1(n10546), .C2(keyinput38), .A(n10545), .ZN(n10552) );
  AOI22_X1 U11589 ( .A1(n10549), .A2(keyinput79), .B1(n10548), .B2(keyinput59), 
        .ZN(n10547) );
  OAI221_X1 U11590 ( .B1(n10549), .B2(keyinput79), .C1(n10548), .C2(keyinput59), .A(n10547), .ZN(n10551) );
  XNOR2_X1 U11591 ( .A(n5213), .B(keyinput11), .ZN(n10550) );
  OR3_X1 U11592 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n10557) );
  AOI22_X1 U11593 ( .A1(n8344), .A2(keyinput83), .B1(keyinput53), .B2(n7234), 
        .ZN(n10553) );
  OAI221_X1 U11594 ( .B1(n8344), .B2(keyinput83), .C1(n7234), .C2(keyinput53), 
        .A(n10553), .ZN(n10556) );
  XNOR2_X1 U11595 ( .A(n10554), .B(keyinput109), .ZN(n10555) );
  NOR3_X1 U11596 ( .A1(n10557), .A2(n10556), .A3(n10555), .ZN(n10558) );
  NAND4_X1 U11597 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n10620) );
  AOI22_X1 U11598 ( .A1(n10564), .A2(keyinput0), .B1(keyinput110), .B2(n10563), 
        .ZN(n10562) );
  OAI221_X1 U11599 ( .B1(n10564), .B2(keyinput0), .C1(n10563), .C2(keyinput110), .A(n10562), .ZN(n10573) );
  XNOR2_X1 U11600 ( .A(n10565), .B(keyinput89), .ZN(n10572) );
  XNOR2_X1 U11601 ( .A(keyinput18), .B(n9709), .ZN(n10571) );
  XNOR2_X1 U11602 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput96), .ZN(n10569)
         );
  XNOR2_X1 U11603 ( .A(SI_30_), .B(keyinput21), .ZN(n10568) );
  XNOR2_X1 U11604 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput88), .ZN(n10567) );
  XNOR2_X1 U11605 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput121), .ZN(n10566) );
  NAND4_X1 U11606 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  NOR4_X1 U11607 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10618) );
  XOR2_X1 U11608 ( .A(n10574), .B(keyinput34), .Z(n10579) );
  XOR2_X1 U11609 ( .A(n5926), .B(keyinput32), .Z(n10578) );
  XOR2_X1 U11610 ( .A(n10575), .B(keyinput106), .Z(n10577) );
  XNOR2_X1 U11611 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput4), .ZN(n10576) );
  NAND4_X1 U11612 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10586) );
  XOR2_X1 U11613 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput51), .Z(n10585) );
  INV_X1 U11614 ( .A(keyinput30), .ZN(n10581) );
  XNOR2_X1 U11615 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput127), .ZN(n10580)
         );
  OAI21_X1 U11616 ( .B1(P2_IR_REG_10__SCAN_IN), .B2(n10581), .A(n10580), .ZN(
        n10584) );
  XNOR2_X1 U11617 ( .A(n10582), .B(keyinput52), .ZN(n10583) );
  NOR4_X1 U11618 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10617) );
  AOI22_X1 U11619 ( .A1(n10588), .A2(keyinput10), .B1(keyinput42), .B2(n5817), 
        .ZN(n10587) );
  OAI221_X1 U11620 ( .B1(n10588), .B2(keyinput10), .C1(n5817), .C2(keyinput42), 
        .A(n10587), .ZN(n10600) );
  AOI22_X1 U11621 ( .A1(n6060), .A2(keyinput26), .B1(keyinput65), .B2(n10590), 
        .ZN(n10589) );
  OAI221_X1 U11622 ( .B1(n6060), .B2(keyinput26), .C1(n10590), .C2(keyinput65), 
        .A(n10589), .ZN(n10599) );
  AOI22_X1 U11623 ( .A1(n10593), .A2(keyinput119), .B1(keyinput82), .B2(n10592), .ZN(n10591) );
  OAI221_X1 U11624 ( .B1(n10593), .B2(keyinput119), .C1(n10592), .C2(
        keyinput82), .A(n10591), .ZN(n10598) );
  XOR2_X1 U11625 ( .A(n10594), .B(keyinput29), .Z(n10596) );
  XNOR2_X1 U11626 ( .A(SI_7_), .B(keyinput103), .ZN(n10595) );
  NAND2_X1 U11627 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  NOR4_X1 U11628 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .ZN(
        n10616) );
  INV_X1 U11629 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U11630 ( .A1(n10603), .A2(keyinput66), .B1(n10602), .B2(keyinput5), 
        .ZN(n10601) );
  OAI221_X1 U11631 ( .B1(n10603), .B2(keyinput66), .C1(n10602), .C2(keyinput5), 
        .A(n10601), .ZN(n10614) );
  AOI22_X1 U11632 ( .A1(n10605), .A2(keyinput22), .B1(n10356), .B2(keyinput23), 
        .ZN(n10604) );
  OAI221_X1 U11633 ( .B1(n10605), .B2(keyinput22), .C1(n10356), .C2(keyinput23), .A(n10604), .ZN(n10613) );
  AOI22_X1 U11634 ( .A1(n5786), .A2(keyinput40), .B1(n10607), .B2(keyinput81), 
        .ZN(n10606) );
  OAI221_X1 U11635 ( .B1(n5786), .B2(keyinput40), .C1(n10607), .C2(keyinput81), 
        .A(n10606), .ZN(n10612) );
  XOR2_X1 U11636 ( .A(n10608), .B(keyinput17), .Z(n10610) );
  XNOR2_X1 U11637 ( .A(SI_6_), .B(keyinput101), .ZN(n10609) );
  NAND2_X1 U11638 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NOR4_X1 U11639 ( .A1(n10614), .A2(n10613), .A3(n10612), .A4(n10611), .ZN(
        n10615) );
  NAND4_X1 U11640 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10619) );
  NOR4_X1 U11641 ( .A1(n10622), .A2(n10621), .A3(n10620), .A4(n10619), .ZN(
        n10623) );
  OAI21_X1 U11642 ( .B1(keyinput30), .B2(n10624), .A(n10623), .ZN(n10627) );
  XNOR2_X1 U11643 ( .A(n10625), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10626) );
  XNOR2_X1 U11644 ( .A(n10627), .B(n10626), .ZN(n10632) );
  NOR2_X1 U11645 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10628), .ZN(n10629) );
  NOR2_X1 U11646 ( .A1(n10630), .A2(n10629), .ZN(n10631) );
  XOR2_X1 U11647 ( .A(n10632), .B(n10631), .Z(ADD_1068_U4) );
  XOR2_X1 U11648 ( .A(n10634), .B(n10633), .Z(ADD_1068_U54) );
  NOR2_X1 U11649 ( .A1(n10636), .A2(n10635), .ZN(n10638) );
  XNOR2_X1 U11650 ( .A(n10638), .B(n10637), .ZN(ADD_1068_U50) );
  AOI21_X1 U11651 ( .B1(n10640), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10639), .ZN(
        n10642) );
  XNOR2_X1 U11652 ( .A(n10642), .B(n10641), .ZN(ADD_1068_U51) );
  XOR2_X1 U11653 ( .A(n10644), .B(n10643), .Z(ADD_1068_U53) );
  XNOR2_X1 U11654 ( .A(n10646), .B(n10645), .ZN(ADD_1068_U52) );
  INV_X2 U4948 ( .A(n9053), .ZN(n6984) );
  CLKBUF_X1 U4999 ( .A(n5154), .Z(n5155) );
  CLKBUF_X1 U5183 ( .A(n6063), .Z(n4553) );
  CLKBUF_X1 U5219 ( .A(n6073), .Z(n6659) );
  CLKBUF_X1 U5676 ( .A(n7788), .Z(n4416) );
endmodule

