

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984;

  INV_X2 U2302 ( .A(n3542), .ZN(n3347) );
  INV_X4 U2303 ( .A(n4770), .ZN(n4893) );
  AND2_X1 U2304 ( .A1(n2482), .A2(n2300), .ZN(n3607) );
  NAND2_X1 U2305 ( .A1(n2329), .A2(n2328), .ZN(n3220) );
  INV_X1 U2306 ( .A(n3556), .ZN(n3548) );
  INV_X1 U2307 ( .A(n3836), .ZN(n4665) );
  NAND2_X1 U2308 ( .A1(n2570), .A2(n2569), .ZN(n3669) );
  OAI21_X1 U2309 ( .B1(n4527), .B2(n2935), .A(n4528), .ZN(n4526) );
  OAI211_X1 U2310 ( .C1(IR_REG_1__SCAN_IN), .C2(IR_REG_31__SCAN_IN), .A(n2335), 
        .B(n2601), .ZN(n3841) );
  NAND4_X1 U2311 ( .A1(n2620), .A2(n2619), .A3(n2618), .A4(n2617), .ZN(n3835)
         );
  AOI21_X1 U2312 ( .B1(n4110), .B2(n4912), .A(n4115), .ZN(n2919) );
  NAND2_X1 U2313 ( .A1(n2555), .A2(n2563), .ZN(n2266) );
  INV_X2 U2314 ( .A(n2555), .ZN(n4483) );
  XNOR2_X2 U2315 ( .A(n2425), .B(IR_REG_2__SCAN_IN), .ZN(n4615) );
  INV_X1 U2316 ( .A(n2496), .ZN(n4143) );
  OAI21_X1 U2317 ( .B1(n4154), .B2(n2305), .A(n2497), .ZN(n2496) );
  OAI21_X1 U2318 ( .B1(n4121), .B2(n2873), .A(n3687), .ZN(n2874) );
  NAND2_X1 U2319 ( .A1(n2499), .A2(n2498), .ZN(n4154) );
  NAND2_X1 U2320 ( .A1(n2514), .A2(n2512), .ZN(n4201) );
  INV_X1 U2321 ( .A(n3018), .ZN(n3062) );
  OAI21_X1 U2322 ( .B1(n2294), .B2(n2774), .A(IR_REG_31__SCAN_IN), .ZN(n2834)
         );
  NAND2_X1 U2323 ( .A1(n2750), .A2(n2749), .ZN(n2774) );
  OAI21_X1 U2324 ( .B1(n2835), .B2(n2387), .A(IR_REG_31__SCAN_IN), .ZN(n2893)
         );
  INV_X8 U2325 ( .A(IR_REG_0__SCAN_IN), .ZN(n4609) );
  AND2_X1 U2326 ( .A1(n4134), .A2(n3686), .ZN(n4121) );
  AND2_X1 U2327 ( .A1(n4811), .A2(n2461), .ZN(n2457) );
  NAND2_X1 U2328 ( .A1(n4812), .A2(n4814), .ZN(n3462) );
  NAND2_X1 U2329 ( .A1(n3461), .A2(n3460), .ZN(n4811) );
  AND2_X1 U2330 ( .A1(n4390), .A2(n3748), .ZN(n4268) );
  NAND2_X1 U2331 ( .A1(n2396), .A2(n2394), .ZN(n2330) );
  AND2_X1 U2332 ( .A1(n4144), .A2(n4125), .ZN(n4127) );
  AND2_X1 U2333 ( .A1(n4152), .A2(n4146), .ZN(n4144) );
  NAND2_X1 U2334 ( .A1(n2724), .A2(n2723), .ZN(n4403) );
  NAND2_X1 U2335 ( .A1(n3613), .A2(n4160), .ZN(n2497) );
  NAND2_X1 U2336 ( .A1(n2664), .A2(n2663), .ZN(n3326) );
  OAI211_X1 U2337 ( .C1(n2452), .C2(n2450), .A(n2326), .B(n3219), .ZN(n3221)
         );
  NAND2_X1 U2338 ( .A1(n2329), .A2(n2455), .ZN(n2326) );
  OAI21_X1 U2339 ( .B1(n2453), .B2(n3160), .A(n3159), .ZN(n2452) );
  OR2_X1 U2340 ( .A1(n3145), .A2(n2454), .ZN(n2453) );
  AOI21_X1 U2341 ( .B1(n2508), .B2(n2506), .A(n2287), .ZN(n2505) );
  NAND2_X1 U2342 ( .A1(n2332), .A2(n3148), .ZN(n3149) );
  NOR2_X1 U2343 ( .A1(n2646), .A2(n2511), .ZN(n2510) );
  NAND2_X1 U2344 ( .A1(n4665), .A2(n3135), .ZN(n3720) );
  NAND4_X1 U2345 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n3836)
         );
  NAND4_X1 U2346 ( .A1(n2629), .A2(n2628), .A3(n2627), .A4(n2626), .ZN(n3834)
         );
  INV_X4 U2347 ( .A(n3555), .ZN(n3249) );
  AND2_X4 U2348 ( .A1(n4483), .A2(n3003), .ZN(n2610) );
  INV_X1 U2349 ( .A(n2563), .ZN(n3003) );
  XNOR2_X1 U2350 ( .A(n2550), .B(n3568), .ZN(n2555) );
  NAND2_X1 U2351 ( .A1(n2554), .A2(n2553), .ZN(n2563) );
  NAND2_X1 U2352 ( .A1(n2553), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U2353 ( .A(n2882), .B(n2545), .ZN(n2998) );
  XNOR2_X1 U2354 ( .A(n2889), .B(IR_REG_26__SCAN_IN), .ZN(n3008) );
  NAND2_X1 U2355 ( .A1(n2886), .A2(IR_REG_31__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U2356 ( .A1(n2734), .A2(IR_REG_31__SCAN_IN), .ZN(n2750) );
  AND3_X1 U2357 ( .A1(n2643), .A2(n2277), .A3(n2538), .ZN(n2544) );
  AND2_X1 U2358 ( .A1(n4609), .A2(n2621), .ZN(n2385) );
  AND2_X1 U2359 ( .A1(n2386), .A2(n2535), .ZN(n2384) );
  INV_X1 U2360 ( .A(IR_REG_1__SCAN_IN), .ZN(n2386) );
  NOR2_X1 U2361 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2534)
         );
  INV_X1 U2362 ( .A(IR_REG_5__SCAN_IN), .ZN(n2535) );
  NOR2_X1 U2363 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2682)
         );
  AND4_X2 U2364 ( .A1(n2599), .A2(n2600), .A3(n2597), .A4(n2598), .ZN(n2604)
         );
  INV_X1 U2365 ( .A(n2333), .ZN(n2267) );
  INV_X2 U2366 ( .A(n2333), .ZN(n3013) );
  NAND2_X1 U2367 ( .A1(n2570), .A2(n2569), .ZN(n2268) );
  NAND2_X1 U2368 ( .A1(n2570), .A2(n2569), .ZN(n2269) );
  OAI21_X2 U2369 ( .B1(n3291), .B2(n2413), .A(n2410), .ZN(n4307) );
  INV_X2 U2370 ( .A(n2266), .ZN(n2270) );
  INV_X2 U2371 ( .A(n2266), .ZN(n2271) );
  INV_X1 U2372 ( .A(IR_REG_13__SCAN_IN), .ZN(n2538) );
  AND2_X1 U2373 ( .A1(n2459), .A2(n2320), .ZN(n2379) );
  AND4_X1 U2374 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n2272)
         );
  NOR2_X1 U2375 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2542)
         );
  NOR2_X1 U2376 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2541)
         );
  NOR2_X1 U2377 ( .A1(n2395), .A2(n3434), .ZN(n2394) );
  INV_X1 U2378 ( .A(n3391), .ZN(n2395) );
  NAND2_X1 U2379 ( .A1(n2372), .A2(n3585), .ZN(n3461) );
  INV_X1 U2380 ( .A(n2510), .ZN(n2506) );
  INV_X1 U2381 ( .A(IR_REG_22__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U2382 ( .A1(n2751), .A2(n2539), .ZN(n2773) );
  INV_X1 U2383 ( .A(IR_REG_16__SCAN_IN), .ZN(n2539) );
  INV_X1 U2384 ( .A(IR_REG_9__SCAN_IN), .ZN(n2687) );
  NAND2_X1 U2385 ( .A1(n3009), .A2(n2397), .ZN(n3019) );
  AND2_X1 U2386 ( .A1(n4484), .A2(n3008), .ZN(n2397) );
  NAND2_X1 U2387 ( .A1(n2845), .A2(n2568), .ZN(n2569) );
  NAND2_X1 U2388 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2533) );
  INV_X1 U2389 ( .A(n2375), .ZN(n2374) );
  OAI21_X1 U2390 ( .B1(n2379), .B2(n2376), .A(n4933), .ZN(n2375) );
  INV_X1 U2391 ( .A(n2377), .ZN(n2376) );
  INV_X1 U2392 ( .A(n3669), .ZN(n3670) );
  OAI21_X1 U2393 ( .B1(n4622), .B2(n4617), .A(n2424), .ZN(n4620) );
  XNOR2_X1 U2394 ( .A(n2930), .B(n2428), .ZN(n4631) );
  INV_X1 U2395 ( .A(n2967), .ZN(n2341) );
  NOR2_X1 U2396 ( .A1(n4634), .A2(n2965), .ZN(n3051) );
  INV_X1 U2397 ( .A(n2544), .ZN(n2734) );
  NOR2_X1 U2398 ( .A1(n4081), .A2(n2951), .ZN(n4097) );
  INV_X1 U2399 ( .A(n4340), .ZN(n4339) );
  NAND2_X1 U2400 ( .A1(n2890), .A2(n3008), .ZN(n3006) );
  INV_X1 U2401 ( .A(n3039), .ZN(n3037) );
  NAND2_X1 U2402 ( .A1(n2883), .A2(n2417), .ZN(n2843) );
  NOR2_X1 U2403 ( .A1(n2502), .A2(IR_REG_25__SCAN_IN), .ZN(n2417) );
  INV_X1 U2404 ( .A(IR_REG_28__SCAN_IN), .ZN(n2503) );
  OR2_X1 U2405 ( .A1(n2774), .A2(n2483), .ZN(n2832) );
  INV_X1 U2406 ( .A(n2484), .ZN(n2483) );
  NAND2_X1 U2407 ( .A1(n4609), .A2(n2386), .ZN(n2601) );
  INV_X1 U2408 ( .A(n2495), .ZN(n2494) );
  OAI21_X1 U2409 ( .B1(n3289), .B2(n2317), .A(n2691), .ZN(n2495) );
  INV_X1 U2410 ( .A(n3147), .ZN(n2332) );
  NOR2_X1 U2411 ( .A1(n2351), .A2(n4582), .ZN(n2350) );
  INV_X1 U2412 ( .A(n2979), .ZN(n2351) );
  NOR2_X1 U2413 ( .A1(n4790), .A2(REG2_REG_13__SCAN_IN), .ZN(n2348) );
  AOI21_X1 U2414 ( .B1(n4571), .B2(n2350), .A(n2345), .ZN(n2981) );
  NAND2_X1 U2415 ( .A1(n2346), .A2(n4063), .ZN(n2345) );
  INV_X1 U2416 ( .A(n2348), .ZN(n2346) );
  OAI21_X1 U2417 ( .B1(n2518), .B2(n4215), .A(n2310), .ZN(n2516) );
  AND2_X1 U2418 ( .A1(n2525), .A2(n2519), .ZN(n2518) );
  NAND2_X1 U2419 ( .A1(n2522), .A2(n2520), .ZN(n2519) );
  NOR2_X1 U2420 ( .A1(n2521), .A2(n4215), .ZN(n2517) );
  INV_X1 U2421 ( .A(n2522), .ZN(n2521) );
  INV_X1 U2422 ( .A(n2516), .ZN(n2515) );
  OR2_X1 U2423 ( .A1(n2795), .A2(n2794), .ZN(n2796) );
  NOR2_X1 U2424 ( .A1(n4827), .A2(n2407), .ZN(n2406) );
  INV_X1 U2425 ( .A(n3673), .ZN(n2407) );
  AOI21_X1 U2426 ( .B1(n3737), .B2(n3738), .A(n2415), .ZN(n2414) );
  INV_X1 U2427 ( .A(n3708), .ZN(n2415) );
  OAI21_X1 U2428 ( .B1(n2491), .B2(n2490), .A(n2488), .ZN(n3186) );
  INV_X1 U2429 ( .A(n2489), .ZN(n2488) );
  OAI22_X1 U2430 ( .A1(n2490), .A2(n2615), .B1(n3103), .B2(n2852), .ZN(n2489)
         );
  NAND2_X1 U2431 ( .A1(n2286), .A2(n2616), .ZN(n2490) );
  INV_X1 U2432 ( .A(n3804), .ZN(n2615) );
  INV_X1 U2433 ( .A(n3115), .ZN(n2491) );
  INV_X1 U2434 ( .A(n2632), .ZN(n2511) );
  INV_X1 U2435 ( .A(n3240), .ZN(n2380) );
  OAI22_X1 U2436 ( .A1(n3220), .A2(n2382), .B1(n2383), .B2(n3218), .ZN(n2327)
         );
  INV_X1 U2437 ( .A(n2392), .ZN(n2391) );
  NAND2_X1 U2438 ( .A1(n3339), .A2(n3338), .ZN(n2477) );
  NAND2_X1 U2439 ( .A1(n2320), .A2(n2378), .ZN(n2377) );
  INV_X1 U2440 ( .A(n3649), .ZN(n2378) );
  NAND2_X1 U2441 ( .A1(n3554), .A2(n3553), .ZN(n2473) );
  NOR2_X1 U2442 ( .A1(n2476), .A2(n3020), .ZN(n3065) );
  NOR2_X1 U2443 ( .A1(n3347), .A2(n3072), .ZN(n2476) );
  OAI21_X1 U2444 ( .B1(n3556), .B2(n3072), .A(n3023), .ZN(n3024) );
  NAND2_X1 U2445 ( .A1(n2331), .A2(n3509), .ZN(n4966) );
  NAND2_X1 U2446 ( .A1(n4953), .A2(n4951), .ZN(n2331) );
  XNOR2_X1 U2447 ( .A(n3063), .B(n3557), .ZN(n3084) );
  NAND2_X1 U2448 ( .A1(n3837), .A2(n3542), .ZN(n3060) );
  XNOR2_X1 U2449 ( .A(n3080), .B(n3545), .ZN(n3097) );
  AOI21_X1 U2450 ( .B1(n2461), .B2(n2460), .A(n2313), .ZN(n2459) );
  INV_X1 U2451 ( .A(n4845), .ZN(n2460) );
  NAND2_X1 U2452 ( .A1(n2457), .A2(n3462), .ZN(n2458) );
  OR2_X1 U2453 ( .A1(n3071), .A2(n3070), .ZN(n3612) );
  AND4_X1 U2454 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n2564), .ZN(n4120)
         );
  NAND2_X1 U2455 ( .A1(n4610), .A2(n2449), .ZN(n2448) );
  NAND2_X1 U2456 ( .A1(n4615), .A2(REG2_REG_2__SCAN_IN), .ZN(n2449) );
  NOR2_X1 U2457 ( .A1(n4635), .A2(n4636), .ZN(n4634) );
  NAND2_X1 U2458 ( .A1(n4504), .A2(n2929), .ZN(n2930) );
  OAI21_X1 U2459 ( .B1(n2343), .B2(n2339), .A(n2279), .ZN(n2338) );
  NOR2_X1 U2460 ( .A1(n4508), .A2(n2969), .ZN(n4521) );
  NAND2_X1 U2461 ( .A1(n2932), .A2(n3053), .ZN(n2933) );
  XNOR2_X1 U2462 ( .A(n4526), .B(n4748), .ZN(n4533) );
  NOR2_X1 U2463 ( .A1(n4533), .A2(n4534), .ZN(n4532) );
  NAND2_X1 U2464 ( .A1(n2446), .A2(n2445), .ZN(n2970) );
  OR2_X1 U2465 ( .A1(n4525), .A2(REG2_REG_7__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U2466 ( .A1(n4521), .A2(n2447), .ZN(n2446) );
  NAND2_X1 U2467 ( .A1(n4525), .A2(REG2_REG_7__SCAN_IN), .ZN(n2447) );
  XNOR2_X1 U2468 ( .A(n2974), .B(n4759), .ZN(n4050) );
  NAND2_X1 U2469 ( .A1(n2434), .A2(n2433), .ZN(n2937) );
  NAND2_X1 U2470 ( .A1(n2435), .A2(REG1_REG_9__SCAN_IN), .ZN(n2433) );
  OAI21_X1 U2471 ( .B1(n2435), .B2(REG1_REG_9__SCAN_IN), .A(n4543), .ZN(n2434)
         );
  OAI21_X1 U2472 ( .B1(n4556), .B2(n2319), .A(n2941), .ZN(n2942) );
  NOR2_X1 U2473 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2537)
         );
  NAND2_X1 U2474 ( .A1(n2437), .A2(n2436), .ZN(n4069) );
  INV_X1 U2475 ( .A(n4071), .ZN(n2436) );
  NAND2_X1 U2476 ( .A1(n4065), .A2(n2946), .ZN(n4074) );
  AND2_X1 U2477 ( .A1(n4069), .A2(n2983), .ZN(n2985) );
  NAND2_X1 U2478 ( .A1(n3375), .A2(n3781), .ZN(n2487) );
  AND2_X1 U2479 ( .A1(n3271), .A2(n3726), .ZN(n3801) );
  AND2_X1 U2480 ( .A1(n3187), .A2(n3722), .ZN(n3803) );
  NOR2_X1 U2481 ( .A1(n4339), .A2(n2370), .ZN(n2369) );
  INV_X1 U2482 ( .A(n3689), .ZN(n2370) );
  NAND2_X1 U2483 ( .A1(n4127), .A2(n3689), .ZN(n4338) );
  INV_X1 U2484 ( .A(n3360), .ZN(n3376) );
  MUX2_X1 U2485 ( .A(IR_REG_31__SCAN_IN), .B(n2552), .S(IR_REG_29__SCAN_IN), 
        .Z(n2554) );
  INV_X1 U2486 ( .A(n2527), .ZN(n2387) );
  NAND2_X1 U2487 ( .A1(n2291), .A2(n2280), .ZN(n2486) );
  INV_X1 U2488 ( .A(IR_REG_15__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U2489 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U2490 ( .A1(n2293), .A2(IR_REG_1__SCAN_IN), .ZN(n2335) );
  AND2_X1 U2491 ( .A1(n2467), .A2(n4974), .ZN(n2466) );
  OAI21_X1 U2492 ( .B1(n3561), .B2(n2469), .A(n2468), .ZN(n2467) );
  NOR2_X1 U2493 ( .A1(n2474), .A2(n2470), .ZN(n2469) );
  NAND2_X1 U2494 ( .A1(n3561), .A2(n2473), .ZN(n2468) );
  NAND2_X1 U2495 ( .A1(n2472), .A2(n2473), .ZN(n2471) );
  INV_X1 U2496 ( .A(n3561), .ZN(n2472) );
  OAI21_X1 U2497 ( .B1(n3538), .B2(n3605), .A(n3537), .ZN(n3539) );
  NAND2_X1 U2498 ( .A1(n4631), .A2(REG1_REG_4__SCAN_IN), .ZN(n4639) );
  XNOR2_X1 U2499 ( .A(n2970), .B(n2675), .ZN(n4539) );
  NAND2_X1 U2500 ( .A1(n4066), .A2(REG1_REG_14__SCAN_IN), .ZN(n4065) );
  NAND2_X1 U2501 ( .A1(n2443), .A2(n2442), .ZN(n2441) );
  NAND2_X1 U2502 ( .A1(n4099), .A2(REG2_REG_18__SCAN_IN), .ZN(n2442) );
  XNOR2_X1 U2503 ( .A(n2955), .B(n2954), .ZN(n2423) );
  NAND2_X1 U2504 ( .A1(n2956), .A2(n2323), .ZN(n2422) );
  NAND2_X1 U2505 ( .A1(n3123), .A2(n4882), .ZN(n4770) );
  INV_X1 U2506 ( .A(n2998), .ZN(n3009) );
  INV_X1 U2507 ( .A(n3436), .ZN(n2393) );
  INV_X1 U2508 ( .A(n2530), .ZN(n2520) );
  NOR2_X1 U2509 ( .A1(n2529), .A2(n2523), .ZN(n2522) );
  INV_X1 U2510 ( .A(n4212), .ZN(n2523) );
  INV_X1 U2511 ( .A(n2324), .ZN(n2383) );
  NOR2_X1 U2512 ( .A1(n2393), .A2(n2390), .ZN(n2389) );
  INV_X1 U2513 ( .A(n3385), .ZN(n2390) );
  OAI21_X1 U2514 ( .B1(n2394), .B2(n2393), .A(n3640), .ZN(n2392) );
  NOR2_X1 U2515 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2568)
         );
  INV_X1 U2516 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4018) );
  INV_X1 U2517 ( .A(n3471), .ZN(n2462) );
  OR2_X1 U2518 ( .A1(n4499), .A2(n2962), .ZN(n2334) );
  INV_X1 U2519 ( .A(n2448), .ZN(n2961) );
  INV_X1 U2520 ( .A(IR_REG_3__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U2521 ( .A1(n2416), .A2(n3751), .ZN(n2872) );
  NAND2_X1 U2522 ( .A1(n4268), .A2(n3747), .ZN(n2416) );
  NAND2_X1 U2523 ( .A1(n4406), .A2(n2409), .ZN(n2408) );
  AOI21_X1 U2524 ( .B1(n2494), .B2(n2317), .A(n2278), .ZN(n2493) );
  AND2_X1 U2525 ( .A1(n3718), .A2(n3824), .ZN(n2895) );
  INV_X1 U2526 ( .A(n4972), .ZN(n3513) );
  NAND2_X1 U2527 ( .A1(n2911), .A2(n4387), .ZN(n2364) );
  OR2_X1 U2528 ( .A1(n4854), .A2(n4855), .ZN(n4386) );
  NAND2_X1 U2529 ( .A1(n2365), .A2(n2861), .ZN(n4319) );
  NOR2_X1 U2530 ( .A1(n4416), .A2(n4423), .ZN(n2365) );
  INV_X1 U2531 ( .A(n4723), .ZN(n4725) );
  NAND2_X1 U2532 ( .A1(n2399), .A2(n2398), .ZN(n4724) );
  NAND2_X1 U2533 ( .A1(n2400), .A2(n3271), .ZN(n2399) );
  INV_X1 U2534 ( .A(n2401), .ZN(n2400) );
  INV_X1 U2535 ( .A(n3214), .ZN(n3103) );
  INV_X1 U2536 ( .A(IR_REG_27__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U2537 ( .A1(n2548), .A2(n2504), .ZN(n2501) );
  AND2_X1 U2538 ( .A1(n2838), .A2(n2528), .ZN(n2527) );
  INV_X1 U2539 ( .A(IR_REG_21__SCAN_IN), .ZN(n2528) );
  NOR2_X1 U2540 ( .A1(n2486), .A2(n2290), .ZN(n2484) );
  OR2_X1 U2541 ( .A1(n2708), .A2(IR_REG_10__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U2542 ( .A1(n2330), .A2(n2303), .ZN(n3444) );
  AND2_X1 U2543 ( .A1(n3670), .A2(DATAI_23_), .ZN(n3599) );
  XNOR2_X1 U2544 ( .A(n3102), .B(n3557), .ZN(n3147) );
  INV_X1 U2545 ( .A(n2473), .ZN(n2470) );
  NOR2_X1 U2546 ( .A1(n3577), .A2(n2475), .ZN(n2474) );
  INV_X1 U2547 ( .A(n3659), .ZN(n2475) );
  AND2_X1 U2548 ( .A1(n3570), .A2(n3248), .ZN(n3259) );
  INV_X1 U2549 ( .A(n2452), .ZN(n2329) );
  NAND2_X1 U2550 ( .A1(n2456), .A2(n3149), .ZN(n2455) );
  INV_X1 U2551 ( .A(n3160), .ZN(n2456) );
  AND2_X1 U2552 ( .A1(n3670), .A2(DATAI_24_), .ZN(n3633) );
  INV_X1 U2553 ( .A(n3149), .ZN(n2454) );
  NAND2_X1 U2554 ( .A1(n3259), .A2(n3260), .ZN(n3303) );
  NAND2_X1 U2555 ( .A1(n3065), .A2(n3021), .ZN(n3025) );
  NAND2_X1 U2556 ( .A1(n3024), .A2(n3025), .ZN(n3067) );
  NOR2_X1 U2557 ( .A1(n2798), .A2(n4018), .ZN(n2807) );
  INV_X1 U2558 ( .A(n2806), .ZN(n2812) );
  NAND2_X1 U2559 ( .A1(n2477), .A2(n2308), .ZN(n3366) );
  NOR2_X1 U2560 ( .A1(n3597), .A2(n2479), .ZN(n2478) );
  INV_X1 U2561 ( .A(n3523), .ZN(n2479) );
  NOR2_X1 U2562 ( .A1(n2301), .A2(n2481), .ZN(n2480) );
  NOR2_X1 U2563 ( .A1(n3606), .A2(n3630), .ZN(n2481) );
  NAND2_X1 U2564 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2426) );
  OAI21_X1 U2565 ( .B1(n4616), .B2(n4625), .A(n4620), .ZN(n2928) );
  XNOR2_X1 U2566 ( .A(n2334), .B(n2963), .ZN(n4635) );
  OR2_X1 U2567 ( .A1(n3051), .A2(n3050), .ZN(n3048) );
  INV_X1 U2568 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3310) );
  OR2_X1 U2569 ( .A1(n4532), .A2(n2936), .ZN(n2435) );
  NAND2_X1 U2570 ( .A1(n4549), .A2(n2972), .ZN(n2974) );
  AOI21_X1 U2571 ( .B1(n4579), .B2(n4576), .A(n2944), .ZN(n2945) );
  NAND2_X1 U2572 ( .A1(n2348), .A2(n2980), .ZN(n2347) );
  NAND2_X1 U2573 ( .A1(n2350), .A2(n2980), .ZN(n2349) );
  NAND2_X1 U2574 ( .A1(n4592), .A2(n2986), .ZN(n4083) );
  NAND2_X1 U2575 ( .A1(n4083), .A2(n4085), .ZN(n4084) );
  NAND2_X1 U2576 ( .A1(n4629), .A2(ADDR_REG_18__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2577 ( .A1(n4197), .A2(n4183), .ZN(n2498) );
  NAND2_X1 U2578 ( .A1(n4171), .A2(n2500), .ZN(n2499) );
  NAND2_X1 U2579 ( .A1(n4161), .A2(n4177), .ZN(n2500) );
  INV_X1 U2580 ( .A(n4151), .ZN(n4160) );
  INV_X1 U2581 ( .A(n2513), .ZN(n2512) );
  OAI21_X1 U2582 ( .B1(n2516), .B2(n2517), .A(n2312), .ZN(n2513) );
  AND2_X1 U2583 ( .A1(n4219), .A2(n2871), .ZN(n4239) );
  AND2_X1 U2584 ( .A1(n2524), .A2(n2526), .ZN(n4258) );
  NAND2_X1 U2585 ( .A1(n2805), .A2(n2530), .ZN(n2524) );
  INV_X1 U2586 ( .A(n2872), .ZN(n4251) );
  AND2_X1 U2587 ( .A1(n3800), .A2(n3799), .ZN(n4292) );
  INV_X1 U2588 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3652) );
  NOR2_X1 U2589 ( .A1(n2780), .A2(n3652), .ZN(n2787) );
  NAND2_X1 U2590 ( .A1(n2767), .A2(REG3_REG_17__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U2591 ( .A1(n2405), .A2(n3675), .ZN(n2404) );
  INV_X1 U2592 ( .A(n2406), .ZN(n2405) );
  NAND2_X1 U2593 ( .A1(n2557), .A2(REG3_REG_15__SCAN_IN), .ZN(n2757) );
  INV_X1 U2594 ( .A(n2743), .ZN(n2557) );
  NOR2_X1 U2595 ( .A1(n2757), .A2(n4590), .ZN(n2767) );
  INV_X1 U2596 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U2597 ( .A1(n2408), .A2(n3673), .ZN(n4826) );
  NAND2_X1 U2598 ( .A1(n4822), .A2(n4825), .ZN(n4854) );
  OR2_X1 U2599 ( .A1(n2736), .A2(n3907), .ZN(n2743) );
  INV_X1 U2600 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U2601 ( .A1(n2487), .A2(n2309), .ZN(n2724) );
  AND2_X1 U2602 ( .A1(n2701), .A2(n2556), .ZN(n2715) );
  AND2_X1 U2603 ( .A1(REG3_REG_10__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2556) );
  AOI21_X1 U2604 ( .B1(n2414), .B2(n2412), .A(n2411), .ZN(n2410) );
  INV_X1 U2605 ( .A(n2414), .ZN(n2413) );
  INV_X1 U2606 ( .A(n3738), .ZN(n2412) );
  NOR2_X1 U2607 ( .A1(n2676), .A2(n3310), .ZN(n2701) );
  INV_X1 U2608 ( .A(n2508), .ZN(n2507) );
  AND2_X1 U2609 ( .A1(n2292), .A2(n2645), .ZN(n2508) );
  NAND2_X1 U2610 ( .A1(n3019), .A2(n3007), .ZN(n3039) );
  NOR2_X1 U2611 ( .A1(n2647), .A2(n3232), .ZN(n2655) );
  NAND2_X1 U2612 ( .A1(n3117), .A2(n2616), .ZN(n3201) );
  NAND2_X1 U2613 ( .A1(n2491), .A2(n2615), .ZN(n3117) );
  NOR2_X1 U2614 ( .A1(n3006), .A2(D_REG_1__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U2615 ( .A1(n3044), .A2(n2895), .ZN(n4906) );
  INV_X1 U2616 ( .A(n4862), .ZN(n4902) );
  AND2_X1 U2617 ( .A1(n3670), .A2(DATAI_26_), .ZN(n4151) );
  NOR2_X1 U2618 ( .A1(n4185), .A2(n4151), .ZN(n4152) );
  OR2_X1 U2619 ( .A1(n4202), .A2(n4183), .ZN(n4185) );
  OR2_X1 U2620 ( .A1(n4211), .A2(n3633), .ZN(n4202) );
  INV_X1 U2621 ( .A(n3633), .ZN(n4203) );
  AND2_X1 U2622 ( .A1(n4259), .A2(n3513), .ZN(n4244) );
  NAND2_X1 U2623 ( .A1(n4244), .A2(n4222), .ZN(n4211) );
  INV_X1 U2624 ( .A(n3599), .ZN(n4222) );
  NOR2_X1 U2625 ( .A1(n2275), .A2(n4958), .ZN(n4259) );
  NOR2_X1 U2626 ( .A1(n4386), .A2(n2364), .ZN(n4897) );
  NOR2_X1 U2627 ( .A1(n4319), .A2(n3588), .ZN(n4822) );
  INV_X1 U2628 ( .A(n2365), .ZN(n4417) );
  NAND2_X1 U2629 ( .A1(n3410), .A2(n3376), .ZN(n4416) );
  AND2_X1 U2630 ( .A1(n4721), .A2(n2362), .ZN(n3410) );
  AND2_X1 U2631 ( .A1(n2273), .A2(n3412), .ZN(n2362) );
  NAND2_X1 U2632 ( .A1(n4721), .A2(n2299), .ZN(n3325) );
  AND2_X1 U2633 ( .A1(n3280), .A2(n3279), .ZN(n4721) );
  INV_X1 U2634 ( .A(n4898), .ZN(n4872) );
  NAND2_X1 U2635 ( .A1(n2633), .A2(n2510), .ZN(n2509) );
  OR2_X1 U2636 ( .A1(n3211), .A2(n3196), .ZN(n3194) );
  NOR2_X1 U2637 ( .A1(n3194), .A2(n3181), .ZN(n3280) );
  NAND2_X1 U2638 ( .A1(n3210), .A2(n3103), .ZN(n3211) );
  NOR2_X1 U2639 ( .A1(n4673), .A2(n3135), .ZN(n3210) );
  NAND2_X1 U2640 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2845) );
  AND2_X1 U2641 ( .A1(n2547), .A2(n2504), .ZN(n2367) );
  NAND2_X1 U2642 ( .A1(n2887), .A2(n2886), .ZN(n2892) );
  INV_X1 U2643 ( .A(n2883), .ZN(n2884) );
  XNOR2_X1 U2644 ( .A(n2839), .B(n2838), .ZN(n2875) );
  NAND2_X1 U2645 ( .A1(n2837), .A2(n2276), .ZN(n3812) );
  INV_X1 U2646 ( .A(n3019), .ZN(n3105) );
  NAND2_X1 U2647 ( .A1(n3445), .A2(n3444), .ZN(n3587) );
  INV_X1 U2648 ( .A(n2482), .ZN(n3595) );
  NAND2_X1 U2649 ( .A1(n4967), .A2(n3523), .ZN(n3596) );
  NAND2_X1 U2650 ( .A1(n2477), .A2(n3343), .ZN(n3368) );
  NAND2_X1 U2651 ( .A1(n2373), .A2(n2377), .ZN(n4932) );
  NAND2_X1 U2652 ( .A1(n2458), .A2(n2379), .ZN(n2373) );
  OAI21_X1 U2653 ( .B1(n2269), .B2(n2603), .A(n2602), .ZN(n4662) );
  AND2_X1 U2654 ( .A1(n3670), .A2(DATAI_21_), .ZN(n4958) );
  NAND2_X1 U2655 ( .A1(n2396), .A2(n3391), .ZN(n3435) );
  NAND2_X1 U2656 ( .A1(n2463), .A2(n3471), .ZN(n3622) );
  NAND2_X1 U2657 ( .A1(n4844), .A2(n4845), .ZN(n2463) );
  INV_X1 U2658 ( .A(n2451), .ZN(n3161) );
  AOI21_X1 U2659 ( .B1(n3146), .B2(n3145), .A(n2454), .ZN(n2451) );
  NAND2_X1 U2660 ( .A1(n3303), .A2(n3302), .ZN(n3339) );
  NAND2_X1 U2661 ( .A1(n2267), .A2(REG2_REG_1__SCAN_IN), .ZN(n2599) );
  AND2_X1 U2662 ( .A1(n3670), .A2(DATAI_20_), .ZN(n4945) );
  NAND2_X1 U2663 ( .A1(n4931), .A2(n3495), .ZN(n4953) );
  NAND2_X1 U2664 ( .A1(n2330), .A2(n3436), .ZN(n3642) );
  AND2_X1 U2665 ( .A1(n3670), .A2(DATAI_22_), .ZN(n4972) );
  INV_X1 U2666 ( .A(n4934), .ZN(n4964) );
  NAND2_X1 U2667 ( .A1(n2458), .A2(n2459), .ZN(n3651) );
  AND2_X1 U2668 ( .A1(n3392), .A2(n3043), .ZN(n3822) );
  NAND4_X1 U2669 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n4180)
         );
  NAND4_X1 U2670 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n4225)
         );
  NAND4_X1 U2671 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n4963)
         );
  NAND2_X1 U2672 ( .A1(n3013), .A2(REG2_REG_2__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U2673 ( .A1(n3013), .A2(REG2_REG_0__SCAN_IN), .ZN(n2607) );
  INV_X2 U2674 ( .A(U4043), .ZN(n3838) );
  XNOR2_X1 U2675 ( .A(n3841), .B(REG2_REG_1__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U2676 ( .A1(n3848), .A2(n3847), .ZN(n3846) );
  NAND2_X1 U2677 ( .A1(n4613), .A2(n4612), .ZN(n4610) );
  XNOR2_X1 U2678 ( .A(n2448), .B(n2960), .ZN(n4500) );
  NAND2_X1 U2679 ( .A1(n4639), .A2(n2931), .ZN(n3055) );
  OAI211_X1 U2680 ( .C1(n3051), .C2(n2281), .A(n2337), .B(n2336), .ZN(n4509)
         );
  INV_X1 U2681 ( .A(n2338), .ZN(n2337) );
  INV_X1 U2682 ( .A(n4521), .ZN(n4520) );
  NAND2_X1 U2683 ( .A1(n4513), .A2(n2934), .ZN(n4527) );
  INV_X1 U2684 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U2685 ( .A1(n4538), .A2(n2971), .ZN(n4550) );
  NAND2_X1 U2686 ( .A1(n4550), .A2(n4551), .ZN(n4549) );
  INV_X1 U2687 ( .A(n2435), .ZN(n4546) );
  NAND2_X1 U2688 ( .A1(n4047), .A2(n2938), .ZN(n4556) );
  XNOR2_X1 U2689 ( .A(n2942), .B(n4782), .ZN(n4567) );
  NOR2_X1 U2690 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U2691 ( .A1(n2735), .A2(n2734), .ZN(n4589) );
  NAND2_X1 U2692 ( .A1(n4571), .A2(n2979), .ZN(n4585) );
  XNOR2_X1 U2693 ( .A(n2945), .B(n2980), .ZN(n4066) );
  NAND2_X1 U2694 ( .A1(n4074), .A2(n2420), .ZN(n4077) );
  NOR2_X1 U2695 ( .A1(n2322), .A2(n2421), .ZN(n2420) );
  NOR2_X1 U2696 ( .A1(n4486), .A2(REG1_REG_15__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U2697 ( .A(n2985), .B(n2984), .ZN(n4593) );
  NAND2_X1 U2698 ( .A1(n4593), .A2(n4591), .ZN(n4592) );
  NOR2_X1 U2699 ( .A1(n4595), .A2(REG1_REG_16__SCAN_IN), .ZN(n4596) );
  INV_X1 U2700 ( .A(n3429), .ZN(n4629) );
  NAND2_X1 U2701 ( .A1(n2432), .A2(n2431), .ZN(n2430) );
  NAND2_X1 U2702 ( .A1(n2948), .A2(n2432), .ZN(n2429) );
  INV_X1 U2703 ( .A(n4082), .ZN(n2432) );
  NAND2_X1 U2704 ( .A1(n4094), .A2(n4095), .ZN(n2361) );
  NOR2_X1 U2705 ( .A1(n2356), .A2(n2355), .ZN(n2354) );
  NAND2_X1 U2706 ( .A1(n2358), .A2(n2357), .ZN(n2356) );
  NOR2_X1 U2707 ( .A1(n4643), .A2(n4103), .ZN(n2355) );
  INV_X1 U2708 ( .A(n4096), .ZN(n2357) );
  NOR2_X1 U2709 ( .A1(n4094), .A2(n4095), .ZN(n4093) );
  INV_X1 U2710 ( .A(n2990), .ZN(n2440) );
  AOI21_X1 U2711 ( .B1(n2419), .B2(n4909), .A(n2284), .ZN(n4347) );
  XNOR2_X1 U2712 ( .A(n4121), .B(n4122), .ZN(n2419) );
  AND2_X1 U2713 ( .A1(n4124), .A2(n4869), .ZN(n2418) );
  NAND2_X1 U2714 ( .A1(n2487), .A2(n2714), .ZN(n4420) );
  INV_X1 U2715 ( .A(n4882), .ZN(n4920) );
  AND2_X1 U2716 ( .A1(n4770), .A2(n3124), .ZN(n4776) );
  XNOR2_X1 U2717 ( .A(n2371), .B(n4107), .ZN(n4435) );
  INV_X1 U2718 ( .A(n2371), .ZN(n4337) );
  NAND2_X2 U2719 ( .A1(n3037), .A2(n3006), .ZN(n4491) );
  INV_X1 U2720 ( .A(IR_REG_29__SCAN_IN), .ZN(n2549) );
  INV_X1 U2721 ( .A(IR_REG_30__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U2722 ( .A1(n2893), .A2(n2546), .ZN(n2881) );
  INV_X1 U2723 ( .A(n3812), .ZN(n3718) );
  XNOR2_X1 U2724 ( .A(n2315), .B(n2786), .ZN(n4099) );
  NAND2_X1 U2725 ( .A1(n2485), .A2(n2291), .ZN(n2785) );
  INV_X1 U2726 ( .A(n2774), .ZN(n2485) );
  NOR2_X1 U2727 ( .A1(n2644), .A2(n2643), .ZN(n4487) );
  NAND2_X1 U2728 ( .A1(IR_REG_31__SCAN_IN), .A2(n2601), .ZN(n2425) );
  NAND2_X1 U2729 ( .A1(n2466), .A2(n2471), .ZN(n2465) );
  NAND2_X1 U2730 ( .A1(n3086), .A2(n3085), .ZN(n3089) );
  NAND2_X1 U2731 ( .A1(n2359), .A2(n2353), .ZN(U3258) );
  OR2_X1 U2732 ( .A1(n2360), .A2(n4093), .ZN(n2359) );
  AND2_X1 U2733 ( .A1(n4102), .A2(n2354), .ZN(n2353) );
  NAND2_X1 U2734 ( .A1(n2361), .A2(n4611), .ZN(n2360) );
  AOI21_X1 U2735 ( .B1(n2423), .B2(n4630), .A(n2422), .ZN(n2444) );
  XNOR2_X1 U2736 ( .A(n2441), .B(n2440), .ZN(n2439) );
  AND2_X1 U2737 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  OR2_X1 U2738 ( .A1(n4113), .A2(n4431), .ZN(n2917) );
  AND2_X1 U2739 ( .A1(n2299), .A2(n3307), .ZN(n2273) );
  AND2_X1 U2740 ( .A1(n2409), .A2(n3675), .ZN(n2274) );
  OR3_X1 U2741 ( .A1(n4386), .A2(n2364), .A3(n2307), .ZN(n2275) );
  INV_X1 U2742 ( .A(n2963), .ZN(n2428) );
  OR2_X1 U2743 ( .A1(n2835), .A2(IR_REG_21__SCAN_IN), .ZN(n2276) );
  AND4_X1 U2744 ( .A1(n2682), .A2(n2537), .A3(n2536), .A4(n2687), .ZN(n2277)
         );
  AND2_X1 U2745 ( .A1(n3830), .A2(n3311), .ZN(n2278) );
  INV_X1 U2746 ( .A(n3050), .ZN(n2343) );
  OR2_X1 U2747 ( .A1(n2967), .A2(n2342), .ZN(n2279) );
  NAND2_X1 U2748 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  OR2_X1 U2749 ( .A1(n3050), .A2(n2342), .ZN(n2281) );
  AND2_X1 U2750 ( .A1(n2466), .A2(n2311), .ZN(n2282) );
  AND2_X1 U2751 ( .A1(n2527), .A2(n2289), .ZN(n2283) );
  OR2_X1 U2752 ( .A1(n4123), .A2(n2418), .ZN(n2284) );
  NAND4_X1 U2753 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n4663)
         );
  OR2_X1 U2754 ( .A1(n2352), .A2(n2981), .ZN(n2285) );
  INV_X1 U2755 ( .A(IR_REG_4__SCAN_IN), .ZN(n4036) );
  OR2_X1 U2756 ( .A1(n3835), .A2(n3214), .ZN(n2286) );
  NAND2_X1 U2757 ( .A1(n3462), .A2(n4811), .ZN(n4844) );
  AND2_X1 U2758 ( .A1(n3832), .A2(n3273), .ZN(n2287) );
  INV_X1 U2759 ( .A(IR_REG_2__SCAN_IN), .ZN(n2621) );
  NOR2_X1 U2760 ( .A1(n4596), .A2(n2948), .ZN(n2288) );
  AND2_X1 U2761 ( .A1(n2546), .A2(n2545), .ZN(n2289) );
  AND2_X1 U2762 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2290)
         );
  NAND2_X1 U2763 ( .A1(n2773), .A2(IR_REG_31__SCAN_IN), .ZN(n2291) );
  INV_X1 U2764 ( .A(IR_REG_25__SCAN_IN), .ZN(n2547) );
  OR2_X1 U2765 ( .A1(n3832), .A2(n3273), .ZN(n2292) );
  AND2_X1 U2766 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2293)
         );
  NAND2_X1 U2767 ( .A1(n2484), .A2(n2540), .ZN(n2294) );
  AND2_X1 U2768 ( .A1(n2625), .A2(n2630), .ZN(n2960) );
  INV_X1 U2769 ( .A(n2960), .ZN(n2927) );
  AND2_X1 U2770 ( .A1(n3048), .A2(n2967), .ZN(n2295) );
  AND2_X1 U2771 ( .A1(n3271), .A2(n3706), .ZN(n2296) );
  INV_X1 U2772 ( .A(n2340), .ZN(n2339) );
  NOR2_X1 U2773 ( .A1(n2341), .A2(n2968), .ZN(n2340) );
  AND2_X1 U2774 ( .A1(n2272), .A2(n2283), .ZN(n2297) );
  AND2_X1 U2775 ( .A1(n2297), .A2(n2544), .ZN(n2883) );
  INV_X1 U2776 ( .A(IR_REG_26__SCAN_IN), .ZN(n2504) );
  NAND4_X1 U2777 ( .A1(n2581), .A2(n2580), .A3(n2579), .A4(n2578), .ZN(n4197)
         );
  OR2_X1 U2778 ( .A1(n4386), .A2(n4391), .ZN(n2298) );
  INV_X1 U2779 ( .A(n4929), .ZN(n4297) );
  INV_X1 U2780 ( .A(n2968), .ZN(n2342) );
  AND2_X1 U2781 ( .A1(n4725), .A2(n3328), .ZN(n2299) );
  INV_X1 U2782 ( .A(n3726), .ZN(n2402) );
  NAND2_X1 U2783 ( .A1(n3530), .A2(n3529), .ZN(n2300) );
  AND2_X1 U2784 ( .A1(n3605), .A2(n3604), .ZN(n2301) );
  INV_X1 U2785 ( .A(IR_REG_24__SCAN_IN), .ZN(n2545) );
  OR3_X1 U2786 ( .A1(n4386), .A2(n2364), .A3(n4929), .ZN(n2302) );
  AND2_X1 U2787 ( .A1(n3436), .A2(n3443), .ZN(n2303) );
  NOR2_X1 U2788 ( .A1(n4899), .A2(n2795), .ZN(n2304) );
  NAND2_X1 U2789 ( .A1(n2643), .A2(n2277), .ZN(n2732) );
  AND2_X1 U2790 ( .A1(n4180), .A2(n4151), .ZN(n2305) );
  AND2_X1 U2791 ( .A1(n2408), .A2(n2406), .ZN(n2306) );
  OR2_X1 U2792 ( .A1(n4929), .A2(n4945), .ZN(n2307) );
  AND2_X1 U2793 ( .A1(n3349), .A2(n3343), .ZN(n2308) );
  AND2_X1 U2794 ( .A1(n2532), .A2(n2714), .ZN(n2309) );
  OR2_X1 U2795 ( .A1(n4963), .A2(n3599), .ZN(n2310) );
  INV_X1 U2796 ( .A(IR_REG_23__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U2797 ( .A1(n3561), .A2(n2474), .ZN(n2311) );
  OR2_X1 U2798 ( .A1(n4195), .A2(n4222), .ZN(n2312) );
  AND2_X1 U2799 ( .A1(n3477), .A2(n3619), .ZN(n2313) );
  NOR2_X1 U2800 ( .A1(n3478), .A2(n2462), .ZN(n2461) );
  AND2_X1 U2801 ( .A1(n2480), .A2(n2300), .ZN(n2314) );
  INV_X1 U2802 ( .A(n2529), .ZN(n2526) );
  OR2_X1 U2803 ( .A1(n2774), .A2(n2486), .ZN(n2315) );
  AND2_X1 U2804 ( .A1(n4721), .A2(n4725), .ZN(n2316) );
  NAND2_X1 U2805 ( .A1(n2883), .A2(n2547), .ZN(n2886) );
  INV_X1 U2806 ( .A(n4405), .ZN(n2409) );
  NAND2_X1 U2807 ( .A1(n2509), .A2(n2645), .ZN(n3270) );
  AND2_X1 U2808 ( .A1(n4729), .A2(n3263), .ZN(n2317) );
  INV_X1 U2809 ( .A(n3707), .ZN(n2411) );
  NOR2_X1 U2810 ( .A1(n3161), .A2(n3160), .ZN(n2318) );
  AND2_X1 U2811 ( .A1(n4554), .A2(REG1_REG_11__SCAN_IN), .ZN(n2319) );
  NAND2_X1 U2812 ( .A1(n4721), .A2(n2273), .ZN(n2363) );
  NAND2_X1 U2813 ( .A1(n3487), .A2(n3486), .ZN(n2320) );
  OR2_X1 U2814 ( .A1(n2886), .A2(n2501), .ZN(n2321) );
  AND2_X1 U2815 ( .A1(n2841), .A2(n3718), .ZN(n3018) );
  AND2_X1 U2816 ( .A1(n4486), .A2(REG1_REG_15__SCAN_IN), .ZN(n2322) );
  OR2_X1 U2817 ( .A1(n4643), .A2(n4732), .ZN(n2323) );
  AND2_X1 U2818 ( .A1(n3700), .A2(n2876), .ZN(n4864) );
  INV_X1 U2819 ( .A(n4864), .ZN(n4909) );
  AND2_X1 U2820 ( .A1(n2764), .A2(n2763), .ZN(n2984) );
  NAND2_X1 U2821 ( .A1(n3069), .A2(n3068), .ZN(n3086) );
  INV_X1 U2822 ( .A(n4611), .ZN(n4633) );
  AND2_X1 U2823 ( .A1(n4495), .A2(n4600), .ZN(n4611) );
  INV_X1 U2824 ( .A(n4183), .ZN(n4177) );
  AND2_X1 U2825 ( .A1(n3670), .A2(DATAI_25_), .ZN(n4183) );
  NAND2_X1 U2826 ( .A1(n3227), .A2(n3228), .ZN(n2324) );
  NAND2_X1 U2827 ( .A1(n3451), .A2(n3452), .ZN(n2325) );
  INV_X1 U2828 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2431) );
  AOI21_X2 U2829 ( .B1(n2327), .B2(n3221), .A(n2380), .ZN(n3572) );
  OR2_X2 U2830 ( .A1(n2455), .A2(n3146), .ZN(n2328) );
  NAND2_X2 U2831 ( .A1(n4966), .A2(n3519), .ZN(n4967) );
  OR2_X2 U2832 ( .A1(n3461), .A2(n3460), .ZN(n4812) );
  NAND2_X2 U2833 ( .A1(n3366), .A2(n3354), .ZN(n3386) );
  NAND2_X1 U2834 ( .A1(n4483), .A2(n2563), .ZN(n2333) );
  INV_X1 U2835 ( .A(n2334), .ZN(n2964) );
  NOR2_X1 U2836 ( .A1(n4500), .A2(n4501), .ZN(n4499) );
  NAND2_X1 U2837 ( .A1(n3051), .A2(n2340), .ZN(n2336) );
  NOR2_X1 U2838 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  INV_X1 U2839 ( .A(n4571), .ZN(n2344) );
  OAI21_X1 U2840 ( .B1(n2349), .B2(n2344), .A(n2347), .ZN(n2352) );
  INV_X1 U2841 ( .A(n2363), .ZN(n3413) );
  NAND2_X1 U2842 ( .A1(n2883), .A2(n2367), .ZN(n2366) );
  NAND2_X1 U2843 ( .A1(n4144), .A2(n2368), .ZN(n2371) );
  AND2_X1 U2844 ( .A1(n2369), .A2(n4125), .ZN(n2368) );
  NAND3_X1 U2845 ( .A1(n3445), .A2(n3444), .A3(n2325), .ZN(n2372) );
  OAI21_X2 U2846 ( .B1(n2458), .B2(n2376), .A(n2374), .ZN(n4931) );
  NAND2_X1 U2847 ( .A1(n2381), .A2(n3221), .ZN(n3239) );
  OAI21_X1 U2848 ( .B1(n3220), .B2(n3219), .A(n3218), .ZN(n2381) );
  OR2_X1 U2849 ( .A1(n2383), .A2(n3219), .ZN(n2382) );
  NAND3_X1 U2850 ( .A1(n2385), .A2(n2384), .A3(n2534), .ZN(n2642) );
  AND2_X1 U2851 ( .A1(n2622), .A2(n2534), .ZN(n2640) );
  NOR2_X1 U2852 ( .A1(IR_REG_2__SCAN_IN), .A2(n2601), .ZN(n2622) );
  NAND2_X1 U2853 ( .A1(n3386), .A2(n3385), .ZN(n2396) );
  NAND2_X1 U2854 ( .A1(n2388), .A2(n2391), .ZN(n3442) );
  NAND2_X1 U2855 ( .A1(n3386), .A2(n2389), .ZN(n2388) );
  NAND2_X2 U2856 ( .A1(n3062), .A2(n3019), .ZN(n3555) );
  NAND2_X1 U2857 ( .A1(n4724), .A2(n3731), .ZN(n2856) );
  NAND2_X1 U2858 ( .A1(n3175), .A2(n2296), .ZN(n2398) );
  OAI21_X1 U2859 ( .B1(n3175), .B2(n2855), .A(n3706), .ZN(n3272) );
  AOI21_X1 U2860 ( .B1(n2855), .B2(n3706), .A(n2402), .ZN(n2401) );
  NAND2_X1 U2861 ( .A1(n4406), .A2(n2274), .ZN(n2403) );
  NAND2_X1 U2862 ( .A1(n2403), .A2(n2404), .ZN(n4866) );
  OAI21_X1 U2863 ( .B1(n3291), .B2(n3737), .A(n3738), .ZN(n3415) );
  INV_X1 U2864 ( .A(n2843), .ZN(n2551) );
  NAND2_X1 U2865 ( .A1(n2843), .A2(IR_REG_31__SCAN_IN), .ZN(n2552) );
  MUX2_X1 U2866 ( .A(REG1_REG_2__SCAN_IN), .B(n4616), .S(n4615), .Z(n2424) );
  NOR2_X2 U2867 ( .A1(n2427), .A2(n2426), .ZN(n4622) );
  MUX2_X1 U2868 ( .A(REG1_REG_1__SCAN_IN), .B(n3842), .S(n3841), .Z(n2427) );
  OAI21_X1 U2869 ( .B1(n4595), .B2(n2430), .A(n2429), .ZN(n4081) );
  AOI211_X2 U2870 ( .C1(n4104), .C2(n3827), .A(n2879), .B(n2878), .ZN(n2880)
         );
  AOI21_X2 U2871 ( .B1(n4155), .B2(n3701), .A(n3772), .ZN(n4135) );
  NAND2_X1 U2872 ( .A1(n3719), .A2(n3717), .ZN(n4668) );
  NAND2_X1 U2873 ( .A1(n2551), .A2(n2549), .ZN(n2553) );
  XNOR2_X1 U2874 ( .A(n2928), .B(n2927), .ZN(n4505) );
  INV_X1 U2875 ( .A(n2437), .ZN(n4072) );
  OR2_X1 U2876 ( .A1(n4059), .A2(n2981), .ZN(n2437) );
  NOR2_X1 U2877 ( .A1(n2285), .A2(n4060), .ZN(n4059) );
  NAND2_X1 U2878 ( .A1(n2444), .A2(n2438), .ZN(U3259) );
  NAND2_X1 U2879 ( .A1(n2439), .A2(n4611), .ZN(n2438) );
  INV_X1 U2880 ( .A(n4093), .ZN(n2443) );
  INV_X1 U2881 ( .A(n3146), .ZN(n2450) );
  NAND2_X1 U2882 ( .A1(n3551), .A2(n2282), .ZN(n2464) );
  OAI211_X1 U2883 ( .C1(n3551), .C2(n2465), .A(n3567), .B(n2464), .ZN(U3217)
         );
  NAND2_X1 U2884 ( .A1(n3551), .A2(n3659), .ZN(n3578) );
  INV_X2 U2885 ( .A(n3347), .ZN(n3392) );
  INV_X2 U2886 ( .A(n3556), .ZN(n3467) );
  NAND2_X1 U2887 ( .A1(n4967), .A2(n2478), .ZN(n2482) );
  NAND2_X1 U2888 ( .A1(n2482), .A2(n2314), .ZN(n3541) );
  NAND3_X1 U2889 ( .A1(n3086), .A2(n3085), .A3(n3087), .ZN(n3099) );
  NAND2_X1 U2890 ( .A1(n3326), .A2(n2494), .ZN(n2492) );
  NAND2_X1 U2891 ( .A1(n2492), .A2(n2493), .ZN(n3414) );
  NAND3_X1 U2892 ( .A1(n2548), .A2(n2504), .A3(n2503), .ZN(n2502) );
  OAI21_X2 U2893 ( .B1(n2633), .B2(n2507), .A(n2505), .ZN(n4733) );
  NAND2_X1 U2894 ( .A1(n2633), .A2(n2632), .ZN(n3174) );
  NAND2_X1 U2895 ( .A1(n2805), .A2(n2515), .ZN(n2514) );
  NOR2_X1 U2896 ( .A1(n4239), .A2(n4213), .ZN(n2525) );
  NAND2_X1 U2897 ( .A1(n2544), .A2(n2272), .ZN(n2835) );
  NAND2_X1 U2898 ( .A1(n2604), .A2(n4662), .ZN(n3719) );
  NAND2_X1 U2899 ( .A1(n4896), .A2(n2304), .ZN(n2797) );
  INV_X2 U2900 ( .A(n4913), .ZN(n4915) );
  OR2_X1 U2901 ( .A1(n2915), .A2(n3120), .ZN(n4913) );
  INV_X1 U2902 ( .A(IR_REG_31__SCAN_IN), .ZN(n2686) );
  AND2_X1 U2903 ( .A1(n2712), .A2(n2721), .ZN(n4554) );
  INV_X1 U2904 ( .A(n4554), .ZN(n2940) );
  AND2_X1 U2905 ( .A1(n4957), .A2(n4945), .ZN(n2529) );
  OR2_X1 U2906 ( .A1(n4957), .A2(n4945), .ZN(n2530) );
  OR2_X1 U2907 ( .A1(n3550), .A2(n3549), .ZN(n2531) );
  INV_X1 U2908 ( .A(DATAI_1_), .ZN(n2603) );
  INV_X2 U2909 ( .A(n4916), .ZN(n4919) );
  OR2_X1 U2910 ( .A1(n4313), .A2(n4423), .ZN(n2532) );
  INV_X1 U2911 ( .A(IR_REG_19__SCAN_IN), .ZN(n2540) );
  NOR2_X1 U2912 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2536)
         );
  INV_X1 U2913 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2939) );
  INV_X1 U2914 ( .A(n3090), .ZN(n3087) );
  AND2_X1 U2915 ( .A1(REG3_REG_22__SCAN_IN), .A2(n2812), .ZN(n2588) );
  NAND2_X1 U2916 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  INV_X1 U2917 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2725) );
  INV_X1 U2918 ( .A(n3273), .ZN(n3279) );
  INV_X1 U2919 ( .A(IR_REG_20__SCAN_IN), .ZN(n2833) );
  INV_X1 U2920 ( .A(n2592), .ZN(n2558) );
  NAND2_X1 U2921 ( .A1(n2588), .A2(REG3_REG_23__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U2922 ( .A1(n4048), .A2(REG1_REG_10__SCAN_IN), .ZN(n4047) );
  AND2_X1 U2923 ( .A1(n4112), .A2(n2821), .ZN(n4128) );
  AND2_X1 U2924 ( .A1(n4830), .A2(n4861), .ZN(n3744) );
  OR2_X1 U2925 ( .A1(n2726), .A2(n2725), .ZN(n2736) );
  AND2_X1 U2926 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2634) );
  INV_X1 U2927 ( .A(n4726), .ZN(n4903) );
  INV_X1 U2928 ( .A(n4901), .ZN(n2911) );
  AND2_X2 U2929 ( .A1(n3720), .A2(n3723), .ZN(n3804) );
  NOR2_X1 U2930 ( .A1(n2684), .A2(n2683), .ZN(n2688) );
  NAND2_X1 U2931 ( .A1(n3522), .A2(n3521), .ZN(n3523) );
  NAND2_X1 U2932 ( .A1(n2268), .A2(n4488), .ZN(n2602) );
  NAND2_X1 U2933 ( .A1(n2558), .A2(REG3_REG_24__SCAN_IN), .ZN(n2583) );
  OR2_X1 U2934 ( .A1(n3071), .A2(n3045), .ZN(n4934) );
  INV_X1 U2935 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3232) );
  AND2_X1 U2936 ( .A1(n4525), .A2(REG1_REG_7__SCAN_IN), .ZN(n2935) );
  INV_X1 U2937 ( .A(n4757), .ZN(n4543) );
  NOR2_X1 U2938 ( .A1(n2943), .A2(n4566), .ZN(n4579) );
  OR2_X1 U2939 ( .A1(n2820), .A2(n2819), .ZN(n4112) );
  AND2_X1 U2940 ( .A1(n2875), .A2(n3812), .ZN(n4644) );
  AND2_X1 U2941 ( .A1(n2867), .A2(n4290), .ZN(n4899) );
  INV_X1 U2942 ( .A(n3455), .ZN(n4825) );
  NAND2_X1 U2943 ( .A1(n2715), .A2(REG3_REG_12__SCAN_IN), .ZN(n2726) );
  OR2_X1 U2944 ( .A1(n2665), .A2(n4535), .ZN(n2676) );
  OR2_X1 U2945 ( .A1(n3044), .A2(n3030), .ZN(n4726) );
  NAND2_X1 U2946 ( .A1(n2840), .A2(n4732), .ZN(n4669) );
  AND2_X1 U2947 ( .A1(n2841), .A2(n4485), .ZN(n4651) );
  NAND2_X1 U2948 ( .A1(n2787), .A2(REG3_REG_19__SCAN_IN), .ZN(n2798) );
  INV_X1 U2949 ( .A(n4846), .ZN(n4974) );
  AND4_X1 U2950 ( .A1(n2825), .A2(n2824), .A3(n2823), .A4(n2822), .ZN(n4140)
         );
  NAND2_X1 U2951 ( .A1(n4505), .A2(REG1_REG_3__SCAN_IN), .ZN(n4504) );
  XNOR2_X1 U2952 ( .A(n2947), .B(n2984), .ZN(n4595) );
  AND2_X1 U2953 ( .A1(n4495), .A2(n4603), .ZN(n4630) );
  AND2_X1 U2954 ( .A1(n2820), .A2(n2562), .ZN(n4141) );
  NAND2_X1 U2955 ( .A1(n2841), .A2(n4644), .ZN(n4898) );
  INV_X1 U2956 ( .A(n4906), .ZN(n4869) );
  NOR2_X1 U2957 ( .A1(n3039), .A2(n3718), .ZN(n3040) );
  INV_X1 U2958 ( .A(n4887), .ZN(n4924) );
  INV_X1 U2959 ( .A(n4886), .ZN(n4981) );
  NAND2_X1 U2960 ( .A1(n4913), .A2(REG1_REG_29__SCAN_IN), .ZN(n2916) );
  OAI22_X1 U2961 ( .A1(n3006), .A2(D_REG_0__SCAN_IN), .B1(n3008), .B2(n3009), 
        .ZN(n3120) );
  INV_X1 U2962 ( .A(n3416), .ZN(n3412) );
  NAND2_X1 U2963 ( .A1(n4669), .A2(n4792), .ZN(n4912) );
  OAI211_X1 U2964 ( .C1(n3119), .C2(n3026), .A(n2909), .B(n2908), .ZN(n2915)
         );
  AND2_X1 U2965 ( .A1(n4651), .A2(n2875), .ZN(n4705) );
  INV_X1 U2966 ( .A(n2875), .ZN(n3824) );
  INV_X1 U2967 ( .A(n4589), .ZN(n4790) );
  AND2_X1 U2968 ( .A1(n2654), .A2(n2684), .ZN(n2968) );
  AND2_X1 U2969 ( .A1(n2894), .A2(STATE_REG_SCAN_IN), .ZN(n3007) );
  OR2_X1 U2970 ( .A1(n3071), .A2(n3031), .ZN(n4846) );
  INV_X1 U2971 ( .A(n4120), .ZN(n4163) );
  NAND4_X1 U2972 ( .A1(n2804), .A2(n2803), .A3(n2802), .A4(n2801), .ZN(n4957)
         );
  NAND2_X1 U2973 ( .A1(n4495), .A2(n3044), .ZN(n4643) );
  OR2_X1 U2974 ( .A1(n4130), .A2(n4898), .ZN(n4886) );
  NAND2_X1 U2975 ( .A1(n3040), .A2(n4705), .ZN(n4882) );
  NAND2_X1 U2976 ( .A1(n4915), .A2(n4872), .ZN(n4431) );
  AND2_X1 U2977 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  NAND2_X1 U2978 ( .A1(n4919), .A2(n4872), .ZN(n4482) );
  OR2_X1 U2979 ( .A1(n2915), .A2(n2910), .ZN(n4916) );
  AND2_X1 U2980 ( .A1(n2891), .A2(n2892), .ZN(n3026) );
  INV_X1 U2981 ( .A(n4732), .ZN(n4485) );
  OR2_X1 U2982 ( .A1(n2690), .A2(n2689), .ZN(n4757) );
  AND2_X1 U2983 ( .A1(n3105), .A2(n3007), .ZN(U4043) );
  OAI21_X1 U2984 ( .B1(n2919), .B2(n4913), .A(n2918), .ZN(U3547) );
  OAI21_X1 U2985 ( .B1(n2919), .B2(n4916), .A(n2914), .ZN(U3515) );
  INV_X1 U2986 ( .A(n2773), .ZN(n2543) );
  NAND2_X1 U2987 ( .A1(n2271), .A2(REG0_REG_27__SCAN_IN), .ZN(n2567) );
  AND2_X4 U2988 ( .A1(n2555), .A2(n3003), .ZN(n2700) );
  NAND2_X1 U2989 ( .A1(n2700), .A2(REG1_REG_27__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U2990 ( .A1(n2634), .A2(REG3_REG_5__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U2991 ( .A1(n2655), .A2(REG3_REG_7__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U2992 ( .A1(n2807), .A2(REG3_REG_21__SCAN_IN), .ZN(n2806) );
  INV_X1 U2993 ( .A(n2583), .ZN(n2560) );
  AND2_X1 U2994 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2559) );
  NAND2_X1 U2995 ( .A1(n2560), .A2(n2559), .ZN(n2573) );
  INV_X1 U2996 ( .A(n2573), .ZN(n2561) );
  NAND2_X1 U2997 ( .A1(n2561), .A2(REG3_REG_27__SCAN_IN), .ZN(n2820) );
  INV_X1 U2998 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U2999 ( .A1(n2573), .A2(n4008), .ZN(n2562) );
  NAND2_X1 U3000 ( .A1(n2610), .A2(n4141), .ZN(n2565) );
  NAND2_X1 U3001 ( .A1(n3013), .A2(REG2_REG_27__SCAN_IN), .ZN(n2564) );
  OR2_X1 U3002 ( .A1(n2845), .A2(n2533), .ZN(n2570) );
  NAND2_X1 U3003 ( .A1(n3670), .A2(DATAI_27_), .ZN(n4146) );
  INV_X1 U3004 ( .A(n4146), .ZN(n4137) );
  NAND2_X1 U3005 ( .A1(n2700), .A2(REG1_REG_26__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U3006 ( .A1(n2270), .A2(REG0_REG_26__SCAN_IN), .ZN(n2576) );
  INV_X1 U3007 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3946) );
  INV_X1 U3008 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2571) );
  OAI21_X1 U3009 ( .B1(n2583), .B2(n3946), .A(n2571), .ZN(n2572) );
  AND2_X1 U3010 ( .A1(n2573), .A2(n2572), .ZN(n3662) );
  NAND2_X1 U3011 ( .A1(n2610), .A2(n3662), .ZN(n2575) );
  NAND2_X1 U3012 ( .A1(n3013), .A2(REG2_REG_26__SCAN_IN), .ZN(n2574) );
  INV_X1 U3013 ( .A(n4180), .ZN(n3613) );
  NAND2_X1 U3014 ( .A1(n2270), .A2(REG0_REG_25__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U3015 ( .A1(n2700), .A2(REG1_REG_25__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U3016 ( .A(n2583), .B(REG3_REG_25__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U3017 ( .A1(n2610), .A2(n4186), .ZN(n2579) );
  NAND2_X1 U3018 ( .A1(n3013), .A2(REG2_REG_25__SCAN_IN), .ZN(n2578) );
  INV_X1 U3019 ( .A(n4197), .ZN(n4161) );
  NAND2_X1 U3020 ( .A1(n2700), .A2(REG1_REG_24__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U3021 ( .A1(n2271), .A2(REG0_REG_24__SCAN_IN), .ZN(n2586) );
  INV_X1 U3022 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U3023 ( .A1(n2592), .A2(n3952), .ZN(n2582) );
  AND2_X1 U3024 ( .A1(n2583), .A2(n2582), .ZN(n3632) );
  NAND2_X1 U3025 ( .A1(n2610), .A2(n3632), .ZN(n2585) );
  NAND2_X1 U3026 ( .A1(n3013), .A2(REG2_REG_24__SCAN_IN), .ZN(n2584) );
  INV_X1 U3027 ( .A(n4225), .ZN(n4178) );
  NAND2_X1 U3028 ( .A1(n2700), .A2(REG1_REG_23__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U3029 ( .A1(n2271), .A2(REG0_REG_23__SCAN_IN), .ZN(n2595) );
  INV_X1 U3030 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2590) );
  INV_X1 U3031 ( .A(n2588), .ZN(n2589) );
  NAND2_X1 U3032 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  AND2_X1 U3033 ( .A1(n2592), .A2(n2591), .ZN(n3598) );
  NAND2_X1 U3034 ( .A1(n2610), .A2(n3598), .ZN(n2594) );
  NAND2_X1 U3035 ( .A1(n2267), .A2(REG2_REG_23__SCAN_IN), .ZN(n2593) );
  INV_X1 U3036 ( .A(n4963), .ZN(n4195) );
  NAND2_X1 U3037 ( .A1(n2700), .A2(REG1_REG_1__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U3038 ( .A1(n2610), .A2(REG3_REG_1__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3039 ( .A1(n2270), .A2(REG0_REG_1__SCAN_IN), .ZN(n2597) );
  INV_X1 U3040 ( .A(n3841), .ZN(n4488) );
  INV_X2 U3041 ( .A(n2604), .ZN(n3837) );
  INV_X1 U3042 ( .A(n4662), .ZN(n4675) );
  NAND2_X1 U3043 ( .A1(n3837), .A2(n4675), .ZN(n3717) );
  NAND2_X1 U3044 ( .A1(n2700), .A2(REG1_REG_0__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U3045 ( .A1(n2610), .A2(REG3_REG_0__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U3046 ( .A1(n2271), .A2(REG0_REG_0__SCAN_IN), .ZN(n2605) );
  INV_X1 U3047 ( .A(DATAI_0_), .ZN(n4599) );
  MUX2_X1 U3048 ( .A(n4599), .B(n4609), .S(n2269), .Z(n4674) );
  INV_X1 U3049 ( .A(n4674), .ZN(n3022) );
  AND2_X1 U3050 ( .A1(n4663), .A2(n3022), .ZN(n4667) );
  NAND2_X1 U3051 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U3052 ( .A1(n3837), .A2(n4662), .ZN(n2609) );
  NAND2_X1 U3053 ( .A1(n4666), .A2(n2609), .ZN(n3115) );
  NAND2_X1 U3054 ( .A1(n2700), .A2(REG1_REG_2__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U3055 ( .A1(n2270), .A2(REG0_REG_2__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3056 ( .A1(n2610), .A2(REG3_REG_2__SCAN_IN), .ZN(n2612) );
  MUX2_X1 U3057 ( .A(DATAI_2_), .B(n4615), .S(n2269), .Z(n3135) );
  INV_X1 U3058 ( .A(n3135), .ZN(n3129) );
  NAND2_X1 U3059 ( .A1(n3836), .A2(n3129), .ZN(n3723) );
  NAND2_X1 U3060 ( .A1(n4665), .A2(n3129), .ZN(n2616) );
  NAND2_X1 U3061 ( .A1(n2271), .A2(REG0_REG_3__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U3062 ( .A1(n3013), .A2(REG2_REG_3__SCAN_IN), .ZN(n2619) );
  INV_X1 U3063 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U3064 ( .A1(n2610), .A2(n4696), .ZN(n2618) );
  NAND2_X1 U3065 ( .A1(n2700), .A2(REG1_REG_3__SCAN_IN), .ZN(n2617) );
  OR2_X1 U3066 ( .A1(n2622), .A2(n2686), .ZN(n2624) );
  INV_X1 U3067 ( .A(n2624), .ZN(n2623) );
  NAND2_X1 U3068 ( .A1(n2623), .A2(IR_REG_3__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3069 ( .A1(n2624), .A2(n4033), .ZN(n2630) );
  MUX2_X1 U3070 ( .A(DATAI_3_), .B(n2960), .S(n2269), .Z(n3214) );
  INV_X1 U3071 ( .A(n3835), .ZN(n2852) );
  NAND2_X1 U3072 ( .A1(n2271), .A2(REG0_REG_4__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3073 ( .A1(n3013), .A2(REG2_REG_4__SCAN_IN), .ZN(n2628) );
  INV_X1 U3074 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4016) );
  XNOR2_X1 U3075 ( .A(n4016), .B(REG3_REG_3__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U3076 ( .A1(n2610), .A2(n3193), .ZN(n2627) );
  NAND2_X1 U3077 ( .A1(n2700), .A2(REG1_REG_4__SCAN_IN), .ZN(n2626) );
  INV_X1 U3078 ( .A(n3834), .ZN(n3177) );
  NAND2_X1 U3079 ( .A1(n2630), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  XNOR2_X1 U3080 ( .A(n2631), .B(IR_REG_4__SCAN_IN), .ZN(n2963) );
  MUX2_X1 U3081 ( .A(DATAI_4_), .B(n2963), .S(n3669), .Z(n3196) );
  NAND2_X1 U3082 ( .A1(n3177), .A2(n3196), .ZN(n2853) );
  INV_X1 U3083 ( .A(n3196), .ZN(n3143) );
  NAND2_X1 U3084 ( .A1(n3834), .A2(n3143), .ZN(n3727) );
  NAND2_X1 U3085 ( .A1(n2853), .A2(n3727), .ZN(n3782) );
  NAND2_X1 U3086 ( .A1(n3186), .A2(n3782), .ZN(n2633) );
  NAND2_X1 U3087 ( .A1(n3834), .A2(n3196), .ZN(n2632) );
  NAND2_X1 U3088 ( .A1(n2700), .A2(REG1_REG_5__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U3089 ( .A1(n2271), .A2(REG0_REG_5__SCAN_IN), .ZN(n2638) );
  OAI21_X1 U3090 ( .B1(n2634), .B2(REG3_REG_5__SCAN_IN), .A(n2647), .ZN(n4327)
         );
  INV_X1 U3091 ( .A(n4327), .ZN(n2635) );
  NAND2_X1 U3092 ( .A1(n2610), .A2(n2635), .ZN(n2637) );
  NAND2_X1 U3093 ( .A1(n3013), .A2(REG2_REG_5__SCAN_IN), .ZN(n2636) );
  NAND4_X1 U3094 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n3833)
         );
  NOR2_X1 U3095 ( .A1(n2640), .A2(n2686), .ZN(n2641) );
  MUX2_X1 U3096 ( .A(n2686), .B(n2641), .S(IR_REG_5__SCAN_IN), .Z(n2644) );
  INV_X1 U3097 ( .A(n2642), .ZN(n2643) );
  MUX2_X1 U3098 ( .A(DATAI_5_), .B(n4487), .S(n3669), .Z(n3181) );
  AND2_X1 U3099 ( .A1(n3833), .A2(n3181), .ZN(n2646) );
  INV_X1 U3100 ( .A(n3833), .ZN(n3275) );
  INV_X1 U3101 ( .A(n3181), .ZN(n3176) );
  NAND2_X1 U3102 ( .A1(n3275), .A2(n3176), .ZN(n2645) );
  NAND2_X1 U3103 ( .A1(n2270), .A2(REG0_REG_6__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3104 ( .A1(n3013), .A2(REG2_REG_6__SCAN_IN), .ZN(n2651) );
  AND2_X1 U3105 ( .A1(n2647), .A2(n3232), .ZN(n2648) );
  NOR2_X1 U3106 ( .A1(n2655), .A2(n2648), .ZN(n4711) );
  NAND2_X1 U3107 ( .A1(n2610), .A2(n4711), .ZN(n2650) );
  NAND2_X1 U3108 ( .A1(n2700), .A2(REG1_REG_6__SCAN_IN), .ZN(n2649) );
  NAND4_X1 U3109 ( .A1(n2652), .A2(n2651), .A3(n2650), .A4(n2649), .ZN(n3832)
         );
  NAND2_X1 U3110 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2653) );
  MUX2_X1 U3111 ( .A(IR_REG_31__SCAN_IN), .B(n2653), .S(IR_REG_6__SCAN_IN), 
        .Z(n2654) );
  OR2_X1 U3112 ( .A1(n2642), .A2(IR_REG_6__SCAN_IN), .ZN(n2684) );
  MUX2_X1 U3113 ( .A(DATAI_6_), .B(n2968), .S(n3669), .Z(n3273) );
  NAND2_X1 U3114 ( .A1(n2271), .A2(REG0_REG_7__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3115 ( .A1(n3013), .A2(REG2_REG_7__SCAN_IN), .ZN(n2660) );
  OR2_X1 U3116 ( .A1(n2655), .A2(REG3_REG_7__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3117 ( .A1(n2665), .A2(n2656), .ZN(n4740) );
  INV_X1 U3118 ( .A(n4740), .ZN(n2657) );
  NAND2_X1 U3119 ( .A1(n2610), .A2(n2657), .ZN(n2659) );
  NAND2_X1 U3120 ( .A1(n2700), .A2(REG1_REG_7__SCAN_IN), .ZN(n2658) );
  NAND4_X1 U3121 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n3831)
         );
  INV_X1 U3122 ( .A(n3831), .ZN(n2662) );
  NAND2_X1 U3123 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2671) );
  XNOR2_X1 U3124 ( .A(n2671), .B(IR_REG_7__SCAN_IN), .ZN(n4525) );
  MUX2_X1 U3125 ( .A(DATAI_7_), .B(n4525), .S(n3669), .Z(n4723) );
  NAND2_X1 U3126 ( .A1(n2662), .A2(n4723), .ZN(n3731) );
  NAND2_X1 U3127 ( .A1(n3831), .A2(n4725), .ZN(n3705) );
  NAND2_X1 U3128 ( .A1(n3731), .A2(n3705), .ZN(n4734) );
  NAND2_X1 U3129 ( .A1(n4733), .A2(n4734), .ZN(n2664) );
  NAND2_X1 U3130 ( .A1(n3831), .A2(n4723), .ZN(n2663) );
  NAND2_X1 U3131 ( .A1(n2271), .A2(REG0_REG_8__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3132 ( .A1(n3013), .A2(REG2_REG_8__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3133 ( .A1(n2665), .A2(n4535), .ZN(n2666) );
  AND2_X1 U3134 ( .A1(n2676), .A2(n2666), .ZN(n4749) );
  NAND2_X1 U3135 ( .A1(n2610), .A2(n4749), .ZN(n2668) );
  NAND2_X1 U3136 ( .A1(n2700), .A2(REG1_REG_8__SCAN_IN), .ZN(n2667) );
  NAND4_X1 U3137 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(n4729)
         );
  INV_X1 U3138 ( .A(n4729), .ZN(n2857) );
  INV_X1 U3139 ( .A(IR_REG_7__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U3140 ( .A1(n2671), .A2(n4038), .ZN(n2672) );
  NAND2_X1 U3141 ( .A1(n2672), .A2(IR_REG_31__SCAN_IN), .ZN(n2674) );
  INV_X1 U3142 ( .A(IR_REG_8__SCAN_IN), .ZN(n2673) );
  XNOR2_X1 U3143 ( .A(n2674), .B(n2673), .ZN(n4748) );
  INV_X1 U3144 ( .A(n4748), .ZN(n2675) );
  MUX2_X1 U3145 ( .A(DATAI_8_), .B(n2675), .S(n3669), .Z(n3263) );
  INV_X1 U3146 ( .A(n3263), .ZN(n3328) );
  NAND2_X1 U3147 ( .A1(n2857), .A2(n3328), .ZN(n3289) );
  NAND2_X1 U31480 ( .A1(n2270), .A2(REG0_REG_9__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U31490 ( .A1(n3013), .A2(REG2_REG_9__SCAN_IN), .ZN(n2680) );
  AND2_X1 U3150 ( .A1(n2676), .A2(n3310), .ZN(n2677) );
  NOR2_X1 U3151 ( .A1(n2701), .A2(n2677), .ZN(n3309) );
  NAND2_X1 U3152 ( .A1(n2610), .A2(n3309), .ZN(n2679) );
  NAND2_X1 U3153 ( .A1(n2700), .A2(REG1_REG_9__SCAN_IN), .ZN(n2678) );
  NAND4_X1 U3154 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n3830)
         );
  INV_X1 U3155 ( .A(n3830), .ZN(n3418) );
  INV_X1 U3156 ( .A(n2682), .ZN(n2683) );
  NOR2_X1 U3157 ( .A1(n2688), .A2(n2686), .ZN(n2685) );
  MUX2_X1 U3158 ( .A(n2686), .B(n2685), .S(IR_REG_9__SCAN_IN), .Z(n2690) );
  NAND2_X1 U3159 ( .A1(n2688), .A2(n2687), .ZN(n2708) );
  INV_X1 U3160 ( .A(n2708), .ZN(n2689) );
  MUX2_X1 U3161 ( .A(DATAI_9_), .B(n4543), .S(n3669), .Z(n3311) );
  INV_X1 U3162 ( .A(n3311), .ZN(n3307) );
  NAND2_X1 U3163 ( .A1(n3418), .A2(n3307), .ZN(n2691) );
  NAND2_X1 U3164 ( .A1(n2700), .A2(REG1_REG_10__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3165 ( .A1(n2271), .A2(REG0_REG_10__SCAN_IN), .ZN(n2695) );
  INV_X1 U3166 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2692) );
  XNOR2_X1 U3167 ( .A(n2701), .B(n2692), .ZN(n4760) );
  NAND2_X1 U3168 ( .A1(n2610), .A2(n4760), .ZN(n2694) );
  NAND2_X1 U3169 ( .A1(n3013), .A2(REG2_REG_10__SCAN_IN), .ZN(n2693) );
  NAND4_X1 U3170 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n3829)
         );
  NAND2_X1 U3171 ( .A1(n2708), .A2(IR_REG_31__SCAN_IN), .ZN(n2697) );
  XNOR2_X1 U3172 ( .A(n2697), .B(IR_REG_10__SCAN_IN), .ZN(n2973) );
  MUX2_X1 U3173 ( .A(DATAI_10_), .B(n2973), .S(n3669), .Z(n3416) );
  AND2_X1 U3174 ( .A1(n3829), .A2(n3416), .ZN(n2699) );
  INV_X1 U3175 ( .A(n3829), .ZN(n3377) );
  NAND2_X1 U3176 ( .A1(n3377), .A2(n3412), .ZN(n2698) );
  OAI21_X1 U3177 ( .B1(n3414), .B2(n2699), .A(n2698), .ZN(n3375) );
  NAND2_X1 U3178 ( .A1(n2700), .A2(REG1_REG_11__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3179 ( .A1(n2271), .A2(REG0_REG_11__SCAN_IN), .ZN(n2706) );
  AOI21_X1 U3180 ( .B1(n2701), .B2(REG3_REG_10__SCAN_IN), .A(
        REG3_REG_11__SCAN_IN), .ZN(n2702) );
  OR2_X1 U3181 ( .A1(n2715), .A2(n2702), .ZN(n4772) );
  INV_X1 U3182 ( .A(n4772), .ZN(n2703) );
  NAND2_X1 U3183 ( .A1(n2610), .A2(n2703), .ZN(n2705) );
  NAND2_X1 U3184 ( .A1(n3013), .A2(REG2_REG_11__SCAN_IN), .ZN(n2704) );
  NAND4_X1 U3185 ( .A1(n2707), .A2(n2706), .A3(n2705), .A4(n2704), .ZN(n4424)
         );
  INV_X1 U3186 ( .A(n4424), .ZN(n2713) );
  NAND2_X1 U3187 ( .A1(n2709), .A2(IR_REG_31__SCAN_IN), .ZN(n2711) );
  INV_X1 U3188 ( .A(IR_REG_11__SCAN_IN), .ZN(n2710) );
  OR2_X1 U3189 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  NAND2_X1 U3190 ( .A1(n2711), .A2(n2710), .ZN(n2721) );
  MUX2_X1 U3191 ( .A(DATAI_11_), .B(n4554), .S(n3669), .Z(n3360) );
  NAND2_X1 U3192 ( .A1(n2713), .A2(n3360), .ZN(n4304) );
  NAND2_X1 U3193 ( .A1(n4424), .A2(n3376), .ZN(n4306) );
  NAND2_X1 U3194 ( .A1(n4304), .A2(n4306), .ZN(n3781) );
  NAND2_X1 U3195 ( .A1(n2713), .A2(n3376), .ZN(n2714) );
  NAND2_X1 U3196 ( .A1(n2270), .A2(REG0_REG_12__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3197 ( .A1(n3013), .A2(REG2_REG_12__SCAN_IN), .ZN(n2719) );
  OR2_X1 U3198 ( .A1(n2715), .A2(REG3_REG_12__SCAN_IN), .ZN(n2716) );
  AND2_X1 U3199 ( .A1(n2726), .A2(n2716), .ZN(n4783) );
  NAND2_X1 U3200 ( .A1(n2610), .A2(n4783), .ZN(n2718) );
  NAND2_X1 U3201 ( .A1(n2700), .A2(REG1_REG_12__SCAN_IN), .ZN(n2717) );
  NAND4_X1 U3202 ( .A1(n2720), .A2(n2719), .A3(n2718), .A4(n2717), .ZN(n4313)
         );
  NAND2_X1 U3203 ( .A1(n2721), .A2(IR_REG_31__SCAN_IN), .ZN(n2722) );
  XNOR2_X1 U3204 ( .A(n2722), .B(IR_REG_12__SCAN_IN), .ZN(n2977) );
  MUX2_X1 U3205 ( .A(DATAI_12_), .B(n2977), .S(n3669), .Z(n4423) );
  NAND2_X1 U3206 ( .A1(n4313), .A2(n4423), .ZN(n2723) );
  NAND2_X1 U3207 ( .A1(n2700), .A2(REG1_REG_13__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3208 ( .A1(n2270), .A2(REG0_REG_13__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3209 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  AND2_X1 U32100 ( .A1(n2736), .A2(n2727), .ZN(n3643) );
  NAND2_X1 U32110 ( .A1(n2610), .A2(n3643), .ZN(n2729) );
  NAND2_X1 U32120 ( .A1(n2267), .A2(REG2_REG_13__SCAN_IN), .ZN(n2728) );
  NAND4_X1 U32130 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .ZN(n4407)
         );
  INV_X1 U32140 ( .A(n4407), .ZN(n4426) );
  NAND2_X1 U32150 ( .A1(n2732), .A2(IR_REG_31__SCAN_IN), .ZN(n2733) );
  MUX2_X1 U32160 ( .A(IR_REG_31__SCAN_IN), .B(n2733), .S(IR_REG_13__SCAN_IN), 
        .Z(n2735) );
  MUX2_X1 U32170 ( .A(DATAI_13_), .B(n4790), .S(n3669), .Z(n4320) );
  INV_X1 U32180 ( .A(n4320), .ZN(n2861) );
  NAND2_X1 U32190 ( .A1(n4426), .A2(n2861), .ZN(n4401) );
  NAND2_X1 U32200 ( .A1(n4403), .A2(n4401), .ZN(n2756) );
  NAND2_X1 U32210 ( .A1(n2271), .A2(REG0_REG_14__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U32220 ( .A1(n3013), .A2(REG2_REG_14__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U32230 ( .A1(n2736), .A2(n3907), .ZN(n2737) );
  AND2_X1 U32240 ( .A1(n2743), .A2(n2737), .ZN(n4800) );
  NAND2_X1 U32250 ( .A1(n2610), .A2(n4800), .ZN(n2739) );
  NAND2_X1 U32260 ( .A1(n2700), .A2(REG1_REG_14__SCAN_IN), .ZN(n2738) );
  NAND4_X1 U32270 ( .A1(n2741), .A2(n2740), .A3(n2739), .A4(n2738), .ZN(n4823)
         );
  INV_X1 U32280 ( .A(n4823), .ZN(n4315) );
  XNOR2_X1 U32290 ( .A(n2750), .B(IR_REG_14__SCAN_IN), .ZN(n4063) );
  MUX2_X1 U32300 ( .A(DATAI_14_), .B(n4063), .S(n3669), .Z(n3588) );
  NAND2_X1 U32310 ( .A1(n4315), .A2(n3588), .ZN(n3673) );
  INV_X1 U32320 ( .A(n3588), .ZN(n4410) );
  NAND2_X1 U32330 ( .A1(n4823), .A2(n4410), .ZN(n3674) );
  NAND2_X1 U32340 ( .A1(n3673), .A2(n3674), .ZN(n4405) );
  NAND2_X1 U32350 ( .A1(n2700), .A2(REG1_REG_15__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U32360 ( .A1(n2271), .A2(REG0_REG_15__SCAN_IN), .ZN(n2747) );
  INV_X1 U32370 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U32380 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  NAND2_X1 U32390 ( .A1(n2757), .A2(n2744), .ZN(n4818) );
  INV_X1 U32400 ( .A(n4818), .ZN(n4835) );
  NAND2_X1 U32410 ( .A1(n2610), .A2(n4835), .ZN(n2746) );
  NAND2_X1 U32420 ( .A1(n3013), .A2(REG2_REG_15__SCAN_IN), .ZN(n2745) );
  NAND4_X1 U32430 ( .A1(n2748), .A2(n2747), .A3(n2746), .A4(n2745), .ZN(n4859)
         );
  XNOR2_X1 U32440 ( .A(n2774), .B(n2751), .ZN(n4486) );
  MUX2_X1 U32450 ( .A(DATAI_15_), .B(n4486), .S(n3669), .Z(n3455) );
  NAND2_X1 U32460 ( .A1(n4859), .A2(n3455), .ZN(n2752) );
  NAND2_X1 U32470 ( .A1(n4407), .A2(n4320), .ZN(n4400) );
  AND3_X1 U32480 ( .A1(n4405), .A2(n2752), .A3(n4400), .ZN(n2755) );
  NAND2_X1 U32490 ( .A1(n4315), .A2(n4410), .ZN(n4819) );
  INV_X1 U32500 ( .A(n2752), .ZN(n2753) );
  OAI22_X1 U32510 ( .A1(n4819), .A2(n2753), .B1(n3455), .B2(n4859), .ZN(n2754)
         );
  AOI21_X2 U32520 ( .B1(n2756), .B2(n2755), .A(n2754), .ZN(n4857) );
  NAND2_X1 U32530 ( .A1(n2700), .A2(REG1_REG_16__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U32540 ( .A1(n2271), .A2(REG0_REG_16__SCAN_IN), .ZN(n2760) );
  AOI21_X1 U32550 ( .B1(n2757), .B2(n4590), .A(n2767), .ZN(n4875) );
  NAND2_X1 U32560 ( .A1(n2610), .A2(n4875), .ZN(n2759) );
  NAND2_X1 U32570 ( .A1(n3013), .A2(REG2_REG_16__SCAN_IN), .ZN(n2758) );
  NAND4_X1 U32580 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n4830)
         );
  OAI21_X1 U32590 ( .B1(n2774), .B2(IR_REG_15__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2762) );
  MUX2_X1 U32600 ( .A(IR_REG_31__SCAN_IN), .B(n2762), .S(IR_REG_16__SCAN_IN), 
        .Z(n2764) );
  OR2_X1 U32610 ( .A1(n2774), .A2(n2773), .ZN(n2763) );
  MUX2_X1 U32620 ( .A(DATAI_16_), .B(n2984), .S(n3669), .Z(n4855) );
  INV_X1 U32630 ( .A(n4855), .ZN(n4861) );
  INV_X1 U32640 ( .A(n3744), .ZN(n2765) );
  INV_X1 U32650 ( .A(n4830), .ZN(n4807) );
  NAND2_X1 U32660 ( .A1(n4807), .A2(n4855), .ZN(n3702) );
  NAND2_X1 U32670 ( .A1(n2765), .A2(n3702), .ZN(n4865) );
  NAND2_X1 U32680 ( .A1(n4857), .A2(n4865), .ZN(n4856) );
  NAND2_X1 U32690 ( .A1(n4830), .A2(n4855), .ZN(n2766) );
  NAND2_X1 U32700 ( .A1(n4856), .A2(n2766), .ZN(n4388) );
  NAND2_X1 U32710 ( .A1(n2271), .A2(REG0_REG_17__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U32720 ( .A1(n3013), .A2(REG2_REG_17__SCAN_IN), .ZN(n2771) );
  OAI21_X1 U32730 ( .B1(n2767), .B2(REG3_REG_17__SCAN_IN), .A(n2780), .ZN(
        n4883) );
  INV_X1 U32740 ( .A(n4883), .ZN(n2768) );
  NAND2_X1 U32750 ( .A1(n2610), .A2(n2768), .ZN(n2770) );
  NAND2_X1 U32760 ( .A1(n2700), .A2(REG1_REG_17__SCAN_IN), .ZN(n2769) );
  NAND4_X1 U32770 ( .A1(n2772), .A2(n2771), .A3(n2770), .A4(n2769), .ZN(n4904)
         );
  INV_X1 U32780 ( .A(n4904), .ZN(n2776) );
  INV_X1 U32790 ( .A(IR_REG_17__SCAN_IN), .ZN(n2775) );
  XNOR2_X1 U32800 ( .A(n2785), .B(n2775), .ZN(n2994) );
  MUX2_X1 U32810 ( .A(DATAI_17_), .B(n2994), .S(n3669), .Z(n4391) );
  INV_X1 U32820 ( .A(n4391), .ZN(n4387) );
  NAND2_X1 U32830 ( .A1(n2776), .A2(n4387), .ZN(n2777) );
  NAND2_X1 U32840 ( .A1(n4388), .A2(n2777), .ZN(n2779) );
  NAND2_X1 U32850 ( .A1(n4904), .A2(n4391), .ZN(n2778) );
  NAND2_X1 U32860 ( .A1(n2779), .A2(n2778), .ZN(n4283) );
  INV_X1 U32870 ( .A(n4283), .ZN(n4896) );
  NAND2_X1 U32880 ( .A1(n2270), .A2(REG0_REG_18__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U32890 ( .A1(n2267), .A2(REG2_REG_18__SCAN_IN), .ZN(n2783) );
  AOI21_X1 U32900 ( .B1(n2780), .B2(n3652), .A(n2787), .ZN(n4921) );
  NAND2_X1 U32910 ( .A1(n2610), .A2(n4921), .ZN(n2782) );
  NAND2_X1 U32920 ( .A1(n2700), .A2(REG1_REG_18__SCAN_IN), .ZN(n2781) );
  NAND4_X1 U32930 ( .A1(n2784), .A2(n2783), .A3(n2782), .A4(n2781), .ZN(n4930)
         );
  INV_X1 U32940 ( .A(n4930), .ZN(n4393) );
  INV_X1 U32950 ( .A(IR_REG_18__SCAN_IN), .ZN(n2786) );
  MUX2_X1 U32960 ( .A(DATAI_18_), .B(n4099), .S(n3669), .Z(n4901) );
  NAND2_X1 U32970 ( .A1(n4393), .A2(n4901), .ZN(n2867) );
  NAND2_X1 U32980 ( .A1(n4930), .A2(n2911), .ZN(n4290) );
  NAND2_X1 U32990 ( .A1(n2700), .A2(REG1_REG_19__SCAN_IN), .ZN(n2792) );
  NAND2_X1 U33000 ( .A1(n2271), .A2(REG0_REG_19__SCAN_IN), .ZN(n2791) );
  OR2_X1 U33010 ( .A1(n2787), .A2(REG3_REG_19__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U33020 ( .A1(n2788), .A2(n2798), .ZN(n4941) );
  INV_X1 U33030 ( .A(n4941), .ZN(n4299) );
  NAND2_X1 U33040 ( .A1(n2610), .A2(n4299), .ZN(n2790) );
  NAND2_X1 U33050 ( .A1(n3013), .A2(REG2_REG_19__SCAN_IN), .ZN(n2789) );
  NAND4_X1 U33060 ( .A1(n2792), .A2(n2791), .A3(n2790), .A4(n2789), .ZN(n4943)
         );
  XNOR2_X2 U33070 ( .A(n2832), .B(IR_REG_19__SCAN_IN), .ZN(n4732) );
  MUX2_X1 U33080 ( .A(DATAI_19_), .B(n4485), .S(n3669), .Z(n4929) );
  AND2_X1 U33090 ( .A1(n4943), .A2(n4929), .ZN(n2795) );
  NAND2_X1 U33100 ( .A1(n4393), .A2(n2911), .ZN(n4284) );
  INV_X1 U33110 ( .A(n4943), .ZN(n4907) );
  NAND2_X1 U33120 ( .A1(n4907), .A2(n4297), .ZN(n2793) );
  AND2_X1 U33130 ( .A1(n4284), .A2(n2793), .ZN(n2794) );
  NAND2_X1 U33140 ( .A1(n2797), .A2(n2796), .ZN(n4266) );
  INV_X1 U33150 ( .A(n4266), .ZN(n2805) );
  NAND2_X1 U33160 ( .A1(n2270), .A2(REG0_REG_20__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U33170 ( .A1(n3013), .A2(REG2_REG_20__SCAN_IN), .ZN(n2803) );
  INV_X1 U33180 ( .A(n2798), .ZN(n2800) );
  INV_X1 U33190 ( .A(n2807), .ZN(n2799) );
  OAI21_X1 U33200 ( .B1(REG3_REG_20__SCAN_IN), .B2(n2800), .A(n2799), .ZN(
        n4948) );
  INV_X1 U33210 ( .A(n4948), .ZN(n4278) );
  NAND2_X1 U33220 ( .A1(n2610), .A2(n4278), .ZN(n2802) );
  NAND2_X1 U33230 ( .A1(n2700), .A2(REG1_REG_20__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U33240 ( .A1(n2271), .A2(REG0_REG_21__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U33250 ( .A1(n3013), .A2(REG2_REG_21__SCAN_IN), .ZN(n2810) );
  OAI21_X1 U33260 ( .B1(REG3_REG_21__SCAN_IN), .B2(n2807), .A(n2806), .ZN(
        n4962) );
  INV_X1 U33270 ( .A(n4962), .ZN(n4260) );
  NAND2_X1 U33280 ( .A1(n2610), .A2(n4260), .ZN(n2809) );
  NAND2_X1 U33290 ( .A1(n2700), .A2(REG1_REG_21__SCAN_IN), .ZN(n2808) );
  NAND4_X1 U33300 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .ZN(n4971)
         );
  NAND2_X1 U33310 ( .A1(n4971), .A2(n4958), .ZN(n4212) );
  NAND2_X1 U33320 ( .A1(n2271), .A2(REG0_REG_22__SCAN_IN), .ZN(n2816) );
  NAND2_X1 U33330 ( .A1(n2700), .A2(REG1_REG_22__SCAN_IN), .ZN(n2815) );
  XNOR2_X1 U33340 ( .A(REG3_REG_22__SCAN_IN), .B(n2812), .ZN(n4978) );
  INV_X1 U33350 ( .A(n4978), .ZN(n4246) );
  NAND2_X1 U33360 ( .A1(n2610), .A2(n4246), .ZN(n2814) );
  NAND2_X1 U33370 ( .A1(n2267), .A2(REG2_REG_22__SCAN_IN), .ZN(n2813) );
  NAND4_X1 U33380 ( .A1(n2816), .A2(n2815), .A3(n2814), .A4(n2813), .ZN(n4949)
         );
  INV_X1 U33390 ( .A(n4949), .ZN(n4223) );
  NAND2_X1 U33400 ( .A1(n4223), .A2(n4972), .ZN(n4219) );
  NAND2_X1 U33410 ( .A1(n4949), .A2(n3513), .ZN(n2871) );
  NOR2_X1 U33420 ( .A1(n4971), .A2(n4958), .ZN(n4213) );
  NOR2_X1 U33430 ( .A1(n4223), .A2(n3513), .ZN(n4215) );
  AOI21_X1 U33440 ( .B1(n3633), .B2(n4225), .A(n4201), .ZN(n2817) );
  AOI21_X2 U33450 ( .B1(n4178), .B2(n4203), .A(n2817), .ZN(n4171) );
  OAI21_X1 U33460 ( .B1(n4137), .B2(n4163), .A(n4143), .ZN(n2818) );
  OAI21_X1 U33470 ( .B1(n4120), .B2(n4146), .A(n2818), .ZN(n4119) );
  NAND2_X1 U33480 ( .A1(n2700), .A2(REG1_REG_28__SCAN_IN), .ZN(n2825) );
  NAND2_X1 U33490 ( .A1(n2271), .A2(REG0_REG_28__SCAN_IN), .ZN(n2824) );
  INV_X1 U33500 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U33510 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  NAND2_X1 U33520 ( .A1(n2610), .A2(n4128), .ZN(n2823) );
  NAND2_X1 U3353 ( .A1(n2267), .A2(REG2_REG_28__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U33540 ( .A1(n3670), .A2(DATAI_28_), .ZN(n4125) );
  INV_X1 U3355 ( .A(n4125), .ZN(n3562) );
  OR2_X1 U3356 ( .A1(n4140), .A2(n3562), .ZN(n3691) );
  NAND2_X1 U3357 ( .A1(n4140), .A2(n3562), .ZN(n3687) );
  NAND2_X1 U3358 ( .A1(n3691), .A2(n3687), .ZN(n4122) );
  INV_X1 U3359 ( .A(n4140), .ZN(n3828) );
  AOI22_X1 U3360 ( .A1(n4119), .A2(n4122), .B1(n3562), .B2(n3828), .ZN(n2831)
         );
  NAND2_X1 U3361 ( .A1(n2700), .A2(REG1_REG_29__SCAN_IN), .ZN(n2830) );
  NAND2_X1 U3362 ( .A1(n2271), .A2(REG0_REG_29__SCAN_IN), .ZN(n2829) );
  INV_X1 U3363 ( .A(n4112), .ZN(n2826) );
  NAND2_X1 U3364 ( .A1(n2610), .A2(n2826), .ZN(n2828) );
  NAND2_X1 U3365 ( .A1(n2267), .A2(REG2_REG_29__SCAN_IN), .ZN(n2827) );
  NAND4_X1 U3366 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .ZN(n4124)
         );
  NAND2_X1 U3367 ( .A1(n3670), .A2(DATAI_29_), .ZN(n3689) );
  XNOR2_X1 U3368 ( .A(n4124), .B(n3689), .ZN(n3794) );
  XNOR2_X1 U3369 ( .A(n2831), .B(n3794), .ZN(n4110) );
  XNOR2_X1 U3370 ( .A(n2834), .B(n2833), .ZN(n2841) );
  NAND2_X1 U3371 ( .A1(n2835), .A2(IR_REG_31__SCAN_IN), .ZN(n2836) );
  MUX2_X1 U3372 ( .A(IR_REG_31__SCAN_IN), .B(n2836), .S(IR_REG_21__SCAN_IN), 
        .Z(n2837) );
  NAND2_X1 U3373 ( .A1(n2276), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  XNOR2_X1 U3374 ( .A(n3018), .B(n2875), .ZN(n2840) );
  INV_X1 U3375 ( .A(n4705), .ZN(n4792) );
  NAND2_X1 U3376 ( .A1(n2321), .A2(IR_REG_31__SCAN_IN), .ZN(n2842) );
  MUX2_X1 U3377 ( .A(IR_REG_31__SCAN_IN), .B(n2842), .S(IR_REG_28__SCAN_IN), 
        .Z(n2844) );
  NAND2_X1 U3378 ( .A1(n2844), .A2(n2843), .ZN(n3044) );
  XNOR2_X1 U3379 ( .A(n2845), .B(IR_REG_27__SCAN_IN), .ZN(n4494) );
  AND2_X1 U3380 ( .A1(n4494), .A2(B_REG_SCAN_IN), .ZN(n2846) );
  NOR2_X1 U3381 ( .A1(n4906), .A2(n2846), .ZN(n4104) );
  NAND2_X1 U3382 ( .A1(n2700), .A2(REG1_REG_30__SCAN_IN), .ZN(n2849) );
  NAND2_X1 U3383 ( .A1(n2267), .A2(REG2_REG_30__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U3384 ( .A1(n2271), .A2(REG0_REG_30__SCAN_IN), .ZN(n2847) );
  NAND3_X1 U3385 ( .A1(n2849), .A2(n2848), .A3(n2847), .ZN(n3827) );
  INV_X1 U3386 ( .A(n2895), .ZN(n3030) );
  INV_X1 U3387 ( .A(n2841), .ZN(n3813) );
  NAND2_X1 U3388 ( .A1(n3813), .A2(n4644), .ZN(n4862) );
  OAI22_X1 U3389 ( .A1(n4140), .A2(n4726), .B1(n3689), .B2(n4862), .ZN(n2879)
         );
  AND2_X1 U3390 ( .A1(n4225), .A2(n4203), .ZN(n4172) );
  NOR2_X1 U3391 ( .A1(n4161), .A2(n4183), .ZN(n2850) );
  NOR2_X1 U3392 ( .A1(n4172), .A2(n2850), .ZN(n3763) );
  NOR2_X1 U3393 ( .A1(n4225), .A2(n4203), .ZN(n3796) );
  NOR2_X1 U3394 ( .A1(n4963), .A2(n4222), .ZN(n4191) );
  NOR2_X1 U3395 ( .A1(n3796), .A2(n4191), .ZN(n3755) );
  INV_X1 U3396 ( .A(n4971), .ZN(n4241) );
  NAND2_X1 U3397 ( .A1(n4241), .A2(n4958), .ZN(n4217) );
  NAND2_X1 U3398 ( .A1(n4219), .A2(n4217), .ZN(n3753) );
  AND2_X1 U3399 ( .A1(n4904), .A2(n4387), .ZN(n4288) );
  NAND2_X1 U3400 ( .A1(n4943), .A2(n4297), .ZN(n3799) );
  NAND2_X1 U3401 ( .A1(n4290), .A2(n3799), .ZN(n2868) );
  NOR2_X1 U3402 ( .A1(n4288), .A2(n2868), .ZN(n3748) );
  INV_X1 U3403 ( .A(n4663), .ZN(n3072) );
  NAND2_X1 U3404 ( .A1(n3072), .A2(n3022), .ZN(n3798) );
  OR2_X1 U3405 ( .A1(n4668), .A2(n3798), .ZN(n4659) );
  NAND2_X1 U3406 ( .A1(n4659), .A2(n3719), .ZN(n2851) );
  NAND2_X1 U3407 ( .A1(n2851), .A2(n3804), .ZN(n3126) );
  NAND2_X1 U3408 ( .A1(n3126), .A2(n3720), .ZN(n3203) );
  NAND2_X1 U3409 ( .A1(n2852), .A2(n3214), .ZN(n3187) );
  NAND2_X1 U3410 ( .A1(n3835), .A2(n3103), .ZN(n3722) );
  NAND2_X1 U3411 ( .A1(n3203), .A2(n3803), .ZN(n3202) );
  AND2_X1 U3412 ( .A1(n3187), .A2(n2853), .ZN(n3729) );
  NAND2_X1 U3413 ( .A1(n3202), .A2(n3729), .ZN(n2854) );
  NAND2_X1 U3414 ( .A1(n2854), .A2(n3727), .ZN(n3175) );
  NAND2_X1 U3415 ( .A1(n3833), .A2(n3176), .ZN(n3725) );
  INV_X1 U3416 ( .A(n3725), .ZN(n2855) );
  NAND2_X1 U3417 ( .A1(n3275), .A2(n3181), .ZN(n3706) );
  NAND2_X1 U3418 ( .A1(n3832), .A2(n3279), .ZN(n3726) );
  INV_X1 U3419 ( .A(n3832), .ZN(n4727) );
  NAND2_X1 U3420 ( .A1(n4727), .A2(n3273), .ZN(n3271) );
  INV_X1 U3421 ( .A(n3271), .ZN(n3732) );
  NAND2_X1 U3422 ( .A1(n2856), .A2(n3705), .ZN(n3327) );
  NAND2_X1 U3423 ( .A1(n2857), .A2(n3263), .ZN(n3739) );
  NAND2_X1 U3424 ( .A1(n3327), .A2(n3739), .ZN(n2858) );
  NAND2_X1 U3425 ( .A1(n4729), .A2(n3328), .ZN(n3703) );
  NAND2_X1 U3426 ( .A1(n2858), .A2(n3703), .ZN(n3291) );
  NAND2_X1 U3427 ( .A1(n3830), .A2(n3307), .ZN(n3704) );
  INV_X1 U3428 ( .A(n3704), .ZN(n3737) );
  NAND2_X1 U3429 ( .A1(n3418), .A2(n3311), .ZN(n3738) );
  NAND2_X1 U3430 ( .A1(n3829), .A2(n3412), .ZN(n3708) );
  NAND2_X1 U3431 ( .A1(n3377), .A2(n3416), .ZN(n3707) );
  INV_X1 U3432 ( .A(n4423), .ZN(n4418) );
  NAND2_X1 U3433 ( .A1(n4313), .A2(n4418), .ZN(n4308) );
  NAND2_X1 U3434 ( .A1(n4407), .A2(n2861), .ZN(n2859) );
  AND2_X1 U3435 ( .A1(n4308), .A2(n2859), .ZN(n2863) );
  AND2_X1 U3436 ( .A1(n2863), .A2(n4306), .ZN(n3709) );
  NAND2_X1 U3437 ( .A1(n4307), .A2(n3709), .ZN(n2865) );
  INV_X1 U3438 ( .A(n4313), .ZN(n2860) );
  NAND2_X1 U3439 ( .A1(n2860), .A2(n4423), .ZN(n4310) );
  NAND2_X1 U3440 ( .A1(n4304), .A2(n4310), .ZN(n2864) );
  NOR2_X1 U3441 ( .A1(n4407), .A2(n2861), .ZN(n2862) );
  AOI21_X1 U3442 ( .B1(n2864), .B2(n2863), .A(n2862), .ZN(n3713) );
  NAND2_X1 U3443 ( .A1(n2865), .A2(n3713), .ZN(n4406) );
  INV_X1 U3444 ( .A(n4859), .ZN(n2866) );
  NAND2_X1 U3445 ( .A1(n2866), .A2(n3455), .ZN(n3677) );
  NAND2_X1 U3446 ( .A1(n4859), .A2(n4825), .ZN(n3675) );
  NAND2_X1 U3447 ( .A1(n3677), .A2(n3675), .ZN(n4827) );
  NOR2_X1 U3448 ( .A1(n4866), .A2(n4865), .ZN(n4863) );
  NOR2_X2 U3449 ( .A1(n4863), .A2(n3744), .ZN(n4390) );
  INV_X1 U3450 ( .A(n4945), .ZN(n3792) );
  NAND2_X1 U3451 ( .A1(n4957), .A2(n3792), .ZN(n3747) );
  NOR2_X1 U3452 ( .A1(n3792), .A2(n4957), .ZN(n2870) );
  INV_X1 U3453 ( .A(n2867), .ZN(n4291) );
  NOR2_X1 U3454 ( .A1(n4904), .A2(n4387), .ZN(n4286) );
  NOR2_X1 U3455 ( .A1(n4291), .A2(n4286), .ZN(n2869) );
  NAND2_X1 U3456 ( .A1(n4907), .A2(n4929), .ZN(n3800) );
  OAI21_X1 U3457 ( .B1(n2869), .B2(n2868), .A(n3800), .ZN(n4267) );
  OAI21_X1 U34580 ( .B1(n2870), .B2(n4267), .A(n3747), .ZN(n3751) );
  INV_X1 U34590 ( .A(n4958), .ZN(n4254) );
  AND2_X1 U3460 ( .A1(n4971), .A2(n4254), .ZN(n4218) );
  NAND2_X1 U3461 ( .A1(n4963), .A2(n4222), .ZN(n3789) );
  NAND2_X1 U3462 ( .A1(n3789), .A2(n2871), .ZN(n3756) );
  AOI21_X1 U3463 ( .B1(n4218), .B2(n4219), .A(n3756), .ZN(n3682) );
  OAI21_X1 U3464 ( .B1(n3753), .B2(n2872), .A(n3682), .ZN(n4193) );
  NAND2_X1 U3465 ( .A1(n3755), .A2(n4193), .ZN(n4174) );
  NAND2_X1 U3466 ( .A1(n3763), .A2(n4174), .ZN(n4155) );
  NOR2_X1 U34670 ( .A1(n4197), .A2(n4177), .ZN(n4157) );
  NOR2_X1 U3468 ( .A1(n4180), .A2(n4160), .ZN(n3771) );
  NOR2_X1 U34690 ( .A1(n4157), .A2(n3771), .ZN(n3701) );
  NAND2_X1 U3470 ( .A1(n4180), .A2(n4160), .ZN(n3694) );
  INV_X1 U34710 ( .A(n3694), .ZN(n3772) );
  XNOR2_X1 U3472 ( .A(n4120), .B(n4146), .ZN(n4142) );
  NAND2_X1 U34730 ( .A1(n4135), .A2(n4142), .ZN(n4134) );
  NAND2_X1 U3474 ( .A1(n4120), .A2(n4137), .ZN(n3686) );
  INV_X1 U34750 ( .A(n3691), .ZN(n2873) );
  XNOR2_X1 U3476 ( .A(n2874), .B(n3794), .ZN(n2877) );
  OR2_X1 U34770 ( .A1(n2841), .A2(n3812), .ZN(n3700) );
  OR2_X1 U3478 ( .A1(n4732), .A2(n2875), .ZN(n2876) );
  NOR2_X1 U34790 ( .A1(n2877), .A2(n4864), .ZN(n2878) );
  INV_X1 U3480 ( .A(n2880), .ZN(n4115) );
  NAND2_X1 U34810 ( .A1(n2881), .A2(IR_REG_31__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3482 ( .A1(n2884), .A2(IR_REG_31__SCAN_IN), .ZN(n2885) );
  MUX2_X1 U34830 ( .A(IR_REG_31__SCAN_IN), .B(n2885), .S(IR_REG_25__SCAN_IN), 
        .Z(n2887) );
  NAND2_X1 U3484 ( .A1(n2892), .A2(n2998), .ZN(n2888) );
  MUX2_X1 U34850 ( .A(n2998), .B(n2888), .S(B_REG_SCAN_IN), .Z(n2890) );
  INV_X1 U3486 ( .A(n3008), .ZN(n2891) );
  AND2_X1 U34870 ( .A1(n4705), .A2(n3812), .ZN(n2896) );
  INV_X1 U3488 ( .A(n2892), .ZN(n4484) );
  XNOR2_X1 U34890 ( .A(n2893), .B(IR_REG_23__SCAN_IN), .ZN(n2921) );
  INV_X1 U3490 ( .A(n2921), .ZN(n2894) );
  NAND2_X1 U34910 ( .A1(n2841), .A2(n4732), .ZN(n3029) );
  NAND2_X1 U3492 ( .A1(n3029), .A2(n2895), .ZN(n3033) );
  NAND2_X1 U34930 ( .A1(n3037), .A2(n3033), .ZN(n3118) );
  NOR2_X1 U3494 ( .A1(n2896), .A2(n3118), .ZN(n2909) );
  NOR4_X1 U34950 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2900) );
  NOR4_X1 U3496 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2899) );
  NOR4_X1 U34970 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2898) );
  NOR4_X1 U3498 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2897) );
  NAND4_X1 U34990 ( .A1(n2900), .A2(n2899), .A3(n2898), .A4(n2897), .ZN(n2906)
         );
  NOR2_X1 U3500 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2904)
         );
  NOR4_X1 U35010 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2903) );
  NOR4_X1 U3502 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U35030 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2901) );
  NAND4_X1 U3504 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .ZN(n2905)
         );
  NOR2_X1 U35050 ( .A1(n2906), .A2(n2905), .ZN(n2907) );
  NOR2_X1 U35060 ( .A1(n3006), .A2(n2907), .ZN(n3027) );
  INV_X1 U35070 ( .A(n3027), .ZN(n2908) );
  INV_X1 U35080 ( .A(n3120), .ZN(n2910) );
  NAND2_X1 U35090 ( .A1(n4675), .A2(n4674), .ZN(n4673) );
  OAI21_X1 U35100 ( .B1(n4127), .B2(n3689), .A(n4338), .ZN(n4113) );
  OR2_X1 U35110 ( .A1(n4113), .A2(n4482), .ZN(n2913) );
  NAND2_X1 U35120 ( .A1(n4916), .A2(REG0_REG_29__SCAN_IN), .ZN(n2912) );
  INV_X2 U35130 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U35140 ( .A1(n3030), .A2(n2921), .ZN(n2920) );
  NOR2_X1 U35150 ( .A1(n3669), .A2(n2920), .ZN(n2924) );
  NAND2_X1 U35160 ( .A1(n2921), .A2(STATE_REG_SCAN_IN), .ZN(n4489) );
  NAND2_X1 U35170 ( .A1(n3039), .A2(n4489), .ZN(n2922) );
  AND2_X1 U35180 ( .A1(n2924), .A2(n2922), .ZN(n4495) );
  INV_X1 U35190 ( .A(n2922), .ZN(n2923) );
  OR2_X1 U35200 ( .A1(n2924), .A2(n2923), .ZN(n3429) );
  AND2_X1 U35210 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4936) );
  AOI21_X1 U35220 ( .B1(n4629), .B2(ADDR_REG_19__SCAN_IN), .A(n4936), .ZN(
        n2956) );
  INV_X1 U35230 ( .A(n4099), .ZN(n4103) );
  INV_X1 U35240 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4914) );
  NOR2_X1 U35250 ( .A1(n2994), .A2(REG1_REG_17__SCAN_IN), .ZN(n2951) );
  INV_X1 U35260 ( .A(n4486), .ZN(n4080) );
  INV_X1 U35270 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U35280 ( .A1(n4487), .A2(REG1_REG_5__SCAN_IN), .ZN(n2932) );
  INV_X1 U35290 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2925) );
  MUX2_X1 U35300 ( .A(n2925), .B(REG1_REG_5__SCAN_IN), .S(n4487), .Z(n2926) );
  INV_X1 U35310 ( .A(n2926), .ZN(n3054) );
  INV_X1 U35320 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4616) );
  INV_X1 U35330 ( .A(n4615), .ZN(n4625) );
  INV_X1 U35340 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4648) );
  INV_X1 U35350 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3842) );
  NOR2_X1 U35360 ( .A1(n3841), .A2(n3842), .ZN(n4617) );
  NAND2_X1 U35370 ( .A1(n2960), .A2(n2928), .ZN(n2929) );
  NAND2_X1 U35380 ( .A1(n2963), .A2(n2930), .ZN(n2931) );
  NAND2_X1 U35390 ( .A1(n3054), .A2(n3055), .ZN(n3053) );
  XNOR2_X1 U35400 ( .A(n2933), .B(n2342), .ZN(n4514) );
  NAND2_X1 U35410 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4514), .ZN(n4513) );
  NAND2_X1 U35420 ( .A1(n2968), .A2(n2933), .ZN(n2934) );
  INV_X1 U35430 ( .A(n4525), .ZN(n4720) );
  INV_X1 U35440 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U35450 ( .A1(n4720), .A2(n4744), .ZN(n4528) );
  NOR2_X1 U35460 ( .A1(n4748), .A2(n4526), .ZN(n2936) );
  INV_X1 U35470 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4534) );
  INV_X1 U35480 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U35490 ( .A1(n2973), .A2(n2937), .ZN(n2938) );
  INV_X1 U35500 ( .A(n2973), .ZN(n4759) );
  XNOR2_X1 U35510 ( .A(n2937), .B(n4759), .ZN(n4048) );
  INV_X1 U35520 ( .A(n2977), .ZN(n4782) );
  NOR2_X1 U35530 ( .A1(n2942), .A2(n4782), .ZN(n2943) );
  INV_X1 U35540 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4568) );
  NAND2_X1 U35550 ( .A1(n4790), .A2(REG1_REG_13__SCAN_IN), .ZN(n4576) );
  INV_X1 U35560 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U35570 ( .A1(n4589), .A2(n4797), .ZN(n4575) );
  INV_X1 U35580 ( .A(n4575), .ZN(n2944) );
  NAND2_X1 U35590 ( .A1(n4063), .A2(n2945), .ZN(n2946) );
  OAI21_X1 U35600 ( .B1(n4080), .B2(n4832), .A(n4077), .ZN(n2947) );
  NOR2_X1 U35610 ( .A1(n2984), .A2(n2947), .ZN(n2948) );
  INV_X1 U35620 ( .A(n2984), .ZN(n4843) );
  INV_X1 U35630 ( .A(n2994), .ZN(n4089) );
  INV_X1 U35640 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2950) );
  INV_X1 U35650 ( .A(n2951), .ZN(n2949) );
  OAI21_X1 U35660 ( .B1(n4089), .B2(n2950), .A(n2949), .ZN(n4082) );
  NAND2_X1 U35670 ( .A1(n4099), .A2(REG1_REG_18__SCAN_IN), .ZN(n2952) );
  OAI211_X1 U35680 ( .C1(n4099), .C2(REG1_REG_18__SCAN_IN), .A(n4097), .B(
        n2952), .ZN(n4101) );
  OAI21_X1 U35690 ( .B1(n4103), .B2(n4914), .A(n4101), .ZN(n2955) );
  INV_X1 U35700 ( .A(REG1_REG_19__SCAN_IN), .ZN(n2953) );
  MUX2_X1 U35710 ( .A(REG1_REG_19__SCAN_IN), .B(n2953), .S(n4732), .Z(n2954)
         );
  INV_X1 U35720 ( .A(n4494), .ZN(n4603) );
  NAND2_X1 U35730 ( .A1(n4554), .A2(REG2_REG_11__SCAN_IN), .ZN(n2976) );
  INV_X1 U35740 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4771) );
  AOI22_X1 U35750 ( .A1(n4554), .A2(REG2_REG_11__SCAN_IN), .B1(n4771), .B2(
        n2940), .ZN(n4562) );
  NAND2_X1 U35760 ( .A1(n4543), .A2(REG2_REG_9__SCAN_IN), .ZN(n2972) );
  INV_X1 U35770 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2957) );
  AOI22_X1 U35780 ( .A1(n4543), .A2(REG2_REG_9__SCAN_IN), .B1(n2957), .B2(
        n4757), .ZN(n4551) );
  INV_X1 U35790 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2958) );
  MUX2_X1 U35800 ( .A(REG2_REG_2__SCAN_IN), .B(n2958), .S(n4615), .Z(n4613) );
  NAND2_X1 U35810 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n4601) );
  INV_X1 U3582 ( .A(n4601), .ZN(n3847) );
  NAND2_X1 U3583 ( .A1(n4488), .A2(REG2_REG_1__SCAN_IN), .ZN(n2959) );
  NAND2_X1 U3584 ( .A1(n3846), .A2(n2959), .ZN(n4612) );
  NOR2_X1 U3585 ( .A1(n2961), .A2(n2927), .ZN(n2962) );
  INV_X1 U3586 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4501) );
  NOR2_X1 U3587 ( .A1(n2964), .A2(n2428), .ZN(n2965) );
  INV_X1 U3588 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4636) );
  NAND2_X1 U3589 ( .A1(n4487), .A2(REG2_REG_5__SCAN_IN), .ZN(n2967) );
  OR2_X1 U3590 ( .A1(n4487), .A2(REG2_REG_5__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3591 ( .A1(n2967), .A2(n2966), .ZN(n3050) );
  NOR2_X1 U3592 ( .A1(n2295), .A2(n2342), .ZN(n2969) );
  INV_X1 U3593 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4510) );
  OR2_X1 U3594 ( .A1(n4748), .A2(n2970), .ZN(n2971) );
  NAND2_X1 U3595 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U3596 ( .A1(n2973), .A2(n2974), .ZN(n2975) );
  NAND2_X1 U3597 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4050), .ZN(n4049) );
  NAND2_X1 U3598 ( .A1(n2975), .A2(n4049), .ZN(n4561) );
  NAND2_X1 U3599 ( .A1(n4562), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U3600 ( .A1(n2976), .A2(n4560), .ZN(n2978) );
  NAND2_X1 U3601 ( .A1(n2977), .A2(n2978), .ZN(n2979) );
  XNOR2_X1 U3602 ( .A(n2978), .B(n4782), .ZN(n4572) );
  NAND2_X1 U3603 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4572), .ZN(n4571) );
  INV_X1 U3604 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4583) );
  NOR2_X1 U3605 ( .A1(n4589), .A2(n4583), .ZN(n4582) );
  INV_X1 U3606 ( .A(n4063), .ZN(n2980) );
  INV_X1 U3607 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U3608 ( .A1(n4486), .A2(REG2_REG_15__SCAN_IN), .ZN(n2983) );
  OR2_X1 U3609 ( .A1(n4486), .A2(REG2_REG_15__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U3610 ( .A1(n2983), .A2(n2982), .ZN(n4071) );
  NAND2_X1 U3611 ( .A1(n2985), .A2(n4843), .ZN(n2986) );
  INV_X1 U3612 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4591) );
  XNOR2_X1 U3613 ( .A(n4089), .B(REG2_REG_17__SCAN_IN), .ZN(n4085) );
  OAI21_X1 U3614 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2994), .A(n4084), .ZN(n4094) );
  INV_X1 U3615 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2988) );
  NOR2_X1 U3616 ( .A1(n4099), .A2(n2988), .ZN(n2987) );
  AOI21_X1 U3617 ( .B1(n2988), .B2(n4099), .A(n2987), .ZN(n4095) );
  INV_X1 U3618 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2989) );
  MUX2_X1 U3619 ( .A(n2989), .B(REG2_REG_19__SCAN_IN), .S(n4732), .Z(n2990) );
  NOR2_X1 U3620 ( .A1(n3044), .A2(n4603), .ZN(n4600) );
  INV_X1 U3621 ( .A(DATAI_14_), .ZN(n2992) );
  NAND2_X1 U3622 ( .A1(n4063), .A2(STATE_REG_SCAN_IN), .ZN(n2991) );
  OAI21_X1 U3623 ( .B1(STATE_REG_SCAN_IN), .B2(n2992), .A(n2991), .ZN(U3338)
         );
  INV_X1 U3624 ( .A(DATAI_21_), .ZN(n3861) );
  NAND2_X1 U3625 ( .A1(n3718), .A2(STATE_REG_SCAN_IN), .ZN(n2993) );
  OAI21_X1 U3626 ( .B1(STATE_REG_SCAN_IN), .B2(n3861), .A(n2993), .ZN(U3331)
         );
  INV_X1 U3627 ( .A(DATAI_17_), .ZN(n2996) );
  NAND2_X1 U3628 ( .A1(n2994), .A2(STATE_REG_SCAN_IN), .ZN(n2995) );
  OAI21_X1 U3629 ( .B1(STATE_REG_SCAN_IN), .B2(n2996), .A(n2995), .ZN(U3335)
         );
  INV_X1 U3630 ( .A(DATAI_22_), .ZN(n3860) );
  NAND2_X1 U3631 ( .A1(n3824), .A2(STATE_REG_SCAN_IN), .ZN(n2997) );
  OAI21_X1 U3632 ( .B1(STATE_REG_SCAN_IN), .B2(n3860), .A(n2997), .ZN(U3330)
         );
  INV_X1 U3633 ( .A(DATAI_24_), .ZN(n3970) );
  MUX2_X1 U3634 ( .A(n3970), .B(n2998), .S(STATE_REG_SCAN_IN), .Z(n2999) );
  INV_X1 U3635 ( .A(n2999), .ZN(U3328) );
  INV_X1 U3636 ( .A(DATAI_18_), .ZN(n3878) );
  NAND2_X1 U3637 ( .A1(n4099), .A2(STATE_REG_SCAN_IN), .ZN(n3000) );
  OAI21_X1 U3638 ( .B1(STATE_REG_SCAN_IN), .B2(n3878), .A(n3000), .ZN(U3334)
         );
  INV_X1 U3639 ( .A(DATAI_26_), .ZN(n3957) );
  NAND2_X1 U3640 ( .A1(n3008), .A2(STATE_REG_SCAN_IN), .ZN(n3001) );
  OAI21_X1 U3641 ( .B1(STATE_REG_SCAN_IN), .B2(n3957), .A(n3001), .ZN(U3326)
         );
  INV_X1 U3642 ( .A(DATAI_20_), .ZN(n3976) );
  NAND2_X1 U3643 ( .A1(n3813), .A2(STATE_REG_SCAN_IN), .ZN(n3002) );
  OAI21_X1 U3644 ( .B1(STATE_REG_SCAN_IN), .B2(n3976), .A(n3002), .ZN(U3332)
         );
  INV_X1 U3645 ( .A(DATAI_29_), .ZN(n3964) );
  NAND2_X1 U3646 ( .A1(n3003), .A2(STATE_REG_SCAN_IN), .ZN(n3004) );
  OAI21_X1 U3647 ( .B1(STATE_REG_SCAN_IN), .B2(n3964), .A(n3004), .ZN(U3323)
         );
  INV_X1 U3648 ( .A(DATAI_28_), .ZN(n3865) );
  INV_X1 U3649 ( .A(n3044), .ZN(n4604) );
  NAND2_X1 U3650 ( .A1(n4604), .A2(STATE_REG_SCAN_IN), .ZN(n3005) );
  OAI21_X1 U3651 ( .B1(STATE_REG_SCAN_IN), .B2(n3865), .A(n3005), .ZN(U3324)
         );
  INV_X1 U3652 ( .A(D_REG_0__SCAN_IN), .ZN(n3011) );
  INV_X1 U3653 ( .A(n3007), .ZN(n3042) );
  NOR3_X1 U3654 ( .A1(n3009), .A2(n3042), .A3(n3008), .ZN(n3010) );
  AOI21_X1 U3655 ( .B1(n4491), .B2(n3011), .A(n3010), .ZN(U3458) );
  NAND2_X1 U3656 ( .A1(n4491), .A2(D_REG_1__SCAN_IN), .ZN(n3012) );
  OAI21_X1 U3657 ( .B1(n4491), .B2(n3026), .A(n3012), .ZN(U3459) );
  NAND2_X1 U3658 ( .A1(n2700), .A2(REG1_REG_31__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U3659 ( .A1(n3013), .A2(REG2_REG_31__SCAN_IN), .ZN(n3015) );
  NAND2_X1 U3660 ( .A1(n2270), .A2(REG0_REG_31__SCAN_IN), .ZN(n3014) );
  AND3_X1 U3661 ( .A1(n3016), .A2(n3015), .A3(n3014), .ZN(n4106) );
  NAND2_X1 U3662 ( .A1(n3838), .A2(DATAO_REG_31__SCAN_IN), .ZN(n3017) );
  OAI21_X1 U3663 ( .B1(n4106), .B2(n3838), .A(n3017), .ZN(U3581) );
  AND2_X2 U3664 ( .A1(n3018), .A2(n3019), .ZN(n3542) );
  NOR2_X1 U3665 ( .A1(n4674), .A2(n3555), .ZN(n3020) );
  NAND2_X1 U3666 ( .A1(n3105), .A2(REG1_REG_0__SCAN_IN), .ZN(n3021) );
  NAND2_X2 U3667 ( .A1(n3249), .A2(n4898), .ZN(n3556) );
  AOI22_X1 U3668 ( .A1(n3022), .A2(n3542), .B1(n3105), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n3023) );
  OAI21_X1 U3669 ( .B1(n3025), .B2(n3024), .A(n3067), .ZN(n4605) );
  NOR2_X1 U3670 ( .A1(n3027), .A2(n3026), .ZN(n3122) );
  NOR2_X1 U3671 ( .A1(n3120), .A2(n3119), .ZN(n3028) );
  NAND2_X1 U3672 ( .A1(n3122), .A2(n3028), .ZN(n3071) );
  NAND2_X1 U3673 ( .A1(n3029), .A2(n4644), .ZN(n3032) );
  NAND3_X1 U3674 ( .A1(n3037), .A2(n3032), .A3(n3030), .ZN(n3031) );
  NAND2_X1 U3675 ( .A1(n3071), .A2(n3032), .ZN(n3034) );
  NAND2_X1 U3676 ( .A1(n3034), .A2(n3033), .ZN(n3106) );
  INV_X1 U3677 ( .A(n3106), .ZN(n3036) );
  NOR2_X1 U3678 ( .A1(n4862), .A2(U3149), .ZN(n3035) );
  NAND2_X1 U3679 ( .A1(n3071), .A2(n3035), .ZN(n3107) );
  NAND3_X1 U3680 ( .A1(n3036), .A2(n3037), .A3(n3107), .ZN(n3093) );
  NAND2_X1 U3681 ( .A1(n3037), .A2(n4902), .ZN(n3038) );
  OR2_X1 U3682 ( .A1(n3071), .A2(n3038), .ZN(n3041) );
  NAND2_X2 U3683 ( .A1(n3041), .A2(n4882), .ZN(n4973) );
  INV_X1 U3684 ( .A(n4973), .ZN(n4808) );
  NAND2_X1 U3685 ( .A1(n4732), .A2(n3824), .ZN(n3061) );
  NOR2_X1 U3686 ( .A1(n3061), .A2(n3042), .ZN(n3043) );
  NAND2_X1 U3687 ( .A1(n3822), .A2(n3044), .ZN(n3045) );
  OAI22_X1 U3688 ( .A1(n4808), .A2(n4674), .B1(n2604), .B2(n4934), .ZN(n3046)
         );
  AOI21_X1 U3689 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3093), .A(n3046), .ZN(n3047)
         );
  OAI21_X1 U3690 ( .B1(n4605), .B2(n4846), .A(n3047), .ZN(U3229) );
  INV_X1 U3691 ( .A(n4487), .ZN(n3058) );
  AND2_X1 U3692 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3168) );
  INV_X1 U3693 ( .A(n3048), .ZN(n3049) );
  AOI211_X1 U3694 ( .C1(n3051), .C2(n3050), .A(n3049), .B(n4633), .ZN(n3052)
         );
  AOI211_X1 U3695 ( .C1(n4629), .C2(ADDR_REG_5__SCAN_IN), .A(n3168), .B(n3052), 
        .ZN(n3057) );
  OAI211_X1 U3696 ( .C1(n3055), .C2(n3054), .A(n4630), .B(n3053), .ZN(n3056)
         );
  OAI211_X1 U3697 ( .C1(n4643), .C2(n3058), .A(n3057), .B(n3056), .ZN(U3245)
         );
  INV_X1 U3698 ( .A(n3093), .ZN(n3077) );
  INV_X1 U3699 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3700 ( .A1(n4662), .A2(n3249), .ZN(n3059) );
  NAND2_X1 U3701 ( .A1(n3060), .A2(n3059), .ZN(n3063) );
  NAND2_X4 U3702 ( .A1(n3062), .A2(n3061), .ZN(n3557) );
  NOR2_X1 U3703 ( .A1(n4675), .A2(n3347), .ZN(n3064) );
  AOI21_X2 U3704 ( .B1(n3837), .B2(n3467), .A(n3064), .ZN(n3082) );
  XNOR2_X1 U3705 ( .A(n3084), .B(n3082), .ZN(n3068) );
  NAND2_X1 U3706 ( .A1(n3065), .A2(n3545), .ZN(n3066) );
  NAND2_X1 U3707 ( .A1(n3067), .A2(n3066), .ZN(n3069) );
  OAI211_X1 U3708 ( .C1(n3068), .C2(n3069), .A(n3086), .B(n4974), .ZN(n3075)
         );
  NAND2_X1 U3709 ( .A1(n3822), .A2(n4604), .ZN(n3070) );
  OAI22_X1 U3710 ( .A1(n3072), .A2(n3612), .B1(n4665), .B2(n4934), .ZN(n3073)
         );
  AOI21_X1 U3711 ( .B1(n4662), .B2(n4973), .A(n3073), .ZN(n3074) );
  OAI211_X1 U3712 ( .C1(n3077), .C2(n3076), .A(n3075), .B(n3074), .ZN(U3219)
         );
  NAND2_X1 U3713 ( .A1(n3836), .A2(n3542), .ZN(n3079) );
  NAND2_X1 U3714 ( .A1(n3135), .A2(n3249), .ZN(n3078) );
  NAND2_X1 U3715 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  NOR2_X1 U3716 ( .A1(n3129), .A2(n3347), .ZN(n3081) );
  AOI21_X1 U3717 ( .B1(n3836), .B2(n3467), .A(n3081), .ZN(n3096) );
  XNOR2_X1 U3718 ( .A(n3097), .B(n3096), .ZN(n3090) );
  INV_X1 U3719 ( .A(n3082), .ZN(n3083) );
  NAND2_X1 U3720 ( .A1(n3084), .A2(n3083), .ZN(n3085) );
  INV_X1 U3721 ( .A(n3099), .ZN(n3088) );
  AOI21_X1 U3722 ( .B1(n3090), .B2(n3089), .A(n3088), .ZN(n3095) );
  INV_X2 U3723 ( .A(n3612), .ZN(n4970) );
  AOI22_X1 U3724 ( .A1(n4964), .A2(n3835), .B1(n4970), .B2(n3837), .ZN(n3091)
         );
  OAI21_X1 U3725 ( .B1(n4808), .B2(n3129), .A(n3091), .ZN(n3092) );
  AOI21_X1 U3726 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3093), .A(n3092), .ZN(n3094)
         );
  OAI21_X1 U3727 ( .B1(n3095), .B2(n4846), .A(n3094), .ZN(U3234) );
  NAND2_X1 U3728 ( .A1(n3097), .A2(n3096), .ZN(n3098) );
  NAND2_X1 U3729 ( .A1(n3099), .A2(n3098), .ZN(n3146) );
  NAND2_X1 U3730 ( .A1(n3835), .A2(n3542), .ZN(n3101) );
  NAND2_X1 U3731 ( .A1(n3214), .A2(n3249), .ZN(n3100) );
  NAND2_X1 U3732 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  NOR2_X1 U3733 ( .A1(n3103), .A2(n3347), .ZN(n3104) );
  AOI21_X1 U3734 ( .B1(n3835), .B2(n3467), .A(n3104), .ZN(n3148) );
  XNOR2_X1 U3735 ( .A(n3147), .B(n3148), .ZN(n3145) );
  XNOR2_X1 U3736 ( .A(n3146), .B(n3145), .ZN(n3113) );
  OAI21_X1 U3737 ( .B1(n3106), .B2(n3105), .A(STATE_REG_SCAN_IN), .ZN(n3109)
         );
  AND2_X1 U3738 ( .A1(n3107), .A2(n4489), .ZN(n3108) );
  AND2_X2 U3739 ( .A1(n3109), .A2(n3108), .ZN(n4979) );
  NOR2_X1 U3740 ( .A1(STATE_REG_SCAN_IN), .A2(n4696), .ZN(n4502) );
  AOI21_X1 U3741 ( .B1(n4964), .B2(n3834), .A(n4502), .ZN(n3111) );
  AOI22_X1 U3742 ( .A1(n4970), .A2(n3836), .B1(n4973), .B2(n3214), .ZN(n3110)
         );
  OAI211_X1 U3743 ( .C1(n4979), .C2(REG3_REG_3__SCAN_IN), .A(n3111), .B(n3110), 
        .ZN(n3112) );
  AOI21_X1 U3744 ( .B1(n3113), .B2(n4974), .A(n3112), .ZN(n3114) );
  INV_X1 U3745 ( .A(n3114), .ZN(U3215) );
  NAND2_X1 U3746 ( .A1(n3115), .A2(n3804), .ZN(n3116) );
  NAND2_X1 U3747 ( .A1(n3117), .A2(n3116), .ZN(n4688) );
  INV_X1 U3748 ( .A(n4688), .ZN(n3139) );
  NOR2_X1 U3749 ( .A1(n3119), .A2(n3118), .ZN(n3121) );
  NAND3_X1 U3750 ( .A1(n3122), .A2(n3121), .A3(n3120), .ZN(n3123) );
  NAND2_X1 U3751 ( .A1(n3018), .A2(n4485), .ZN(n4111) );
  INV_X1 U3752 ( .A(n4111), .ZN(n3124) );
  INV_X1 U3753 ( .A(n4776), .ZN(n4325) );
  NAND3_X1 U3754 ( .A1(n2615), .A2(n3719), .A3(n4659), .ZN(n3125) );
  NAND2_X1 U3755 ( .A1(n3126), .A2(n3125), .ZN(n3131) );
  NAND2_X1 U3756 ( .A1(n3835), .A2(n4869), .ZN(n3128) );
  NAND2_X1 U3757 ( .A1(n3837), .A2(n4903), .ZN(n3127) );
  OAI211_X1 U3758 ( .C1(n4862), .C2(n3129), .A(n3128), .B(n3127), .ZN(n3130)
         );
  AOI21_X1 U3759 ( .B1(n3131), .B2(n4909), .A(n3130), .ZN(n3133) );
  INV_X1 U3760 ( .A(n4669), .ZN(n4769) );
  NAND2_X1 U3761 ( .A1(n4688), .A2(n4769), .ZN(n3132) );
  NAND2_X1 U3762 ( .A1(n3133), .A2(n3132), .ZN(n4687) );
  MUX2_X1 U3763 ( .A(n4687), .B(REG2_REG_2__SCAN_IN), .S(n4893), .Z(n3134) );
  INV_X1 U3764 ( .A(n3134), .ZN(n3138) );
  NAND2_X1 U3765 ( .A1(n4770), .A2(n4732), .ZN(n4130) );
  AND2_X1 U3766 ( .A1(n4673), .A2(n3135), .ZN(n3136) );
  NOR2_X1 U3767 ( .A1(n3210), .A2(n3136), .ZN(n4691) );
  AOI22_X1 U3768 ( .A1(n4981), .A2(n4691), .B1(REG3_REG_2__SCAN_IN), .B2(n4920), .ZN(n3137) );
  OAI211_X1 U3769 ( .C1(n3139), .C2(n4325), .A(n3138), .B(n3137), .ZN(U3288)
         );
  NAND2_X1 U3770 ( .A1(n3834), .A2(n3542), .ZN(n3141) );
  NAND2_X1 U3771 ( .A1(n3196), .A2(n3249), .ZN(n3140) );
  NAND2_X1 U3772 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  XNOR2_X1 U3773 ( .A(n3142), .B(n3545), .ZN(n3155) );
  NOR2_X1 U3774 ( .A1(n3143), .A2(n3347), .ZN(n3144) );
  AOI21_X1 U3775 ( .B1(n3834), .B2(n3467), .A(n3144), .ZN(n3156) );
  XNOR2_X1 U3776 ( .A(n3155), .B(n3156), .ZN(n3160) );
  AOI211_X1 U3777 ( .C1(n3160), .C2(n3161), .A(n4846), .B(n2318), .ZN(n3154)
         );
  INV_X1 U3778 ( .A(n3193), .ZN(n3152) );
  NOR2_X1 U3779 ( .A1(STATE_REG_SCAN_IN), .A2(n4016), .ZN(n4628) );
  AOI21_X1 U3780 ( .B1(n4964), .B2(n3833), .A(n4628), .ZN(n3151) );
  AOI22_X1 U3781 ( .A1(n4970), .A2(n3835), .B1(n4973), .B2(n3196), .ZN(n3150)
         );
  OAI211_X1 U3782 ( .C1(n4979), .C2(n3152), .A(n3151), .B(n3150), .ZN(n3153)
         );
  OR2_X1 U3783 ( .A1(n3154), .A2(n3153), .ZN(U3227) );
  INV_X1 U3784 ( .A(n3155), .ZN(n3158) );
  INV_X1 U3785 ( .A(n3156), .ZN(n3157) );
  NAND2_X1 U3786 ( .A1(n3158), .A2(n3157), .ZN(n3159) );
  NAND2_X1 U3787 ( .A1(n3833), .A2(n3542), .ZN(n3163) );
  NAND2_X1 U3788 ( .A1(n3181), .A2(n3249), .ZN(n3162) );
  NAND2_X1 U3789 ( .A1(n3163), .A2(n3162), .ZN(n3164) );
  XNOR2_X1 U3790 ( .A(n3164), .B(n3557), .ZN(n3218) );
  NAND2_X1 U3791 ( .A1(n3833), .A2(n3548), .ZN(n3166) );
  NAND2_X1 U3792 ( .A1(n3181), .A2(n3542), .ZN(n3165) );
  NAND2_X1 U3793 ( .A1(n3166), .A2(n3165), .ZN(n3219) );
  XNOR2_X1 U3794 ( .A(n3218), .B(n3219), .ZN(n3167) );
  XNOR2_X1 U3795 ( .A(n3220), .B(n3167), .ZN(n3172) );
  AOI21_X1 U3796 ( .B1(n4970), .B2(n3834), .A(n3168), .ZN(n3170) );
  AOI22_X1 U3797 ( .A1(n4964), .A2(n3832), .B1(n4973), .B2(n3181), .ZN(n3169)
         );
  OAI211_X1 U3798 ( .C1(n4979), .C2(n4327), .A(n3170), .B(n3169), .ZN(n3171)
         );
  AOI21_X1 U3799 ( .B1(n3172), .B2(n4974), .A(n3171), .ZN(n3173) );
  INV_X1 U3800 ( .A(n3173), .ZN(U3224) );
  NAND2_X1 U3801 ( .A1(n3706), .A2(n3725), .ZN(n3780) );
  XOR2_X1 U3802 ( .A(n3174), .B(n3780), .Z(n4326) );
  XOR2_X1 U3803 ( .A(n3780), .B(n3175), .Z(n3180) );
  OAI22_X1 U3804 ( .A1(n3177), .A2(n4726), .B1(n3176), .B2(n4862), .ZN(n3178)
         );
  AOI21_X1 U3805 ( .B1(n4869), .B2(n3832), .A(n3178), .ZN(n3179) );
  OAI21_X1 U3806 ( .B1(n3180), .B2(n4864), .A(n3179), .ZN(n4329) );
  AOI21_X1 U3807 ( .B1(n4326), .B2(n4912), .A(n4329), .ZN(n3185) );
  AND2_X1 U3808 ( .A1(n3194), .A2(n3181), .ZN(n3182) );
  NOR2_X1 U3809 ( .A1(n3280), .A2(n3182), .ZN(n4330) );
  INV_X1 U3810 ( .A(n4482), .ZN(n4692) );
  AOI22_X1 U3811 ( .A1(n4330), .A2(n4692), .B1(REG0_REG_5__SCAN_IN), .B2(n4916), .ZN(n3183) );
  OAI21_X1 U3812 ( .B1(n3185), .B2(n4916), .A(n3183), .ZN(U3477) );
  INV_X1 U3813 ( .A(n4431), .ZN(n4689) );
  AOI22_X1 U3814 ( .A1(n4330), .A2(n4689), .B1(REG1_REG_5__SCAN_IN), .B2(n4913), .ZN(n3184) );
  OAI21_X1 U3815 ( .B1(n3185), .B2(n4913), .A(n3184), .ZN(U3523) );
  XNOR2_X1 U3816 ( .A(n3186), .B(n3782), .ZN(n3197) );
  NAND2_X1 U3817 ( .A1(n3202), .A2(n3187), .ZN(n3188) );
  XOR2_X1 U3818 ( .A(n3782), .B(n3188), .Z(n3191) );
  AOI22_X1 U3819 ( .A1(n3835), .A2(n4903), .B1(n3196), .B2(n4902), .ZN(n3189)
         );
  OAI21_X1 U3820 ( .B1(n3275), .B2(n4906), .A(n3189), .ZN(n3190) );
  AOI21_X1 U3821 ( .B1(n3191), .B2(n4909), .A(n3190), .ZN(n3192) );
  OAI21_X1 U3822 ( .B1(n3197), .B2(n4669), .A(n3192), .ZN(n4703) );
  AOI21_X1 U3823 ( .B1(n3193), .B2(n4920), .A(n4703), .ZN(n3200) );
  INV_X1 U3824 ( .A(n3194), .ZN(n3195) );
  AOI211_X1 U3825 ( .C1(n3196), .C2(n3211), .A(n4898), .B(n3195), .ZN(n4704)
         );
  INV_X1 U3826 ( .A(n4130), .ZN(n4923) );
  AOI22_X1 U3827 ( .A1(n4704), .A2(n4923), .B1(REG2_REG_4__SCAN_IN), .B2(n4893), .ZN(n3199) );
  INV_X1 U3828 ( .A(n3197), .ZN(n4706) );
  NAND2_X1 U3829 ( .A1(n4706), .A2(n4776), .ZN(n3198) );
  OAI211_X1 U3830 ( .C1(n3200), .C2(n4893), .A(n3199), .B(n3198), .ZN(U3286)
         );
  XNOR2_X1 U3831 ( .A(n3201), .B(n3803), .ZN(n3205) );
  INV_X1 U3832 ( .A(n3205), .ZN(n4698) );
  OAI21_X1 U3833 ( .B1(n3803), .B2(n3203), .A(n3202), .ZN(n3208) );
  AOI22_X1 U3834 ( .A1(n3834), .A2(n4869), .B1(n4902), .B2(n3214), .ZN(n3204)
         );
  OAI21_X1 U3835 ( .B1(n4665), .B2(n4726), .A(n3204), .ZN(n3207) );
  NOR2_X1 U3836 ( .A1(n3205), .A2(n4669), .ZN(n3206) );
  AOI211_X1 U3837 ( .C1(n4909), .C2(n3208), .A(n3207), .B(n3206), .ZN(n4701)
         );
  INV_X1 U3838 ( .A(n4701), .ZN(n3209) );
  AOI21_X1 U3839 ( .B1(n4705), .B2(n4698), .A(n3209), .ZN(n3217) );
  INV_X1 U3840 ( .A(n3210), .ZN(n3213) );
  INV_X1 U3841 ( .A(n3211), .ZN(n3212) );
  AOI21_X1 U3842 ( .B1(n3214), .B2(n3213), .A(n3212), .ZN(n4697) );
  AOI22_X1 U3843 ( .A1(n4697), .A2(n4689), .B1(REG1_REG_3__SCAN_IN), .B2(n4913), .ZN(n3215) );
  OAI21_X1 U3844 ( .B1(n3217), .B2(n4913), .A(n3215), .ZN(U3521) );
  AOI22_X1 U3845 ( .A1(n4697), .A2(n4692), .B1(REG0_REG_3__SCAN_IN), .B2(n4916), .ZN(n3216) );
  OAI21_X1 U3846 ( .B1(n3217), .B2(n4916), .A(n3216), .ZN(U3473) );
  NAND2_X1 U3847 ( .A1(n3832), .A2(n3542), .ZN(n3223) );
  NAND2_X1 U3848 ( .A1(n3273), .A2(n3249), .ZN(n3222) );
  NAND2_X1 U3849 ( .A1(n3223), .A2(n3222), .ZN(n3224) );
  XNOR2_X1 U3850 ( .A(n3224), .B(n3557), .ZN(n3227) );
  NAND2_X1 U3851 ( .A1(n3832), .A2(n3548), .ZN(n3226) );
  NAND2_X1 U3852 ( .A1(n3273), .A2(n3542), .ZN(n3225) );
  NAND2_X1 U3853 ( .A1(n3226), .A2(n3225), .ZN(n3228) );
  INV_X1 U3854 ( .A(n3227), .ZN(n3230) );
  INV_X1 U3855 ( .A(n3228), .ZN(n3229) );
  NAND2_X1 U3856 ( .A1(n3230), .A2(n3229), .ZN(n3240) );
  NAND2_X1 U3857 ( .A1(n2324), .A2(n3240), .ZN(n3231) );
  XNOR2_X1 U3858 ( .A(n3239), .B(n3231), .ZN(n3237) );
  INV_X1 U3859 ( .A(n4711), .ZN(n3235) );
  NOR2_X1 U3860 ( .A1(STATE_REG_SCAN_IN), .A2(n3232), .ZN(n4511) );
  AOI21_X1 U3861 ( .B1(n4964), .B2(n3831), .A(n4511), .ZN(n3234) );
  AOI22_X1 U3862 ( .A1(n4970), .A2(n3833), .B1(n4973), .B2(n3273), .ZN(n3233)
         );
  OAI211_X1 U3863 ( .C1(n4979), .C2(n3235), .A(n3234), .B(n3233), .ZN(n3236)
         );
  AOI21_X1 U3864 ( .B1(n3237), .B2(n4974), .A(n3236), .ZN(n3238) );
  INV_X1 U3865 ( .A(n3238), .ZN(U3236) );
  NAND2_X1 U3866 ( .A1(n3831), .A2(n3392), .ZN(n3242) );
  NAND2_X1 U3867 ( .A1(n4723), .A2(n3249), .ZN(n3241) );
  NAND2_X1 U3868 ( .A1(n3242), .A2(n3241), .ZN(n3243) );
  XNOR2_X1 U3869 ( .A(n3243), .B(n3557), .ZN(n3247) );
  NOR2_X1 U3870 ( .A1(n4725), .A2(n3347), .ZN(n3244) );
  AOI21_X1 U3871 ( .B1(n3831), .B2(n3467), .A(n3244), .ZN(n3245) );
  XNOR2_X1 U3872 ( .A(n3247), .B(n3245), .ZN(n3571) );
  NAND2_X1 U3873 ( .A1(n3572), .A2(n3571), .ZN(n3570) );
  INV_X1 U3874 ( .A(n3245), .ZN(n3246) );
  NAND2_X1 U3875 ( .A1(n3247), .A2(n3246), .ZN(n3248) );
  NAND2_X1 U3876 ( .A1(n4729), .A2(n3392), .ZN(n3251) );
  NAND2_X1 U3877 ( .A1(n3263), .A2(n3249), .ZN(n3250) );
  NAND2_X1 U3878 ( .A1(n3251), .A2(n3250), .ZN(n3252) );
  XNOR2_X1 U3879 ( .A(n3252), .B(n3557), .ZN(n3255) );
  NAND2_X1 U3880 ( .A1(n4729), .A2(n3548), .ZN(n3254) );
  NAND2_X1 U3881 ( .A1(n3263), .A2(n3392), .ZN(n3253) );
  NAND2_X1 U3882 ( .A1(n3254), .A2(n3253), .ZN(n3256) );
  NAND2_X1 U3883 ( .A1(n3255), .A2(n3256), .ZN(n3260) );
  INV_X1 U3884 ( .A(n3303), .ZN(n3262) );
  INV_X1 U3885 ( .A(n3255), .ZN(n3258) );
  INV_X1 U3886 ( .A(n3256), .ZN(n3257) );
  NAND2_X1 U3887 ( .A1(n3258), .A2(n3257), .ZN(n3302) );
  AOI21_X1 U3888 ( .B1(n3302), .B2(n3260), .A(n3259), .ZN(n3261) );
  AOI21_X1 U3889 ( .B1(n3262), .B2(n3302), .A(n3261), .ZN(n3269) );
  INV_X1 U3890 ( .A(n4749), .ZN(n3266) );
  AOI22_X1 U3891 ( .A1(n4964), .A2(n3830), .B1(REG3_REG_8__SCAN_IN), .B2(U3149), .ZN(n3265) );
  AOI22_X1 U3892 ( .A1(n4970), .A2(n3831), .B1(n4973), .B2(n3263), .ZN(n3264)
         );
  OAI211_X1 U3893 ( .C1(n4979), .C2(n3266), .A(n3265), .B(n3264), .ZN(n3267)
         );
  INV_X1 U3894 ( .A(n3267), .ZN(n3268) );
  OAI21_X1 U3895 ( .B1(n3269), .B2(n4846), .A(n3268), .ZN(U3218) );
  XNOR2_X1 U3896 ( .A(n3270), .B(n3801), .ZN(n4712) );
  XNOR2_X1 U3897 ( .A(n3272), .B(n3801), .ZN(n3278) );
  AOI22_X1 U3898 ( .A1(n3831), .A2(n4869), .B1(n4902), .B2(n3273), .ZN(n3274)
         );
  OAI21_X1 U3899 ( .B1(n3275), .B2(n4726), .A(n3274), .ZN(n3277) );
  NOR2_X1 U3900 ( .A1(n4712), .A2(n4669), .ZN(n3276) );
  AOI211_X1 U3901 ( .C1(n3278), .C2(n4909), .A(n3277), .B(n3276), .ZN(n4718)
         );
  OAI21_X1 U3902 ( .B1(n4712), .B2(n4792), .A(n4718), .ZN(n3287) );
  NOR2_X1 U3903 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  OR2_X1 U3904 ( .A1(n4721), .A2(n3281), .ZN(n4713) );
  INV_X1 U3905 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3282) );
  OAI22_X1 U3906 ( .A1(n4713), .A2(n4482), .B1(n4919), .B2(n3282), .ZN(n3283)
         );
  AOI21_X1 U3907 ( .B1(n3287), .B2(n4919), .A(n3283), .ZN(n3284) );
  INV_X1 U3908 ( .A(n3284), .ZN(U3479) );
  INV_X1 U3909 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3285) );
  OAI22_X1 U3910 ( .A1(n4713), .A2(n4431), .B1(n4915), .B2(n3285), .ZN(n3286)
         );
  AOI21_X1 U3911 ( .B1(n3287), .B2(n4915), .A(n3286), .ZN(n3288) );
  INV_X1 U3912 ( .A(n3288), .ZN(U3524) );
  OAI21_X1 U3913 ( .B1(n3326), .B2(n2317), .A(n3289), .ZN(n3290) );
  AND2_X1 U3914 ( .A1(n3738), .A2(n3704), .ZN(n3802) );
  XNOR2_X1 U3915 ( .A(n3290), .B(n3802), .ZN(n3296) );
  XOR2_X1 U3916 ( .A(n3802), .B(n3291), .Z(n3294) );
  AOI22_X1 U3917 ( .A1(n4729), .A2(n4903), .B1(n4902), .B2(n3311), .ZN(n3292)
         );
  OAI21_X1 U3918 ( .B1(n3377), .B2(n4906), .A(n3292), .ZN(n3293) );
  AOI21_X1 U3919 ( .B1(n3294), .B2(n4909), .A(n3293), .ZN(n3295) );
  OAI21_X1 U3920 ( .B1(n3296), .B2(n4669), .A(n3295), .ZN(n3318) );
  INV_X1 U3921 ( .A(n3318), .ZN(n3301) );
  INV_X1 U3922 ( .A(n3296), .ZN(n3319) );
  INV_X1 U3923 ( .A(n3325), .ZN(n3297) );
  OAI21_X1 U3924 ( .B1(n3297), .B2(n3307), .A(n2363), .ZN(n3324) );
  AOI22_X1 U3925 ( .A1(n4893), .A2(REG2_REG_9__SCAN_IN), .B1(n3309), .B2(n4920), .ZN(n3298) );
  OAI21_X1 U3926 ( .B1(n3324), .B2(n4886), .A(n3298), .ZN(n3299) );
  AOI21_X1 U3927 ( .B1(n3319), .B2(n4776), .A(n3299), .ZN(n3300) );
  OAI21_X1 U3928 ( .B1(n3301), .B2(n4893), .A(n3300), .ZN(U3281) );
  NAND2_X1 U3929 ( .A1(n3830), .A2(n3392), .ZN(n3305) );
  NAND2_X1 U3930 ( .A1(n3311), .A2(n3249), .ZN(n3304) );
  NAND2_X1 U3931 ( .A1(n3305), .A2(n3304), .ZN(n3306) );
  XNOR2_X1 U3932 ( .A(n3306), .B(n3557), .ZN(n3340) );
  NOR2_X1 U3933 ( .A1(n3307), .A2(n3347), .ZN(n3308) );
  AOI21_X1 U3934 ( .B1(n3830), .B2(n3467), .A(n3308), .ZN(n3341) );
  XNOR2_X1 U3935 ( .A(n3340), .B(n3341), .ZN(n3338) );
  XNOR2_X1 U3936 ( .A(n3339), .B(n3338), .ZN(n3316) );
  INV_X1 U3937 ( .A(n3309), .ZN(n3314) );
  NOR2_X1 U3938 ( .A1(STATE_REG_SCAN_IN), .A2(n3310), .ZN(n4547) );
  AOI21_X1 U3939 ( .B1(n4964), .B2(n3829), .A(n4547), .ZN(n3313) );
  AOI22_X1 U3940 ( .A1(n4970), .A2(n4729), .B1(n4973), .B2(n3311), .ZN(n3312)
         );
  OAI211_X1 U3941 ( .C1(n4979), .C2(n3314), .A(n3313), .B(n3312), .ZN(n3315)
         );
  AOI21_X1 U3942 ( .B1(n3316), .B2(n4974), .A(n3315), .ZN(n3317) );
  INV_X1 U3943 ( .A(n3317), .ZN(U3228) );
  AOI21_X1 U3944 ( .B1(n4705), .B2(n3319), .A(n3318), .ZN(n3321) );
  MUX2_X1 U3945 ( .A(n4542), .B(n3321), .S(n4915), .Z(n3320) );
  OAI21_X1 U3946 ( .B1(n4431), .B2(n3324), .A(n3320), .ZN(U3527) );
  INV_X1 U3947 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3322) );
  MUX2_X1 U3948 ( .A(n3322), .B(n3321), .S(n4919), .Z(n3323) );
  OAI21_X1 U3949 ( .B1(n3324), .B2(n4482), .A(n3323), .ZN(U3485) );
  OAI21_X1 U3950 ( .B1(n2316), .B2(n3328), .A(n3325), .ZN(n4750) );
  INV_X1 U3951 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U3952 ( .A1(n3739), .A2(n3703), .ZN(n3779) );
  XOR2_X1 U3953 ( .A(n3779), .B(n3326), .Z(n4752) );
  XOR2_X1 U3954 ( .A(n3779), .B(n3327), .Z(n3331) );
  OAI22_X1 U3955 ( .A1(n3418), .A2(n4906), .B1(n3328), .B2(n4862), .ZN(n3329)
         );
  AOI21_X1 U3956 ( .B1(n4903), .B2(n3831), .A(n3329), .ZN(n3330) );
  OAI21_X1 U3957 ( .B1(n3331), .B2(n4864), .A(n3330), .ZN(n3332) );
  AOI21_X1 U3958 ( .B1(n4752), .B2(n4769), .A(n3332), .ZN(n4755) );
  INV_X1 U3959 ( .A(n4755), .ZN(n3333) );
  AOI21_X1 U3960 ( .B1(n4705), .B2(n4752), .A(n3333), .ZN(n3336) );
  MUX2_X1 U3961 ( .A(n3334), .B(n3336), .S(n4919), .Z(n3335) );
  OAI21_X1 U3962 ( .B1(n4750), .B2(n4482), .A(n3335), .ZN(U3483) );
  MUX2_X1 U3963 ( .A(n4534), .B(n3336), .S(n4915), .Z(n3337) );
  OAI21_X1 U3964 ( .B1(n4750), .B2(n4431), .A(n3337), .ZN(U3526) );
  INV_X1 U3965 ( .A(n3340), .ZN(n3342) );
  NAND2_X1 U3966 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  NAND2_X1 U3967 ( .A1(n3829), .A2(n3392), .ZN(n3345) );
  NAND2_X1 U3968 ( .A1(n3416), .A2(n3249), .ZN(n3344) );
  NAND2_X1 U3969 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  XNOR2_X1 U3970 ( .A(n3346), .B(n3545), .ZN(n3350) );
  NOR2_X1 U3971 ( .A1(n3412), .A2(n3347), .ZN(n3348) );
  AOI21_X1 U3972 ( .B1(n3829), .B2(n3467), .A(n3348), .ZN(n3351) );
  XNOR2_X1 U3973 ( .A(n3350), .B(n3351), .ZN(n3369) );
  INV_X1 U3974 ( .A(n3369), .ZN(n3349) );
  INV_X1 U3975 ( .A(n3350), .ZN(n3353) );
  INV_X1 U3976 ( .A(n3351), .ZN(n3352) );
  NAND2_X1 U3977 ( .A1(n3353), .A2(n3352), .ZN(n3354) );
  NAND2_X1 U3978 ( .A1(n4424), .A2(n3542), .ZN(n3356) );
  NAND2_X1 U3979 ( .A1(n3360), .A2(n3249), .ZN(n3355) );
  NAND2_X1 U3980 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  XNOR2_X1 U3981 ( .A(n3357), .B(n3545), .ZN(n3387) );
  NOR2_X1 U3982 ( .A1(n3376), .A2(n3347), .ZN(n3358) );
  AOI21_X1 U3983 ( .B1(n4424), .B2(n3467), .A(n3358), .ZN(n3388) );
  XNOR2_X1 U3984 ( .A(n3387), .B(n3388), .ZN(n3359) );
  XNOR2_X1 U3985 ( .A(n3386), .B(n3359), .ZN(n3364) );
  AND2_X1 U3986 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4558) );
  AOI21_X1 U3987 ( .B1(n4964), .B2(n4313), .A(n4558), .ZN(n3362) );
  AOI22_X1 U3988 ( .A1(n4970), .A2(n3829), .B1(n4973), .B2(n3360), .ZN(n3361)
         );
  OAI211_X1 U3989 ( .C1(n4979), .C2(n4772), .A(n3362), .B(n3361), .ZN(n3363)
         );
  AOI21_X1 U3990 ( .B1(n3364), .B2(n4974), .A(n3363), .ZN(n3365) );
  INV_X1 U3991 ( .A(n3365), .ZN(U3233) );
  INV_X1 U3992 ( .A(n3366), .ZN(n3367) );
  AOI211_X1 U3993 ( .C1(n3369), .C2(n3368), .A(n4846), .B(n3367), .ZN(n3374)
         );
  INV_X1 U3994 ( .A(n4760), .ZN(n3372) );
  AND2_X1 U3995 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4054) );
  AOI21_X1 U3996 ( .B1(n4970), .B2(n3830), .A(n4054), .ZN(n3371) );
  AOI22_X1 U3997 ( .A1(n4964), .A2(n4424), .B1(n4973), .B2(n3416), .ZN(n3370)
         );
  OAI211_X1 U3998 ( .C1(n4979), .C2(n3372), .A(n3371), .B(n3370), .ZN(n3373)
         );
  OR2_X1 U3999 ( .A1(n3374), .A2(n3373), .ZN(U3214) );
  OAI21_X1 U4000 ( .B1(n3410), .B2(n3376), .A(n4416), .ZN(n4774) );
  XNOR2_X1 U4001 ( .A(n3375), .B(n3781), .ZN(n4777) );
  XNOR2_X1 U4002 ( .A(n4307), .B(n3781), .ZN(n3380) );
  OAI22_X1 U4003 ( .A1(n3377), .A2(n4726), .B1(n4862), .B2(n3376), .ZN(n3378)
         );
  AOI21_X1 U4004 ( .B1(n4869), .B2(n4313), .A(n3378), .ZN(n3379) );
  OAI21_X1 U4005 ( .B1(n3380), .B2(n4864), .A(n3379), .ZN(n4768) );
  AOI21_X1 U4006 ( .B1(n4912), .B2(n4777), .A(n4768), .ZN(n3382) );
  MUX2_X1 U4007 ( .A(n2939), .B(n3382), .S(n4915), .Z(n3381) );
  OAI21_X1 U4008 ( .B1(n4431), .B2(n4774), .A(n3381), .ZN(U3529) );
  INV_X1 U4009 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3383) );
  MUX2_X1 U4010 ( .A(n3383), .B(n3382), .S(n4919), .Z(n3384) );
  OAI21_X1 U4011 ( .B1(n4774), .B2(n4482), .A(n3384), .ZN(U3489) );
  NAND2_X1 U4012 ( .A1(n3387), .A2(n3388), .ZN(n3385) );
  INV_X1 U4013 ( .A(n3387), .ZN(n3390) );
  INV_X1 U4014 ( .A(n3388), .ZN(n3389) );
  NAND2_X1 U4015 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NAND2_X1 U4016 ( .A1(n4313), .A2(n3392), .ZN(n3394) );
  NAND2_X1 U4017 ( .A1(n4423), .A2(n3249), .ZN(n3393) );
  NAND2_X1 U4018 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  XNOR2_X1 U4019 ( .A(n3395), .B(n3557), .ZN(n3398) );
  NAND2_X1 U4020 ( .A1(n4313), .A2(n3548), .ZN(n3397) );
  NAND2_X1 U4021 ( .A1(n4423), .A2(n3542), .ZN(n3396) );
  NAND2_X1 U4022 ( .A1(n3397), .A2(n3396), .ZN(n3399) );
  AND2_X1 U4023 ( .A1(n3398), .A2(n3399), .ZN(n3434) );
  INV_X1 U4024 ( .A(n3434), .ZN(n3402) );
  INV_X1 U4025 ( .A(n3398), .ZN(n3401) );
  INV_X1 U4026 ( .A(n3399), .ZN(n3400) );
  NAND2_X1 U4027 ( .A1(n3401), .A2(n3400), .ZN(n3436) );
  NAND2_X1 U4028 ( .A1(n3402), .A2(n3436), .ZN(n3403) );
  XNOR2_X1 U4029 ( .A(n3435), .B(n3403), .ZN(n3408) );
  INV_X1 U4030 ( .A(n4783), .ZN(n3406) );
  INV_X1 U4031 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3947) );
  NOR2_X1 U4032 ( .A1(STATE_REG_SCAN_IN), .A2(n3947), .ZN(n4569) );
  AOI21_X1 U4033 ( .B1(n4964), .B2(n4407), .A(n4569), .ZN(n3405) );
  AOI22_X1 U4034 ( .A1(n4970), .A2(n4424), .B1(n4973), .B2(n4423), .ZN(n3404)
         );
  OAI211_X1 U4035 ( .C1(n4979), .C2(n3406), .A(n3405), .B(n3404), .ZN(n3407)
         );
  AOI21_X1 U4036 ( .B1(n3408), .B2(n4974), .A(n3407), .ZN(n3409) );
  INV_X1 U4037 ( .A(n3409), .ZN(U3221) );
  INV_X1 U4038 ( .A(n3410), .ZN(n3411) );
  OAI21_X1 U4039 ( .B1(n3413), .B2(n3412), .A(n3411), .ZN(n4761) );
  INV_X1 U4040 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4041 ( .A1(n3707), .A2(n3708), .ZN(n3774) );
  XNOR2_X1 U4042 ( .A(n3414), .B(n3774), .ZN(n3419) );
  INV_X1 U40430 ( .A(n3419), .ZN(n4763) );
  XOR2_X1 U4044 ( .A(n3774), .B(n3415), .Z(n3422) );
  AOI22_X1 U4045 ( .A1(n4424), .A2(n4869), .B1(n3416), .B2(n4902), .ZN(n3417)
         );
  OAI21_X1 U4046 ( .B1(n3418), .B2(n4726), .A(n3417), .ZN(n3421) );
  NOR2_X1 U4047 ( .A1(n3419), .A2(n4669), .ZN(n3420) );
  AOI211_X1 U4048 ( .C1(n3422), .C2(n4909), .A(n3421), .B(n3420), .ZN(n4766)
         );
  INV_X1 U4049 ( .A(n4766), .ZN(n3423) );
  AOI21_X1 U4050 ( .B1(n4705), .B2(n4763), .A(n3423), .ZN(n3426) );
  MUX2_X1 U4051 ( .A(n3424), .B(n3426), .S(n4915), .Z(n3425) );
  OAI21_X1 U4052 ( .B1(n4761), .B2(n4431), .A(n3425), .ZN(U3528) );
  INV_X1 U4053 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3427) );
  MUX2_X1 U4054 ( .A(n3427), .B(n3426), .S(n4919), .Z(n3428) );
  OAI21_X1 U4055 ( .B1(n4761), .B2(n4482), .A(n3428), .ZN(U3487) );
  AND2_X1 U4056 ( .A1(n3429), .A2(n3838), .ZN(U3148) );
  NOR2_X1 U4057 ( .A1(n4203), .A2(n3347), .ZN(n3430) );
  AOI21_X1 U4058 ( .B1(n4225), .B2(n3548), .A(n3430), .ZN(n3630) );
  NAND2_X1 U4059 ( .A1(n4225), .A2(n3392), .ZN(n3432) );
  NAND2_X1 U4060 ( .A1(n3633), .A2(n3249), .ZN(n3431) );
  NAND2_X1 U4061 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  XNOR2_X1 U4062 ( .A(n3433), .B(n3545), .ZN(n3606) );
  NAND2_X1 U4063 ( .A1(n4407), .A2(n3392), .ZN(n3438) );
  NAND2_X1 U4064 ( .A1(n4320), .A2(n3249), .ZN(n3437) );
  NAND2_X1 U4065 ( .A1(n3438), .A2(n3437), .ZN(n3439) );
  XNOR2_X1 U4066 ( .A(n3439), .B(n3545), .ZN(n3640) );
  NAND2_X1 U4067 ( .A1(n4407), .A2(n3548), .ZN(n3441) );
  NAND2_X1 U4068 ( .A1(n4320), .A2(n3392), .ZN(n3440) );
  NAND2_X1 U4069 ( .A1(n3441), .A2(n3440), .ZN(n3639) );
  NAND2_X1 U4070 ( .A1(n3442), .A2(n3639), .ZN(n3445) );
  INV_X1 U4071 ( .A(n3640), .ZN(n3443) );
  NAND2_X1 U4072 ( .A1(n4823), .A2(n3392), .ZN(n3447) );
  NAND2_X1 U4073 ( .A1(n3588), .A2(n3249), .ZN(n3446) );
  NAND2_X1 U4074 ( .A1(n3447), .A2(n3446), .ZN(n3448) );
  XNOR2_X1 U4075 ( .A(n3448), .B(n3557), .ZN(n3451) );
  NAND2_X1 U4076 ( .A1(n4823), .A2(n3548), .ZN(n3450) );
  NAND2_X1 U4077 ( .A1(n3588), .A2(n3392), .ZN(n3449) );
  NAND2_X1 U4078 ( .A1(n3450), .A2(n3449), .ZN(n3452) );
  INV_X1 U4079 ( .A(n3451), .ZN(n3454) );
  INV_X1 U4080 ( .A(n3452), .ZN(n3453) );
  NAND2_X1 U4081 ( .A1(n3454), .A2(n3453), .ZN(n3585) );
  NAND2_X1 U4082 ( .A1(n4859), .A2(n3392), .ZN(n3457) );
  NAND2_X1 U4083 ( .A1(n3455), .A2(n3249), .ZN(n3456) );
  NAND2_X1 U4084 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  XNOR2_X1 U4085 ( .A(n3458), .B(n3545), .ZN(n3460) );
  NOR2_X1 U4086 ( .A1(n4825), .A2(n3347), .ZN(n3459) );
  AOI21_X1 U4087 ( .B1(n4859), .B2(n3548), .A(n3459), .ZN(n4814) );
  NAND2_X1 U4088 ( .A1(n4830), .A2(n3392), .ZN(n3464) );
  NAND2_X1 U4089 ( .A1(n4855), .A2(n3249), .ZN(n3463) );
  NAND2_X1 U4090 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  XNOR2_X1 U4091 ( .A(n3465), .B(n3557), .ZN(n3468) );
  NOR2_X1 U4092 ( .A1(n4861), .A2(n3347), .ZN(n3466) );
  AOI21_X1 U4093 ( .B1(n4830), .B2(n3467), .A(n3466), .ZN(n3469) );
  XNOR2_X1 U4094 ( .A(n3468), .B(n3469), .ZN(n4845) );
  INV_X1 U4095 ( .A(n3468), .ZN(n3470) );
  NAND2_X1 U4096 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  NAND2_X1 U4097 ( .A1(n4904), .A2(n3392), .ZN(n3473) );
  NAND2_X1 U4098 ( .A1(n4391), .A2(n3249), .ZN(n3472) );
  NAND2_X1 U4099 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  XNOR2_X1 U4100 ( .A(n3474), .B(n3545), .ZN(n3620) );
  NOR2_X1 U4101 ( .A1(n4387), .A2(n3347), .ZN(n3475) );
  AOI21_X1 U4102 ( .B1(n4904), .B2(n3548), .A(n3475), .ZN(n3476) );
  AND2_X1 U4103 ( .A1(n3620), .A2(n3476), .ZN(n3478) );
  INV_X1 U4104 ( .A(n3620), .ZN(n3477) );
  INV_X1 U4105 ( .A(n3476), .ZN(n3619) );
  NAND2_X1 U4106 ( .A1(n4930), .A2(n3392), .ZN(n3480) );
  NAND2_X1 U4107 ( .A1(n4901), .A2(n3249), .ZN(n3479) );
  NAND2_X1 U4108 ( .A1(n3480), .A2(n3479), .ZN(n3481) );
  XNOR2_X1 U4109 ( .A(n3481), .B(n3557), .ZN(n3487) );
  INV_X1 U4110 ( .A(n3487), .ZN(n3485) );
  NAND2_X1 U4111 ( .A1(n4930), .A2(n3548), .ZN(n3483) );
  NAND2_X1 U4112 ( .A1(n4901), .A2(n3392), .ZN(n3482) );
  NAND2_X1 U4113 ( .A1(n3483), .A2(n3482), .ZN(n3486) );
  INV_X1 U4114 ( .A(n3486), .ZN(n3484) );
  NAND2_X1 U4115 ( .A1(n3485), .A2(n3484), .ZN(n3649) );
  NAND2_X1 U4116 ( .A1(n4943), .A2(n3392), .ZN(n3489) );
  NAND2_X1 U4117 ( .A1(n4929), .A2(n3249), .ZN(n3488) );
  NAND2_X1 U4118 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  XNOR2_X1 U4119 ( .A(n3490), .B(n3557), .ZN(n3492) );
  NOR2_X1 U4120 ( .A1(n4297), .A2(n3347), .ZN(n3491) );
  AOI21_X1 U4121 ( .B1(n4943), .B2(n3548), .A(n3491), .ZN(n3493) );
  XNOR2_X1 U4122 ( .A(n3492), .B(n3493), .ZN(n4933) );
  INV_X1 U4123 ( .A(n3492), .ZN(n3494) );
  NAND2_X1 U4124 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  NAND2_X1 U4125 ( .A1(n4957), .A2(n3392), .ZN(n3497) );
  NAND2_X1 U4126 ( .A1(n4945), .A2(n3249), .ZN(n3496) );
  NAND2_X1 U4127 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  XNOR2_X1 U4128 ( .A(n3498), .B(n3557), .ZN(n3501) );
  NAND2_X1 U4129 ( .A1(n4957), .A2(n3548), .ZN(n3500) );
  NAND2_X1 U4130 ( .A1(n4945), .A2(n3392), .ZN(n3499) );
  NAND2_X1 U4131 ( .A1(n3500), .A2(n3499), .ZN(n3502) );
  NAND2_X1 U4132 ( .A1(n3501), .A2(n3502), .ZN(n4951) );
  INV_X1 U4133 ( .A(n3501), .ZN(n3504) );
  INV_X1 U4134 ( .A(n3502), .ZN(n3503) );
  NAND2_X1 U4135 ( .A1(n3504), .A2(n3503), .ZN(n4950) );
  NAND2_X1 U4136 ( .A1(n4971), .A2(n3392), .ZN(n3506) );
  NAND2_X1 U4137 ( .A1(n4958), .A2(n3249), .ZN(n3505) );
  NAND2_X1 U4138 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  XNOR2_X1 U4139 ( .A(n3507), .B(n3545), .ZN(n3515) );
  NOR2_X1 U4140 ( .A1(n4254), .A2(n3347), .ZN(n3508) );
  AOI21_X1 U4141 ( .B1(n4971), .B2(n3548), .A(n3508), .ZN(n3516) );
  NAND2_X1 U4142 ( .A1(n3515), .A2(n3516), .ZN(n4954) );
  AND2_X1 U4143 ( .A1(n4950), .A2(n4954), .ZN(n3509) );
  NAND2_X1 U4144 ( .A1(n4949), .A2(n3392), .ZN(n3511) );
  NAND2_X1 U4145 ( .A1(n4972), .A2(n3249), .ZN(n3510) );
  NAND2_X1 U4146 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  XNOR2_X1 U4147 ( .A(n3512), .B(n3557), .ZN(n3520) );
  NOR2_X1 U4148 ( .A1(n3513), .A2(n3347), .ZN(n3514) );
  AOI21_X1 U4149 ( .B1(n4949), .B2(n3548), .A(n3514), .ZN(n3521) );
  XNOR2_X1 U4150 ( .A(n3520), .B(n3521), .ZN(n4968) );
  INV_X1 U4151 ( .A(n3515), .ZN(n3518) );
  INV_X1 U4152 ( .A(n3516), .ZN(n3517) );
  NAND2_X1 U4153 ( .A1(n3518), .A2(n3517), .ZN(n4965) );
  AND2_X1 U4154 ( .A1(n4968), .A2(n4965), .ZN(n3519) );
  INV_X1 U4155 ( .A(n3520), .ZN(n3522) );
  NOR2_X1 U4156 ( .A1(n4222), .A2(n3347), .ZN(n3524) );
  AOI21_X1 U4157 ( .B1(n4963), .B2(n3548), .A(n3524), .ZN(n3528) );
  NAND2_X1 U4158 ( .A1(n4963), .A2(n3392), .ZN(n3526) );
  NAND2_X1 U4159 ( .A1(n3599), .A2(n3249), .ZN(n3525) );
  NAND2_X1 U4160 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  XNOR2_X1 U4161 ( .A(n3527), .B(n3557), .ZN(n3530) );
  XOR2_X1 U4162 ( .A(n3528), .B(n3530), .Z(n3597) );
  INV_X1 U4163 ( .A(n3528), .ZN(n3529) );
  NAND2_X1 U4164 ( .A1(n4197), .A2(n3392), .ZN(n3532) );
  NAND2_X1 U4165 ( .A1(n4183), .A2(n3249), .ZN(n3531) );
  NAND2_X1 U4166 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  XNOR2_X1 U4167 ( .A(n3533), .B(n3557), .ZN(n3605) );
  NAND2_X1 U4168 ( .A1(n4197), .A2(n3548), .ZN(n3535) );
  NAND2_X1 U4169 ( .A1(n4183), .A2(n3392), .ZN(n3534) );
  NAND2_X1 U4170 ( .A1(n3535), .A2(n3534), .ZN(n3604) );
  INV_X1 U4171 ( .A(n3604), .ZN(n3536) );
  AOI21_X1 U4172 ( .B1(n3606), .B2(n3630), .A(n3536), .ZN(n3538) );
  NAND3_X1 U4173 ( .A1(n3606), .A2(n3630), .A3(n3536), .ZN(n3537) );
  INV_X1 U4174 ( .A(n3539), .ZN(n3540) );
  NAND2_X1 U4175 ( .A1(n3541), .A2(n3540), .ZN(n3661) );
  NAND2_X1 U4176 ( .A1(n4180), .A2(n3542), .ZN(n3544) );
  NAND2_X1 U4177 ( .A1(n4151), .A2(n3249), .ZN(n3543) );
  NAND2_X1 U4178 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  XNOR2_X1 U4179 ( .A(n3546), .B(n3545), .ZN(n3550) );
  NOR2_X1 U4180 ( .A1(n4160), .A2(n3347), .ZN(n3547) );
  AOI21_X1 U4181 ( .B1(n4180), .B2(n3548), .A(n3547), .ZN(n3549) );
  NAND2_X1 U4182 ( .A1(n3661), .A2(n2531), .ZN(n3551) );
  NAND2_X1 U4183 ( .A1(n3550), .A2(n3549), .ZN(n3659) );
  OAI22_X1 U4184 ( .A1(n4120), .A2(n3347), .B1(n4146), .B2(n3555), .ZN(n3552)
         );
  XNOR2_X1 U4185 ( .A(n3552), .B(n3557), .ZN(n3554) );
  OAI22_X1 U4186 ( .A1(n4120), .A2(n3556), .B1(n4146), .B2(n3347), .ZN(n3553)
         );
  XNOR2_X1 U4187 ( .A(n3554), .B(n3553), .ZN(n3577) );
  OAI22_X1 U4188 ( .A1(n4140), .A2(n3347), .B1(n3555), .B2(n4125), .ZN(n3560)
         );
  OAI22_X1 U4189 ( .A1(n4140), .A2(n3556), .B1(n3347), .B2(n4125), .ZN(n3558)
         );
  XNOR2_X1 U4190 ( .A(n3558), .B(n3557), .ZN(n3559) );
  XOR2_X1 U4191 ( .A(n3560), .B(n3559), .Z(n3561) );
  INV_X1 U4192 ( .A(n4128), .ZN(n3565) );
  AOI22_X1 U4193 ( .A1(n4970), .A2(n4163), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3564) );
  AOI22_X1 U4194 ( .A1(n4964), .A2(n4124), .B1(n4973), .B2(n3562), .ZN(n3563)
         );
  OAI211_X1 U4195 ( .C1(n4979), .C2(n3565), .A(n3564), .B(n3563), .ZN(n3566)
         );
  INV_X1 U4196 ( .A(n3566), .ZN(n3567) );
  NAND3_X1 U4197 ( .A1(n3568), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3569) );
  INV_X1 U4198 ( .A(DATAI_31_), .ZN(n3668) );
  OAI22_X1 U4199 ( .A1(n2553), .A2(n3569), .B1(STATE_REG_SCAN_IN), .B2(n3668), 
        .ZN(U3321) );
  OAI211_X1 U4200 ( .C1(n3572), .C2(n3571), .A(n3570), .B(n4974), .ZN(n3576)
         );
  INV_X1 U4201 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4007) );
  NOR2_X1 U4202 ( .A1(STATE_REG_SCAN_IN), .A2(n4007), .ZN(n4517) );
  AOI21_X1 U4203 ( .B1(n4964), .B2(n4729), .A(n4517), .ZN(n3575) );
  AOI22_X1 U4204 ( .A1(n4970), .A2(n3832), .B1(n4973), .B2(n4723), .ZN(n3574)
         );
  OR2_X1 U4205 ( .A1(n4979), .A2(n4740), .ZN(n3573) );
  NAND4_X1 U4206 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(U3210)
         );
  XNOR2_X1 U4207 ( .A(n3578), .B(n3577), .ZN(n3584) );
  INV_X1 U4208 ( .A(n4141), .ZN(n3581) );
  AOI22_X1 U4209 ( .A1(n3828), .A2(n4964), .B1(n4137), .B2(n4973), .ZN(n3580)
         );
  AOI22_X1 U4210 ( .A1(n4970), .A2(n4180), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3579) );
  OAI211_X1 U4211 ( .C1(n4979), .C2(n3581), .A(n3580), .B(n3579), .ZN(n3582)
         );
  INV_X1 U4212 ( .A(n3582), .ZN(n3583) );
  OAI21_X1 U4213 ( .B1(n3584), .B2(n4846), .A(n3583), .ZN(U3211) );
  NAND2_X1 U4214 ( .A1(n2325), .A2(n3585), .ZN(n3586) );
  XNOR2_X1 U4215 ( .A(n3587), .B(n3586), .ZN(n3593) );
  INV_X1 U4216 ( .A(n4800), .ZN(n3591) );
  NOR2_X1 U4217 ( .A1(n3907), .A2(STATE_REG_SCAN_IN), .ZN(n4057) );
  AOI21_X1 U4218 ( .B1(n4970), .B2(n4407), .A(n4057), .ZN(n3590) );
  AOI22_X1 U4219 ( .A1(n4964), .A2(n4859), .B1(n4973), .B2(n3588), .ZN(n3589)
         );
  OAI211_X1 U4220 ( .C1(n4979), .C2(n3591), .A(n3590), .B(n3589), .ZN(n3592)
         );
  AOI21_X1 U4221 ( .B1(n3593), .B2(n4974), .A(n3592), .ZN(n3594) );
  INV_X1 U4222 ( .A(n3594), .ZN(U3212) );
  AOI211_X1 U4223 ( .C1(n3597), .C2(n3596), .A(n4846), .B(n3595), .ZN(n3603)
         );
  INV_X1 U4224 ( .A(n3598), .ZN(n4228) );
  AOI22_X1 U4225 ( .A1(n4970), .A2(n4949), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3601) );
  AOI22_X1 U4226 ( .A1(n4964), .A2(n4225), .B1(n4973), .B2(n3599), .ZN(n3600)
         );
  OAI211_X1 U4227 ( .C1(n4979), .C2(n4228), .A(n3601), .B(n3600), .ZN(n3602)
         );
  OR2_X1 U4228 ( .A1(n3603), .A2(n3602), .ZN(U3213) );
  NOR2_X1 U4229 ( .A1(n3605), .A2(n3604), .ZN(n3608) );
  INV_X1 U4230 ( .A(n3608), .ZN(n3611) );
  OR2_X1 U4231 ( .A1(n3607), .A2(n3606), .ZN(n3629) );
  NAND2_X1 U4232 ( .A1(n3607), .A2(n3606), .ZN(n3628) );
  OAI21_X1 U4233 ( .B1(n2301), .B2(n3608), .A(n3628), .ZN(n3609) );
  AOI21_X1 U4234 ( .B1(n3630), .B2(n3629), .A(n3609), .ZN(n3610) );
  AOI21_X1 U4235 ( .B1(n3661), .B2(n3611), .A(n3610), .ZN(n3618) );
  INV_X1 U4236 ( .A(n4979), .ZN(n3616) );
  OAI22_X1 U4237 ( .A1(n4178), .A2(n3612), .B1(STATE_REG_SCAN_IN), .B2(n3946), 
        .ZN(n3615) );
  OAI22_X1 U4238 ( .A1(n4808), .A2(n4177), .B1(n3613), .B2(n4934), .ZN(n3614)
         );
  AOI211_X1 U4239 ( .C1(n4186), .C2(n3616), .A(n3615), .B(n3614), .ZN(n3617)
         );
  OAI21_X1 U4240 ( .B1(n3618), .B2(n4846), .A(n3617), .ZN(U3222) );
  XNOR2_X1 U4241 ( .A(n3620), .B(n3619), .ZN(n3621) );
  XNOR2_X1 U4242 ( .A(n3622), .B(n3621), .ZN(n3626) );
  INV_X1 U4243 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3919) );
  NOR2_X1 U4244 ( .A1(STATE_REG_SCAN_IN), .A2(n3919), .ZN(n4087) );
  AOI21_X1 U4245 ( .B1(n4970), .B2(n4830), .A(n4087), .ZN(n3624) );
  AOI22_X1 U4246 ( .A1(n4964), .A2(n4930), .B1(n4973), .B2(n4391), .ZN(n3623)
         );
  OAI211_X1 U4247 ( .C1(n4979), .C2(n4883), .A(n3624), .B(n3623), .ZN(n3625)
         );
  AOI21_X1 U4248 ( .B1(n3626), .B2(n4974), .A(n3625), .ZN(n3627) );
  INV_X1 U4249 ( .A(n3627), .ZN(U3225) );
  NAND2_X1 U4250 ( .A1(n3629), .A2(n3628), .ZN(n3631) );
  XNOR2_X1 U4251 ( .A(n3631), .B(n3630), .ZN(n3638) );
  INV_X1 U4252 ( .A(n3632), .ZN(n4205) );
  AOI22_X1 U4253 ( .A1(n4970), .A2(n4963), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3635) );
  AOI22_X1 U4254 ( .A1(n4964), .A2(n4197), .B1(n4973), .B2(n3633), .ZN(n3634)
         );
  OAI211_X1 U4255 ( .C1(n4979), .C2(n4205), .A(n3635), .B(n3634), .ZN(n3636)
         );
  INV_X1 U4256 ( .A(n3636), .ZN(n3637) );
  OAI21_X1 U4257 ( .B1(n3638), .B2(n4846), .A(n3637), .ZN(U3226) );
  XNOR2_X1 U4258 ( .A(n3640), .B(n3639), .ZN(n3641) );
  XNOR2_X1 U4259 ( .A(n3642), .B(n3641), .ZN(n3647) );
  INV_X1 U4260 ( .A(n3643), .ZN(n4321) );
  NOR2_X1 U4261 ( .A1(STATE_REG_SCAN_IN), .A2(n2725), .ZN(n4580) );
  AOI21_X1 U4262 ( .B1(n4964), .B2(n4823), .A(n4580), .ZN(n3645) );
  AOI22_X1 U4263 ( .A1(n4970), .A2(n4313), .B1(n4973), .B2(n4320), .ZN(n3644)
         );
  OAI211_X1 U4264 ( .C1(n4979), .C2(n4321), .A(n3645), .B(n3644), .ZN(n3646)
         );
  AOI21_X1 U4265 ( .B1(n3647), .B2(n4974), .A(n3646), .ZN(n3648) );
  INV_X1 U4266 ( .A(n3648), .ZN(U3231) );
  NAND2_X1 U4267 ( .A1(n2320), .A2(n3649), .ZN(n3650) );
  XNOR2_X1 U4268 ( .A(n3651), .B(n3650), .ZN(n3657) );
  INV_X1 U4269 ( .A(n4921), .ZN(n3655) );
  NOR2_X1 U4270 ( .A1(STATE_REG_SCAN_IN), .A2(n3652), .ZN(n4096) );
  AOI21_X1 U4271 ( .B1(n4970), .B2(n4904), .A(n4096), .ZN(n3654) );
  AOI22_X1 U4272 ( .A1(n4964), .A2(n4943), .B1(n4973), .B2(n4901), .ZN(n3653)
         );
  OAI211_X1 U4273 ( .C1(n4979), .C2(n3655), .A(n3654), .B(n3653), .ZN(n3656)
         );
  AOI21_X1 U4274 ( .B1(n3657), .B2(n4974), .A(n3656), .ZN(n3658) );
  INV_X1 U4275 ( .A(n3658), .ZN(U3235) );
  NAND2_X1 U4276 ( .A1(n2531), .A2(n3659), .ZN(n3660) );
  XNOR2_X1 U4277 ( .A(n3661), .B(n3660), .ZN(n3667) );
  INV_X1 U4278 ( .A(n3662), .ZN(n4166) );
  AOI22_X1 U4279 ( .A1(n4163), .A2(n4964), .B1(n4151), .B2(n4973), .ZN(n3664)
         );
  AOI22_X1 U4280 ( .A1(n4970), .A2(n4197), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3663) );
  OAI211_X1 U4281 ( .C1(n4979), .C2(n4166), .A(n3664), .B(n3663), .ZN(n3665)
         );
  INV_X1 U4282 ( .A(n3665), .ZN(n3666) );
  OAI21_X1 U4283 ( .B1(n3667), .B2(n4846), .A(n3666), .ZN(U3237) );
  NOR2_X1 U4284 ( .A1(n3669), .A2(n3668), .ZN(n4107) );
  NAND2_X1 U4285 ( .A1(n4106), .A2(n4107), .ZN(n3672) );
  NAND2_X1 U4286 ( .A1(n3670), .A2(DATAI_30_), .ZN(n4340) );
  NAND2_X1 U4287 ( .A1(n3827), .A2(n4340), .ZN(n3671) );
  NAND2_X1 U4288 ( .A1(n3672), .A2(n3671), .ZN(n3773) );
  NAND2_X1 U4289 ( .A1(n3677), .A2(n3673), .ZN(n3711) );
  AND2_X1 U4290 ( .A1(n3675), .A2(n3674), .ZN(n3740) );
  INV_X1 U4291 ( .A(n3740), .ZN(n3676) );
  NAND2_X1 U4292 ( .A1(n3677), .A2(n3676), .ZN(n3715) );
  OAI21_X1 U4293 ( .B1(n4406), .B2(n3711), .A(n3715), .ZN(n3679) );
  INV_X1 U4294 ( .A(n3747), .ZN(n3678) );
  AOI211_X1 U4295 ( .C1(n3702), .C2(n3679), .A(n3678), .B(n3744), .ZN(n3681)
         );
  INV_X1 U4296 ( .A(n3751), .ZN(n3680) );
  AOI211_X1 U4297 ( .C1(n3748), .C2(n3681), .A(n3680), .B(n3753), .ZN(n3684)
         );
  INV_X1 U4298 ( .A(n3682), .ZN(n3683) );
  OAI21_X1 U4299 ( .B1(n3684), .B2(n3683), .A(n3755), .ZN(n3688) );
  OR2_X1 U4300 ( .A1(n4106), .A2(n4107), .ZN(n3767) );
  OAI21_X1 U4301 ( .B1(n4340), .B2(n3827), .A(n3767), .ZN(n3778) );
  INV_X1 U4302 ( .A(n3778), .ZN(n3685) );
  OAI21_X1 U4303 ( .B1(n4124), .B2(n3689), .A(n3685), .ZN(n3692) );
  NAND2_X1 U4304 ( .A1(n3687), .A2(n3686), .ZN(n3693) );
  AOI211_X1 U4305 ( .C1(n3763), .C2(n3688), .A(n3692), .B(n3693), .ZN(n3696)
         );
  NAND2_X1 U4306 ( .A1(n4124), .A2(n3689), .ZN(n3690) );
  AND2_X1 U4307 ( .A1(n3691), .A2(n3690), .ZN(n3758) );
  AOI21_X1 U4308 ( .B1(n3693), .B2(n3758), .A(n3692), .ZN(n3766) );
  NAND3_X1 U4309 ( .A1(n4142), .A2(n3758), .A3(n3694), .ZN(n3695) );
  AOI22_X1 U4310 ( .A1(n3701), .A2(n3696), .B1(n3766), .B2(n3695), .ZN(n3697)
         );
  AOI21_X1 U4311 ( .B1(n4339), .B2(n4106), .A(n3697), .ZN(n3698) );
  AOI21_X1 U4312 ( .B1(n4107), .B2(n3773), .A(n3698), .ZN(n3699) );
  XNOR2_X1 U4313 ( .A(n3699), .B(n4732), .ZN(n3821) );
  INV_X1 U4314 ( .A(n3700), .ZN(n3820) );
  INV_X1 U4315 ( .A(n3701), .ZN(n3764) );
  INV_X1 U4316 ( .A(n3702), .ZN(n3750) );
  NAND3_X1 U4317 ( .A1(n3705), .A2(n3704), .A3(n3703), .ZN(n3735) );
  NOR3_X1 U4318 ( .A1(n3735), .A2(n2402), .A3(n3706), .ZN(n3710) );
  AND2_X1 U4319 ( .A1(n3709), .A2(n3708), .ZN(n3741) );
  OAI21_X1 U4320 ( .B1(n3710), .B2(n2411), .A(n3741), .ZN(n3714) );
  INV_X1 U4321 ( .A(n3711), .ZN(n3712) );
  NAND3_X1 U4322 ( .A1(n3714), .A2(n3713), .A3(n3712), .ZN(n3716) );
  NAND2_X1 U4323 ( .A1(n3716), .A2(n3715), .ZN(n3746) );
  INV_X1 U4324 ( .A(n3798), .ZN(n4660) );
  NAND2_X1 U4325 ( .A1(n4663), .A2(n4674), .ZN(n3797) );
  OAI211_X1 U4326 ( .C1(n4660), .C2(n3718), .A(n3797), .B(n3717), .ZN(n3721)
         );
  NAND3_X1 U4327 ( .A1(n3721), .A2(n3720), .A3(n3719), .ZN(n3724) );
  NAND3_X1 U4328 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3730) );
  NAND3_X1 U4329 ( .A1(n3727), .A2(n3726), .A3(n3725), .ZN(n3728) );
  AOI21_X1 U4330 ( .B1(n3730), .B2(n3729), .A(n3728), .ZN(n3734) );
  INV_X1 U4331 ( .A(n3731), .ZN(n3733) );
  NOR3_X1 U4332 ( .A1(n3734), .A2(n3733), .A3(n3732), .ZN(n3736) );
  NOR2_X1 U4333 ( .A1(n3736), .A2(n3735), .ZN(n3743) );
  AOI21_X1 U4334 ( .B1(n3739), .B2(n3738), .A(n3737), .ZN(n3742) );
  OAI211_X1 U4335 ( .C1(n3743), .C2(n3742), .A(n3741), .B(n3740), .ZN(n3745)
         );
  AOI21_X1 U4336 ( .B1(n3746), .B2(n3745), .A(n3744), .ZN(n3749) );
  OAI211_X1 U4337 ( .C1(n3750), .C2(n3749), .A(n3748), .B(n3747), .ZN(n3752)
         );
  AOI21_X1 U4338 ( .B1(n3752), .B2(n3751), .A(n4218), .ZN(n3754) );
  NOR2_X1 U4339 ( .A1(n3754), .A2(n3753), .ZN(n3757) );
  OAI21_X1 U4340 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n3762) );
  NOR2_X1 U4341 ( .A1(n4120), .A2(n4137), .ZN(n3760) );
  INV_X1 U4342 ( .A(n3758), .ZN(n3759) );
  NOR4_X1 U4343 ( .A1(n3760), .A2(n3772), .A3(n3759), .A4(n3773), .ZN(n3761)
         );
  OAI221_X1 U4344 ( .B1(n3764), .B2(n3763), .C1(n3764), .C2(n3762), .A(n3761), 
        .ZN(n3765) );
  INV_X1 U4345 ( .A(n3765), .ZN(n3769) );
  AOI21_X1 U4346 ( .B1(n3773), .B2(n3767), .A(n3766), .ZN(n3768) );
  OAI21_X1 U4347 ( .B1(n3769), .B2(n3768), .A(n2841), .ZN(n3814) );
  INV_X1 U4348 ( .A(n3814), .ZN(n3811) );
  INV_X1 U4349 ( .A(n4218), .ZN(n3770) );
  NAND2_X1 U4350 ( .A1(n3770), .A2(n4217), .ZN(n4257) );
  OR2_X1 U4351 ( .A1(n3772), .A2(n3771), .ZN(n4159) );
  NOR2_X1 U4352 ( .A1(n4257), .A2(n4159), .ZN(n3777) );
  INV_X1 U4353 ( .A(n3773), .ZN(n3776) );
  NOR4_X1 U4354 ( .A1(n4865), .A2(n4827), .A3(n4405), .A4(n3774), .ZN(n3775)
         );
  NAND4_X1 U4355 ( .A1(n3777), .A2(n4239), .A3(n3776), .A4(n3775), .ZN(n3788)
         );
  AND2_X1 U4356 ( .A1(n4401), .A2(n4400), .ZN(n4312) );
  NOR2_X1 U4357 ( .A1(n4312), .A2(n3778), .ZN(n3786) );
  NAND2_X1 U4358 ( .A1(n4310), .A2(n4308), .ZN(n4421) );
  NOR2_X1 U4359 ( .A1(n4421), .A2(n3779), .ZN(n3785) );
  NOR2_X1 U4360 ( .A1(n3781), .A2(n3780), .ZN(n3784) );
  NOR2_X1 U4361 ( .A1(n4734), .A2(n3782), .ZN(n3783) );
  NAND4_X1 U4362 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3787)
         );
  NOR2_X1 U4363 ( .A1(n3788), .A2(n3787), .ZN(n3809) );
  INV_X1 U4364 ( .A(n3789), .ZN(n3790) );
  NOR2_X1 U4365 ( .A1(n4191), .A2(n3790), .ZN(n4220) );
  INV_X1 U4366 ( .A(n4122), .ZN(n3791) );
  NOR2_X1 U4367 ( .A1(n4286), .A2(n4288), .ZN(n4389) );
  NAND4_X1 U4368 ( .A1(n4220), .A2(n3791), .A3(n4389), .A4(n4899), .ZN(n3795)
         );
  XNOR2_X1 U4369 ( .A(n4957), .B(n3792), .ZN(n4269) );
  INV_X1 U4370 ( .A(n4269), .ZN(n4265) );
  XNOR2_X1 U4371 ( .A(n4197), .B(n4183), .ZN(n4175) );
  NAND2_X1 U4372 ( .A1(n4265), .A2(n4175), .ZN(n3793) );
  NOR3_X1 U4373 ( .A1(n3795), .A2(n3794), .A3(n3793), .ZN(n3808) );
  NOR2_X1 U4374 ( .A1(n3796), .A2(n4172), .ZN(n4200) );
  INV_X1 U4375 ( .A(n4668), .ZN(n4661) );
  AND2_X1 U4376 ( .A1(n3798), .A2(n3797), .ZN(n4647) );
  NAND4_X1 U4377 ( .A1(n4200), .A2(n4661), .A3(n4647), .A4(n4292), .ZN(n3806)
         );
  NAND4_X1 U4378 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  NOR2_X1 U4379 ( .A1(n3806), .A2(n3805), .ZN(n3807) );
  NAND4_X1 U4380 ( .A1(n3809), .A2(n3808), .A3(n4142), .A4(n3807), .ZN(n3816)
         );
  AOI21_X1 U4381 ( .B1(n3816), .B2(n3812), .A(n2841), .ZN(n3810) );
  NOR2_X1 U4382 ( .A1(n3811), .A2(n3810), .ZN(n3818) );
  NAND2_X1 U4383 ( .A1(n3813), .A2(n3812), .ZN(n3815) );
  OAI21_X1 U4384 ( .B1(n3816), .B2(n3815), .A(n3814), .ZN(n3817) );
  MUX2_X1 U4385 ( .A(n3818), .B(n3817), .S(n4732), .Z(n3819) );
  AOI21_X1 U4386 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3826) );
  NAND2_X1 U4387 ( .A1(n4600), .A2(n3822), .ZN(n3823) );
  OAI211_X1 U4388 ( .C1(n3824), .C2(n4489), .A(n3823), .B(B_REG_SCAN_IN), .ZN(
        n3825) );
  OAI21_X1 U4389 ( .B1(n3826), .B2(n4489), .A(n3825), .ZN(U3239) );
  MUX2_X1 U4390 ( .A(n3827), .B(DATAO_REG_30__SCAN_IN), .S(n3838), .Z(U3580)
         );
  MUX2_X1 U4391 ( .A(n4124), .B(DATAO_REG_29__SCAN_IN), .S(n3838), .Z(U3579)
         );
  MUX2_X1 U4392 ( .A(DATAO_REG_28__SCAN_IN), .B(n3828), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4393 ( .A(DATAO_REG_27__SCAN_IN), .B(n4163), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4394 ( .A(n4180), .B(DATAO_REG_26__SCAN_IN), .S(n3838), .Z(U3576)
         );
  MUX2_X1 U4395 ( .A(n4197), .B(DATAO_REG_25__SCAN_IN), .S(n3838), .Z(U3575)
         );
  MUX2_X1 U4396 ( .A(n4225), .B(DATAO_REG_24__SCAN_IN), .S(n3838), .Z(U3574)
         );
  MUX2_X1 U4397 ( .A(n4963), .B(DATAO_REG_23__SCAN_IN), .S(n3838), .Z(U3573)
         );
  MUX2_X1 U4398 ( .A(n4949), .B(DATAO_REG_22__SCAN_IN), .S(n3838), .Z(U3572)
         );
  MUX2_X1 U4399 ( .A(n4971), .B(DATAO_REG_21__SCAN_IN), .S(n3838), .Z(U3571)
         );
  MUX2_X1 U4400 ( .A(n4957), .B(DATAO_REG_20__SCAN_IN), .S(n3838), .Z(U3570)
         );
  MUX2_X1 U4401 ( .A(n4943), .B(DATAO_REG_19__SCAN_IN), .S(n3838), .Z(U3569)
         );
  MUX2_X1 U4402 ( .A(n4930), .B(DATAO_REG_18__SCAN_IN), .S(n3838), .Z(U3568)
         );
  MUX2_X1 U4403 ( .A(n4904), .B(DATAO_REG_17__SCAN_IN), .S(n3838), .Z(U3567)
         );
  MUX2_X1 U4404 ( .A(n4830), .B(DATAO_REG_16__SCAN_IN), .S(n3838), .Z(U3566)
         );
  MUX2_X1 U4405 ( .A(n4859), .B(DATAO_REG_15__SCAN_IN), .S(n3838), .Z(U3565)
         );
  MUX2_X1 U4406 ( .A(n4823), .B(DATAO_REG_14__SCAN_IN), .S(n3838), .Z(U3564)
         );
  MUX2_X1 U4407 ( .A(n4407), .B(DATAO_REG_13__SCAN_IN), .S(n3838), .Z(U3563)
         );
  MUX2_X1 U4408 ( .A(n4313), .B(DATAO_REG_12__SCAN_IN), .S(n3838), .Z(U3562)
         );
  MUX2_X1 U4409 ( .A(n4424), .B(DATAO_REG_11__SCAN_IN), .S(n3838), .Z(U3561)
         );
  MUX2_X1 U4410 ( .A(n3829), .B(DATAO_REG_10__SCAN_IN), .S(n3838), .Z(U3560)
         );
  MUX2_X1 U4411 ( .A(n3830), .B(DATAO_REG_9__SCAN_IN), .S(n3838), .Z(U3559) );
  MUX2_X1 U4412 ( .A(n4729), .B(DATAO_REG_8__SCAN_IN), .S(n3838), .Z(U3558) );
  MUX2_X1 U4413 ( .A(n3831), .B(DATAO_REG_7__SCAN_IN), .S(n3838), .Z(U3557) );
  MUX2_X1 U4414 ( .A(n3832), .B(DATAO_REG_6__SCAN_IN), .S(n3838), .Z(U3556) );
  MUX2_X1 U4415 ( .A(n3833), .B(DATAO_REG_5__SCAN_IN), .S(n3838), .Z(U3555) );
  MUX2_X1 U4416 ( .A(n3834), .B(DATAO_REG_4__SCAN_IN), .S(n3838), .Z(U3554) );
  MUX2_X1 U4417 ( .A(n3835), .B(DATAO_REG_3__SCAN_IN), .S(n3838), .Z(U3553) );
  MUX2_X1 U4418 ( .A(n3836), .B(DATAO_REG_2__SCAN_IN), .S(n3838), .Z(U3552) );
  MUX2_X1 U4419 ( .A(n3837), .B(DATAO_REG_1__SCAN_IN), .S(n3838), .Z(U3551) );
  MUX2_X1 U4420 ( .A(n4663), .B(DATAO_REG_0__SCAN_IN), .S(n3838), .Z(U3550) );
  NOR2_X1 U4421 ( .A1(STATE_REG_SCAN_IN), .A2(n3076), .ZN(n3840) );
  NOR2_X1 U4422 ( .A1(n4643), .A2(n3841), .ZN(n3839) );
  AOI211_X1 U4423 ( .C1(n4629), .C2(ADDR_REG_1__SCAN_IN), .A(n3840), .B(n3839), 
        .ZN(n3851) );
  NOR2_X1 U4424 ( .A1(n4609), .A2(n4648), .ZN(n3845) );
  MUX2_X1 U4425 ( .A(n3842), .B(REG1_REG_1__SCAN_IN), .S(n3841), .Z(n3844) );
  INV_X1 U4426 ( .A(n4622), .ZN(n3843) );
  OAI211_X1 U4427 ( .C1(n3845), .C2(n3844), .A(n4630), .B(n3843), .ZN(n3850)
         );
  OAI211_X1 U4428 ( .C1(n3848), .C2(n3847), .A(n4611), .B(n3846), .ZN(n3849)
         );
  NAND3_X1 U4429 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(U3241) );
  XOR2_X1 U4430 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_127), .Z(n4046) );
  INV_X1 U4431 ( .A(IR_REG_6__SCAN_IN), .ZN(n3853) );
  OAI22_X1 U4432 ( .A1(n3853), .A2(keyinput_125), .B1(keyinput_124), .B2(
        IR_REG_5__SCAN_IN), .ZN(n3852) );
  AOI221_X1 U4433 ( .B1(n3853), .B2(keyinput_125), .C1(IR_REG_5__SCAN_IN), 
        .C2(keyinput_124), .A(n3852), .ZN(n3941) );
  INV_X1 U4434 ( .A(keyinput_123), .ZN(n3939) );
  INV_X1 U4435 ( .A(keyinput_122), .ZN(n3937) );
  OAI22_X1 U4436 ( .A1(n2725), .A2(keyinput_118), .B1(keyinput_121), .B2(
        IR_REG_2__SCAN_IN), .ZN(n3854) );
  AOI221_X1 U4437 ( .B1(n2725), .B2(keyinput_118), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_121), .A(n3854), .ZN(n3935) );
  OAI22_X1 U4438 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_119), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput_120), .ZN(n3855) );
  AOI221_X1 U4439 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_119), .C1(
        keyinput_120), .C2(IR_REG_1__SCAN_IN), .A(n3855), .ZN(n3934) );
  OAI22_X1 U4440 ( .A1(n4007), .A2(keyinput_97), .B1(REG3_REG_27__SCAN_IN), 
        .B2(keyinput_98), .ZN(n3856) );
  AOI221_X1 U4441 ( .B1(n4007), .B2(keyinput_97), .C1(keyinput_98), .C2(
        REG3_REG_27__SCAN_IN), .A(n3856), .ZN(n3912) );
  INV_X1 U4442 ( .A(keyinput_96), .ZN(n3905) );
  INV_X1 U4443 ( .A(keyinput_95), .ZN(n3903) );
  INV_X1 U4444 ( .A(keyinput_94), .ZN(n3901) );
  INV_X1 U4445 ( .A(DATAI_2_), .ZN(n3899) );
  INV_X1 U4446 ( .A(DATAI_3_), .ZN(n4695) );
  OAI22_X1 U4447 ( .A1(n4695), .A2(keyinput_92), .B1(DATAI_4_), .B2(
        keyinput_91), .ZN(n3857) );
  AOI221_X1 U4448 ( .B1(n4695), .B2(keyinput_92), .C1(keyinput_91), .C2(
        DATAI_4_), .A(n3857), .ZN(n3897) );
  INV_X1 U4449 ( .A(DATAI_5_), .ZN(n3995) );
  INV_X1 U4450 ( .A(keyinput_90), .ZN(n3895) );
  INV_X1 U4451 ( .A(DATAI_7_), .ZN(n4719) );
  AOI22_X1 U4452 ( .A1(DATAI_8_), .A2(keyinput_87), .B1(n4719), .B2(
        keyinput_88), .ZN(n3858) );
  OAI221_X1 U4453 ( .B1(DATAI_8_), .B2(keyinput_87), .C1(n4719), .C2(
        keyinput_88), .A(n3858), .ZN(n3893) );
  AOI22_X1 U4454 ( .A1(n3861), .A2(keyinput_74), .B1(n3860), .B2(keyinput_73), 
        .ZN(n3859) );
  OAI221_X1 U4455 ( .B1(n3861), .B2(keyinput_74), .C1(n3860), .C2(keyinput_73), 
        .A(n3859), .ZN(n3875) );
  INV_X1 U4456 ( .A(DATAI_25_), .ZN(n3968) );
  OAI22_X1 U4457 ( .A1(n3968), .A2(keyinput_70), .B1(keyinput_72), .B2(
        DATAI_23_), .ZN(n3862) );
  AOI221_X1 U4458 ( .B1(n3968), .B2(keyinput_70), .C1(DATAI_23_), .C2(
        keyinput_72), .A(n3862), .ZN(n3872) );
  INV_X1 U4459 ( .A(keyinput_69), .ZN(n3870) );
  OAI22_X1 U4460 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        DATAI_31_), .ZN(n3863) );
  AOI221_X1 U4461 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n3863), .ZN(n3867) );
  INV_X1 U4462 ( .A(DATAI_27_), .ZN(n3960) );
  AOI22_X1 U4463 ( .A1(n3960), .A2(keyinput_68), .B1(n3865), .B2(keyinput_67), 
        .ZN(n3864) );
  OAI221_X1 U4464 ( .B1(n3960), .B2(keyinput_68), .C1(n3865), .C2(keyinput_67), 
        .A(n3864), .ZN(n3866) );
  AOI211_X1 U4465 ( .C1(keyinput_66), .C2(DATAI_29_), .A(n3867), .B(n3866), 
        .ZN(n3868) );
  OAI21_X1 U4466 ( .B1(keyinput_66), .B2(DATAI_29_), .A(n3868), .ZN(n3869) );
  OAI221_X1 U4467 ( .B1(DATAI_26_), .B2(n3870), .C1(n3957), .C2(keyinput_69), 
        .A(n3869), .ZN(n3871) );
  OAI211_X1 U4468 ( .C1(DATAI_24_), .C2(keyinput_71), .A(n3872), .B(n3871), 
        .ZN(n3873) );
  AOI21_X1 U4469 ( .B1(DATAI_24_), .B2(keyinput_71), .A(n3873), .ZN(n3874) );
  OAI22_X1 U4470 ( .A1(keyinput_75), .A2(n3976), .B1(n3875), .B2(n3874), .ZN(
        n3876) );
  AOI21_X1 U4471 ( .B1(keyinput_75), .B2(n3976), .A(n3876), .ZN(n3883) );
  INV_X1 U4472 ( .A(DATAI_19_), .ZN(n3977) );
  XOR2_X1 U4473 ( .A(n3977), .B(keyinput_76), .Z(n3882) );
  INV_X1 U4474 ( .A(DATAI_15_), .ZN(n3979) );
  AOI22_X1 U4475 ( .A1(n3979), .A2(keyinput_80), .B1(n3878), .B2(keyinput_77), 
        .ZN(n3877) );
  OAI221_X1 U4476 ( .B1(n3979), .B2(keyinput_80), .C1(n3878), .C2(keyinput_77), 
        .A(n3877), .ZN(n3881) );
  AOI22_X1 U4477 ( .A1(DATAI_16_), .A2(keyinput_79), .B1(DATAI_17_), .B2(
        keyinput_78), .ZN(n3879) );
  OAI221_X1 U4478 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(DATAI_17_), .C2(
        keyinput_78), .A(n3879), .ZN(n3880) );
  AOI211_X1 U4479 ( .C1(n3883), .C2(n3882), .A(n3881), .B(n3880), .ZN(n3890)
         );
  INV_X1 U4480 ( .A(DATAI_11_), .ZN(n4767) );
  OAI22_X1 U4481 ( .A1(n4767), .A2(keyinput_84), .B1(DATAI_12_), .B2(
        keyinput_83), .ZN(n3884) );
  AOI221_X1 U4482 ( .B1(n4767), .B2(keyinput_84), .C1(keyinput_83), .C2(
        DATAI_12_), .A(n3884), .ZN(n3889) );
  AOI22_X1 U4483 ( .A1(DATAI_13_), .A2(keyinput_82), .B1(DATAI_14_), .B2(
        keyinput_81), .ZN(n3885) );
  OAI221_X1 U4484 ( .B1(DATAI_13_), .B2(keyinput_82), .C1(DATAI_14_), .C2(
        keyinput_81), .A(n3885), .ZN(n3888) );
  AOI22_X1 U4485 ( .A1(DATAI_9_), .A2(keyinput_86), .B1(DATAI_10_), .B2(
        keyinput_85), .ZN(n3886) );
  OAI221_X1 U4486 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(DATAI_10_), .C2(
        keyinput_85), .A(n3886), .ZN(n3887) );
  AOI221_X1 U4487 ( .B1(n3890), .B2(n3889), .C1(n3888), .C2(n3889), .A(n3887), 
        .ZN(n3892) );
  NAND2_X1 U4488 ( .A1(DATAI_6_), .A2(keyinput_89), .ZN(n3891) );
  OAI221_X1 U4489 ( .B1(n3893), .B2(n3892), .C1(DATAI_6_), .C2(keyinput_89), 
        .A(n3891), .ZN(n3894) );
  OAI221_X1 U4490 ( .B1(DATAI_5_), .B2(keyinput_90), .C1(n3995), .C2(n3895), 
        .A(n3894), .ZN(n3896) );
  AOI22_X1 U4491 ( .A1(keyinput_93), .A2(n3899), .B1(n3897), .B2(n3896), .ZN(
        n3898) );
  OAI21_X1 U4492 ( .B1(n3899), .B2(keyinput_93), .A(n3898), .ZN(n3900) );
  OAI221_X1 U4493 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(n2603), .C2(n3901), 
        .A(n3900), .ZN(n3902) );
  OAI221_X1 U4494 ( .B1(DATAI_0_), .B2(keyinput_95), .C1(n4599), .C2(n3903), 
        .A(n3902), .ZN(n3904) );
  OAI221_X1 U4495 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_96), .C1(U3149), .C2(
        n3905), .A(n3904), .ZN(n3911) );
  AOI22_X1 U4496 ( .A1(n3907), .A2(keyinput_99), .B1(n4696), .B2(keyinput_102), 
        .ZN(n3906) );
  OAI221_X1 U4497 ( .B1(n3907), .B2(keyinput_99), .C1(n4696), .C2(keyinput_102), .A(n3906), .ZN(n3910) );
  AOI22_X1 U4498 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_100), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_101), .ZN(n3908) );
  OAI221_X1 U4499 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_100), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_101), .A(n3908), .ZN(n3909) );
  AOI211_X1 U4500 ( .C1(n3912), .C2(n3911), .A(n3910), .B(n3909), .ZN(n3932)
         );
  AOI22_X1 U4501 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_104), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_103), .ZN(n3913) );
  OAI221_X1 U4502 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_104), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_103), .A(n3913), .ZN(n3931) );
  OAI22_X1 U4503 ( .A1(n3947), .A2(keyinput_108), .B1(n3946), .B2(keyinput_109), .ZN(n3914) );
  AOI221_X1 U4504 ( .B1(n3947), .B2(keyinput_108), .C1(keyinput_109), .C2(
        n3946), .A(n3914), .ZN(n3917) );
  OAI22_X1 U4505 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_117), .B1(
        keyinput_106), .B2(REG3_REG_1__SCAN_IN), .ZN(n3915) );
  AOI221_X1 U4506 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_117), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_106), .A(n3915), .ZN(n3916) );
  OAI211_X1 U4507 ( .C1(n3919), .C2(keyinput_112), .A(n3917), .B(n3916), .ZN(
        n3918) );
  AOI21_X1 U4508 ( .B1(n3919), .B2(keyinput_112), .A(n3918), .ZN(n3930) );
  AOI22_X1 U4509 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_110), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_115), .ZN(n3920) );
  OAI221_X1 U4510 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_110), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_115), .A(n3920), .ZN(n3928) );
  AOI22_X1 U4511 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_107), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput_111), .ZN(n3921) );
  OAI221_X1 U4512 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_107), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_111), .A(n3921), .ZN(n3927) );
  AOI22_X1 U4513 ( .A1(n4016), .A2(keyinput_114), .B1(keyinput_105), .B2(n4535), .ZN(n3922) );
  OAI221_X1 U4514 ( .B1(n4016), .B2(keyinput_114), .C1(n4535), .C2(
        keyinput_105), .A(n3922), .ZN(n3926) );
  INV_X1 U4515 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4516 ( .A1(n3924), .A2(keyinput_116), .B1(n3952), .B2(keyinput_113), .ZN(n3923) );
  OAI221_X1 U4517 ( .B1(n3924), .B2(keyinput_116), .C1(n3952), .C2(
        keyinput_113), .A(n3923), .ZN(n3925) );
  NOR4_X1 U4518 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3929)
         );
  OAI211_X1 U4519 ( .C1(n3932), .C2(n3931), .A(n3930), .B(n3929), .ZN(n3933)
         );
  NAND3_X1 U4520 ( .A1(n3935), .A2(n3934), .A3(n3933), .ZN(n3936) );
  OAI221_X1 U4521 ( .B1(IR_REG_3__SCAN_IN), .B2(n3937), .C1(n4033), .C2(
        keyinput_122), .A(n3936), .ZN(n3938) );
  OAI221_X1 U4522 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_123), .C1(n4036), 
        .C2(n3939), .A(n3938), .ZN(n3940) );
  OAI211_X1 U4523 ( .C1(IR_REG_7__SCAN_IN), .C2(keyinput_126), .A(n3941), .B(
        n3940), .ZN(n3942) );
  AOI21_X1 U4524 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_126), .A(n3942), .ZN(
        n4045) );
  INV_X1 U4525 ( .A(keyinput_59), .ZN(n4037) );
  INV_X1 U4526 ( .A(keyinput_58), .ZN(n4034) );
  OAI22_X1 U4527 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_41), .B1(keyinput_52), .B2(REG3_REG_0__SCAN_IN), .ZN(n3943) );
  AOI221_X1 U4528 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_41), .C1(
        REG3_REG_0__SCAN_IN), .C2(keyinput_52), .A(n3943), .ZN(n4026) );
  OAI22_X1 U4529 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_47), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_48), .ZN(n3944) );
  AOI221_X1 U4530 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_47), .C1(
        keyinput_48), .C2(REG3_REG_17__SCAN_IN), .A(n3944), .ZN(n4025) );
  OAI22_X1 U4531 ( .A1(n3947), .A2(keyinput_44), .B1(n3946), .B2(keyinput_45), 
        .ZN(n3945) );
  AOI221_X1 U4532 ( .B1(n3947), .B2(keyinput_44), .C1(keyinput_45), .C2(n3946), 
        .A(n3945), .ZN(n3950) );
  OAI22_X1 U4533 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_51), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_43), .ZN(n3948) );
  AOI221_X1 U4534 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_51), .C1(
        keyinput_43), .C2(REG3_REG_21__SCAN_IN), .A(n3948), .ZN(n3949) );
  OAI211_X1 U4535 ( .C1(n3952), .C2(keyinput_49), .A(n3950), .B(n3949), .ZN(
        n3951) );
  AOI21_X1 U4536 ( .B1(n3952), .B2(keyinput_49), .A(n3951), .ZN(n4024) );
  OAI22_X1 U4537 ( .A1(n2819), .A2(keyinput_40), .B1(keyinput_39), .B2(
        REG3_REG_19__SCAN_IN), .ZN(n3953) );
  AOI221_X1 U4538 ( .B1(n2819), .B2(keyinput_40), .C1(REG3_REG_19__SCAN_IN), 
        .C2(keyinput_39), .A(n3953), .ZN(n4022) );
  INV_X1 U4539 ( .A(keyinput_32), .ZN(n4005) );
  INV_X1 U4540 ( .A(keyinput_31), .ZN(n4003) );
  INV_X1 U4541 ( .A(keyinput_30), .ZN(n4001) );
  INV_X1 U4542 ( .A(DATAI_4_), .ZN(n4702) );
  AOI22_X1 U4543 ( .A1(DATAI_3_), .A2(keyinput_28), .B1(n4702), .B2(
        keyinput_27), .ZN(n3954) );
  OAI221_X1 U4544 ( .B1(DATAI_3_), .B2(keyinput_28), .C1(n4702), .C2(
        keyinput_27), .A(n3954), .ZN(n3998) );
  INV_X1 U4545 ( .A(keyinput_26), .ZN(n3996) );
  INV_X1 U4546 ( .A(DATAI_12_), .ZN(n4781) );
  AOI22_X1 U4547 ( .A1(n4781), .A2(keyinput_19), .B1(keyinput_20), .B2(n4767), 
        .ZN(n3955) );
  OAI221_X1 U4548 ( .B1(n4781), .B2(keyinput_19), .C1(n4767), .C2(keyinput_20), 
        .A(n3955), .ZN(n3989) );
  OAI22_X1 U4549 ( .A1(DATAI_14_), .A2(keyinput_17), .B1(keyinput_18), .B2(
        DATAI_13_), .ZN(n3956) );
  AOI221_X1 U4550 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(DATAI_13_), .C2(
        keyinput_18), .A(n3956), .ZN(n3988) );
  XOR2_X1 U4551 ( .A(n3957), .B(keyinput_5), .Z(n3966) );
  OAI22_X1 U4552 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        DATAI_31_), .ZN(n3958) );
  AOI221_X1 U4553 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n3958), .ZN(n3963) );
  OAI22_X1 U4554 ( .A1(n3960), .A2(keyinput_4), .B1(keyinput_3), .B2(DATAI_28_), .ZN(n3959) );
  AOI221_X1 U4555 ( .B1(n3960), .B2(keyinput_4), .C1(DATAI_28_), .C2(
        keyinput_3), .A(n3959), .ZN(n3961) );
  OAI21_X1 U4556 ( .B1(n3964), .B2(keyinput_2), .A(n3961), .ZN(n3962) );
  AOI211_X1 U4557 ( .C1(n3964), .C2(keyinput_2), .A(n3963), .B(n3962), .ZN(
        n3965) );
  OAI22_X1 U4558 ( .A1(n3966), .A2(n3965), .B1(n3968), .B2(keyinput_6), .ZN(
        n3967) );
  AOI21_X1 U4559 ( .B1(n3968), .B2(keyinput_6), .A(n3967), .ZN(n3974) );
  OAI22_X1 U4560 ( .A1(n3970), .A2(keyinput_7), .B1(keyinput_8), .B2(DATAI_23_), .ZN(n3969) );
  AOI221_X1 U4561 ( .B1(n3970), .B2(keyinput_7), .C1(DATAI_23_), .C2(
        keyinput_8), .A(n3969), .ZN(n3973) );
  AOI22_X1 U4562 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(DATAI_22_), .B2(
        keyinput_9), .ZN(n3971) );
  OAI221_X1 U4563 ( .B1(DATAI_21_), .B2(keyinput_10), .C1(DATAI_22_), .C2(
        keyinput_9), .A(n3971), .ZN(n3972) );
  AOI21_X1 U4564 ( .B1(n3974), .B2(n3973), .A(n3972), .ZN(n3984) );
  AOI22_X1 U4565 ( .A1(n3977), .A2(keyinput_12), .B1(n3976), .B2(keyinput_11), 
        .ZN(n3975) );
  OAI221_X1 U4566 ( .B1(n3977), .B2(keyinput_12), .C1(n3976), .C2(keyinput_11), 
        .A(n3975), .ZN(n3983) );
  INV_X1 U4567 ( .A(DATAI_16_), .ZN(n4842) );
  OAI22_X1 U4568 ( .A1(n4842), .A2(keyinput_15), .B1(n3979), .B2(keyinput_16), 
        .ZN(n3978) );
  AOI221_X1 U4569 ( .B1(n4842), .B2(keyinput_15), .C1(keyinput_16), .C2(n3979), 
        .A(n3978), .ZN(n3982) );
  OAI22_X1 U4570 ( .A1(DATAI_18_), .A2(keyinput_13), .B1(DATAI_17_), .B2(
        keyinput_14), .ZN(n3980) );
  AOI221_X1 U4571 ( .B1(DATAI_18_), .B2(keyinput_13), .C1(keyinput_14), .C2(
        DATAI_17_), .A(n3980), .ZN(n3981) );
  OAI211_X1 U4572 ( .C1(n3984), .C2(n3983), .A(n3982), .B(n3981), .ZN(n3987)
         );
  INV_X1 U4573 ( .A(DATAI_9_), .ZN(n4756) );
  OAI22_X1 U4574 ( .A1(n4756), .A2(keyinput_22), .B1(DATAI_10_), .B2(
        keyinput_21), .ZN(n3985) );
  AOI221_X1 U4575 ( .B1(n4756), .B2(keyinput_22), .C1(keyinput_21), .C2(
        DATAI_10_), .A(n3985), .ZN(n3986) );
  OAI221_X1 U4576 ( .B1(n3989), .B2(n3988), .C1(n3989), .C2(n3987), .A(n3986), 
        .ZN(n3993) );
  INV_X1 U4577 ( .A(DATAI_8_), .ZN(n4747) );
  OAI22_X1 U4578 ( .A1(n4747), .A2(keyinput_23), .B1(n4719), .B2(keyinput_24), 
        .ZN(n3990) );
  AOI221_X1 U4579 ( .B1(n4747), .B2(keyinput_23), .C1(keyinput_24), .C2(n4719), 
        .A(n3990), .ZN(n3992) );
  NOR2_X1 U4580 ( .A1(DATAI_6_), .A2(keyinput_25), .ZN(n3991) );
  AOI221_X1 U4581 ( .B1(n3993), .B2(n3992), .C1(keyinput_25), .C2(DATAI_6_), 
        .A(n3991), .ZN(n3994) );
  AOI221_X1 U4582 ( .B1(DATAI_5_), .B2(n3996), .C1(n3995), .C2(keyinput_26), 
        .A(n3994), .ZN(n3997) );
  OAI22_X1 U4583 ( .A1(n3998), .A2(n3997), .B1(keyinput_29), .B2(DATAI_2_), 
        .ZN(n3999) );
  AOI21_X1 U4584 ( .B1(keyinput_29), .B2(DATAI_2_), .A(n3999), .ZN(n4000) );
  AOI221_X1 U4585 ( .B1(DATAI_1_), .B2(n4001), .C1(n2603), .C2(keyinput_30), 
        .A(n4000), .ZN(n4002) );
  AOI221_X1 U4586 ( .B1(DATAI_0_), .B2(n4003), .C1(n4599), .C2(keyinput_31), 
        .A(n4002), .ZN(n4004) );
  AOI221_X1 U4587 ( .B1(STATE_REG_SCAN_IN), .B2(n4005), .C1(U3149), .C2(
        keyinput_32), .A(n4004), .ZN(n4014) );
  AOI22_X1 U4588 ( .A1(n4008), .A2(keyinput_34), .B1(n4007), .B2(keyinput_33), 
        .ZN(n4006) );
  OAI221_X1 U4589 ( .B1(n4008), .B2(keyinput_34), .C1(n4007), .C2(keyinput_33), 
        .A(n4006), .ZN(n4013) );
  OAI22_X1 U4590 ( .A1(n4696), .A2(keyinput_38), .B1(keyinput_35), .B2(
        REG3_REG_14__SCAN_IN), .ZN(n4009) );
  AOI221_X1 U4591 ( .B1(n4696), .B2(keyinput_38), .C1(REG3_REG_14__SCAN_IN), 
        .C2(keyinput_35), .A(n4009), .ZN(n4012) );
  OAI22_X1 U4592 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_37), .B1(
        keyinput_36), .B2(REG3_REG_23__SCAN_IN), .ZN(n4010) );
  AOI221_X1 U4593 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_37), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_36), .A(n4010), .ZN(n4011) );
  OAI211_X1 U4594 ( .C1(n4014), .C2(n4013), .A(n4012), .B(n4011), .ZN(n4021)
         );
  AOI22_X1 U4595 ( .A1(n4590), .A2(keyinput_46), .B1(n4016), .B2(keyinput_50), 
        .ZN(n4015) );
  OAI221_X1 U4596 ( .B1(n4590), .B2(keyinput_46), .C1(n4016), .C2(keyinput_50), 
        .A(n4015), .ZN(n4020) );
  AOI22_X1 U4597 ( .A1(n3076), .A2(keyinput_42), .B1(n4018), .B2(keyinput_53), 
        .ZN(n4017) );
  OAI221_X1 U4598 ( .B1(n3076), .B2(keyinput_42), .C1(n4018), .C2(keyinput_53), 
        .A(n4017), .ZN(n4019) );
  AOI211_X1 U4599 ( .C1(n4022), .C2(n4021), .A(n4020), .B(n4019), .ZN(n4023)
         );
  NAND4_X1 U4600 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4031)
         );
  OAI22_X1 U4601 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_55), .B1(
        REG3_REG_13__SCAN_IN), .B2(keyinput_54), .ZN(n4027) );
  AOI221_X1 U4602 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_55), .C1(keyinput_54), 
        .C2(REG3_REG_13__SCAN_IN), .A(n4027), .ZN(n4030) );
  XOR2_X1 U4603 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .Z(n4029) );
  XNOR2_X1 U4604 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n4028) );
  NAND4_X1 U4605 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  OAI221_X1 U4606 ( .B1(IR_REG_3__SCAN_IN), .B2(n4034), .C1(n4033), .C2(
        keyinput_58), .A(n4032), .ZN(n4035) );
  OAI221_X1 U4607 ( .B1(IR_REG_4__SCAN_IN), .B2(n4037), .C1(n4036), .C2(
        keyinput_59), .A(n4035), .ZN(n4042) );
  XNOR2_X1 U4608 ( .A(n4038), .B(keyinput_62), .ZN(n4041) );
  XOR2_X1 U4609 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .Z(n4040) );
  XNOR2_X1 U4610 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4039) );
  NAND4_X1 U4611 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4044)
         );
  XNOR2_X1 U4612 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n4043) );
  OAI211_X1 U4613 ( .C1(n4046), .C2(n4045), .A(n4044), .B(n4043), .ZN(n4056)
         );
  OAI211_X1 U4614 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4048), .A(n4630), .B(n4047), .ZN(n4052) );
  OAI211_X1 U4615 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4050), .A(n4611), .B(n4049), .ZN(n4051) );
  OAI211_X1 U4616 ( .C1(n4643), .C2(n4759), .A(n4052), .B(n4051), .ZN(n4053)
         );
  AOI211_X1 U4617 ( .C1(n4629), .C2(ADDR_REG_10__SCAN_IN), .A(n4054), .B(n4053), .ZN(n4055) );
  XOR2_X1 U4618 ( .A(n4056), .B(n4055), .Z(U3250) );
  INV_X1 U4619 ( .A(n4643), .ZN(n4064) );
  AOI21_X1 U4620 ( .B1(n4629), .B2(ADDR_REG_14__SCAN_IN), .A(n4057), .ZN(n4058) );
  INV_X1 U4621 ( .A(n4058), .ZN(n4062) );
  AOI211_X1 U4622 ( .C1(n4060), .C2(n2285), .A(n4059), .B(n4633), .ZN(n4061)
         );
  AOI211_X1 U4623 ( .C1(n4064), .C2(n4063), .A(n4062), .B(n4061), .ZN(n4068)
         );
  OAI211_X1 U4624 ( .C1(n4066), .C2(REG1_REG_14__SCAN_IN), .A(n4630), .B(n4065), .ZN(n4067) );
  NAND2_X1 U4625 ( .A1(n4068), .A2(n4067), .ZN(U3254) );
  AND2_X1 U4626 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4810) );
  INV_X1 U4627 ( .A(n4069), .ZN(n4070) );
  AOI211_X1 U4628 ( .C1(n4072), .C2(n4071), .A(n4070), .B(n4633), .ZN(n4073)
         );
  AOI211_X1 U4629 ( .C1(n4629), .C2(ADDR_REG_15__SCAN_IN), .A(n4810), .B(n4073), .ZN(n4079) );
  AOI21_X1 U4630 ( .B1(n4486), .B2(n4832), .A(n4074), .ZN(n4075) );
  OAI21_X1 U4631 ( .B1(n4832), .B2(n4486), .A(n4075), .ZN(n4076) );
  NAND3_X1 U4632 ( .A1(n4630), .A2(n4077), .A3(n4076), .ZN(n4078) );
  OAI211_X1 U4633 ( .C1(n4080), .C2(n4643), .A(n4079), .B(n4078), .ZN(U3255)
         );
  AOI21_X1 U4634 ( .B1(n2288), .B2(n4082), .A(n4081), .ZN(n4092) );
  INV_X1 U4635 ( .A(n4630), .ZN(n4565) );
  AOI221_X1 U4636 ( .B1(n4085), .B2(n4084), .C1(n4083), .C2(n4084), .A(n4633), 
        .ZN(n4086) );
  OR2_X1 U4637 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  AOI21_X1 U4638 ( .B1(n4629), .B2(ADDR_REG_17__SCAN_IN), .A(n4088), .ZN(n4091) );
  OR2_X1 U4639 ( .A1(n4643), .A2(n4089), .ZN(n4090) );
  OAI211_X1 U4640 ( .C1(n4092), .C2(n4565), .A(n4091), .B(n4090), .ZN(U3257)
         );
  AOI21_X1 U4641 ( .B1(n4099), .B2(n4914), .A(n4097), .ZN(n4098) );
  OAI21_X1 U4642 ( .B1(n4914), .B2(n4099), .A(n4098), .ZN(n4100) );
  NAND3_X1 U4643 ( .A1(n4630), .A2(n4101), .A3(n4100), .ZN(n4102) );
  INV_X1 U4644 ( .A(n4104), .ZN(n4105) );
  NOR2_X1 U4645 ( .A1(n4106), .A2(n4105), .ZN(n4342) );
  AOI21_X1 U4646 ( .B1(n4107), .B2(n4902), .A(n4342), .ZN(n4432) );
  NOR2_X1 U4647 ( .A1(n4432), .A2(n4893), .ZN(n4108) );
  AOI21_X1 U4648 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4893), .A(n4108), .ZN(n4109) );
  OAI21_X1 U4649 ( .B1(n4435), .B2(n4886), .A(n4109), .ZN(U3260) );
  INV_X1 U4650 ( .A(n4110), .ZN(n4118) );
  NAND2_X1 U4651 ( .A1(n4669), .A2(n4111), .ZN(n4735) );
  NAND2_X1 U4652 ( .A1(n4770), .A2(n4735), .ZN(n4887) );
  OAI22_X1 U4653 ( .A1(n4113), .A2(n4886), .B1(n4112), .B2(n4882), .ZN(n4114)
         );
  OAI21_X1 U4654 ( .B1(n4115), .B2(n4114), .A(n4770), .ZN(n4117) );
  NAND2_X1 U4655 ( .A1(n4893), .A2(REG2_REG_29__SCAN_IN), .ZN(n4116) );
  OAI211_X1 U4656 ( .C1(n4118), .C2(n4887), .A(n4117), .B(n4116), .ZN(U3354)
         );
  XNOR2_X1 U4657 ( .A(n4119), .B(n4122), .ZN(n4348) );
  OAI22_X1 U4658 ( .A1(n4120), .A2(n4726), .B1(n4862), .B2(n4125), .ZN(n4123)
         );
  INV_X1 U4659 ( .A(n4347), .ZN(n4132) );
  OAI21_X1 U4660 ( .B1(n4144), .B2(n4125), .A(n4872), .ZN(n4126) );
  OR2_X1 U4661 ( .A1(n4127), .A2(n4126), .ZN(n4346) );
  AOI22_X1 U4662 ( .A1(n4893), .A2(REG2_REG_28__SCAN_IN), .B1(n4128), .B2(
        n4920), .ZN(n4129) );
  OAI21_X1 U4663 ( .B1(n4346), .B2(n4130), .A(n4129), .ZN(n4131) );
  AOI21_X1 U4664 ( .B1(n4132), .B2(n4770), .A(n4131), .ZN(n4133) );
  OAI21_X1 U4665 ( .B1(n4348), .B2(n4887), .A(n4133), .ZN(U3262) );
  OAI21_X1 U4666 ( .B1(n4142), .B2(n4135), .A(n4134), .ZN(n4136) );
  NAND2_X1 U4667 ( .A1(n4136), .A2(n4909), .ZN(n4139) );
  AOI22_X1 U4668 ( .A1(n4180), .A2(n4903), .B1(n4137), .B2(n4902), .ZN(n4138)
         );
  OAI211_X1 U4669 ( .C1(n4140), .C2(n4906), .A(n4139), .B(n4138), .ZN(n4349)
         );
  AOI21_X1 U4670 ( .B1(n4141), .B2(n4920), .A(n4349), .ZN(n4150) );
  XNOR2_X1 U4671 ( .A(n4143), .B(n4142), .ZN(n4350) );
  NAND2_X1 U4672 ( .A1(n4350), .A2(n4924), .ZN(n4149) );
  INV_X1 U4673 ( .A(n4144), .ZN(n4145) );
  OAI21_X1 U4674 ( .B1(n4152), .B2(n4146), .A(n4145), .ZN(n4443) );
  INV_X1 U4675 ( .A(n4443), .ZN(n4147) );
  AOI22_X1 U4676 ( .A1(n4147), .A2(n4981), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4893), .ZN(n4148) );
  OAI211_X1 U4677 ( .C1(n4893), .C2(n4150), .A(n4149), .B(n4148), .ZN(U3263)
         );
  AND2_X1 U4678 ( .A1(n4185), .A2(n4151), .ZN(n4153) );
  OR2_X1 U4679 ( .A1(n4153), .A2(n4152), .ZN(n4447) );
  XOR2_X1 U4680 ( .A(n4159), .B(n4154), .Z(n4354) );
  NAND2_X1 U4681 ( .A1(n4354), .A2(n4924), .ZN(n4170) );
  INV_X1 U4682 ( .A(n4155), .ZN(n4156) );
  NOR2_X1 U4683 ( .A1(n4157), .A2(n4156), .ZN(n4158) );
  XOR2_X1 U4684 ( .A(n4159), .B(n4158), .Z(n4165) );
  OAI22_X1 U4685 ( .A1(n4161), .A2(n4726), .B1(n4160), .B2(n4862), .ZN(n4162)
         );
  AOI21_X1 U4686 ( .B1(n4869), .B2(n4163), .A(n4162), .ZN(n4164) );
  OAI21_X1 U4687 ( .B1(n4165), .B2(n4864), .A(n4164), .ZN(n4353) );
  INV_X1 U4688 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4167) );
  OAI22_X1 U4689 ( .A1(n4770), .A2(n4167), .B1(n4166), .B2(n4882), .ZN(n4168)
         );
  AOI21_X1 U4690 ( .B1(n4353), .B2(n4770), .A(n4168), .ZN(n4169) );
  OAI211_X1 U4691 ( .C1(n4447), .C2(n4886), .A(n4170), .B(n4169), .ZN(U3264)
         );
  XNOR2_X1 U4692 ( .A(n4171), .B(n4175), .ZN(n4358) );
  INV_X1 U4693 ( .A(n4358), .ZN(n4190) );
  INV_X1 U4694 ( .A(n4172), .ZN(n4173) );
  NAND2_X1 U4695 ( .A1(n4174), .A2(n4173), .ZN(n4176) );
  XNOR2_X1 U4696 ( .A(n4176), .B(n4175), .ZN(n4182) );
  OAI22_X1 U4697 ( .A1(n4178), .A2(n4726), .B1(n4862), .B2(n4177), .ZN(n4179)
         );
  AOI21_X1 U4698 ( .B1(n4869), .B2(n4180), .A(n4179), .ZN(n4181) );
  OAI21_X1 U4699 ( .B1(n4182), .B2(n4864), .A(n4181), .ZN(n4357) );
  NAND2_X1 U4700 ( .A1(n4202), .A2(n4183), .ZN(n4184) );
  NAND2_X1 U4701 ( .A1(n4185), .A2(n4184), .ZN(n4451) );
  AOI22_X1 U4702 ( .A1(n4893), .A2(REG2_REG_25__SCAN_IN), .B1(n4186), .B2(
        n4920), .ZN(n4187) );
  OAI21_X1 U4703 ( .B1(n4451), .B2(n4886), .A(n4187), .ZN(n4188) );
  AOI21_X1 U4704 ( .B1(n4357), .B2(n4770), .A(n4188), .ZN(n4189) );
  OAI21_X1 U4705 ( .B1(n4190), .B2(n4887), .A(n4189), .ZN(U3265) );
  INV_X1 U4706 ( .A(n4191), .ZN(n4192) );
  NAND2_X1 U4707 ( .A1(n4193), .A2(n4192), .ZN(n4194) );
  XOR2_X1 U4708 ( .A(n4200), .B(n4194), .Z(n4199) );
  OAI22_X1 U4709 ( .A1(n4195), .A2(n4726), .B1(n4862), .B2(n4203), .ZN(n4196)
         );
  AOI21_X1 U4710 ( .B1(n4869), .B2(n4197), .A(n4196), .ZN(n4198) );
  OAI21_X1 U4711 ( .B1(n4199), .B2(n4864), .A(n4198), .ZN(n4361) );
  INV_X1 U4712 ( .A(n4361), .ZN(n4210) );
  XNOR2_X1 U4713 ( .A(n4201), .B(n4200), .ZN(n4362) );
  INV_X1 U4714 ( .A(n4211), .ZN(n4204) );
  OAI21_X1 U4715 ( .B1(n4204), .B2(n4203), .A(n4202), .ZN(n4455) );
  NOR2_X1 U4716 ( .A1(n4455), .A2(n4886), .ZN(n4208) );
  INV_X1 U4717 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4206) );
  OAI22_X1 U4718 ( .A1(n4770), .A2(n4206), .B1(n4205), .B2(n4882), .ZN(n4207)
         );
  AOI211_X1 U4719 ( .C1(n4362), .C2(n4924), .A(n4208), .B(n4207), .ZN(n4209)
         );
  OAI21_X1 U4720 ( .B1(n4210), .B2(n4893), .A(n4209), .ZN(U3266) );
  OAI21_X1 U4721 ( .B1(n4244), .B2(n4222), .A(n4211), .ZN(n4459) );
  OAI21_X1 U4722 ( .B1(n4258), .B2(n4213), .A(n4212), .ZN(n4236) );
  INV_X1 U4723 ( .A(n4236), .ZN(n4214) );
  NOR2_X1 U4724 ( .A1(n4214), .A2(n4239), .ZN(n4233) );
  NOR2_X1 U4725 ( .A1(n4233), .A2(n4215), .ZN(n4216) );
  XOR2_X1 U4726 ( .A(n4220), .B(n4216), .Z(n4366) );
  NAND2_X1 U4727 ( .A1(n4366), .A2(n4924), .ZN(n4232) );
  OAI21_X1 U4728 ( .B1(n4218), .B2(n4251), .A(n4217), .ZN(n4238) );
  NAND2_X1 U4729 ( .A1(n4239), .A2(n4238), .ZN(n4237) );
  NAND2_X1 U4730 ( .A1(n4219), .A2(n4237), .ZN(n4221) );
  XOR2_X1 U4731 ( .A(n4221), .B(n4220), .Z(n4227) );
  OAI22_X1 U4732 ( .A1(n4223), .A2(n4726), .B1(n4222), .B2(n4862), .ZN(n4224)
         );
  AOI21_X1 U4733 ( .B1(n4869), .B2(n4225), .A(n4224), .ZN(n4226) );
  OAI21_X1 U4734 ( .B1(n4227), .B2(n4864), .A(n4226), .ZN(n4365) );
  INV_X1 U4735 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4229) );
  OAI22_X1 U4736 ( .A1(n4770), .A2(n4229), .B1(n4228), .B2(n4882), .ZN(n4230)
         );
  AOI21_X1 U4737 ( .B1(n4365), .B2(n4770), .A(n4230), .ZN(n4231) );
  OAI211_X1 U4738 ( .C1(n4459), .C2(n4886), .A(n4232), .B(n4231), .ZN(U3267)
         );
  INV_X1 U4739 ( .A(n4239), .ZN(n4235) );
  INV_X1 U4740 ( .A(n4233), .ZN(n4234) );
  OAI21_X1 U4741 ( .B1(n4236), .B2(n4235), .A(n4234), .ZN(n4373) );
  OAI21_X1 U4742 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(n4243) );
  AOI22_X1 U4743 ( .A1(n4963), .A2(n4869), .B1(n4902), .B2(n4972), .ZN(n4240)
         );
  OAI21_X1 U4744 ( .B1(n4241), .B2(n4726), .A(n4240), .ZN(n4242) );
  AOI21_X1 U4745 ( .B1(n4243), .B2(n4909), .A(n4242), .ZN(n4372) );
  INV_X1 U4746 ( .A(n4244), .ZN(n4370) );
  INV_X1 U4747 ( .A(n4259), .ZN(n4245) );
  NAND2_X1 U4748 ( .A1(n4245), .A2(n4972), .ZN(n4369) );
  NAND3_X1 U4749 ( .A1(n4370), .A2(n4981), .A3(n4369), .ZN(n4248) );
  AOI22_X1 U4750 ( .A1(n4893), .A2(REG2_REG_22__SCAN_IN), .B1(n4920), .B2(
        n4246), .ZN(n4247) );
  OAI211_X1 U4751 ( .C1(n4893), .C2(n4372), .A(n4248), .B(n4247), .ZN(n4249)
         );
  INV_X1 U4752 ( .A(n4249), .ZN(n4250) );
  OAI21_X1 U4753 ( .B1(n4373), .B2(n4887), .A(n4250), .ZN(U3268) );
  XNOR2_X1 U4754 ( .A(n4251), .B(n4257), .ZN(n4256) );
  NAND2_X1 U4755 ( .A1(n4957), .A2(n4903), .ZN(n4253) );
  NAND2_X1 U4756 ( .A1(n4949), .A2(n4869), .ZN(n4252) );
  OAI211_X1 U4757 ( .C1(n4862), .C2(n4254), .A(n4253), .B(n4252), .ZN(n4255)
         );
  AOI21_X1 U4758 ( .B1(n4256), .B2(n4909), .A(n4255), .ZN(n4376) );
  XNOR2_X1 U4759 ( .A(n4258), .B(n4257), .ZN(n4374) );
  AOI21_X1 U4760 ( .B1(n4958), .B2(n2275), .A(n4259), .ZN(n4463) );
  INV_X1 U4761 ( .A(n4463), .ZN(n4262) );
  AOI22_X1 U4762 ( .A1(n4893), .A2(REG2_REG_21__SCAN_IN), .B1(n4260), .B2(
        n4920), .ZN(n4261) );
  OAI21_X1 U4763 ( .B1(n4262), .B2(n4886), .A(n4261), .ZN(n4263) );
  AOI21_X1 U4764 ( .B1(n4374), .B2(n4924), .A(n4263), .ZN(n4264) );
  OAI21_X1 U4765 ( .B1(n4376), .B2(n4893), .A(n4264), .ZN(U3269) );
  XNOR2_X1 U4766 ( .A(n4266), .B(n4265), .ZN(n4276) );
  NOR2_X1 U4767 ( .A1(n4268), .A2(n4267), .ZN(n4270) );
  XNOR2_X1 U4768 ( .A(n4270), .B(n4269), .ZN(n4271) );
  NAND2_X1 U4769 ( .A1(n4271), .A2(n4909), .ZN(n4273) );
  AOI22_X1 U4770 ( .A1(n4971), .A2(n4869), .B1(n4945), .B2(n4902), .ZN(n4272)
         );
  OAI211_X1 U4771 ( .C1(n4907), .C2(n4726), .A(n4273), .B(n4272), .ZN(n4274)
         );
  INV_X1 U4772 ( .A(n4274), .ZN(n4275) );
  OAI21_X1 U4773 ( .B1(n4276), .B2(n4669), .A(n4275), .ZN(n4379) );
  INV_X1 U4774 ( .A(n4379), .ZN(n4282) );
  INV_X1 U4775 ( .A(n4276), .ZN(n4380) );
  NAND2_X1 U4776 ( .A1(n2302), .A2(n4945), .ZN(n4277) );
  NAND2_X1 U4777 ( .A1(n2275), .A2(n4277), .ZN(n4468) );
  AOI22_X1 U4778 ( .A1(n4893), .A2(REG2_REG_20__SCAN_IN), .B1(n4278), .B2(
        n4920), .ZN(n4279) );
  OAI21_X1 U4779 ( .B1(n4468), .B2(n4886), .A(n4279), .ZN(n4280) );
  AOI21_X1 U4780 ( .B1(n4380), .B2(n4776), .A(n4280), .ZN(n4281) );
  OAI21_X1 U4781 ( .B1(n4282), .B2(n4893), .A(n4281), .ZN(U3270) );
  OR2_X1 U4782 ( .A1(n4283), .A2(n4899), .ZN(n4894) );
  NAND2_X1 U4783 ( .A1(n4894), .A2(n4284), .ZN(n4285) );
  XOR2_X1 U4784 ( .A(n4292), .B(n4285), .Z(n4384) );
  INV_X1 U4785 ( .A(n4384), .ZN(n4303) );
  INV_X1 U4786 ( .A(n4390), .ZN(n4289) );
  INV_X1 U4787 ( .A(n4286), .ZN(n4287) );
  OAI21_X1 U4788 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n4900) );
  OAI21_X1 U4789 ( .B1(n4900), .B2(n4291), .A(n4290), .ZN(n4293) );
  XNOR2_X1 U4790 ( .A(n4293), .B(n4292), .ZN(n4296) );
  OAI22_X1 U4791 ( .A1(n4393), .A2(n4726), .B1(n4297), .B2(n4862), .ZN(n4294)
         );
  AOI21_X1 U4792 ( .B1(n4869), .B2(n4957), .A(n4294), .ZN(n4295) );
  OAI21_X1 U4793 ( .B1(n4296), .B2(n4864), .A(n4295), .ZN(n4383) );
  OR2_X1 U4794 ( .A1(n4897), .A2(n4297), .ZN(n4298) );
  NAND2_X1 U4795 ( .A1(n2302), .A2(n4298), .ZN(n4472) );
  AOI22_X1 U4796 ( .A1(n4893), .A2(REG2_REG_19__SCAN_IN), .B1(n4299), .B2(
        n4920), .ZN(n4300) );
  OAI21_X1 U4797 ( .B1(n4472), .B2(n4886), .A(n4300), .ZN(n4301) );
  AOI21_X1 U4798 ( .B1(n4383), .B2(n4770), .A(n4301), .ZN(n4302) );
  OAI21_X1 U4799 ( .B1(n4303), .B2(n4887), .A(n4302), .ZN(U3271) );
  XNOR2_X1 U4800 ( .A(n4403), .B(n4312), .ZN(n4793) );
  INV_X1 U4801 ( .A(n4304), .ZN(n4305) );
  AOI21_X1 U4802 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(n4422) );
  INV_X1 U4803 ( .A(n4308), .ZN(n4309) );
  AOI21_X1 U4804 ( .B1(n4422), .B2(n4310), .A(n4309), .ZN(n4311) );
  XOR2_X1 U4805 ( .A(n4312), .B(n4311), .Z(n4317) );
  AOI22_X1 U4806 ( .A1(n4313), .A2(n4903), .B1(n4320), .B2(n4902), .ZN(n4314)
         );
  OAI21_X1 U4807 ( .B1(n4315), .B2(n4906), .A(n4314), .ZN(n4316) );
  AOI21_X1 U4808 ( .B1(n4317), .B2(n4909), .A(n4316), .ZN(n4318) );
  OAI21_X1 U4809 ( .B1(n4793), .B2(n4669), .A(n4318), .ZN(n4794) );
  NAND2_X1 U4810 ( .A1(n4794), .A2(n4770), .ZN(n4324) );
  INV_X1 U4811 ( .A(n4319), .ZN(n4399) );
  AOI21_X1 U4812 ( .B1(n4320), .B2(n4417), .A(n4399), .ZN(n4796) );
  OAI22_X1 U4813 ( .A1(n4770), .A2(n4583), .B1(n4321), .B2(n4882), .ZN(n4322)
         );
  AOI21_X1 U4814 ( .B1(n4796), .B2(n4981), .A(n4322), .ZN(n4323) );
  OAI211_X1 U4815 ( .C1(n4793), .C2(n4325), .A(n4324), .B(n4323), .ZN(U3277)
         );
  NAND2_X1 U4816 ( .A1(n4326), .A2(n4924), .ZN(n4334) );
  NOR2_X1 U4817 ( .A1(n4327), .A2(n4882), .ZN(n4328) );
  AOI21_X1 U4818 ( .B1(n4893), .B2(REG2_REG_5__SCAN_IN), .A(n4328), .ZN(n4333)
         );
  NAND2_X1 U4819 ( .A1(n4329), .A2(n4770), .ZN(n4332) );
  NAND2_X1 U4820 ( .A1(n4330), .A2(n4981), .ZN(n4331) );
  NAND4_X1 U4821 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(U3285)
         );
  NOR2_X1 U4822 ( .A1(n4432), .A2(n4913), .ZN(n4335) );
  AOI21_X1 U4823 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4913), .A(n4335), .ZN(n4336) );
  OAI21_X1 U4824 ( .B1(n4435), .B2(n4431), .A(n4336), .ZN(U3549) );
  INV_X1 U4825 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4345) );
  AOI21_X1 U4826 ( .B1(n4339), .B2(n4338), .A(n4337), .ZN(n4982) );
  NAND2_X1 U4827 ( .A1(n4982), .A2(n4689), .ZN(n4344) );
  NOR2_X1 U4828 ( .A1(n4340), .A2(n4862), .ZN(n4341) );
  OR2_X1 U4829 ( .A1(n4342), .A2(n4341), .ZN(n4980) );
  NAND2_X1 U4830 ( .A1(n4980), .A2(n4915), .ZN(n4343) );
  OAI211_X1 U4831 ( .C1(n4915), .C2(n4345), .A(n4344), .B(n4343), .ZN(U3548)
         );
  INV_X1 U4832 ( .A(n4912), .ZN(n4858) );
  OAI211_X1 U4833 ( .C1(n4348), .C2(n4858), .A(n4347), .B(n4346), .ZN(n4439)
         );
  MUX2_X1 U4834 ( .A(REG1_REG_28__SCAN_IN), .B(n4439), .S(n4915), .Z(U3546) );
  INV_X1 U4835 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4351) );
  AOI21_X1 U4836 ( .B1(n4350), .B2(n4912), .A(n4349), .ZN(n4440) );
  MUX2_X1 U4837 ( .A(n4351), .B(n4440), .S(n4915), .Z(n4352) );
  OAI21_X1 U4838 ( .B1(n4431), .B2(n4443), .A(n4352), .ZN(U3545) );
  INV_X1 U4839 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4355) );
  AOI21_X1 U4840 ( .B1(n4354), .B2(n4912), .A(n4353), .ZN(n4444) );
  MUX2_X1 U4841 ( .A(n4355), .B(n4444), .S(n4915), .Z(n4356) );
  OAI21_X1 U4842 ( .B1(n4431), .B2(n4447), .A(n4356), .ZN(U3544) );
  INV_X1 U4843 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4359) );
  AOI21_X1 U4844 ( .B1(n4358), .B2(n4912), .A(n4357), .ZN(n4448) );
  MUX2_X1 U4845 ( .A(n4359), .B(n4448), .S(n4915), .Z(n4360) );
  OAI21_X1 U4846 ( .B1(n4431), .B2(n4451), .A(n4360), .ZN(U3543) );
  INV_X1 U4847 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4363) );
  AOI21_X1 U4848 ( .B1(n4362), .B2(n4912), .A(n4361), .ZN(n4452) );
  MUX2_X1 U4849 ( .A(n4363), .B(n4452), .S(n4915), .Z(n4364) );
  OAI21_X1 U4850 ( .B1(n4431), .B2(n4455), .A(n4364), .ZN(U3542) );
  INV_X1 U4851 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4367) );
  AOI21_X1 U4852 ( .B1(n4366), .B2(n4912), .A(n4365), .ZN(n4456) );
  MUX2_X1 U4853 ( .A(n4367), .B(n4456), .S(n4915), .Z(n4368) );
  OAI21_X1 U4854 ( .B1(n4431), .B2(n4459), .A(n4368), .ZN(U3541) );
  NAND3_X1 U4855 ( .A1(n4370), .A2(n4872), .A3(n4369), .ZN(n4371) );
  OAI211_X1 U4856 ( .C1(n4373), .C2(n4858), .A(n4372), .B(n4371), .ZN(n4460)
         );
  MUX2_X1 U4857 ( .A(REG1_REG_22__SCAN_IN), .B(n4460), .S(n4915), .Z(U3540) );
  NAND2_X1 U4858 ( .A1(n4374), .A2(n4912), .ZN(n4375) );
  NAND2_X1 U4859 ( .A1(n4376), .A2(n4375), .ZN(n4461) );
  MUX2_X1 U4860 ( .A(REG1_REG_21__SCAN_IN), .B(n4461), .S(n4915), .Z(n4377) );
  AOI21_X1 U4861 ( .B1(n4689), .B2(n4463), .A(n4377), .ZN(n4378) );
  INV_X1 U4862 ( .A(n4378), .ZN(U3539) );
  INV_X1 U4863 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4381) );
  AOI21_X1 U4864 ( .B1(n4705), .B2(n4380), .A(n4379), .ZN(n4465) );
  MUX2_X1 U4865 ( .A(n4381), .B(n4465), .S(n4915), .Z(n4382) );
  OAI21_X1 U4866 ( .B1(n4431), .B2(n4468), .A(n4382), .ZN(U3538) );
  AOI21_X1 U4867 ( .B1(n4912), .B2(n4384), .A(n4383), .ZN(n4469) );
  MUX2_X1 U4868 ( .A(n2953), .B(n4469), .S(n4915), .Z(n4385) );
  OAI21_X1 U4869 ( .B1(n4431), .B2(n4472), .A(n4385), .ZN(U3537) );
  INV_X1 U4870 ( .A(n4386), .ZN(n4853) );
  OAI21_X1 U4871 ( .B1(n4853), .B2(n4387), .A(n2298), .ZN(n4885) );
  XNOR2_X1 U4872 ( .A(n4388), .B(n4389), .ZN(n4884) );
  XNOR2_X1 U4873 ( .A(n4390), .B(n4389), .ZN(n4395) );
  AOI22_X1 U4874 ( .A1(n4830), .A2(n4903), .B1(n4391), .B2(n4902), .ZN(n4392)
         );
  OAI21_X1 U4875 ( .B1(n4393), .B2(n4906), .A(n4392), .ZN(n4394) );
  AOI21_X1 U4876 ( .B1(n4395), .B2(n4909), .A(n4394), .ZN(n4892) );
  INV_X1 U4877 ( .A(n4892), .ZN(n4396) );
  AOI21_X1 U4878 ( .B1(n4884), .B2(n4912), .A(n4396), .ZN(n4473) );
  MUX2_X1 U4879 ( .A(n2950), .B(n4473), .S(n4915), .Z(n4397) );
  OAI21_X1 U4880 ( .B1(n4431), .B2(n4885), .A(n4397), .ZN(U3535) );
  INV_X1 U4881 ( .A(n4822), .ZN(n4398) );
  OAI21_X1 U4882 ( .B1(n4399), .B2(n4410), .A(n4398), .ZN(n4801) );
  INV_X1 U4883 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4414) );
  INV_X1 U4884 ( .A(n4400), .ZN(n4402) );
  OAI21_X1 U4885 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(n4404) );
  NAND2_X1 U4886 ( .A1(n4404), .A2(n4405), .ZN(n4820) );
  OAI21_X1 U4887 ( .B1(n4404), .B2(n4405), .A(n4820), .ZN(n4803) );
  XNOR2_X1 U4888 ( .A(n4406), .B(n2409), .ZN(n4412) );
  NAND2_X1 U4889 ( .A1(n4859), .A2(n4869), .ZN(n4409) );
  NAND2_X1 U4890 ( .A1(n4407), .A2(n4903), .ZN(n4408) );
  OAI211_X1 U4891 ( .C1(n4862), .C2(n4410), .A(n4409), .B(n4408), .ZN(n4411)
         );
  AOI21_X1 U4892 ( .B1(n4412), .B2(n4909), .A(n4411), .ZN(n4806) );
  INV_X1 U4893 ( .A(n4806), .ZN(n4413) );
  AOI21_X1 U4894 ( .B1(n4803), .B2(n4912), .A(n4413), .ZN(n4476) );
  MUX2_X1 U4895 ( .A(n4414), .B(n4476), .S(n4915), .Z(n4415) );
  OAI21_X1 U4896 ( .B1(n4801), .B2(n4431), .A(n4415), .ZN(U3532) );
  INV_X1 U4897 ( .A(n4416), .ZN(n4419) );
  OAI21_X1 U4898 ( .B1(n4419), .B2(n4418), .A(n4417), .ZN(n4784) );
  XNOR2_X1 U4899 ( .A(n4420), .B(n4421), .ZN(n4786) );
  XNOR2_X1 U4900 ( .A(n4422), .B(n4421), .ZN(n4428) );
  AOI22_X1 U4901 ( .A1(n4424), .A2(n4903), .B1(n4423), .B2(n4902), .ZN(n4425)
         );
  OAI21_X1 U4902 ( .B1(n4426), .B2(n4906), .A(n4425), .ZN(n4427) );
  AOI21_X1 U4903 ( .B1(n4428), .B2(n4909), .A(n4427), .ZN(n4789) );
  INV_X1 U4904 ( .A(n4789), .ZN(n4429) );
  AOI21_X1 U4905 ( .B1(n4912), .B2(n4786), .A(n4429), .ZN(n4479) );
  MUX2_X1 U4906 ( .A(n4568), .B(n4479), .S(n4915), .Z(n4430) );
  OAI21_X1 U4907 ( .B1(n4784), .B2(n4431), .A(n4430), .ZN(U3530) );
  NOR2_X1 U4908 ( .A1(n4432), .A2(n4916), .ZN(n4433) );
  AOI21_X1 U4909 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4916), .A(n4433), .ZN(n4434) );
  OAI21_X1 U4910 ( .B1(n4435), .B2(n4482), .A(n4434), .ZN(U3517) );
  INV_X1 U4911 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U4912 ( .A1(n4982), .A2(n4692), .ZN(n4437) );
  NAND2_X1 U4913 ( .A1(n4980), .A2(n4919), .ZN(n4436) );
  OAI211_X1 U4914 ( .C1(n4919), .C2(n4438), .A(n4437), .B(n4436), .ZN(U3516)
         );
  MUX2_X1 U4915 ( .A(REG0_REG_28__SCAN_IN), .B(n4439), .S(n4919), .Z(U3514) );
  INV_X1 U4916 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4441) );
  MUX2_X1 U4917 ( .A(n4441), .B(n4440), .S(n4919), .Z(n4442) );
  OAI21_X1 U4918 ( .B1(n4443), .B2(n4482), .A(n4442), .ZN(U3513) );
  INV_X1 U4919 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4445) );
  MUX2_X1 U4920 ( .A(n4445), .B(n4444), .S(n4919), .Z(n4446) );
  OAI21_X1 U4921 ( .B1(n4447), .B2(n4482), .A(n4446), .ZN(U3512) );
  INV_X1 U4922 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4449) );
  MUX2_X1 U4923 ( .A(n4449), .B(n4448), .S(n4919), .Z(n4450) );
  OAI21_X1 U4924 ( .B1(n4451), .B2(n4482), .A(n4450), .ZN(U3511) );
  INV_X1 U4925 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4453) );
  MUX2_X1 U4926 ( .A(n4453), .B(n4452), .S(n4919), .Z(n4454) );
  OAI21_X1 U4927 ( .B1(n4455), .B2(n4482), .A(n4454), .ZN(U3510) );
  INV_X1 U4928 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4457) );
  MUX2_X1 U4929 ( .A(n4457), .B(n4456), .S(n4919), .Z(n4458) );
  OAI21_X1 U4930 ( .B1(n4459), .B2(n4482), .A(n4458), .ZN(U3509) );
  MUX2_X1 U4931 ( .A(REG0_REG_22__SCAN_IN), .B(n4460), .S(n4919), .Z(U3508) );
  MUX2_X1 U4932 ( .A(REG0_REG_21__SCAN_IN), .B(n4461), .S(n4919), .Z(n4462) );
  AOI21_X1 U4933 ( .B1(n4463), .B2(n4692), .A(n4462), .ZN(n4464) );
  INV_X1 U4934 ( .A(n4464), .ZN(U3507) );
  INV_X1 U4935 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U4936 ( .A(n4466), .B(n4465), .S(n4919), .Z(n4467) );
  OAI21_X1 U4937 ( .B1(n4468), .B2(n4482), .A(n4467), .ZN(U3506) );
  INV_X1 U4938 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U4939 ( .A(n4470), .B(n4469), .S(n4919), .Z(n4471) );
  OAI21_X1 U4940 ( .B1(n4472), .B2(n4482), .A(n4471), .ZN(U3505) );
  INV_X1 U4941 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U4942 ( .A(n4474), .B(n4473), .S(n4919), .Z(n4475) );
  OAI21_X1 U4943 ( .B1(n4885), .B2(n4482), .A(n4475), .ZN(U3501) );
  INV_X1 U4944 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4477) );
  MUX2_X1 U4945 ( .A(n4477), .B(n4476), .S(n4919), .Z(n4478) );
  OAI21_X1 U4946 ( .B1(n4801), .B2(n4482), .A(n4478), .ZN(U3495) );
  INV_X1 U4947 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4480) );
  MUX2_X1 U4948 ( .A(n4480), .B(n4479), .S(n4919), .Z(n4481) );
  OAI21_X1 U4949 ( .B1(n4784), .B2(n4482), .A(n4481), .ZN(U3491) );
  MUX2_X1 U4950 ( .A(DATAI_30_), .B(n4483), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4951 ( .A(n4494), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4952 ( .A(n4484), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4953 ( .A(DATAI_19_), .B(n4485), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4954 ( .A(DATAI_15_), .B(n4486), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U4955 ( .A(DATAI_5_), .B(n4487), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U4956 ( .A(n4615), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4957 ( .A(n4488), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4958 ( .A(DATAI_23_), .ZN(n4490) );
  OAI21_X1 U4959 ( .B1(STATE_REG_SCAN_IN), .B2(n4490), .A(n4489), .ZN(U3329)
         );
  AND2_X1 U4960 ( .A1(D_REG_2__SCAN_IN), .A2(n4491), .ZN(U3320) );
  AND2_X1 U4961 ( .A1(D_REG_3__SCAN_IN), .A2(n4491), .ZN(U3319) );
  AND2_X1 U4962 ( .A1(D_REG_4__SCAN_IN), .A2(n4491), .ZN(U3318) );
  AND2_X1 U4963 ( .A1(D_REG_5__SCAN_IN), .A2(n4491), .ZN(U3317) );
  AND2_X1 U4964 ( .A1(D_REG_6__SCAN_IN), .A2(n4491), .ZN(U3316) );
  AND2_X1 U4965 ( .A1(D_REG_7__SCAN_IN), .A2(n4491), .ZN(U3315) );
  AND2_X1 U4966 ( .A1(D_REG_8__SCAN_IN), .A2(n4491), .ZN(U3314) );
  AND2_X1 U4967 ( .A1(D_REG_9__SCAN_IN), .A2(n4491), .ZN(U3313) );
  AND2_X1 U4968 ( .A1(D_REG_10__SCAN_IN), .A2(n4491), .ZN(U3312) );
  AND2_X1 U4969 ( .A1(D_REG_11__SCAN_IN), .A2(n4491), .ZN(U3311) );
  AND2_X1 U4970 ( .A1(D_REG_12__SCAN_IN), .A2(n4491), .ZN(U3310) );
  AND2_X1 U4971 ( .A1(D_REG_13__SCAN_IN), .A2(n4491), .ZN(U3309) );
  AND2_X1 U4972 ( .A1(D_REG_14__SCAN_IN), .A2(n4491), .ZN(U3308) );
  AND2_X1 U4973 ( .A1(D_REG_15__SCAN_IN), .A2(n4491), .ZN(U3307) );
  AND2_X1 U4974 ( .A1(D_REG_16__SCAN_IN), .A2(n4491), .ZN(U3306) );
  AND2_X1 U4975 ( .A1(D_REG_17__SCAN_IN), .A2(n4491), .ZN(U3305) );
  AND2_X1 U4976 ( .A1(D_REG_18__SCAN_IN), .A2(n4491), .ZN(U3304) );
  AND2_X1 U4977 ( .A1(D_REG_19__SCAN_IN), .A2(n4491), .ZN(U3303) );
  AND2_X1 U4978 ( .A1(D_REG_20__SCAN_IN), .A2(n4491), .ZN(U3302) );
  AND2_X1 U4979 ( .A1(D_REG_21__SCAN_IN), .A2(n4491), .ZN(U3301) );
  AND2_X1 U4980 ( .A1(D_REG_22__SCAN_IN), .A2(n4491), .ZN(U3300) );
  AND2_X1 U4981 ( .A1(D_REG_23__SCAN_IN), .A2(n4491), .ZN(U3299) );
  AND2_X1 U4982 ( .A1(D_REG_24__SCAN_IN), .A2(n4491), .ZN(U3298) );
  AND2_X1 U4983 ( .A1(D_REG_25__SCAN_IN), .A2(n4491), .ZN(U3297) );
  AND2_X1 U4984 ( .A1(D_REG_26__SCAN_IN), .A2(n4491), .ZN(U3296) );
  AND2_X1 U4985 ( .A1(D_REG_27__SCAN_IN), .A2(n4491), .ZN(U3295) );
  AND2_X1 U4986 ( .A1(D_REG_28__SCAN_IN), .A2(n4491), .ZN(U3294) );
  AND2_X1 U4987 ( .A1(D_REG_29__SCAN_IN), .A2(n4491), .ZN(U3293) );
  AND2_X1 U4988 ( .A1(D_REG_30__SCAN_IN), .A2(n4491), .ZN(U3292) );
  AND2_X1 U4989 ( .A1(D_REG_31__SCAN_IN), .A2(n4491), .ZN(U3291) );
  INV_X1 U4990 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U4991 ( .A1(n4494), .A2(n4657), .ZN(n4492) );
  NAND2_X1 U4992 ( .A1(n4604), .A2(n4492), .ZN(n4608) );
  INV_X1 U4993 ( .A(n4608), .ZN(n4493) );
  OAI211_X1 U4994 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4494), .A(n4493), .B(n4495), 
        .ZN(n4498) );
  AOI22_X1 U4995 ( .A1(n4495), .A2(n4608), .B1(n4630), .B2(n4648), .ZN(n4497)
         );
  AOI22_X1 U4996 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4629), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4496) );
  OAI221_X1 U4997 ( .B1(IR_REG_0__SCAN_IN), .B2(n4498), .C1(n4609), .C2(n4497), 
        .A(n4496), .ZN(U3240) );
  AOI211_X1 U4998 ( .C1(n4501), .C2(n4500), .A(n4499), .B(n4633), .ZN(n4503)
         );
  AOI211_X1 U4999 ( .C1(n4629), .C2(ADDR_REG_3__SCAN_IN), .A(n4503), .B(n4502), 
        .ZN(n4507) );
  OAI211_X1 U5000 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4505), .A(n4630), .B(n4504), 
        .ZN(n4506) );
  OAI211_X1 U5001 ( .C1(n4643), .C2(n2927), .A(n4507), .B(n4506), .ZN(U3243)
         );
  AOI211_X1 U5002 ( .C1(n4510), .C2(n4509), .A(n4508), .B(n4633), .ZN(n4512)
         );
  AOI211_X1 U5003 ( .C1(n4629), .C2(ADDR_REG_6__SCAN_IN), .A(n4512), .B(n4511), 
        .ZN(n4516) );
  OAI211_X1 U5004 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4514), .A(n4630), .B(n4513), 
        .ZN(n4515) );
  OAI211_X1 U5005 ( .C1(n4643), .C2(n2342), .A(n4516), .B(n4515), .ZN(U3246)
         );
  AOI21_X1 U5006 ( .B1(n4629), .B2(ADDR_REG_7__SCAN_IN), .A(n4517), .ZN(n4531)
         );
  NAND3_X1 U5007 ( .A1(n4527), .A2(n4630), .A3(REG1_REG_7__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U5008 ( .A1(n4518), .A2(n4643), .ZN(n4524) );
  INV_X1 U5009 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5010 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4521), .B1(n4520), .B2(n4519), .ZN(n4522) );
  XOR2_X1 U5011 ( .A(n4720), .B(n4522), .Z(n4523) );
  AOI22_X1 U5012 ( .A1(n4525), .A2(n4524), .B1(n4611), .B2(n4523), .ZN(n4530)
         );
  OAI211_X1 U5013 ( .C1(n4528), .C2(n4527), .A(n4630), .B(n4526), .ZN(n4529)
         );
  NAND3_X1 U5014 ( .A1(n4531), .A2(n4530), .A3(n4529), .ZN(U3247) );
  AOI211_X1 U5015 ( .C1(n4534), .C2(n4533), .A(n4532), .B(n4565), .ZN(n4537)
         );
  NOR2_X1 U5016 ( .A1(STATE_REG_SCAN_IN), .A2(n4535), .ZN(n4536) );
  AOI211_X1 U5017 ( .C1(n4629), .C2(ADDR_REG_8__SCAN_IN), .A(n4537), .B(n4536), 
        .ZN(n4541) );
  OAI211_X1 U5018 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4539), .A(n4611), .B(n4538), 
        .ZN(n4540) );
  OAI211_X1 U5019 ( .C1(n4643), .C2(n4748), .A(n4541), .B(n4540), .ZN(U3248)
         );
  AOI22_X1 U5020 ( .A1(n4543), .A2(n4542), .B1(REG1_REG_9__SCAN_IN), .B2(n4757), .ZN(n4545) );
  OAI21_X1 U5021 ( .B1(n4546), .B2(n4545), .A(n4630), .ZN(n4544) );
  AOI21_X1 U5022 ( .B1(n4546), .B2(n4545), .A(n4544), .ZN(n4548) );
  AOI211_X1 U5023 ( .C1(n4629), .C2(ADDR_REG_9__SCAN_IN), .A(n4548), .B(n4547), 
        .ZN(n4553) );
  OAI211_X1 U5024 ( .C1(n4551), .C2(n4550), .A(n4611), .B(n4549), .ZN(n4552)
         );
  OAI211_X1 U5025 ( .C1(n4643), .C2(n4757), .A(n4553), .B(n4552), .ZN(U3249)
         );
  AOI22_X1 U5026 ( .A1(n4554), .A2(REG1_REG_11__SCAN_IN), .B1(n2939), .B2(
        n2940), .ZN(n4557) );
  OAI21_X1 U5027 ( .B1(n4557), .B2(n4556), .A(n4630), .ZN(n4555) );
  AOI21_X1 U5028 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(n4559) );
  AOI211_X1 U5029 ( .C1(n4629), .C2(ADDR_REG_11__SCAN_IN), .A(n4559), .B(n4558), .ZN(n4564) );
  OAI211_X1 U5030 ( .C1(n4562), .C2(n4561), .A(n4611), .B(n4560), .ZN(n4563)
         );
  OAI211_X1 U5031 ( .C1(n4643), .C2(n2940), .A(n4564), .B(n4563), .ZN(U3251)
         );
  AOI211_X1 U5032 ( .C1(n4568), .C2(n4567), .A(n4566), .B(n4565), .ZN(n4570)
         );
  AOI211_X1 U5033 ( .C1(n4629), .C2(ADDR_REG_12__SCAN_IN), .A(n4570), .B(n4569), .ZN(n4574) );
  OAI211_X1 U5034 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4572), .A(n4611), .B(n4571), .ZN(n4573) );
  OAI211_X1 U5035 ( .C1(n4643), .C2(n4782), .A(n4574), .B(n4573), .ZN(U3252)
         );
  NAND2_X1 U5036 ( .A1(n4576), .A2(n4575), .ZN(n4578) );
  OAI21_X1 U5037 ( .B1(n4579), .B2(n4578), .A(n4630), .ZN(n4577) );
  AOI21_X1 U5038 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n4581) );
  AOI211_X1 U5039 ( .C1(n4629), .C2(ADDR_REG_13__SCAN_IN), .A(n4581), .B(n4580), .ZN(n4588) );
  AOI21_X1 U5040 ( .B1(n4589), .B2(n4583), .A(n4582), .ZN(n4586) );
  AOI21_X1 U5041 ( .B1(n4586), .B2(n4585), .A(n4633), .ZN(n4584) );
  OAI21_X1 U5042 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n4587) );
  OAI211_X1 U5043 ( .C1(n4643), .C2(n4589), .A(n4588), .B(n4587), .ZN(U3253)
         );
  NOR2_X1 U5044 ( .A1(STATE_REG_SCAN_IN), .A2(n4590), .ZN(n4849) );
  AOI221_X1 U5045 ( .B1(n4593), .B2(n4592), .C1(n4591), .C2(n4592), .A(n4633), 
        .ZN(n4594) );
  AOI211_X1 U5046 ( .C1(n4629), .C2(ADDR_REG_16__SCAN_IN), .A(n4849), .B(n4594), .ZN(n4598) );
  OAI221_X1 U5047 ( .B1(n4596), .B2(REG1_REG_16__SCAN_IN), .C1(n4596), .C2(
        n4595), .A(n4630), .ZN(n4597) );
  OAI211_X1 U5048 ( .C1(n4643), .C2(n4843), .A(n4598), .B(n4597), .ZN(U3256)
         );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n4609), .B1(n4599), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5050 ( .A(n4600), .ZN(n4602) );
  OAI21_X1 U5051 ( .B1(n4602), .B2(n4601), .A(U4043), .ZN(n4607) );
  AND3_X1 U5052 ( .A1(n4605), .A2(n4604), .A3(n4603), .ZN(n4606) );
  AOI211_X1 U5053 ( .C1(n4609), .C2(n4608), .A(n4607), .B(n4606), .ZN(n4637)
         );
  OAI211_X1 U5054 ( .C1(n4613), .C2(n4612), .A(n4611), .B(n4610), .ZN(n4614)
         );
  INV_X1 U5055 ( .A(n4614), .ZN(n4627) );
  AOI22_X1 U5056 ( .A1(n4629), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4624) );
  MUX2_X1 U5057 ( .A(n4616), .B(REG1_REG_2__SCAN_IN), .S(n4615), .Z(n4619) );
  INV_X1 U5058 ( .A(n4617), .ZN(n4618) );
  NAND2_X1 U5059 ( .A1(n4619), .A2(n4618), .ZN(n4621) );
  OAI211_X1 U5060 ( .C1(n4622), .C2(n4621), .A(n4630), .B(n4620), .ZN(n4623)
         );
  OAI211_X1 U5061 ( .C1(n4643), .C2(n4625), .A(n4624), .B(n4623), .ZN(n4626)
         );
  OR3_X1 U5062 ( .A1(n4637), .A2(n4627), .A3(n4626), .ZN(U3242) );
  AOI21_X1 U5063 ( .B1(n4629), .B2(ADDR_REG_4__SCAN_IN), .A(n4628), .ZN(n4642)
         );
  OAI21_X1 U5064 ( .B1(REG1_REG_4__SCAN_IN), .B2(n4631), .A(n4630), .ZN(n4632)
         );
  INV_X1 U5065 ( .A(n4632), .ZN(n4640) );
  AOI211_X1 U5066 ( .C1(n4636), .C2(n4635), .A(n4634), .B(n4633), .ZN(n4638)
         );
  AOI211_X1 U5067 ( .C1(n4640), .C2(n4639), .A(n4638), .B(n4637), .ZN(n4641)
         );
  OAI211_X1 U5068 ( .C1(n2428), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3244)
         );
  INV_X1 U5069 ( .A(n4647), .ZN(n4655) );
  INV_X1 U5070 ( .A(n4644), .ZN(n4645) );
  NOR2_X1 U5071 ( .A1(n4674), .A2(n4645), .ZN(n4654) );
  NOR2_X1 U5072 ( .A1(n4769), .A2(n4909), .ZN(n4646) );
  OAI22_X1 U5073 ( .A1(n4647), .A2(n4646), .B1(n2604), .B2(n4906), .ZN(n4652)
         );
  AOI211_X1 U5074 ( .C1(n4705), .C2(n4655), .A(n4654), .B(n4652), .ZN(n4650)
         );
  AOI22_X1 U5075 ( .A1(n4915), .A2(n4650), .B1(n4648), .B2(n4913), .ZN(U3518)
         );
  INV_X1 U5076 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5077 ( .A1(n4919), .A2(n4650), .B1(n4649), .B2(n4916), .ZN(U3467)
         );
  INV_X1 U5078 ( .A(n4651), .ZN(n4653) );
  AOI21_X1 U5079 ( .B1(n4654), .B2(n4653), .A(n4652), .ZN(n4658) );
  AOI22_X1 U5080 ( .A1(n4655), .A2(n4776), .B1(REG3_REG_0__SCAN_IN), .B2(n4920), .ZN(n4656) );
  OAI221_X1 U5081 ( .B1(n4893), .B2(n4658), .C1(n4770), .C2(n4657), .A(n4656), 
        .ZN(U3290) );
  OAI21_X1 U5082 ( .B1(n4661), .B2(n4660), .A(n4659), .ZN(n4672) );
  AOI22_X1 U5083 ( .A1(n4663), .A2(n4903), .B1(n4662), .B2(n4902), .ZN(n4664)
         );
  OAI21_X1 U5084 ( .B1(n4665), .B2(n4906), .A(n4664), .ZN(n4671) );
  OAI21_X1 U5085 ( .B1(n4668), .B2(n4667), .A(n4666), .ZN(n4680) );
  NOR2_X1 U5086 ( .A1(n4680), .A2(n4669), .ZN(n4670) );
  AOI211_X1 U5087 ( .C1(n4909), .C2(n4672), .A(n4671), .B(n4670), .ZN(n4686)
         );
  INV_X1 U5088 ( .A(n4686), .ZN(n4677) );
  OAI21_X1 U5089 ( .B1(n4675), .B2(n4674), .A(n4673), .ZN(n4681) );
  OAI22_X1 U5090 ( .A1(n4680), .A2(n4792), .B1(n4898), .B2(n4681), .ZN(n4676)
         );
  NOR2_X1 U5091 ( .A1(n4677), .A2(n4676), .ZN(n4679) );
  AOI22_X1 U5092 ( .A1(n4915), .A2(n4679), .B1(n3842), .B2(n4913), .ZN(U3519)
         );
  INV_X1 U5093 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5094 ( .A1(n4919), .A2(n4679), .B1(n4678), .B2(n4916), .ZN(U3469)
         );
  AOI22_X1 U5095 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4920), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4893), .ZN(n4685) );
  INV_X1 U5096 ( .A(n4680), .ZN(n4683) );
  INV_X1 U5097 ( .A(n4681), .ZN(n4682) );
  AOI22_X1 U5098 ( .A1(n4683), .A2(n4776), .B1(n4981), .B2(n4682), .ZN(n4684)
         );
  OAI211_X1 U5099 ( .C1(n4893), .C2(n4686), .A(n4685), .B(n4684), .ZN(U3289)
         );
  AOI21_X1 U5100 ( .B1(n4705), .B2(n4688), .A(n4687), .ZN(n4694) );
  AOI22_X1 U5101 ( .A1(n4689), .A2(n4691), .B1(n4913), .B2(REG1_REG_2__SCAN_IN), .ZN(n4690) );
  OAI21_X1 U5102 ( .B1(n4694), .B2(n4913), .A(n4690), .ZN(U3520) );
  AOI22_X1 U5103 ( .A1(n4692), .A2(n4691), .B1(REG0_REG_2__SCAN_IN), .B2(n4916), .ZN(n4693) );
  OAI21_X1 U5104 ( .B1(n4694), .B2(n4916), .A(n4693), .ZN(U3471) );
  AOI22_X1 U5105 ( .A1(STATE_REG_SCAN_IN), .A2(n2927), .B1(n4695), .B2(U3149), 
        .ZN(U3349) );
  AOI22_X1 U5106 ( .A1(n4893), .A2(REG2_REG_3__SCAN_IN), .B1(n4920), .B2(n4696), .ZN(n4700) );
  AOI22_X1 U5107 ( .A1(n4698), .A2(n4776), .B1(n4981), .B2(n4697), .ZN(n4699)
         );
  OAI211_X1 U5108 ( .C1(n4893), .C2(n4701), .A(n4700), .B(n4699), .ZN(U3287)
         );
  AOI22_X1 U5109 ( .A1(STATE_REG_SCAN_IN), .A2(n2428), .B1(n4702), .B2(U3149), 
        .ZN(U3348) );
  AOI211_X1 U5110 ( .C1(n4706), .C2(n4705), .A(n4704), .B(n4703), .ZN(n4709)
         );
  INV_X1 U5111 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5112 ( .A1(n4915), .A2(n4709), .B1(n4707), .B2(n4913), .ZN(U3522)
         );
  INV_X1 U5113 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5114 ( .A1(n4919), .A2(n4709), .B1(n4708), .B2(n4916), .ZN(U3475)
         );
  INV_X1 U5115 ( .A(DATAI_6_), .ZN(n4710) );
  AOI22_X1 U5116 ( .A1(STATE_REG_SCAN_IN), .A2(n2342), .B1(n4710), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5117 ( .A1(n4711), .A2(n4920), .B1(REG2_REG_6__SCAN_IN), .B2(n4893), .ZN(n4717) );
  INV_X1 U5118 ( .A(n4712), .ZN(n4715) );
  INV_X1 U5119 ( .A(n4713), .ZN(n4714) );
  AOI22_X1 U5120 ( .A1(n4715), .A2(n4776), .B1(n4981), .B2(n4714), .ZN(n4716)
         );
  OAI211_X1 U5121 ( .C1(n4893), .C2(n4718), .A(n4717), .B(n4716), .ZN(U3284)
         );
  AOI22_X1 U5122 ( .A1(STATE_REG_SCAN_IN), .A2(n4720), .B1(n4719), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5123 ( .A(n4721), .ZN(n4722) );
  AOI211_X1 U5124 ( .C1(n4723), .C2(n4722), .A(n4898), .B(n2316), .ZN(n4742)
         );
  XOR2_X1 U5125 ( .A(n4734), .B(n4724), .Z(n4731) );
  OAI22_X1 U5126 ( .A1(n4727), .A2(n4726), .B1(n4725), .B2(n4862), .ZN(n4728)
         );
  AOI21_X1 U5127 ( .B1(n4869), .B2(n4729), .A(n4728), .ZN(n4730) );
  OAI21_X1 U5128 ( .B1(n4731), .B2(n4864), .A(n4730), .ZN(n4741) );
  AOI211_X1 U5129 ( .C1(n4732), .C2(n4742), .A(n4893), .B(n4741), .ZN(n4737)
         );
  XOR2_X1 U5130 ( .A(n4734), .B(n4733), .Z(n4743) );
  NAND2_X1 U5131 ( .A1(n4743), .A2(n4735), .ZN(n4736) );
  NAND2_X1 U5132 ( .A1(n4737), .A2(n4736), .ZN(n4738) );
  OAI21_X1 U5133 ( .B1(REG2_REG_7__SCAN_IN), .B2(n4770), .A(n4738), .ZN(n4739)
         );
  OAI21_X1 U5134 ( .B1(n4740), .B2(n4882), .A(n4739), .ZN(U3283) );
  AOI211_X1 U5135 ( .C1(n4743), .C2(n4912), .A(n4742), .B(n4741), .ZN(n4746)
         );
  AOI22_X1 U5136 ( .A1(n4915), .A2(n4746), .B1(n4744), .B2(n4913), .ZN(U3525)
         );
  INV_X1 U5137 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5138 ( .A1(n4919), .A2(n4746), .B1(n4745), .B2(n4916), .ZN(U3481)
         );
  AOI22_X1 U5139 ( .A1(STATE_REG_SCAN_IN), .A2(n4748), .B1(n4747), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5140 ( .A1(n4749), .A2(n4920), .B1(REG2_REG_8__SCAN_IN), .B2(n4893), .ZN(n4754) );
  INV_X1 U5141 ( .A(n4750), .ZN(n4751) );
  AOI22_X1 U5142 ( .A1(n4752), .A2(n4776), .B1(n4981), .B2(n4751), .ZN(n4753)
         );
  OAI211_X1 U5143 ( .C1(n4893), .C2(n4755), .A(n4754), .B(n4753), .ZN(U3282)
         );
  AOI22_X1 U5144 ( .A1(STATE_REG_SCAN_IN), .A2(n4757), .B1(n4756), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5145 ( .A(DATAI_10_), .ZN(n4758) );
  AOI22_X1 U5146 ( .A1(STATE_REG_SCAN_IN), .A2(n4759), .B1(n4758), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5147 ( .A1(n4760), .A2(n4920), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4893), .ZN(n4765) );
  INV_X1 U5148 ( .A(n4761), .ZN(n4762) );
  AOI22_X1 U5149 ( .A1(n4763), .A2(n4776), .B1(n4981), .B2(n4762), .ZN(n4764)
         );
  OAI211_X1 U5150 ( .C1(n4893), .C2(n4766), .A(n4765), .B(n4764), .ZN(U3280)
         );
  AOI22_X1 U5151 ( .A1(STATE_REG_SCAN_IN), .A2(n2940), .B1(n4767), .B2(U3149), 
        .ZN(U3341) );
  AOI21_X1 U5152 ( .B1(n4769), .B2(n4777), .A(n4768), .ZN(n4780) );
  OAI22_X1 U5153 ( .A1(n4772), .A2(n4882), .B1(n4771), .B2(n4770), .ZN(n4773)
         );
  INV_X1 U5154 ( .A(n4773), .ZN(n4779) );
  INV_X1 U5155 ( .A(n4774), .ZN(n4775) );
  AOI22_X1 U5156 ( .A1(n4777), .A2(n4776), .B1(n4981), .B2(n4775), .ZN(n4778)
         );
  OAI211_X1 U5157 ( .C1(n4893), .C2(n4780), .A(n4779), .B(n4778), .ZN(U3279)
         );
  AOI22_X1 U5158 ( .A1(STATE_REG_SCAN_IN), .A2(n4782), .B1(n4781), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5159 ( .A1(n4783), .A2(n4920), .B1(REG2_REG_12__SCAN_IN), .B2(
        n4893), .ZN(n4788) );
  INV_X1 U5160 ( .A(n4784), .ZN(n4785) );
  AOI22_X1 U5161 ( .A1(n4786), .A2(n4924), .B1(n4981), .B2(n4785), .ZN(n4787)
         );
  OAI211_X1 U5162 ( .C1(n4893), .C2(n4789), .A(n4788), .B(n4787), .ZN(U3278)
         );
  OAI22_X1 U5163 ( .A1(U3149), .A2(n4790), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4791) );
  INV_X1 U5164 ( .A(n4791), .ZN(U3339) );
  NOR2_X1 U5165 ( .A1(n4793), .A2(n4792), .ZN(n4795) );
  AOI211_X1 U5166 ( .C1(n4872), .C2(n4796), .A(n4795), .B(n4794), .ZN(n4799)
         );
  AOI22_X1 U5167 ( .A1(n4915), .A2(n4799), .B1(n4797), .B2(n4913), .ZN(U3531)
         );
  INV_X1 U5168 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5169 ( .A1(n4919), .A2(n4799), .B1(n4798), .B2(n4916), .ZN(U3493)
         );
  AOI22_X1 U5170 ( .A1(n4800), .A2(n4920), .B1(REG2_REG_14__SCAN_IN), .B2(
        n4893), .ZN(n4805) );
  INV_X1 U5171 ( .A(n4801), .ZN(n4802) );
  AOI22_X1 U5172 ( .A1(n4803), .A2(n4924), .B1(n4981), .B2(n4802), .ZN(n4804)
         );
  OAI211_X1 U5173 ( .C1(n4893), .C2(n4806), .A(n4805), .B(n4804), .ZN(U3276)
         );
  OAI22_X1 U5174 ( .A1(n4825), .A2(n4808), .B1(n4807), .B2(n4934), .ZN(n4809)
         );
  AOI211_X1 U5175 ( .C1(n4970), .C2(n4823), .A(n4810), .B(n4809), .ZN(n4817)
         );
  NAND2_X1 U5176 ( .A1(n4812), .A2(n4811), .ZN(n4813) );
  XOR2_X1 U5177 ( .A(n4814), .B(n4813), .Z(n4815) );
  NAND2_X1 U5178 ( .A1(n4815), .A2(n4974), .ZN(n4816) );
  OAI211_X1 U5179 ( .C1(n4979), .C2(n4818), .A(n4817), .B(n4816), .ZN(U3238)
         );
  NAND2_X1 U5180 ( .A1(n4820), .A2(n4819), .ZN(n4821) );
  XNOR2_X1 U5181 ( .A(n4821), .B(n4827), .ZN(n4838) );
  OAI21_X1 U5182 ( .B1(n4822), .B2(n4825), .A(n4854), .ZN(n4836) );
  NAND2_X1 U5183 ( .A1(n4823), .A2(n4903), .ZN(n4824) );
  OAI21_X1 U5184 ( .B1(n4825), .B2(n4862), .A(n4824), .ZN(n4829) );
  AOI211_X1 U5185 ( .C1(n4827), .C2(n4826), .A(n4864), .B(n2306), .ZN(n4828)
         );
  AOI211_X1 U5186 ( .C1(n4869), .C2(n4830), .A(n4829), .B(n4828), .ZN(n4841)
         );
  OAI21_X1 U5187 ( .B1(n4898), .B2(n4836), .A(n4841), .ZN(n4831) );
  AOI21_X1 U5188 ( .B1(n4912), .B2(n4838), .A(n4831), .ZN(n4834) );
  AOI22_X1 U5189 ( .A1(n4915), .A2(n4834), .B1(n4832), .B2(n4913), .ZN(U3533)
         );
  INV_X1 U5190 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5191 ( .A1(n4919), .A2(n4834), .B1(n4833), .B2(n4916), .ZN(U3497)
         );
  AOI22_X1 U5192 ( .A1(n4835), .A2(n4920), .B1(REG2_REG_15__SCAN_IN), .B2(
        n4893), .ZN(n4840) );
  INV_X1 U5193 ( .A(n4836), .ZN(n4837) );
  AOI22_X1 U5194 ( .A1(n4838), .A2(n4924), .B1(n4981), .B2(n4837), .ZN(n4839)
         );
  OAI211_X1 U5195 ( .C1(n4893), .C2(n4841), .A(n4840), .B(n4839), .ZN(U3275)
         );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4843), .B1(n4842), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5197 ( .A(n4875), .ZN(n4852) );
  AOI22_X1 U5198 ( .A1(n4964), .A2(n4904), .B1(n4973), .B2(n4855), .ZN(n4851)
         );
  XOR2_X1 U5199 ( .A(n4845), .B(n4844), .Z(n4847) );
  NOR2_X1 U5200 ( .A1(n4847), .A2(n4846), .ZN(n4848) );
  AOI211_X1 U5201 ( .C1(n4970), .C2(n4859), .A(n4849), .B(n4848), .ZN(n4850)
         );
  OAI211_X1 U5202 ( .C1(n4979), .C2(n4852), .A(n4851), .B(n4850), .ZN(U3223)
         );
  AOI21_X1 U5203 ( .B1(n4855), .B2(n4854), .A(n4853), .ZN(n4877) );
  OAI21_X1 U5204 ( .B1(n4857), .B2(n4865), .A(n4856), .ZN(n4876) );
  NOR2_X1 U5205 ( .A1(n4876), .A2(n4858), .ZN(n4871) );
  NAND2_X1 U5206 ( .A1(n4859), .A2(n4903), .ZN(n4860) );
  OAI21_X1 U5207 ( .B1(n4862), .B2(n4861), .A(n4860), .ZN(n4868) );
  AOI211_X1 U5208 ( .C1(n4866), .C2(n4865), .A(n4864), .B(n4863), .ZN(n4867)
         );
  AOI211_X1 U5209 ( .C1(n4869), .C2(n4904), .A(n4868), .B(n4867), .ZN(n4881)
         );
  INV_X1 U5210 ( .A(n4881), .ZN(n4870) );
  AOI211_X1 U5211 ( .C1(n4872), .C2(n4877), .A(n4871), .B(n4870), .ZN(n4874)
         );
  AOI22_X1 U5212 ( .A1(n4915), .A2(n4874), .B1(n2431), .B2(n4913), .ZN(U3534)
         );
  INV_X1 U5213 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4873) );
  AOI22_X1 U5214 ( .A1(n4919), .A2(n4874), .B1(n4873), .B2(n4916), .ZN(U3499)
         );
  AOI22_X1 U5215 ( .A1(n4875), .A2(n4920), .B1(REG2_REG_16__SCAN_IN), .B2(
        n4893), .ZN(n4880) );
  INV_X1 U5216 ( .A(n4876), .ZN(n4878) );
  AOI22_X1 U5217 ( .A1(n4878), .A2(n4924), .B1(n4981), .B2(n4877), .ZN(n4879)
         );
  OAI211_X1 U5218 ( .C1(n4893), .C2(n4881), .A(n4880), .B(n4879), .ZN(U3274)
         );
  NOR2_X1 U5219 ( .A1(n4883), .A2(n4882), .ZN(n4890) );
  INV_X1 U5220 ( .A(n4884), .ZN(n4888) );
  OAI22_X1 U5221 ( .A1(n4888), .A2(n4887), .B1(n4886), .B2(n4885), .ZN(n4889)
         );
  AOI211_X1 U5222 ( .C1(n4893), .C2(REG2_REG_17__SCAN_IN), .A(n4890), .B(n4889), .ZN(n4891) );
  OAI21_X1 U5223 ( .B1(n4893), .B2(n4892), .A(n4891), .ZN(U3273) );
  INV_X1 U5224 ( .A(n4899), .ZN(n4895) );
  OAI21_X1 U5225 ( .B1(n4896), .B2(n4895), .A(n4894), .ZN(n4925) );
  AOI211_X1 U5226 ( .C1(n4901), .C2(n2298), .A(n4898), .B(n4897), .ZN(n4922)
         );
  XNOR2_X1 U5227 ( .A(n4900), .B(n4899), .ZN(n4910) );
  AOI22_X1 U5228 ( .A1(n4904), .A2(n4903), .B1(n4902), .B2(n4901), .ZN(n4905)
         );
  OAI21_X1 U5229 ( .B1(n4907), .B2(n4906), .A(n4905), .ZN(n4908) );
  AOI21_X1 U5230 ( .B1(n4910), .B2(n4909), .A(n4908), .ZN(n4928) );
  INV_X1 U5231 ( .A(n4928), .ZN(n4911) );
  AOI211_X1 U5232 ( .C1(n4912), .C2(n4925), .A(n4922), .B(n4911), .ZN(n4918)
         );
  AOI22_X1 U5233 ( .A1(n4915), .A2(n4918), .B1(n4914), .B2(n4913), .ZN(U3536)
         );
  INV_X1 U5234 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4917) );
  AOI22_X1 U5235 ( .A1(n4919), .A2(n4918), .B1(n4917), .B2(n4916), .ZN(U3503)
         );
  AOI22_X1 U5236 ( .A1(n4921), .A2(n4920), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4893), .ZN(n4927) );
  AOI22_X1 U5237 ( .A1(n4925), .A2(n4924), .B1(n4923), .B2(n4922), .ZN(n4926)
         );
  OAI211_X1 U5238 ( .C1(n4893), .C2(n4928), .A(n4927), .B(n4926), .ZN(U3272)
         );
  AOI22_X1 U5239 ( .A1(n4970), .A2(n4930), .B1(n4973), .B2(n4929), .ZN(n4940)
         );
  OAI21_X1 U5240 ( .B1(n4933), .B2(n4932), .A(n4931), .ZN(n4938) );
  INV_X1 U5241 ( .A(n4957), .ZN(n4935) );
  NOR2_X1 U5242 ( .A1(n4935), .A2(n4934), .ZN(n4937) );
  AOI211_X1 U5243 ( .C1(n4938), .C2(n4974), .A(n4937), .B(n4936), .ZN(n4939)
         );
  OAI211_X1 U5244 ( .C1(n4979), .C2(n4941), .A(n4940), .B(n4939), .ZN(U3216)
         );
  AOI22_X1 U5245 ( .A1(n4964), .A2(n4971), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4947) );
  NAND2_X1 U5246 ( .A1(n4951), .A2(n4950), .ZN(n4942) );
  XOR2_X1 U5247 ( .A(n4942), .B(n4953), .Z(n4944) );
  AOI222_X1 U5248 ( .A1(n4973), .A2(n4945), .B1(n4974), .B2(n4944), .C1(n4943), 
        .C2(n4970), .ZN(n4946) );
  OAI211_X1 U5249 ( .C1(n4979), .C2(n4948), .A(n4947), .B(n4946), .ZN(U3230)
         );
  AOI22_X1 U5250 ( .A1(n4964), .A2(n4949), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4961) );
  INV_X1 U5251 ( .A(n4950), .ZN(n4952) );
  OAI21_X1 U5252 ( .B1(n4953), .B2(n4952), .A(n4951), .ZN(n4956) );
  NAND2_X1 U5253 ( .A1(n4965), .A2(n4954), .ZN(n4955) );
  XNOR2_X1 U5254 ( .A(n4956), .B(n4955), .ZN(n4959) );
  AOI222_X1 U5255 ( .A1(n4959), .A2(n4974), .B1(n4973), .B2(n4958), .C1(n4957), 
        .C2(n4970), .ZN(n4960) );
  OAI211_X1 U5256 ( .C1(n4979), .C2(n4962), .A(n4961), .B(n4960), .ZN(U3220)
         );
  AOI22_X1 U5257 ( .A1(n4964), .A2(n4963), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n4977) );
  AND2_X1 U5258 ( .A1(n4966), .A2(n4965), .ZN(n4969) );
  OAI21_X1 U5259 ( .B1(n4969), .B2(n4968), .A(n4967), .ZN(n4975) );
  AOI222_X1 U5260 ( .A1(n4975), .A2(n4974), .B1(n4973), .B2(n4972), .C1(n4971), 
        .C2(n4970), .ZN(n4976) );
  OAI211_X1 U5261 ( .C1(n4979), .C2(n4978), .A(n4977), .B(n4976), .ZN(U3232)
         );
  INV_X1 U5262 ( .A(n4980), .ZN(n4984) );
  AOI22_X1 U5263 ( .A1(n4982), .A2(n4981), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4893), .ZN(n4983) );
  OAI21_X1 U5264 ( .B1(n4893), .B2(n4984), .A(n4983), .ZN(U3261) );
  INV_X1 U2301 ( .A(n3557), .ZN(n3545) );
endmodule

