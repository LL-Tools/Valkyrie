

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6405, n6406, n6407, n6409, n6410, n6411, n6412, n6413, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6424, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15375;

  NAND2_X1 U7152 ( .A1(n13053), .A2(n11967), .ZN(n13122) );
  NAND2_X1 U7153 ( .A1(n7121), .A2(n6444), .ZN(n13049) );
  INV_X4 U7154 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OR2_X1 U7155 ( .A1(n14132), .A2(n14140), .ZN(n14130) );
  NAND2_X1 U7156 ( .A1(n14129), .A2(n13982), .ZN(n14113) );
  NAND2_X1 U7157 ( .A1(n7118), .A2(n6442), .ZN(n13030) );
  NAND2_X1 U7158 ( .A1(n13491), .A2(n13503), .ZN(n13490) );
  OAI21_X1 U7159 ( .B1(n10705), .B2(n10704), .A(n11998), .ZN(n10706) );
  CLKBUF_X2 U7160 ( .A(n10254), .Z(n12122) );
  INV_X2 U7162 ( .A(n8455), .ZN(n9005) );
  NAND2_X2 U7163 ( .A1(n9560), .A2(n11541), .ZN(n12047) );
  NAND2_X1 U7164 ( .A1(n8626), .A2(n8625), .ZN(n8652) );
  BUF_X1 U7165 ( .A(n8360), .Z(n8980) );
  AND2_X1 U7167 ( .A1(n8299), .A2(n8348), .ZN(n8360) );
  BUF_X4 U7168 ( .A(n11713), .Z(n6412) );
  INV_X1 U7169 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9639) );
  INV_X1 U7171 ( .A(n15375), .ZN(n6405) );
  AOI21_X1 U7172 ( .B1(n14030), .B2(n14039), .A(n13990), .ZN(n14017) );
  NAND2_X1 U7173 ( .A1(n10342), .A2(n10341), .ZN(n10886) );
  OR2_X1 U7174 ( .A1(n8320), .A2(n13671), .ZN(n8322) );
  AOI21_X1 U7175 ( .B1(n6950), .B2(n6952), .A(n6543), .ZN(n6947) );
  INV_X1 U7176 ( .A(n9090), .ZN(n8771) );
  INV_X1 U7177 ( .A(n9007), .ZN(n8772) );
  INV_X1 U7178 ( .A(n9563), .ZN(n12129) );
  OR2_X1 U7180 ( .A1(n15100), .A2(n15099), .ZN(n15102) );
  OR2_X1 U7181 ( .A1(n12585), .A2(n12584), .ZN(n12613) );
  NAND2_X2 U7182 ( .A1(n8140), .A2(n6412), .ZN(n12299) );
  INV_X1 U7183 ( .A(n11101), .ZN(n11972) );
  CLKBUF_X3 U7184 ( .A(n8411), .Z(n6409) );
  AND2_X1 U7185 ( .A1(n7031), .A2(n10538), .ZN(n10717) );
  NAND2_X1 U7186 ( .A1(n13490), .A2(n7547), .ZN(n13478) );
  INV_X1 U7187 ( .A(n10541), .ZN(n14995) );
  BUF_X1 U7189 ( .A(n8306), .Z(n8679) );
  INV_X1 U7190 ( .A(n6411), .ZN(n7606) );
  OAI211_X2 U7191 ( .C1(n9090), .C2(n13151), .A(n8333), .B(n8332), .ZN(n9053)
         );
  INV_X1 U7192 ( .A(n8360), .ZN(n9012) );
  CLKBUF_X2 U7193 ( .A(n8389), .Z(n9017) );
  INV_X1 U7194 ( .A(n10369), .ZN(n8318) );
  NAND2_X1 U7195 ( .A1(n11776), .A2(n11775), .ZN(n14038) );
  NAND2_X1 U7196 ( .A1(n9222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9223) );
  INV_X1 U7197 ( .A(n8348), .ZN(n13676) );
  XNOR2_X1 U7198 ( .A(n9223), .B(n9122), .ZN(n11870) );
  INV_X1 U7199 ( .A(n12521), .ZN(P3_U3897) );
  XNOR2_X1 U7200 ( .A(n8322), .B(n8321), .ZN(n9093) );
  AND2_X1 U7201 ( .A1(n7241), .A2(n13294), .ZN(n6406) );
  OR2_X1 U7202 ( .A1(n12142), .A2(n15179), .ZN(n8242) );
  OR2_X2 U7203 ( .A1(n10891), .A2(n6939), .ZN(n6938) );
  INV_X2 U7204 ( .A(n11541), .ZN(n11863) );
  AND2_X2 U7205 ( .A1(n6800), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14380) );
  INV_X1 U7206 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U7207 ( .A1(n9093), .A2(n9094), .ZN(n6407) );
  NAND2_X2 U7208 ( .A1(n9093), .A2(n9094), .ZN(n9090) );
  INV_X2 U7209 ( .A(n8126), .ZN(n11019) );
  AOI21_X2 U7210 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8396) );
  XNOR2_X2 U7211 ( .A(n8372), .B(SI_1_), .ZN(n8375) );
  OAI21_X2 U7212 ( .B1(n8679), .B2(n7136), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8311) );
  BUF_X2 U7214 ( .A(n8411), .Z(n6410) );
  OAI222_X1 U7216 ( .A1(n13686), .A2(n12000), .B1(P2_U3088), .B2(n8299), .C1(
        n13688), .C2(n11999), .ZN(P2_U3297) );
  NOR2_X2 U7217 ( .A1(n10027), .A2(n15190), .ZN(n10026) );
  NAND2_X2 U7218 ( .A1(n6973), .A2(n9780), .ZN(n10027) );
  BUF_X8 U7219 ( .A(n11713), .Z(n6411) );
  INV_X4 U7220 ( .A(n8330), .ZN(n11713) );
  OAI211_X2 U7221 ( .C1(n12299), .C2(SI_9_), .A(n7760), .B(n7759), .ZN(n12391)
         );
  CLKBUF_X2 U7222 ( .A(n13145), .Z(n6413) );
  NAND2_X1 U7223 ( .A1(n8305), .A2(n8304), .ZN(n13145) );
  XNOR2_X2 U7224 ( .A(n9125), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9262) );
  CLKBUF_X1 U7226 ( .A(n14653), .Z(n6415) );
  XNOR2_X1 U7227 ( .A(n9233), .B(n9232), .ZN(n14653) );
  BUF_X1 U7229 ( .A(n9811), .Z(n6417) );
  CLKBUF_X1 U7230 ( .A(n9811), .Z(n6418) );
  XNOR2_X1 U7231 ( .A(n7596), .B(n7598), .ZN(n9811) );
  AND2_X2 U7232 ( .A1(n12617), .A2(n12616), .ZN(n12640) );
  INV_X2 U7233 ( .A(n10946), .ZN(n9649) );
  NAND2_X2 U7234 ( .A1(n8315), .A2(n9087), .ZN(n10946) );
  AOI21_X2 U7235 ( .B1(n6953), .B2(n6955), .A(n6951), .ZN(n6950) );
  XNOR2_X2 U7236 ( .A(n13836), .B(n11542), .ZN(n11877) );
  NAND2_X1 U7237 ( .A1(n7112), .A2(n7111), .ZN(n13019) );
  INV_X1 U7238 ( .A(n7648), .ZN(n7561) );
  NAND2_X2 U7240 ( .A1(n7568), .A2(n6458), .ZN(n8101) );
  NAND3_X2 U7241 ( .A1(n6688), .A2(n6691), .A3(n7632), .ZN(n6689) );
  NOR2_X2 U7242 ( .A1(n12615), .A2(n12614), .ZN(n12636) );
  XNOR2_X2 U7243 ( .A(n12635), .B(n12641), .ZN(n12614) );
  NOR2_X2 U7244 ( .A1(n15369), .A2(n14384), .ZN(n14437) );
  XNOR2_X2 U7245 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14379) );
  XNOR2_X2 U7246 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14375), .ZN(n14387) );
  NAND2_X2 U7247 ( .A1(n9829), .A2(n10035), .ZN(n9850) );
  NOR2_X1 U7248 ( .A1(n14847), .A2(n14463), .ZN(n14462) );
  AOI211_X2 U7249 ( .C1(n15106), .C2(n12641), .A(n12632), .B(n12631), .ZN(
        n12633) );
  OR2_X1 U7250 ( .A1(n12710), .A2(n12713), .ZN(n7415) );
  CLKBUF_X2 U7251 ( .A(n13582), .Z(n6879) );
  NAND2_X1 U7252 ( .A1(n6808), .A2(n11743), .ZN(n14073) );
  OAI21_X1 U7253 ( .B1(n12845), .B2(n7281), .A(n7278), .ZN(n12818) );
  NAND2_X1 U7254 ( .A1(n13975), .A2(n13974), .ZN(n14582) );
  NAND2_X1 U7255 ( .A1(n6703), .A2(n12408), .ZN(n11278) );
  NAND2_X1 U7256 ( .A1(n11634), .A2(n11633), .ZN(n14303) );
  NOR2_X1 U7257 ( .A1(n11319), .A2(n11318), .ZN(n12534) );
  OAI21_X1 U7258 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(n10902) );
  NAND2_X1 U7259 ( .A1(n12341), .A2(n12351), .ZN(n8225) );
  NOR2_X1 U7260 ( .A1(n13527), .A2(n10621), .ZN(n10616) );
  INV_X1 U7261 ( .A(n15001), .ZN(n7032) );
  OR2_X1 U7262 ( .A1(n9784), .A2(n9783), .ZN(n10165) );
  OAI211_X1 U7263 ( .C1(n8455), .C2(n9930), .A(n8426), .B(n6490), .ZN(n10541)
         );
  AND3_X2 U7264 ( .A1(n7243), .A2(n8377), .A3(n6483), .ZN(n9052) );
  INV_X4 U7265 ( .A(n11844), .ZN(n11867) );
  INV_X1 U7266 ( .A(n8842), .ZN(n6420) );
  INV_X4 U7267 ( .A(n8842), .ZN(n9046) );
  NOR2_X1 U7268 ( .A1(n10856), .A2(n15161), .ZN(n12357) );
  OR2_X1 U7269 ( .A1(n9053), .A2(n13530), .ZN(n13527) );
  INV_X2 U7270 ( .A(n11542), .ZN(n11552) );
  INV_X4 U7271 ( .A(n11574), .ZN(n11844) );
  INV_X1 U7272 ( .A(n13834), .ZN(n10253) );
  INV_X1 U7273 ( .A(n13833), .ZN(n6845) );
  NAND3_X4 U7274 ( .A1(n9560), .A2(n11863), .A3(n14718), .ZN(n10184) );
  AND2_X1 U7276 ( .A1(n7619), .A2(n7620), .ZN(n7634) );
  NAND3_X2 U7277 ( .A1(n9262), .A2(n9258), .A3(n14320), .ZN(n9560) );
  INV_X1 U7278 ( .A(n9925), .ZN(n10072) );
  INV_X2 U7279 ( .A(n11715), .ZN(n11659) );
  NAND2_X2 U7280 ( .A1(n11531), .A2(n14314), .ZN(n9944) );
  INV_X2 U7281 ( .A(n9796), .ZN(n12675) );
  INV_X2 U7282 ( .A(n9276), .ZN(n14314) );
  NAND2_X1 U7283 ( .A1(n7013), .A2(n7011), .ZN(n14331) );
  NAND2_X1 U7284 ( .A1(n6411), .A2(P3_U3151), .ZN(n12997) );
  NAND2_X1 U7285 ( .A1(n6881), .A2(n6880), .ZN(n7649) );
  NAND4_X1 U7286 ( .A1(n8284), .A2(n8417), .A3(n8288), .A4(n7454), .ZN(n8306)
         );
  NOR2_X1 U7287 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9113) );
  INV_X2 U7288 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U7289 ( .A1(n6669), .A2(n9049), .ZN(n9106) );
  NAND2_X2 U7290 ( .A1(n12270), .A2(n12271), .ZN(n12269) );
  NAND2_X1 U7291 ( .A1(n12148), .A2(n8242), .ZN(n8274) );
  AOI21_X1 U7292 ( .B1(n12895), .B2(n15141), .A(n12716), .ZN(n12717) );
  NAND2_X1 U7293 ( .A1(n6768), .A2(n13496), .ZN(n13549) );
  NAND2_X1 U7294 ( .A1(n8018), .A2(n8026), .ZN(n7340) );
  OAI21_X1 U7295 ( .B1(n14048), .B2(n7153), .A(n6431), .ZN(n13997) );
  OAI21_X1 U7296 ( .B1(n12713), .B2(n6467), .A(n12712), .ZN(n12895) );
  OAI21_X1 U7297 ( .B1(n12711), .B2(n12484), .A(n12482), .ZN(n12496) );
  OR2_X1 U7298 ( .A1(n8786), .A2(n8785), .ZN(n8802) );
  AOI21_X1 U7299 ( .B1(n7058), .B2(n7057), .A(n6538), .ZN(n7056) );
  AND2_X1 U7300 ( .A1(n7068), .A2(n13313), .ZN(n13396) );
  INV_X1 U7301 ( .A(n14202), .ZN(n6419) );
  NAND2_X1 U7302 ( .A1(n14066), .A2(n14065), .ZN(n14064) );
  NAND2_X1 U7303 ( .A1(n7123), .A2(n11955), .ZN(n13074) );
  AND2_X1 U7304 ( .A1(n6976), .A2(n7190), .ZN(n6804) );
  NAND2_X1 U7305 ( .A1(n8979), .A2(n8978), .ZN(n13558) );
  NAND2_X2 U7306 ( .A1(n11808), .A2(n11807), .ZN(n14205) );
  NAND2_X1 U7307 ( .A1(n7125), .A2(n7126), .ZN(n13097) );
  NAND2_X2 U7308 ( .A1(n11793), .A2(n11792), .ZN(n14026) );
  NAND2_X2 U7309 ( .A1(n9009), .A2(n9008), .ZN(n13568) );
  OR2_X1 U7310 ( .A1(n8724), .A2(n7460), .ZN(n6640) );
  XNOR2_X1 U7311 ( .A(n8976), .B(n8975), .ZN(n13678) );
  XNOR2_X1 U7312 ( .A(n9004), .B(n9003), .ZN(n13681) );
  XNOR2_X1 U7313 ( .A(n13582), .B(n13284), .ZN(n13379) );
  NAND2_X1 U7314 ( .A1(n12747), .A2(n12465), .ZN(n12751) );
  NAND2_X1 U7315 ( .A1(n13308), .A2(n6767), .ZN(n13438) );
  NAND2_X1 U7316 ( .A1(n11757), .A2(n11756), .ZN(n14220) );
  NAND2_X1 U7317 ( .A1(n12766), .A2(n7544), .ZN(n12747) );
  NAND2_X1 U7318 ( .A1(n7391), .A2(n7393), .ZN(n9004) );
  NAND2_X1 U7319 ( .A1(n14643), .A2(n14645), .ZN(n14650) );
  NAND2_X1 U7320 ( .A1(n6677), .A2(n6499), .ZN(n12766) );
  NAND2_X1 U7321 ( .A1(n8070), .A2(n8069), .ZN(n8238) );
  NAND2_X2 U7322 ( .A1(n8871), .A2(n8870), .ZN(n13587) );
  NAND2_X1 U7323 ( .A1(n7392), .A2(n7398), .ZN(n7391) );
  NAND2_X1 U7324 ( .A1(n11741), .A2(n9005), .ZN(n8871) );
  NAND2_X1 U7325 ( .A1(n6777), .A2(n6776), .ZN(n14645) );
  INV_X1 U7326 ( .A(n14422), .ZN(n6777) );
  OAI21_X1 U7327 ( .B1(n12789), .B2(n12454), .A(n12317), .ZN(n12779) );
  AND2_X1 U7328 ( .A1(n14325), .A2(n11715), .ZN(n13986) );
  NAND2_X1 U7329 ( .A1(n12863), .A2(n12429), .ZN(n12845) );
  NAND2_X1 U7330 ( .A1(n8852), .A2(n8851), .ZN(n13410) );
  NAND2_X1 U7331 ( .A1(n6908), .A2(n6907), .ZN(n12211) );
  NAND2_X1 U7332 ( .A1(n12878), .A2(n12877), .ZN(n12876) );
  NAND2_X1 U7333 ( .A1(n7052), .A2(n7051), .ZN(n13298) );
  NAND2_X1 U7334 ( .A1(n6849), .A2(n8849), .ZN(n8866) );
  OAI21_X1 U7335 ( .B1(n14582), .B2(n13976), .A(n13977), .ZN(n14158) );
  XNOR2_X1 U7336 ( .A(n12046), .B(n12045), .ZN(n13812) );
  NAND2_X1 U7337 ( .A1(n6799), .A2(n6798), .ZN(n6834) );
  NAND2_X1 U7338 ( .A1(n11698), .A2(n11697), .ZN(n14292) );
  OAI21_X1 U7339 ( .B1(n11278), .B2(n8231), .A(n12413), .ZN(n11401) );
  NAND2_X1 U7340 ( .A1(n7326), .A2(n7325), .ZN(n12241) );
  NAND2_X1 U7341 ( .A1(n15118), .A2(n11328), .ZN(n6760) );
  NAND2_X1 U7342 ( .A1(n8829), .A2(n6574), .ZN(n7370) );
  NAND2_X1 U7343 ( .A1(n13776), .A2(n13775), .ZN(n14542) );
  INV_X1 U7344 ( .A(n14421), .ZN(n6776) );
  NAND2_X1 U7345 ( .A1(n6988), .A2(n6987), .ZN(n15118) );
  NAND2_X1 U7346 ( .A1(n8826), .A2(n8825), .ZN(n8829) );
  NAND3_X1 U7347 ( .A1(n6941), .A2(n6940), .A3(n6938), .ZN(n10893) );
  NOR2_X1 U7348 ( .A1(n15044), .A2(n7108), .ZN(n7107) );
  NOR2_X1 U7349 ( .A1(n15037), .A2(n7108), .ZN(n7106) );
  NOR2_X1 U7350 ( .A1(n11207), .A2(n11208), .ZN(n11206) );
  NAND2_X1 U7351 ( .A1(n7185), .A2(n6501), .ZN(n10891) );
  OAI211_X1 U7352 ( .C1(n6666), .C2(n6629), .A(n6525), .B(n6628), .ZN(n6630)
         );
  NAND2_X1 U7353 ( .A1(n11149), .A2(n11148), .ZN(n14606) );
  NAND2_X1 U7354 ( .A1(n10742), .A2(n10741), .ZN(n10744) );
  XNOR2_X1 U7355 ( .A(n10886), .B(n14443), .ZN(n10343) );
  NAND2_X1 U7356 ( .A1(n14459), .A2(n14405), .ZN(n14406) );
  NAND2_X1 U7357 ( .A1(n10516), .A2(n10515), .ZN(n10785) );
  NAND2_X1 U7358 ( .A1(n10597), .A2(n10596), .ZN(n10966) );
  NAND2_X1 U7359 ( .A1(n7193), .A2(n7192), .ZN(n10342) );
  OAI21_X1 U7360 ( .B1(n13738), .B2(n13736), .A(n13734), .ZN(n10516) );
  OAI21_X1 U7361 ( .B1(n6736), .B2(n6735), .A(n6733), .ZN(n7092) );
  NOR2_X1 U7362 ( .A1(n9835), .A2(n9836), .ZN(n9895) );
  NAND2_X1 U7363 ( .A1(n6805), .A2(n6492), .ZN(n6986) );
  AOI21_X1 U7364 ( .B1(n10902), .B2(n10901), .A(n10900), .ZN(n15109) );
  NAND2_X1 U7365 ( .A1(n10536), .A2(n10544), .ZN(n10535) );
  OAI22_X1 U7366 ( .A1(n8407), .A2(n6636), .B1(n8406), .B2(n8405), .ZN(n8433)
         );
  NAND2_X1 U7367 ( .A1(n10576), .A2(n10575), .ZN(n11609) );
  NAND2_X1 U7368 ( .A1(n6761), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U7369 ( .A1(n6930), .A2(n9834), .ZN(n6929) );
  NAND2_X1 U7370 ( .A1(n10071), .A2(n10070), .ZN(n10125) );
  CLKBUF_X1 U7371 ( .A(n13543), .Z(n14941) );
  NAND2_X1 U7372 ( .A1(n7187), .A2(n7186), .ZN(n6930) );
  NAND2_X1 U7373 ( .A1(n8541), .A2(n8540), .ZN(n15038) );
  NAND2_X1 U7374 ( .A1(n9729), .A2(n9730), .ZN(n10191) );
  CLKBUF_X1 U7375 ( .A(n8558), .Z(n6784) );
  AND2_X1 U7376 ( .A1(n10842), .A2(n8177), .ZN(n7431) );
  NAND2_X1 U7377 ( .A1(n8498), .A2(n8497), .ZN(n15020) );
  NAND2_X1 U7378 ( .A1(n8513), .A2(n8512), .ZN(n15029) );
  NAND2_X1 U7379 ( .A1(n14979), .A2(n9754), .ZN(n14938) );
  NAND2_X2 U7380 ( .A1(n9909), .A2(n14698), .ZN(n14700) );
  INV_X1 U7381 ( .A(n13540), .ZN(n13538) );
  CLKBUF_X3 U7382 ( .A(n7654), .Z(n7851) );
  BUF_X4 U7383 ( .A(n8842), .Z(n6426) );
  NAND2_X1 U7384 ( .A1(n9832), .A2(n9831), .ZN(n7543) );
  INV_X1 U7385 ( .A(n11976), .ZN(n11101) );
  OAI22_X1 U7386 ( .A1(n9817), .A2(n9844), .B1(n9816), .B2(n9830), .ZN(n10162)
         );
  AND2_X1 U7387 ( .A1(n9782), .A2(n10163), .ZN(n9784) );
  NAND4_X1 U7388 ( .A1(n8366), .A2(n8365), .A3(n8364), .A4(n8363), .ZN(n13144)
         );
  NAND4_X1 U7389 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n13143)
         );
  NAND3_X1 U7390 ( .A1(n7644), .A2(n6773), .A3(n7645), .ZN(n15144) );
  BUF_X1 U7391 ( .A(n8167), .Z(n12349) );
  NAND4_X2 U7392 ( .A1(n7661), .A2(n7660), .A3(n7659), .A4(n7658), .ZN(n10856)
         );
  INV_X4 U7393 ( .A(n10184), .ZN(n9562) );
  AOI21_X1 U7394 ( .B1(n9424), .B2(n15345), .A(n6529), .ZN(n12987) );
  XNOR2_X1 U7395 ( .A(n14338), .B(n7024), .ZN(n14389) );
  INV_X2 U7396 ( .A(n8361), .ZN(n9010) );
  INV_X1 U7397 ( .A(n8100), .ZN(n12014) );
  NAND2_X1 U7398 ( .A1(n7025), .A2(n14337), .ZN(n14338) );
  AND4_X2 U7399 ( .A1(n9615), .A2(n9612), .A3(n9613), .A4(n9614), .ZN(n10185)
         );
  NAND2_X1 U7400 ( .A1(n7464), .A2(n7462), .ZN(n13838) );
  AND2_X1 U7401 ( .A1(n7572), .A2(n7571), .ZN(n8100) );
  AND2_X2 U7402 ( .A1(n11529), .A2(n7619), .ZN(n6457) );
  XNOR2_X1 U7403 ( .A(n7587), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12687) );
  INV_X1 U7404 ( .A(n10163), .ZN(n9831) );
  OR2_X1 U7405 ( .A1(n9779), .A2(n10035), .ZN(n6973) );
  INV_X1 U7406 ( .A(n6698), .ZN(n7619) );
  INV_X1 U7407 ( .A(n11532), .ZN(n9258) );
  INV_X1 U7408 ( .A(n7620), .ZN(n11529) );
  MUX2_X1 U7409 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8314), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8315) );
  OR2_X1 U7410 ( .A1(n7675), .A2(n7674), .ZN(n10163) );
  AND2_X1 U7411 ( .A1(n7594), .A2(n7593), .ZN(n9860) );
  XNOR2_X1 U7412 ( .A(n6899), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7620) );
  XNOR2_X1 U7413 ( .A(n9124), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14320) );
  OR2_X1 U7414 ( .A1(n6827), .A2(n9159), .ZN(n9125) );
  XNOR2_X1 U7415 ( .A(n9236), .B(P1_IR_REG_20__SCAN_IN), .ZN(n11869) );
  XNOR2_X1 U7416 ( .A(n9221), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14326) );
  NOR2_X1 U7417 ( .A1(n6460), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9075) );
  OR2_X1 U7418 ( .A1(n7803), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U7419 ( .A1(n8296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8297) );
  BUF_X1 U7420 ( .A(n14317), .Z(n6424) );
  INV_X2 U7421 ( .A(n14310), .ZN(n11530) );
  XNOR2_X1 U7422 ( .A(n14331), .B(n7010), .ZN(n14376) );
  AOI21_X1 U7423 ( .B1(n7095), .B2(n7097), .A(n7094), .ZN(n7093) );
  XNOR2_X1 U7424 ( .A(n8474), .B(SI_5_), .ZN(n8471) );
  OAI21_X1 U7425 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9245) );
  NOR2_X1 U7426 ( .A1(n9220), .A2(n7527), .ZN(n6827) );
  MUX2_X1 U7427 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7602), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7605) );
  NAND2_X1 U7428 ( .A1(n12989), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U7429 ( .B1(n9220), .B2(n7528), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9124) );
  NAND2_X1 U7430 ( .A1(n6821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9233) );
  AND2_X2 U7431 ( .A1(n7648), .A2(n7183), .ZN(n10005) );
  NOR2_X1 U7432 ( .A1(n7591), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7673) );
  INV_X2 U7433 ( .A(n9207), .ZN(n6421) );
  NAND2_X1 U7434 ( .A1(n9235), .A2(n6709), .ZN(n9220) );
  NOR2_X1 U7435 ( .A1(n6465), .A2(n7456), .ZN(n7455) );
  AND2_X1 U7436 ( .A1(n9157), .A2(n9160), .ZN(n9237) );
  INV_X1 U7437 ( .A(n7649), .ZN(n7183) );
  INV_X1 U7438 ( .A(n8306), .ZN(n8292) );
  AND2_X1 U7439 ( .A1(n9120), .A2(n9157), .ZN(n9235) );
  NAND2_X1 U7440 ( .A1(n7530), .A2(n6498), .ZN(n7528) );
  NAND2_X2 U7441 ( .A1(n7626), .A2(n7627), .ZN(n10050) );
  INV_X1 U7443 ( .A(n7918), .ZN(n7094) );
  AND3_X1 U7444 ( .A1(n6687), .A2(n7672), .A3(n6686), .ZN(n7565) );
  AND2_X1 U7445 ( .A1(n7458), .A2(n9084), .ZN(n6836) );
  AND2_X1 U7446 ( .A1(n9118), .A2(n9119), .ZN(n7159) );
  AND4_X1 U7447 ( .A1(n8290), .A2(n8289), .A3(n8317), .A4(n7141), .ZN(n8291)
         );
  NAND2_X1 U7448 ( .A1(n7646), .A2(n7559), .ZN(n7648) );
  AND4_X1 U7449 ( .A1(n8282), .A2(n8281), .A3(n8280), .A4(n8476), .ZN(n8284)
         );
  INV_X1 U7450 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n15324) );
  INV_X1 U7451 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14487) );
  INV_X1 U7452 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13252) );
  INV_X1 U7453 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9084) );
  INV_X1 U7454 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9118) );
  INV_X1 U7455 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9160) );
  INV_X4 U7456 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7457 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9238) );
  INV_X1 U7458 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8561) );
  NOR2_X1 U7459 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8280) );
  NOR2_X1 U7460 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8281) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8282) );
  NOR2_X1 U7462 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7564) );
  NOR2_X1 U7463 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7563) );
  NOR2_X1 U7464 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7562) );
  INV_X1 U7465 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7598) );
  NOR2_X1 U7466 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7574) );
  INV_X1 U7467 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8123) );
  INV_X1 U7468 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7577) );
  INV_X1 U7469 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7578) );
  INV_X1 U7470 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8476) );
  INV_X2 U7471 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7472 ( .A1(n6974), .A2(n12553), .ZN(n12578) );
  NAND2_X1 U7473 ( .A1(n12799), .A2(n12804), .ZN(n12798) );
  AND2_X1 U7474 ( .A1(n11715), .A2(n6411), .ZN(n6422) );
  AND2_X1 U7475 ( .A1(n11715), .A2(n6411), .ZN(n11660) );
  NAND2_X1 U7476 ( .A1(n6702), .A2(n12345), .ZN(n7255) );
  XNOR2_X1 U7478 ( .A(n9231), .B(n9270), .ZN(n14317) );
  AND2_X2 U7479 ( .A1(n8326), .A2(n8283), .ZN(n8417) );
  AND2_X2 U7480 ( .A1(n6660), .A2(n6659), .ZN(n8326) );
  OR2_X1 U7481 ( .A1(n9895), .A2(n9896), .ZN(n7193) );
  AND2_X1 U7482 ( .A1(n9277), .A2(n9279), .ZN(n6791) );
  OR2_X2 U7483 ( .A1(n14203), .A2(n14609), .ZN(n6963) );
  NAND2_X1 U7484 ( .A1(n8299), .A2(n13676), .ZN(n8361) );
  NOR2_X1 U7485 ( .A1(n10893), .A2(n10894), .ZN(n11305) );
  NAND2_X2 U7486 ( .A1(n6407), .A2(n7606), .ZN(n8400) );
  NOR2_X2 U7487 ( .A1(n14631), .A2(n14632), .ZN(n14630) );
  XNOR2_X2 U7488 ( .A(n14335), .B(n7026), .ZN(n14375) );
  OAI21_X1 U7489 ( .B1(n9090), .B2(n6659), .A(n8352), .ZN(n13530) );
  OAI21_X2 U7490 ( .B1(n11381), .B2(n11380), .A(n11382), .ZN(n11383) );
  NOR2_X2 U7491 ( .A1(n13485), .A2(n13618), .ZN(n6771) );
  NOR2_X2 U7492 ( .A1(n14462), .A2(n14408), .ZN(n14466) );
  XNOR2_X2 U7493 ( .A(n8311), .B(n8310), .ZN(n8951) );
  OAI21_X2 U7494 ( .B1(n10535), .B2(n6462), .A(n7044), .ZN(n10444) );
  NOR2_X1 U7495 ( .A1(n15363), .A2(n15364), .ZN(n15362) );
  NAND2_X1 U7496 ( .A1(n8303), .A2(n8348), .ZN(n8389) );
  XNOR2_X2 U7497 ( .A(n8336), .B(n8343), .ZN(n8299) );
  NAND2_X2 U7498 ( .A1(n13670), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U7499 ( .A1(n7337), .A2(n7336), .ZN(n7335) );
  AND2_X1 U7500 ( .A1(n7847), .A2(n7576), .ZN(n7336) );
  NAND2_X1 U7501 ( .A1(n8866), .A2(n8865), .ZN(n8869) );
  XNOR2_X1 U7502 ( .A(n12904), .B(n12152), .ZN(n12465) );
  NAND2_X1 U7503 ( .A1(n6879), .A2(n13284), .ZN(n7221) );
  NAND2_X1 U7504 ( .A1(n13279), .A2(n7204), .ZN(n7202) );
  AND2_X1 U7505 ( .A1(n8307), .A2(n7141), .ZN(n7140) );
  INV_X1 U7506 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U7507 ( .A1(n8935), .A2(n8934), .ZN(n8976) );
  NAND2_X1 U7508 ( .A1(n7391), .A2(n7389), .ZN(n8935) );
  NOR2_X1 U7509 ( .A1(n7390), .A2(n8933), .ZN(n7389) );
  AND2_X1 U7510 ( .A1(n7379), .A2(n8602), .ZN(n7378) );
  NAND2_X1 U7511 ( .A1(n12262), .A2(n7934), .ZN(n12157) );
  NAND2_X1 U7512 ( .A1(n6916), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7185) );
  INV_X1 U7513 ( .A(n10343), .ZN(n6916) );
  NAND2_X1 U7514 ( .A1(n6685), .A2(n6807), .ZN(n12710) );
  NAND2_X1 U7515 ( .A1(n8238), .A2(n12736), .ZN(n6807) );
  NAND2_X1 U7516 ( .A1(n13558), .A2(n13124), .ZN(n13324) );
  NAND2_X1 U7517 ( .A1(n7061), .A2(n7063), .ZN(n13378) );
  AOI21_X1 U7518 ( .B1(n7064), .B2(n7066), .A(n13285), .ZN(n7063) );
  NAND2_X1 U7519 ( .A1(n13409), .A2(n7064), .ZN(n7061) );
  INV_X1 U7520 ( .A(n11660), .ZN(n11857) );
  AOI21_X1 U7521 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14357), .A(n14356), .ZN(
        n14415) );
  NOR2_X1 U7522 ( .A1(n14369), .A2(n14370), .ZN(n14356) );
  NAND2_X1 U7523 ( .A1(n11844), .A2(n13743), .ZN(n6844) );
  NAND2_X1 U7524 ( .A1(n8334), .A2(n8335), .ZN(n6649) );
  INV_X1 U7525 ( .A(n11623), .ZN(n6846) );
  NOR2_X1 U7526 ( .A1(n11630), .A2(n11648), .ZN(n7486) );
  NAND2_X1 U7527 ( .A1(n6633), .A2(n8575), .ZN(n6632) );
  MUX2_X1 U7528 ( .A(n13988), .B(n14073), .S(n11867), .Z(n11744) );
  AND2_X1 U7529 ( .A1(n7590), .A2(n7589), .ZN(n7811) );
  NAND2_X1 U7530 ( .A1(n7303), .A2(n7302), .ZN(n11067) );
  INV_X1 U7531 ( .A(n11888), .ZN(n7302) );
  INV_X1 U7532 ( .A(n11065), .ZN(n7303) );
  INV_X1 U7533 ( .A(n8653), .ZN(n7365) );
  NAND2_X1 U7534 ( .A1(n12251), .A2(n8008), .ZN(n8017) );
  INV_X1 U7535 ( .A(n7811), .ZN(n12006) );
  AND2_X1 U7536 ( .A1(n11465), .A2(n6891), .ZN(n6890) );
  NAND2_X1 U7537 ( .A1(n12240), .A2(n6892), .ZN(n6891) );
  OR2_X1 U7538 ( .A1(n10005), .A2(n10267), .ZN(n6926) );
  NAND2_X1 U7539 ( .A1(n6925), .A2(n9826), .ZN(n6924) );
  NAND2_X1 U7540 ( .A1(n12900), .A2(n12749), .ZN(n12470) );
  OR2_X1 U7541 ( .A1(n12900), .A2(n12749), .ZN(n12474) );
  AND2_X1 U7542 ( .A1(n12453), .A2(n12801), .ZN(n12454) );
  OR2_X1 U7543 ( .A1(n12453), .A2(n12801), .ZN(n12317) );
  OAI21_X1 U7544 ( .B1(n7436), .B2(n7434), .A(n8192), .ZN(n7433) );
  OR2_X1 U7545 ( .A1(n12977), .A2(n12828), .ZN(n8192) );
  OR2_X1 U7546 ( .A1(n8190), .A2(n8191), .ZN(n12437) );
  OR2_X1 U7547 ( .A1(n14499), .A2(n12511), .ZN(n12418) );
  INV_X1 U7548 ( .A(n7429), .ZN(n6681) );
  AOI21_X1 U7549 ( .B1(n7431), .B2(n12378), .A(n6520), .ZN(n7429) );
  INV_X1 U7550 ( .A(n8158), .ZN(n6852) );
  INV_X1 U7551 ( .A(n7783), .ZN(n7089) );
  OAI21_X1 U7552 ( .B1(n7073), .B2(n7077), .A(n6511), .ZN(n7072) );
  INV_X1 U7553 ( .A(n7074), .ZN(n7073) );
  NOR2_X1 U7554 ( .A1(n11243), .A2(n15054), .ZN(n7036) );
  NAND2_X1 U7555 ( .A1(n11863), .A2(n9282), .ZN(n9724) );
  INV_X1 U7556 ( .A(n13836), .ZN(n11556) );
  XNOR2_X1 U7557 ( .A(n14026), .B(n11873), .ZN(n14018) );
  AND2_X1 U7558 ( .A1(n9281), .A2(n11860), .ZN(n11541) );
  NAND2_X1 U7559 ( .A1(n10279), .A2(n11883), .ZN(n7172) );
  NAND2_X1 U7560 ( .A1(n7172), .A2(n7171), .ZN(n10554) );
  AND2_X1 U7561 ( .A1(n11884), .A2(n10280), .ZN(n7171) );
  NAND2_X1 U7562 ( .A1(n8890), .A2(n8889), .ZN(n8908) );
  NAND2_X1 U7563 ( .A1(n8869), .A2(n8868), .ZN(n8888) );
  NAND2_X1 U7564 ( .A1(n9126), .A2(n7532), .ZN(n7531) );
  OR2_X1 U7565 ( .A1(n8828), .A2(n7371), .ZN(n7369) );
  NAND2_X1 U7566 ( .A1(n8766), .A2(SI_18_), .ZN(n7387) );
  INV_X1 U7567 ( .A(n8532), .ZN(n8533) );
  XNOR2_X1 U7568 ( .A(n8510), .B(SI_7_), .ZN(n8508) );
  NAND2_X1 U7569 ( .A1(n7159), .A2(n9130), .ZN(n9224) );
  NAND2_X1 U7570 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7012), .ZN(n7011) );
  INV_X1 U7571 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7012) );
  NAND2_X1 U7572 ( .A1(n14375), .A2(n14336), .ZN(n7025) );
  NAND2_X1 U7573 ( .A1(n7836), .A2(n12512), .ZN(n6892) );
  INV_X1 U7574 ( .A(n12220), .ZN(n6898) );
  AND2_X1 U7575 ( .A1(n7321), .A2(n6884), .ZN(n6883) );
  NAND2_X1 U7576 ( .A1(n6886), .A2(n6888), .ZN(n6884) );
  NOR2_X1 U7577 ( .A1(n12233), .A2(n7329), .ZN(n7328) );
  INV_X1 U7578 ( .A(n7952), .ZN(n7329) );
  NOR2_X1 U7579 ( .A1(n6539), .A2(n6786), .ZN(n6785) );
  INV_X1 U7580 ( .A(n12326), .ZN(n6788) );
  XNOR2_X1 U7581 ( .A(n6697), .B(n12687), .ZN(n6696) );
  NAND2_X1 U7582 ( .A1(n6695), .A2(n6694), .ZN(n6697) );
  AOI21_X1 U7583 ( .B1(n6459), .B2(n12495), .A(n6445), .ZN(n6694) );
  NAND2_X1 U7584 ( .A1(n12496), .A2(n6459), .ZN(n6695) );
  NAND2_X1 U7585 ( .A1(n7084), .A2(n6737), .ZN(n12489) );
  AND2_X1 U7586 ( .A1(n6738), .A2(n12295), .ZN(n6737) );
  INV_X1 U7587 ( .A(n6929), .ZN(n9893) );
  NAND2_X1 U7588 ( .A1(n6986), .A2(n6985), .ZN(n10328) );
  INV_X1 U7589 ( .A(n9879), .ZN(n6985) );
  INV_X1 U7590 ( .A(n10886), .ZN(n10887) );
  OR2_X1 U7591 ( .A1(n8197), .A2(n12749), .ZN(n7556) );
  OAI21_X1 U7592 ( .B1(n8234), .B2(n7284), .A(n7282), .ZN(n8237) );
  INV_X1 U7593 ( .A(n7283), .ZN(n7282) );
  NAND2_X1 U7594 ( .A1(n12798), .A2(n7538), .ZN(n12789) );
  OR2_X1 U7595 ( .A1(n12973), .A2(n12816), .ZN(n7538) );
  OR2_X1 U7596 ( .A1(n12237), .A2(n12816), .ZN(n12450) );
  NAND2_X1 U7597 ( .A1(n11279), .A2(n12406), .ZN(n8183) );
  NAND2_X1 U7598 ( .A1(n10759), .A2(n8226), .ZN(n10840) );
  NAND2_X1 U7599 ( .A1(n10315), .A2(n12377), .ZN(n10760) );
  NAND2_X1 U7600 ( .A1(n10760), .A2(n12378), .ZN(n10759) );
  NAND2_X1 U7601 ( .A1(n8203), .A2(n8202), .ZN(n8255) );
  INV_X1 U7602 ( .A(n12299), .ZN(n7948) );
  INV_X1 U7603 ( .A(n8068), .ZN(n12296) );
  AND2_X1 U7604 ( .A1(n6519), .A2(n6684), .ZN(n6683) );
  INV_X1 U7605 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U7606 ( .A1(n8160), .A2(n8159), .ZN(n8201) );
  AND2_X1 U7607 ( .A1(n7351), .A2(n7578), .ZN(n7350) );
  AND2_X1 U7608 ( .A1(n7972), .A2(n11681), .ZN(n7091) );
  NAND2_X1 U7609 ( .A1(n7876), .A2(n7875), .ZN(n7879) );
  NAND2_X1 U7610 ( .A1(n7879), .A2(n7878), .ZN(n7904) );
  OR2_X1 U7611 ( .A1(n7781), .A2(n6718), .ZN(n7085) );
  INV_X1 U7612 ( .A(n7088), .ZN(n6718) );
  OAI21_X1 U7613 ( .B1(n7700), .B2(n6723), .A(n6721), .ZN(n7731) );
  INV_X1 U7614 ( .A(n6724), .ZN(n6723) );
  AOI21_X1 U7615 ( .B1(n6724), .B2(n6722), .A(n6534), .ZN(n6721) );
  NOR2_X1 U7616 ( .A1(n7716), .A2(n6725), .ZN(n6724) );
  AND2_X1 U7617 ( .A1(n7113), .A2(n6521), .ZN(n6440) );
  AND2_X1 U7618 ( .A1(n6440), .A2(n13020), .ZN(n7111) );
  NAND2_X1 U7619 ( .A1(n8963), .A2(n8962), .ZN(n13555) );
  AOI21_X1 U7620 ( .B1(n7056), .B2(n7059), .A(n13323), .ZN(n7054) );
  AOI21_X1 U7621 ( .B1(n7215), .B2(n7213), .A(n6536), .ZN(n7212) );
  INV_X1 U7622 ( .A(n6464), .ZN(n7213) );
  AOI21_X1 U7623 ( .B1(n7200), .B2(n7198), .A(n6516), .ZN(n7197) );
  INV_X1 U7624 ( .A(n7204), .ZN(n7198) );
  NAND2_X1 U7625 ( .A1(n13424), .A2(n6488), .ZN(n13409) );
  AOI22_X1 U7626 ( .A1(n13438), .A2(n13437), .B1(n13604), .B2(n13310), .ZN(
        n13426) );
  OR2_X1 U7627 ( .A1(n13439), .A2(n13310), .ZN(n7204) );
  NOR2_X1 U7628 ( .A1(n11040), .A2(n7228), .ZN(n7227) );
  INV_X1 U7629 ( .A(n8291), .ZN(n7456) );
  NAND2_X1 U7630 ( .A1(n8309), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U7631 ( .A1(n11856), .A2(n11855), .ZN(n11871) );
  MUX2_X1 U7632 ( .A(n11910), .B(n11909), .S(n11908), .Z(n11911) );
  NAND2_X1 U7633 ( .A1(n11826), .A2(n11825), .ZN(n14202) );
  INV_X1 U7634 ( .A(n6953), .ZN(n6952) );
  NAND2_X1 U7635 ( .A1(n6623), .A2(n7158), .ZN(n6622) );
  INV_X1 U7636 ( .A(n7307), .ZN(n7306) );
  OAI21_X1 U7637 ( .B1(n7309), .B2(n7310), .A(n13989), .ZN(n7307) );
  NAND2_X1 U7638 ( .A1(n14064), .A2(n13954), .ZN(n14050) );
  NOR2_X1 U7639 ( .A1(n11884), .A2(n11883), .ZN(n7287) );
  XNOR2_X1 U7640 ( .A(n14202), .B(n13998), .ZN(n13992) );
  NOR2_X1 U7641 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6709) );
  NAND2_X1 U7642 ( .A1(n6833), .A2(n6834), .ZN(n14419) );
  OAI21_X1 U7643 ( .B1(n14650), .B2(n14649), .A(n7018), .ZN(n7017) );
  INV_X1 U7644 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7018) );
  INV_X1 U7645 ( .A(n7347), .ZN(n7346) );
  OAI21_X1 U7646 ( .B1(n7348), .B2(n10676), .A(n7762), .ZN(n7347) );
  INV_X1 U7647 ( .A(n12697), .ZN(n12726) );
  NAND2_X1 U7648 ( .A1(n13678), .A2(n11791), .ZN(n11808) );
  NAND2_X1 U7649 ( .A1(n14650), .A2(n14649), .ZN(n14648) );
  NAND2_X1 U7650 ( .A1(n6841), .A2(n7498), .ZN(n11581) );
  NAND2_X1 U7651 ( .A1(n11575), .A2(n11577), .ZN(n7498) );
  OR2_X1 U7652 ( .A1(n11575), .A2(n11577), .ZN(n7497) );
  NAND2_X1 U7653 ( .A1(n8359), .A2(n6643), .ZN(n6642) );
  NOR2_X1 U7654 ( .A1(n6855), .A2(n6637), .ZN(n6636) );
  INV_X1 U7655 ( .A(n8489), .ZN(n6631) );
  NAND2_X1 U7656 ( .A1(n6667), .A2(n7453), .ZN(n6666) );
  NAND2_X1 U7657 ( .A1(n8461), .A2(n6447), .ZN(n7453) );
  NOR2_X1 U7658 ( .A1(n6486), .A2(n6631), .ZN(n6629) );
  NAND2_X1 U7659 ( .A1(n11620), .A2(n11621), .ZN(n7471) );
  NAND2_X1 U7660 ( .A1(n8526), .A2(n8527), .ZN(n8525) );
  INV_X1 U7661 ( .A(n7486), .ZN(n7482) );
  MUX2_X1 U7662 ( .A(n13985), .B(n13986), .S(n11867), .Z(n11716) );
  AND2_X1 U7663 ( .A1(n7478), .A2(n11702), .ZN(n7477) );
  OR2_X1 U7664 ( .A1(n8669), .A2(n8668), .ZN(n6658) );
  NAND2_X1 U7665 ( .A1(n11744), .A2(n7491), .ZN(n7490) );
  INV_X1 U7666 ( .A(n11745), .ZN(n7491) );
  INV_X1 U7667 ( .A(n8763), .ZN(n6639) );
  NAND2_X1 U7668 ( .A1(n6451), .A2(n6570), .ZN(n7461) );
  INV_X1 U7669 ( .A(n8762), .ZN(n6850) );
  OAI21_X1 U7670 ( .B1(n8723), .B2(n8722), .A(n6453), .ZN(n7460) );
  INV_X1 U7671 ( .A(n11777), .ZN(n6813) );
  INV_X1 U7672 ( .A(n12468), .ZN(n6795) );
  XNOR2_X1 U7673 ( .A(n14326), .B(n14471), .ZN(n11537) );
  INV_X1 U7674 ( .A(n8804), .ZN(n6652) );
  NAND2_X1 U7675 ( .A1(n6743), .A2(n12483), .ZN(n6742) );
  NAND2_X1 U7676 ( .A1(n12472), .A2(n12471), .ZN(n6743) );
  NAND2_X1 U7677 ( .A1(n12476), .A2(n12487), .ZN(n6741) );
  OAI21_X1 U7678 ( .B1(n10050), .B2(n9827), .A(n6435), .ZN(n6925) );
  INV_X1 U7679 ( .A(n11034), .ZN(n7229) );
  NAND2_X1 U7680 ( .A1(n11839), .A2(n11536), .ZN(n11827) );
  INV_X1 U7681 ( .A(n8960), .ZN(n7410) );
  AOI21_X1 U7682 ( .B1(n8907), .B2(n7401), .A(n7400), .ZN(n7399) );
  INV_X1 U7683 ( .A(n8931), .ZN(n7400) );
  AOI21_X1 U7684 ( .B1(n8907), .B2(n8894), .A(SI_26_), .ZN(n7402) );
  NAND2_X1 U7685 ( .A1(n8583), .A2(n8582), .ZN(n8602) );
  INV_X1 U7686 ( .A(n8553), .ZN(n8554) );
  AOI21_X1 U7687 ( .B1(n8490), .B2(n8493), .A(n8508), .ZN(n7357) );
  OAI21_X1 U7688 ( .B1(n6411), .B2(n9176), .A(n6871), .ZN(n8492) );
  NAND2_X1 U7689 ( .A1(n6412), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6871) );
  NOR2_X1 U7690 ( .A1(n7935), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7963) );
  AND2_X1 U7691 ( .A1(n7736), .A2(n9889), .ZN(n7746) );
  NOR2_X1 U7692 ( .A1(n11206), .A2(n7779), .ZN(n7797) );
  NAND2_X1 U7693 ( .A1(n12302), .A2(n12690), .ZN(n6746) );
  INV_X1 U7694 ( .A(n15120), .ZN(n6987) );
  OR2_X1 U7695 ( .A1(n12330), .A2(n8026), .ZN(n12329) );
  NAND2_X1 U7696 ( .A1(n12783), .A2(n12461), .ZN(n7261) );
  OAI21_X1 U7697 ( .B1(n7285), .B2(n7284), .A(n8235), .ZN(n7283) );
  INV_X1 U7698 ( .A(n8189), .ZN(n6679) );
  INV_X1 U7699 ( .A(n7438), .ZN(n7437) );
  AOI21_X1 U7700 ( .B1(n7421), .B2(n7423), .A(n7420), .ZN(n7419) );
  OR2_X1 U7701 ( .A1(n14504), .A2(n12512), .ZN(n12414) );
  INV_X1 U7702 ( .A(n8227), .ZN(n7273) );
  OR2_X1 U7703 ( .A1(n7771), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U7704 ( .A1(n10807), .A2(n10650), .ZN(n12344) );
  NOR2_X1 U7705 ( .A1(n12804), .A2(n7286), .ZN(n7285) );
  INV_X1 U7706 ( .A(n12445), .ZN(n7286) );
  NAND2_X1 U7707 ( .A1(n10840), .A2(n8227), .ZN(n7277) );
  AND2_X1 U7708 ( .A1(n6456), .A2(n8065), .ZN(n6720) );
  AND2_X1 U7709 ( .A1(n7566), .A2(n7577), .ZN(n7351) );
  AND2_X1 U7710 ( .A1(n7095), .A2(n6734), .ZN(n6733) );
  NAND2_X1 U7711 ( .A1(n7859), .A2(n7875), .ZN(n6734) );
  INV_X1 U7712 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n6687) );
  INV_X1 U7713 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U7714 ( .A1(n6716), .A2(n7663), .ZN(n6715) );
  INV_X1 U7715 ( .A(n7610), .ZN(n6716) );
  AND2_X1 U7716 ( .A1(n9028), .A2(n7441), .ZN(n7440) );
  NAND2_X1 U7717 ( .A1(n8927), .A2(n7442), .ZN(n7441) );
  OAI21_X1 U7718 ( .B1(n8922), .B2(n8923), .A(n7443), .ZN(n7442) );
  NAND2_X1 U7719 ( .A1(n8884), .A2(n8885), .ZN(n7446) );
  INV_X1 U7720 ( .A(n8299), .ZN(n8303) );
  NAND2_X1 U7721 ( .A1(n8910), .A2(n8909), .ZN(n13582) );
  NAND2_X1 U7722 ( .A1(n11043), .A2(n15047), .ZN(n11192) );
  NOR2_X1 U7723 ( .A1(n10935), .A2(n15038), .ZN(n11043) );
  XNOR2_X1 U7724 ( .A(n13143), .B(n14783), .ZN(n10152) );
  AND2_X1 U7725 ( .A1(n8293), .A2(n8294), .ZN(n6837) );
  INV_X1 U7726 ( .A(n14065), .ZN(n7310) );
  NAND2_X1 U7727 ( .A1(n13984), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U7728 ( .A1(n11380), .A2(n11624), .ZN(n7176) );
  OR2_X1 U7729 ( .A1(n12036), .A2(n14553), .ZN(n11629) );
  NOR2_X1 U7730 ( .A1(n11352), .A2(n12036), .ZN(n7003) );
  INV_X1 U7731 ( .A(n13957), .ZN(n7152) );
  AND2_X1 U7732 ( .A1(n7155), .A2(n13959), .ZN(n7154) );
  AOI21_X1 U7733 ( .B1(n11069), .B2(n6971), .A(n6515), .ZN(n6970) );
  INV_X1 U7734 ( .A(n11066), .ZN(n6971) );
  OR2_X1 U7735 ( .A1(n11067), .A2(n11889), .ZN(n6969) );
  AOI21_X1 U7736 ( .B1(n7363), .B2(n7365), .A(n7361), .ZN(n7360) );
  INV_X1 U7737 ( .A(n8703), .ZN(n7361) );
  AOI21_X1 U7738 ( .B1(n8579), .B2(n7382), .A(n6524), .ZN(n7381) );
  INV_X1 U7739 ( .A(n8557), .ZN(n7382) );
  XNOR2_X1 U7740 ( .A(n8492), .B(SI_6_), .ZN(n8490) );
  NAND2_X1 U7741 ( .A1(n6945), .A2(n8475), .ZN(n6878) );
  INV_X1 U7742 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7026) );
  INV_X1 U7743 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7024) );
  OAI21_X1 U7744 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14348), .A(n14347), .ZN(
        n14373) );
  NAND2_X1 U7745 ( .A1(n8015), .A2(n8014), .ZN(n8018) );
  AND2_X1 U7746 ( .A1(n12219), .A2(n12195), .ZN(n6896) );
  AND2_X1 U7747 ( .A1(n8064), .A2(n8063), .ZN(n12193) );
  AND2_X1 U7748 ( .A1(n12202), .A2(n7322), .ZN(n7321) );
  OR2_X1 U7749 ( .A1(n12280), .A2(n7323), .ZN(n7322) );
  INV_X1 U7750 ( .A(n7874), .ZN(n7323) );
  AND2_X1 U7751 ( .A1(n12195), .A2(n8045), .ZN(n12220) );
  NAND2_X1 U7752 ( .A1(n8017), .A2(n8016), .ZN(n12219) );
  NOR2_X1 U7753 ( .A1(n10627), .A2(n7342), .ZN(n7341) );
  INV_X1 U7754 ( .A(n7668), .ZN(n7342) );
  NAND2_X1 U7755 ( .A1(n12157), .A2(n12158), .ZN(n7953) );
  NAND2_X1 U7756 ( .A1(n7797), .A2(n7796), .ZN(n11457) );
  NAND2_X1 U7757 ( .A1(n7317), .A2(n10650), .ZN(n10810) );
  XNOR2_X1 U7758 ( .A(n7654), .B(n12349), .ZN(n7655) );
  INV_X1 U7759 ( .A(n12213), .ZN(n6907) );
  INV_X1 U7760 ( .A(n6890), .ZN(n6888) );
  AOI21_X1 U7761 ( .B1(n6890), .B2(n6887), .A(n6441), .ZN(n6886) );
  INV_X1 U7762 ( .A(n6892), .ZN(n6887) );
  NOR2_X1 U7763 ( .A1(n9875), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9776) );
  OR2_X1 U7764 ( .A1(n7561), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7182) );
  OAI21_X1 U7765 ( .B1(n7649), .B2(n7561), .A(P3_REG2_REG_2__SCAN_IN), .ZN(
        n7181) );
  INV_X1 U7766 ( .A(n9990), .ZN(n7186) );
  INV_X1 U7767 ( .A(n9897), .ZN(n7192) );
  NAND2_X1 U7768 ( .A1(n10328), .A2(n10327), .ZN(n6984) );
  NOR2_X1 U7769 ( .A1(n10915), .A2(n15343), .ZN(n11325) );
  XNOR2_X1 U7770 ( .A(n6760), .B(n14455), .ZN(n11329) );
  NAND2_X1 U7771 ( .A1(n7267), .A2(n12754), .ZN(n7264) );
  AND2_X1 U7772 ( .A1(n7269), .A2(n6473), .ZN(n7267) );
  INV_X1 U7773 ( .A(n7270), .ZN(n7269) );
  OAI21_X1 U7774 ( .B1(n12739), .B2(n12327), .A(n12470), .ZN(n7270) );
  AND2_X1 U7775 ( .A1(n6473), .A2(n12471), .ZN(n12727) );
  NAND2_X1 U7776 ( .A1(n6701), .A2(n7258), .ZN(n12753) );
  AOI21_X1 U7777 ( .B1(n12762), .B2(n7260), .A(n7259), .ZN(n7258) );
  NAND2_X1 U7778 ( .A1(n12783), .A2(n7256), .ZN(n6701) );
  INV_X1 U7779 ( .A(n12460), .ZN(n7260) );
  OR2_X1 U7780 ( .A1(n12961), .A2(n8026), .ZN(n7544) );
  NAND2_X1 U7781 ( .A1(n12779), .A2(n8193), .ZN(n6677) );
  OR2_X1 U7782 ( .A1(n12977), .A2(n12800), .ZN(n12445) );
  NAND2_X1 U7783 ( .A1(n12450), .A2(n12449), .ZN(n12804) );
  AOI21_X1 U7784 ( .B1(n7280), .B2(n12837), .A(n7279), .ZN(n7278) );
  INV_X1 U7785 ( .A(n12437), .ZN(n7279) );
  NAND2_X1 U7786 ( .A1(n12845), .A2(n12844), .ZN(n12843) );
  NAND2_X1 U7787 ( .A1(n11229), .A2(n8230), .ZN(n6703) );
  NAND2_X1 U7788 ( .A1(n8181), .A2(n8180), .ZN(n11279) );
  AND2_X1 U7789 ( .A1(n12314), .A2(n6479), .ZN(n7425) );
  NAND2_X1 U7790 ( .A1(n10949), .A2(n7427), .ZN(n7426) );
  AOI21_X1 U7791 ( .B1(n11462), .B2(n11202), .A(n7428), .ZN(n7427) );
  INV_X1 U7792 ( .A(n8179), .ZN(n7428) );
  OAI21_X1 U7793 ( .B1(n10317), .B2(n7430), .A(n6680), .ZN(n10950) );
  AOI21_X1 U7794 ( .B1(n7431), .B2(n6682), .A(n6681), .ZN(n6680) );
  INV_X1 U7795 ( .A(n8174), .ZN(n6682) );
  NAND2_X1 U7796 ( .A1(n10950), .A2(n12310), .ZN(n10949) );
  AND2_X1 U7797 ( .A1(n10754), .A2(n8177), .ZN(n10843) );
  NAND2_X1 U7798 ( .A1(n8176), .A2(n8175), .ZN(n10754) );
  INV_X1 U7799 ( .A(n10756), .ZN(n8176) );
  AND2_X1 U7800 ( .A1(n12377), .A2(n12376), .ZN(n12373) );
  NAND2_X1 U7801 ( .A1(n10214), .A2(n6496), .ZN(n10422) );
  NAND2_X1 U7802 ( .A1(n12487), .A2(n8142), .ZN(n12873) );
  NAND2_X1 U7803 ( .A1(n10854), .A2(n7424), .ZN(n10214) );
  NOR2_X1 U7804 ( .A1(n12366), .A2(n6840), .ZN(n7424) );
  INV_X1 U7805 ( .A(n8171), .ZN(n6840) );
  NAND2_X1 U7806 ( .A1(n12360), .A2(n12365), .ZN(n12356) );
  NAND2_X1 U7807 ( .A1(n8224), .A2(n12344), .ZN(n10804) );
  NAND2_X1 U7808 ( .A1(n8034), .A2(n8033), .ZN(n12904) );
  NAND2_X1 U7809 ( .A1(n8234), .A2(n7285), .ZN(n12922) );
  NAND2_X1 U7810 ( .A1(n8160), .A2(n6731), .ZN(n6730) );
  NOR2_X1 U7811 ( .A1(n7099), .A2(n6732), .ZN(n6731) );
  INV_X1 U7812 ( .A(n8159), .ZN(n6732) );
  NAND2_X1 U7813 ( .A1(n6600), .A2(n11522), .ZN(n7099) );
  NAND2_X1 U7814 ( .A1(n6730), .A2(n7098), .ZN(n11524) );
  NAND2_X1 U7815 ( .A1(n7617), .A2(n12989), .ZN(n6698) );
  MUX2_X1 U7816 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7616), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7617) );
  OAI21_X1 U7817 ( .B1(n8082), .B2(n8081), .A(n8083), .ZN(n8158) );
  NAND2_X1 U7818 ( .A1(n8047), .A2(n8032), .ZN(n8046) );
  OAI21_X1 U7819 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8028) );
  NAND2_X1 U7820 ( .A1(n7993), .A2(n7992), .ZN(n8011) );
  OR2_X1 U7821 ( .A1(n7956), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U7822 ( .A1(n7956), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U7823 ( .A1(n6736), .A2(n7860), .ZN(n7876) );
  NAND2_X1 U7824 ( .A1(n7844), .A2(n6739), .ZN(n7843) );
  OR2_X1 U7825 ( .A1(n7823), .A2(n11059), .ZN(n6739) );
  AOI21_X1 U7826 ( .B1(n7088), .B2(n7087), .A(n6581), .ZN(n7086) );
  INV_X1 U7827 ( .A(n7780), .ZN(n7087) );
  NAND2_X1 U7828 ( .A1(n7764), .A2(n7763), .ZN(n6719) );
  XNOR2_X1 U7829 ( .A(n9183), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U7830 ( .A1(n7677), .A2(n7676), .ZN(n7679) );
  XNOR2_X1 U7831 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7699) );
  NAND2_X1 U7832 ( .A1(n9138), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U7833 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7663) );
  NAND2_X1 U7834 ( .A1(n7609), .A2(n7608), .ZN(n7651) );
  NAND2_X1 U7835 ( .A1(n9152), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7608) );
  XNOR2_X1 U7836 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7650) );
  BUF_X1 U7837 ( .A(n7646), .Z(n9828) );
  OR2_X1 U7838 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  AND2_X1 U7839 ( .A1(n10875), .A2(n10817), .ZN(n7117) );
  NAND2_X1 U7840 ( .A1(n13030), .A2(n11935), .ZN(n13086) );
  NOR2_X1 U7841 ( .A1(n13343), .A2(n13555), .ZN(n13328) );
  NAND2_X1 U7842 ( .A1(n13328), .A2(n13552), .ZN(n13260) );
  XNOR2_X1 U7843 ( .A(n13555), .B(n9050), .ZN(n13325) );
  INV_X1 U7844 ( .A(n7029), .ZN(n13355) );
  NAND2_X1 U7845 ( .A1(n7219), .A2(n7221), .ZN(n7218) );
  NAND2_X1 U7846 ( .A1(n13395), .A2(n7222), .ZN(n7220) );
  AND2_X1 U7847 ( .A1(n13395), .A2(n13313), .ZN(n7067) );
  NAND2_X1 U7848 ( .A1(n13587), .A2(n13056), .ZN(n7222) );
  AND2_X1 U7849 ( .A1(n7196), .A2(n6549), .ZN(n13282) );
  OR2_X1 U7850 ( .A1(n13436), .A2(n7201), .ZN(n7196) );
  INV_X1 U7851 ( .A(n7079), .ZN(n7078) );
  AOI21_X1 U7852 ( .B1(n7077), .B2(n7079), .A(n7075), .ZN(n7074) );
  INV_X1 U7853 ( .A(n13305), .ZN(n7075) );
  NOR2_X1 U7854 ( .A1(n13623), .A2(n13128), .ZN(n7079) );
  NOR2_X1 U7855 ( .A1(n13272), .A2(n7254), .ZN(n7253) );
  INV_X1 U7856 ( .A(n13270), .ZN(n7254) );
  NAND2_X1 U7857 ( .A1(n7251), .A2(n13273), .ZN(n7250) );
  OR2_X1 U7858 ( .A1(n13272), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U7859 ( .A1(n13271), .A2(n13270), .ZN(n7252) );
  OR2_X1 U7860 ( .A1(n13301), .A2(n13511), .ZN(n7547) );
  NOR2_X1 U7861 ( .A1(n13478), .A2(n13479), .ZN(n13477) );
  INV_X1 U7862 ( .A(n13302), .ZN(n13479) );
  NOR2_X1 U7863 ( .A1(n6568), .A2(n7206), .ZN(n7205) );
  OR2_X1 U7864 ( .A1(n11512), .A2(n13132), .ZN(n7051) );
  NAND2_X1 U7865 ( .A1(n11185), .A2(n11175), .ZN(n7232) );
  OR2_X1 U7866 ( .A1(n10746), .A2(n15029), .ZN(n10935) );
  NAND2_X1 U7867 ( .A1(n10717), .A2(n7030), .ZN(n10746) );
  NOR2_X1 U7868 ( .A1(n15020), .A2(n10720), .ZN(n7030) );
  NAND2_X1 U7869 ( .A1(n10717), .A2(n15011), .ZN(n10716) );
  NAND2_X1 U7870 ( .A1(n7239), .A2(n10392), .ZN(n10725) );
  NAND2_X1 U7871 ( .A1(n10393), .A2(n10394), .ZN(n7239) );
  OAI211_X1 U7872 ( .C1(n10609), .C2(n7195), .A(n10152), .B(n7194), .ZN(n10545) );
  OR2_X1 U7873 ( .A1(n10610), .A2(n7195), .ZN(n7194) );
  INV_X1 U7874 ( .A(n10151), .ZN(n7195) );
  NAND2_X1 U7875 ( .A1(n10609), .A2(n10610), .ZN(n10608) );
  OR2_X1 U7876 ( .A1(n14978), .A2(n9752), .ZN(n10366) );
  NAND2_X1 U7877 ( .A1(n13681), .A2(n9005), .ZN(n9009) );
  INV_X1 U7878 ( .A(n13373), .ZN(n13574) );
  AND2_X1 U7879 ( .A1(n9769), .A2(n9760), .ZN(n15053) );
  INV_X1 U7880 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U7881 ( .A1(n8320), .A2(n8321), .ZN(n8296) );
  NAND2_X1 U7882 ( .A1(n9077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8324) );
  AND2_X1 U7883 ( .A1(n9075), .A2(n9088), .ZN(n9083) );
  INV_X1 U7884 ( .A(n7139), .ZN(n7137) );
  NOR2_X1 U7885 ( .A1(n8679), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8707) );
  INV_X1 U7886 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8283) );
  AND2_X1 U7887 ( .A1(n13802), .A2(n7506), .ZN(n7505) );
  OR2_X1 U7888 ( .A1(n13727), .A2(n7507), .ZN(n7506) );
  INV_X1 U7889 ( .A(n12115), .ZN(n7507) );
  NAND2_X1 U7890 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  INV_X1 U7891 ( .A(n10186), .ZN(n10189) );
  AOI21_X1 U7892 ( .B1(n7510), .B2(n7512), .A(n6509), .ZN(n7509) );
  INV_X1 U7893 ( .A(n10252), .ZN(n6708) );
  AOI21_X1 U7894 ( .B1(n13838), .B2(n9562), .A(n9561), .ZN(n9567) );
  OR2_X1 U7895 ( .A1(n9563), .A2(n9906), .ZN(n6778) );
  AOI22_X1 U7896 ( .A1(n7516), .A2(n10503), .B1(n10504), .B2(n10505), .ZN(
        n13738) );
  NAND2_X1 U7897 ( .A1(n14544), .A2(n12035), .ZN(n12046) );
  INV_X1 U7898 ( .A(n11818), .ZN(n11706) );
  OR2_X1 U7899 ( .A1(n11818), .A2(n10051), .ZN(n9602) );
  OR2_X1 U7900 ( .A1(n6802), .A2(n9599), .ZN(n9600) );
  NAND2_X1 U7901 ( .A1(n13962), .A2(n14272), .ZN(n13929) );
  AND2_X1 U7902 ( .A1(n14044), .A2(n6994), .ZN(n13962) );
  AND2_X1 U7903 ( .A1(n6995), .A2(n6419), .ZN(n6994) );
  NAND2_X1 U7904 ( .A1(n14044), .A2(n6995), .ZN(n14003) );
  NAND2_X1 U7905 ( .A1(n14048), .A2(n13957), .ZN(n14041) );
  NAND2_X1 U7906 ( .A1(n7311), .A2(n7310), .ZN(n7308) );
  INV_X1 U7907 ( .A(n14061), .ZN(n7311) );
  INV_X1 U7908 ( .A(n7308), .ZN(n14060) );
  AND2_X1 U7909 ( .A1(n14080), .A2(n13952), .ZN(n14066) );
  OAI21_X1 U7910 ( .B1(n14093), .B2(n14095), .A(n13950), .ZN(n14082) );
  NAND2_X1 U7911 ( .A1(n7294), .A2(n7292), .ZN(n14078) );
  NOR2_X1 U7912 ( .A1(n14081), .A2(n7293), .ZN(n7292) );
  INV_X1 U7913 ( .A(n7296), .ZN(n7293) );
  OR2_X1 U7914 ( .A1(n14292), .A2(n13983), .ZN(n7301) );
  NAND2_X1 U7915 ( .A1(n14122), .A2(n13945), .ZN(n14108) );
  OAI21_X1 U7916 ( .B1(n14156), .B2(n6615), .A(n6612), .ZN(n14122) );
  INV_X1 U7917 ( .A(n7162), .ZN(n6615) );
  AND2_X1 U7918 ( .A1(n7160), .A2(n6613), .ZN(n6612) );
  NAND2_X1 U7919 ( .A1(n7162), .A2(n6614), .ZN(n6613) );
  AND2_X1 U7920 ( .A1(n14146), .A2(n13941), .ZN(n7162) );
  NAND2_X1 U7921 ( .A1(n14156), .A2(n14160), .ZN(n13942) );
  NAND2_X1 U7922 ( .A1(n6611), .A2(n7173), .ZN(n11379) );
  NAND2_X1 U7923 ( .A1(n7176), .A2(n11629), .ZN(n7173) );
  NAND2_X1 U7924 ( .A1(n11160), .A2(n6609), .ZN(n6611) );
  NOR2_X1 U7925 ( .A1(n7174), .A2(n6610), .ZN(n6609) );
  INV_X1 U7926 ( .A(n7176), .ZN(n7175) );
  INV_X1 U7927 ( .A(n11893), .ZN(n11380) );
  NOR2_X1 U7928 ( .A1(n11150), .A2(n14469), .ZN(n7005) );
  NAND2_X1 U7929 ( .A1(n7005), .A2(n7004), .ZN(n11352) );
  INV_X1 U7930 ( .A(n14606), .ZN(n7004) );
  INV_X1 U7931 ( .A(n6616), .ZN(n10978) );
  OAI21_X1 U7932 ( .B1(n10976), .B2(n10975), .A(n6526), .ZN(n6616) );
  OAI21_X1 U7933 ( .B1(n10966), .B2(n10965), .A(n10967), .ZN(n11065) );
  XNOR2_X1 U7934 ( .A(n14756), .B(n11258), .ZN(n7146) );
  AND2_X1 U7935 ( .A1(n10554), .A2(n10553), .ZN(n14678) );
  NAND2_X1 U7936 ( .A1(n14678), .A2(n14677), .ZN(n14676) );
  AOI21_X1 U7937 ( .B1(n7290), .B2(n10593), .A(n6513), .ZN(n7289) );
  INV_X1 U7938 ( .A(n10272), .ZN(n7290) );
  NAND2_X1 U7939 ( .A1(n10077), .A2(n10076), .ZN(n10271) );
  AND3_X1 U7940 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U7941 ( .A1(n6838), .A2(n10091), .ZN(n6627) );
  NAND2_X1 U7942 ( .A1(n6617), .A2(n11544), .ZN(n14695) );
  NAND2_X1 U7943 ( .A1(n9924), .A2(n11877), .ZN(n6617) );
  NAND2_X1 U7944 ( .A1(n9954), .A2(n9953), .ZN(n14704) );
  AND2_X1 U7945 ( .A1(n11715), .A2(n7606), .ZN(n9925) );
  NAND2_X1 U7946 ( .A1(n11859), .A2(n11858), .ZN(n13922) );
  INV_X1 U7947 ( .A(n14609), .ZN(n14762) );
  NOR2_X1 U7948 ( .A1(n14326), .A2(n11869), .ZN(n7534) );
  NAND2_X1 U7949 ( .A1(n11870), .A2(n7533), .ZN(n9569) );
  AND2_X1 U7950 ( .A1(n9270), .A2(n9232), .ZN(n7492) );
  NAND2_X1 U7951 ( .A1(n8976), .A2(n6429), .ZN(n7403) );
  AOI21_X1 U7952 ( .B1(n6429), .B2(n7408), .A(n6604), .ZN(n7404) );
  NAND2_X1 U7953 ( .A1(n14305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9271) );
  XNOR2_X1 U7954 ( .A(n8948), .B(n6598), .ZN(n11834) );
  NAND2_X1 U7955 ( .A1(n7405), .A2(n7406), .ZN(n8948) );
  OR2_X1 U7956 ( .A1(n8976), .A2(n7408), .ZN(n7405) );
  AND2_X1 U7957 ( .A1(n9227), .A2(n9225), .ZN(n6625) );
  AND2_X1 U7958 ( .A1(n9226), .A2(n9228), .ZN(n6624) );
  XNOR2_X1 U7959 ( .A(n8908), .B(n8907), .ZN(n11754) );
  OAI21_X1 U7960 ( .B1(n9220), .B2(n7531), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7535) );
  NAND2_X1 U7961 ( .A1(n7530), .A2(n9123), .ZN(n7527) );
  XNOR2_X1 U7962 ( .A(n8886), .B(n8887), .ZN(n11741) );
  NAND2_X1 U7963 ( .A1(n8829), .A2(n8828), .ZN(n8848) );
  AND3_X1 U7964 ( .A1(n7514), .A2(n7513), .A3(n6478), .ZN(n9120) );
  XNOR2_X1 U7965 ( .A(n8678), .B(n8677), .ZN(n11337) );
  XNOR2_X1 U7966 ( .A(n6878), .B(n8490), .ZN(n10073) );
  XNOR2_X1 U7967 ( .A(n6753), .B(n14379), .ZN(n14382) );
  INV_X1 U7968 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7010) );
  NOR2_X1 U7969 ( .A1(n14409), .A2(n14352), .ZN(n14372) );
  AND2_X1 U7970 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14411), .ZN(n14352) );
  AND2_X1 U7971 ( .A1(n14638), .A2(n14640), .ZN(n14422) );
  INV_X1 U7972 ( .A(n15144), .ZN(n10802) );
  NAND2_X1 U7973 ( .A1(n8164), .A2(n8163), .ZN(n12011) );
  AND4_X1 U7974 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n10758)
         );
  AND4_X1 U7975 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n12181)
         );
  NAND2_X1 U7976 ( .A1(n8050), .A2(n8049), .ZN(n12900) );
  NAND2_X1 U7977 ( .A1(n7320), .A2(n7874), .ZN(n12201) );
  NAND2_X1 U7978 ( .A1(n12279), .A2(n12280), .ZN(n7320) );
  NAND2_X1 U7979 ( .A1(n7886), .A2(n7885), .ZN(n12938) );
  OR2_X1 U7980 ( .A1(n9503), .A2(n8068), .ZN(n7886) );
  NAND2_X1 U7981 ( .A1(n10526), .A2(n10525), .ZN(n10524) );
  NAND2_X1 U7982 ( .A1(n7961), .A2(n7960), .ZN(n12237) );
  OR2_X1 U7983 ( .A1(n12016), .A2(n8068), .ZN(n7961) );
  NAND2_X1 U7984 ( .A1(n8151), .A2(n8150), .ZN(n12281) );
  NAND2_X1 U7985 ( .A1(n6696), .A2(n7263), .ZN(n6792) );
  XNOR2_X1 U7986 ( .A(n6785), .B(n12499), .ZN(n12501) );
  AND2_X1 U7987 ( .A1(n6539), .A2(n12489), .ZN(n6744) );
  AND2_X1 U7988 ( .A1(n7970), .A2(n7969), .ZN(n12816) );
  INV_X1 U7989 ( .A(n12181), .ZN(n11202) );
  NAND4_X1 U7990 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n12515)
         );
  NAND4_X1 U7991 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n12516)
         );
  INV_X1 U7992 ( .A(n10758), .ZN(n12517) );
  INV_X1 U7993 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U7994 ( .A1(n15085), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15084) );
  INV_X1 U7995 ( .A(n9814), .ZN(n10035) );
  OAI22_X1 U7996 ( .A1(n10023), .A2(n10022), .B1(n10035), .B2(n9815), .ZN(
        n9845) );
  INV_X1 U7997 ( .A(n9787), .ZN(n6761) );
  AOI21_X1 U7998 ( .B1(n6942), .B2(n15093), .A(n6537), .ZN(n6940) );
  NAND2_X1 U7999 ( .A1(n10891), .A2(n6495), .ZN(n6941) );
  NAND2_X1 U8000 ( .A1(n7179), .A2(n6593), .ZN(n6918) );
  NOR2_X1 U8001 ( .A1(n12686), .A2(n7191), .ZN(n7190) );
  AND2_X1 U8002 ( .A1(n15106), .A2(n12687), .ZN(n7191) );
  AND2_X1 U8003 ( .A1(n12673), .A2(n12665), .ZN(n6977) );
  NAND2_X1 U8004 ( .A1(n6983), .A2(n6599), .ZN(n6978) );
  NAND2_X1 U8005 ( .A1(n6983), .A2(n6601), .ZN(n6979) );
  XNOR2_X1 U8006 ( .A(n12685), .B(n7189), .ZN(n7188) );
  INV_X1 U8007 ( .A(n12684), .ZN(n7189) );
  AND2_X1 U8008 ( .A1(n6934), .A2(n6932), .ZN(n12685) );
  NOR2_X1 U8009 ( .A1(n12682), .A2(n6933), .ZN(n6932) );
  AND2_X1 U8010 ( .A1(n12300), .A2(n7082), .ZN(n14492) );
  NAND2_X1 U8011 ( .A1(n12297), .A2(n12296), .ZN(n7082) );
  AOI21_X1 U8012 ( .B1(n8223), .B2(n12854), .A(n8222), .ZN(n12148) );
  AND2_X1 U8013 ( .A1(n7415), .A2(n7417), .ZN(n12696) );
  AND2_X1 U8014 ( .A1(n6856), .A2(n7415), .ZN(n12718) );
  NAND2_X1 U8015 ( .A1(n12710), .A2(n12713), .ZN(n6856) );
  NAND2_X1 U8016 ( .A1(n7912), .A2(n7911), .ZN(n12934) );
  NAND2_X1 U8017 ( .A1(n7850), .A2(n7849), .ZN(n14499) );
  OR2_X1 U8018 ( .A1(n15199), .A2(n12896), .ZN(n6875) );
  INV_X1 U8019 ( .A(n12011), .ZN(n12948) );
  NAND2_X1 U8020 ( .A1(n7101), .A2(n8200), .ZN(n11520) );
  NAND2_X1 U8021 ( .A1(n7102), .A2(n6600), .ZN(n7101) );
  XNOR2_X1 U8022 ( .A(n8099), .B(n15324), .ZN(n12331) );
  INV_X1 U8023 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U8024 ( .A1(n8564), .A2(n8563), .ZN(n13024) );
  AND2_X1 U8025 ( .A1(n7112), .A2(n6440), .ZN(n13021) );
  NAND2_X1 U8026 ( .A1(n8774), .A2(n8773), .ZN(n13618) );
  NAND2_X1 U8027 ( .A1(n13678), .A2(n9005), .ZN(n8979) );
  NAND2_X1 U8028 ( .A1(n13094), .A2(n11943), .ZN(n13044) );
  NAND2_X1 U8029 ( .A1(n8812), .A2(n8811), .ZN(n13439) );
  NAND2_X1 U8030 ( .A1(n8611), .A2(n8610), .ZN(n11243) );
  NOR2_X1 U8031 ( .A1(n9099), .A2(n9098), .ZN(n6854) );
  NAND2_X1 U8032 ( .A1(n6653), .A2(n6670), .ZN(n6669) );
  INV_X1 U8033 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U8034 ( .B1(n13247), .B2(n13246), .A(n14930), .ZN(n6780) );
  NAND2_X1 U8035 ( .A1(n7053), .A2(n7056), .ZN(n13342) );
  OR2_X1 U8036 ( .A1(n13365), .A2(n7059), .ZN(n7053) );
  NAND2_X1 U8037 ( .A1(n8831), .A2(n8830), .ZN(n13598) );
  OAI21_X1 U8038 ( .B1(n10744), .B2(n7050), .A(n7048), .ZN(n11039) );
  NAND2_X1 U8039 ( .A1(n10930), .A2(n10929), .ZN(n10932) );
  OAI21_X1 U8040 ( .B1(n8679), .B2(n7139), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6676) );
  NAND2_X1 U8041 ( .A1(n6972), .A2(n10080), .ZN(n11587) );
  NAND2_X1 U8042 ( .A1(n11262), .A2(n11261), .ZN(n11439) );
  NAND2_X1 U8043 ( .A1(n6704), .A2(n12108), .ZN(n13726) );
  NAND2_X1 U8044 ( .A1(n13708), .A2(n12074), .ZN(n13768) );
  NAND2_X1 U8045 ( .A1(n12020), .A2(n7546), .ZN(n13776) );
  OR2_X1 U8046 ( .A1(n12019), .A2(n12018), .ZN(n7546) );
  OAI21_X1 U8047 ( .B1(n11871), .B2(n6764), .A(n6512), .ZN(n6812) );
  NAND2_X1 U8048 ( .A1(n11908), .A2(n6765), .ZN(n6764) );
  INV_X1 U8049 ( .A(n11906), .ZN(n6765) );
  AND2_X1 U8050 ( .A1(n9677), .A2(n9471), .ZN(n11061) );
  NAND2_X1 U8051 ( .A1(n6953), .A2(n6949), .ZN(n14010) );
  AND2_X1 U8052 ( .A1(n6756), .A2(n6584), .ZN(n14208) );
  NAND2_X1 U8053 ( .A1(n14002), .A2(n14751), .ZN(n6756) );
  NAND2_X1 U8054 ( .A1(n6619), .A2(n6618), .ZN(n14022) );
  OAI21_X1 U8055 ( .B1(n6622), .B2(n14570), .A(n6621), .ZN(n6618) );
  NAND2_X1 U8056 ( .A1(n10558), .A2(n10557), .ZN(n14688) );
  NAND2_X1 U8057 ( .A1(n7166), .A2(n7167), .ZN(n6962) );
  XNOR2_X1 U8058 ( .A(n13961), .B(n13992), .ZN(n7169) );
  AND2_X1 U8059 ( .A1(n7150), .A2(n7147), .ZN(n13961) );
  AOI21_X1 U8060 ( .B1(n6431), .B2(n7149), .A(n7148), .ZN(n7147) );
  AND2_X1 U8061 ( .A1(n6963), .A2(n6998), .ZN(n7166) );
  NOR2_X1 U8062 ( .A1(n14200), .A2(n6999), .ZN(n6998) );
  NAND2_X1 U8063 ( .A1(n7002), .A2(n7000), .ZN(n6999) );
  AOI21_X1 U8064 ( .B1(n7166), .B2(n14570), .A(n14763), .ZN(n7165) );
  NAND2_X1 U8065 ( .A1(n13681), .A2(n11791), .ZN(n11793) );
  NOR2_X1 U8066 ( .A1(n14211), .A2(n14210), .ZN(n14274) );
  NAND2_X1 U8067 ( .A1(n14461), .A2(n14460), .ZN(n14459) );
  XNOR2_X1 U8068 ( .A(n14406), .B(n14407), .ZN(n14463) );
  INV_X1 U8069 ( .A(n14635), .ZN(n6798) );
  NAND2_X1 U8070 ( .A1(n14419), .A2(n14420), .ZN(n14641) );
  NAND2_X1 U8071 ( .A1(n14641), .A2(n14642), .ZN(n14638) );
  NAND2_X1 U8072 ( .A1(n6775), .A2(n6774), .ZN(n14640) );
  INV_X1 U8073 ( .A(n14420), .ZN(n6774) );
  INV_X1 U8074 ( .A(n14419), .ZN(n6775) );
  NAND2_X1 U8075 ( .A1(n14422), .A2(n14421), .ZN(n14646) );
  NAND2_X1 U8076 ( .A1(n14646), .A2(n14647), .ZN(n14643) );
  NAND2_X1 U8077 ( .A1(n14478), .A2(n14425), .ZN(n14485) );
  OAI21_X1 U8078 ( .B1(n14485), .B2(n14484), .A(n7023), .ZN(n7022) );
  INV_X1 U8079 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U8080 ( .A1(n11588), .A2(n7501), .ZN(n7500) );
  NAND3_X1 U8081 ( .A1(n8357), .A2(n8358), .A3(n8356), .ZN(n6648) );
  NAND2_X1 U8082 ( .A1(n11598), .A2(n11600), .ZN(n7475) );
  INV_X1 U8083 ( .A(n8406), .ZN(n6637) );
  NAND2_X1 U8084 ( .A1(n11610), .A2(n11612), .ZN(n7473) );
  INV_X1 U8085 ( .A(n8433), .ZN(n8436) );
  NOR2_X1 U8086 ( .A1(n11891), .A2(n7469), .ZN(n7468) );
  NOR2_X1 U8087 ( .A1(n11620), .A2(n11621), .ZN(n7469) );
  NAND2_X1 U8088 ( .A1(n6630), .A2(n7450), .ZN(n8526) );
  NAND2_X1 U8089 ( .A1(n8507), .A2(n6448), .ZN(n7450) );
  NAND2_X1 U8090 ( .A1(n6631), .A2(n6486), .ZN(n6628) );
  NOR2_X1 U8091 ( .A1(n11647), .A2(n7484), .ZN(n7483) );
  OAI21_X1 U8092 ( .B1(n7537), .B2(n7486), .A(n7485), .ZN(n7484) );
  NAND2_X1 U8093 ( .A1(n11630), .A2(n11648), .ZN(n7485) );
  NAND2_X1 U8094 ( .A1(n6634), .A2(n6504), .ZN(n8577) );
  NAND2_X1 U8095 ( .A1(n8577), .A2(n8576), .ZN(n6633) );
  NOR2_X1 U8096 ( .A1(n11687), .A2(n11684), .ZN(n7480) );
  NAND2_X1 U8097 ( .A1(n11687), .A2(n11684), .ZN(n7479) );
  NAND2_X1 U8098 ( .A1(n7480), .A2(n7479), .ZN(n7478) );
  AOI21_X1 U8099 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n6665) );
  OAI21_X1 U8100 ( .B1(n8601), .B2(n8600), .A(n6532), .ZN(n6664) );
  NAND2_X1 U8101 ( .A1(n6814), .A2(n7493), .ZN(n11731) );
  NAND2_X1 U8102 ( .A1(n11716), .A2(n7494), .ZN(n7493) );
  INV_X1 U8103 ( .A(n8693), .ZN(n7459) );
  INV_X1 U8104 ( .A(n12739), .ZN(n6794) );
  NAND2_X1 U8105 ( .A1(n6671), .A2(n6641), .ZN(n8784) );
  NAND2_X1 U8106 ( .A1(n6640), .A2(n6638), .ZN(n6641) );
  AND2_X1 U8107 ( .A1(n6639), .A2(n7461), .ZN(n6638) );
  NAND2_X1 U8108 ( .A1(n11794), .A2(n7496), .ZN(n7495) );
  AOI21_X1 U8109 ( .B1(n11778), .B2(n11779), .A(n6813), .ZN(n6843) );
  AND2_X1 U8110 ( .A1(n8894), .A2(SI_26_), .ZN(n7401) );
  NOR2_X1 U8111 ( .A1(n7866), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U8112 ( .A1(n7445), .A2(n7444), .ZN(n7443) );
  INV_X1 U8113 ( .A(n8884), .ZN(n7444) );
  INV_X1 U8114 ( .A(n8885), .ZN(n7445) );
  OAI21_X1 U8115 ( .B1(n6651), .B2(n6650), .A(n7451), .ZN(n6663) );
  NAND2_X1 U8116 ( .A1(n7452), .A2(n6575), .ZN(n7451) );
  INV_X1 U8117 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7458) );
  INV_X1 U8118 ( .A(n7393), .ZN(n7390) );
  INV_X1 U8119 ( .A(n7401), .ZN(n7395) );
  NOR2_X1 U8120 ( .A1(n8766), .A2(SI_18_), .ZN(n7386) );
  NOR2_X1 U8121 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  INV_X1 U8122 ( .A(n8749), .ZN(n7385) );
  INV_X1 U8123 ( .A(n7364), .ZN(n7363) );
  OAI21_X1 U8124 ( .B1(n7554), .B2(n7365), .A(n7536), .ZN(n7364) );
  INV_X1 U8125 ( .A(n8670), .ZN(n8698) );
  NAND2_X1 U8126 ( .A1(n8627), .A2(n14450), .ZN(n8653) );
  INV_X1 U8127 ( .A(n8603), .ZN(n7380) );
  NAND2_X1 U8128 ( .A1(n8605), .A2(n9191), .ZN(n8625) );
  NAND2_X1 U8129 ( .A1(n14333), .A2(n14334), .ZN(n14335) );
  NOR2_X1 U8130 ( .A1(n7812), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U8131 ( .A1(n6763), .A2(n6762), .ZN(n7629) );
  INV_X1 U8132 ( .A(n9151), .ZN(n6762) );
  INV_X1 U8133 ( .A(n8068), .ZN(n6763) );
  AND2_X1 U8134 ( .A1(n7963), .A2(n7962), .ZN(n7981) );
  AND2_X1 U8135 ( .A1(n7887), .A2(n12203), .ZN(n7898) );
  NAND2_X1 U8136 ( .A1(n6742), .A2(n6741), .ZN(n12477) );
  INV_X1 U8137 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7337) );
  INV_X1 U8138 ( .A(n12645), .ZN(n6937) );
  OR2_X1 U8139 ( .A1(n8255), .A2(n8210), .ZN(n12494) );
  OR2_X1 U8140 ( .A1(n12011), .A2(n12715), .ZN(n12482) );
  OR2_X1 U8141 ( .A1(n8199), .A2(n12726), .ZN(n12478) );
  NOR2_X1 U8142 ( .A1(n8035), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8052) );
  NOR2_X1 U8143 ( .A1(n12767), .A2(n7257), .ZN(n7256) );
  INV_X1 U8144 ( .A(n12461), .ZN(n7257) );
  INV_X1 U8145 ( .A(n12329), .ZN(n7259) );
  OR2_X1 U8146 ( .A1(n8000), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8019) );
  INV_X1 U8147 ( .A(n12450), .ZN(n7284) );
  AOI21_X1 U8148 ( .B1(n11402), .B2(n7422), .A(n6518), .ZN(n7421) );
  INV_X1 U8149 ( .A(n8182), .ZN(n7422) );
  OR2_X1 U8150 ( .A1(n7790), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U8151 ( .A1(n7746), .A2(n7745), .ZN(n7771) );
  NAND2_X1 U8152 ( .A1(n6605), .A2(n11522), .ZN(n7098) );
  INV_X1 U8153 ( .A(n8200), .ZN(n7100) );
  INV_X1 U8154 ( .A(n11521), .ZN(n7103) );
  INV_X1 U8155 ( .A(n7875), .ZN(n6735) );
  INV_X1 U8156 ( .A(n7096), .ZN(n7095) );
  OAI21_X1 U8157 ( .B1(n7878), .B2(n7097), .A(n7916), .ZN(n7096) );
  INV_X1 U8158 ( .A(n7903), .ZN(n7097) );
  INV_X1 U8159 ( .A(n7858), .ZN(n6736) );
  NAND2_X1 U8160 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U8161 ( .A1(n7823), .A2(n11059), .ZN(n7844) );
  INV_X1 U8162 ( .A(n7701), .ZN(n6725) );
  AND2_X1 U8163 ( .A1(n9179), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7716) );
  INV_X1 U8164 ( .A(n7699), .ZN(n6722) );
  AND2_X1 U8165 ( .A1(n8439), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8462) );
  OR2_X1 U8166 ( .A1(n13558), .A2(n13124), .ZN(n9051) );
  NOR2_X1 U8167 ( .A1(n13450), .A2(n13439), .ZN(n7039) );
  INV_X1 U8168 ( .A(n7253), .ZN(n7245) );
  OR2_X1 U8169 ( .A1(n8756), .A2(n8755), .ZN(n8776) );
  INV_X1 U8170 ( .A(n11513), .ZN(n7206) );
  INV_X1 U8171 ( .A(n11177), .ZN(n7231) );
  NOR2_X1 U8172 ( .A1(n11031), .A2(n7229), .ZN(n7228) );
  NOR2_X1 U8173 ( .A1(n7229), .A2(n7225), .ZN(n7224) );
  INV_X1 U8174 ( .A(n10924), .ZN(n7225) );
  INV_X1 U8175 ( .A(n13136), .ZN(n11172) );
  INV_X1 U8176 ( .A(n10723), .ZN(n7238) );
  NOR2_X1 U8177 ( .A1(n7238), .A2(n7237), .ZN(n7236) );
  INV_X1 U8178 ( .A(n10394), .ZN(n7237) );
  INV_X1 U8179 ( .A(n7037), .ZN(n13412) );
  NAND2_X1 U8180 ( .A1(n8292), .A2(n8291), .ZN(n8312) );
  INV_X1 U8181 ( .A(n12060), .ZN(n7512) );
  NAND2_X1 U8182 ( .A1(n13812), .A2(n6710), .ZN(n6711) );
  AND2_X1 U8183 ( .A1(n13811), .A2(n12053), .ZN(n6710) );
  AND2_X1 U8184 ( .A1(n13792), .A2(n7511), .ZN(n7510) );
  OR2_X1 U8185 ( .A1(n13752), .A2(n7512), .ZN(n7511) );
  NAND2_X1 U8186 ( .A1(n9560), .A2(n11863), .ZN(n9563) );
  INV_X1 U8187 ( .A(n6802), .ZN(n6626) );
  NOR2_X1 U8188 ( .A1(n6996), .A2(n14205), .ZN(n6995) );
  INV_X1 U8189 ( .A(n6997), .ZN(n6996) );
  NAND2_X1 U8190 ( .A1(n14039), .A2(n6957), .ZN(n6955) );
  NOR2_X1 U8191 ( .A1(n14038), .A2(n14026), .ZN(n6997) );
  INV_X1 U8192 ( .A(n14160), .ZN(n6614) );
  AND2_X1 U8193 ( .A1(n14126), .A2(n6474), .ZN(n7160) );
  NOR2_X1 U8194 ( .A1(n14584), .A2(n14303), .ZN(n14138) );
  NAND2_X1 U8195 ( .A1(n11161), .A2(n11629), .ZN(n7174) );
  INV_X1 U8196 ( .A(n11159), .ZN(n6610) );
  NOR2_X1 U8197 ( .A1(n14183), .A2(n11609), .ZN(n10982) );
  NOR2_X1 U8198 ( .A1(n14687), .A2(n14688), .ZN(n6751) );
  INV_X1 U8199 ( .A(n7313), .ZN(n7312) );
  OAI21_X1 U8200 ( .B1(n7314), .B2(n9955), .A(n9956), .ZN(n7313) );
  NAND2_X1 U8201 ( .A1(n13835), .A2(n6990), .ZN(n11555) );
  NAND2_X1 U8202 ( .A1(n9596), .A2(n11546), .ZN(n11540) );
  INV_X1 U8203 ( .A(n7154), .ZN(n7153) );
  NOR2_X1 U8204 ( .A1(n11161), .A2(n6968), .ZN(n6967) );
  INV_X1 U8205 ( .A(n6970), .ZN(n6968) );
  NAND2_X1 U8206 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  NAND2_X1 U8207 ( .A1(n11068), .A2(n11069), .ZN(n11158) );
  AOI21_X1 U8208 ( .B1(n7409), .B2(n7407), .A(n6596), .ZN(n7406) );
  INV_X1 U8209 ( .A(n8938), .ZN(n7407) );
  AND2_X1 U8210 ( .A1(n7396), .A2(n7394), .ZN(n7393) );
  NAND2_X1 U8211 ( .A1(n7402), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U8212 ( .A1(n7399), .A2(n7395), .ZN(n7394) );
  INV_X1 U8213 ( .A(n8894), .ZN(n7397) );
  INV_X1 U8214 ( .A(n8908), .ZN(n7392) );
  NOR2_X1 U8215 ( .A1(n7375), .A2(SI_24_), .ZN(n7374) );
  INV_X1 U8216 ( .A(n8868), .ZN(n7375) );
  AND2_X1 U8217 ( .A1(n7369), .A2(n8847), .ZN(n7367) );
  NAND2_X1 U8218 ( .A1(n8810), .A2(n8809), .ZN(n8826) );
  NAND2_X1 U8219 ( .A1(n8675), .A2(SI_15_), .ZN(n8701) );
  XNOR2_X1 U8220 ( .A(n8556), .B(SI_9_), .ZN(n8553) );
  XNOR2_X1 U8221 ( .A(n8535), .B(SI_8_), .ZN(n8532) );
  AOI21_X1 U8222 ( .B1(n7357), .B2(n7358), .A(n6523), .ZN(n7355) );
  INV_X1 U8223 ( .A(n8493), .ZN(n7358) );
  OAI21_X1 U8224 ( .B1(n11713), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n6877), .ZN(
        n8451) );
  OR2_X1 U8225 ( .A1(n8330), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6877) );
  INV_X1 U8226 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U8227 ( .A1(n8376), .A2(n9152), .ZN(n6866) );
  NAND2_X1 U8228 ( .A1(n14346), .A2(n14345), .ZN(n14401) );
  AOI21_X1 U8229 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14350), .A(n14349), .ZN(
        n14351) );
  NOR2_X1 U8230 ( .A1(n14374), .A2(n14373), .ZN(n14349) );
  OR2_X1 U8231 ( .A1(n7837), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7866) );
  AOI21_X1 U8232 ( .B1(n8098), .B2(n8079), .A(n12004), .ZN(n6906) );
  INV_X1 U8233 ( .A(n6906), .ZN(n6904) );
  NAND2_X1 U8234 ( .A1(n7340), .A2(n12219), .ZN(n6897) );
  NAND2_X1 U8235 ( .A1(n10997), .A2(n7349), .ZN(n7348) );
  INV_X1 U8236 ( .A(n7551), .ZN(n7349) );
  NAND2_X1 U8237 ( .A1(n7971), .A2(n12816), .ZN(n12167) );
  NAND2_X1 U8238 ( .A1(n7683), .A2(n7682), .ZN(n7691) );
  INV_X1 U8239 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7682) );
  INV_X1 U8240 ( .A(n12500), .ZN(n7263) );
  NAND2_X1 U8241 ( .A1(n12498), .A2(n12690), .ZN(n7083) );
  NAND2_X1 U8242 ( .A1(n14492), .A2(n12507), .ZN(n7081) );
  NOR2_X1 U8243 ( .A1(n12326), .A2(n12325), .ZN(n12497) );
  AND4_X1 U8244 ( .A1(n7638), .A2(n7637), .A3(n7636), .A4(n7635), .ZN(n9869)
         );
  OR2_X1 U8245 ( .A1(n10050), .A2(n9827), .ZN(n6928) );
  AND2_X1 U8246 ( .A1(n6928), .A2(n6435), .ZN(n10039) );
  NAND2_X1 U8247 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n6921), .ZN(n7548) );
  NOR2_X1 U8248 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n6921) );
  NOR2_X1 U8249 ( .A1(n10039), .A2(n7184), .ZN(n10009) );
  INV_X1 U8250 ( .A(n6984), .ZN(n10909) );
  INV_X1 U8251 ( .A(n6942), .ZN(n6939) );
  NOR2_X1 U8252 ( .A1(n6943), .A2(n14449), .ZN(n6942) );
  INV_X1 U8253 ( .A(n10892), .ZN(n6943) );
  NOR2_X1 U8254 ( .A1(n10904), .A2(n10905), .ZN(n11315) );
  NAND2_X1 U8255 ( .A1(n15123), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U8256 ( .A1(n12535), .A2(n6591), .ZN(n12556) );
  AOI21_X1 U8257 ( .B1(n9796), .B2(n12567), .A(n6454), .ZN(n6867) );
  NAND2_X1 U8258 ( .A1(n7337), .A2(n7847), .ZN(n7333) );
  OR2_X1 U8259 ( .A1(n12605), .A2(n12604), .ZN(n12617) );
  NAND2_X1 U8260 ( .A1(n12643), .A2(n6937), .ZN(n6935) );
  NAND2_X1 U8261 ( .A1(n6982), .A2(n12673), .ZN(n6981) );
  NAND2_X1 U8262 ( .A1(n12638), .A2(n12665), .ZN(n6982) );
  INV_X1 U8263 ( .A(n6935), .ZN(n6933) );
  OR2_X1 U8264 ( .A1(n12619), .A2(n6936), .ZN(n6934) );
  NAND2_X1 U8265 ( .A1(n6937), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6936) );
  AND2_X1 U8266 ( .A1(n8134), .A2(n8133), .ZN(n12688) );
  NAND2_X1 U8267 ( .A1(n7266), .A2(n6473), .ZN(n7265) );
  NAND2_X1 U8268 ( .A1(n6745), .A2(n12471), .ZN(n7266) );
  OR2_X1 U8269 ( .A1(n8019), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U8270 ( .A1(n12763), .A2(n12762), .ZN(n12765) );
  NAND2_X1 U8271 ( .A1(n7261), .A2(n12460), .ZN(n12763) );
  OAI21_X1 U8272 ( .B1(n12836), .B2(n7436), .A(n6533), .ZN(n12799) );
  NAND2_X1 U8273 ( .A1(n7435), .A2(n6679), .ZN(n6678) );
  INV_X1 U8274 ( .A(n7433), .ZN(n7432) );
  OR2_X1 U8275 ( .A1(n12824), .A2(n7436), .ZN(n12813) );
  NAND2_X1 U8276 ( .A1(n12836), .A2(n8189), .ZN(n12825) );
  NOR2_X1 U8277 ( .A1(n12825), .A2(n12826), .ZN(n12824) );
  AND2_X1 U8278 ( .A1(n12422), .A2(n12429), .ZN(n12859) );
  NAND2_X1 U8279 ( .A1(n8186), .A2(n8187), .ZN(n12852) );
  OAI21_X1 U8280 ( .B1(n11401), .B2(n11402), .A(n12418), .ZN(n12878) );
  AND2_X1 U8281 ( .A1(n12423), .A2(n12861), .ZN(n12877) );
  OAI21_X1 U8282 ( .B1(n8183), .B2(n7423), .A(n7421), .ZN(n12870) );
  AND2_X1 U8283 ( .A1(n7272), .A2(n8229), .ZN(n7271) );
  NAND2_X1 U8284 ( .A1(n7274), .A2(n7273), .ZN(n7272) );
  NAND2_X1 U8285 ( .A1(n10422), .A2(n8173), .ZN(n10319) );
  NAND2_X1 U8286 ( .A1(n6693), .A2(n12341), .ZN(n10853) );
  INV_X1 U8287 ( .A(n12356), .ZN(n12307) );
  NAND2_X1 U8288 ( .A1(n8166), .A2(n8165), .ZN(n9863) );
  OAI21_X1 U8289 ( .B1(n12338), .B2(n15140), .A(n12344), .ZN(n6702) );
  NAND2_X1 U8290 ( .A1(n15142), .A2(n10380), .ZN(n15139) );
  OR2_X1 U8291 ( .A1(n12299), .A2(SI_2_), .ZN(n7652) );
  OR2_X1 U8292 ( .A1(n11199), .A2(n8068), .ZN(n8070) );
  NAND2_X1 U8293 ( .A1(n7979), .A2(n7978), .ZN(n12453) );
  OR2_X1 U8294 ( .A1(n10249), .A2(n8068), .ZN(n7979) );
  NAND2_X1 U8295 ( .A1(n7926), .A2(n7925), .ZN(n8190) );
  OR2_X1 U8296 ( .A1(n9682), .A2(n8068), .ZN(n7926) );
  AND2_X1 U8297 ( .A1(n12771), .A2(n12893), .ZN(n15179) );
  NAND2_X1 U8298 ( .A1(n7277), .A2(n8228), .ZN(n10955) );
  OAI211_X1 U8299 ( .C1(n8140), .C2(n10335), .A(n7735), .B(n7734), .ZN(n12384)
         );
  OAI21_X1 U8300 ( .B1(n7098), .B2(n6729), .A(n12291), .ZN(n6728) );
  NAND2_X1 U8301 ( .A1(n8065), .A2(n11742), .ZN(n7105) );
  OR2_X1 U8302 ( .A1(n7569), .A2(n12990), .ZN(n7570) );
  OAI21_X1 U8303 ( .B1(n7843), .B2(n9465), .A(n7844), .ZN(n7856) );
  BUF_X1 U8304 ( .A(n7805), .Z(n7806) );
  XNOR2_X1 U8305 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7763) );
  INV_X1 U8306 ( .A(n7729), .ZN(n7730) );
  XNOR2_X1 U8307 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7753) );
  INV_X1 U8308 ( .A(n7663), .ZN(n6717) );
  AND2_X1 U8309 ( .A1(n6715), .A2(n7612), .ZN(n6714) );
  NAND2_X1 U8310 ( .A1(n9143), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7612) );
  XNOR2_X1 U8311 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7676) );
  NAND2_X1 U8312 ( .A1(n12990), .A2(n7559), .ZN(n6880) );
  NAND2_X1 U8313 ( .A1(n7647), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8314 ( .A1(n8331), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U8315 ( .A1(n8499), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8515) );
  NOR2_X1 U8316 ( .A1(n10482), .A2(n10483), .ZN(n7132) );
  OR2_X1 U8317 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  NOR2_X1 U8318 ( .A1(n8776), .A2(n8775), .ZN(n8814) );
  NOR2_X1 U8319 ( .A1(n8874), .A2(n8873), .ZN(n8913) );
  AND2_X1 U8320 ( .A1(n11966), .A2(n11964), .ZN(n13050) );
  NOR2_X1 U8321 ( .A1(n8712), .A2(n8711), .ZN(n8738) );
  NAND2_X1 U8322 ( .A1(n13097), .A2(n11953), .ZN(n7123) );
  AND2_X1 U8323 ( .A1(n13097), .A2(n6547), .ZN(n13071) );
  OR2_X1 U8324 ( .A1(n11954), .A2(n13010), .ZN(n7124) );
  INV_X1 U8325 ( .A(n7126), .ZN(n7122) );
  AND2_X1 U8326 ( .A1(n11960), .A2(n11959), .ZN(n13072) );
  NAND2_X1 U8327 ( .A1(n7133), .A2(n7131), .ZN(n7135) );
  AND2_X1 U8328 ( .A1(n8613), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U8329 ( .A1(n8635), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8658) );
  NOR2_X1 U8330 ( .A1(n13311), .A2(n13496), .ZN(n7126) );
  NOR2_X1 U8331 ( .A1(n8591), .A2(n9541), .ZN(n8613) );
  AND2_X1 U8332 ( .A1(n8462), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8499) );
  INV_X1 U8333 ( .A(n8912), .ZN(n8899) );
  NAND2_X1 U8334 ( .A1(n8316), .A2(n10946), .ZN(n9651) );
  AND2_X1 U8335 ( .A1(n7439), .A2(n9044), .ZN(n6851) );
  AND2_X1 U8336 ( .A1(n7440), .A2(n8992), .ZN(n7439) );
  INV_X1 U8337 ( .A(n6410), .ZN(n8964) );
  NAND2_X1 U8338 ( .A1(n13162), .A2(n13161), .ZN(n13172) );
  NAND2_X1 U8339 ( .A1(n9338), .A2(n9337), .ZN(n14816) );
  NAND2_X1 U8340 ( .A1(n9343), .A2(n9342), .ZN(n13192) );
  OR2_X1 U8341 ( .A1(n14836), .A2(n14835), .ZN(n14838) );
  INV_X1 U8342 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8287) );
  INV_X1 U8343 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8286) );
  XNOR2_X1 U8344 ( .A(n13218), .B(n13219), .ZN(n14875) );
  NAND2_X1 U8345 ( .A1(n14875), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14874) );
  XNOR2_X1 U8346 ( .A(n13221), .B(n13231), .ZN(n14886) );
  NAND2_X1 U8347 ( .A1(n14886), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14885) );
  INV_X1 U8348 ( .A(n7140), .ZN(n7138) );
  NOR2_X1 U8349 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14918), .ZN(n14919) );
  NAND2_X1 U8350 ( .A1(n8950), .A2(n8949), .ZN(n13253) );
  INV_X1 U8351 ( .A(n13320), .ZN(n7057) );
  NAND2_X1 U8352 ( .A1(n6771), .A2(n6770), .ZN(n13450) );
  INV_X1 U8353 ( .A(n7039), .ZN(n13440) );
  OR2_X1 U8354 ( .A1(n13449), .A2(n13309), .ZN(n6767) );
  OAI21_X1 U8355 ( .B1(n13504), .B2(n7246), .A(n7244), .ZN(n13458) );
  INV_X1 U8356 ( .A(n7248), .ZN(n7246) );
  AOI21_X1 U8357 ( .B1(n7248), .B2(n7245), .A(n6487), .ZN(n7244) );
  NOR2_X1 U8358 ( .A1(n7250), .A2(n13275), .ZN(n7248) );
  NAND2_X1 U8359 ( .A1(n11427), .A2(n7036), .ZN(n7035) );
  NOR2_X1 U8360 ( .A1(n11192), .A2(n7034), .ZN(n11248) );
  INV_X1 U8361 ( .A(n7036), .ZN(n7034) );
  AOI21_X1 U8362 ( .B1(n7048), .B2(n7050), .A(n6484), .ZN(n7046) );
  NAND2_X1 U8363 ( .A1(n7226), .A2(n11034), .ZN(n11171) );
  NAND2_X1 U8364 ( .A1(n11032), .A2(n11031), .ZN(n7226) );
  INV_X1 U8365 ( .A(n10929), .ZN(n7050) );
  NAND2_X1 U8366 ( .A1(n10925), .A2(n10924), .ZN(n11032) );
  NAND2_X1 U8367 ( .A1(n10744), .A2(n10743), .ZN(n10930) );
  INV_X1 U8368 ( .A(n7045), .ZN(n7044) );
  OAI21_X1 U8369 ( .B1(n6462), .B2(n10388), .A(n10443), .ZN(n7045) );
  AND2_X1 U8370 ( .A1(n7032), .A2(n14995), .ZN(n7031) );
  NAND2_X1 U8371 ( .A1(n10545), .A2(n10543), .ZN(n10390) );
  NAND2_X1 U8372 ( .A1(n10538), .A2(n14995), .ZN(n10537) );
  NAND2_X1 U8373 ( .A1(n9090), .A2(n13690), .ZN(n8352) );
  AND2_X1 U8374 ( .A1(n13555), .A2(n15053), .ZN(n7240) );
  INV_X1 U8375 ( .A(n13439), .ZN(n13604) );
  NAND2_X1 U8376 ( .A1(n7207), .A2(n11513), .ZN(n13264) );
  NAND2_X1 U8377 ( .A1(n10608), .A2(n10151), .ZN(n10153) );
  INV_X1 U8378 ( .A(n7108), .ZN(n15064) );
  OR2_X1 U8379 ( .A1(n9661), .A2(n9660), .ZN(n9764) );
  INV_X1 U8380 ( .A(n7457), .ZN(n7027) );
  OR2_X1 U8381 ( .A1(n9079), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9081) );
  OR2_X1 U8382 ( .A1(n8495), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8538) );
  OR2_X1 U8383 ( .A1(n8479), .A2(n8478), .ZN(n8481) );
  INV_X1 U8384 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8416) );
  INV_X1 U8385 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8386 ( .A1(n6829), .A2(n10784), .ZN(n6828) );
  INV_X1 U8387 ( .A(n10786), .ZN(n6829) );
  INV_X1 U8388 ( .A(n14019), .ZN(n13960) );
  INV_X1 U8389 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U8390 ( .A1(n11720), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11735) );
  INV_X1 U8391 ( .A(n7522), .ZN(n7521) );
  INV_X1 U8392 ( .A(n9724), .ZN(n12039) );
  NAND2_X1 U8393 ( .A1(n13766), .A2(n6502), .ZN(n13716) );
  NAND2_X1 U8394 ( .A1(n11646), .A2(n11645), .ZN(n13749) );
  NAND2_X1 U8395 ( .A1(n11346), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11386) );
  OR2_X1 U8396 ( .A1(n10284), .A2(n10283), .ZN(n10566) );
  OR2_X1 U8397 ( .A1(n10566), .A2(n10565), .ZN(n10578) );
  XNOR2_X1 U8398 ( .A(n9725), .B(n9724), .ZN(n10187) );
  OAI22_X1 U8399 ( .A1(n11552), .A2(n9563), .B1(n11556), .B2(n12047), .ZN(
        n9725) );
  NAND2_X1 U8400 ( .A1(n13751), .A2(n13752), .ZN(n13750) );
  NOR2_X1 U8401 ( .A1(n11072), .A2(n11071), .ZN(n11153) );
  AND2_X1 U8402 ( .A1(n11153), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11346) );
  AOI21_X1 U8403 ( .B1(n13922), .B2(n11867), .A(n7353), .ZN(n7352) );
  NAND2_X1 U8404 ( .A1(n14268), .A2(n11868), .ZN(n7354) );
  NOR2_X1 U8405 ( .A1(n11867), .A2(n11868), .ZN(n7353) );
  INV_X1 U8406 ( .A(n6802), .ZN(n11817) );
  INV_X1 U8407 ( .A(n7465), .ZN(n7464) );
  OAI22_X1 U8408 ( .A1(n6802), .A2(n9478), .B1(n11820), .B2(n9284), .ZN(n7465)
         );
  NOR2_X1 U8409 ( .A1(n6491), .A2(n7463), .ZN(n7462) );
  AND3_X1 U8410 ( .A1(n9275), .A2(n9276), .A3(P1_REG3_REG_0__SCAN_IN), .ZN(
        n7463) );
  NAND2_X1 U8411 ( .A1(n14030), .A2(n6954), .ZN(n6949) );
  INV_X1 U8412 ( .A(n6955), .ZN(n6954) );
  AND2_X1 U8413 ( .A1(n6958), .A2(n14018), .ZN(n6956) );
  AOI21_X1 U8414 ( .B1(n14017), .B2(n14762), .A(n7155), .ZN(n6621) );
  NAND2_X1 U8415 ( .A1(n6620), .A2(n6750), .ZN(n6619) );
  AND2_X1 U8416 ( .A1(n6839), .A2(n7155), .ZN(n6750) );
  NAND2_X1 U8417 ( .A1(n14016), .A2(n14762), .ZN(n6839) );
  NAND2_X1 U8418 ( .A1(n14044), .A2(n14280), .ZN(n14035) );
  INV_X1 U8419 ( .A(n11735), .ZN(n11736) );
  NAND2_X1 U8420 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11736), .ZN(n11748) );
  INV_X1 U8421 ( .A(n6992), .ZN(n14083) );
  AOI21_X1 U8422 ( .B1(n7298), .B2(n7297), .A(n6517), .ZN(n7296) );
  INV_X1 U8423 ( .A(n7301), .ZN(n7297) );
  NAND2_X1 U8424 ( .A1(n14097), .A2(n14238), .ZN(n14098) );
  AND2_X1 U8425 ( .A1(n11674), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11688) );
  NOR2_X1 U8426 ( .A1(n14130), .A2(n14292), .ZN(n14097) );
  AND2_X1 U8427 ( .A1(n11663), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U8428 ( .A1(n13942), .A2(n13941), .ZN(n14142) );
  NOR2_X1 U8429 ( .A1(n11636), .A2(n11635), .ZN(n11663) );
  OR2_X1 U8430 ( .A1(n11386), .A2(n11385), .ZN(n11636) );
  AND2_X1 U8431 ( .A1(n7003), .A2(n13973), .ZN(n14585) );
  NAND2_X1 U8432 ( .A1(n14585), .A2(n14591), .ZN(n14584) );
  INV_X1 U8433 ( .A(n13936), .ZN(n14569) );
  NAND2_X1 U8434 ( .A1(n11379), .A2(n11378), .ZN(n13934) );
  INV_X1 U8435 ( .A(n7003), .ZN(n11384) );
  OR2_X1 U8436 ( .A1(n10969), .A2(n10968), .ZN(n11072) );
  NOR2_X1 U8437 ( .A1(n10578), .A2(n10577), .ZN(n10585) );
  NAND2_X1 U8438 ( .A1(n6751), .A2(n6993), .ZN(n14183) );
  INV_X1 U8439 ( .A(n6751), .ZN(n14689) );
  NAND2_X1 U8440 ( .A1(n10277), .A2(n10278), .ZN(n14687) );
  NOR2_X1 U8441 ( .A1(n10083), .A2(n10082), .ZN(n10095) );
  NOR2_X1 U8442 ( .A1(n10122), .A2(n11587), .ZN(n10277) );
  NAND2_X1 U8443 ( .A1(n9957), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U8444 ( .A1(n10123), .A2(n10138), .ZN(n10122) );
  AND2_X1 U8445 ( .A1(n14731), .A2(n14710), .ZN(n10116) );
  AND2_X1 U8446 ( .A1(n10116), .A2(n10065), .ZN(n10123) );
  AND2_X1 U8447 ( .A1(n11552), .A2(n6989), .ZN(n14710) );
  AND2_X1 U8448 ( .A1(n6990), .A2(n9908), .ZN(n6989) );
  NAND2_X1 U8449 ( .A1(n11540), .A2(n11547), .ZN(n9924) );
  INV_X1 U8450 ( .A(n11877), .ZN(n9951) );
  NAND2_X1 U8451 ( .A1(n11552), .A2(n9908), .ZN(n14706) );
  INV_X1 U8452 ( .A(n7157), .ZN(n7156) );
  NAND2_X1 U8453 ( .A1(n7154), .A2(n7152), .ZN(n7151) );
  OAI21_X1 U8454 ( .B1(n14018), .B2(n7158), .A(n6481), .ZN(n7157) );
  AND2_X1 U8455 ( .A1(n7153), .A2(n6470), .ZN(n7149) );
  NOR2_X1 U8456 ( .A1(n14205), .A2(n13960), .ZN(n7148) );
  NAND2_X1 U8457 ( .A1(n14202), .A2(n14755), .ZN(n7002) );
  AND2_X1 U8458 ( .A1(n6573), .A2(n7001), .ZN(n7000) );
  INV_X1 U8459 ( .A(n14201), .ZN(n7001) );
  NAND2_X1 U8460 ( .A1(n11683), .A2(n11682), .ZN(n14132) );
  NAND2_X1 U8461 ( .A1(n11342), .A2(n11341), .ZN(n12036) );
  NOR2_X1 U8462 ( .A1(n7146), .A2(n7145), .ZN(n7144) );
  INV_X1 U8463 ( .A(n10559), .ZN(n7145) );
  NAND2_X1 U8464 ( .A1(n14676), .A2(n10559), .ZN(n14180) );
  NAND2_X1 U8465 ( .A1(n7172), .A2(n10280), .ZN(n10281) );
  AND2_X1 U8466 ( .A1(n14707), .A2(n14184), .ZN(n9687) );
  AND2_X1 U8467 ( .A1(n9264), .A2(n9263), .ZN(n13966) );
  MUX2_X1 U8468 ( .A(n13842), .B(n14327), .S(n11715), .Z(n9906) );
  NAND2_X1 U8469 ( .A1(n15268), .A2(n9798), .ZN(n6922) );
  INV_X1 U8470 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7529) );
  INV_X1 U8471 ( .A(n7531), .ZN(n7530) );
  NAND2_X1 U8472 ( .A1(n9220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U8473 ( .A(n7388), .B(SI_18_), .ZN(n8767) );
  NAND2_X1 U8474 ( .A1(n8750), .A2(n8749), .ZN(n7388) );
  OAI21_X1 U8475 ( .B1(n6784), .B2(n8578), .A(n7381), .ZN(n8604) );
  OR2_X1 U8476 ( .A1(n9643), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9196) );
  XNOR2_X1 U8477 ( .A(n8580), .B(n8578), .ZN(n10560) );
  NAND2_X1 U8478 ( .A1(n6784), .A2(n8557), .ZN(n8580) );
  OR2_X1 U8479 ( .A1(n9186), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9643) );
  NAND2_X1 U8480 ( .A1(n6944), .A2(n8493), .ZN(n8509) );
  NAND2_X1 U8481 ( .A1(n6878), .A2(n8491), .ZN(n6944) );
  INV_X1 U8482 ( .A(n8490), .ZN(n8491) );
  XNOR2_X1 U8483 ( .A(n8451), .B(SI_4_), .ZN(n8449) );
  NAND2_X1 U8484 ( .A1(n9130), .A2(n9118), .ZN(n9139) );
  NAND2_X1 U8485 ( .A1(n14330), .A2(n7014), .ZN(n14378) );
  NAND2_X1 U8486 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7015), .ZN(n7014) );
  INV_X1 U8487 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7015) );
  XNOR2_X1 U8488 ( .A(n14389), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14391) );
  NOR2_X1 U8489 ( .A1(n15355), .A2(n14388), .ZN(n14390) );
  NAND2_X1 U8490 ( .A1(n14340), .A2(n14339), .ZN(n14395) );
  NOR2_X1 U8491 ( .A1(n15362), .A2(n14400), .ZN(n14403) );
  OAI21_X1 U8492 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14355), .A(n14354), .ZN(
        n14370) );
  OR2_X1 U8493 ( .A1(n12241), .A2(n12240), .ZN(n6889) );
  INV_X1 U8494 ( .A(n7340), .ZN(n7339) );
  NAND2_X1 U8495 ( .A1(n8013), .A2(n8012), .ZN(n12330) );
  AND2_X1 U8496 ( .A1(n6910), .A2(n6528), .ZN(n10526) );
  OR2_X1 U8497 ( .A1(n10431), .A2(n10758), .ZN(n7723) );
  AND2_X1 U8498 ( .A1(n10677), .A2(n10676), .ZN(n10683) );
  AND2_X1 U8499 ( .A1(n7327), .A2(n11457), .ZN(n12184) );
  NAND2_X1 U8500 ( .A1(n11456), .A2(n12181), .ZN(n7327) );
  AND2_X1 U8501 ( .A1(n12193), .A2(n6894), .ZN(n6893) );
  NAND2_X1 U8502 ( .A1(n6898), .A2(n12195), .ZN(n6894) );
  INV_X1 U8503 ( .A(n7343), .ZN(n6911) );
  AOI21_X1 U8504 ( .B1(n7321), .B2(n7323), .A(n6477), .ZN(n7318) );
  NOR2_X1 U8505 ( .A1(n10683), .A2(n7551), .ZN(n10996) );
  OR2_X1 U8506 ( .A1(n10683), .A2(n7348), .ZN(n10995) );
  CLKBUF_X1 U8507 ( .A(n12165), .Z(n12166) );
  NAND2_X1 U8508 ( .A1(n7345), .A2(n7344), .ZN(n12253) );
  NAND2_X1 U8509 ( .A1(n7995), .A2(n7994), .ZN(n12257) );
  NAND2_X1 U8510 ( .A1(n12211), .A2(n7330), .ZN(n12262) );
  NOR2_X1 U8511 ( .A1(n12260), .A2(n7331), .ZN(n7330) );
  INV_X1 U8512 ( .A(n7914), .ZN(n7331) );
  NAND2_X1 U8513 ( .A1(n12211), .A2(n7914), .ZN(n12261) );
  AND2_X1 U8514 ( .A1(n8060), .A2(n8059), .ZN(n12749) );
  INV_X1 U8515 ( .A(n12289), .ZN(n12272) );
  OR2_X1 U8516 ( .A1(n12502), .A2(n8145), .ZN(n12285) );
  OR2_X1 U8517 ( .A1(n12241), .A2(n6888), .ZN(n6882) );
  OR2_X1 U8518 ( .A1(n9399), .A2(n8068), .ZN(n7865) );
  INV_X1 U8519 ( .A(n12506), .ZN(n6748) );
  NAND2_X1 U8520 ( .A1(n8095), .A2(n8094), .ZN(n12697) );
  NOR2_X1 U8521 ( .A1(n6433), .A2(n6466), .ZN(n6773) );
  NAND2_X1 U8522 ( .A1(n7657), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6691) );
  INV_X1 U8523 ( .A(n9869), .ZN(n15142) );
  AND2_X1 U8524 ( .A1(P3_U3151), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8525 ( .A1(n6928), .A2(n9826), .ZN(n10040) );
  OR2_X1 U8526 ( .A1(n10036), .A2(n15188), .ZN(n10038) );
  NAND2_X1 U8527 ( .A1(n10038), .A2(n7548), .ZN(n10007) );
  INV_X1 U8528 ( .A(n7187), .ZN(n9991) );
  INV_X1 U8529 ( .A(n6930), .ZN(n9989) );
  INV_X1 U8530 ( .A(n7193), .ZN(n9898) );
  XNOR2_X1 U8531 ( .A(n6984), .B(n14443), .ZN(n10329) );
  INV_X1 U8532 ( .A(n7185), .ZN(n10888) );
  INV_X1 U8533 ( .A(n10891), .ZN(n15094) );
  INV_X1 U8534 ( .A(n6988), .ZN(n15121) );
  NOR2_X1 U8535 ( .A1(n11305), .A2(n11306), .ZN(n15117) );
  INV_X1 U8536 ( .A(n7179), .ZN(n15115) );
  INV_X1 U8537 ( .A(n6760), .ZN(n12522) );
  NAND2_X1 U8538 ( .A1(n7269), .A2(n7268), .ZN(n12728) );
  OR2_X1 U8539 ( .A1(n12754), .A2(n12739), .ZN(n7268) );
  AND2_X1 U8540 ( .A1(n12754), .A2(n12327), .ZN(n12740) );
  NAND2_X1 U8541 ( .A1(n12922), .A2(n12450), .ZN(n12791) );
  NAND2_X1 U8542 ( .A1(n8234), .A2(n12445), .ZN(n12805) );
  NAND2_X1 U8543 ( .A1(n12843), .A2(n12433), .ZN(n12830) );
  NAND2_X1 U8544 ( .A1(n8183), .A2(n8182), .ZN(n11403) );
  NAND2_X1 U8545 ( .A1(n7826), .A2(n7825), .ZN(n14504) );
  AND2_X1 U8546 ( .A1(n7426), .A2(n6479), .ZN(n11230) );
  NAND2_X1 U8547 ( .A1(n10949), .A2(n8179), .ZN(n11086) );
  NAND2_X1 U8548 ( .A1(n10754), .A2(n7431), .ZN(n10841) );
  AND2_X1 U8549 ( .A1(n10214), .A2(n8172), .ZN(n10424) );
  NAND2_X1 U8550 ( .A1(n10414), .A2(n10262), .ZN(n12885) );
  NAND2_X1 U8551 ( .A1(n10854), .A2(n8171), .ZN(n10216) );
  OR2_X1 U8552 ( .A1(n10239), .A2(n10238), .ZN(n12883) );
  NAND2_X1 U8553 ( .A1(n11405), .A2(n10239), .ZN(n15154) );
  INV_X1 U8554 ( .A(n11405), .ZN(n15151) );
  INV_X1 U8555 ( .A(n12330), .ZN(n12961) );
  INV_X1 U8556 ( .A(n12237), .ZN(n12973) );
  NAND2_X1 U8557 ( .A1(n7950), .A2(n7949), .ZN(n12977) );
  INV_X1 U8558 ( .A(n8190), .ZN(n12982) );
  OR3_X1 U8559 ( .A1(n12942), .A2(n12941), .A3(n12940), .ZN(n12984) );
  AND3_X1 U8560 ( .A1(n7722), .A2(n7721), .A3(n7720), .ZN(n10434) );
  OAI21_X1 U8561 ( .B1(n6730), .B2(n6729), .A(n6727), .ZN(n12294) );
  INV_X1 U8562 ( .A(n6728), .ZN(n6727) );
  NAND2_X1 U8563 ( .A1(n6471), .A2(n7615), .ZN(n12989) );
  NAND2_X1 U8564 ( .A1(n11524), .A2(n11525), .ZN(n12292) );
  XNOR2_X1 U8565 ( .A(n8201), .B(n8162), .ZN(n12998) );
  OAI21_X1 U8566 ( .B1(n8046), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8047), .ZN(
        n8066) );
  MUX2_X1 U8567 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7567), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7568) );
  NAND2_X1 U8568 ( .A1(n7571), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U8569 ( .A1(n7972), .A2(n7957), .ZN(n7958) );
  NAND2_X1 U8570 ( .A1(n7904), .A2(n7903), .ZN(n7917) );
  AND2_X1 U8571 ( .A1(n7338), .A2(n6437), .ZN(n7846) );
  NAND2_X1 U8572 ( .A1(n7085), .A2(n7086), .ZN(n7820) );
  NAND2_X1 U8573 ( .A1(n7090), .A2(n7783), .ZN(n7799) );
  NAND2_X1 U8574 ( .A1(n7781), .A2(n7780), .ZN(n7090) );
  NAND2_X1 U8575 ( .A1(n6726), .A2(n7701), .ZN(n7717) );
  NAND2_X1 U8576 ( .A1(n7700), .A2(n7699), .ZN(n6726) );
  NAND2_X1 U8577 ( .A1(n7611), .A2(n7610), .ZN(n7664) );
  NAND2_X1 U8578 ( .A1(n7648), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7662) );
  MUX2_X1 U8579 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7625), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n7627) );
  NAND2_X1 U8580 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7625) );
  NAND2_X1 U8581 ( .A1(n13122), .A2(n11971), .ZN(n13002) );
  NOR2_X1 U8582 ( .A1(n13001), .A2(n7110), .ZN(n7109) );
  INV_X1 U8583 ( .A(n11971), .ZN(n7110) );
  AND2_X1 U8584 ( .A1(n11296), .A2(n11291), .ZN(n11292) );
  NAND2_X1 U8585 ( .A1(n7133), .A2(n7130), .ZN(n14779) );
  INV_X1 U8586 ( .A(n7132), .ZN(n7130) );
  NAND2_X1 U8587 ( .A1(n8710), .A2(n8709), .ZN(n14536) );
  NOR2_X1 U8588 ( .A1(n13068), .A2(n14529), .ZN(n7120) );
  OR2_X1 U8589 ( .A1(n13068), .A2(n11927), .ZN(n7119) );
  NAND2_X1 U8590 ( .A1(n11925), .A2(n11924), .ZN(n14532) );
  AND2_X1 U8591 ( .A1(n7135), .A2(n7134), .ZN(n11993) );
  INV_X1 U8592 ( .A(n7128), .ZN(n7134) );
  NOR2_X1 U8593 ( .A1(n10828), .A2(n7115), .ZN(n7114) );
  INV_X1 U8594 ( .A(n7117), .ZN(n7115) );
  NAND2_X1 U8595 ( .A1(n7116), .A2(n6497), .ZN(n7113) );
  NAND2_X1 U8596 ( .A1(n10818), .A2(n7117), .ZN(n10871) );
  NAND2_X1 U8597 ( .A1(n11939), .A2(n13088), .ZN(n13094) );
  AND2_X1 U8598 ( .A1(n7118), .A2(n6436), .ZN(n13104) );
  INV_X1 U8599 ( .A(n13109), .ZN(n14782) );
  NAND2_X1 U8600 ( .A1(n9759), .A2(n9758), .ZN(n14777) );
  INV_X1 U8601 ( .A(n14777), .ZN(n14788) );
  NAND2_X1 U8602 ( .A1(n8682), .A2(n8681), .ZN(n13640) );
  NOR2_X1 U8603 ( .A1(n8302), .A2(n8301), .ZN(n8305) );
  NOR2_X1 U8604 ( .A1(n8361), .A2(n8300), .ZN(n8301) );
  NAND2_X1 U8605 ( .A1(n8351), .A2(n8350), .ZN(n13146) );
  NAND2_X1 U8606 ( .A1(n13151), .A2(n13545), .ZN(n6781) );
  OR2_X1 U8607 ( .A1(n13151), .A2(n13545), .ZN(n6782) );
  AOI21_X1 U8608 ( .B1(n14848), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14852), .ZN(
        n9540) );
  XNOR2_X1 U8609 ( .A(n13260), .B(n6769), .ZN(n6768) );
  INV_X1 U8610 ( .A(n13253), .ZN(n13552) );
  INV_X1 U8611 ( .A(n13325), .ZN(n13326) );
  AND2_X1 U8612 ( .A1(n7060), .A2(n6475), .ZN(n13354) );
  NAND2_X1 U8613 ( .A1(n7060), .A2(n7058), .ZN(n13564) );
  AND2_X1 U8614 ( .A1(n13356), .A2(n13355), .ZN(n13566) );
  OAI21_X1 U8615 ( .B1(n13392), .B2(n7214), .A(n7212), .ZN(n13352) );
  INV_X1 U8616 ( .A(n7216), .ZN(n13366) );
  NAND2_X1 U8617 ( .A1(n7217), .A2(n7218), .ZN(n13367) );
  NAND2_X1 U8618 ( .A1(n13392), .A2(n6464), .ZN(n7217) );
  NAND2_X1 U8619 ( .A1(n7062), .A2(n7064), .ZN(n13380) );
  NAND2_X1 U8620 ( .A1(n7069), .A2(n7065), .ZN(n7062) );
  OAI21_X1 U8621 ( .B1(n13392), .B2(n13395), .A(n7222), .ZN(n13377) );
  NAND2_X1 U8622 ( .A1(n7069), .A2(n13312), .ZN(n7068) );
  NAND2_X1 U8623 ( .A1(n7196), .A2(n7197), .ZN(n13406) );
  NAND2_X1 U8624 ( .A1(n7199), .A2(n7204), .ZN(n13421) );
  OR2_X1 U8625 ( .A1(n13436), .A2(n13279), .ZN(n7199) );
  OAI21_X1 U8626 ( .B1(n13478), .B2(n7076), .A(n7074), .ZN(n13448) );
  NOR2_X1 U8627 ( .A1(n13477), .A2(n7079), .ZN(n13463) );
  NAND2_X1 U8628 ( .A1(n7249), .A2(n7247), .ZN(n13461) );
  INV_X1 U8629 ( .A(n7250), .ZN(n7247) );
  NAND2_X1 U8630 ( .A1(n13504), .A2(n7253), .ZN(n7249) );
  OAI21_X1 U8631 ( .B1(n13504), .B2(n13271), .A(n13270), .ZN(n13474) );
  NAND2_X1 U8632 ( .A1(n8737), .A2(n8736), .ZN(n13628) );
  NAND2_X1 U8633 ( .A1(n8657), .A2(n8656), .ZN(n11512) );
  NAND2_X1 U8634 ( .A1(n7232), .A2(n11177), .ZN(n11241) );
  INV_X1 U8635 ( .A(n13533), .ZN(n13518) );
  NAND2_X1 U8636 ( .A1(n10535), .A2(n10388), .ZN(n10441) );
  OR2_X1 U8637 ( .A1(n14974), .A2(n9675), .ZN(n15078) );
  OAI21_X1 U8638 ( .B1(n15022), .B2(n13557), .A(n13563), .ZN(n13654) );
  AND2_X1 U8639 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  AND2_X1 U8640 ( .A1(n13560), .A2(n13559), .ZN(n13561) );
  NOR2_X1 U8641 ( .A1(n14944), .A2(n14976), .ZN(n14969) );
  NOR2_X1 U8642 ( .A1(n9764), .A2(P2_U3088), .ZN(n14979) );
  NOR2_X1 U8643 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6635) );
  OR2_X1 U8644 ( .A1(n9083), .A2(n13671), .ZN(n9085) );
  NAND2_X1 U8645 ( .A1(n7137), .A2(n8317), .ZN(n7136) );
  INV_X1 U8646 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9383) );
  INV_X1 U8647 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9211) );
  INV_X1 U8648 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9179) );
  INV_X1 U8649 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9164) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9147) );
  INV_X1 U8651 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9143) );
  INV_X1 U8652 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U8653 ( .A1(n10791), .A2(n10790), .ZN(n11006) );
  AOI21_X1 U8654 ( .B1(n7505), .B2(n7507), .A(n6508), .ZN(n7503) );
  NAND2_X1 U8655 ( .A1(n14542), .A2(n12031), .ZN(n14544) );
  NAND2_X1 U8656 ( .A1(n11728), .A2(n11727), .ZN(n14232) );
  OR2_X1 U8657 ( .A1(n11256), .A2(n11255), .ZN(n7541) );
  NAND2_X1 U8658 ( .A1(n10191), .A2(n10190), .ZN(n10193) );
  NAND2_X1 U8659 ( .A1(n6870), .A2(n6869), .ZN(n13708) );
  INV_X1 U8660 ( .A(n13706), .ZN(n6869) );
  NAND2_X1 U8661 ( .A1(n11006), .A2(n7522), .ZN(n11009) );
  NOR2_X1 U8662 ( .A1(n9726), .A2(n9626), .ZN(n9630) );
  NAND2_X1 U8663 ( .A1(n13766), .A2(n12081), .ZN(n13718) );
  AND2_X1 U8664 ( .A1(n11484), .A2(n6446), .ZN(n7523) );
  NAND2_X1 U8665 ( .A1(n11741), .A2(n11791), .ZN(n6808) );
  NAND2_X1 U8666 ( .A1(n6708), .A2(n7515), .ZN(n6707) );
  AND2_X1 U8667 ( .A1(n13805), .A2(n14572), .ZN(n13794) );
  AND2_X1 U8668 ( .A1(n7518), .A2(n6713), .ZN(n11122) );
  NAND2_X1 U8669 ( .A1(n13750), .A2(n12060), .ZN(n13793) );
  NAND2_X1 U8670 ( .A1(n13812), .A2(n13811), .ZN(n14555) );
  INV_X1 U8671 ( .A(n14559), .ZN(n13810) );
  INV_X1 U8672 ( .A(n11918), .ZN(n6811) );
  NAND4_X1 U8673 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n13833)
         );
  OR2_X1 U8674 ( .A1(n11797), .A2(n9597), .ZN(n9603) );
  OR2_X1 U8675 ( .A1(n11820), .A2(n9598), .ZN(n9601) );
  OR2_X1 U8676 ( .A1(n11820), .A2(n9309), .ZN(n9278) );
  NAND2_X1 U8677 ( .A1(n6443), .A2(n14707), .ZN(n14193) );
  NAND2_X1 U8678 ( .A1(n7308), .A2(n7305), .ZN(n14051) );
  NAND2_X1 U8679 ( .A1(n7295), .A2(n7298), .ZN(n14094) );
  NAND2_X1 U8680 ( .A1(n14113), .A2(n7301), .ZN(n7295) );
  NAND2_X1 U8681 ( .A1(n13942), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U8682 ( .A1(n11662), .A2(n11661), .ZN(n14153) );
  NAND2_X1 U8683 ( .A1(n7177), .A2(n7175), .ZN(n11374) );
  INV_X1 U8684 ( .A(n7005), .ZN(n11152) );
  NAND2_X1 U8685 ( .A1(n7288), .A2(n7289), .ZN(n14686) );
  NAND2_X1 U8686 ( .A1(n7291), .A2(n10272), .ZN(n10594) );
  NAND2_X1 U8687 ( .A1(n10271), .A2(n10270), .ZN(n7291) );
  NAND2_X1 U8688 ( .A1(n7170), .A2(n10075), .ZN(n11578) );
  NAND2_X1 U8689 ( .A1(n10073), .A2(n11791), .ZN(n7170) );
  NAND2_X1 U8690 ( .A1(n9942), .A2(n9941), .ZN(n13743) );
  NAND2_X1 U8691 ( .A1(n7315), .A2(n9955), .ZN(n10111) );
  INV_X1 U8692 ( .A(n9906), .ZN(n9584) );
  INV_X1 U8693 ( .A(n14101), .ZN(n14702) );
  NAND2_X1 U8694 ( .A1(n11063), .A2(n11062), .ZN(n14469) );
  NAND2_X1 U8695 ( .A1(n10963), .A2(n10962), .ZN(n11613) );
  AND2_X1 U8696 ( .A1(n14193), .A2(n14196), .ZN(n14265) );
  AND2_X1 U8697 ( .A1(n11837), .A2(n11836), .ZN(n14272) );
  NAND2_X1 U8698 ( .A1(n14208), .A2(n6754), .ZN(n14273) );
  INV_X1 U8699 ( .A(n6755), .ZN(n6754) );
  OAI21_X1 U8700 ( .B1(n14209), .B2(n14609), .A(n14207), .ZN(n6755) );
  INV_X1 U8701 ( .A(n6790), .ZN(n6789) );
  OAI21_X1 U8702 ( .B1(n14217), .B2(n14609), .A(n14216), .ZN(n6790) );
  NOR3_X1 U8703 ( .A1(n15316), .A2(n15315), .A3(n6922), .ZN(n15318) );
  AND2_X1 U8704 ( .A1(n7492), .A2(n7143), .ZN(n7142) );
  INV_X1 U8705 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7143) );
  XNOR2_X1 U8706 ( .A(n8943), .B(n8942), .ZN(n13669) );
  NAND2_X1 U8707 ( .A1(n7403), .A2(n7404), .ZN(n8943) );
  NAND2_X1 U8708 ( .A1(n7316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9231) );
  OR2_X1 U8709 ( .A1(n7535), .A2(n9123), .ZN(n6859) );
  NOR2_X1 U8710 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6858) );
  CLKBUF_X1 U8711 ( .A(n14326), .Z(n6831) );
  NAND2_X1 U8712 ( .A1(n6816), .A2(n7606), .ZN(n11714) );
  NAND2_X1 U8713 ( .A1(n9235), .A2(n9121), .ZN(n9222) );
  INV_X1 U8714 ( .A(n11869), .ZN(n11860) );
  INV_X1 U8715 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9380) );
  INV_X1 U8716 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9216) );
  INV_X1 U8717 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9197) );
  INV_X1 U8718 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U8719 ( .A(n8450), .B(n8449), .ZN(n9930) );
  AOI21_X1 U8720 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14386), .A(n15365), .ZN(
        n15357) );
  XNOR2_X1 U8721 ( .A(n14390), .B(n6872), .ZN(n15360) );
  INV_X1 U8722 ( .A(n14391), .ZN(n6872) );
  NAND2_X1 U8723 ( .A1(n15360), .A2(n15359), .ZN(n15358) );
  XNOR2_X1 U8724 ( .A(n14398), .B(n14399), .ZN(n15363) );
  XNOR2_X1 U8725 ( .A(n14403), .B(n7019), .ZN(n14461) );
  INV_X1 U8726 ( .A(n14404), .ZN(n7019) );
  NAND2_X1 U8727 ( .A1(n14466), .A2(n14465), .ZN(n14464) );
  NAND2_X1 U8728 ( .A1(n7008), .A2(n14464), .ZN(n14627) );
  OAI21_X1 U8729 ( .B1(n14466), .B2(n14465), .A(n7009), .ZN(n7008) );
  INV_X1 U8730 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U8731 ( .A1(n14627), .A2(n14628), .ZN(n14626) );
  NAND2_X1 U8732 ( .A1(n7006), .A2(n14626), .ZN(n14631) );
  OAI21_X1 U8733 ( .B1(n14627), .B2(n14628), .A(n7007), .ZN(n7006) );
  INV_X1 U8734 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7007) );
  INV_X1 U8735 ( .A(n14423), .ZN(n7016) );
  NAND2_X1 U8736 ( .A1(n7557), .A2(n10252), .ZN(n7516) );
  NAND2_X1 U8737 ( .A1(n10524), .A2(n7668), .ZN(n10626) );
  OR2_X1 U8738 ( .A1(n12505), .A2(n12504), .ZN(n6747) );
  AOI21_X1 U8739 ( .B1(n15106), .B2(P3_IR_REG_0__SCAN_IN), .A(n6923), .ZN(
        n15089) );
  OAI21_X1 U8740 ( .B1(n15085), .B2(P3_IR_REG_0__SCAN_IN), .A(n15084), .ZN(
        n15086) );
  INV_X1 U8741 ( .A(n6805), .ZN(n9877) );
  NAND2_X1 U8742 ( .A1(n6919), .A2(n6918), .ZN(n11307) );
  NAND2_X1 U8743 ( .A1(n7188), .A2(n12546), .ZN(n6931) );
  INV_X1 U8744 ( .A(n6861), .ZN(n6860) );
  OAI22_X1 U8745 ( .A1(n12948), .A2(n12933), .B1(n15199), .B2(n12892), .ZN(
        n6861) );
  INV_X1 U8746 ( .A(n6874), .ZN(n6873) );
  OAI21_X1 U8747 ( .B1(n12951), .B2(n12933), .A(n6875), .ZN(n6874) );
  AND2_X1 U8748 ( .A1(n8258), .A2(n7552), .ZN(n8259) );
  INV_X1 U8749 ( .A(n6864), .ZN(n6863) );
  OAI22_X1 U8750 ( .A1(n12948), .A2(n12981), .B1(n15185), .B2(n12947), .ZN(
        n6864) );
  NAND2_X1 U8751 ( .A1(n6759), .A2(n6757), .ZN(P3_U3454) );
  AOI21_X1 U8752 ( .B1(n8199), .B2(n8256), .A(n6758), .ZN(n6757) );
  OR2_X1 U8753 ( .A1(n12949), .A2(n15187), .ZN(n6759) );
  NOR2_X1 U8754 ( .A1(n15185), .A2(n12950), .ZN(n6758) );
  OAI21_X1 U8755 ( .B1(n12995), .B2(n14451), .A(n6699), .ZN(P3_U3266) );
  AOI21_X1 U8756 ( .B1(n7619), .B2(P3_STATE_REG_SCAN_IN), .A(n6700), .ZN(n6699) );
  NOR2_X1 U8757 ( .A1(n12997), .A2(n12996), .ZN(n6700) );
  NAND2_X1 U8758 ( .A1(n6668), .A2(n6854), .ZN(n6853) );
  AND2_X1 U8759 ( .A1(n13245), .A2(n6779), .ZN(n13248) );
  NAND2_X1 U8760 ( .A1(n6602), .A2(n6810), .ZN(n6809) );
  INV_X1 U8761 ( .A(n11917), .ZN(n6810) );
  AOI211_X1 U8762 ( .C1(n14200), .C2(n14711), .A(n13995), .B(n13994), .ZN(
        n13996) );
  AND2_X1 U8763 ( .A1(n7167), .A2(n6573), .ZN(n14204) );
  OR2_X1 U8764 ( .A1(n14772), .A2(n6960), .ZN(n6959) );
  INV_X1 U8765 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6960) );
  AND2_X1 U8766 ( .A1(n6835), .A2(n6819), .ZN(n6818) );
  NAND2_X1 U8767 ( .A1(n6820), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U8768 ( .A1(n14026), .A2(n14263), .ZN(n6835) );
  NAND2_X1 U8769 ( .A1(n14763), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7168) );
  AOI21_X1 U8770 ( .B1(n14026), .B2(n6824), .A(n6823), .ZN(n6822) );
  NOR2_X1 U8771 ( .A1(n14764), .A2(n14275), .ZN(n6823) );
  INV_X1 U8772 ( .A(n6834), .ZN(n14634) );
  INV_X1 U8773 ( .A(n14640), .ZN(n14639) );
  INV_X1 U8774 ( .A(n14645), .ZN(n14644) );
  NAND2_X1 U8775 ( .A1(n14486), .A2(n6766), .ZN(n14433) );
  OR2_X1 U8776 ( .A1(n14485), .A2(n14484), .ZN(n6766) );
  XNOR2_X1 U8777 ( .A(n14490), .B(n14489), .ZN(n7020) );
  NAND2_X2 U8778 ( .A1(n8951), .A2(n9760), .ZN(n10303) );
  OR2_X1 U8779 ( .A1(n14795), .A2(n13133), .ZN(n6428) );
  AND2_X1 U8780 ( .A1(n7406), .A2(n6598), .ZN(n6429) );
  INV_X2 U8781 ( .A(n9796), .ZN(n12626) );
  AND2_X1 U8782 ( .A1(n7517), .A2(n10190), .ZN(n6430) );
  INV_X1 U8783 ( .A(n11870), .ZN(n9281) );
  INV_X1 U8784 ( .A(n11402), .ZN(n7423) );
  AND2_X1 U8785 ( .A1(n7151), .A2(n7156), .ZN(n6431) );
  AND2_X1 U8786 ( .A1(n7339), .A2(n12219), .ZN(n6432) );
  XNOR2_X1 U8787 ( .A(n11587), .B(n10787), .ZN(n10270) );
  INV_X1 U8788 ( .A(n10270), .ZN(n11883) );
  NAND2_X1 U8789 ( .A1(n14038), .A2(n13958), .ZN(n7158) );
  AND2_X1 U8790 ( .A1(n7634), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8791 ( .A1(n8754), .A2(n8753), .ZN(n13623) );
  NOR2_X1 U8792 ( .A1(n10458), .A2(n10445), .ZN(n6434) );
  INV_X1 U8793 ( .A(n7059), .ZN(n7058) );
  NAND2_X1 U8794 ( .A1(n13353), .A2(n6475), .ZN(n7059) );
  AND2_X1 U8795 ( .A1(n9826), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6435) );
  AND2_X1 U8796 ( .A1(n7119), .A2(n6514), .ZN(n6436) );
  AND2_X1 U8797 ( .A1(n7565), .A2(n7801), .ZN(n6437) );
  XNOR2_X1 U8798 ( .A(n13568), .B(n13286), .ZN(n13321) );
  INV_X1 U8799 ( .A(n13321), .ZN(n13353) );
  INV_X1 U8800 ( .A(n12826), .ZN(n7434) );
  AND2_X1 U8801 ( .A1(n9276), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6438) );
  AND4_X1 U8802 ( .A1(n7416), .A2(n12713), .A3(n12727), .A4(n12322), .ZN(n6439) );
  AND2_X1 U8803 ( .A1(n7852), .A2(n12511), .ZN(n6441) );
  AND2_X1 U8804 ( .A1(n6436), .A2(n13103), .ZN(n6442) );
  INV_X1 U8805 ( .A(n14795), .ZN(n11427) );
  NAND2_X1 U8806 ( .A1(n8633), .A2(n8632), .ZN(n14795) );
  AOI21_X1 U8807 ( .B1(n7519), .B2(n7520), .A(n6541), .ZN(n7518) );
  XOR2_X1 U8808 ( .A(n13922), .B(n13929), .Z(n6443) );
  INV_X1 U8809 ( .A(n7077), .ZN(n7076) );
  AOI21_X1 U8810 ( .B1(n7078), .B2(n13479), .A(n13306), .ZN(n7077) );
  INV_X1 U8811 ( .A(n12498), .ZN(n12945) );
  NAND2_X1 U8812 ( .A1(n7084), .A2(n12295), .ZN(n12498) );
  AND2_X1 U8813 ( .A1(n13072), .A2(n6510), .ZN(n6444) );
  OR2_X1 U8814 ( .A1(n7067), .A2(n13315), .ZN(n7064) );
  AND2_X1 U8815 ( .A1(n6539), .A2(n12498), .ZN(n6445) );
  INV_X1 U8816 ( .A(n7436), .ZN(n7435) );
  NAND2_X1 U8817 ( .A1(n12817), .A2(n7437), .ZN(n7436) );
  OR2_X1 U8818 ( .A1(n11477), .A2(n11476), .ZN(n6446) );
  AND2_X1 U8819 ( .A1(n8459), .A2(n8458), .ZN(n6447) );
  AND2_X1 U8820 ( .A1(n8505), .A2(n8504), .ZN(n6448) );
  INV_X1 U8821 ( .A(n13558), .ZN(n7028) );
  INV_X1 U8822 ( .A(n14492), .ZN(n12302) );
  AND2_X1 U8823 ( .A1(n7027), .A2(n8291), .ZN(n6449) );
  OR2_X1 U8824 ( .A1(n13410), .A2(n7203), .ZN(n6450) );
  NAND2_X1 U8825 ( .A1(n11529), .A2(n6698), .ZN(n8057) );
  NAND2_X1 U8826 ( .A1(n8747), .A2(n8746), .ZN(n6451) );
  INV_X1 U8827 ( .A(n12690), .ZN(n6738) );
  AND2_X1 U8828 ( .A1(n11160), .A2(n11159), .ZN(n6452) );
  OR2_X1 U8829 ( .A1(n6451), .A2(n6570), .ZN(n6453) );
  INV_X1 U8830 ( .A(n8199), .ZN(n12951) );
  NAND2_X1 U8831 ( .A1(n8086), .A2(n8085), .ZN(n8199) );
  INV_X1 U8832 ( .A(n15125), .ZN(n6983) );
  AND2_X1 U8833 ( .A1(n12675), .A2(n12540), .ZN(n6454) );
  INV_X1 U8834 ( .A(n7409), .ZN(n7408) );
  AOI21_X1 U8835 ( .B1(n8975), .B2(n8938), .A(n7410), .ZN(n7409) );
  OR2_X1 U8836 ( .A1(n8868), .A2(n7376), .ZN(n6455) );
  AND2_X1 U8837 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8029), .ZN(n6456) );
  INV_X2 U8839 ( .A(n9944), .ZN(n11707) );
  INV_X2 U8840 ( .A(n11136), .ZN(n13529) );
  OR2_X1 U8841 ( .A1(n7571), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6458) );
  AND2_X1 U8842 ( .A1(n12497), .A2(n6746), .ZN(n6459) );
  OR2_X1 U8843 ( .A1(n8312), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8844 ( .A1(n13768), .A2(n13767), .ZN(n13766) );
  INV_X1 U8845 ( .A(n7634), .ZN(n7827) );
  INV_X2 U8846 ( .A(n7827), .ZN(n8090) );
  NOR2_X1 U8847 ( .A1(n14073), .A2(n13988), .ZN(n6461) );
  AND2_X1 U8848 ( .A1(n13141), .A2(n15001), .ZN(n6462) );
  NAND2_X1 U8849 ( .A1(n12965), .A2(n8007), .ZN(n6463) );
  INV_X1 U8850 ( .A(n14018), .ZN(n7155) );
  AND2_X1 U8851 ( .A1(n7221), .A2(n7222), .ZN(n6464) );
  OR2_X1 U8852 ( .A1(n7457), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6465) );
  AND2_X1 U8853 ( .A1(n7657), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6466) );
  INV_X1 U8854 ( .A(n14038), .ZN(n14280) );
  AND2_X1 U8855 ( .A1(n7264), .A2(n7265), .ZN(n6467) );
  NAND2_X1 U8856 ( .A1(n14044), .A2(n6997), .ZN(n6468) );
  INV_X1 U8857 ( .A(n8127), .ZN(n6848) );
  OR2_X1 U8858 ( .A1(n8577), .A2(n8576), .ZN(n6469) );
  NAND2_X1 U8859 ( .A1(n6719), .A2(n7765), .ZN(n7781) );
  OR2_X1 U8860 ( .A1(n13921), .A2(n14019), .ZN(n6470) );
  AND4_X1 U8861 ( .A1(n6683), .A2(n6912), .A3(n7561), .A4(n7411), .ZN(n6471)
         );
  OR2_X1 U8862 ( .A1(n11818), .A2(n9910), .ZN(n6472) );
  NAND2_X1 U8863 ( .A1(n12101), .A2(n12100), .ZN(n13759) );
  NAND2_X1 U8864 ( .A1(n8238), .A2(n12714), .ZN(n6473) );
  NAND2_X1 U8865 ( .A1(n14153), .A2(n13943), .ZN(n6474) );
  OR2_X1 U8866 ( .A1(n13373), .A2(n13318), .ZN(n6475) );
  INV_X1 U8867 ( .A(n8578), .ZN(n8579) );
  XNOR2_X1 U8868 ( .A(n8581), .B(SI_10_), .ZN(n8578) );
  AND2_X1 U8869 ( .A1(n8101), .A2(n8100), .ZN(n6476) );
  AND2_X1 U8870 ( .A1(n7896), .A2(n12839), .ZN(n6477) );
  XNOR2_X1 U8871 ( .A(n14205), .B(n13960), .ZN(n14009) );
  INV_X1 U8872 ( .A(n14009), .ZN(n6951) );
  XNOR2_X1 U8873 ( .A(n11565), .B(n10253), .ZN(n11880) );
  INV_X1 U8874 ( .A(n11880), .ZN(n7314) );
  XNOR2_X1 U8875 ( .A(n15144), .B(n8167), .ZN(n12339) );
  NAND2_X1 U8876 ( .A1(n8946), .A2(n8945), .ZN(n9033) );
  INV_X1 U8877 ( .A(n9033), .ZN(n6769) );
  INV_X1 U8878 ( .A(n12310), .ZN(n7276) );
  NAND2_X1 U8879 ( .A1(n8791), .A2(n8790), .ZN(n13449) );
  INV_X1 U8880 ( .A(n13449), .ZN(n6770) );
  NAND2_X1 U8881 ( .A1(n9927), .A2(n9928), .ZN(n14705) );
  INV_X1 U8882 ( .A(n13095), .ZN(n7125) );
  AND4_X1 U8883 ( .A1(n9160), .A2(n9238), .A3(n9239), .A4(n9117), .ZN(n6478)
         );
  OR2_X1 U8884 ( .A1(n11462), .A2(n11202), .ZN(n6479) );
  OR2_X1 U8885 ( .A1(n14268), .A2(n14300), .ZN(n6480) );
  NAND2_X1 U8886 ( .A1(n8018), .A2(n12219), .ZN(n12149) );
  OR2_X1 U8887 ( .A1(n14276), .A2(n13999), .ZN(n6481) );
  OR2_X1 U8888 ( .A1(n12948), .A2(n12715), .ZN(n6482) );
  INV_X1 U8889 ( .A(n11795), .ZN(n7496) );
  OR2_X1 U8890 ( .A1(n9090), .A2(n13159), .ZN(n6483) );
  INV_X1 U8891 ( .A(n11589), .ZN(n7501) );
  AND2_X1 U8892 ( .A1(n15038), .A2(n13137), .ZN(n6484) );
  INV_X1 U8893 ( .A(n12518), .ZN(n10437) );
  NAND2_X1 U8894 ( .A1(n7865), .A2(n7864), .ZN(n12879) );
  INV_X1 U8895 ( .A(n12879), .ZN(n7420) );
  NOR2_X1 U8896 ( .A1(n10722), .A2(n10458), .ZN(n6485) );
  AND2_X1 U8897 ( .A1(n8488), .A2(n8487), .ZN(n6486) );
  INV_X1 U8898 ( .A(n10828), .ZN(n7116) );
  MUX2_X1 U8899 ( .A(n13985), .B(n13986), .S(n11844), .Z(n11717) );
  INV_X1 U8900 ( .A(n11717), .ZN(n7494) );
  AND2_X1 U8901 ( .A1(n13618), .A2(n13274), .ZN(n6487) );
  OR2_X1 U8902 ( .A1(n7038), .A2(n13311), .ZN(n6488) );
  AND4_X1 U8903 ( .A1(n7578), .A2(n7577), .A3(n7576), .A4(n8123), .ZN(n6489)
         );
  OR2_X1 U8904 ( .A1(n9090), .A2(n14809), .ZN(n6490) );
  INV_X1 U8905 ( .A(n13598), .ZN(n7038) );
  NOR2_X1 U8906 ( .A1(n9944), .A2(n9285), .ZN(n6491) );
  OR2_X1 U8907 ( .A1(n9894), .A2(n9876), .ZN(n6492) );
  NOR2_X1 U8908 ( .A1(n12642), .A2(n12643), .ZN(n6493) );
  AND2_X1 U8909 ( .A1(n7294), .A2(n7296), .ZN(n6494) );
  OAI21_X1 U8910 ( .B1(n11844), .B2(n6845), .A(n6844), .ZN(n11576) );
  INV_X1 U8911 ( .A(n11576), .ZN(n11577) );
  AND2_X1 U8912 ( .A1(n10890), .A2(n14449), .ZN(n6495) );
  AND2_X1 U8913 ( .A1(n10423), .A2(n8172), .ZN(n6496) );
  AND2_X1 U8914 ( .A1(n10826), .A2(n10820), .ZN(n6497) );
  AND2_X1 U8915 ( .A1(n9123), .A2(n7529), .ZN(n6498) );
  INV_X1 U8916 ( .A(n8405), .ZN(n6855) );
  AND2_X1 U8917 ( .A1(n12767), .A2(n6463), .ZN(n6499) );
  INV_X1 U8918 ( .A(n12767), .ZN(n12762) );
  NAND2_X1 U8919 ( .A1(n12329), .A2(n8194), .ZN(n12767) );
  OR2_X1 U8920 ( .A1(n11990), .A2(n10702), .ZN(n6500) );
  OR2_X1 U8921 ( .A1(n10910), .A2(n10887), .ZN(n6501) );
  INV_X1 U8922 ( .A(n13944), .ZN(n14126) );
  INV_X1 U8923 ( .A(n7066), .ZN(n7065) );
  NAND2_X1 U8924 ( .A1(n7070), .A2(n13312), .ZN(n7066) );
  AND2_X1 U8925 ( .A1(n12083), .A2(n12081), .ZN(n6502) );
  OR2_X1 U8926 ( .A1(n14268), .A2(n14259), .ZN(n6503) );
  OR2_X1 U8927 ( .A1(n8551), .A2(n8552), .ZN(n6504) );
  AND2_X1 U8928 ( .A1(n12703), .A2(n7417), .ZN(n6505) );
  OR2_X1 U8929 ( .A1(n11588), .A2(n7501), .ZN(n6506) );
  AND2_X1 U8930 ( .A1(n9031), .A2(n9032), .ZN(n6507) );
  AND2_X1 U8931 ( .A1(n12121), .A2(n12120), .ZN(n6508) );
  AND2_X1 U8932 ( .A1(n12066), .A2(n12065), .ZN(n6509) );
  NAND2_X1 U8933 ( .A1(n11954), .A2(n13010), .ZN(n6510) );
  INV_X1 U8934 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7559) );
  INV_X1 U8935 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8317) );
  INV_X1 U8936 ( .A(n6689), .ZN(n10650) );
  OR2_X1 U8937 ( .A1(n6770), .A2(n13307), .ZN(n6511) );
  NOR2_X1 U8938 ( .A1(n11912), .A2(n11911), .ZN(n6512) );
  NOR2_X1 U8939 ( .A1(n14737), .A2(n13830), .ZN(n6513) );
  OR2_X1 U8940 ( .A1(n8238), .A2(n12714), .ZN(n12471) );
  OR2_X1 U8941 ( .A1(n11931), .A2(n11930), .ZN(n6514) );
  NOR2_X1 U8942 ( .A1(n14469), .A2(n13825), .ZN(n6515) );
  NOR2_X1 U8943 ( .A1(n13598), .A2(n13311), .ZN(n6516) );
  NOR2_X1 U8944 ( .A1(n13986), .A2(n13985), .ZN(n6517) );
  NOR2_X1 U8945 ( .A1(n14499), .A2(n12874), .ZN(n6518) );
  NAND2_X1 U8946 ( .A1(n12482), .A2(n8239), .ZN(n12703) );
  INV_X1 U8947 ( .A(n12703), .ZN(n7416) );
  AND4_X1 U8948 ( .A1(n7601), .A2(n7600), .A3(n7599), .A4(n7598), .ZN(n6519)
         );
  AND2_X1 U8949 ( .A1(n12390), .A2(n12515), .ZN(n6520) );
  AND2_X1 U8950 ( .A1(n9828), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7184) );
  NAND2_X1 U8951 ( .A1(n11097), .A2(n11096), .ZN(n6521) );
  AND3_X1 U8952 ( .A1(n9601), .A2(n9600), .A3(n9602), .ZN(n6522) );
  AND2_X1 U8953 ( .A1(n8510), .A2(SI_7_), .ZN(n6523) );
  AND2_X1 U8954 ( .A1(n8581), .A2(SI_10_), .ZN(n6524) );
  OR2_X1 U8955 ( .A1(n8507), .A2(n6448), .ZN(n6525) );
  NAND2_X1 U8956 ( .A1(n11609), .A2(n10977), .ZN(n6526) );
  NAND2_X1 U8957 ( .A1(n7909), .A2(n7566), .ZN(n6527) );
  NAND2_X1 U8958 ( .A1(n7362), .A2(n8653), .ZN(n8697) );
  NAND2_X1 U8959 ( .A1(n7656), .A2(n10802), .ZN(n6528) );
  AND2_X1 U8960 ( .A1(n6848), .A2(n11019), .ZN(n6529) );
  AND2_X1 U8961 ( .A1(n11243), .A2(n11242), .ZN(n6530) );
  NOR2_X1 U8962 ( .A1(n14060), .A2(n6461), .ZN(n6531) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9176) );
  INV_X1 U8964 ( .A(n7281), .ZN(n7280) );
  NAND2_X1 U8965 ( .A1(n12826), .A2(n12433), .ZN(n7281) );
  NAND2_X1 U8966 ( .A1(n8622), .A2(n8623), .ZN(n6532) );
  NAND2_X1 U8967 ( .A1(n6897), .A2(n12220), .ZN(n12192) );
  AND2_X1 U8968 ( .A1(n12437), .A2(n12440), .ZN(n12826) );
  AND2_X1 U8969 ( .A1(n7432), .A2(n6678), .ZN(n6533) );
  AND2_X1 U8970 ( .A1(n9176), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6534) );
  OR2_X1 U8971 ( .A1(n7494), .A2(n11716), .ZN(n6535) );
  INV_X1 U8972 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9181) );
  NOR2_X1 U8973 ( .A1(n13574), .A2(n13318), .ZN(n6536) );
  INV_X1 U8974 ( .A(n7431), .ZN(n7430) );
  INV_X1 U8975 ( .A(n13323), .ZN(n13341) );
  NAND2_X1 U8976 ( .A1(n13324), .A2(n9051), .ZN(n13323) );
  NOR2_X1 U8977 ( .A1(n11324), .A2(n10892), .ZN(n6537) );
  AND2_X1 U8978 ( .A1(n13568), .A2(n13286), .ZN(n6538) );
  NAND2_X1 U8979 ( .A1(n7083), .A2(n7081), .ZN(n6539) );
  AND2_X1 U8980 ( .A1(n14795), .A2(n13133), .ZN(n6540) );
  AND2_X1 U8981 ( .A1(n11115), .A2(n11114), .ZN(n6541) );
  INV_X1 U8982 ( .A(n13990), .ZN(n6958) );
  NAND2_X1 U8983 ( .A1(n7354), .A2(n7352), .ZN(n11908) );
  INV_X1 U8984 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10016) );
  AND2_X1 U8985 ( .A1(n8927), .A2(n7446), .ZN(n6542) );
  AND2_X1 U8986 ( .A1(n14205), .A2(n14019), .ZN(n6543) );
  INV_X1 U8987 ( .A(n12323), .ZN(n6787) );
  AND2_X1 U8988 ( .A1(n11953), .A2(n7124), .ZN(n6544) );
  OR2_X1 U8989 ( .A1(n8140), .A2(n10050), .ZN(n6545) );
  AND2_X1 U8990 ( .A1(n7381), .A2(n7380), .ZN(n6546) );
  AND2_X1 U8991 ( .A1(n11953), .A2(n11954), .ZN(n6547) );
  OR2_X1 U8992 ( .A1(n6447), .A2(n8461), .ZN(n6548) );
  AND2_X1 U8993 ( .A1(n7197), .A2(n6450), .ZN(n6549) );
  OR2_X1 U8994 ( .A1(n8693), .A2(n8695), .ZN(n6550) );
  OR2_X1 U8995 ( .A1(n13955), .A2(n6461), .ZN(n7309) );
  INV_X1 U8996 ( .A(n7309), .ZN(n7305) );
  AND2_X1 U8997 ( .A1(n12128), .A2(n12127), .ZN(n6551) );
  INV_X1 U8998 ( .A(n13991), .ZN(n6957) );
  INV_X1 U8999 ( .A(n13973), .ZN(n14598) );
  AND2_X1 U9000 ( .A1(n11377), .A2(n11376), .ZN(n13973) );
  AND2_X1 U9001 ( .A1(n7179), .A2(n7178), .ZN(n6552) );
  AND2_X1 U9002 ( .A1(n9830), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6553) );
  AND2_X1 U9003 ( .A1(n12478), .A2(n12701), .ZN(n12713) );
  AND2_X1 U9004 ( .A1(n10503), .A2(n10252), .ZN(n6554) );
  AND2_X1 U9005 ( .A1(n8992), .A2(n6507), .ZN(n6555) );
  INV_X1 U9006 ( .A(n7049), .ZN(n7048) );
  OAI21_X1 U9007 ( .B1(n10743), .B2(n7050), .A(n10931), .ZN(n7049) );
  AND2_X1 U9008 ( .A1(n6431), .A2(n6470), .ZN(n6556) );
  OR2_X1 U9009 ( .A1(n7496), .A2(n11794), .ZN(n6557) );
  NOR2_X1 U9010 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n6558) );
  OR2_X1 U9011 ( .A1(n7459), .A2(n8694), .ZN(n6559) );
  OR2_X1 U9012 ( .A1(n11600), .A2(n11598), .ZN(n6560) );
  INV_X1 U9013 ( .A(n7299), .ZN(n7298) );
  NAND2_X1 U9014 ( .A1(n14095), .A2(n7300), .ZN(n7299) );
  OR2_X1 U9015 ( .A1(n11610), .A2(n11612), .ZN(n6561) );
  AND2_X1 U9016 ( .A1(n11944), .A2(n11943), .ZN(n6562) );
  AND2_X1 U9017 ( .A1(n6677), .A2(n6463), .ZN(n6563) );
  OR2_X1 U9018 ( .A1(n7449), .A2(n7448), .ZN(n6564) );
  INV_X1 U9019 ( .A(n13955), .ZN(n14052) );
  NAND2_X1 U9020 ( .A1(n12951), .A2(n12726), .ZN(n7417) );
  NOR2_X1 U9021 ( .A1(n13554), .A2(n7240), .ZN(n6565) );
  NAND2_X1 U9022 ( .A1(n13568), .A2(n13322), .ZN(n6566) );
  AND2_X1 U9023 ( .A1(n7161), .A2(n6474), .ZN(n6567) );
  INV_X1 U9024 ( .A(n10503), .ZN(n7515) );
  INV_X1 U9025 ( .A(n7201), .ZN(n7200) );
  NAND2_X1 U9026 ( .A1(n13280), .A2(n7202), .ZN(n7201) );
  INV_X1 U9027 ( .A(n13315), .ZN(n7070) );
  AND2_X1 U9028 ( .A1(n13587), .A2(n13314), .ZN(n13315) );
  AND2_X1 U9029 ( .A1(n13640), .A2(n13509), .ZN(n6568) );
  INV_X1 U9030 ( .A(n7215), .ZN(n7214) );
  AND2_X1 U9031 ( .A1(n7218), .A2(n7216), .ZN(n7215) );
  INV_X1 U9032 ( .A(n7275), .ZN(n7274) );
  NAND2_X1 U9033 ( .A1(n7276), .A2(n8228), .ZN(n7275) );
  INV_X1 U9034 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7141) );
  NOR2_X1 U9035 ( .A1(n7798), .A2(n7089), .ZN(n7088) );
  NOR2_X1 U9036 ( .A1(n11010), .A2(n7521), .ZN(n7520) );
  AND3_X1 U9037 ( .A1(n9110), .A2(n6853), .A3(n9109), .ZN(P2_U3328) );
  XNOR2_X1 U9038 ( .A(n6676), .B(n8317), .ZN(n10369) );
  INV_X1 U9039 ( .A(n14073), .ZN(n6991) );
  INV_X1 U9040 ( .A(n13281), .ZN(n7203) );
  NOR2_X1 U9041 ( .A1(n8679), .A2(n7138), .ZN(n8731) );
  AND2_X1 U9042 ( .A1(n8745), .A2(n8744), .ZN(n6570) );
  AND2_X1 U9043 ( .A1(n8284), .A2(n8417), .ZN(n8559) );
  XNOR2_X1 U9044 ( .A(n12516), .B(n12384), .ZN(n12378) );
  INV_X1 U9045 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13671) );
  AND2_X1 U9046 ( .A1(n6437), .A2(n7334), .ZN(n7881) );
  INV_X1 U9047 ( .A(n14443), .ZN(n10910) );
  NAND2_X1 U9048 ( .A1(n6889), .A2(n6892), .ZN(n11464) );
  NAND2_X1 U9049 ( .A1(n6882), .A2(n6886), .ZN(n12279) );
  OR2_X1 U9050 ( .A1(n12182), .A2(n12246), .ZN(n6571) );
  OR2_X1 U9051 ( .A1(n14280), .A2(n14300), .ZN(n6572) );
  NAND2_X1 U9052 ( .A1(n7953), .A2(n7952), .ZN(n12231) );
  NAND2_X1 U9053 ( .A1(n14019), .A2(n14572), .ZN(n6573) );
  AND2_X1 U9054 ( .A1(n8042), .A2(n8041), .ZN(n12152) );
  AND2_X1 U9055 ( .A1(n8828), .A2(n7371), .ZN(n6574) );
  AND2_X1 U9056 ( .A1(n8822), .A2(n8821), .ZN(n6575) );
  AND2_X1 U9057 ( .A1(n6969), .A2(n6970), .ZN(n6576) );
  INV_X1 U9058 ( .A(n6771), .ZN(n13464) );
  INV_X1 U9059 ( .A(n7177), .ZN(n11344) );
  NAND2_X1 U9060 ( .A1(n6452), .A2(n11161), .ZN(n7177) );
  OR2_X1 U9061 ( .A1(n14280), .A2(n14259), .ZN(n6577) );
  AND2_X1 U9062 ( .A1(n12843), .A2(n7280), .ZN(n6578) );
  AND2_X1 U9063 ( .A1(n7118), .A2(n7119), .ZN(n6579) );
  OR2_X1 U9064 ( .A1(n7452), .A2(n6575), .ZN(n6580) );
  AND2_X1 U9065 ( .A1(n9211), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6581) );
  AND2_X1 U9066 ( .A1(n7086), .A2(n7819), .ZN(n6582) );
  OR2_X1 U9067 ( .A1(n13299), .A2(n13300), .ZN(n6583) );
  AND2_X1 U9068 ( .A1(n14001), .A2(n14000), .ZN(n6584) );
  NOR2_X1 U9069 ( .A1(n12824), .A2(n7438), .ZN(n6585) );
  OR2_X1 U9070 ( .A1(n7386), .A2(n7387), .ZN(n6586) );
  AND2_X1 U9071 ( .A1(n6571), .A2(n12181), .ZN(n6587) );
  AND2_X1 U9072 ( .A1(n7524), .A2(n6446), .ZN(n6588) );
  INV_X1 U9073 ( .A(n14772), .ZN(n6820) );
  INV_X1 U9074 ( .A(n14300), .ZN(n6824) );
  AND2_X1 U9075 ( .A1(n7277), .A2(n7274), .ZN(n6589) );
  NAND2_X1 U9076 ( .A1(n10818), .A2(n7114), .ZN(n7112) );
  NAND2_X1 U9077 ( .A1(n10785), .A2(n6828), .ZN(n10791) );
  OR2_X1 U9078 ( .A1(n11192), .A2(n15054), .ZN(n6590) );
  NAND2_X1 U9079 ( .A1(n6857), .A2(n6859), .ZN(n11532) );
  NAND2_X1 U9080 ( .A1(n10317), .A2(n8174), .ZN(n10756) );
  NAND2_X1 U9081 ( .A1(n14753), .A2(n10572), .ZN(n10976) );
  AND2_X1 U9082 ( .A1(n12536), .A2(n6867), .ZN(n6591) );
  AND2_X1 U9083 ( .A1(n11006), .A2(n7520), .ZN(n6592) );
  AND2_X1 U9084 ( .A1(n7178), .A2(n12532), .ZN(n6593) );
  OR2_X1 U9085 ( .A1(n7402), .A2(n7399), .ZN(n7398) );
  OR2_X1 U9086 ( .A1(n9220), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6594) );
  AND2_X1 U9087 ( .A1(n7112), .A2(n7113), .ZN(n6595) );
  AND2_X1 U9088 ( .A1(n8939), .A2(n12996), .ZN(n6596) );
  AND2_X1 U9089 ( .A1(n6455), .A2(n8887), .ZN(n6597) );
  INV_X1 U9090 ( .A(n13837), .ZN(n9732) );
  XOR2_X1 U9091 ( .A(n8940), .B(SI_30_), .Z(n6598) );
  NAND2_X1 U9092 ( .A1(n7605), .A2(n7604), .ZN(n8139) );
  INV_X1 U9093 ( .A(n12638), .ZN(n6806) );
  INV_X1 U9094 ( .A(n13508), .ZN(n13116) );
  AND2_X1 U9095 ( .A1(n6981), .A2(n6980), .ZN(n6599) );
  OR2_X1 U9096 ( .A1(n8977), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6600) );
  AND2_X1 U9097 ( .A1(n6806), .A2(n12666), .ZN(n6601) );
  INV_X1 U9098 ( .A(n12687), .ZN(n12499) );
  XNOR2_X1 U9099 ( .A(n8324), .B(n8323), .ZN(n9094) );
  OR3_X1 U9100 ( .A1(n11916), .A2(n14165), .A3(n11915), .ZN(n6602) );
  INV_X1 U9101 ( .A(n15020), .ZN(n7033) );
  NAND2_X1 U9102 ( .A1(n10563), .A2(n10562), .ZN(n14756) );
  INV_X1 U9103 ( .A(n14756), .ZN(n6993) );
  INV_X1 U9104 ( .A(n6831), .ZN(n7533) );
  AND2_X1 U9105 ( .A1(n10524), .A2(n7341), .ZN(n6603) );
  AND2_X1 U9106 ( .A1(n8940), .A2(SI_30_), .ZN(n6604) );
  OR2_X1 U9107 ( .A1(n7103), .A2(n7100), .ZN(n6605) );
  AND2_X1 U9108 ( .A1(n11755), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6606) );
  INV_X1 U9109 ( .A(SI_22_), .ZN(n7371) );
  INV_X1 U9110 ( .A(SI_24_), .ZN(n7376) );
  NAND2_X2 U9111 ( .A1(n11870), .A2(n7534), .ZN(n14718) );
  INV_X1 U9112 ( .A(n14718), .ZN(n14707) );
  INV_X1 U9113 ( .A(n11525), .ZN(n6729) );
  NOR2_X1 U9114 ( .A1(n10009), .A2(n10010), .ZN(n6607) );
  OR2_X1 U9115 ( .A1(n14318), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6608) );
  NAND4_X1 U9116 ( .A1(n9240), .A2(n9229), .A3(n7142), .A4(n9230), .ZN(n14305)
         );
  NAND2_X2 U9117 ( .A1(n9280), .A2(n11536), .ZN(n14751) );
  NAND2_X1 U9118 ( .A1(n11064), .A2(n11889), .ZN(n11160) );
  NAND2_X1 U9119 ( .A1(n10093), .A2(n10092), .ZN(n10279) );
  NAND2_X1 U9120 ( .A1(n14676), .A2(n7144), .ZN(n14753) );
  NAND2_X2 U9121 ( .A1(n6522), .A2(n9603), .ZN(n13836) );
  NAND2_X4 U9122 ( .A1(n9275), .A2(n9276), .ZN(n11818) );
  XNOR2_X2 U9123 ( .A(n9273), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9276) );
  XNOR2_X2 U9124 ( .A(n9271), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9275) );
  OR2_X2 U9125 ( .A1(n14050), .A2(n14052), .ZN(n14048) );
  NAND2_X1 U9126 ( .A1(n6622), .A2(n14751), .ZN(n6620) );
  NAND2_X1 U9127 ( .A1(n14041), .A2(n13959), .ZN(n6623) );
  AND3_X2 U9128 ( .A1(n6478), .A2(n6625), .A3(n6624), .ZN(n9229) );
  AND2_X2 U9129 ( .A1(n7514), .A2(n7513), .ZN(n9240) );
  AND2_X1 U9130 ( .A1(n9116), .A2(n9115), .ZN(n7513) );
  INV_X1 U9131 ( .A(n6868), .ZN(n7514) );
  NAND2_X1 U9132 ( .A1(n11531), .A2(n6438), .ZN(n9277) );
  NAND2_X4 U9133 ( .A1(n11531), .A2(n9276), .ZN(n6802) );
  NAND2_X1 U9134 ( .A1(n6626), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U9135 ( .A1(n6626), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U9136 ( .A1(n6627), .A2(n10124), .ZN(n10093) );
  XNOR2_X1 U9137 ( .A(n6627), .B(n10124), .ZN(n10129) );
  NAND2_X1 U9138 ( .A1(n6469), .A2(n6632), .ZN(n8601) );
  NAND3_X1 U9139 ( .A1(n8531), .A2(n6564), .A3(n8530), .ZN(n6634) );
  NAND2_X1 U9140 ( .A1(n8320), .A2(n6635), .ZN(n13670) );
  NAND2_X1 U9141 ( .A1(n6640), .A2(n7461), .ZN(n8764) );
  AOI21_X1 U9142 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n8786) );
  NAND2_X1 U9143 ( .A1(n6644), .A2(n6642), .ZN(n8383) );
  INV_X1 U9144 ( .A(n6649), .ZN(n6643) );
  NAND2_X1 U9145 ( .A1(n6647), .A2(n6645), .ZN(n6644) );
  NAND2_X1 U9146 ( .A1(n8355), .A2(n6646), .ZN(n6645) );
  NAND2_X1 U9147 ( .A1(n8842), .A2(n6413), .ZN(n6646) );
  NAND2_X1 U9148 ( .A1(n6649), .A2(n6648), .ZN(n6647) );
  OAI21_X1 U9149 ( .B1(n8802), .B2(n8801), .A(n6580), .ZN(n6650) );
  AOI21_X1 U9150 ( .B1(n8802), .B2(n8801), .A(n6652), .ZN(n6651) );
  NAND2_X1 U9151 ( .A1(n6654), .A2(n6851), .ZN(n6653) );
  NAND3_X1 U9152 ( .A1(n6656), .A2(n6655), .A3(n6542), .ZN(n6654) );
  NAND2_X1 U9153 ( .A1(n6661), .A2(n8845), .ZN(n6655) );
  NAND2_X1 U9154 ( .A1(n6662), .A2(n8843), .ZN(n6656) );
  NAND2_X1 U9155 ( .A1(n6657), .A2(n6559), .ZN(n8723) );
  NAND3_X1 U9156 ( .A1(n6673), .A2(n6550), .A3(n6658), .ZN(n6657) );
  NAND2_X1 U9157 ( .A1(n8651), .A2(n8650), .ZN(n8669) );
  INV_X2 U9158 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6659) );
  INV_X1 U9159 ( .A(n6663), .ZN(n6661) );
  NAND2_X1 U9160 ( .A1(n6663), .A2(n8844), .ZN(n6662) );
  OAI22_X1 U9161 ( .A1(n6665), .A2(n6664), .B1(n8622), .B2(n8623), .ZN(n8646)
         );
  NAND3_X1 U9162 ( .A1(n8438), .A2(n6548), .A3(n8437), .ZN(n6667) );
  INV_X1 U9163 ( .A(n9106), .ZN(n6668) );
  AND2_X1 U9164 ( .A1(n9045), .A2(n7447), .ZN(n6670) );
  NAND2_X1 U9165 ( .A1(n6672), .A2(n6850), .ZN(n6671) );
  NAND2_X1 U9166 ( .A1(n8764), .A2(n8763), .ZN(n6672) );
  NAND2_X1 U9167 ( .A1(n6675), .A2(n6674), .ZN(n6673) );
  INV_X1 U9168 ( .A(n8667), .ZN(n6674) );
  NAND2_X1 U9169 ( .A1(n8669), .A2(n8668), .ZN(n6675) );
  NAND4_X1 U9170 ( .A1(n6912), .A2(n7561), .A3(n7411), .A4(n6519), .ZN(n7603)
         );
  NAND2_X1 U9171 ( .A1(n7415), .A2(n6505), .ZN(n12695) );
  NAND2_X1 U9172 ( .A1(n12724), .A2(n8198), .ZN(n6685) );
  INV_X1 U9173 ( .A(n12870), .ZN(n8185) );
  AND2_X1 U9174 ( .A1(n7631), .A2(n6690), .ZN(n6688) );
  NAND3_X1 U9175 ( .A1(n11529), .A2(n7619), .A3(P3_REG1_REG_1__SCAN_IN), .ZN(
        n6690) );
  NAND2_X1 U9176 ( .A1(n6692), .A2(n7630), .ZN(n10807) );
  AND2_X1 U9177 ( .A1(n7629), .A2(n6545), .ZN(n6692) );
  NAND2_X1 U9178 ( .A1(n10852), .A2(n12360), .ZN(n10213) );
  NAND2_X1 U9179 ( .A1(n10853), .A2(n12307), .ZN(n10852) );
  NAND2_X1 U9180 ( .A1(n10409), .A2(n12304), .ZN(n6693) );
  AND2_X2 U9181 ( .A1(n6698), .A2(n7620), .ZN(n7657) );
  OR2_X2 U9182 ( .A1(n12753), .A2(n12465), .ZN(n12754) );
  NAND2_X1 U9183 ( .A1(n10316), .A2(n12373), .ZN(n10315) );
  OAI21_X1 U9184 ( .B1(n6702), .B2(n12345), .A(n7255), .ZN(n10263) );
  OR2_X2 U9185 ( .A1(n12818), .A2(n8233), .ZN(n8234) );
  NAND2_X1 U9186 ( .A1(n13726), .A2(n7505), .ZN(n7502) );
  NAND2_X1 U9187 ( .A1(n13759), .A2(n13760), .ZN(n6704) );
  NAND3_X1 U9188 ( .A1(n6705), .A2(n6706), .A3(n6707), .ZN(n10505) );
  NAND2_X1 U9189 ( .A1(n7557), .A2(n6554), .ZN(n6705) );
  NAND3_X1 U9190 ( .A1(n6430), .A2(n10191), .A3(n7515), .ZN(n6706) );
  NAND2_X1 U9191 ( .A1(n10191), .A2(n6430), .ZN(n7557) );
  OAI211_X1 U9192 ( .C1(n12048), .C2(n6712), .A(n6711), .B(n7510), .ZN(n7508)
         );
  INV_X1 U9193 ( .A(n12053), .ZN(n6712) );
  NAND2_X1 U9194 ( .A1(n14560), .A2(n12053), .ZN(n13751) );
  NAND2_X1 U9195 ( .A1(n12048), .A2(n14555), .ZN(n14560) );
  NAND3_X1 U9196 ( .A1(n6713), .A2(n7518), .A3(n11121), .ZN(n11257) );
  NAND3_X1 U9197 ( .A1(n10785), .A2(n7520), .A3(n6828), .ZN(n6713) );
  OAI21_X1 U9198 ( .B1(n7611), .B2(n6717), .A(n6714), .ZN(n7677) );
  NAND2_X1 U9199 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U9200 ( .A1(n8030), .A2(n6456), .ZN(n8047) );
  AOI21_X1 U9201 ( .B1(n8030), .B2(n6720), .A(n6606), .ZN(n7104) );
  NAND2_X1 U9202 ( .A1(n7731), .A2(n7730), .ZN(n7733) );
  NAND2_X1 U9203 ( .A1(n12303), .A2(n12489), .ZN(n12326) );
  NAND2_X1 U9204 ( .A1(n7955), .A2(n7954), .ZN(n7956) );
  XNOR2_X1 U9205 ( .A(n12294), .B(n12293), .ZN(n12988) );
  NAND2_X1 U9206 ( .A1(n7921), .A2(n7920), .ZN(n7943) );
  NAND2_X1 U9207 ( .A1(n6740), .A2(n6747), .ZN(P3_U3296) );
  OAI21_X1 U9208 ( .B1(n6796), .B2(n6832), .A(n6748), .ZN(n6740) );
  AOI21_X1 U9209 ( .B1(n12490), .B2(n12497), .A(n6744), .ZN(n12491) );
  NAND2_X1 U9210 ( .A1(n12998), .A2(n12296), .ZN(n8164) );
  NAND2_X1 U9211 ( .A1(n7976), .A2(n7975), .ZN(n7993) );
  NAND2_X1 U9212 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  NOR2_X1 U9213 ( .A1(n9624), .A2(n9625), .ZN(n9726) );
  NAND2_X1 U9214 ( .A1(n13934), .A2(n13933), .ZN(n13936) );
  NAND2_X1 U9215 ( .A1(n9939), .A2(n9938), .ZN(n10090) );
  NAND2_X1 U9216 ( .A1(n7269), .A2(n12739), .ZN(n6745) );
  XNOR2_X1 U9217 ( .A(n8066), .B(n8048), .ZN(n11130) );
  AND2_X2 U9218 ( .A1(n11555), .A2(n11558), .ZN(n14694) );
  NAND2_X1 U9219 ( .A1(n7502), .A2(n7503), .ZN(n13691) );
  AOI21_X1 U9220 ( .B1(n13691), .B2(n13692), .A(n6551), .ZN(n12135) );
  NAND2_X1 U9221 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  NAND2_X1 U9222 ( .A1(n13939), .A2(n13938), .ZN(n14156) );
  NAND2_X1 U9223 ( .A1(n9929), .A2(n11558), .ZN(n10112) );
  NAND2_X1 U9224 ( .A1(n13784), .A2(n12093), .ZN(n13698) );
  NAND2_X1 U9225 ( .A1(n13716), .A2(n12086), .ZN(n13785) );
  NAND2_X1 U9226 ( .A1(n11257), .A2(n7541), .ZN(n11262) );
  NAND2_X1 U9227 ( .A1(n9630), .A2(n9629), .ZN(n9728) );
  NAND2_X1 U9228 ( .A1(n12988), .A2(n12296), .ZN(n7084) );
  INV_X1 U9229 ( .A(n10790), .ZN(n7519) );
  NAND2_X1 U9230 ( .A1(n6749), .A2(n6809), .ZN(P1_U3242) );
  OAI21_X1 U9231 ( .B1(n11913), .B2(n6812), .A(n6811), .ZN(n6749) );
  OAI21_X1 U9232 ( .B1(n6842), .B2(n6843), .A(n7495), .ZN(n11811) );
  NAND3_X1 U9233 ( .A1(n7542), .A2(n11564), .A3(n11563), .ZN(n11568) );
  OR2_X1 U9234 ( .A1(n11701), .A2(n11702), .ZN(n6815) );
  OAI21_X2 U9235 ( .B1(n8396), .B2(n8397), .A(n8399), .ZN(n8421) );
  NAND2_X1 U9236 ( .A1(n6962), .A2(n14772), .ZN(n6961) );
  NAND2_X1 U9237 ( .A1(n7508), .A2(n7509), .ZN(n13707) );
  NAND2_X1 U9238 ( .A1(n14219), .A2(n6577), .ZN(P1_U3554) );
  NAND2_X1 U9239 ( .A1(n14279), .A2(n6572), .ZN(P1_U3522) );
  NAND2_X1 U9240 ( .A1(n14267), .A2(n6480), .ZN(P1_U3527) );
  NAND2_X1 U9241 ( .A1(n14195), .A2(n6503), .ZN(P1_U3559) );
  NAND2_X1 U9242 ( .A1(n6992), .A2(n6991), .ZN(n14045) );
  NAND2_X1 U9243 ( .A1(n14138), .A2(n13920), .ZN(n14140) );
  NAND2_X1 U9244 ( .A1(n6789), .A2(n6752), .ZN(n14277) );
  NAND2_X1 U9245 ( .A1(n14212), .A2(n14751), .ZN(n6752) );
  OAI21_X2 U9246 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14385), .A(n14436), .ZN(
        n15366) );
  NOR2_X1 U9247 ( .A1(n14458), .A2(n14457), .ZN(n14456) );
  INV_X1 U9248 ( .A(n14380), .ZN(n6753) );
  NAND2_X1 U9249 ( .A1(n14485), .A2(n14484), .ZN(n14486) );
  AOI21_X2 U9250 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(n14413), .A(n14630), .ZN(
        n14636) );
  XNOR2_X1 U9251 ( .A(n6783), .B(n13993), .ZN(n14203) );
  NAND2_X1 U9252 ( .A1(n8425), .A2(n8424), .ZN(n8450) );
  INV_X1 U9253 ( .A(n7166), .ZN(n7164) );
  NAND2_X1 U9254 ( .A1(n8748), .A2(n7545), .ZN(n8750) );
  OAI21_X2 U9255 ( .B1(n8788), .B2(n8787), .A(n8789), .ZN(n8808) );
  AND3_X2 U9256 ( .A1(n7265), .A2(n7264), .A3(n12713), .ZN(n12711) );
  OAI21_X1 U9257 ( .B1(n12718), .B2(n15149), .A(n12717), .ZN(n12894) );
  NAND2_X1 U9258 ( .A1(n10007), .A2(n10008), .ZN(n10006) );
  NOR2_X1 U9259 ( .A1(n14498), .A2(n12551), .ZN(n12580) );
  NOR2_X1 U9260 ( .A1(n10911), .A2(n10912), .ZN(n15100) );
  NOR2_X1 U9261 ( .A1(n12523), .A2(n12524), .ZN(n12526) );
  INV_X1 U9262 ( .A(n9828), .ZN(n7626) );
  INV_X1 U9263 ( .A(n6975), .ZN(n6803) );
  NAND2_X2 U9264 ( .A1(n8140), .A2(n7606), .ZN(n8068) );
  NAND2_X1 U9265 ( .A1(n10855), .A2(n12356), .ZN(n10854) );
  NAND2_X1 U9266 ( .A1(n12735), .A2(n12739), .ZN(n12734) );
  AOI21_X1 U9267 ( .B1(n12891), .B2(n15177), .A(n12890), .ZN(n12946) );
  NAND2_X1 U9268 ( .A1(n10804), .A2(n15139), .ZN(n8166) );
  NAND2_X1 U9269 ( .A1(n8185), .A2(n7420), .ZN(n8186) );
  NAND2_X1 U9270 ( .A1(n6689), .A2(n10801), .ZN(n8224) );
  NAND2_X1 U9271 ( .A1(n7413), .A2(n7412), .ZN(n7558) );
  INV_X1 U9272 ( .A(n6471), .ZN(n7604) );
  NAND2_X1 U9273 ( .A1(n12838), .A2(n12837), .ZN(n12836) );
  NAND2_X1 U9274 ( .A1(n7356), .A2(n7355), .ZN(n8534) );
  NAND2_X1 U9275 ( .A1(n8537), .A2(n8536), .ZN(n8555) );
  INV_X2 U9276 ( .A(n8376), .ZN(n8330) );
  NAND2_X1 U9277 ( .A1(n7489), .A2(n11745), .ZN(n7488) );
  NOR2_X2 U9278 ( .A1(n14456), .A2(n14396), .ZN(n14398) );
  XNOR2_X1 U9279 ( .A(n14424), .B(n7016), .ZN(n14479) );
  AOI22_X1 U9280 ( .A1(n13298), .A2(n13297), .B1(n13296), .B2(n13509), .ZN(
        n13515) );
  INV_X1 U9281 ( .A(n10152), .ZN(n10383) );
  INV_X1 U9282 ( .A(n11412), .ZN(n6801) );
  NOR2_X1 U9283 ( .A1(n15371), .A2(n15370), .ZN(n15369) );
  AOI21_X2 U9284 ( .B1(n11186), .B2(n11169), .A(n11168), .ZN(n11239) );
  NAND3_X2 U9285 ( .A1(n6472), .A2(n9278), .A3(n6791), .ZN(n13837) );
  OAI21_X2 U9286 ( .B1(n7288), .B2(n14677), .A(n6964), .ZN(n14176) );
  NAND2_X1 U9287 ( .A1(n7037), .A2(n13283), .ZN(n13400) );
  NAND2_X1 U9288 ( .A1(n7029), .A2(n7028), .ZN(n13343) );
  NAND2_X1 U9289 ( .A1(n7039), .A2(n7038), .ZN(n13430) );
  AND2_X2 U9290 ( .A1(n10616), .A2(n10385), .ZN(n10538) );
  NAND2_X1 U9291 ( .A1(n7558), .A2(n8225), .ZN(n10410) );
  NOR2_X2 U9292 ( .A1(n6772), .A2(n7579), .ZN(n7411) );
  NAND2_X1 U9293 ( .A1(n6489), .A2(n7337), .ZN(n6772) );
  NAND2_X1 U9294 ( .A1(n14416), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U9295 ( .A1(n14392), .A2(n15358), .ZN(n14393) );
  XNOR2_X1 U9296 ( .A(n14382), .B(n14383), .ZN(n15370) );
  NAND2_X1 U9297 ( .A1(n6961), .A2(n6959), .ZN(P1_U3557) );
  OAI22_X1 U9298 ( .A1(n12047), .A2(n9906), .B1(n13842), .B2(n9560), .ZN(n9561) );
  NAND3_X1 U9299 ( .A1(n9566), .A2(n9565), .A3(n6778), .ZN(n9628) );
  OAI22_X1 U9300 ( .A1(n9732), .A2(n12047), .B1(n9563), .B2(n14717), .ZN(n9623) );
  NAND3_X1 U9301 ( .A1(n6782), .A2(n6781), .A3(n9332), .ZN(n13154) );
  NAND2_X1 U9302 ( .A1(n6947), .A2(n6948), .ZN(n6783) );
  NAND2_X1 U9303 ( .A1(n7359), .A2(n7360), .ZN(n8725) );
  NAND2_X1 U9304 ( .A1(n8555), .A2(n8554), .ZN(n8558) );
  NAND2_X1 U9305 ( .A1(n8473), .A2(n8472), .ZN(n6945) );
  NAND2_X1 U9306 ( .A1(n8727), .A2(n8726), .ZN(n8748) );
  NAND2_X1 U9307 ( .A1(n7377), .A2(n7378), .ZN(n8624) );
  NAND3_X1 U9308 ( .A1(n6788), .A2(n6787), .A3(n6439), .ZN(n6786) );
  NAND2_X1 U9309 ( .A1(n7242), .A2(n13288), .ZN(n7241) );
  NAND2_X1 U9310 ( .A1(n7220), .A2(n13285), .ZN(n7219) );
  NAND2_X1 U9311 ( .A1(n13336), .A2(n13323), .ZN(n13338) );
  NAND2_X1 U9312 ( .A1(n6852), .A2(n6608), .ZN(n8160) );
  NAND2_X4 U9313 ( .A1(n14314), .A2(n9275), .ZN(n11820) );
  NAND2_X1 U9314 ( .A1(n13785), .A2(n13786), .ZN(n13784) );
  OAI21_X1 U9315 ( .B1(n14274), .B2(n6820), .A(n6818), .ZN(P1_U3555) );
  NAND2_X1 U9316 ( .A1(n6792), .A2(n7262), .ZN(n6832) );
  AOI21_X1 U9317 ( .B1(n7856), .B2(n7855), .A(n7854), .ZN(n7858) );
  NAND2_X1 U9318 ( .A1(n7957), .A2(n7091), .ZN(n7973) );
  NAND2_X1 U9319 ( .A1(n7085), .A2(n6582), .ZN(n7822) );
  NAND3_X1 U9320 ( .A1(n12473), .A2(n12727), .A3(n12474), .ZN(n12475) );
  OR2_X1 U9321 ( .A1(n6793), .A2(n12469), .ZN(n12473) );
  OAI21_X1 U9322 ( .B1(n12491), .B2(n15150), .A(n6797), .ZN(n6796) );
  NAND2_X1 U9323 ( .A1(n12491), .A2(n12492), .ZN(n6797) );
  INV_X1 U9324 ( .A(n14636), .ZN(n6799) );
  NAND2_X1 U9325 ( .A1(n10387), .A2(n10386), .ZN(n10536) );
  AOI21_X2 U9326 ( .B1(n6801), .B2(n6428), .A(n6540), .ZN(n11504) );
  NOR2_X1 U9327 ( .A1(n11329), .A2(n14508), .ZN(n12523) );
  NAND3_X1 U9328 ( .A1(n6804), .A2(n6803), .A3(n6931), .ZN(P3_U3201) );
  INV_X1 U9329 ( .A(n6986), .ZN(n9880) );
  XNOR2_X1 U9330 ( .A(n12639), .B(n6806), .ZN(n12664) );
  NAND2_X1 U9331 ( .A1(n8166), .A2(n7414), .ZN(n7413) );
  XNOR2_X1 U9332 ( .A(n8808), .B(SI_20_), .ZN(n8807) );
  INV_X1 U9333 ( .A(n8846), .ZN(n6816) );
  NAND3_X1 U9334 ( .A1(n6535), .A2(n11703), .A3(n6815), .ZN(n6814) );
  OAI21_X2 U9335 ( .B1(n8908), .B2(n8907), .A(n8894), .ZN(n8932) );
  NAND2_X1 U9336 ( .A1(n13338), .A2(n6817), .ZN(n13287) );
  NAND3_X1 U9337 ( .A1(n7368), .A2(n7370), .A3(n7369), .ZN(n8846) );
  NAND2_X1 U9338 ( .A1(n11765), .A2(n11764), .ZN(n11778) );
  NOR2_X2 U9339 ( .A1(n6913), .A2(n7648), .ZN(n7805) );
  NAND3_X1 U9340 ( .A1(n7801), .A2(n7560), .A3(n7565), .ZN(n6913) );
  NAND2_X1 U9341 ( .A1(n7028), .A2(n13124), .ZN(n6817) );
  NAND3_X1 U9342 ( .A1(n9240), .A2(n9230), .A3(n9229), .ZN(n6821) );
  NAND2_X1 U9343 ( .A1(n7604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7616) );
  OAI21_X1 U9344 ( .B1(n14274), .B2(n14763), .A(n6822), .ZN(P1_U3523) );
  NAND2_X1 U9345 ( .A1(n12695), .A2(n6482), .ZN(n8211) );
  NAND2_X1 U9346 ( .A1(n13698), .A2(n13699), .ZN(n12101) );
  NOR2_X2 U9347 ( .A1(n12527), .A2(n12528), .ZN(n12568) );
  NOR2_X2 U9348 ( .A1(n6917), .A2(n6920), .ZN(n12527) );
  NOR2_X1 U9349 ( .A1(n9854), .A2(n6553), .ZN(n9832) );
  NOR2_X1 U9350 ( .A1(n12571), .A2(n12572), .ZN(n12598) );
  XNOR2_X1 U9351 ( .A(n12596), .B(n12597), .ZN(n12571) );
  XOR2_X2 U9352 ( .A(n12640), .B(n12651), .Z(n12619) );
  NAND2_X1 U9353 ( .A1(n6915), .A2(n7543), .ZN(n6914) );
  INV_X1 U9354 ( .A(n10010), .ZN(n7180) );
  NAND3_X1 U9355 ( .A1(n6826), .A2(n6825), .A3(n7488), .ZN(n7487) );
  NAND2_X1 U9356 ( .A1(n11734), .A2(n11733), .ZN(n6825) );
  NAND2_X1 U9357 ( .A1(n11730), .A2(n11729), .ZN(n6826) );
  NAND2_X1 U9358 ( .A1(n11504), .A2(n7540), .ZN(n7052) );
  NAND2_X1 U9359 ( .A1(n13513), .A2(n6583), .ZN(n13491) );
  AOI21_X2 U9360 ( .B1(n10446), .B2(n6485), .A(n6434), .ZN(n10742) );
  NAND2_X2 U9361 ( .A1(n13378), .A2(n13317), .ZN(n13365) );
  OAI21_X1 U9362 ( .B1(n7047), .B2(n7049), .A(n7046), .ZN(n11041) );
  NAND3_X1 U9363 ( .A1(n8186), .A2(n12860), .A3(n8187), .ZN(n12851) );
  INV_X1 U9364 ( .A(n13707), .ZN(n6870) );
  INV_X1 U9366 ( .A(n10194), .ZN(n7517) );
  XNOR2_X1 U9367 ( .A(n6830), .B(n9724), .ZN(n10250) );
  OAI22_X1 U9368 ( .A1(n6990), .A2(n9563), .B1(n10185), .B2(n12047), .ZN(n6830) );
  INV_X1 U9369 ( .A(n12047), .ZN(n10254) );
  AND2_X1 U9370 ( .A1(n9624), .A2(n9625), .ZN(n9626) );
  NOR2_X1 U9371 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9114) );
  NAND2_X1 U9372 ( .A1(n10430), .A2(n7723), .ZN(n10677) );
  NAND2_X1 U9373 ( .A1(n7319), .A2(n7318), .ZN(n12210) );
  OR2_X2 U9374 ( .A1(n7797), .A2(n7796), .ZN(n11456) );
  NAND2_X1 U9375 ( .A1(n8097), .A2(n8098), .ZN(n12005) );
  NAND2_X1 U9376 ( .A1(n6895), .A2(n6893), .ZN(n12197) );
  NAND2_X1 U9377 ( .A1(n14479), .A2(n15294), .ZN(n14478) );
  NAND2_X1 U9378 ( .A1(n7017), .A2(n14648), .ZN(n14424) );
  NAND2_X1 U9379 ( .A1(n14378), .A2(n14377), .ZN(n7013) );
  NAND2_X1 U9380 ( .A1(n7679), .A2(n7678), .ZN(n7700) );
  NOR2_X1 U9381 ( .A1(n6827), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U9382 ( .A1(n7022), .A2(n14486), .ZN(n7021) );
  XNOR2_X1 U9383 ( .A(n7021), .B(n7020), .ZN(SUB_1596_U4) );
  AND2_X2 U9384 ( .A1(n7455), .A2(n8292), .ZN(n8320) );
  AOI21_X1 U9385 ( .B1(n13478), .B2(n7074), .A(n7072), .ZN(n7071) );
  INV_X1 U9386 ( .A(n10744), .ZN(n7047) );
  NAND2_X1 U9387 ( .A1(n7055), .A2(n7054), .ZN(n13340) );
  NAND2_X1 U9388 ( .A1(n10006), .A2(n9778), .ZN(n9779) );
  NAND3_X1 U9389 ( .A1(n6837), .A2(n6836), .A3(n8295), .ZN(n7457) );
  NAND2_X1 U9390 ( .A1(n9849), .A2(n9781), .ZN(n9782) );
  NAND2_X1 U9391 ( .A1(n10090), .A2(n10089), .ZN(n6838) );
  OAI22_X2 U9392 ( .A1(n11878), .A2(n9610), .B1(n13837), .B2(n9609), .ZN(n9952) );
  NAND2_X1 U9393 ( .A1(n11383), .A2(n11892), .ZN(n13975) );
  NAND2_X1 U9394 ( .A1(n14704), .A2(n14703), .ZN(n7315) );
  NAND2_X1 U9395 ( .A1(n13980), .A2(n13979), .ZN(n14144) );
  INV_X1 U9396 ( .A(n14127), .ZN(n6966) );
  NAND2_X1 U9397 ( .A1(n14176), .A2(n7146), .ZN(n10597) );
  NOR3_X1 U9398 ( .A1(n11866), .A2(n11872), .A3(n11905), .ZN(n11913) );
  NAND2_X1 U9399 ( .A1(n10319), .A2(n10318), .ZN(n10317) );
  NAND2_X1 U9400 ( .A1(n11816), .A2(n11815), .ZN(n11847) );
  NAND2_X1 U9401 ( .A1(n11619), .A2(n11618), .ZN(n7466) );
  NAND2_X1 U9402 ( .A1(n7470), .A2(n7468), .ZN(n6847) );
  NAND2_X1 U9403 ( .A1(n6847), .A2(n6846), .ZN(n11627) );
  NAND2_X1 U9404 ( .A1(n7504), .A2(n12115), .ZN(n13801) );
  NAND3_X1 U9405 ( .A1(n7497), .A2(n11573), .A3(n11572), .ZN(n6841) );
  NAND2_X1 U9406 ( .A1(n11782), .A2(n6557), .ZN(n6842) );
  NAND2_X1 U9407 ( .A1(n13685), .A2(n9005), .ZN(n8897) );
  NAND4_X1 U9408 ( .A1(n14487), .A2(n7041), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7040) );
  NAND3_X1 U9409 ( .A1(n13556), .A2(n6406), .A3(n6565), .ZN(n13653) );
  INV_X1 U9410 ( .A(n8471), .ZN(n8472) );
  NAND4_X1 U9411 ( .A1(n11228), .A2(n13252), .A3(n7043), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U9412 ( .A1(n12987), .A2(n6476), .ZN(n7590) );
  AOI21_X2 U9413 ( .B1(n7585), .B2(n11131), .A(n6848), .ZN(n9424) );
  NAND3_X1 U9414 ( .A1(n7368), .A2(n7370), .A3(n7367), .ZN(n6849) );
  NAND2_X1 U9415 ( .A1(n10432), .A2(n10431), .ZN(n10430) );
  INV_X1 U9416 ( .A(n12210), .ZN(n6908) );
  NAND2_X1 U9417 ( .A1(n7997), .A2(n7996), .ZN(n7345) );
  NAND2_X1 U9418 ( .A1(n6885), .A2(n6883), .ZN(n7319) );
  NAND2_X1 U9419 ( .A1(n7806), .A2(n7411), .ZN(n7597) );
  OAI21_X1 U9420 ( .B1(n7169), .B2(n7164), .A(n7165), .ZN(n7163) );
  NAND2_X1 U9421 ( .A1(n12734), .A2(n7556), .ZN(n12724) );
  AOI21_X1 U9422 ( .B1(n15164), .B2(n12895), .A(n12894), .ZN(n12949) );
  NAND2_X2 U9423 ( .A1(n8319), .A2(n8318), .ZN(n8842) );
  NAND2_X1 U9424 ( .A1(n12501), .A2(n6476), .ZN(n7262) );
  NAND2_X1 U9425 ( .A1(n6862), .A2(n6860), .ZN(P3_U3487) );
  OR2_X1 U9426 ( .A1(n12946), .A2(n15196), .ZN(n6862) );
  NAND2_X1 U9427 ( .A1(n6865), .A2(n6863), .ZN(P3_U3455) );
  OR2_X1 U9428 ( .A1(n12946), .A2(n15187), .ZN(n6865) );
  OAI21_X2 U9429 ( .B1(n8376), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6866), .ZN(
        n8372) );
  OAI21_X1 U9430 ( .B1(n8046), .B2(n7105), .A(n7104), .ZN(n8082) );
  NAND2_X1 U9431 ( .A1(n10078), .A2(n11791), .ZN(n6972) );
  NAND4_X1 U9432 ( .A1(n9212), .A2(n9113), .A3(n9639), .A4(n9114), .ZN(n6868)
         );
  NAND2_X1 U9433 ( .A1(n7215), .A2(n13321), .ZN(n7211) );
  XNOR2_X1 U9434 ( .A(n8932), .B(n8895), .ZN(n13685) );
  INV_X1 U9435 ( .A(n7208), .ZN(n13336) );
  XNOR2_X2 U9436 ( .A(n13373), .B(n13318), .ZN(n7216) );
  NAND2_X1 U9437 ( .A1(n7733), .A2(n7732), .ZN(n7754) );
  NAND2_X1 U9438 ( .A1(n7080), .A2(n7756), .ZN(n7764) );
  NAND2_X1 U9439 ( .A1(n7754), .A2(n7753), .ZN(n7080) );
  NAND2_X1 U9440 ( .A1(n7946), .A2(n7945), .ZN(n7955) );
  INV_X1 U9441 ( .A(n7640), .ZN(n7607) );
  NAND2_X1 U9442 ( .A1(n6876), .A2(n6873), .ZN(P3_U3486) );
  OR2_X1 U9443 ( .A1(n12949), .A2(n15196), .ZN(n6876) );
  NAND2_X1 U9444 ( .A1(n13948), .A2(n13947), .ZN(n14093) );
  NAND2_X1 U9445 ( .A1(n8421), .A2(n8420), .ZN(n8425) );
  AND2_X2 U9446 ( .A1(n7042), .A2(n7040), .ZN(n8376) );
  NAND2_X1 U9447 ( .A1(n8454), .A2(n8453), .ZN(n8473) );
  NAND2_X1 U9448 ( .A1(n8624), .A2(n7553), .ZN(n8626) );
  XNOR2_X1 U9449 ( .A(n13287), .B(n13325), .ZN(n7242) );
  OAI21_X1 U9450 ( .B1(n7212), .B2(n13353), .A(n6566), .ZN(n7210) );
  INV_X1 U9451 ( .A(n7210), .ZN(n7209) );
  NOR2_X2 U9452 ( .A1(n10164), .A2(n9784), .ZN(n9994) );
  NOR2_X2 U9453 ( .A1(n10165), .A2(n10221), .ZN(n10164) );
  OAI21_X1 U9454 ( .B1(n10026), .B2(n9847), .A(n9846), .ZN(n9849) );
  NOR2_X2 U9455 ( .A1(n12637), .A2(n12636), .ZN(n12639) );
  NOR2_X1 U9456 ( .A1(n12580), .A2(n12581), .ZN(n12585) );
  OR2_X2 U9457 ( .A1(n12526), .A2(n12540), .ZN(n6974) );
  NAND2_X1 U9458 ( .A1(n12241), .A2(n6886), .ZN(n6885) );
  NAND2_X1 U9459 ( .A1(n7340), .A2(n6896), .ZN(n6895) );
  NOR2_X2 U9460 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7646) );
  NAND2_X1 U9461 ( .A1(n12269), .A2(n8080), .ZN(n8097) );
  OAI211_X1 U9462 ( .C1(n12269), .C2(n6905), .A(n6902), .B(n6900), .ZN(n12013)
         );
  OAI22_X1 U9463 ( .A1(n6904), .A2(n6901), .B1(n12007), .B2(n6906), .ZN(n6900)
         );
  NOR2_X1 U9464 ( .A1(n12007), .A2(n8098), .ZN(n6901) );
  NAND2_X1 U9465 ( .A1(n12269), .A2(n6903), .ZN(n6902) );
  NOR2_X1 U9466 ( .A1(n12007), .A2(n6904), .ZN(n6903) );
  NAND2_X1 U9467 ( .A1(n8098), .A2(n12007), .ZN(n6905) );
  NAND2_X1 U9468 ( .A1(n10646), .A2(n10647), .ZN(n6910) );
  OAI21_X1 U9469 ( .B1(n7341), .B2(n6911), .A(n6909), .ZN(n10635) );
  NAND4_X1 U9470 ( .A1(n6910), .A2(n10525), .A3(n6528), .A4(n7343), .ZN(n6909)
         );
  OAI21_X2 U9471 ( .B1(n10677), .B2(n7348), .A(n7346), .ZN(n11207) );
  INV_X1 U9472 ( .A(n6913), .ZN(n6912) );
  NOR2_X1 U9473 ( .A1(n6914), .A2(n9798), .ZN(n10166) );
  AND2_X1 U9474 ( .A1(n6914), .A2(n9798), .ZN(n10167) );
  INV_X1 U9475 ( .A(n9833), .ZN(n6915) );
  NAND2_X1 U9476 ( .A1(n6918), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6917) );
  INV_X1 U9477 ( .A(n6920), .ZN(n6919) );
  AOI21_X2 U9478 ( .B1(n7179), .B2(n7178), .A(n12532), .ZN(n6920) );
  NAND2_X1 U9479 ( .A1(n7180), .A2(n6924), .ZN(n6927) );
  NAND2_X1 U9480 ( .A1(n6927), .A2(n6926), .ZN(n9829) );
  XNOR2_X2 U9481 ( .A(n6929), .B(n9883), .ZN(n9835) );
  NOR2_X1 U9482 ( .A1(n12619), .A2(n12618), .ZN(n12642) );
  NAND2_X1 U9483 ( .A1(n6934), .A2(n6935), .ZN(n12683) );
  NAND2_X1 U9484 ( .A1(n10891), .A2(n10890), .ZN(n15091) );
  AND2_X1 U9485 ( .A1(n15091), .A2(n10892), .ZN(n11304) );
  NAND2_X1 U9486 ( .A1(n6946), .A2(n6950), .ZN(n14008) );
  OR2_X1 U9487 ( .A1(n14030), .A2(n6952), .ZN(n6946) );
  NAND2_X1 U9488 ( .A1(n14030), .A2(n6950), .ZN(n6948) );
  OR2_X2 U9489 ( .A1(n6956), .A2(n13991), .ZN(n6953) );
  INV_X1 U9490 ( .A(n6965), .ZN(n6964) );
  OAI21_X1 U9491 ( .B1(n14677), .B2(n7289), .A(n10595), .ZN(n6965) );
  OAI21_X2 U9492 ( .B1(n14144), .B2(n14146), .A(n13981), .ZN(n14127) );
  NAND2_X1 U9493 ( .A1(n6969), .A2(n6967), .ZN(n11336) );
  XNOR2_X1 U9494 ( .A(n8422), .B(SI_3_), .ZN(n8420) );
  MUX2_X1 U9495 ( .A(n9143), .B(n9141), .S(n8330), .Z(n8422) );
  INV_X1 U9496 ( .A(n6974), .ZN(n12550) );
  OAI21_X1 U9497 ( .B1(n12639), .B2(n6979), .A(n6978), .ZN(n6975) );
  NAND3_X1 U9498 ( .A1(n12639), .A2(n6983), .A3(n6977), .ZN(n6976) );
  NAND2_X1 U9499 ( .A1(n12666), .A2(n12665), .ZN(n6980) );
  XNOR2_X2 U9500 ( .A(n9876), .B(n9894), .ZN(n9787) );
  NOR2_X2 U9501 ( .A1(n9992), .A2(n9786), .ZN(n9876) );
  NOR2_X2 U9502 ( .A1(n9994), .A2(n9993), .ZN(n9992) );
  AND2_X2 U9503 ( .A1(n12613), .A2(n12612), .ZN(n12635) );
  NOR2_X2 U9504 ( .A1(n10329), .A2(n10882), .ZN(n10911) );
  OR2_X2 U9505 ( .A1(n11325), .A2(n11326), .ZN(n6988) );
  XNOR2_X2 U9506 ( .A(n11323), .B(n11324), .ZN(n10915) );
  NOR2_X2 U9508 ( .A1(n14098), .A2(n14232), .ZN(n6992) );
  NAND2_X1 U9509 ( .A1(n8292), .A2(n6449), .ZN(n9077) );
  NOR2_X2 U9510 ( .A1(n13368), .A2(n13568), .ZN(n7029) );
  NAND2_X1 U9511 ( .A1(n13646), .A2(n11418), .ZN(n11506) );
  NOR2_X2 U9512 ( .A1(n11192), .A2(n7035), .ZN(n11418) );
  NOR2_X2 U9513 ( .A1(n13430), .A2(n13410), .ZN(n7037) );
  INV_X1 U9514 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7043) );
  INV_X1 U9515 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7041) );
  NAND2_X1 U9516 ( .A1(n13365), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U9517 ( .A1(n13365), .A2(n13320), .ZN(n7060) );
  INV_X1 U9518 ( .A(n13409), .ZN(n7069) );
  INV_X1 U9519 ( .A(n7071), .ZN(n13308) );
  NAND2_X1 U9520 ( .A1(n7973), .A2(n7972), .ZN(n7976) );
  NAND2_X1 U9521 ( .A1(n7092), .A2(n7093), .ZN(n7921) );
  INV_X1 U9522 ( .A(n8201), .ZN(n7102) );
  NAND2_X2 U9523 ( .A1(n9652), .A2(n10369), .ZN(n7108) );
  NAND2_X4 U9524 ( .A1(n7108), .A2(n8354), .ZN(n11976) );
  NAND2_X1 U9525 ( .A1(n15059), .A2(n7108), .ZN(n14999) );
  OR2_X1 U9526 ( .A1(n15028), .A2(n7108), .ZN(n15034) );
  NAND2_X1 U9527 ( .A1(n13122), .A2(n7109), .ZN(n13006) );
  NAND2_X1 U9528 ( .A1(n13094), .A2(n6562), .ZN(n13042) );
  NAND2_X1 U9529 ( .A1(n11925), .A2(n7120), .ZN(n7118) );
  OAI21_X1 U9530 ( .B1(n13095), .B2(n7122), .A(n6544), .ZN(n7121) );
  NAND2_X1 U9531 ( .A1(n7128), .A2(n6500), .ZN(n7127) );
  OR2_X1 U9532 ( .A1(n10492), .A2(n10493), .ZN(n7128) );
  NAND3_X1 U9533 ( .A1(n7129), .A2(n7127), .A3(n11991), .ZN(n11998) );
  NAND3_X1 U9534 ( .A1(n6500), .A2(n7131), .A3(n7133), .ZN(n7129) );
  NOR2_X1 U9535 ( .A1(n14778), .A2(n7132), .ZN(n7131) );
  OR2_X1 U9536 ( .A1(n10485), .A2(n10484), .ZN(n7133) );
  INV_X1 U9537 ( .A(n7135), .ZN(n14776) );
  NAND4_X1 U9538 ( .A1(n9240), .A2(n9230), .A3(n9229), .A4(n7492), .ZN(n9272)
         );
  NAND2_X1 U9539 ( .A1(n14048), .A2(n6556), .ZN(n7150) );
  NOR2_X4 U9540 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9130) );
  NAND2_X1 U9541 ( .A1(n7169), .A2(n14751), .ZN(n7167) );
  NAND2_X1 U9542 ( .A1(n7163), .A2(n7168), .ZN(P1_U3525) );
  NOR2_X1 U9543 ( .A1(n11344), .A2(n11343), .ZN(n11345) );
  OR2_X2 U9544 ( .A1(n15117), .A2(n15116), .ZN(n7179) );
  OAI21_X2 U9545 ( .B1(n7649), .B2(n7182), .A(n7181), .ZN(n10010) );
  OR2_X2 U9546 ( .A1(n10166), .A2(n9833), .ZN(n7187) );
  INV_X2 U9547 ( .A(n9275), .ZN(n11531) );
  NOR2_X4 U9548 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9212) );
  NOR2_X2 U9549 ( .A1(n10025), .A2(n9810), .ZN(n10024) );
  NAND2_X1 U9550 ( .A1(n11510), .A2(n11509), .ZN(n7207) );
  NAND2_X1 U9551 ( .A1(n7207), .A2(n7205), .ZN(n13266) );
  OAI21_X1 U9552 ( .B1(n13392), .B2(n7211), .A(n7209), .ZN(n7208) );
  NAND2_X1 U9553 ( .A1(n7223), .A2(n7227), .ZN(n11174) );
  NAND2_X1 U9554 ( .A1(n10925), .A2(n7224), .ZN(n7223) );
  NAND2_X1 U9555 ( .A1(n7232), .A2(n7230), .ZN(n11245) );
  NOR2_X1 U9556 ( .A1(n7231), .A2(n6530), .ZN(n7230) );
  NAND2_X1 U9557 ( .A1(n7235), .A2(n7233), .ZN(n10727) );
  INV_X1 U9558 ( .A(n7234), .ZN(n7233) );
  OAI21_X1 U9559 ( .B1(n10392), .B2(n7238), .A(n10722), .ZN(n7234) );
  NAND2_X1 U9560 ( .A1(n10393), .A2(n7236), .ZN(n7235) );
  INV_X1 U9561 ( .A(n9052), .ZN(n10621) );
  XNOR2_X1 U9562 ( .A(n13144), .B(n9052), .ZN(n10604) );
  OR2_X1 U9563 ( .A1(n8455), .A2(n9604), .ZN(n7243) );
  NAND2_X1 U9564 ( .A1(n7255), .A2(n12340), .ZN(n10409) );
  OAI21_X1 U9565 ( .B1(n10840), .B2(n7275), .A(n7271), .ZN(n11089) );
  NAND3_X1 U9566 ( .A1(n7805), .A2(n7411), .A3(n6558), .ZN(n7595) );
  NAND2_X1 U9567 ( .A1(n10271), .A2(n7287), .ZN(n7288) );
  OR2_X2 U9568 ( .A1(n14113), .A2(n7299), .ZN(n7294) );
  OAI21_X1 U9569 ( .B1(n14113), .B2(n13984), .A(n7301), .ZN(n14096) );
  NAND2_X1 U9570 ( .A1(n14061), .A2(n7305), .ZN(n7304) );
  OAI21_X2 U9572 ( .B1(n7315), .B2(n7314), .A(n7312), .ZN(n10069) );
  NAND4_X1 U9573 ( .A1(n9240), .A2(n9230), .A3(n9232), .A4(n9229), .ZN(n7316)
         );
  INV_X2 U9574 ( .A(n7811), .ZN(n7654) );
  INV_X1 U9575 ( .A(n7633), .ZN(n7317) );
  XNOR2_X1 U9576 ( .A(n7811), .B(n10807), .ZN(n7633) );
  NAND2_X1 U9577 ( .A1(n11456), .A2(n6587), .ZN(n7325) );
  NAND2_X1 U9578 ( .A1(n11457), .A2(n7818), .ZN(n7324) );
  NAND2_X1 U9579 ( .A1(n7324), .A2(n6571), .ZN(n7326) );
  NAND2_X1 U9580 ( .A1(n7953), .A2(n7328), .ZN(n12165) );
  NAND2_X1 U9581 ( .A1(n12165), .A2(n12167), .ZN(n7989) );
  NOR2_X1 U9582 ( .A1(n7591), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U9583 ( .A1(n6437), .A2(n7332), .ZN(n7862) );
  NOR2_X1 U9584 ( .A1(n7591), .A2(n7333), .ZN(n7332) );
  NOR2_X1 U9585 ( .A1(n7591), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U9586 ( .A1(n7670), .A2(n10641), .ZN(n7343) );
  CLKBUF_X1 U9587 ( .A(n8008), .Z(n7344) );
  NAND3_X1 U9588 ( .A1(n7345), .A2(n8008), .A3(n8007), .ZN(n12251) );
  NAND2_X1 U9589 ( .A1(n7999), .A2(n7998), .ZN(n8008) );
  AND2_X1 U9590 ( .A1(n7909), .A2(n7351), .ZN(n7569) );
  NAND2_X1 U9591 ( .A1(n7909), .A2(n7350), .ZN(n7571) );
  NAND2_X1 U9592 ( .A1(n6878), .A2(n7357), .ZN(n7356) );
  NAND2_X1 U9593 ( .A1(n8652), .A2(n7363), .ZN(n7359) );
  NAND2_X1 U9594 ( .A1(n8652), .A2(n7554), .ZN(n7362) );
  INV_X1 U9595 ( .A(n8829), .ZN(n7366) );
  NAND2_X1 U9596 ( .A1(n7366), .A2(SI_22_), .ZN(n7368) );
  NAND3_X1 U9597 ( .A1(n7373), .A2(n6597), .A3(n7372), .ZN(n8890) );
  NAND2_X1 U9598 ( .A1(n8869), .A2(n7374), .ZN(n7372) );
  OR2_X2 U9599 ( .A1(n8869), .A2(n7376), .ZN(n7373) );
  NAND3_X1 U9600 ( .A1(n7373), .A2(n6455), .A3(n7372), .ZN(n8886) );
  NAND2_X1 U9601 ( .A1(n8558), .A2(n6546), .ZN(n7377) );
  NAND3_X1 U9602 ( .A1(n7381), .A2(n8578), .A3(n7380), .ZN(n7379) );
  NAND2_X1 U9603 ( .A1(n8750), .A2(n7384), .ZN(n7383) );
  NAND2_X1 U9604 ( .A1(n7383), .A2(n6586), .ZN(n8788) );
  OAI21_X1 U9605 ( .B1(n8976), .B2(n8975), .A(n8938), .ZN(n8961) );
  NAND2_X1 U9606 ( .A1(n12345), .A2(n8168), .ZN(n7412) );
  AND2_X1 U9607 ( .A1(n8168), .A2(n8165), .ZN(n7414) );
  NAND2_X1 U9608 ( .A1(n7418), .A2(n7419), .ZN(n8184) );
  NAND2_X1 U9609 ( .A1(n8183), .A2(n7421), .ZN(n7418) );
  NAND2_X1 U9610 ( .A1(n12851), .A2(n8188), .ZN(n12838) );
  NAND2_X1 U9611 ( .A1(n7426), .A2(n7425), .ZN(n8181) );
  AND2_X1 U9612 ( .A1(n12982), .A2(n8191), .ZN(n7438) );
  NAND2_X1 U9613 ( .A1(n9044), .A2(n6555), .ZN(n7447) );
  INV_X1 U9614 ( .A(n8552), .ZN(n7448) );
  INV_X1 U9615 ( .A(n8551), .ZN(n7449) );
  INV_X1 U9616 ( .A(n8823), .ZN(n7452) );
  NAND3_X1 U9617 ( .A1(n8284), .A2(n8417), .A3(n8288), .ZN(n8654) );
  NAND2_X1 U9618 ( .A1(n8646), .A2(n8647), .ZN(n8645) );
  NAND3_X1 U9619 ( .A1(n7464), .A2(n7462), .A3(n9584), .ZN(n11535) );
  NAND3_X1 U9620 ( .A1(n7467), .A2(n7466), .A3(n7471), .ZN(n7470) );
  NAND2_X1 U9621 ( .A1(n11615), .A2(n11614), .ZN(n7467) );
  NAND2_X1 U9622 ( .A1(n7472), .A2(n7473), .ZN(n11616) );
  NAND3_X1 U9623 ( .A1(n11608), .A2(n6561), .A3(n11607), .ZN(n7472) );
  NAND2_X1 U9624 ( .A1(n7474), .A2(n7475), .ZN(n11603) );
  NAND3_X1 U9625 ( .A1(n11597), .A2(n6560), .A3(n11596), .ZN(n7474) );
  OAI21_X1 U9626 ( .B1(n11685), .B2(n7480), .A(n7479), .ZN(n11701) );
  NAND2_X1 U9627 ( .A1(n7476), .A2(n7477), .ZN(n11700) );
  NAND2_X1 U9628 ( .A1(n11685), .A2(n7479), .ZN(n7476) );
  NAND2_X1 U9629 ( .A1(n11628), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U9630 ( .A1(n7481), .A2(n7483), .ZN(n11657) );
  NAND2_X1 U9631 ( .A1(n7487), .A2(n7490), .ZN(n11760) );
  INV_X1 U9632 ( .A(n11744), .ZN(n7489) );
  NAND3_X1 U9633 ( .A1(n11586), .A2(n11585), .A3(n6506), .ZN(n7499) );
  NAND2_X1 U9634 ( .A1(n7499), .A2(n7500), .ZN(n11592) );
  NAND2_X1 U9635 ( .A1(n13726), .A2(n13727), .ZN(n7504) );
  NAND2_X1 U9636 ( .A1(n9116), .A2(n9212), .ZN(n9641) );
  OR2_X1 U9637 ( .A1(n11007), .A2(n11008), .ZN(n7522) );
  NAND2_X1 U9638 ( .A1(n11439), .A2(n7525), .ZN(n7524) );
  NAND2_X1 U9639 ( .A1(n7524), .A2(n7523), .ZN(n12020) );
  NAND2_X1 U9640 ( .A1(n11439), .A2(n11438), .ZN(n11440) );
  INV_X1 U9641 ( .A(n7524), .ZN(n11478) );
  NOR2_X1 U9642 ( .A1(n11441), .A2(n7526), .ZN(n7525) );
  INV_X1 U9643 ( .A(n11438), .ZN(n7526) );
  INV_X1 U9644 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9645 ( .A1(n13086), .A2(n11938), .ZN(n11939) );
  OAI21_X1 U9646 ( .B1(n11100), .B2(n11099), .A(n13019), .ZN(n11135) );
  OAI21_X2 U9647 ( .B1(n11288), .B2(n11287), .A(n11286), .ZN(n14790) );
  XNOR2_X1 U9648 ( .A(n11976), .B(n9053), .ZN(n10304) );
  CLKBUF_X1 U9649 ( .A(n12157), .Z(n12159) );
  XNOR2_X1 U9650 ( .A(n13997), .B(n6951), .ZN(n14002) );
  NOR2_X2 U9651 ( .A1(n13520), .A2(n13628), .ZN(n13498) );
  NAND2_X2 U9652 ( .A1(n11827), .A2(n11538), .ZN(n11574) );
  NAND2_X1 U9653 ( .A1(n8848), .A2(SI_22_), .ZN(n8849) );
  INV_X1 U9654 ( .A(n13922), .ZN(n14268) );
  OAI22_X1 U9655 ( .A1(n11847), .A2(n11846), .B1(n11852), .B2(n11851), .ZN(
        n11843) );
  AOI21_X2 U9656 ( .B1(n10309), .B2(n10308), .A(n10355), .ZN(n10485) );
  NAND2_X1 U9657 ( .A1(n11245), .A2(n11244), .ZN(n11417) );
  INV_X1 U9658 ( .A(n7557), .ZN(n10192) );
  INV_X1 U9659 ( .A(n8140), .ZN(n9789) );
  AOI21_X1 U9660 ( .B1(n11417), .B2(n11416), .A(n11415), .ZN(n11510) );
  INV_X1 U9661 ( .A(n10604), .ZN(n10609) );
  XNOR2_X1 U9662 ( .A(n8961), .B(n8960), .ZN(n13675) );
  NOR2_X1 U9663 ( .A1(n9224), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9157) );
  OAI22_X1 U9664 ( .A1(n10184), .A2(n9732), .B1(n14717), .B2(n12047), .ZN(
        n9625) );
  NAND2_X1 U9665 ( .A1(n6407), .A2(n6411), .ZN(n8371) );
  INV_X1 U9666 ( .A(n12933), .ZN(n8275) );
  OR2_X1 U9667 ( .A1(n15187), .A2(n15173), .ZN(n12981) );
  INV_X1 U9668 ( .A(n12981), .ZN(n8256) );
  AND2_X1 U9669 ( .A1(n8696), .A2(n8701), .ZN(n7536) );
  OR2_X1 U9670 ( .A1(n11629), .A2(n11867), .ZN(n7537) );
  OR2_X1 U9671 ( .A1(n15047), .A2(n11172), .ZN(n7539) );
  OR2_X1 U9672 ( .A1(n13646), .A2(n11511), .ZN(n7540) );
  AND3_X1 U9673 ( .A1(n11562), .A2(n11561), .A3(n11560), .ZN(n7542) );
  AND2_X1 U9674 ( .A1(n8749), .A2(n8730), .ZN(n7545) );
  NOR3_X1 U9675 ( .A1(n9769), .A2(n6427), .A3(n9094), .ZN(n7549) );
  NOR2_X1 U9676 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7550) );
  AND2_X1 U9677 ( .A1(n7744), .A2(n12516), .ZN(n7551) );
  INV_X1 U9678 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7560) );
  OR2_X1 U9679 ( .A1(n15185), .A2(n8257), .ZN(n7552) );
  AND2_X1 U9680 ( .A1(n8625), .A2(n8607), .ZN(n7553) );
  INV_X1 U9681 ( .A(n13316), .ZN(n13284) );
  AND2_X1 U9682 ( .A1(n8653), .A2(n8629), .ZN(n7554) );
  INV_X1 U9683 ( .A(n8225), .ZN(n12304) );
  INV_X1 U9684 ( .A(n11884), .ZN(n10593) );
  AND2_X1 U9685 ( .A1(n8726), .A2(n8706), .ZN(n7555) );
  INV_X1 U9686 ( .A(n12856), .ZN(n12829) );
  NAND2_X1 U9687 ( .A1(n8077), .A2(n8076), .ZN(n12736) );
  INV_X1 U9688 ( .A(n12736), .ZN(n12714) );
  INV_X1 U9689 ( .A(n12768), .ZN(n8007) );
  MUX2_X1 U9690 ( .A(n11540), .B(n11539), .S(n11574), .Z(n11551) );
  NAND2_X1 U9691 ( .A1(n6420), .A2(n9053), .ZN(n8355) );
  INV_X1 U9692 ( .A(n8384), .ZN(n8385) );
  INV_X1 U9693 ( .A(n8506), .ZN(n8507) );
  OAI21_X1 U9694 ( .B1(n11654), .B2(n11653), .A(n11652), .ZN(n11655) );
  INV_X1 U9695 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8285) );
  AND4_X1 U9696 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8561), .ZN(n8288)
         );
  NAND2_X1 U9697 ( .A1(n12955), .A2(n12714), .ZN(n8198) );
  NAND2_X1 U9698 ( .A1(n8028), .A2(n8027), .ZN(n8030) );
  INV_X1 U9699 ( .A(n14272), .ZN(n11899) );
  INV_X1 U9700 ( .A(n11624), .ZN(n11343) );
  INV_X1 U9701 ( .A(n12510), .ZN(n8026) );
  INV_X1 U9702 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9889) );
  INV_X1 U9703 ( .A(n12516), .ZN(n12385) );
  OR2_X1 U9704 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  INV_X1 U9705 ( .A(n10187), .ZN(n10188) );
  NAND2_X1 U9706 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  INV_X1 U9707 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10082) );
  INV_X1 U9708 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9270) );
  AOI21_X1 U9709 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(n8703) );
  NOR2_X1 U9710 ( .A1(n7710), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7736) );
  OR2_X1 U9711 ( .A1(n7761), .A2(n12515), .ZN(n7762) );
  INV_X1 U9712 ( .A(n12006), .ZN(n10808) );
  NOR2_X1 U9713 ( .A1(n8087), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8134) );
  OR2_X1 U9714 ( .A1(n8071), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U9715 ( .A1(n7898), .A2(n7897), .ZN(n7927) );
  NAND2_X1 U9716 ( .A1(n7829), .A2(n7828), .ZN(n7837) );
  INV_X1 U9717 ( .A(n15093), .ZN(n10890) );
  NOR2_X1 U9718 ( .A1(n12599), .A2(n12598), .ZN(n12605) );
  NAND2_X1 U9719 ( .A1(n12494), .A2(n12324), .ZN(n12323) );
  NOR2_X1 U9720 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7683) );
  INV_X1 U9721 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9722 ( .A1(n9147), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7678) );
  AND2_X1 U9723 ( .A1(n13038), .A2(n11934), .ZN(n11935) );
  OR2_X1 U9724 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  AND2_X1 U9725 ( .A1(n8965), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8982) );
  OR2_X1 U9726 ( .A1(n8658), .A2(n11299), .ZN(n8684) );
  NOR2_X1 U9727 ( .A1(n8515), .A2(n8514), .ZN(n8543) );
  NOR2_X1 U9728 ( .A1(n13292), .A2(n13291), .ZN(n13293) );
  AND2_X1 U9729 ( .A1(n14540), .A2(n14541), .ZN(n12031) );
  INV_X1 U9730 ( .A(n13719), .ZN(n12083) );
  INV_X1 U9731 ( .A(n11434), .ZN(n11437) );
  OR2_X1 U9732 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  INV_X1 U9733 ( .A(n14205), .ZN(n13921) );
  INV_X1 U9734 ( .A(n14097), .ZN(n14115) );
  INV_X1 U9735 ( .A(n14153), .ZN(n13920) );
  NAND2_X1 U9736 ( .A1(n8888), .A2(SI_24_), .ZN(n8889) );
  OR2_X1 U9737 ( .A1(n8808), .A2(n12015), .ZN(n8809) );
  NAND2_X1 U9738 ( .A1(n8534), .A2(n8533), .ZN(n8537) );
  NAND2_X1 U9739 ( .A1(n8450), .A2(n8449), .ZN(n8454) );
  INV_X1 U9740 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15224) );
  NAND2_X1 U9741 ( .A1(n14402), .A2(n14401), .ZN(n14347) );
  XNOR2_X1 U9742 ( .A(n7654), .B(n15161), .ZN(n7667) );
  NAND2_X1 U9743 ( .A1(n7981), .A2(n7980), .ZN(n8000) );
  NAND2_X1 U9744 ( .A1(n7667), .A2(n10856), .ZN(n7668) );
  OR2_X1 U9745 ( .A1(n7927), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7935) );
  OR2_X1 U9746 ( .A1(n7691), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7710) );
  OR2_X1 U9747 ( .A1(n12688), .A2(n8135), .ZN(n12705) );
  INV_X1 U9748 ( .A(n12873), .ZN(n15145) );
  NOR2_X1 U9749 ( .A1(n9788), .A2(n8130), .ZN(n12881) );
  INV_X1 U9750 ( .A(n15143), .ZN(n12875) );
  AND2_X1 U9751 ( .A1(n8241), .A2(n8270), .ZN(n12771) );
  INV_X1 U9752 ( .A(n12854), .ZN(n15149) );
  NAND2_X1 U9753 ( .A1(n7943), .A2(n7942), .ZN(n7946) );
  AND2_X1 U9754 ( .A1(n7821), .A2(n7800), .ZN(n7819) );
  OR2_X1 U9755 ( .A1(n8566), .A2(n8565), .ZN(n8591) );
  OR2_X1 U9756 ( .A1(n8684), .A2(n8683), .ZN(n8712) );
  INV_X1 U9757 ( .A(n14529), .ZN(n11924) );
  OR2_X1 U9758 ( .A1(n13087), .A2(n11937), .ZN(n11938) );
  AND2_X1 U9759 ( .A1(n13131), .A2(n13529), .ZN(n11497) );
  AND2_X1 U9760 ( .A1(n8832), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8853) );
  AND2_X1 U9761 ( .A1(n8814), .A2(n8813), .ZN(n8832) );
  AND2_X1 U9762 ( .A1(n14832), .A2(n14831), .ZN(n14834) );
  OR2_X1 U9763 ( .A1(n9973), .A2(n9972), .ZN(n13227) );
  INV_X1 U9764 ( .A(n13129), .ZN(n13511) );
  AND2_X1 U9765 ( .A1(n15054), .A2(n13135), .ZN(n11168) );
  AND2_X1 U9766 ( .A1(n9757), .A2(n6427), .ZN(n13254) );
  INV_X1 U9767 ( .A(n13024), .ZN(n15047) );
  OR2_X1 U9768 ( .A1(n14933), .A2(n9649), .ZN(n15059) );
  NAND2_X1 U9769 ( .A1(n11437), .A2(n11436), .ZN(n11438) );
  INV_X1 U9770 ( .A(n11871), .ZN(n11866) );
  AND2_X1 U9771 ( .A1(n11688), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11704) );
  AND2_X1 U9772 ( .A1(n9738), .A2(n9706), .ZN(n9707) );
  NAND2_X1 U9773 ( .A1(n13998), .A2(n14575), .ZN(n14001) );
  AND2_X1 U9774 ( .A1(n9260), .A2(n9259), .ZN(n9684) );
  NAND2_X1 U9775 ( .A1(n8602), .A2(n8585), .ZN(n8603) );
  AOI22_X1 U9776 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14342), .B1(n14395), .B2(
        n14341), .ZN(n14344) );
  OAI21_X1 U9777 ( .B1(n12951), .B2(n12278), .A(n8154), .ZN(n8155) );
  OR2_X1 U9778 ( .A1(n15151), .A2(n8132), .ZN(n12287) );
  AOI21_X1 U9779 ( .B1(n12705), .B2(n8090), .A(n8138), .ZN(n12715) );
  INV_X1 U9780 ( .A(n6457), .ZN(n8207) );
  AND4_X1 U9781 ( .A1(n7817), .A2(n7816), .A3(n7815), .A4(n7814), .ZN(n12246)
         );
  NAND2_X1 U9782 ( .A1(n8214), .A2(n12500), .ZN(n12854) );
  INV_X1 U9783 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10267) );
  INV_X1 U9784 ( .A(n12881), .ZN(n11405) );
  NAND2_X1 U9785 ( .A1(n8255), .A2(n8256), .ZN(n8258) );
  INV_X1 U9786 ( .A(n15184), .ZN(n15173) );
  AND2_X1 U9787 ( .A1(n12331), .A2(n8101), .ZN(n15184) );
  INV_X1 U9788 ( .A(n15179), .ZN(n15177) );
  OR2_X1 U9789 ( .A1(n8244), .A2(n8243), .ZN(n8254) );
  INV_X1 U9790 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7847) );
  AND2_X1 U9791 ( .A1(n9771), .A2(n9770), .ZN(n14534) );
  AND2_X1 U9792 ( .A1(n13112), .A2(n11966), .ZN(n11967) );
  INV_X1 U9793 ( .A(n14853), .ZN(n14917) );
  INV_X1 U9794 ( .A(n10303), .ZN(n13496) );
  INV_X1 U9795 ( .A(n13276), .ZN(n13457) );
  AND2_X1 U9796 ( .A1(n13543), .A2(n10369), .ZN(n13535) );
  AND2_X1 U9797 ( .A1(n9654), .A2(n9653), .ZN(n15057) );
  INV_X1 U9798 ( .A(n14999), .ZN(n15022) );
  INV_X1 U9799 ( .A(n15057), .ZN(n15026) );
  AOI21_X1 U9800 ( .B1(n9657), .B2(n11361), .A(n13689), .ZN(n14944) );
  AND2_X1 U9801 ( .A1(n9659), .A2(n9658), .ZN(n10365) );
  AND2_X1 U9802 ( .A1(n8496), .A2(n8538), .ZN(n9545) );
  OR2_X1 U9803 ( .A1(n9737), .A2(n9705), .ZN(n9738) );
  AND2_X1 U9804 ( .A1(n9686), .A2(n9685), .ZN(n13967) );
  AND2_X1 U9805 ( .A1(n9560), .A2(n9199), .ZN(n9580) );
  AND2_X1 U9806 ( .A1(n9794), .A2(n9793), .ZN(n15082) );
  INV_X1 U9807 ( .A(n12904), .ZN(n12759) );
  INV_X1 U9808 ( .A(n12287), .ZN(n12278) );
  INV_X1 U9809 ( .A(n15106), .ZN(n15122) );
  OR2_X1 U9810 ( .A1(n9838), .A2(n9837), .ZN(n15136) );
  OR2_X1 U9811 ( .A1(n9838), .A2(n9796), .ZN(n15125) );
  AND2_X1 U9812 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  INV_X1 U9813 ( .A(n15199), .ZN(n15196) );
  INV_X1 U9814 ( .A(n8238), .ZN(n12955) );
  AND2_X1 U9815 ( .A1(n8254), .A2(n8253), .ZN(n15187) );
  NAND2_X1 U9816 ( .A1(n9790), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12986) );
  AND2_X1 U9817 ( .A1(n9353), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14923) );
  OR2_X1 U9818 ( .A1(n8743), .A2(n8742), .ZN(n13129) );
  INV_X1 U9819 ( .A(n13535), .ZN(n13500) );
  INV_X1 U9820 ( .A(n13542), .ZN(n13524) );
  AND4_X1 U9821 ( .A1(n15035), .A2(n15034), .A3(n15033), .A4(n15032), .ZN(
        n15074) );
  INV_X1 U9822 ( .A(n15066), .ZN(n15065) );
  CLKBUF_X1 U9823 ( .A(n14969), .Z(n14973) );
  INV_X1 U9824 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9465) );
  INV_X1 U9825 ( .A(n13749), .ZN(n14591) );
  INV_X1 U9826 ( .A(n13986), .ZN(n14238) );
  INV_X1 U9827 ( .A(n14564), .ZN(n13821) );
  NAND2_X1 U9828 ( .A1(n13967), .A2(n9688), .ZN(n14763) );
  INV_X1 U9829 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11059) );
  AND3_X2 U9830 ( .A1(n7564), .A2(n7563), .A3(n7562), .ZN(n7801) );
  AND2_X2 U9831 ( .A1(n7881), .A2(n7550), .ZN(n7909) );
  INV_X1 U9832 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7566) );
  MUX2_X1 U9833 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7570), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7572) );
  NOR2_X1 U9834 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7575) );
  INV_X1 U9835 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7573) );
  NAND4_X1 U9836 ( .A1(n7575), .A2(n7574), .A3(n15324), .A4(n7573), .ZN(n7579)
         );
  INV_X1 U9837 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9838 ( .A1(n7597), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7580) );
  MUX2_X1 U9839 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7580), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7581) );
  OR2_X1 U9840 ( .A1(n7597), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7582) );
  AND2_X1 U9841 ( .A1(n7581), .A2(n7582), .ZN(n8126) );
  XNOR2_X1 U9842 ( .A(n11019), .B(P3_B_REG_SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9843 ( .A1(n7582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7583) );
  MUX2_X1 U9844 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7583), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7584) );
  AND2_X1 U9845 ( .A1(n7595), .A2(n7584), .ZN(n8125) );
  INV_X1 U9846 ( .A(n8125), .ZN(n11131) );
  NAND2_X1 U9847 ( .A1(n7595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7586) );
  XNOR2_X1 U9848 ( .A(n7586), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8127) );
  INV_X1 U9849 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n15345) );
  NAND2_X1 U9850 ( .A1(n6527), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7587) );
  NAND2_X1 U9851 ( .A1(n8101), .A2(n12687), .ZN(n7588) );
  NAND2_X1 U9852 ( .A1(n7588), .A2(n12014), .ZN(n7589) );
  NAND2_X1 U9853 ( .A1(n7591), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7592) );
  MUX2_X1 U9854 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7592), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7594) );
  INV_X1 U9855 ( .A(n7673), .ZN(n7593) );
  OAI21_X2 U9856 ( .B1(n7595), .B2(P3_IR_REG_26__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7596) );
  INV_X1 U9857 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7601) );
  INV_X1 U9858 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7600) );
  INV_X1 U9859 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U9860 ( .A1(n7603), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7602) );
  NAND2_X4 U9861 ( .A1(n6416), .A2(n8139), .ZN(n8140) );
  XNOR2_X1 U9862 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7628) );
  NAND2_X1 U9863 ( .A1(n7628), .A2(n7607), .ZN(n7609) );
  INV_X1 U9864 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U9865 ( .A1(n7651), .A2(n7650), .ZN(n7611) );
  XNOR2_X1 U9866 ( .A(n7677), .B(n7676), .ZN(n9173) );
  OR2_X1 U9867 ( .A1(n8068), .A2(n9173), .ZN(n7614) );
  OR2_X1 U9868 ( .A1(n12299), .A2(SI_4_), .ZN(n7613) );
  OAI211_X1 U9869 ( .C1(n9860), .C2(n8140), .A(n7614), .B(n7613), .ZN(n8170)
         );
  XNOR2_X1 U9870 ( .A(n7851), .B(n8170), .ZN(n7669) );
  INV_X1 U9871 ( .A(n7669), .ZN(n7670) );
  INV_X2 U9872 ( .A(n8057), .ZN(n8215) );
  NAND2_X1 U9873 ( .A1(n8215), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7624) );
  INV_X1 U9874 ( .A(n7683), .ZN(n7684) );
  NAND2_X1 U9875 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7618) );
  NAND2_X1 U9876 ( .A1(n7684), .A2(n7618), .ZN(n10860) );
  NAND2_X1 U9877 ( .A1(n7634), .A2(n10860), .ZN(n7623) );
  NAND2_X1 U9878 ( .A1(n6457), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9879 ( .A1(n7657), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7621) );
  NAND4_X1 U9880 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n12520)
         );
  INV_X1 U9881 ( .A(n12520), .ZN(n10641) );
  INV_X1 U9882 ( .A(SI_1_), .ZN(n9150) );
  OR2_X1 U9883 ( .A1(n12299), .A2(n9150), .ZN(n7630) );
  XNOR2_X1 U9884 ( .A(n7640), .B(n7628), .ZN(n9151) );
  INV_X1 U9885 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15160) );
  OR2_X1 U9886 ( .A1(n8057), .A2(n15160), .ZN(n7632) );
  NAND2_X1 U9887 ( .A1(n7634), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U9888 ( .A1(n7633), .A2(n6689), .ZN(n7643) );
  NAND2_X1 U9889 ( .A1(n7634), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9890 ( .A1(n6457), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7637) );
  INV_X1 U9891 ( .A(n8057), .ZN(n7890) );
  NAND2_X1 U9892 ( .A1(n8215), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9893 ( .A1(n7657), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9894 ( .A1(n8376), .A2(SI_0_), .ZN(n9144) );
  MUX2_X1 U9895 ( .A(n15268), .B(n9144), .S(n8140), .Z(n7642) );
  INV_X1 U9896 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U9897 ( .A1(n9267), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7639) );
  AND2_X1 U9898 ( .A1(n7640), .A2(n7639), .ZN(n9146) );
  OR2_X1 U9899 ( .A1(n8068), .A2(n9146), .ZN(n7641) );
  NAND2_X1 U9900 ( .A1(n7642), .A2(n7641), .ZN(n10380) );
  NAND2_X1 U9901 ( .A1(n9869), .A2(n10380), .ZN(n15140) );
  NAND2_X1 U9902 ( .A1(n7851), .A2(n15140), .ZN(n10806) );
  NAND4_X1 U9903 ( .A1(n10810), .A2(n7643), .A3(n15139), .A4(n10806), .ZN(
        n10805) );
  NAND2_X1 U9904 ( .A1(n10805), .A2(n10810), .ZN(n10646) );
  NAND2_X1 U9905 ( .A1(n7890), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U9906 ( .A1(n6457), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7644) );
  NOR2_X1 U9907 ( .A1(n7646), .A2(n12990), .ZN(n7647) );
  XNOR2_X1 U9908 ( .A(n7651), .B(n7650), .ZN(n9165) );
  OR2_X1 U9909 ( .A1(n8068), .A2(n9165), .ZN(n7653) );
  OAI211_X1 U9910 ( .C1(n10005), .C2(n8140), .A(n7653), .B(n7652), .ZN(n8167)
         );
  XOR2_X1 U9911 ( .A(n15144), .B(n7655), .Z(n10647) );
  INV_X1 U9912 ( .A(n7655), .ZN(n7656) );
  NAND2_X1 U9913 ( .A1(n7890), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7661) );
  INV_X1 U9914 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U9915 ( .A1(n7634), .A2(n10532), .ZN(n7660) );
  NAND2_X1 U9916 ( .A1(n6457), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U9917 ( .A1(n7657), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7658) );
  XNOR2_X1 U9918 ( .A(n7662), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9814) );
  XNOR2_X1 U9919 ( .A(n7664), .B(n7663), .ZN(n9169) );
  OR2_X1 U9920 ( .A1(n8068), .A2(n9169), .ZN(n7666) );
  OR2_X1 U9921 ( .A1(n12299), .A2(SI_3_), .ZN(n7665) );
  OAI211_X1 U9922 ( .C1(n9814), .C2(n8140), .A(n7666), .B(n7665), .ZN(n15161)
         );
  XOR2_X1 U9923 ( .A(n10856), .B(n7667), .Z(n10525) );
  INV_X1 U9924 ( .A(n10856), .ZN(n10631) );
  XNOR2_X1 U9925 ( .A(n7669), .B(n12520), .ZN(n10627) );
  NOR2_X1 U9926 ( .A1(n7673), .A2(n12990), .ZN(n7671) );
  MUX2_X1 U9927 ( .A(n12990), .B(n7671), .S(P3_IR_REG_5__SCAN_IN), .Z(n7675)
         );
  INV_X1 U9928 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9929 ( .A1(n7673), .A2(n7672), .ZN(n7803) );
  INV_X1 U9930 ( .A(n7803), .ZN(n7674) );
  XNOR2_X1 U9931 ( .A(n7700), .B(n7699), .ZN(n9171) );
  OR2_X1 U9932 ( .A1(n8068), .A2(n9171), .ZN(n7681) );
  OR2_X1 U9933 ( .A1(n12299), .A2(SI_5_), .ZN(n7680) );
  OAI211_X1 U9934 ( .C1(n9831), .C2(n8140), .A(n7681), .B(n7680), .ZN(n10222)
         );
  XNOR2_X1 U9935 ( .A(n7851), .B(n10222), .ZN(n7690) );
  NAND2_X1 U9936 ( .A1(n8215), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9937 ( .A1(n7684), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9938 ( .A1(n7691), .A2(n7685), .ZN(n10643) );
  NAND2_X1 U9939 ( .A1(n8090), .A2(n10643), .ZN(n7688) );
  NAND2_X1 U9940 ( .A1(n6457), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9941 ( .A1(n7657), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7686) );
  NAND4_X1 U9942 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .ZN(n12519)
         );
  XNOR2_X1 U9943 ( .A(n7690), .B(n12519), .ZN(n10636) );
  OAI22_X1 U9944 ( .A1(n10635), .A2(n10636), .B1(n7690), .B2(n12519), .ZN(
        n10472) );
  INV_X1 U9945 ( .A(n10472), .ZN(n7706) );
  NAND2_X1 U9946 ( .A1(n8215), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9947 ( .A1(n7691), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9948 ( .A1(n7710), .A2(n7692), .ZN(n10478) );
  NAND2_X1 U9949 ( .A1(n8090), .A2(n10478), .ZN(n7695) );
  NAND2_X1 U9950 ( .A1(n6457), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U9951 ( .A1(n8216), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7693) );
  NAND4_X1 U9952 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7693), .ZN(n12518)
         );
  NAND2_X1 U9953 ( .A1(n7803), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7698) );
  INV_X1 U9954 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7697) );
  XNOR2_X1 U9955 ( .A(n7698), .B(n7697), .ZN(n10004) );
  NAND2_X1 U9956 ( .A1(n9164), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U9957 ( .A(n9179), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U9958 ( .A(n7717), .B(n7702), .ZN(n9154) );
  OR2_X1 U9959 ( .A1(n8068), .A2(n9154), .ZN(n7704) );
  INV_X1 U9960 ( .A(SI_6_), .ZN(n9153) );
  OR2_X1 U9961 ( .A1(n12299), .A2(n9153), .ZN(n7703) );
  OAI211_X1 U9962 ( .C1(n8140), .C2(n10004), .A(n7704), .B(n7703), .ZN(n10468)
         );
  XNOR2_X1 U9963 ( .A(n7851), .B(n10468), .ZN(n7707) );
  XOR2_X1 U9964 ( .A(n12518), .B(n7707), .Z(n10475) );
  INV_X1 U9965 ( .A(n10475), .ZN(n7705) );
  NAND2_X1 U9966 ( .A1(n7706), .A2(n7705), .ZN(n10473) );
  INV_X1 U9967 ( .A(n7707), .ZN(n7708) );
  NAND2_X1 U9968 ( .A1(n12518), .A2(n7708), .ZN(n7709) );
  NAND2_X1 U9969 ( .A1(n10473), .A2(n7709), .ZN(n10432) );
  INV_X1 U9970 ( .A(n7736), .ZN(n7737) );
  NAND2_X1 U9971 ( .A1(n7710), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U9972 ( .A1(n7737), .A2(n7711), .ZN(n10687) );
  NAND2_X1 U9973 ( .A1(n8090), .A2(n10687), .ZN(n7715) );
  NAND2_X1 U9974 ( .A1(n6457), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U9975 ( .A1(n8215), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9976 ( .A1(n8216), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7712) );
  XNOR2_X1 U9977 ( .A(n7731), .B(n7729), .ZN(n9167) );
  OR2_X1 U9978 ( .A1(n8068), .A2(n9167), .ZN(n7722) );
  OR2_X1 U9979 ( .A1(n12299), .A2(SI_7_), .ZN(n7721) );
  NAND2_X1 U9980 ( .A1(n7724), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7719) );
  INV_X1 U9981 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7718) );
  XNOR2_X1 U9982 ( .A(n7719), .B(n7718), .ZN(n9883) );
  INV_X1 U9983 ( .A(n9883), .ZN(n9894) );
  OR2_X1 U9984 ( .A1(n8140), .A2(n9894), .ZN(n7720) );
  NAND2_X1 U9985 ( .A1(n10758), .A2(n10434), .ZN(n12377) );
  INV_X1 U9986 ( .A(n10434), .ZN(n10689) );
  NAND2_X1 U9987 ( .A1(n12517), .A2(n10689), .ZN(n12376) );
  XNOR2_X1 U9988 ( .A(n12373), .B(n7851), .ZN(n10431) );
  NOR2_X1 U9989 ( .A1(n7724), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7727) );
  OR2_X1 U9990 ( .A1(n7727), .A2(n12990), .ZN(n7725) );
  INV_X1 U9991 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7726) );
  MUX2_X1 U9992 ( .A(n7725), .B(P3_IR_REG_31__SCAN_IN), .S(n7726), .Z(n7728)
         );
  NAND2_X1 U9993 ( .A1(n7727), .A2(n7726), .ZN(n7766) );
  NAND2_X1 U9994 ( .A1(n7728), .A2(n7766), .ZN(n10335) );
  NAND2_X1 U9995 ( .A1(n9183), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U9996 ( .A(n7754), .B(n7753), .ZN(n9148) );
  OR2_X1 U9997 ( .A1(n8068), .A2(n9148), .ZN(n7735) );
  INV_X1 U9998 ( .A(SI_8_), .ZN(n9149) );
  OR2_X1 U9999 ( .A1(n12299), .A2(n9149), .ZN(n7734) );
  XNOR2_X1 U10000 ( .A(n7851), .B(n12384), .ZN(n7743) );
  NAND2_X1 U10001 ( .A1(n8215), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7742) );
  INV_X1 U10002 ( .A(n7746), .ZN(n7747) );
  NAND2_X1 U10003 ( .A1(n7737), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10004 ( .A1(n7747), .A2(n7738), .ZN(n10761) );
  NAND2_X1 U10005 ( .A1(n8090), .A2(n10761), .ZN(n7741) );
  NAND2_X1 U10006 ( .A1(n6457), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10007 ( .A1(n8216), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7739) );
  XNOR2_X1 U10008 ( .A(n7743), .B(n12516), .ZN(n10676) );
  INV_X1 U10009 ( .A(n7743), .ZN(n7744) );
  NAND2_X1 U10010 ( .A1(n8216), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U10011 ( .A1(n6457), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7751) );
  INV_X1 U10012 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10013 ( .A1(n7747), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10014 ( .A1(n7771), .A2(n7748), .ZN(n10847) );
  NAND2_X1 U10015 ( .A1(n8090), .A2(n10847), .ZN(n7750) );
  NAND2_X1 U10016 ( .A1(n8215), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7749) );
  INV_X1 U10017 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10018 ( .A1(n7755), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7756) );
  XNOR2_X1 U10019 ( .A(n7764), .B(n7763), .ZN(n14440) );
  NAND2_X1 U10020 ( .A1(n14440), .A2(n12296), .ZN(n7760) );
  NAND2_X1 U10021 ( .A1(n7766), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7758) );
  INV_X1 U10022 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7757) );
  XNOR2_X1 U10023 ( .A(n7758), .B(n7757), .ZN(n14443) );
  OR2_X1 U10024 ( .A1(n8140), .A2(n10910), .ZN(n7759) );
  XNOR2_X1 U10025 ( .A(n7851), .B(n12391), .ZN(n7761) );
  XOR2_X1 U10026 ( .A(n12515), .B(n7761), .Z(n10997) );
  NAND2_X1 U10027 ( .A1(n9197), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7765) );
  XNOR2_X1 U10028 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7780) );
  XNOR2_X1 U10029 ( .A(n7781), .B(n7780), .ZN(n9155) );
  NAND2_X1 U10030 ( .A1(n9155), .A2(n12296), .ZN(n7770) );
  INV_X1 U10031 ( .A(SI_10_), .ZN(n9156) );
  OR2_X1 U10032 ( .A1(n7766), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U10033 ( .A1(n7785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7768) );
  INV_X1 U10034 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7767) );
  XNOR2_X1 U10035 ( .A(n7768), .B(n7767), .ZN(n15095) );
  AOI22_X1 U10036 ( .A1(n7948), .A2(n9156), .B1(n9789), .B2(n15095), .ZN(n7769) );
  NAND2_X1 U10037 ( .A1(n7770), .A2(n7769), .ZN(n8178) );
  XNOR2_X1 U10038 ( .A(n7851), .B(n8178), .ZN(n7777) );
  NAND2_X1 U10039 ( .A1(n8215), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10040 ( .A1(n7771), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10041 ( .A1(n7790), .A2(n7772), .ZN(n11200) );
  NAND2_X1 U10042 ( .A1(n8090), .A2(n11200), .ZN(n7775) );
  NAND2_X1 U10043 ( .A1(n6457), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10044 ( .A1(n8216), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7773) );
  NAND4_X1 U10045 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n12514) );
  XNOR2_X1 U10046 ( .A(n7777), .B(n12514), .ZN(n11208) );
  INV_X1 U10047 ( .A(n7777), .ZN(n7778) );
  INV_X1 U10048 ( .A(n12514), .ZN(n11455) );
  NOR2_X1 U10049 ( .A1(n7778), .A2(n11455), .ZN(n7779) );
  INV_X1 U10050 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U10051 ( .A1(n7782), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7783) );
  XNOR2_X1 U10052 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7784) );
  XNOR2_X1 U10053 ( .A(n7799), .B(n7784), .ZN(n14444) );
  NAND2_X1 U10054 ( .A1(n14444), .A2(n12296), .ZN(n7789) );
  INV_X1 U10055 ( .A(SI_11_), .ZN(n8582) );
  OAI21_X1 U10056 ( .B1(n7785), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7787) );
  INV_X1 U10057 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7786) );
  XNOR2_X1 U10058 ( .A(n7787), .B(n7786), .ZN(n14449) );
  AOI22_X1 U10059 ( .A1(n7948), .A2(n8582), .B1(n9789), .B2(n14449), .ZN(n7788) );
  NAND2_X1 U10060 ( .A1(n7789), .A2(n7788), .ZN(n14513) );
  XOR2_X1 U10061 ( .A(n14513), .B(n7851), .Z(n7796) );
  NAND2_X1 U10062 ( .A1(n7790), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10063 ( .A1(n7812), .A2(n7791), .ZN(n11451) );
  NAND2_X1 U10064 ( .A1(n8090), .A2(n11451), .ZN(n7795) );
  NAND2_X1 U10065 ( .A1(n6457), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10066 ( .A1(n8216), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U10067 ( .A1(n8215), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7792) );
  AND2_X1 U10068 ( .A1(n9216), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10069 ( .A1(n9380), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10070 ( .A1(n9383), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U10071 ( .A(n7820), .B(n7819), .ZN(n9189) );
  NAND2_X1 U10072 ( .A1(n9189), .A2(n12296), .ZN(n7810) );
  INV_X1 U10073 ( .A(n7801), .ZN(n7802) );
  OAI21_X1 U10074 ( .B1(n7803), .B2(n7802), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7804) );
  MUX2_X1 U10075 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7804), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7808) );
  INV_X1 U10076 ( .A(n7806), .ZN(n7807) );
  NAND2_X1 U10077 ( .A1(n7808), .A2(n7807), .ZN(n15123) );
  INV_X1 U10078 ( .A(n15123), .ZN(n11312) );
  AOI22_X1 U10079 ( .A1(n7948), .A2(SI_12_), .B1(n9789), .B2(n11312), .ZN(
        n7809) );
  NAND2_X1 U10080 ( .A1(n7810), .A2(n7809), .ZN(n14512) );
  XNOR2_X1 U10081 ( .A(n14512), .B(n12006), .ZN(n12182) );
  INV_X1 U10082 ( .A(n7829), .ZN(n7830) );
  NAND2_X1 U10083 ( .A1(n7812), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10084 ( .A1(n7830), .A2(n7813), .ZN(n12177) );
  NAND2_X1 U10085 ( .A1(n8090), .A2(n12177), .ZN(n7817) );
  NAND2_X1 U10086 ( .A1(n6457), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10087 ( .A1(n8216), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10088 ( .A1(n8215), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10089 ( .A1(n12182), .A2(n12246), .ZN(n7818) );
  XNOR2_X1 U10090 ( .A(n7843), .B(n9465), .ZN(n14452) );
  NAND2_X1 U10091 ( .A1(n14452), .A2(n12296), .ZN(n7826) );
  INV_X1 U10092 ( .A(SI_13_), .ZN(n14450) );
  OR2_X1 U10093 ( .A1(n7806), .A2(n12990), .ZN(n7824) );
  XNOR2_X1 U10094 ( .A(n7824), .B(n7337), .ZN(n14455) );
  AOI22_X1 U10095 ( .A1(n7948), .A2(n14450), .B1(n9789), .B2(n14455), .ZN(
        n7825) );
  XNOR2_X1 U10096 ( .A(n14504), .B(n12006), .ZN(n7836) );
  NAND2_X1 U10097 ( .A1(n8216), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10098 ( .A1(n6457), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7834) );
  INV_X1 U10099 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U10100 ( .A1(n7830), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10101 ( .A1(n7837), .A2(n7831), .ZN(n12242) );
  NAND2_X1 U10102 ( .A1(n8090), .A2(n12242), .ZN(n7833) );
  NAND2_X1 U10103 ( .A1(n8215), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7832) );
  NAND4_X1 U10104 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n12512) );
  XNOR2_X1 U10105 ( .A(n7836), .B(n12512), .ZN(n12240) );
  INV_X1 U10106 ( .A(n12512), .ZN(n11468) );
  NAND2_X1 U10107 ( .A1(n7657), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10108 ( .A1(n6457), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U10109 ( .A1(n7837), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10110 ( .A1(n7866), .A2(n7838), .ZN(n11471) );
  NAND2_X1 U10111 ( .A1(n8090), .A2(n11471), .ZN(n7840) );
  NAND2_X1 U10112 ( .A1(n7890), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7839) );
  NAND4_X1 U10113 ( .A1(n7842), .A2(n7841), .A3(n7840), .A4(n7839), .ZN(n12511) );
  INV_X1 U10114 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U10115 ( .A1(n9679), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7853) );
  INV_X1 U10116 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U10117 ( .A1(n9681), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7845) );
  AND2_X1 U10118 ( .A1(n7853), .A2(n7845), .ZN(n7855) );
  XNOR2_X1 U10119 ( .A(n7856), .B(n7855), .ZN(n9218) );
  NAND2_X1 U10120 ( .A1(n9218), .A2(n12296), .ZN(n7850) );
  INV_X1 U10121 ( .A(SI_14_), .ZN(n9217) );
  OR2_X1 U10122 ( .A1(n7846), .A2(n12990), .ZN(n7848) );
  XNOR2_X1 U10123 ( .A(n7848), .B(n7847), .ZN(n12530) );
  AOI22_X1 U10124 ( .A1(n7948), .A2(n9217), .B1(n9789), .B2(n12530), .ZN(n7849) );
  XNOR2_X1 U10125 ( .A(n14499), .B(n7851), .ZN(n7852) );
  XOR2_X1 U10126 ( .A(n12511), .B(n7852), .Z(n11465) );
  INV_X1 U10127 ( .A(n12511), .ZN(n12874) );
  INV_X1 U10128 ( .A(n7853), .ZN(n7854) );
  INV_X1 U10129 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U10130 ( .A1(n11338), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7875) );
  INV_X1 U10131 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U10132 ( .A1(n9713), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U10133 ( .A1(n7875), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10134 ( .A1(n7858), .A2(n7859), .ZN(n7861) );
  INV_X1 U10135 ( .A(n7859), .ZN(n7860) );
  NAND2_X1 U10136 ( .A1(n7861), .A2(n7876), .ZN(n9399) );
  NAND2_X1 U10137 ( .A1(n7862), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7863) );
  XNOR2_X1 U10138 ( .A(n7863), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U10139 ( .A1(n7948), .A2(SI_15_), .B1(n9789), .B2(n12597), .ZN(
        n7864) );
  XNOR2_X1 U10140 ( .A(n12879), .B(n12006), .ZN(n7872) );
  INV_X1 U10141 ( .A(n7887), .ZN(n7888) );
  NAND2_X1 U10142 ( .A1(n7866), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10143 ( .A1(n7888), .A2(n7867), .ZN(n12880) );
  NAND2_X1 U10144 ( .A1(n12880), .A2(n8090), .ZN(n7871) );
  NAND2_X1 U10145 ( .A1(n7890), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10146 ( .A1(n6457), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10147 ( .A1(n7657), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7868) );
  NAND4_X1 U10148 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n12855) );
  XNOR2_X1 U10149 ( .A(n7872), .B(n12855), .ZN(n12280) );
  INV_X1 U10150 ( .A(n7872), .ZN(n7873) );
  NAND2_X1 U10151 ( .A1(n7873), .A2(n12855), .ZN(n7874) );
  INV_X1 U10152 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U10153 ( .A1(n9646), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7903) );
  INV_X1 U10154 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U10155 ( .A1(n9648), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7877) );
  AND2_X1 U10156 ( .A1(n7903), .A2(n7877), .ZN(n7878) );
  OR2_X1 U10157 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U10158 ( .A1(n7904), .A2(n7880), .ZN(n9503) );
  INV_X1 U10159 ( .A(n7881), .ZN(n7883) );
  NAND2_X1 U10160 ( .A1(n7883), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7882) );
  MUX2_X1 U10161 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7882), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n7884) );
  OR2_X1 U10162 ( .A1(n7883), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7906) );
  AND2_X1 U10163 ( .A1(n7884), .A2(n7906), .ZN(n12602) );
  AOI22_X1 U10164 ( .A1(n7948), .A2(SI_16_), .B1(n9789), .B2(n12602), .ZN(
        n7885) );
  XNOR2_X1 U10165 ( .A(n12938), .B(n12006), .ZN(n7895) );
  INV_X1 U10166 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12589) );
  INV_X1 U10167 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12203) );
  INV_X1 U10168 ( .A(n7898), .ZN(n7899) );
  NAND2_X1 U10169 ( .A1(n7888), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10170 ( .A1(n7899), .A2(n7889), .ZN(n12864) );
  NAND2_X1 U10171 ( .A1(n12864), .A2(n8090), .ZN(n7894) );
  NAND2_X1 U10172 ( .A1(n7890), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10173 ( .A1(n7657), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7891) );
  AND2_X1 U10174 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  OAI211_X1 U10175 ( .C1(n8207), .C2(n12589), .A(n7894), .B(n7893), .ZN(n12839) );
  XNOR2_X1 U10176 ( .A(n7895), .B(n12839), .ZN(n12202) );
  INV_X1 U10177 ( .A(n7895), .ZN(n7896) );
  INV_X1 U10178 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12615) );
  INV_X1 U10179 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10180 ( .A1(n7899), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10181 ( .A1(n7927), .A2(n7900), .ZN(n12846) );
  NAND2_X1 U10182 ( .A1(n12846), .A2(n8090), .ZN(n7902) );
  AOI22_X1 U10183 ( .A1(n8215), .A2(P3_REG0_REG_17__SCAN_IN), .B1(n8216), .B2(
        P3_REG2_REG_17__SCAN_IN), .ZN(n7901) );
  OAI211_X1 U10184 ( .C1(n8207), .C2(n12615), .A(n7902), .B(n7901), .ZN(n12856) );
  INV_X1 U10185 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U10186 ( .A1(n9721), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7918) );
  INV_X1 U10187 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U10188 ( .A1(n9722), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10189 ( .A1(n7918), .A2(n7905), .ZN(n7915) );
  XNOR2_X1 U10190 ( .A(n7917), .B(n7915), .ZN(n9635) );
  NAND2_X1 U10191 ( .A1(n9635), .A2(n12296), .ZN(n7912) );
  NAND2_X1 U10192 ( .A1(n7906), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7907) );
  MUX2_X1 U10193 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7907), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7908) );
  INV_X1 U10194 ( .A(n7908), .ZN(n7910) );
  NOR2_X1 U10195 ( .A1(n7910), .A2(n7909), .ZN(n12641) );
  AOI22_X1 U10196 ( .A1(n7948), .A2(SI_17_), .B1(n9789), .B2(n12641), .ZN(
        n7911) );
  XNOR2_X1 U10197 ( .A(n12934), .B(n12006), .ZN(n7913) );
  XOR2_X1 U10198 ( .A(n12856), .B(n7913), .Z(n12213) );
  NAND2_X1 U10199 ( .A1(n7913), .A2(n12829), .ZN(n7914) );
  INV_X1 U10200 ( .A(n7915), .ZN(n7916) );
  INV_X1 U10201 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U10202 ( .A1(n10063), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7942) );
  INV_X1 U10203 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U10204 ( .A1(n10060), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7919) );
  AND2_X1 U10205 ( .A1(n7942), .A2(n7919), .ZN(n7920) );
  OR2_X1 U10206 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  NAND2_X1 U10207 ( .A1(n7943), .A2(n7922), .ZN(n9682) );
  INV_X1 U10208 ( .A(n7909), .ZN(n7923) );
  NAND2_X1 U10209 ( .A1(n7923), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7924) );
  XNOR2_X1 U10210 ( .A(n7924), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U10211 ( .A1(n7948), .A2(SI_18_), .B1(n9789), .B2(n12668), .ZN(
        n7925) );
  XNOR2_X1 U10212 ( .A(n8190), .B(n12006), .ZN(n7932) );
  NAND2_X1 U10213 ( .A1(n7927), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U10214 ( .A1(n7935), .A2(n7928), .ZN(n12831) );
  INV_X1 U10215 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n15280) );
  NAND2_X1 U10216 ( .A1(n8215), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10217 ( .A1(n8216), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7929) );
  OAI211_X1 U10218 ( .C1(n15280), .C2(n8207), .A(n7930), .B(n7929), .ZN(n7931)
         );
  AOI21_X1 U10219 ( .B1(n12831), .B2(n8090), .A(n7931), .ZN(n8191) );
  XNOR2_X1 U10220 ( .A(n7932), .B(n8191), .ZN(n12260) );
  INV_X1 U10221 ( .A(n7932), .ZN(n7933) );
  INV_X1 U10222 ( .A(n8191), .ZN(n12840) );
  NAND2_X1 U10223 ( .A1(n7933), .A2(n12840), .ZN(n7934) );
  INV_X1 U10224 ( .A(n7963), .ZN(n7964) );
  NAND2_X1 U10225 ( .A1(n7935), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10226 ( .A1(n7964), .A2(n7936), .ZN(n12819) );
  NAND2_X1 U10227 ( .A1(n12819), .A2(n8090), .ZN(n7941) );
  INV_X1 U10228 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12928) );
  NAND2_X1 U10229 ( .A1(n8215), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10230 ( .A1(n8216), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7937) );
  OAI211_X1 U10231 ( .C1(n12928), .C2(n8207), .A(n7938), .B(n7937), .ZN(n7939)
         );
  INV_X1 U10232 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U10233 ( .A1(n7941), .A2(n7940), .ZN(n12800) );
  INV_X1 U10234 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U10235 ( .A1(n10210), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7954) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n15215) );
  NAND2_X1 U10237 ( .A1(n15215), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7944) );
  AND2_X1 U10238 ( .A1(n7954), .A2(n7944), .ZN(n7945) );
  OR2_X1 U10239 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NAND2_X1 U10240 ( .A1(n7955), .A2(n7947), .ZN(n9751) );
  NAND2_X1 U10241 ( .A1(n9751), .A2(n12296), .ZN(n7950) );
  INV_X1 U10242 ( .A(SI_19_), .ZN(n9750) );
  AOI22_X1 U10243 ( .A1(n7948), .A2(n9750), .B1(n12499), .B2(n9789), .ZN(n7949) );
  XNOR2_X1 U10244 ( .A(n12977), .B(n12006), .ZN(n7951) );
  XOR2_X1 U10245 ( .A(n12800), .B(n7951), .Z(n12158) );
  NAND2_X1 U10246 ( .A1(n7951), .A2(n12800), .ZN(n7952) );
  NAND2_X1 U10247 ( .A1(n7958), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10248 ( .A1(n7973), .A2(n7959), .ZN(n12016) );
  INV_X1 U10249 ( .A(SI_20_), .ZN(n12015) );
  OR2_X1 U10250 ( .A1(n12299), .A2(n12015), .ZN(n7960) );
  XNOR2_X1 U10251 ( .A(n12237), .B(n12006), .ZN(n7971) );
  INV_X1 U10252 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7962) );
  INV_X1 U10253 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U10254 ( .A1(n7964), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10255 ( .A1(n7982), .A2(n7965), .ZN(n12808) );
  NAND2_X1 U10256 ( .A1(n12808), .A2(n8090), .ZN(n7970) );
  INV_X1 U10257 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12924) );
  NAND2_X1 U10258 ( .A1(n7890), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10259 ( .A1(n8216), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7966) );
  OAI211_X1 U10260 ( .C1(n12924), .C2(n8207), .A(n7967), .B(n7966), .ZN(n7968)
         );
  INV_X1 U10261 ( .A(n7968), .ZN(n7969) );
  OAI21_X1 U10262 ( .B1(n7971), .B2(n12816), .A(n12167), .ZN(n12233) );
  INV_X1 U10263 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U10264 ( .A1(n11696), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7992) );
  INV_X1 U10265 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U10266 ( .A1(n15225), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7974) );
  AND2_X1 U10267 ( .A1(n7992), .A2(n7974), .ZN(n7975) );
  OR2_X1 U10268 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NAND2_X1 U10269 ( .A1(n7993), .A2(n7977), .ZN(n10249) );
  INV_X1 U10270 ( .A(SI_21_), .ZN(n10248) );
  OR2_X1 U10271 ( .A1(n12299), .A2(n10248), .ZN(n7978) );
  XNOR2_X1 U10272 ( .A(n12453), .B(n12006), .ZN(n7990) );
  INV_X1 U10273 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10274 ( .A1(n7982), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10275 ( .A1(n8000), .A2(n7983), .ZN(n12793) );
  NAND2_X1 U10276 ( .A1(n12793), .A2(n8090), .ZN(n7988) );
  INV_X1 U10277 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U10278 ( .A1(n7890), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10279 ( .A1(n8216), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7984) );
  OAI211_X1 U10280 ( .C1(n12918), .C2(n8207), .A(n7985), .B(n7984), .ZN(n7986)
         );
  INV_X1 U10281 ( .A(n7986), .ZN(n7987) );
  NAND2_X1 U10282 ( .A1(n7988), .A2(n7987), .ZN(n12801) );
  XNOR2_X1 U10283 ( .A(n7990), .B(n12801), .ZN(n12168) );
  NAND2_X1 U10284 ( .A1(n7989), .A2(n12168), .ZN(n12170) );
  INV_X1 U10285 ( .A(n12801), .ZN(n12781) );
  NAND2_X1 U10286 ( .A1(n7990), .A2(n12781), .ZN(n7991) );
  NAND2_X1 U10287 ( .A1(n12170), .A2(n7991), .ZN(n7999) );
  INV_X1 U10288 ( .A(n7999), .ZN(n7997) );
  INV_X1 U10289 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10948) );
  XNOR2_X1 U10290 ( .A(n10948), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8010) );
  XNOR2_X1 U10291 ( .A(n8011), .B(n8010), .ZN(n10361) );
  NAND2_X1 U10292 ( .A1(n10361), .A2(n12296), .ZN(n7995) );
  OR2_X1 U10293 ( .A1(n12299), .A2(n7371), .ZN(n7994) );
  XNOR2_X1 U10294 ( .A(n12257), .B(n12006), .ZN(n7998) );
  INV_X1 U10295 ( .A(n7998), .ZN(n7996) );
  NAND2_X1 U10296 ( .A1(n8000), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10297 ( .A1(n8019), .A2(n8001), .ZN(n12784) );
  NAND2_X1 U10298 ( .A1(n12784), .A2(n8090), .ZN(n8006) );
  INV_X1 U10299 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U10300 ( .A1(n8215), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10301 ( .A1(n8216), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8002) );
  OAI211_X1 U10302 ( .C1(n12914), .C2(n8207), .A(n8003), .B(n8002), .ZN(n8004)
         );
  INV_X1 U10303 ( .A(n8004), .ZN(n8005) );
  NAND2_X1 U10304 ( .A1(n8006), .A2(n8005), .ZN(n12768) );
  INV_X1 U10305 ( .A(n8017), .ZN(n8015) );
  NAND2_X1 U10306 ( .A1(n10948), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8009) );
  XNOR2_X1 U10307 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8027) );
  XNOR2_X1 U10308 ( .A(n8028), .B(n8027), .ZN(n10711) );
  NAND2_X1 U10309 ( .A1(n10711), .A2(n12296), .ZN(n8013) );
  INV_X1 U10310 ( .A(SI_23_), .ZN(n10713) );
  OR2_X1 U10311 ( .A1(n12299), .A2(n10713), .ZN(n8012) );
  XNOR2_X1 U10312 ( .A(n12330), .B(n12006), .ZN(n8016) );
  INV_X1 U10313 ( .A(n8016), .ZN(n8014) );
  NAND2_X1 U10314 ( .A1(n8019), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10315 ( .A1(n8035), .A2(n8020), .ZN(n12773) );
  NAND2_X1 U10316 ( .A1(n12773), .A2(n8090), .ZN(n8025) );
  INV_X1 U10317 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12910) );
  NAND2_X1 U10318 ( .A1(n8215), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10319 ( .A1(n8216), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8021) );
  OAI211_X1 U10320 ( .C1(n12910), .C2(n8207), .A(n8022), .B(n8021), .ZN(n8023)
         );
  INV_X1 U10321 ( .A(n8023), .ZN(n8024) );
  NAND2_X1 U10322 ( .A1(n8025), .A2(n8024), .ZN(n12510) );
  INV_X1 U10323 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U10324 ( .A1(n11055), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8029) );
  INV_X1 U10325 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U10326 ( .A1(n8031), .A2(n11237), .ZN(n8032) );
  INV_X1 U10327 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11742) );
  XNOR2_X1 U10328 ( .A(n8046), .B(n11742), .ZN(n11017) );
  NAND2_X1 U10329 ( .A1(n11017), .A2(n12296), .ZN(n8034) );
  OR2_X1 U10330 ( .A1(n12299), .A2(n7376), .ZN(n8033) );
  XNOR2_X1 U10331 ( .A(n12904), .B(n12006), .ZN(n8043) );
  INV_X1 U10332 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U10333 ( .A1(n8035), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10334 ( .A1(n8053), .A2(n8036), .ZN(n12757) );
  NAND2_X1 U10335 ( .A1(n12757), .A2(n8090), .ZN(n8042) );
  INV_X1 U10336 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10337 ( .A1(n8216), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10338 ( .A1(n8215), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8037) );
  OAI211_X1 U10339 ( .C1(n8207), .C2(n8039), .A(n8038), .B(n8037), .ZN(n8040)
         );
  INV_X1 U10340 ( .A(n8040), .ZN(n8041) );
  NAND2_X1 U10341 ( .A1(n8043), .A2(n12152), .ZN(n12195) );
  INV_X1 U10342 ( .A(n8043), .ZN(n8044) );
  NAND2_X1 U10343 ( .A1(n8044), .A2(n8195), .ZN(n8045) );
  INV_X1 U10344 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11363) );
  XNOR2_X1 U10345 ( .A(n11363), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10346 ( .A1(n11130), .A2(n12296), .ZN(n8050) );
  INV_X1 U10347 ( .A(SI_25_), .ZN(n15313) );
  OR2_X1 U10348 ( .A1(n12299), .A2(n15313), .ZN(n8049) );
  XNOR2_X1 U10349 ( .A(n12900), .B(n12006), .ZN(n8061) );
  INV_X1 U10350 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10351 ( .A1(n8052), .A2(n8051), .ZN(n8071) );
  NAND2_X1 U10352 ( .A1(n8053), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10353 ( .A1(n8071), .A2(n8054), .ZN(n12742) );
  NAND2_X1 U10354 ( .A1(n12742), .A2(n8090), .ZN(n8060) );
  INV_X1 U10355 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U10356 ( .A1(n6457), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U10357 ( .A1(n8216), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8055) );
  OAI211_X1 U10358 ( .C1(n8057), .C2(n15325), .A(n8056), .B(n8055), .ZN(n8058)
         );
  INV_X1 U10359 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U10360 ( .A1(n8061), .A2(n12749), .ZN(n8064) );
  INV_X1 U10361 ( .A(n8061), .ZN(n8062) );
  INV_X1 U10362 ( .A(n12749), .ZN(n12509) );
  NAND2_X1 U10363 ( .A1(n8062), .A2(n12509), .ZN(n8063) );
  NAND2_X1 U10364 ( .A1(n12197), .A2(n8064), .ZN(n12270) );
  NAND2_X1 U10365 ( .A1(n11363), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8065) );
  INV_X1 U10366 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11755) );
  INV_X1 U10367 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13687) );
  INV_X1 U10368 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14321) );
  AOI22_X1 U10369 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13687), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14321), .ZN(n8067) );
  XNOR2_X1 U10370 ( .A(n8082), .B(n8067), .ZN(n11199) );
  INV_X1 U10371 ( .A(SI_26_), .ZN(n11198) );
  OR2_X1 U10372 ( .A1(n12299), .A2(n11198), .ZN(n8069) );
  XNOR2_X1 U10373 ( .A(n8238), .B(n10808), .ZN(n8078) );
  NAND2_X1 U10374 ( .A1(n8071), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8072) );
  NAND2_X1 U10375 ( .A1(n8087), .A2(n8072), .ZN(n12729) );
  NAND2_X1 U10376 ( .A1(n12729), .A2(n8090), .ZN(n8077) );
  INV_X1 U10377 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n15227) );
  NAND2_X1 U10378 ( .A1(n8216), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10379 ( .A1(n7890), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8073) );
  OAI211_X1 U10380 ( .C1(n8207), .C2(n15227), .A(n8074), .B(n8073), .ZN(n8075)
         );
  INV_X1 U10381 ( .A(n8075), .ZN(n8076) );
  NOR2_X1 U10382 ( .A1(n8078), .A2(n12736), .ZN(n8079) );
  AOI21_X1 U10383 ( .B1(n8078), .B2(n12736), .A(n8079), .ZN(n12271) );
  INV_X1 U10384 ( .A(n8079), .ZN(n8080) );
  AND2_X1 U10385 ( .A1(n14321), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10386 ( .A1(n13687), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8083) );
  INV_X1 U10387 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9006) );
  INV_X1 U10388 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U10389 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n9006), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14318), .ZN(n8084) );
  XNOR2_X1 U10390 ( .A(n8158), .B(n8084), .ZN(n12001) );
  NAND2_X1 U10391 ( .A1(n12001), .A2(n12296), .ZN(n8086) );
  INV_X1 U10392 ( .A(SI_27_), .ZN(n12002) );
  OR2_X1 U10393 ( .A1(n12299), .A2(n12002), .ZN(n8085) );
  XNOR2_X1 U10394 ( .A(n8199), .B(n10808), .ZN(n8096) );
  INV_X1 U10395 ( .A(n8134), .ZN(n8089) );
  NAND2_X1 U10396 ( .A1(n8087), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10397 ( .A1(n8089), .A2(n8088), .ZN(n12719) );
  NAND2_X1 U10398 ( .A1(n12719), .A2(n8090), .ZN(n8095) );
  INV_X1 U10399 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12896) );
  NAND2_X1 U10400 ( .A1(n8215), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10401 ( .A1(n8216), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8091) );
  OAI211_X1 U10402 ( .C1(n8207), .C2(n12896), .A(n8092), .B(n8091), .ZN(n8093)
         );
  INV_X1 U10403 ( .A(n8093), .ZN(n8094) );
  NOR2_X1 U10404 ( .A1(n8096), .A2(n12697), .ZN(n12004) );
  AOI21_X1 U10405 ( .B1(n8096), .B2(n12697), .A(n12004), .ZN(n8098) );
  OAI21_X1 U10406 ( .B1(n8097), .B2(n8098), .A(n12005), .ZN(n8129) );
  NAND2_X1 U10407 ( .A1(n6458), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8099) );
  OAI21_X1 U10408 ( .B1(n12331), .B2(n8100), .A(n12687), .ZN(n8102) );
  NAND2_X1 U10409 ( .A1(n8102), .A2(n8101), .ZN(n8105) );
  NAND2_X1 U10410 ( .A1(n8101), .A2(n12014), .ZN(n8103) );
  NAND2_X1 U10411 ( .A1(n12331), .A2(n8103), .ZN(n8104) );
  NAND2_X1 U10412 ( .A1(n8105), .A2(n8104), .ZN(n8246) );
  NAND2_X1 U10413 ( .A1(n8246), .A2(n15173), .ZN(n9868) );
  INV_X1 U10414 ( .A(n12987), .ZN(n8121) );
  INV_X1 U10415 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10416 ( .A1(n9424), .A2(n8106), .ZN(n8108) );
  NAND2_X1 U10417 ( .A1(n6848), .A2(n11131), .ZN(n8107) );
  NAND2_X1 U10418 ( .A1(n8108), .A2(n8107), .ZN(n10231) );
  OR2_X1 U10419 ( .A1(n8121), .A2(n10231), .ZN(n8262) );
  INV_X1 U10420 ( .A(n8262), .ZN(n8120) );
  INV_X1 U10421 ( .A(n9424), .ZN(n8119) );
  NOR2_X1 U10422 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .ZN(
        n15336) );
  NOR4_X1 U10423 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8111) );
  NOR4_X1 U10424 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8110) );
  NOR4_X1 U10425 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8109) );
  NAND4_X1 U10426 ( .A1(n15336), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8117) );
  NOR4_X1 U10427 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8115) );
  NOR4_X1 U10428 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8114) );
  NOR4_X1 U10429 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8113) );
  NOR4_X1 U10430 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8112) );
  NAND4_X1 U10431 ( .A1(n8115), .A2(n8114), .A3(n8113), .A4(n8112), .ZN(n8116)
         );
  NOR2_X1 U10432 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  OR2_X1 U10433 ( .A1(n8119), .A2(n8118), .ZN(n8263) );
  NAND2_X1 U10434 ( .A1(n8120), .A2(n8263), .ZN(n8243) );
  AND2_X1 U10435 ( .A1(n8121), .A2(n10231), .ZN(n8261) );
  AND2_X1 U10436 ( .A1(n8261), .A2(n8263), .ZN(n8245) );
  INV_X1 U10437 ( .A(n8245), .ZN(n8145) );
  INV_X1 U10438 ( .A(n12331), .ZN(n12503) );
  AND2_X1 U10439 ( .A1(n12503), .A2(n12687), .ZN(n8212) );
  AND2_X1 U10440 ( .A1(n6476), .A2(n8212), .ZN(n8248) );
  INV_X1 U10441 ( .A(n8248), .ZN(n8122) );
  OAI22_X1 U10442 ( .A1(n9868), .A2(n8243), .B1(n8145), .B2(n8122), .ZN(n8128)
         );
  OAI21_X1 U10443 ( .B1(n6458), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8124) );
  XNOR2_X1 U10444 ( .A(n8123), .B(n8124), .ZN(n9790) );
  AND3_X1 U10445 ( .A1(n8125), .A2(n8126), .A3(n8127), .ZN(n8144) );
  OR2_X1 U10446 ( .A1(n12986), .A2(n8144), .ZN(n9788) );
  INV_X1 U10447 ( .A(n9788), .ZN(n8251) );
  NAND2_X1 U10448 ( .A1(n8128), .A2(n8251), .ZN(n12289) );
  NAND2_X1 U10449 ( .A1(n8129), .A2(n12272), .ZN(n8157) );
  NAND2_X1 U10450 ( .A1(n12014), .A2(n12687), .ZN(n15150) );
  INV_X1 U10451 ( .A(n15150), .ZN(n12493) );
  NAND2_X1 U10452 ( .A1(n15184), .A2(n12493), .ZN(n8130) );
  INV_X1 U10453 ( .A(n8243), .ZN(n8247) );
  NAND2_X1 U10454 ( .A1(n15184), .A2(n8247), .ZN(n8131) );
  NOR2_X1 U10455 ( .A1(n9788), .A2(n8131), .ZN(n8132) );
  INV_X1 U10456 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8133) );
  NOR2_X1 U10457 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  INV_X1 U10458 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U10459 ( .A1(n8216), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10460 ( .A1(n8215), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8136) );
  OAI211_X1 U10461 ( .C1(n8207), .C2(n12892), .A(n8137), .B(n8136), .ZN(n8138)
         );
  INV_X1 U10462 ( .A(n12715), .ZN(n12508) );
  NAND2_X1 U10463 ( .A1(n12014), .A2(n12499), .ZN(n8266) );
  NOR2_X1 U10464 ( .A1(n9788), .A2(n8266), .ZN(n8143) );
  INV_X1 U10465 ( .A(n6417), .ZN(n9796) );
  INV_X1 U10466 ( .A(n8139), .ZN(n9795) );
  NAND2_X1 U10467 ( .A1(n9796), .A2(n9795), .ZN(n9837) );
  NAND2_X1 U10468 ( .A1(n8140), .A2(n9837), .ZN(n8142) );
  NOR2_X1 U10469 ( .A1(n12873), .A2(n8145), .ZN(n8141) );
  AND2_X2 U10470 ( .A1(n8143), .A2(n8141), .ZN(n12282) );
  NOR2_X2 U10471 ( .A1(n12483), .A2(n8142), .ZN(n15143) );
  NAND2_X1 U10472 ( .A1(n8143), .A2(n15143), .ZN(n12502) );
  NAND2_X1 U10473 ( .A1(n8143), .A2(n12487), .ZN(n8244) );
  OR2_X1 U10474 ( .A1(n8244), .A2(n8245), .ZN(n8151) );
  NAND2_X1 U10475 ( .A1(n8246), .A2(n8243), .ZN(n8148) );
  INV_X1 U10476 ( .A(n8144), .ZN(n9128) );
  AND2_X1 U10477 ( .A1(n9790), .A2(n9128), .ZN(n8147) );
  NAND2_X1 U10478 ( .A1(n8248), .A2(n8145), .ZN(n8146) );
  NAND2_X1 U10479 ( .A1(n12487), .A2(n8266), .ZN(n8271) );
  NAND4_X1 U10480 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n8271), .ZN(n8149)
         );
  NAND2_X1 U10481 ( .A1(n8149), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8150) );
  AOI22_X1 U10482 ( .A1(n12719), .A2(n12281), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8152) );
  OAI21_X1 U10483 ( .B1(n12714), .B2(n12285), .A(n8152), .ZN(n8153) );
  AOI21_X1 U10484 ( .B1(n12508), .B2(n12282), .A(n8153), .ZN(n8154) );
  INV_X1 U10485 ( .A(n8155), .ZN(n8156) );
  NAND2_X1 U10486 ( .A1(n8157), .A2(n8156), .ZN(P3_U3154) );
  NAND2_X1 U10487 ( .A1(n14318), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8159) );
  INV_X1 U10488 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8977) );
  INV_X1 U10489 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U10490 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8977), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14315), .ZN(n8161) );
  INV_X1 U10491 ( .A(n8161), .ZN(n8162) );
  INV_X1 U10492 ( .A(SI_28_), .ZN(n13000) );
  OR2_X1 U10493 ( .A1(n12299), .A2(n13000), .ZN(n8163) );
  INV_X1 U10494 ( .A(n10807), .ZN(n10801) );
  NAND2_X1 U10495 ( .A1(n10650), .A2(n10801), .ZN(n8165) );
  NAND2_X1 U10496 ( .A1(n10802), .A2(n12349), .ZN(n8168) );
  INV_X1 U10497 ( .A(n12357), .ZN(n12341) );
  NAND2_X1 U10498 ( .A1(n10856), .A2(n15161), .ZN(n12351) );
  INV_X1 U10499 ( .A(n15161), .ZN(n10528) );
  NAND2_X1 U10500 ( .A1(n10528), .A2(n10856), .ZN(n8169) );
  NAND2_X1 U10501 ( .A1(n10410), .A2(n8169), .ZN(n10855) );
  INV_X1 U10502 ( .A(n8170), .ZN(n15167) );
  NAND2_X1 U10503 ( .A1(n10641), .A2(n15167), .ZN(n12360) );
  NAND2_X1 U10504 ( .A1(n12520), .A2(n8170), .ZN(n12365) );
  NAND2_X1 U10505 ( .A1(n15167), .A2(n12520), .ZN(n8171) );
  INV_X1 U10506 ( .A(n12519), .ZN(n10471) );
  INV_X1 U10507 ( .A(n10222), .ZN(n10638) );
  NAND2_X1 U10508 ( .A1(n10471), .A2(n10638), .ZN(n12368) );
  NAND2_X1 U10509 ( .A1(n12519), .A2(n10222), .ZN(n12361) );
  AND2_X2 U10510 ( .A1(n12368), .A2(n12361), .ZN(n12366) );
  NAND2_X1 U10511 ( .A1(n10471), .A2(n10222), .ZN(n8172) );
  NAND2_X1 U10512 ( .A1(n10437), .A2(n10468), .ZN(n12369) );
  INV_X1 U10513 ( .A(n10468), .ZN(n15172) );
  NAND2_X1 U10514 ( .A1(n15172), .A2(n12518), .ZN(n12374) );
  NAND2_X1 U10515 ( .A1(n12369), .A2(n12374), .ZN(n10423) );
  NAND2_X1 U10516 ( .A1(n12518), .A2(n10468), .ZN(n8173) );
  INV_X1 U10517 ( .A(n12373), .ZN(n10318) );
  NAND2_X1 U10518 ( .A1(n12517), .A2(n10434), .ZN(n8174) );
  INV_X1 U10519 ( .A(n12378), .ZN(n8175) );
  INV_X1 U10520 ( .A(n12384), .ZN(n12383) );
  NAND2_X1 U10521 ( .A1(n12385), .A2(n12383), .ZN(n8177) );
  XNOR2_X1 U10522 ( .A(n12515), .B(n12391), .ZN(n10842) );
  INV_X1 U10523 ( .A(n12391), .ZN(n12390) );
  OR2_X1 U10524 ( .A1(n12514), .A2(n8178), .ZN(n12397) );
  NAND2_X1 U10525 ( .A1(n8178), .A2(n12514), .ZN(n12398) );
  NAND2_X1 U10526 ( .A1(n12397), .A2(n12398), .ZN(n12310) );
  INV_X1 U10527 ( .A(n8178), .ZN(n15183) );
  NAND2_X1 U10528 ( .A1(n15183), .A2(n12514), .ZN(n8179) );
  INV_X1 U10529 ( .A(n14513), .ZN(n11462) );
  OR2_X1 U10530 ( .A1(n14512), .A2(n12246), .ZN(n12407) );
  NAND2_X1 U10531 ( .A1(n14512), .A2(n12246), .ZN(n12408) );
  NAND2_X1 U10532 ( .A1(n12407), .A2(n12408), .ZN(n12314) );
  INV_X1 U10533 ( .A(n12246), .ZN(n12513) );
  NAND2_X1 U10534 ( .A1(n14512), .A2(n12513), .ZN(n8180) );
  NAND2_X1 U10535 ( .A1(n14504), .A2(n12512), .ZN(n12413) );
  NAND2_X1 U10536 ( .A1(n12414), .A2(n12413), .ZN(n12406) );
  OR2_X1 U10537 ( .A1(n14504), .A2(n11468), .ZN(n8182) );
  NAND2_X1 U10538 ( .A1(n14499), .A2(n12511), .ZN(n12420) );
  NAND2_X1 U10539 ( .A1(n12418), .A2(n12420), .ZN(n11402) );
  INV_X1 U10540 ( .A(n12855), .ZN(n12206) );
  NAND2_X1 U10541 ( .A1(n8184), .A2(n12206), .ZN(n8187) );
  INV_X1 U10542 ( .A(n12839), .ZN(n12872) );
  OR2_X1 U10543 ( .A1(n12938), .A2(n12872), .ZN(n12422) );
  NAND2_X1 U10544 ( .A1(n12938), .A2(n12872), .ZN(n12429) );
  INV_X1 U10545 ( .A(n12938), .ZN(n12866) );
  NAND2_X1 U10546 ( .A1(n12938), .A2(n12839), .ZN(n8188) );
  OR2_X1 U10547 ( .A1(n12934), .A2(n12829), .ZN(n12434) );
  NAND2_X1 U10548 ( .A1(n12934), .A2(n12829), .ZN(n12433) );
  NAND2_X1 U10549 ( .A1(n12434), .A2(n12433), .ZN(n12837) );
  INV_X1 U10550 ( .A(n12934), .ZN(n12848) );
  NAND2_X1 U10551 ( .A1(n12934), .A2(n12856), .ZN(n8189) );
  NAND2_X1 U10552 ( .A1(n8190), .A2(n8191), .ZN(n12440) );
  NAND2_X1 U10553 ( .A1(n12977), .A2(n12800), .ZN(n12446) );
  NAND2_X1 U10554 ( .A1(n12445), .A2(n12446), .ZN(n12817) );
  INV_X1 U10555 ( .A(n12800), .ZN(n12828) );
  NAND2_X1 U10556 ( .A1(n12237), .A2(n12816), .ZN(n12449) );
  NAND2_X1 U10557 ( .A1(n12257), .A2(n12768), .ZN(n8193) );
  INV_X1 U10558 ( .A(n12257), .ZN(n12965) );
  NAND2_X1 U10559 ( .A1(n12330), .A2(n8026), .ZN(n8194) );
  INV_X1 U10560 ( .A(n12152), .ZN(n8195) );
  NAND2_X1 U10561 ( .A1(n12904), .A2(n8195), .ZN(n8196) );
  NAND2_X1 U10562 ( .A1(n12751), .A2(n8196), .ZN(n12735) );
  NAND2_X2 U10563 ( .A1(n12474), .A2(n12470), .ZN(n12739) );
  INV_X1 U10564 ( .A(n12900), .ZN(n8197) );
  NAND2_X1 U10565 ( .A1(n8199), .A2(n12726), .ZN(n12701) );
  NAND2_X1 U10566 ( .A1(n12011), .A2(n12715), .ZN(n8239) );
  NAND2_X1 U10567 ( .A1(n8977), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U10568 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11521) );
  XNOR2_X1 U10569 ( .A(n11520), .B(n11521), .ZN(n12994) );
  NAND2_X1 U10570 ( .A1(n12994), .A2(n12296), .ZN(n8203) );
  INV_X1 U10571 ( .A(SI_29_), .ZN(n12996) );
  OR2_X1 U10572 ( .A1(n12299), .A2(n12996), .ZN(n8202) );
  NAND2_X1 U10573 ( .A1(n12688), .A2(n8090), .ZN(n10246) );
  INV_X1 U10574 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10575 ( .A1(n8216), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10576 ( .A1(n7890), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8204) );
  OAI211_X1 U10577 ( .C1(n8207), .C2(n8206), .A(n8205), .B(n8204), .ZN(n8208)
         );
  INV_X1 U10578 ( .A(n8208), .ZN(n8209) );
  NAND2_X1 U10579 ( .A1(n10246), .A2(n8209), .ZN(n12698) );
  INV_X1 U10580 ( .A(n12698), .ZN(n8210) );
  NAND2_X1 U10581 ( .A1(n8255), .A2(n8210), .ZN(n12324) );
  XNOR2_X1 U10582 ( .A(n8211), .B(n6787), .ZN(n8223) );
  INV_X1 U10583 ( .A(n8212), .ZN(n8214) );
  INV_X1 U10584 ( .A(n8101), .ZN(n8213) );
  NAND2_X1 U10585 ( .A1(n8213), .A2(n8100), .ZN(n12500) );
  NAND2_X1 U10586 ( .A1(n6457), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U10587 ( .A1(n8215), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10588 ( .A1(n8216), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8217) );
  AND3_X1 U10589 ( .A1(n8219), .A2(n8218), .A3(n8217), .ZN(n8220) );
  AND2_X1 U10590 ( .A1(n10246), .A2(n8220), .ZN(n12301) );
  NAND2_X1 U10591 ( .A1(n9795), .A2(P3_B_REG_SCAN_IN), .ZN(n8221) );
  NAND2_X1 U10592 ( .A1(n15145), .A2(n8221), .ZN(n12689) );
  OAI22_X1 U10593 ( .A1(n12715), .A2(n12875), .B1(n12301), .B2(n12689), .ZN(
        n8222) );
  INV_X1 U10594 ( .A(n8224), .ZN(n12338) );
  INV_X1 U10595 ( .A(n12339), .ZN(n12345) );
  INV_X1 U10596 ( .A(n12349), .ZN(n10648) );
  NAND2_X1 U10597 ( .A1(n10802), .A2(n10648), .ZN(n12340) );
  NAND2_X1 U10598 ( .A1(n10213), .A2(n12366), .ZN(n10212) );
  NAND2_X1 U10599 ( .A1(n10212), .A2(n12368), .ZN(n10420) );
  INV_X1 U10600 ( .A(n10423), .ZN(n12305) );
  NAND2_X1 U10601 ( .A1(n10420), .A2(n12305), .ZN(n10419) );
  NAND2_X1 U10602 ( .A1(n10419), .A2(n12369), .ZN(n10316) );
  NAND2_X1 U10603 ( .A1(n12385), .A2(n12384), .ZN(n8226) );
  NAND2_X1 U10604 ( .A1(n12515), .A2(n12391), .ZN(n8227) );
  INV_X1 U10605 ( .A(n12515), .ZN(n11205) );
  NAND2_X1 U10606 ( .A1(n11205), .A2(n12390), .ZN(n8228) );
  OR2_X1 U10607 ( .A1(n14513), .A2(n11202), .ZN(n12402) );
  NAND2_X1 U10608 ( .A1(n14513), .A2(n11202), .ZN(n12403) );
  NAND2_X1 U10609 ( .A1(n12402), .A2(n12403), .ZN(n12399) );
  INV_X1 U10610 ( .A(n12398), .ZN(n11088) );
  NOR2_X1 U10611 ( .A1(n12399), .A2(n11088), .ZN(n8229) );
  NAND2_X1 U10612 ( .A1(n11089), .A2(n12402), .ZN(n11229) );
  INV_X1 U10613 ( .A(n12314), .ZN(n8230) );
  INV_X1 U10614 ( .A(n12414), .ZN(n8231) );
  OR2_X1 U10615 ( .A1(n12879), .A2(n12206), .ZN(n12423) );
  NAND2_X1 U10616 ( .A1(n12879), .A2(n12206), .ZN(n12861) );
  NAND2_X1 U10617 ( .A1(n12876), .A2(n12861), .ZN(n8232) );
  NAND2_X1 U10618 ( .A1(n8232), .A2(n12859), .ZN(n12863) );
  INV_X1 U10619 ( .A(n12837), .ZN(n12844) );
  INV_X1 U10620 ( .A(n12446), .ZN(n8233) );
  NAND2_X1 U10621 ( .A1(n12453), .A2(n12781), .ZN(n8235) );
  OR2_X1 U10622 ( .A1(n12453), .A2(n12781), .ZN(n8236) );
  NAND2_X1 U10623 ( .A1(n8237), .A2(n8236), .ZN(n12783) );
  NAND2_X1 U10624 ( .A1(n12257), .A2(n8007), .ZN(n12461) );
  OR2_X1 U10625 ( .A1(n12257), .A2(n8007), .ZN(n12460) );
  NAND2_X1 U10626 ( .A1(n12904), .A2(n12152), .ZN(n12327) );
  NAND2_X1 U10627 ( .A1(n8239), .A2(n12701), .ZN(n12484) );
  XOR2_X1 U10628 ( .A(n12496), .B(n12323), .Z(n12142) );
  OR2_X1 U10629 ( .A1(n9868), .A2(n8266), .ZN(n8241) );
  NOR2_X1 U10630 ( .A1(n12014), .A2(n12687), .ZN(n8240) );
  NAND2_X1 U10631 ( .A1(n12503), .A2(n8240), .ZN(n8270) );
  NAND2_X1 U10632 ( .A1(n12331), .A2(n12493), .ZN(n12893) );
  NAND2_X1 U10633 ( .A1(n8246), .A2(n8245), .ZN(n8250) );
  NAND2_X1 U10634 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  NAND2_X1 U10635 ( .A1(n8250), .A2(n8249), .ZN(n8252) );
  NAND2_X1 U10636 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  INV_X2 U10637 ( .A(n15187), .ZN(n15185) );
  NAND2_X1 U10638 ( .A1(n8274), .A2(n15185), .ZN(n8260) );
  INV_X1 U10639 ( .A(n8255), .ZN(n12144) );
  INV_X1 U10640 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U10641 ( .A1(n8260), .A2(n8259), .ZN(P3_U3456) );
  INV_X1 U10642 ( .A(n8261), .ZN(n8264) );
  NAND3_X1 U10643 ( .A1(n8264), .A2(n8263), .A3(n8262), .ZN(n8265) );
  NOR2_X1 U10644 ( .A1(n9788), .A2(n8265), .ZN(n10236) );
  NAND2_X1 U10645 ( .A1(n15184), .A2(n12014), .ZN(n8268) );
  NAND2_X1 U10646 ( .A1(n12503), .A2(n12499), .ZN(n8267) );
  INV_X1 U10647 ( .A(n8266), .ZN(n12492) );
  AOI21_X1 U10648 ( .B1(n8268), .B2(n8267), .A(n12492), .ZN(n8269) );
  OAI21_X1 U10649 ( .B1(n8269), .B2(n12487), .A(n10231), .ZN(n8273) );
  NAND2_X1 U10650 ( .A1(n8270), .A2(n12483), .ZN(n10233) );
  NAND2_X1 U10651 ( .A1(n8271), .A2(n10233), .ZN(n10232) );
  INV_X1 U10652 ( .A(n10231), .ZN(n12985) );
  NAND2_X1 U10653 ( .A1(n10232), .A2(n12985), .ZN(n8272) );
  AND3_X2 U10654 ( .A1(n10236), .A2(n8273), .A3(n8272), .ZN(n15199) );
  NAND2_X1 U10655 ( .A1(n8274), .A2(n15199), .ZN(n8279) );
  NAND2_X1 U10656 ( .A1(n15199), .A2(n15184), .ZN(n12933) );
  NAND2_X1 U10657 ( .A1(n8255), .A2(n8275), .ZN(n8277) );
  OR2_X1 U10658 ( .A1(n15199), .A2(n8206), .ZN(n8276) );
  NAND2_X1 U10659 ( .A1(n8279), .A2(n8278), .ZN(P3_U3488) );
  INV_X1 U10660 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13531) );
  NOR2_X1 U10661 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8290) );
  NOR2_X1 U10662 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8289) );
  NOR2_X1 U10663 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8295) );
  INV_X1 U10664 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8294) );
  INV_X1 U10665 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8293) );
  INV_X1 U10666 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8321) );
  XNOR2_X2 U10667 ( .A(n8297), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10668 ( .A1(n8360), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8298) );
  OAI21_X1 U10669 ( .B1(n13531), .B2(n8389), .A(n8298), .ZN(n8302) );
  INV_X1 U10670 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8300) );
  INV_X1 U10671 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13545) );
  OR2_X1 U10672 ( .A1(n6410), .A2(n13545), .ZN(n8304) );
  INV_X1 U10673 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8307) );
  INV_X1 U10674 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8308) );
  INV_X1 U10675 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8733) );
  AND2_X1 U10676 ( .A1(n8308), .A2(n8733), .ZN(n8309) );
  INV_X1 U10677 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10678 ( .A1(n8312), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8313) );
  XNOR2_X1 U10679 ( .A(n8313), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U10680 ( .A1(n8951), .A2(n9674), .ZN(n8353) );
  INV_X1 U10681 ( .A(n8353), .ZN(n8316) );
  NAND2_X1 U10682 ( .A1(n6460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8314) );
  INV_X1 U10683 ( .A(n9075), .ZN(n9087) );
  INV_X1 U10684 ( .A(n9651), .ZN(n8319) );
  NAND2_X1 U10685 ( .A1(n6413), .A2(n6420), .ZN(n8335) );
  INV_X1 U10686 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10687 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8325) );
  MUX2_X1 U10688 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8325), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8328) );
  INV_X1 U10689 ( .A(n8326), .ZN(n8327) );
  NAND2_X1 U10690 ( .A1(n8328), .A2(n8327), .ZN(n13151) );
  INV_X1 U10691 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9133) );
  AND2_X1 U10692 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8329) );
  NAND2_X1 U10693 ( .A1(n8330), .A2(n8329), .ZN(n9269) );
  OAI21_X1 U10694 ( .B1(n9144), .B2(n8331), .A(n9269), .ZN(n8374) );
  XNOR2_X1 U10695 ( .A(n8374), .B(n8375), .ZN(n9585) );
  OR2_X1 U10696 ( .A1(n8371), .A2(n9585), .ZN(n8333) );
  OR2_X1 U10697 ( .A1(n8400), .A2(n9152), .ZN(n8332) );
  NAND2_X1 U10698 ( .A1(n9053), .A2(n8842), .ZN(n8334) );
  AOI22_X1 U10699 ( .A1(n8343), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n8341) );
  INV_X1 U10700 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10701 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8337) );
  OAI21_X1 U10702 ( .B1(n8338), .B2(P2_IR_REG_30__SCAN_IN), .A(n8337), .ZN(
        n8339) );
  NAND2_X1 U10703 ( .A1(n8336), .A2(n8339), .ZN(n8340) );
  OAI21_X1 U10704 ( .B1(n8336), .B2(n8341), .A(n8340), .ZN(n8342) );
  NAND2_X1 U10705 ( .A1(n8342), .A2(n13676), .ZN(n8351) );
  AOI22_X1 U10706 ( .A1(n8343), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n8347) );
  INV_X1 U10707 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U10708 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n8344) );
  OAI21_X1 U10709 ( .B1(n9416), .B2(P2_IR_REG_30__SCAN_IN), .A(n8344), .ZN(
        n8345) );
  NAND2_X1 U10710 ( .A1(n8336), .A2(n8345), .ZN(n8346) );
  OAI21_X1 U10711 ( .B1(n8336), .B2(n8347), .A(n8346), .ZN(n8349) );
  NAND2_X1 U10712 ( .A1(n8349), .A2(n8348), .ZN(n8350) );
  XNOR2_X1 U10713 ( .A(n9144), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13690) );
  INV_X1 U10714 ( .A(n13530), .ZN(n10305) );
  NAND2_X1 U10715 ( .A1(n13146), .A2(n10305), .ZN(n9054) );
  INV_X1 U10716 ( .A(n9054), .ZN(n9767) );
  NAND2_X1 U10717 ( .A1(n9767), .A2(n6420), .ZN(n8358) );
  BUF_X1 U10718 ( .A(n8353), .Z(n8354) );
  OAI211_X1 U10719 ( .C1(n9649), .C2(n10369), .A(n9054), .B(n8316), .ZN(n8356)
         );
  INV_X1 U10720 ( .A(n13146), .ZN(n10350) );
  AND2_X1 U10721 ( .A1(n10350), .A2(n13530), .ZN(n13539) );
  NAND2_X1 U10722 ( .A1(n13539), .A2(n8842), .ZN(n8357) );
  AND3_X1 U10723 ( .A1(n8358), .A2(n8357), .A3(n8356), .ZN(n8359) );
  NAND2_X1 U10724 ( .A1(n8360), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8366) );
  INV_X1 U10725 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10619) );
  OR2_X1 U10726 ( .A1(n8389), .A2(n10619), .ZN(n8365) );
  INV_X1 U10727 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9331) );
  OR2_X1 U10728 ( .A1(n6409), .A2(n9331), .ZN(n8364) );
  INV_X1 U10729 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8362) );
  OR2_X1 U10730 ( .A1(n8361), .A2(n8362), .ZN(n8363) );
  NAND2_X1 U10731 ( .A1(n13144), .A2(n6426), .ZN(n8379) );
  NOR2_X1 U10732 ( .A1(n8326), .A2(n13671), .ZN(n8367) );
  MUX2_X1 U10733 ( .A(n13671), .B(n8367), .S(P2_IR_REG_2__SCAN_IN), .Z(n8368)
         );
  INV_X1 U10734 ( .A(n8368), .ZN(n8370) );
  INV_X1 U10735 ( .A(n8417), .ZN(n8369) );
  NAND2_X1 U10736 ( .A1(n8370), .A2(n8369), .ZN(n13159) );
  NOR2_X1 U10737 ( .A1(n8372), .A2(n9150), .ZN(n8373) );
  MUX2_X1 U10738 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8376), .Z(n8398) );
  XNOR2_X1 U10739 ( .A(n8398), .B(SI_2_), .ZN(n8397) );
  XNOR2_X1 U10740 ( .A(n8396), .B(n8397), .ZN(n9604) );
  OR2_X1 U10741 ( .A1(n8400), .A2(n9138), .ZN(n8377) );
  NAND2_X1 U10742 ( .A1(n9046), .A2(n10621), .ZN(n8378) );
  NAND2_X1 U10743 ( .A1(n8379), .A2(n8378), .ZN(n8384) );
  NAND2_X1 U10744 ( .A1(n8383), .A2(n8384), .ZN(n8382) );
  AOI22_X1 U10745 ( .A1(n13144), .A2(n9046), .B1(n10621), .B2(n6426), .ZN(
        n8380) );
  INV_X1 U10746 ( .A(n8380), .ZN(n8381) );
  NAND2_X1 U10747 ( .A1(n8382), .A2(n8381), .ZN(n8388) );
  INV_X1 U10748 ( .A(n8383), .ZN(n8386) );
  NAND2_X1 U10749 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  NAND2_X1 U10750 ( .A1(n8388), .A2(n8387), .ZN(n8407) );
  NAND2_X1 U10751 ( .A1(n8980), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8394) );
  OR2_X1 U10752 ( .A1(n8389), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8393) );
  INV_X1 U10753 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9333) );
  OR2_X1 U10754 ( .A1(n6410), .A2(n9333), .ZN(n8392) );
  INV_X1 U10755 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10756 ( .A1(n8361), .A2(n8390), .ZN(n8391) );
  NAND2_X1 U10757 ( .A1(n13143), .A2(n9046), .ZN(n8404) );
  OR2_X1 U10758 ( .A1(n8417), .A2(n13671), .ZN(n8395) );
  XNOR2_X1 U10759 ( .A(n8395), .B(n8416), .ZN(n13174) );
  NAND2_X1 U10760 ( .A1(n8398), .A2(SI_2_), .ZN(n8399) );
  INV_X1 U10761 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9141) );
  XNOR2_X1 U10762 ( .A(n8421), .B(n8420), .ZN(n9926) );
  OR2_X1 U10763 ( .A1(n8455), .A2(n9926), .ZN(n8402) );
  BUF_X4 U10764 ( .A(n8400), .Z(n9007) );
  OR2_X1 U10765 ( .A1(n9007), .A2(n9143), .ZN(n8401) );
  OAI211_X1 U10766 ( .C1(n9090), .C2(n13174), .A(n8402), .B(n8401), .ZN(n14783) );
  NAND2_X1 U10767 ( .A1(n14783), .A2(n6426), .ZN(n8403) );
  NAND2_X1 U10768 ( .A1(n8404), .A2(n8403), .ZN(n8406) );
  AOI22_X1 U10769 ( .A1(n13143), .A2(n6426), .B1(n9046), .B2(n14783), .ZN(
        n8405) );
  NAND2_X1 U10770 ( .A1(n9010), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8415) );
  INV_X1 U10771 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9358) );
  OR2_X1 U10772 ( .A1(n9012), .A2(n9358), .ZN(n8414) );
  AND2_X1 U10773 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8439) );
  INV_X1 U10774 ( .A(n8439), .ZN(n8441) );
  INV_X1 U10775 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8409) );
  INV_X1 U10776 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10777 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  NAND2_X1 U10778 ( .A1(n8441), .A2(n8410), .ZN(n10539) );
  OR2_X1 U10779 ( .A1(n9017), .A2(n10539), .ZN(n8413) );
  INV_X1 U10780 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9336) );
  OR2_X1 U10781 ( .A1(n6410), .A2(n9336), .ZN(n8412) );
  NAND4_X2 U10782 ( .A1(n8415), .A2(n8414), .A3(n8413), .A4(n8412), .ZN(n13142) );
  NAND2_X1 U10783 ( .A1(n13142), .A2(n6426), .ZN(n8428) );
  NAND2_X1 U10784 ( .A1(n8417), .A2(n8416), .ZN(n8479) );
  NAND2_X1 U10785 ( .A1(n8479), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8418) );
  INV_X1 U10786 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U10787 ( .A1(n8418), .A2(n8477), .ZN(n8447) );
  OR2_X1 U10788 ( .A1(n8418), .A2(n8477), .ZN(n8419) );
  NAND2_X1 U10789 ( .A1(n8447), .A2(n8419), .ZN(n14809) );
  INV_X1 U10790 ( .A(n8422), .ZN(n8423) );
  NAND2_X1 U10791 ( .A1(n8423), .A2(SI_3_), .ZN(n8424) );
  OR2_X1 U10792 ( .A1(n9007), .A2(n9147), .ZN(n8426) );
  NAND2_X1 U10793 ( .A1(n9046), .A2(n10541), .ZN(n8427) );
  NAND2_X1 U10794 ( .A1(n8428), .A2(n8427), .ZN(n8434) );
  NAND2_X1 U10795 ( .A1(n8433), .A2(n8434), .ZN(n8432) );
  NAND2_X1 U10796 ( .A1(n13142), .A2(n9046), .ZN(n8430) );
  NAND2_X1 U10797 ( .A1(n10541), .A2(n6426), .ZN(n8429) );
  NAND2_X1 U10798 ( .A1(n8430), .A2(n8429), .ZN(n8431) );
  NAND2_X1 U10799 ( .A1(n8432), .A2(n8431), .ZN(n8438) );
  INV_X1 U10800 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U10801 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  NAND2_X1 U10802 ( .A1(n9010), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8446) );
  INV_X1 U10803 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9361) );
  OR2_X1 U10804 ( .A1(n9012), .A2(n9361), .ZN(n8445) );
  INV_X1 U10805 ( .A(n8462), .ZN(n8464) );
  INV_X1 U10806 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10807 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  NAND2_X1 U10808 ( .A1(n8464), .A2(n8442), .ZN(n11987) );
  OR2_X1 U10809 ( .A1(n9017), .A2(n11987), .ZN(n8444) );
  INV_X1 U10810 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10402) );
  OR2_X1 U10811 ( .A1(n6410), .A2(n10402), .ZN(n8443) );
  NAND4_X1 U10812 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n13141) );
  NAND2_X1 U10813 ( .A1(n13141), .A2(n9046), .ZN(n8459) );
  NAND2_X1 U10814 ( .A1(n8447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U10815 ( .A(n8448), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14819) );
  AOI22_X1 U10816 ( .A1(n8772), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8771), .B2(
        n14819), .ZN(n8457) );
  INV_X1 U10817 ( .A(n8451), .ZN(n8452) );
  NAND2_X1 U10818 ( .A1(n8452), .A2(SI_4_), .ZN(n8453) );
  MUX2_X1 U10819 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6411), .Z(n8474) );
  XNOR2_X1 U10820 ( .A(n8473), .B(n8471), .ZN(n9940) );
  NAND2_X1 U10821 ( .A1(n9940), .A2(n9005), .ZN(n8456) );
  NAND2_X1 U10822 ( .A1(n8457), .A2(n8456), .ZN(n15001) );
  NAND2_X1 U10823 ( .A1(n15001), .A2(n6426), .ZN(n8458) );
  NAND2_X1 U10824 ( .A1(n13141), .A2(n6426), .ZN(n8460) );
  OAI21_X1 U10825 ( .B1(n7032), .B2(n8842), .A(n8460), .ZN(n8461) );
  NAND2_X1 U10826 ( .A1(n9010), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8470) );
  INV_X1 U10827 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9364) );
  OR2_X1 U10828 ( .A1(n9012), .A2(n9364), .ZN(n8469) );
  INV_X1 U10829 ( .A(n8499), .ZN(n8466) );
  INV_X1 U10830 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10831 ( .A1(n8464), .A2(n8463), .ZN(n8465) );
  NAND2_X1 U10832 ( .A1(n8466), .A2(n8465), .ZN(n10718) );
  OR2_X1 U10833 ( .A1(n9017), .A2(n10718), .ZN(n8468) );
  INV_X1 U10834 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9341) );
  OR2_X1 U10835 ( .A1(n6409), .A2(n9341), .ZN(n8467) );
  NAND4_X1 U10836 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n13140) );
  NAND2_X1 U10837 ( .A1(n13140), .A2(n6426), .ZN(n8488) );
  NAND2_X1 U10838 ( .A1(n8474), .A2(SI_5_), .ZN(n8475) );
  NAND2_X1 U10839 ( .A1(n10073), .A2(n9005), .ZN(n8486) );
  NAND2_X1 U10840 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  NAND2_X1 U10841 ( .A1(n8481), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8480) );
  MUX2_X1 U10842 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8480), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8484) );
  INV_X1 U10843 ( .A(n8481), .ZN(n8483) );
  INV_X1 U10844 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10845 ( .A1(n8483), .A2(n8482), .ZN(n8495) );
  NAND2_X1 U10846 ( .A1(n8484), .A2(n8495), .ZN(n13188) );
  INV_X1 U10847 ( .A(n13188), .ZN(n13183) );
  AOI22_X1 U10848 ( .A1(n8772), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8771), .B2(
        n13183), .ZN(n8485) );
  NAND2_X1 U10849 ( .A1(n8486), .A2(n8485), .ZN(n10720) );
  NAND2_X1 U10850 ( .A1(n10720), .A2(n9046), .ZN(n8487) );
  AOI22_X1 U10851 ( .A1(n9046), .A2(n13140), .B1(n10720), .B2(n6426), .ZN(
        n8489) );
  NAND2_X1 U10852 ( .A1(n8492), .A2(SI_6_), .ZN(n8493) );
  MUX2_X1 U10853 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6411), .Z(n8510) );
  XNOR2_X1 U10854 ( .A(n8509), .B(n8508), .ZN(n10078) );
  NAND2_X1 U10855 ( .A1(n10078), .A2(n9005), .ZN(n8498) );
  NAND2_X1 U10856 ( .A1(n8495), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8494) );
  MUX2_X1 U10857 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8494), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8496) );
  AOI22_X1 U10858 ( .A1(n8772), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8771), .B2(
        n9545), .ZN(n8497) );
  NAND2_X1 U10859 ( .A1(n15020), .A2(n6426), .ZN(n8505) );
  NAND2_X1 U10860 ( .A1(n9010), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8503) );
  INV_X1 U10861 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9367) );
  OR2_X1 U10862 ( .A1(n9012), .A2(n9367), .ZN(n8502) );
  OAI21_X1 U10863 ( .B1(n8499), .B2(P2_REG3_REG_7__SCAN_IN), .A(n8515), .ZN(
        n10769) );
  OR2_X1 U10864 ( .A1(n9017), .A2(n10769), .ZN(n8501) );
  INV_X1 U10865 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9344) );
  OR2_X1 U10866 ( .A1(n6409), .A2(n9344), .ZN(n8500) );
  NAND4_X1 U10867 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(n13139) );
  NAND2_X1 U10868 ( .A1(n13139), .A2(n9046), .ZN(n8504) );
  AOI22_X1 U10869 ( .A1(n15020), .A2(n9046), .B1(n13139), .B2(n6426), .ZN(
        n8506) );
  MUX2_X1 U10870 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6412), .Z(n8535) );
  XNOR2_X1 U10871 ( .A(n8534), .B(n8532), .ZN(n10273) );
  NAND2_X1 U10872 ( .A1(n10273), .A2(n9005), .ZN(n8513) );
  NAND2_X1 U10873 ( .A1(n8538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8511) );
  XNOR2_X1 U10874 ( .A(n8511), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U10875 ( .A1(n8772), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8771), .B2(
        n13203), .ZN(n8512) );
  NAND2_X1 U10876 ( .A1(n15029), .A2(n9046), .ZN(n8522) );
  NAND2_X1 U10877 ( .A1(n9010), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8520) );
  INV_X1 U10878 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9546) );
  OR2_X1 U10879 ( .A1(n9012), .A2(n9546), .ZN(n8519) );
  INV_X1 U10880 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8514) );
  AND2_X1 U10881 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  OR2_X1 U10882 ( .A1(n8516), .A2(n8543), .ZN(n10870) );
  OR2_X1 U10883 ( .A1(n9017), .A2(n10870), .ZN(n8518) );
  INV_X1 U10884 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10748) );
  OR2_X1 U10885 ( .A1(n6409), .A2(n10748), .ZN(n8517) );
  NAND4_X1 U10886 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n13138) );
  NAND2_X1 U10887 ( .A1(n13138), .A2(n6426), .ZN(n8521) );
  NAND2_X1 U10888 ( .A1(n8522), .A2(n8521), .ZN(n8527) );
  INV_X1 U10889 ( .A(n13138), .ZN(n10923) );
  NAND2_X1 U10890 ( .A1(n15029), .A2(n8842), .ZN(n8523) );
  OAI21_X1 U10891 ( .B1(n10923), .B2(n8842), .A(n8523), .ZN(n8524) );
  NAND2_X1 U10892 ( .A1(n8525), .A2(n8524), .ZN(n8531) );
  INV_X1 U10893 ( .A(n8526), .ZN(n8529) );
  INV_X1 U10894 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10895 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U10896 ( .A1(n8535), .A2(SI_8_), .ZN(n8536) );
  MUX2_X1 U10897 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6411), .Z(n8556) );
  XNOR2_X1 U10898 ( .A(n8555), .B(n8553), .ZN(n10555) );
  NAND2_X1 U10899 ( .A1(n10555), .A2(n9005), .ZN(n8541) );
  OAI21_X1 U10900 ( .B1(n8538), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10901 ( .A(n8539), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U10902 ( .A1(n8772), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8771), .B2(
        n9550), .ZN(n8540) );
  NAND2_X1 U10903 ( .A1(n15038), .A2(n6426), .ZN(n8550) );
  NAND2_X1 U10904 ( .A1(n8980), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8548) );
  INV_X1 U10905 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8542) );
  OR2_X1 U10906 ( .A1(n8361), .A2(n8542), .ZN(n8547) );
  NAND2_X1 U10907 ( .A1(n8543), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8566) );
  OR2_X1 U10908 ( .A1(n8543), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10909 ( .A1(n8566), .A2(n8544), .ZN(n10937) );
  OR2_X1 U10910 ( .A1(n9017), .A2(n10937), .ZN(n8546) );
  INV_X1 U10911 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10938) );
  OR2_X1 U10912 ( .A1(n6410), .A2(n10938), .ZN(n8545) );
  NAND4_X1 U10913 ( .A1(n8548), .A2(n8547), .A3(n8546), .A4(n8545), .ZN(n13137) );
  NAND2_X1 U10914 ( .A1(n13137), .A2(n9046), .ZN(n8549) );
  NAND2_X1 U10915 ( .A1(n8550), .A2(n8549), .ZN(n8552) );
  AOI22_X1 U10916 ( .A1(n15038), .A2(n9046), .B1(n13137), .B2(n6426), .ZN(
        n8551) );
  NAND2_X1 U10917 ( .A1(n8556), .A2(SI_9_), .ZN(n8557) );
  MUX2_X1 U10918 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6412), .Z(n8581) );
  NAND2_X1 U10919 ( .A1(n10560), .A2(n9005), .ZN(n8564) );
  NOR2_X1 U10920 ( .A1(n8559), .A2(n13671), .ZN(n8560) );
  MUX2_X1 U10921 ( .A(n13671), .B(n8560), .S(P2_IR_REG_10__SCAN_IN), .Z(n8562)
         );
  AND2_X1 U10922 ( .A1(n8559), .A2(n8561), .ZN(n8586) );
  NOR2_X1 U10923 ( .A1(n8562), .A2(n8586), .ZN(n14848) );
  AOI22_X1 U10924 ( .A1(n8772), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8771), 
        .B2(n14848), .ZN(n8563) );
  NAND2_X1 U10925 ( .A1(n13024), .A2(n9046), .ZN(n8573) );
  NAND2_X1 U10926 ( .A1(n9010), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8571) );
  INV_X1 U10927 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9551) );
  OR2_X1 U10928 ( .A1(n9012), .A2(n9551), .ZN(n8570) );
  INV_X1 U10929 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10930 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U10931 ( .A1(n8591), .A2(n8567), .ZN(n13025) );
  OR2_X1 U10932 ( .A1(n9017), .A2(n13025), .ZN(n8569) );
  INV_X1 U10933 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11044) );
  OR2_X1 U10934 ( .A1(n6409), .A2(n11044), .ZN(n8568) );
  NAND4_X1 U10935 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(n13136) );
  NAND2_X1 U10936 ( .A1(n13136), .A2(n8842), .ZN(n8572) );
  NAND2_X1 U10937 ( .A1(n8573), .A2(n8572), .ZN(n8576) );
  NAND2_X1 U10938 ( .A1(n13024), .A2(n6426), .ZN(n8574) );
  OAI21_X1 U10939 ( .B1(n11172), .B2(n8842), .A(n8574), .ZN(n8575) );
  MUX2_X1 U10940 ( .A(n9216), .B(n9211), .S(n6412), .Z(n8583) );
  INV_X1 U10941 ( .A(n8583), .ZN(n8584) );
  NAND2_X1 U10942 ( .A1(n8584), .A2(SI_11_), .ZN(n8585) );
  XNOR2_X1 U10943 ( .A(n8604), .B(n8603), .ZN(n10573) );
  NAND2_X1 U10944 ( .A1(n10573), .A2(n9005), .ZN(n8589) );
  INV_X1 U10945 ( .A(n8586), .ZN(n8608) );
  NAND2_X1 U10946 ( .A1(n8608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8587) );
  XNOR2_X1 U10947 ( .A(n8587), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U10948 ( .A1(n8772), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8771), 
        .B2(n9975), .ZN(n8588) );
  NAND2_X2 U10949 ( .A1(n8589), .A2(n8588), .ZN(n15054) );
  NAND2_X1 U10950 ( .A1(n15054), .A2(n8842), .ZN(n8598) );
  NAND2_X1 U10951 ( .A1(n8980), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8596) );
  INV_X1 U10952 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8590) );
  OR2_X1 U10953 ( .A1(n8361), .A2(n8590), .ZN(n8595) );
  INV_X1 U10954 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9541) );
  AND2_X1 U10955 ( .A1(n8591), .A2(n9541), .ZN(n8592) );
  OR2_X1 U10956 ( .A1(n8592), .A2(n8613), .ZN(n11188) );
  OR2_X1 U10957 ( .A1(n9017), .A2(n11188), .ZN(n8594) );
  INV_X1 U10958 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11191) );
  OR2_X1 U10959 ( .A1(n6410), .A2(n11191), .ZN(n8593) );
  NAND4_X1 U10960 ( .A1(n8596), .A2(n8595), .A3(n8594), .A4(n8593), .ZN(n13135) );
  NAND2_X1 U10961 ( .A1(n13135), .A2(n9046), .ZN(n8597) );
  NAND2_X1 U10962 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  AOI22_X1 U10963 ( .A1(n15054), .A2(n9046), .B1(n13135), .B2(n6426), .ZN(
        n8599) );
  MUX2_X1 U10964 ( .A(n9380), .B(n9383), .S(n6411), .Z(n8605) );
  INV_X1 U10965 ( .A(SI_12_), .ZN(n9191) );
  INV_X1 U10966 ( .A(n8605), .ZN(n8606) );
  NAND2_X1 U10967 ( .A1(n8606), .A2(SI_12_), .ZN(n8607) );
  XNOR2_X1 U10968 ( .A(n8624), .B(n7553), .ZN(n10960) );
  NAND2_X1 U10969 ( .A1(n10960), .A2(n9005), .ZN(n8611) );
  OR2_X1 U10970 ( .A1(n8608), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U10971 ( .A1(n8630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U10972 ( .A(n8609), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14861) );
  AOI22_X1 U10973 ( .A1(n8772), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8771), 
        .B2(n14861), .ZN(n8610) );
  NAND2_X1 U10974 ( .A1(n11243), .A2(n9046), .ZN(n8621) );
  NAND2_X1 U10975 ( .A1(n9010), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8619) );
  INV_X1 U10976 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8612) );
  OR2_X1 U10977 ( .A1(n9012), .A2(n8612), .ZN(n8618) );
  NOR2_X1 U10978 ( .A1(n8613), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8614) );
  OR2_X1 U10979 ( .A1(n8635), .A2(n8614), .ZN(n11179) );
  OR2_X1 U10980 ( .A1(n9017), .A2(n11179), .ZN(n8617) );
  INV_X1 U10981 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8615) );
  OR2_X1 U10982 ( .A1(n6410), .A2(n8615), .ZN(n8616) );
  NAND4_X1 U10983 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n13134) );
  NAND2_X1 U10984 ( .A1(n13134), .A2(n6426), .ZN(n8620) );
  NAND2_X1 U10985 ( .A1(n8621), .A2(n8620), .ZN(n8623) );
  AOI22_X1 U10986 ( .A1(n11243), .A2(n6426), .B1(n9046), .B2(n13134), .ZN(
        n8622) );
  MUX2_X1 U10987 ( .A(n11059), .B(n9465), .S(n6411), .Z(n8627) );
  INV_X1 U10988 ( .A(n8627), .ZN(n8628) );
  NAND2_X1 U10989 ( .A1(n8628), .A2(SI_13_), .ZN(n8629) );
  XNOR2_X1 U10990 ( .A(n8652), .B(n7554), .ZN(n11058) );
  NAND2_X1 U10991 ( .A1(n11058), .A2(n9005), .ZN(n8633) );
  OAI21_X1 U10992 ( .B1(n8630), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8631) );
  XNOR2_X1 U10993 ( .A(n8631), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U10994 ( .A1(n8772), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8771), 
        .B2(n9976), .ZN(n8632) );
  NAND2_X1 U10995 ( .A1(n14795), .A2(n6426), .ZN(n8642) );
  NAND2_X1 U10996 ( .A1(n8980), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8640) );
  INV_X1 U10997 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8634) );
  OR2_X1 U10998 ( .A1(n8361), .A2(n8634), .ZN(n8639) );
  OR2_X1 U10999 ( .A1(n8635), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U11000 ( .A1(n8658), .A2(n8636), .ZN(n14798) );
  OR2_X1 U11001 ( .A1(n9017), .A2(n14798), .ZN(n8638) );
  INV_X1 U11002 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13217) );
  OR2_X1 U11003 ( .A1(n6409), .A2(n13217), .ZN(n8637) );
  NAND4_X1 U11004 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n13133) );
  NAND2_X1 U11005 ( .A1(n13133), .A2(n9046), .ZN(n8641) );
  NAND2_X1 U11006 ( .A1(n8642), .A2(n8641), .ZN(n8647) );
  INV_X1 U11007 ( .A(n13133), .ZN(n11413) );
  NAND2_X1 U11008 ( .A1(n14795), .A2(n9046), .ZN(n8643) );
  OAI21_X1 U11009 ( .B1(n11413), .B2(n9046), .A(n8643), .ZN(n8644) );
  NAND2_X1 U11010 ( .A1(n8645), .A2(n8644), .ZN(n8651) );
  INV_X1 U11011 ( .A(n8646), .ZN(n8649) );
  INV_X1 U11012 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U11013 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  XNOR2_X1 U11014 ( .A(n8697), .B(SI_14_), .ZN(n8671) );
  MUX2_X1 U11015 ( .A(n9679), .B(n9681), .S(n6412), .Z(n8670) );
  XNOR2_X1 U11016 ( .A(n8671), .B(n8670), .ZN(n11146) );
  NAND2_X1 U11017 ( .A1(n11146), .A2(n9005), .ZN(n8657) );
  NAND2_X1 U11018 ( .A1(n8654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8655) );
  XNOR2_X1 U11019 ( .A(n8655), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U11020 ( .A1(n8772), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8771), 
        .B2(n14876), .ZN(n8656) );
  NAND2_X1 U11021 ( .A1(n11512), .A2(n9046), .ZN(n8666) );
  NAND2_X1 U11022 ( .A1(n8980), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8664) );
  INV_X1 U11023 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U11024 ( .A1(n8658), .A2(n11299), .ZN(n8659) );
  NAND2_X1 U11025 ( .A1(n8684), .A2(n8659), .ZN(n11420) );
  OR2_X1 U11026 ( .A1(n9017), .A2(n11420), .ZN(n8663) );
  INV_X1 U11027 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11419) );
  OR2_X1 U11028 ( .A1(n6409), .A2(n11419), .ZN(n8662) );
  INV_X1 U11029 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8660) );
  OR2_X1 U11030 ( .A1(n8361), .A2(n8660), .ZN(n8661) );
  NAND4_X1 U11031 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n13132) );
  NAND2_X1 U11032 ( .A1(n13132), .A2(n6426), .ZN(n8665) );
  NAND2_X1 U11033 ( .A1(n8666), .A2(n8665), .ZN(n8668) );
  AOI22_X1 U11034 ( .A1(n11512), .A2(n6426), .B1(n9046), .B2(n13132), .ZN(
        n8667) );
  NAND2_X1 U11035 ( .A1(n8671), .A2(n8698), .ZN(n8674) );
  INV_X1 U11036 ( .A(n8697), .ZN(n8672) );
  NAND2_X1 U11037 ( .A1(n8672), .A2(SI_14_), .ZN(n8673) );
  NAND2_X1 U11038 ( .A1(n8674), .A2(n8673), .ZN(n8678) );
  MUX2_X1 U11039 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6412), .Z(n8675) );
  INV_X1 U11040 ( .A(n8675), .ZN(n8676) );
  INV_X1 U11041 ( .A(SI_15_), .ZN(n9400) );
  NAND2_X1 U11042 ( .A1(n8676), .A2(n9400), .ZN(n8699) );
  NAND2_X1 U11043 ( .A1(n8701), .A2(n8699), .ZN(n8677) );
  NAND2_X1 U11044 ( .A1(n11337), .A2(n9005), .ZN(n8682) );
  NAND2_X1 U11045 ( .A1(n8679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U11046 ( .A(n8680), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U11047 ( .A1(n8772), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8771), 
        .B2(n14884), .ZN(n8681) );
  NAND2_X1 U11048 ( .A1(n13640), .A2(n6426), .ZN(n8691) );
  NAND2_X1 U11049 ( .A1(n9010), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8689) );
  INV_X1 U11050 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13233) );
  OR2_X1 U11051 ( .A1(n9012), .A2(n13233), .ZN(n8688) );
  INV_X1 U11052 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11053 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  NAND2_X1 U11054 ( .A1(n8712), .A2(n8685), .ZN(n11516) );
  OR2_X1 U11055 ( .A1(n9017), .A2(n11516), .ZN(n8687) );
  INV_X1 U11056 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11507) );
  OR2_X1 U11057 ( .A1(n6409), .A2(n11507), .ZN(n8686) );
  NAND4_X1 U11058 ( .A1(n8689), .A2(n8688), .A3(n8687), .A4(n8686), .ZN(n13131) );
  NAND2_X1 U11059 ( .A1(n13131), .A2(n9046), .ZN(n8690) );
  NAND2_X1 U11060 ( .A1(n8691), .A2(n8690), .ZN(n8694) );
  INV_X1 U11061 ( .A(n13131), .ZN(n13509) );
  NAND2_X1 U11062 ( .A1(n13640), .A2(n9046), .ZN(n8692) );
  OAI21_X1 U11063 ( .B1(n13509), .B2(n9046), .A(n8692), .ZN(n8693) );
  INV_X1 U11064 ( .A(n8694), .ZN(n8695) );
  NAND2_X1 U11065 ( .A1(n8698), .A2(SI_14_), .ZN(n8696) );
  NOR2_X1 U11066 ( .A1(n8698), .A2(SI_14_), .ZN(n8702) );
  INV_X1 U11067 ( .A(n8699), .ZN(n8700) );
  MUX2_X1 U11068 ( .A(n9646), .B(n9648), .S(n6411), .Z(n8704) );
  INV_X1 U11069 ( .A(SI_16_), .ZN(n9504) );
  NAND2_X1 U11070 ( .A1(n8704), .A2(n9504), .ZN(n8726) );
  INV_X1 U11071 ( .A(n8704), .ZN(n8705) );
  NAND2_X1 U11072 ( .A1(n8705), .A2(SI_16_), .ZN(n8706) );
  XNOR2_X1 U11073 ( .A(n8725), .B(n7555), .ZN(n11375) );
  NAND2_X1 U11074 ( .A1(n11375), .A2(n9005), .ZN(n8710) );
  OR2_X1 U11075 ( .A1(n8707), .A2(n13671), .ZN(n8708) );
  XNOR2_X1 U11076 ( .A(n8708), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U11077 ( .A1(n8772), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8771), 
        .B2(n13235), .ZN(n8709) );
  NAND2_X1 U11078 ( .A1(n14536), .A2(n9046), .ZN(n8720) );
  INV_X1 U11079 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8711) );
  AND2_X1 U11080 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  OR2_X1 U11081 ( .A1(n8713), .A2(n8738), .ZN(n14538) );
  INV_X1 U11082 ( .A(n14538), .ZN(n8714) );
  INV_X1 U11083 ( .A(n9017), .ZN(n8855) );
  NAND2_X1 U11084 ( .A1(n8714), .A2(n8855), .ZN(n8718) );
  NAND2_X1 U11085 ( .A1(n8980), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8717) );
  INV_X1 U11086 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13516) );
  OR2_X1 U11087 ( .A1(n6409), .A2(n13516), .ZN(n8716) );
  INV_X1 U11088 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n15228) );
  OR2_X1 U11089 ( .A1(n8361), .A2(n15228), .ZN(n8715) );
  NAND4_X1 U11090 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n13130) );
  NAND2_X1 U11091 ( .A1(n13130), .A2(n6426), .ZN(n8719) );
  NAND2_X1 U11092 ( .A1(n8720), .A2(n8719), .ZN(n8722) );
  AOI22_X1 U11093 ( .A1(n14536), .A2(n6426), .B1(n9046), .B2(n13130), .ZN(
        n8721) );
  AOI21_X1 U11094 ( .B1(n8723), .B2(n8722), .A(n8721), .ZN(n8724) );
  NAND2_X1 U11095 ( .A1(n8725), .A2(n7555), .ZN(n8727) );
  MUX2_X1 U11096 ( .A(n9721), .B(n9722), .S(n6411), .Z(n8728) );
  INV_X1 U11097 ( .A(SI_17_), .ZN(n9636) );
  NAND2_X1 U11098 ( .A1(n8728), .A2(n9636), .ZN(n8749) );
  INV_X1 U11099 ( .A(n8728), .ZN(n8729) );
  NAND2_X1 U11100 ( .A1(n8729), .A2(SI_17_), .ZN(n8730) );
  XNOR2_X1 U11101 ( .A(n8748), .B(n7545), .ZN(n11643) );
  NAND2_X1 U11102 ( .A1(n11643), .A2(n9005), .ZN(n8737) );
  NOR2_X1 U11103 ( .A1(n8731), .A2(n13671), .ZN(n8732) );
  MUX2_X1 U11104 ( .A(n13671), .B(n8732), .S(P2_IR_REG_17__SCAN_IN), .Z(n8735)
         );
  NAND2_X1 U11105 ( .A1(n8731), .A2(n8733), .ZN(n8751) );
  INV_X1 U11106 ( .A(n8751), .ZN(n8734) );
  NOR2_X1 U11107 ( .A1(n8735), .A2(n8734), .ZN(n14905) );
  AOI22_X1 U11108 ( .A1(n8772), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8771), 
        .B2(n14905), .ZN(n8736) );
  NAND2_X1 U11109 ( .A1(n13628), .A2(n6426), .ZN(n8745) );
  NAND2_X1 U11110 ( .A1(n8738), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8756) );
  OR2_X1 U11111 ( .A1(n8738), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11112 ( .A1(n8756), .A2(n8739), .ZN(n13492) );
  NAND2_X1 U11113 ( .A1(n9010), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8740) );
  OAI21_X1 U11114 ( .B1(n13492), .B2(n9017), .A(n8740), .ZN(n8743) );
  INV_X1 U11115 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U11116 ( .A1(n8964), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8741) );
  OAI21_X1 U11117 ( .B1(n13236), .B2(n9012), .A(n8741), .ZN(n8742) );
  NAND2_X1 U11118 ( .A1(n13129), .A2(n9046), .ZN(n8744) );
  NAND2_X1 U11119 ( .A1(n13628), .A2(n9046), .ZN(n8747) );
  NAND2_X1 U11120 ( .A1(n13129), .A2(n6426), .ZN(n8746) );
  MUX2_X1 U11121 ( .A(n10063), .B(n10060), .S(n6411), .Z(n8765) );
  XNOR2_X1 U11122 ( .A(n8767), .B(n8765), .ZN(n11631) );
  NAND2_X1 U11123 ( .A1(n11631), .A2(n9005), .ZN(n8754) );
  NAND2_X1 U11124 ( .A1(n8751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8752) );
  XNOR2_X1 U11125 ( .A(n8752), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U11126 ( .A1(n8772), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8771), 
        .B2(n13239), .ZN(n8753) );
  NAND2_X1 U11127 ( .A1(n13623), .A2(n9046), .ZN(n8761) );
  INV_X1 U11128 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11129 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U11130 ( .A1(n8776), .A2(n8757), .ZN(n13480) );
  AOI22_X1 U11131 ( .A1(n8980), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9010), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8759) );
  INV_X1 U11132 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13481) );
  OR2_X1 U11133 ( .A1(n6410), .A2(n13481), .ZN(n8758) );
  OAI211_X1 U11134 ( .C1(n13480), .C2(n9017), .A(n8759), .B(n8758), .ZN(n13128) );
  NAND2_X1 U11135 ( .A1(n13128), .A2(n6426), .ZN(n8760) );
  NAND2_X1 U11136 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  AOI22_X1 U11137 ( .A1(n13623), .A2(n6426), .B1(n9046), .B2(n13128), .ZN(
        n8762) );
  INV_X1 U11138 ( .A(n8765), .ZN(n8766) );
  MUX2_X1 U11139 ( .A(n10210), .B(n15215), .S(n6412), .Z(n8768) );
  NAND2_X1 U11140 ( .A1(n8768), .A2(n9750), .ZN(n8789) );
  INV_X1 U11141 ( .A(n8768), .ZN(n8769) );
  NAND2_X1 U11142 ( .A1(n8769), .A2(SI_19_), .ZN(n8770) );
  NAND2_X1 U11143 ( .A1(n8789), .A2(n8770), .ZN(n8787) );
  XNOR2_X1 U11144 ( .A(n8788), .B(n8787), .ZN(n11658) );
  NAND2_X1 U11145 ( .A1(n11658), .A2(n9005), .ZN(n8774) );
  AOI22_X1 U11146 ( .A1(n8772), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8318), 
        .B2(n8771), .ZN(n8773) );
  NAND2_X1 U11147 ( .A1(n13618), .A2(n6426), .ZN(n8781) );
  INV_X1 U11148 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8775) );
  AND2_X1 U11149 ( .A1(n8776), .A2(n8775), .ZN(n8777) );
  OR2_X1 U11150 ( .A1(n8777), .A2(n8814), .ZN(n13465) );
  AOI22_X1 U11151 ( .A1(n8980), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9010), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n8779) );
  INV_X1 U11152 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13469) );
  OR2_X1 U11153 ( .A1(n6410), .A2(n13469), .ZN(n8778) );
  OAI211_X1 U11154 ( .C1(n13465), .C2(n9017), .A(n8779), .B(n8778), .ZN(n13127) );
  NAND2_X1 U11155 ( .A1(n13127), .A2(n9046), .ZN(n8780) );
  NAND2_X1 U11156 ( .A1(n8781), .A2(n8780), .ZN(n8783) );
  AOI22_X1 U11157 ( .A1(n13618), .A2(n9046), .B1(n13127), .B2(n6426), .ZN(
        n8782) );
  NOR2_X1 U11158 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  INV_X1 U11159 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11681) );
  INV_X1 U11160 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10686) );
  MUX2_X1 U11161 ( .A(n11681), .B(n10686), .S(n6412), .Z(n8805) );
  XNOR2_X1 U11162 ( .A(n8807), .B(n8805), .ZN(n11680) );
  NAND2_X1 U11163 ( .A1(n11680), .A2(n9005), .ZN(n8791) );
  OR2_X1 U11164 ( .A1(n9007), .A2(n10686), .ZN(n8790) );
  NAND2_X1 U11165 ( .A1(n13449), .A2(n9046), .ZN(n8800) );
  INV_X1 U11166 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8792) );
  XNOR2_X1 U11167 ( .A(n8814), .B(n8792), .ZN(n13083) );
  NAND2_X1 U11168 ( .A1(n13083), .A2(n8855), .ZN(n8798) );
  INV_X1 U11169 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11170 ( .A1(n9010), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11171 ( .A1(n8964), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8793) );
  OAI211_X1 U11172 ( .C1(n9012), .C2(n8795), .A(n8794), .B(n8793), .ZN(n8796)
         );
  INV_X1 U11173 ( .A(n8796), .ZN(n8797) );
  NAND2_X1 U11174 ( .A1(n8798), .A2(n8797), .ZN(n13309) );
  NAND2_X1 U11175 ( .A1(n13309), .A2(n8842), .ZN(n8799) );
  NAND2_X1 U11176 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  INV_X1 U11177 ( .A(n13309), .ZN(n13307) );
  NAND2_X1 U11178 ( .A1(n13449), .A2(n8842), .ZN(n8803) );
  OAI21_X1 U11179 ( .B1(n13307), .B2(n8842), .A(n8803), .ZN(n8804) );
  INV_X1 U11180 ( .A(n8805), .ZN(n8806) );
  NAND2_X1 U11181 ( .A1(n8807), .A2(n8806), .ZN(n8810) );
  MUX2_X1 U11182 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6412), .Z(n8827) );
  XNOR2_X1 U11183 ( .A(n8827), .B(SI_21_), .ZN(n8824) );
  XNOR2_X1 U11184 ( .A(n8826), .B(n8824), .ZN(n11695) );
  NAND2_X1 U11185 ( .A1(n11695), .A2(n9005), .ZN(n8812) );
  OR2_X1 U11186 ( .A1(n9007), .A2(n15225), .ZN(n8811) );
  NAND2_X1 U11187 ( .A1(n13439), .A2(n6426), .ZN(n8822) );
  AND2_X1 U11188 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8813) );
  AOI21_X1 U11189 ( .B1(n8814), .B2(P2_REG3_REG_20__SCAN_IN), .A(
        P2_REG3_REG_21__SCAN_IN), .ZN(n8815) );
  OR2_X1 U11190 ( .A1(n8832), .A2(n8815), .ZN(n13442) );
  INV_X1 U11191 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11192 ( .A1(n9010), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11193 ( .A1(n8964), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8816) );
  OAI211_X1 U11194 ( .C1(n9012), .C2(n8818), .A(n8817), .B(n8816), .ZN(n8819)
         );
  INV_X1 U11195 ( .A(n8819), .ZN(n8820) );
  OAI21_X1 U11196 ( .B1(n13442), .B2(n9017), .A(n8820), .ZN(n13126) );
  NAND2_X1 U11197 ( .A1(n13126), .A2(n9046), .ZN(n8821) );
  AOI22_X1 U11198 ( .A1(n13439), .A2(n9046), .B1(n13126), .B2(n6426), .ZN(
        n8823) );
  INV_X1 U11199 ( .A(n8824), .ZN(n8825) );
  NAND2_X1 U11200 ( .A1(n8827), .A2(SI_21_), .ZN(n8828) );
  MUX2_X1 U11201 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6411), .Z(n8847) );
  XNOR2_X1 U11202 ( .A(n8846), .B(n8847), .ZN(n10945) );
  NAND2_X1 U11203 ( .A1(n10945), .A2(n9005), .ZN(n8831) );
  OR2_X1 U11204 ( .A1(n9007), .A2(n10948), .ZN(n8830) );
  NAND2_X1 U11205 ( .A1(n13598), .A2(n9046), .ZN(n8840) );
  NOR2_X1 U11206 ( .A1(n8832), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8833) );
  OR2_X1 U11207 ( .A1(n8853), .A2(n8833), .ZN(n13427) );
  INV_X1 U11208 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11209 ( .A1(n9010), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11210 ( .A1(n8964), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8834) );
  OAI211_X1 U11211 ( .C1(n9012), .C2(n8836), .A(n8835), .B(n8834), .ZN(n8837)
         );
  INV_X1 U11212 ( .A(n8837), .ZN(n8838) );
  OAI21_X1 U11213 ( .B1(n13427), .B2(n9017), .A(n8838), .ZN(n13125) );
  NAND2_X1 U11214 ( .A1(n13125), .A2(n8842), .ZN(n8839) );
  NAND2_X1 U11215 ( .A1(n8840), .A2(n8839), .ZN(n8844) );
  INV_X1 U11216 ( .A(n13125), .ZN(n13311) );
  NAND2_X1 U11217 ( .A1(n13598), .A2(n8842), .ZN(n8841) );
  OAI21_X1 U11218 ( .B1(n13311), .B2(n8842), .A(n8841), .ZN(n8843) );
  INV_X1 U11219 ( .A(n8844), .ZN(n8845) );
  INV_X1 U11220 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11726) );
  MUX2_X1 U11221 ( .A(n11726), .B(n11055), .S(n6412), .Z(n8864) );
  INV_X1 U11222 ( .A(n8864), .ZN(n8867) );
  XNOR2_X1 U11223 ( .A(n8867), .B(SI_23_), .ZN(n8850) );
  XNOR2_X1 U11224 ( .A(n8866), .B(n8850), .ZN(n11725) );
  NAND2_X1 U11225 ( .A1(n11725), .A2(n9005), .ZN(n8852) );
  OR2_X1 U11226 ( .A1(n9007), .A2(n11055), .ZN(n8851) );
  NAND2_X1 U11227 ( .A1(n13410), .A2(n6426), .ZN(n8863) );
  OR2_X1 U11228 ( .A1(n8853), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11229 ( .A1(n8853), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8874) );
  AND2_X1 U11230 ( .A1(n8854), .A2(n8874), .ZN(n13415) );
  NAND2_X1 U11231 ( .A1(n13415), .A2(n8855), .ZN(n8861) );
  INV_X1 U11232 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U11233 ( .A1(n9010), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U11234 ( .A1(n8964), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8856) );
  OAI211_X1 U11235 ( .C1(n9012), .C2(n8858), .A(n8857), .B(n8856), .ZN(n8859)
         );
  INV_X1 U11236 ( .A(n8859), .ZN(n8860) );
  NAND2_X1 U11237 ( .A1(n8861), .A2(n8860), .ZN(n13281) );
  NAND2_X1 U11238 ( .A1(n13281), .A2(n9046), .ZN(n8862) );
  NAND2_X1 U11239 ( .A1(n8863), .A2(n8862), .ZN(n8885) );
  NAND2_X1 U11240 ( .A1(n8864), .A2(n10713), .ZN(n8865) );
  NAND2_X1 U11241 ( .A1(n8867), .A2(SI_23_), .ZN(n8868) );
  MUX2_X1 U11242 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6411), .Z(n8887) );
  OR2_X1 U11243 ( .A1(n9007), .A2(n11237), .ZN(n8870) );
  NAND2_X1 U11244 ( .A1(n9010), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8880) );
  INV_X1 U11245 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8872) );
  OR2_X1 U11246 ( .A1(n9012), .A2(n8872), .ZN(n8879) );
  INV_X1 U11247 ( .A(n8874), .ZN(n8876) );
  INV_X1 U11248 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8873) );
  INV_X1 U11249 ( .A(n8913), .ZN(n8875) );
  OAI21_X1 U11250 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8876), .A(n8875), .ZN(
        n13397) );
  OR2_X1 U11251 ( .A1(n9017), .A2(n13397), .ZN(n8878) );
  INV_X1 U11252 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13398) );
  OR2_X1 U11253 ( .A1(n6410), .A2(n13398), .ZN(n8877) );
  NAND4_X1 U11254 ( .A1(n8880), .A2(n8879), .A3(n8878), .A4(n8877), .ZN(n13314) );
  AND2_X1 U11255 ( .A1(n13314), .A2(n6426), .ZN(n8881) );
  AOI21_X1 U11256 ( .B1(n13587), .B2(n9046), .A(n8881), .ZN(n8923) );
  NAND2_X1 U11257 ( .A1(n13587), .A2(n6426), .ZN(n8883) );
  NAND2_X1 U11258 ( .A1(n13314), .A2(n9046), .ZN(n8882) );
  NAND2_X1 U11259 ( .A1(n8883), .A2(n8882), .ZN(n8922) );
  AOI22_X1 U11260 ( .A1(n13410), .A2(n9046), .B1(n13281), .B2(n6426), .ZN(
        n8884) );
  MUX2_X1 U11261 ( .A(n11755), .B(n11363), .S(n6411), .Z(n8891) );
  NAND2_X1 U11262 ( .A1(n8891), .A2(n15313), .ZN(n8894) );
  INV_X1 U11263 ( .A(n8891), .ZN(n8892) );
  NAND2_X1 U11264 ( .A1(n8892), .A2(SI_25_), .ZN(n8893) );
  NAND2_X1 U11265 ( .A1(n8894), .A2(n8893), .ZN(n8907) );
  MUX2_X1 U11266 ( .A(n14321), .B(n13687), .S(n6412), .Z(n8931) );
  XNOR2_X1 U11267 ( .A(n8931), .B(SI_26_), .ZN(n8895) );
  OR2_X1 U11268 ( .A1(n9007), .A2(n13687), .ZN(n8896) );
  NAND2_X4 U11269 ( .A1(n8897), .A2(n8896), .ZN(n13373) );
  NAND2_X1 U11270 ( .A1(n9010), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8903) );
  INV_X1 U11271 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8898) );
  OR2_X1 U11272 ( .A1(n9012), .A2(n8898), .ZN(n8902) );
  NAND2_X1 U11273 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n8913), .ZN(n8912) );
  NAND2_X1 U11274 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8899), .ZN(n9014) );
  OAI21_X1 U11275 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8899), .A(n9014), .ZN(
        n13370) );
  OR2_X1 U11276 ( .A1(n9017), .A2(n13370), .ZN(n8901) );
  INV_X1 U11277 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13369) );
  OR2_X1 U11278 ( .A1(n6409), .A2(n13369), .ZN(n8900) );
  NAND4_X1 U11279 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n13318) );
  AND2_X1 U11280 ( .A1(n13318), .A2(n6426), .ZN(n8904) );
  AOI21_X1 U11281 ( .B1(n13373), .B2(n9046), .A(n8904), .ZN(n8995) );
  NAND2_X1 U11282 ( .A1(n13373), .A2(n6426), .ZN(n8906) );
  NAND2_X1 U11283 ( .A1(n13318), .A2(n9046), .ZN(n8905) );
  NAND2_X1 U11284 ( .A1(n8906), .A2(n8905), .ZN(n8996) );
  NAND2_X1 U11285 ( .A1(n11754), .A2(n9005), .ZN(n8910) );
  OR2_X1 U11286 ( .A1(n9007), .A2(n11363), .ZN(n8909) );
  NAND2_X1 U11287 ( .A1(n9010), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8918) );
  INV_X1 U11288 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8911) );
  OR2_X1 U11289 ( .A1(n9012), .A2(n8911), .ZN(n8917) );
  OAI21_X1 U11290 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8913), .A(n8912), .ZN(
        n13384) );
  OR2_X1 U11291 ( .A1(n9017), .A2(n13384), .ZN(n8916) );
  INV_X1 U11292 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8914) );
  OR2_X1 U11293 ( .A1(n6409), .A2(n8914), .ZN(n8915) );
  NAND4_X1 U11294 ( .A1(n8918), .A2(n8917), .A3(n8916), .A4(n8915), .ZN(n13316) );
  AND2_X1 U11295 ( .A1(n13316), .A2(n9046), .ZN(n8919) );
  AOI21_X1 U11296 ( .B1(n6879), .B2(n6426), .A(n8919), .ZN(n8994) );
  NAND2_X1 U11297 ( .A1(n6879), .A2(n9046), .ZN(n8921) );
  NAND2_X1 U11298 ( .A1(n13316), .A2(n6426), .ZN(n8920) );
  NAND2_X1 U11299 ( .A1(n8921), .A2(n8920), .ZN(n8993) );
  INV_X1 U11300 ( .A(n8922), .ZN(n8925) );
  INV_X1 U11301 ( .A(n8923), .ZN(n8924) );
  OAI22_X1 U11302 ( .A1(n8994), .A2(n8993), .B1(n8925), .B2(n8924), .ZN(n8926)
         );
  AOI21_X1 U11303 ( .B1(n8995), .B2(n8996), .A(n8926), .ZN(n8927) );
  INV_X1 U11304 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U11305 ( .A1(n8964), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11306 ( .A1(n9010), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8928) );
  OAI211_X1 U11307 ( .C1(n9012), .C2(n8930), .A(n8929), .B(n8928), .ZN(n13257)
         );
  MUX2_X1 U11308 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6412), .Z(n9001) );
  NOR2_X1 U11309 ( .A1(n9001), .A2(SI_27_), .ZN(n8933) );
  NAND2_X1 U11310 ( .A1(n9001), .A2(SI_27_), .ZN(n8934) );
  MUX2_X1 U11311 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6411), .Z(n8936) );
  XNOR2_X1 U11312 ( .A(n8936), .B(SI_28_), .ZN(n8975) );
  INV_X1 U11313 ( .A(n8936), .ZN(n8937) );
  NAND2_X1 U11314 ( .A1(n8937), .A2(n13000), .ZN(n8938) );
  INV_X1 U11315 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14312) );
  INV_X1 U11316 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13677) );
  MUX2_X1 U11317 ( .A(n14312), .B(n13677), .S(n6412), .Z(n8939) );
  XNOR2_X1 U11318 ( .A(n8939), .B(SI_29_), .ZN(n8960) );
  MUX2_X1 U11319 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6411), .Z(n8940) );
  MUX2_X1 U11320 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6412), .Z(n8941) );
  XNOR2_X1 U11321 ( .A(n8941), .B(SI_31_), .ZN(n8942) );
  NAND2_X1 U11322 ( .A1(n13669), .A2(n9005), .ZN(n8946) );
  INV_X1 U11323 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8944) );
  OR2_X1 U11324 ( .A1(n9007), .A2(n8944), .ZN(n8945) );
  MUX2_X1 U11325 ( .A(n13257), .B(n9046), .S(n9033), .Z(n8947) );
  NAND2_X1 U11326 ( .A1(n13257), .A2(n9046), .ZN(n9048) );
  NAND2_X1 U11327 ( .A1(n8947), .A2(n9048), .ZN(n8974) );
  NAND2_X1 U11328 ( .A1(n11834), .A2(n9005), .ZN(n8950) );
  INV_X1 U11329 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12000) );
  OR2_X1 U11330 ( .A1(n9007), .A2(n12000), .ZN(n8949) );
  NAND2_X1 U11331 ( .A1(n13257), .A2(n6426), .ZN(n8952) );
  NAND2_X1 U11332 ( .A1(n8951), .A2(n8318), .ZN(n14933) );
  OR2_X1 U11333 ( .A1(n14933), .A2(n10946), .ZN(n9103) );
  NAND2_X1 U11334 ( .A1(n8951), .A2(n10369), .ZN(n9769) );
  NAND4_X1 U11335 ( .A1(n8952), .A2(n9674), .A3(n9103), .A4(n9769), .ZN(n8956)
         );
  INV_X1 U11336 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11337 ( .A1(n8964), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11338 ( .A1(n9010), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U11339 ( .C1(n9012), .C2(n8955), .A(n8954), .B(n8953), .ZN(n13290)
         );
  AND2_X1 U11340 ( .A1(n8956), .A2(n13290), .ZN(n8957) );
  AOI21_X1 U11341 ( .B1(n13253), .B2(n9046), .A(n8957), .ZN(n9042) );
  NAND2_X1 U11342 ( .A1(n13253), .A2(n8842), .ZN(n8959) );
  NAND2_X1 U11343 ( .A1(n13290), .A2(n9046), .ZN(n8958) );
  NAND2_X1 U11344 ( .A1(n8959), .A2(n8958), .ZN(n9041) );
  NAND2_X1 U11345 ( .A1(n13675), .A2(n9005), .ZN(n8963) );
  OR2_X1 U11346 ( .A1(n9007), .A2(n13677), .ZN(n8962) );
  NAND2_X1 U11347 ( .A1(n8980), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11348 ( .A1(n8964), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8968) );
  INV_X1 U11349 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15341) );
  OR2_X1 U11350 ( .A1(n8361), .A2(n15341), .ZN(n8967) );
  INV_X1 U11351 ( .A(n9014), .ZN(n8965) );
  NAND2_X1 U11352 ( .A1(n8982), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13329) );
  OR2_X1 U11353 ( .A1(n9017), .A2(n13329), .ZN(n8966) );
  NAND4_X1 U11354 ( .A1(n8969), .A2(n8968), .A3(n8967), .A4(n8966), .ZN(n13123) );
  AND2_X1 U11355 ( .A1(n13123), .A2(n6426), .ZN(n8970) );
  AOI21_X1 U11356 ( .B1(n13555), .B2(n9046), .A(n8970), .ZN(n9039) );
  NAND2_X1 U11357 ( .A1(n13555), .A2(n8842), .ZN(n8972) );
  NAND2_X1 U11358 ( .A1(n13123), .A2(n9046), .ZN(n8971) );
  NAND2_X1 U11359 ( .A1(n8972), .A2(n8971), .ZN(n9038) );
  OAI22_X1 U11360 ( .A1(n9042), .A2(n9041), .B1(n9039), .B2(n9038), .ZN(n8973)
         );
  NAND2_X1 U11361 ( .A1(n8974), .A2(n8973), .ZN(n9044) );
  OR2_X1 U11362 ( .A1(n9007), .A2(n8977), .ZN(n8978) );
  NAND2_X1 U11363 ( .A1(n8980), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8988) );
  INV_X1 U11364 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8981) );
  OR2_X1 U11365 ( .A1(n8361), .A2(n8981), .ZN(n8987) );
  INV_X1 U11366 ( .A(n8982), .ZN(n9016) );
  INV_X1 U11367 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11368 ( .A1(n9016), .A2(n8983), .ZN(n8984) );
  NAND2_X1 U11369 ( .A1(n13329), .A2(n8984), .ZN(n13345) );
  OR2_X1 U11370 ( .A1(n9017), .A2(n13345), .ZN(n8986) );
  INV_X1 U11371 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13346) );
  OR2_X1 U11372 ( .A1(n6409), .A2(n13346), .ZN(n8985) );
  NAND4_X1 U11373 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n13124) );
  AND2_X1 U11374 ( .A1(n13124), .A2(n9046), .ZN(n8989) );
  AOI21_X1 U11375 ( .B1(n13558), .B2(n6426), .A(n8989), .ZN(n9035) );
  NAND2_X1 U11376 ( .A1(n13558), .A2(n9046), .ZN(n8991) );
  NAND2_X1 U11377 ( .A1(n13124), .A2(n6426), .ZN(n8990) );
  NAND2_X1 U11378 ( .A1(n8991), .A2(n8990), .ZN(n9034) );
  NAND2_X1 U11379 ( .A1(n9035), .A2(n9034), .ZN(n8992) );
  AND2_X1 U11380 ( .A1(n8994), .A2(n8993), .ZN(n8998) );
  INV_X1 U11381 ( .A(n8995), .ZN(n8997) );
  OR2_X1 U11382 ( .A1(n8998), .A2(n8997), .ZN(n9000) );
  INV_X1 U11383 ( .A(n8996), .ZN(n8999) );
  AOI22_X1 U11384 ( .A1(n9000), .A2(n8999), .B1(n8998), .B2(n8997), .ZN(n9027)
         );
  INV_X1 U11385 ( .A(n9001), .ZN(n9002) );
  XNOR2_X1 U11386 ( .A(n9002), .B(SI_27_), .ZN(n9003) );
  OR2_X1 U11387 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  NAND2_X1 U11388 ( .A1(n9010), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9022) );
  INV_X1 U11389 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9011) );
  OR2_X1 U11390 ( .A1(n9012), .A2(n9011), .ZN(n9021) );
  INV_X1 U11391 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U11392 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  NAND2_X1 U11393 ( .A1(n9016), .A2(n9015), .ZN(n13357) );
  OR2_X1 U11394 ( .A1(n9017), .A2(n13357), .ZN(n9020) );
  INV_X1 U11395 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9018) );
  OR2_X1 U11396 ( .A1(n6410), .A2(n9018), .ZN(n9019) );
  NAND4_X1 U11397 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n13286) );
  AND2_X1 U11398 ( .A1(n13286), .A2(n9046), .ZN(n9023) );
  AOI21_X1 U11399 ( .B1(n13568), .B2(n8842), .A(n9023), .ZN(n9029) );
  NAND2_X1 U11400 ( .A1(n13568), .A2(n9046), .ZN(n9025) );
  NAND2_X1 U11401 ( .A1(n13286), .A2(n8842), .ZN(n9024) );
  NAND2_X1 U11402 ( .A1(n9025), .A2(n9024), .ZN(n9030) );
  NAND2_X1 U11403 ( .A1(n9029), .A2(n9030), .ZN(n9026) );
  AND2_X1 U11404 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  INV_X1 U11405 ( .A(n9029), .ZN(n9032) );
  INV_X1 U11406 ( .A(n9030), .ZN(n9031) );
  XNOR2_X1 U11407 ( .A(n9033), .B(n13257), .ZN(n9071) );
  INV_X1 U11408 ( .A(n9034), .ZN(n9037) );
  INV_X1 U11409 ( .A(n9035), .ZN(n9036) );
  AOI22_X1 U11410 ( .A1(n9039), .A2(n9038), .B1(n9037), .B2(n9036), .ZN(n9040)
         );
  NAND2_X1 U11411 ( .A1(n9071), .A2(n9040), .ZN(n9043) );
  AOI22_X1 U11412 ( .A1(n9044), .A2(n9043), .B1(n9042), .B2(n9041), .ZN(n9045)
         );
  OR2_X1 U11413 ( .A1(n9046), .A2(n13257), .ZN(n9047) );
  MUX2_X1 U11414 ( .A(n9048), .B(n9047), .S(n9033), .Z(n9049) );
  INV_X1 U11415 ( .A(n13123), .ZN(n9050) );
  INV_X1 U11416 ( .A(n13314), .ZN(n13056) );
  XNOR2_X2 U11417 ( .A(n13587), .B(n13056), .ZN(n13395) );
  XNOR2_X1 U11418 ( .A(n13598), .B(n13311), .ZN(n13425) );
  OR2_X1 U11419 ( .A1(n13410), .A2(n13281), .ZN(n13313) );
  NAND2_X1 U11420 ( .A1(n13410), .A2(n13281), .ZN(n13312) );
  AND2_X1 U11421 ( .A1(n13313), .A2(n13312), .ZN(n13408) );
  INV_X1 U11422 ( .A(n13126), .ZN(n13310) );
  XNOR2_X1 U11423 ( .A(n13439), .B(n13310), .ZN(n13437) );
  XNOR2_X1 U11424 ( .A(n13449), .B(n13307), .ZN(n13276) );
  INV_X1 U11425 ( .A(n13128), .ZN(n13303) );
  XNOR2_X1 U11426 ( .A(n13623), .B(n13303), .ZN(n13302) );
  OR2_X1 U11427 ( .A1(n13618), .A2(n13127), .ZN(n13305) );
  NAND2_X1 U11428 ( .A1(n13618), .A2(n13127), .ZN(n13304) );
  NAND2_X1 U11429 ( .A1(n13305), .A2(n13304), .ZN(n13462) );
  XNOR2_X1 U11430 ( .A(n13628), .B(n13511), .ZN(n13503) );
  INV_X1 U11431 ( .A(n13130), .ZN(n13300) );
  XNOR2_X1 U11432 ( .A(n14536), .B(n13300), .ZN(n13514) );
  INV_X1 U11433 ( .A(n13134), .ZN(n11242) );
  XNOR2_X1 U11434 ( .A(n11243), .B(n11242), .ZN(n11178) );
  OR2_X1 U11435 ( .A1(n14795), .A2(n11413), .ZN(n11414) );
  NAND2_X1 U11436 ( .A1(n14795), .A2(n11413), .ZN(n11416) );
  NAND2_X1 U11437 ( .A1(n11414), .A2(n11416), .ZN(n11246) );
  INV_X1 U11438 ( .A(n13135), .ZN(n11176) );
  XNOR2_X1 U11439 ( .A(n15054), .B(n11176), .ZN(n11187) );
  XNOR2_X2 U11440 ( .A(n13145), .B(n9053), .ZN(n13540) );
  INV_X1 U11441 ( .A(n13539), .ZN(n9055) );
  NAND2_X1 U11442 ( .A1(n9055), .A2(n9054), .ZN(n14932) );
  NOR2_X1 U11443 ( .A1(n14932), .A2(n8951), .ZN(n9056) );
  NAND4_X1 U11444 ( .A1(n10152), .A2(n10609), .A3(n13540), .A4(n9056), .ZN(
        n9058) );
  INV_X1 U11445 ( .A(n13141), .ZN(n10442) );
  NAND2_X1 U11446 ( .A1(n10442), .A2(n15001), .ZN(n10723) );
  NAND2_X1 U11447 ( .A1(n13141), .A2(n7032), .ZN(n9057) );
  NAND2_X1 U11448 ( .A1(n10723), .A2(n9057), .ZN(n10395) );
  XNOR2_X1 U11449 ( .A(n13142), .B(n14995), .ZN(n10544) );
  NOR3_X1 U11450 ( .A1(n9058), .A2(n10395), .A3(n10544), .ZN(n9059) );
  XNOR2_X1 U11451 ( .A(n15029), .B(n13138), .ZN(n10921) );
  XNOR2_X1 U11452 ( .A(n15020), .B(n13139), .ZN(n10458) );
  XNOR2_X1 U11453 ( .A(n13140), .B(n10720), .ZN(n10722) );
  NAND4_X1 U11454 ( .A1(n9059), .A2(n10921), .A3(n10458), .A4(n10722), .ZN(
        n9060) );
  XNOR2_X1 U11455 ( .A(n13024), .B(n11172), .ZN(n11040) );
  INV_X1 U11456 ( .A(n13137), .ZN(n11033) );
  XNOR2_X1 U11457 ( .A(n15038), .B(n11033), .ZN(n10931) );
  OR4_X1 U11458 ( .A1(n11187), .A2(n9060), .A3(n11040), .A4(n10931), .ZN(n9061) );
  OR4_X1 U11459 ( .A1(n13514), .A2(n11178), .A3(n11246), .A4(n9061), .ZN(n9062) );
  NOR2_X1 U11460 ( .A1(n13503), .A2(n9062), .ZN(n9063) );
  XNOR2_X1 U11461 ( .A(n13640), .B(n13131), .ZN(n13295) );
  XNOR2_X1 U11462 ( .A(n11512), .B(n13132), .ZN(n11509) );
  NAND4_X1 U11463 ( .A1(n13462), .A2(n9063), .A3(n13295), .A4(n11509), .ZN(
        n9064) );
  OR4_X1 U11464 ( .A1(n13437), .A2(n13276), .A3(n13302), .A4(n9064), .ZN(n9065) );
  OR4_X1 U11465 ( .A1(n13395), .A2(n13425), .A3(n13408), .A4(n9065), .ZN(n9066) );
  NOR2_X1 U11466 ( .A1(n13379), .A2(n9066), .ZN(n9067) );
  NAND4_X1 U11467 ( .A1(n13323), .A2(n9067), .A3(n13321), .A4(n7216), .ZN(
        n9068) );
  NOR2_X1 U11468 ( .A1(n13325), .A2(n9068), .ZN(n9070) );
  XNOR2_X1 U11469 ( .A(n13253), .B(n13290), .ZN(n9069) );
  NAND3_X1 U11470 ( .A1(n9071), .A2(n9070), .A3(n9069), .ZN(n9072) );
  XNOR2_X1 U11471 ( .A(n9072), .B(n8318), .ZN(n9073) );
  INV_X1 U11472 ( .A(n9674), .ZN(n10674) );
  NAND2_X1 U11473 ( .A1(n9073), .A2(n10674), .ZN(n9104) );
  INV_X1 U11474 ( .A(n14933), .ZN(n9074) );
  NOR2_X1 U11475 ( .A1(n9104), .A2(n9074), .ZN(n9099) );
  INV_X1 U11476 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U11477 ( .A1(n9083), .A2(n9084), .ZN(n9079) );
  NAND2_X1 U11478 ( .A1(n9081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9076) );
  MUX2_X1 U11479 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9076), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9078) );
  NAND2_X1 U11480 ( .A1(n9078), .A2(n9077), .ZN(n13689) );
  NAND2_X1 U11481 ( .A1(n9079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9080) );
  MUX2_X1 U11482 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9080), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9082) );
  NAND2_X1 U11483 ( .A1(n9082), .A2(n9081), .ZN(n11361) );
  XNOR2_X1 U11484 ( .A(n9085), .B(n9084), .ZN(n11236) );
  OR2_X1 U11485 ( .A1(n11361), .A2(n11236), .ZN(n9086) );
  NOR2_X1 U11486 ( .A1(n13689), .A2(n9086), .ZN(n9661) );
  NAND2_X1 U11487 ( .A1(n9087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U11488 ( .A(n9089), .B(n9088), .ZN(n9095) );
  NAND2_X1 U11489 ( .A1(n9661), .A2(n9095), .ZN(n9092) );
  INV_X1 U11490 ( .A(n9095), .ZN(n9660) );
  NAND2_X1 U11491 ( .A1(n9649), .A2(n9674), .ZN(n10144) );
  OAI21_X1 U11492 ( .B1(n9660), .B2(n10144), .A(n9090), .ZN(n9091) );
  AND2_X1 U11493 ( .A1(n9092), .A2(n9091), .ZN(n9353) );
  OR2_X1 U11494 ( .A1(n9095), .A2(P2_U3088), .ZN(n11053) );
  OAI21_X1 U11495 ( .B1(n11053), .B2(n9649), .A(P2_B_REG_SCAN_IN), .ZN(n9096)
         );
  AOI21_X1 U11496 ( .B1(n14923), .B2(n7549), .A(n9096), .ZN(n9108) );
  OAI211_X1 U11497 ( .C1(n8318), .C2(n10674), .A(n9651), .B(n9769), .ZN(n9097)
         );
  OR2_X1 U11498 ( .A1(n9108), .A2(n9097), .ZN(n9098) );
  INV_X1 U11499 ( .A(n9108), .ZN(n9102) );
  INV_X1 U11500 ( .A(n8951), .ZN(n9100) );
  NAND3_X1 U11501 ( .A1(n9100), .A2(n8318), .A3(n9674), .ZN(n9101) );
  AND4_X1 U11502 ( .A1(n9104), .A2(n9103), .A3(n9102), .A4(n9101), .ZN(n9105)
         );
  NAND2_X1 U11503 ( .A1(n9106), .A2(n9105), .ZN(n9110) );
  INV_X1 U11504 ( .A(n11053), .ZN(n9107) );
  OR2_X1 U11505 ( .A1(n9108), .A2(n9107), .ZN(n9109) );
  INV_X1 U11506 ( .A(n9661), .ZN(n9112) );
  NOR3_X1 U11507 ( .A1(n9112), .A2(n9660), .A3(P2_U3088), .ZN(P2_U3947) );
  NOR2_X1 U11508 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9115) );
  NOR2_X1 U11509 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n9116) );
  INV_X2 U11510 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9239) );
  INV_X1 U11511 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9117) );
  INV_X1 U11512 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9119) );
  INV_X1 U11513 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9121) );
  INV_X1 U11514 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9122) );
  INV_X1 U11515 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9126) );
  INV_X1 U11516 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9123) );
  NAND2_X1 U11517 ( .A1(n6594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9127) );
  XNOR2_X1 U11518 ( .A(n9127), .B(n9126), .ZN(n10175) );
  AND2_X1 U11519 ( .A1(n10175), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9199) );
  INV_X1 U11520 ( .A(n9199), .ZN(n9202) );
  NOR2_X1 U11521 ( .A1(n9560), .A2(n9202), .ZN(P1_U4016) );
  OR2_X2 U11522 ( .A1(n12986), .A2(n9128), .ZN(n12521) );
  AND2_X1 U11523 ( .A1(n6412), .A2(P1_U3086), .ZN(n9207) );
  NOR2_X1 U11524 ( .A1(n6411), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14310) );
  NAND2_X1 U11525 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9129) );
  MUX2_X1 U11526 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9129), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9132) );
  INV_X1 U11527 ( .A(n9130), .ZN(n9131) );
  NAND2_X1 U11528 ( .A1(n9132), .A2(n9131), .ZN(n9587) );
  OAI222_X1 U11529 ( .A1(n6421), .A2(n9133), .B1(n11530), .B2(n9585), .C1(
        n9587), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U11530 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9159) );
  NOR2_X1 U11531 ( .A1(n9130), .A2(n9159), .ZN(n9134) );
  MUX2_X1 U11532 ( .A(n9159), .B(n9134), .S(P1_IR_REG_2__SCAN_IN), .Z(n9136)
         );
  INV_X1 U11533 ( .A(n9139), .ZN(n9135) );
  NOR2_X1 U11534 ( .A1(n9136), .A2(n9135), .ZN(n9606) );
  INV_X1 U11535 ( .A(n9606), .ZN(n13850) );
  INV_X1 U11536 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9137) );
  OAI222_X1 U11537 ( .A1(n13850), .A2(P1_U3086), .B1(n11530), .B2(n9604), .C1(
        n9137), .C2(n6421), .ZN(P1_U3353) );
  NOR2_X1 U11538 ( .A1(n6411), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13683) );
  INV_X1 U11539 ( .A(n13683), .ZN(n13686) );
  AND2_X1 U11540 ( .A1(n6412), .A2(P2_U3088), .ZN(n11052) );
  INV_X2 U11541 ( .A(n11052), .ZN(n13688) );
  OAI222_X1 U11542 ( .A1(n13686), .A2(n9138), .B1(n13688), .B2(n9604), .C1(
        P2_U3088), .C2(n13159), .ZN(P2_U3325) );
  NAND2_X1 U11543 ( .A1(n9139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9140) );
  XNOR2_X1 U11544 ( .A(n9140), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13863) );
  INV_X1 U11545 ( .A(n13863), .ZN(n9142) );
  OAI222_X1 U11546 ( .A1(n9142), .A2(P1_U3086), .B1(n11530), .B2(n9926), .C1(
        n9141), .C2(n6421), .ZN(P1_U3352) );
  OAI222_X1 U11547 ( .A1(n13686), .A2(n9143), .B1(n13688), .B2(n9926), .C1(
        P2_U3088), .C2(n13174), .ZN(P2_U3324) );
  NOR2_X1 U11548 ( .A1(n6412), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14446) );
  INV_X1 U11549 ( .A(n14446), .ZN(n14451) );
  MUX2_X1 U11550 ( .A(n9144), .B(n15268), .S(P3_STATE_REG_SCAN_IN), .Z(n9145)
         );
  OAI21_X1 U11551 ( .B1(n9146), .B2(n14451), .A(n9145), .ZN(P3_U3295) );
  OAI222_X1 U11552 ( .A1(n13686), .A2(n9147), .B1(n13688), .B2(n9930), .C1(
        P2_U3088), .C2(n14809), .ZN(P2_U3323) );
  OAI222_X1 U11553 ( .A1(P3_U3151), .A2(n10335), .B1(n12997), .B2(n9149), .C1(
        n14451), .C2(n9148), .ZN(P3_U3287) );
  OAI222_X1 U11554 ( .A1(n14451), .A2(n9151), .B1(n12997), .B2(n9150), .C1(
        P3_U3151), .C2(n10050), .ZN(P3_U3294) );
  CLKBUF_X1 U11555 ( .A(n13686), .Z(n11238) );
  OAI222_X1 U11556 ( .A1(n11238), .A2(n9152), .B1(n13688), .B2(n9585), .C1(
        P2_U3088), .C2(n13151), .ZN(P2_U3326) );
  OAI222_X1 U11557 ( .A1(n10004), .A2(P3_U3151), .B1(n14451), .B2(n9154), .C1(
        n9153), .C2(n12997), .ZN(P3_U3289) );
  OAI222_X1 U11558 ( .A1(P3_U3151), .A2(n15095), .B1(n12997), .B2(n9156), .C1(
        n14451), .C2(n9155), .ZN(P3_U3285) );
  NOR2_X1 U11559 ( .A1(n9157), .A2(n9159), .ZN(n9158) );
  MUX2_X1 U11560 ( .A(n9159), .B(n9158), .S(P1_IR_REG_5__SCAN_IN), .Z(n9161)
         );
  OR2_X1 U11561 ( .A1(n9161), .A2(n9237), .ZN(n13898) );
  INV_X1 U11562 ( .A(n9940), .ZN(n9163) );
  INV_X1 U11563 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9162) );
  OAI222_X1 U11564 ( .A1(n13898), .A2(P1_U3086), .B1(n11530), .B2(n9163), .C1(
        n9162), .C2(n6421), .ZN(P1_U3350) );
  INV_X1 U11565 ( .A(n14819), .ZN(n14827) );
  OAI222_X1 U11566 ( .A1(n13686), .A2(n9164), .B1(n13688), .B2(n9163), .C1(
        P2_U3088), .C2(n14827), .ZN(P2_U3322) );
  INV_X1 U11567 ( .A(n12997), .ZN(n14445) );
  AOI222_X1 U11568 ( .A1(n9165), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10005), .C1(SI_2_), .C2(n14445), .ZN(n9166) );
  INV_X1 U11569 ( .A(n9166), .ZN(P3_U3293) );
  AOI222_X1 U11570 ( .A1(n9167), .A2(n14446), .B1(n9894), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_7_), .C2(n14445), .ZN(n9168) );
  INV_X1 U11571 ( .A(n9168), .ZN(P3_U3288) );
  AOI222_X1 U11572 ( .A1(n9169), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9814), .C1(SI_3_), .C2(n14445), .ZN(n9170) );
  INV_X1 U11573 ( .A(n9170), .ZN(P3_U3292) );
  AOI222_X1 U11574 ( .A1(n9171), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9831), .C1(SI_5_), .C2(n14445), .ZN(n9172) );
  INV_X1 U11575 ( .A(n9172), .ZN(P3_U3290) );
  AOI222_X1 U11576 ( .A1(n9173), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9860), .C1(SI_4_), .C2(n14445), .ZN(n9174) );
  INV_X1 U11577 ( .A(n9174), .ZN(P3_U3291) );
  OR2_X1 U11578 ( .A1(n9237), .A2(n9159), .ZN(n9175) );
  XNOR2_X1 U11579 ( .A(n9175), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10074) );
  INV_X1 U11580 ( .A(n10074), .ZN(n9177) );
  INV_X1 U11581 ( .A(n10073), .ZN(n9178) );
  OAI222_X1 U11582 ( .A1(n9177), .A2(P1_U3086), .B1(n11530), .B2(n9178), .C1(
        n9176), .C2(n6421), .ZN(P1_U3349) );
  OAI222_X1 U11583 ( .A1(n13686), .A2(n9179), .B1(n13688), .B2(n9178), .C1(
        P2_U3088), .C2(n13188), .ZN(P2_U3321) );
  NAND2_X1 U11584 ( .A1(n9224), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U11585 ( .A(n9180), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13880) );
  INV_X1 U11586 ( .A(n13880), .ZN(n9314) );
  OAI222_X1 U11587 ( .A1(n9314), .A2(P1_U3086), .B1(n11530), .B2(n9930), .C1(
        n9181), .C2(n6421), .ZN(P1_U3351) );
  NAND2_X1 U11588 ( .A1(n9237), .A2(n9239), .ZN(n9186) );
  NAND2_X1 U11589 ( .A1(n9186), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9182) );
  XNOR2_X1 U11590 ( .A(n9182), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10079) );
  INV_X1 U11591 ( .A(n10079), .ZN(n9501) );
  INV_X1 U11592 ( .A(n10078), .ZN(n9184) );
  OAI222_X1 U11593 ( .A1(n9501), .A2(P1_U3086), .B1(n11530), .B2(n9184), .C1(
        n9183), .C2(n6421), .ZN(P1_U3348) );
  INV_X1 U11594 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9185) );
  INV_X1 U11595 ( .A(n9545), .ZN(n9375) );
  OAI222_X1 U11596 ( .A1(n11238), .A2(n9185), .B1(n13688), .B2(n9184), .C1(
        P2_U3088), .C2(n9375), .ZN(P2_U3320) );
  INV_X1 U11597 ( .A(n10273), .ZN(n9193) );
  NAND2_X1 U11598 ( .A1(n9643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9187) );
  XNOR2_X1 U11599 ( .A(n9187), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U11600 ( .A1(n10274), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9207), .ZN(n9188) );
  OAI21_X1 U11601 ( .B1(n9193), .B2(n11530), .A(n9188), .ZN(P1_U3347) );
  INV_X1 U11602 ( .A(n9189), .ZN(n9190) );
  OAI222_X1 U11603 ( .A1(P3_U3151), .A2(n15123), .B1(n12997), .B2(n9191), .C1(
        n14451), .C2(n9190), .ZN(P3_U3283) );
  INV_X1 U11604 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9194) );
  INV_X1 U11605 ( .A(n13203), .ZN(n9192) );
  OAI222_X1 U11606 ( .A1(n11238), .A2(n9194), .B1(n13688), .B2(n9193), .C1(
        P2_U3088), .C2(n9192), .ZN(P2_U3319) );
  INV_X1 U11607 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9195) );
  INV_X1 U11608 ( .A(n10555), .ZN(n9198) );
  INV_X1 U11609 ( .A(n9550), .ZN(n14842) );
  OAI222_X1 U11610 ( .A1(n11238), .A2(n9195), .B1(n13688), .B2(n9198), .C1(
        P2_U3088), .C2(n14842), .ZN(P2_U3318) );
  NAND2_X1 U11611 ( .A1(n9196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11612 ( .A(n9214), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10556) );
  INV_X1 U11613 ( .A(n10556), .ZN(n9389) );
  OAI222_X1 U11614 ( .A1(n9389), .A2(P1_U3086), .B1(n11530), .B2(n9198), .C1(
        n9197), .C2(n6421), .ZN(P1_U3346) );
  NAND2_X1 U11615 ( .A1(n11532), .A2(P1_B_REG_SCAN_IN), .ZN(n9201) );
  INV_X1 U11616 ( .A(P1_B_REG_SCAN_IN), .ZN(n13923) );
  NAND2_X1 U11617 ( .A1(n9258), .A2(n13923), .ZN(n9200) );
  OAI211_X1 U11618 ( .C1(n9262), .C2(n9201), .A(n14320), .B(n9200), .ZN(n9261)
         );
  INV_X1 U11620 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9203) );
  NOR2_X1 U11621 ( .A1(n14320), .A2(n9202), .ZN(n11533) );
  INV_X1 U11622 ( .A(n9262), .ZN(n11360) );
  AOI22_X1 U11623 ( .A1(n6405), .A2(n9203), .B1(n11533), .B2(n11360), .ZN(
        P1_U3446) );
  INV_X1 U11624 ( .A(n10560), .ZN(n9210) );
  INV_X1 U11625 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U11626 ( .A1(n9214), .A2(n9204), .ZN(n9205) );
  NAND2_X1 U11627 ( .A1(n9205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9206) );
  XNOR2_X1 U11628 ( .A(n9206), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U11629 ( .A1(n10561), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9207), .ZN(n9208) );
  OAI21_X1 U11630 ( .B1(n9210), .B2(n11530), .A(n9208), .ZN(P1_U3345) );
  INV_X1 U11631 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n15344) );
  INV_X1 U11632 ( .A(n14848), .ZN(n9209) );
  OAI222_X1 U11633 ( .A1(n11238), .A2(n15344), .B1(n13688), .B2(n9210), .C1(
        P2_U3088), .C2(n9209), .ZN(P2_U3317) );
  INV_X1 U11634 ( .A(n10573), .ZN(n9215) );
  INV_X1 U11635 ( .A(n9975), .ZN(n9544) );
  OAI222_X1 U11636 ( .A1(n11238), .A2(n9211), .B1(n13688), .B2(n9215), .C1(
        P2_U3088), .C2(n9544), .ZN(P2_U3316) );
  OR2_X1 U11637 ( .A1(n9212), .A2(n9159), .ZN(n9213) );
  NAND2_X1 U11638 ( .A1(n9214), .A2(n9213), .ZN(n9377) );
  XNOR2_X1 U11639 ( .A(n9377), .B(n9639), .ZN(n10574) );
  INV_X1 U11640 ( .A(n10574), .ZN(n9509) );
  OAI222_X1 U11641 ( .A1(n6421), .A2(n9216), .B1(n11530), .B2(n9215), .C1(
        P1_U3086), .C2(n9509), .ZN(P1_U3344) );
  OAI222_X1 U11642 ( .A1(n12530), .A2(P3_U3151), .B1(n14451), .B2(n9218), .C1(
        n9217), .C2(n12997), .ZN(P3_U3281) );
  INV_X1 U11643 ( .A(n9580), .ZN(n9568) );
  INV_X1 U11644 ( .A(n10175), .ZN(n9219) );
  NAND2_X1 U11645 ( .A1(n9219), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11918) );
  NAND2_X1 U11646 ( .A1(n9568), .A2(n11918), .ZN(n9308) );
  NAND2_X1 U11647 ( .A1(n6831), .A2(n9281), .ZN(n11862) );
  INV_X1 U11648 ( .A(n11862), .ZN(n9572) );
  INV_X1 U11649 ( .A(n9224), .ZN(n9230) );
  NOR2_X1 U11650 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9228) );
  NOR2_X1 U11651 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9227) );
  NOR2_X1 U11652 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9226) );
  NOR2_X1 U11653 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9225) );
  INV_X1 U11654 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9232) );
  AOI21_X1 U11656 ( .B1(n9572), .B2(n10175), .A(n11659), .ZN(n9307) );
  INV_X1 U11657 ( .A(n9307), .ZN(n9234) );
  AND2_X1 U11658 ( .A1(n9308), .A2(n9234), .ZN(n14655) );
  CLKBUF_X2 U11659 ( .A(P1_U4016), .Z(n13844) );
  NOR2_X1 U11660 ( .A1(n14655), .A2(n13844), .ZN(P1_U3085) );
  INV_X1 U11661 ( .A(n9235), .ZN(n9244) );
  NAND2_X1 U11662 ( .A1(n9244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9236) );
  INV_X1 U11663 ( .A(n9237), .ZN(n9243) );
  NAND3_X1 U11664 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(n9242) );
  XNOR2_X1 U11665 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_19__SCAN_IN), .ZN(
        n9241) );
  NAND2_X1 U11666 ( .A1(n9245), .A2(n9244), .ZN(n14471) );
  AND2_X1 U11667 ( .A1(n11860), .A2(n14471), .ZN(n9246) );
  OR2_X1 U11668 ( .A1(n11862), .A2(n9246), .ZN(n10176) );
  NAND2_X1 U11669 ( .A1(n9580), .A2(n10176), .ZN(n9576) );
  NOR4_X1 U11670 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9255) );
  NOR4_X1 U11671 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9254) );
  OR4_X1 U11672 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9252) );
  NOR4_X1 U11673 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9250) );
  NOR4_X1 U11674 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9249) );
  NOR4_X1 U11675 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9248) );
  NOR4_X1 U11676 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9247) );
  NAND4_X1 U11677 ( .A1(n9250), .A2(n9249), .A3(n9248), .A4(n9247), .ZN(n9251)
         );
  NOR4_X1 U11678 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9252), .A4(n9251), .ZN(n9253) );
  AND3_X1 U11679 ( .A1(n9255), .A2(n9254), .A3(n9253), .ZN(n9256) );
  OR2_X1 U11680 ( .A1(n9261), .A2(n9256), .ZN(n9559) );
  INV_X1 U11681 ( .A(n9559), .ZN(n9257) );
  NOR2_X1 U11682 ( .A1(n9576), .A2(n9257), .ZN(n9686) );
  OR2_X1 U11683 ( .A1(n9261), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9260) );
  OR2_X1 U11684 ( .A1(n9258), .A2(n14320), .ZN(n9259) );
  INV_X1 U11685 ( .A(n14471), .ZN(n14184) );
  INV_X1 U11686 ( .A(n9687), .ZN(n9574) );
  AND2_X1 U11687 ( .A1(n9684), .A2(n9574), .ZN(n9266) );
  OR2_X1 U11688 ( .A1(n9261), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9264) );
  OR2_X1 U11689 ( .A1(n14320), .A2(n9262), .ZN(n9263) );
  INV_X1 U11690 ( .A(n13966), .ZN(n9265) );
  AND3_X2 U11691 ( .A1(n9686), .A2(n9266), .A3(n9265), .ZN(n14772) );
  INV_X1 U11692 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9478) );
  INV_X1 U11693 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13842) );
  INV_X1 U11694 ( .A(SI_0_), .ZN(n15326) );
  OAI21_X1 U11695 ( .B1(n6412), .B2(n15326), .A(n9267), .ZN(n9268) );
  NAND2_X1 U11696 ( .A1(n9269), .A2(n9268), .ZN(n14327) );
  INV_X1 U11697 ( .A(n6424), .ZN(n13841) );
  OR2_X1 U11698 ( .A1(n11862), .A2(n13841), .ZN(n11394) );
  INV_X2 U11699 ( .A(n11394), .ZN(n14575) );
  NAND2_X1 U11700 ( .A1(n9272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9273) );
  INV_X1 U11701 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9274) );
  OR2_X1 U11702 ( .A1(n9944), .A2(n9274), .ZN(n9279) );
  INV_X1 U11703 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9910) );
  INV_X1 U11704 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9309) );
  INV_X1 U11705 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U11706 ( .A1(n6831), .A2(n14184), .ZN(n9280) );
  NAND2_X1 U11707 ( .A1(n9281), .A2(n11869), .ZN(n11536) );
  INV_X1 U11708 ( .A(n14751), .ZN(n14570) );
  NAND2_X1 U11709 ( .A1(n14326), .A2(n14471), .ZN(n9282) );
  NAND2_X1 U11710 ( .A1(n11541), .A2(n6831), .ZN(n9283) );
  NAND2_X1 U11711 ( .A1(n12130), .A2(n9283), .ZN(n14609) );
  INV_X1 U11712 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9284) );
  INV_X1 U11713 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11714 ( .A1(n13838), .A2(n9584), .ZN(n9905) );
  OR2_X1 U11715 ( .A1(n13838), .A2(n9584), .ZN(n9286) );
  NAND2_X1 U11716 ( .A1(n9905), .A2(n9286), .ZN(n11876) );
  AOI21_X1 U11717 ( .B1(n14570), .B2(n14609), .A(n11876), .ZN(n9287) );
  AOI21_X1 U11718 ( .B1(n14575), .B2(n13837), .A(n9287), .ZN(n10227) );
  OAI21_X1 U11719 ( .B1(n9906), .B2(n9569), .A(n10227), .ZN(n9689) );
  NAND2_X1 U11720 ( .A1(n14772), .A2(n9689), .ZN(n9288) );
  OAI21_X1 U11721 ( .B1(n14772), .B2(n9478), .A(n9288), .ZN(P1_U3528) );
  INV_X1 U11722 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9599) );
  MUX2_X1 U11723 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9599), .S(n9606), .Z(n13847) );
  MUX2_X1 U11724 ( .A(n9289), .B(P1_REG1_REG_1__SCAN_IN), .S(n9587), .Z(n9291)
         );
  AND2_X1 U11725 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9290) );
  NAND2_X1 U11726 ( .A1(n9291), .A2(n9290), .ZN(n9480) );
  OAI21_X1 U11727 ( .B1(n9289), .B2(n9587), .A(n9480), .ZN(n13846) );
  NAND2_X1 U11728 ( .A1(n13847), .A2(n13846), .ZN(n13866) );
  NAND2_X1 U11729 ( .A1(n9606), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13865) );
  NAND2_X1 U11730 ( .A1(n13866), .A2(n13865), .ZN(n9293) );
  INV_X1 U11731 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U11732 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9611), .S(n13863), .Z(n9292) );
  NAND2_X1 U11733 ( .A1(n9293), .A2(n9292), .ZN(n13883) );
  NAND2_X1 U11734 ( .A1(n13863), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13882) );
  NAND2_X1 U11735 ( .A1(n13883), .A2(n13882), .ZN(n9295) );
  INV_X1 U11736 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U11737 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9933), .S(n13880), .Z(n9294) );
  NAND2_X1 U11738 ( .A1(n9295), .A2(n9294), .ZN(n13885) );
  NAND2_X1 U11739 ( .A1(n13880), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9296) );
  AND2_X1 U11740 ( .A1(n13885), .A2(n9296), .ZN(n13894) );
  INV_X1 U11741 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9967) );
  MUX2_X1 U11742 ( .A(n9967), .B(P1_REG1_REG_5__SCAN_IN), .S(n13898), .Z(
        n13895) );
  NAND2_X1 U11743 ( .A1(n13894), .A2(n13895), .ZN(n13893) );
  NAND2_X1 U11744 ( .A1(n13898), .A2(n9967), .ZN(n9297) );
  NAND2_X1 U11745 ( .A1(n13893), .A2(n9297), .ZN(n9457) );
  INV_X1 U11746 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U11747 ( .A(n10135), .B(P1_REG1_REG_6__SCAN_IN), .S(n10074), .Z(
        n9456) );
  OR2_X1 U11748 ( .A1(n9457), .A2(n9456), .ZN(n9491) );
  NAND2_X1 U11749 ( .A1(n10074), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11750 ( .A1(n9491), .A2(n9490), .ZN(n9300) );
  INV_X1 U11751 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9298) );
  MUX2_X1 U11752 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9298), .S(n10079), .Z(n9299) );
  NAND2_X1 U11753 ( .A1(n9300), .A2(n9299), .ZN(n9493) );
  NAND2_X1 U11754 ( .A1(n10079), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9301) );
  AND2_X1 U11755 ( .A1(n9493), .A2(n9301), .ZN(n9523) );
  MUX2_X1 U11756 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10094), .S(n10274), .Z(
        n9524) );
  NAND2_X1 U11757 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  OR2_X1 U11758 ( .A1(n10274), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11759 ( .A1(n9522), .A2(n9304), .ZN(n9302) );
  INV_X1 U11760 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15311) );
  MUX2_X1 U11761 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15311), .S(n10556), .Z(
        n9303) );
  NAND2_X1 U11762 ( .A1(n9302), .A2(n9303), .ZN(n9391) );
  INV_X1 U11763 ( .A(n9303), .ZN(n9305) );
  NAND3_X1 U11764 ( .A1(n9522), .A2(n9305), .A3(n9304), .ZN(n9306) );
  AND2_X1 U11765 ( .A1(n9391), .A2(n9306), .ZN(n9327) );
  NAND2_X1 U11766 ( .A1(n9308), .A2(n9307), .ZN(n14657) );
  INV_X1 U11767 ( .A(n14653), .ZN(n11914) );
  OR2_X1 U11768 ( .A1(n14657), .A2(n11914), .ZN(n14669) );
  INV_X1 U11769 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9598) );
  MUX2_X1 U11770 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9598), .S(n9606), .Z(n13853) );
  MUX2_X1 U11771 ( .A(n9309), .B(P1_REG2_REG_1__SCAN_IN), .S(n9587), .Z(n9310)
         );
  AND2_X1 U11772 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9473) );
  NAND2_X1 U11773 ( .A1(n9310), .A2(n9473), .ZN(n9474) );
  OAI21_X1 U11774 ( .B1(n9309), .B2(n9587), .A(n9474), .ZN(n13852) );
  NAND2_X1 U11775 ( .A1(n13853), .A2(n13852), .ZN(n13861) );
  NAND2_X1 U11776 ( .A1(n9606), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U11777 ( .A1(n13861), .A2(n13860), .ZN(n9312) );
  INV_X1 U11778 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14699) );
  MUX2_X1 U11779 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14699), .S(n13863), .Z(
        n9311) );
  NAND2_X1 U11780 ( .A1(n9312), .A2(n9311), .ZN(n13876) );
  NAND2_X1 U11781 ( .A1(n13863), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13875) );
  INV_X1 U11782 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9313) );
  MUX2_X1 U11783 ( .A(n9313), .B(P1_REG2_REG_4__SCAN_IN), .S(n13880), .Z(
        n13874) );
  AOI21_X1 U11784 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(n13873) );
  NOR2_X1 U11785 ( .A1(n9314), .A2(n9313), .ZN(n13897) );
  INV_X1 U11786 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U11787 ( .A(n9946), .B(P1_REG2_REG_5__SCAN_IN), .S(n13898), .Z(n9315) );
  OAI21_X1 U11788 ( .B1(n13873), .B2(n13897), .A(n9315), .ZN(n13903) );
  INV_X1 U11789 ( .A(n13898), .ZN(n13892) );
  NAND2_X1 U11790 ( .A1(n13892), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9459) );
  INV_X1 U11791 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9316) );
  MUX2_X1 U11792 ( .A(n9316), .B(P1_REG2_REG_6__SCAN_IN), .S(n10074), .Z(n9458) );
  AOI21_X1 U11793 ( .B1(n13903), .B2(n9459), .A(n9458), .ZN(n9461) );
  AOI21_X1 U11794 ( .B1(n10074), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9461), .ZN(
        n9495) );
  INV_X1 U11795 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9317) );
  MUX2_X1 U11796 ( .A(n9317), .B(P1_REG2_REG_7__SCAN_IN), .S(n10079), .Z(n9494) );
  NOR2_X1 U11797 ( .A1(n9495), .A2(n9494), .ZN(n9529) );
  NOR2_X1 U11798 ( .A1(n9501), .A2(n9317), .ZN(n9528) );
  INV_X1 U11799 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U11800 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10097), .S(n10274), .Z(
        n9527) );
  OAI21_X1 U11801 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9526) );
  NAND2_X1 U11802 ( .A1(n10274), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9321) );
  INV_X1 U11803 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9318) );
  MUX2_X1 U11804 ( .A(n9318), .B(P1_REG2_REG_9__SCAN_IN), .S(n10556), .Z(n9320) );
  AOI21_X1 U11805 ( .B1(n9526), .B2(n9321), .A(n9320), .ZN(n9404) );
  INV_X1 U11806 ( .A(n9404), .ZN(n9323) );
  OR2_X1 U11807 ( .A1(n6424), .A2(n6415), .ZN(n9319) );
  OR2_X1 U11808 ( .A1(n14657), .A2(n9319), .ZN(n14663) );
  INV_X1 U11809 ( .A(n14663), .ZN(n13914) );
  NAND3_X1 U11810 ( .A1(n9526), .A2(n9321), .A3(n9320), .ZN(n9322) );
  NAND3_X1 U11811 ( .A1(n9323), .A2(n13914), .A3(n9322), .ZN(n9326) );
  OR2_X1 U11812 ( .A1(n14657), .A2(n13841), .ZN(n13849) );
  INV_X1 U11813 ( .A(n13849), .ZN(n14666) );
  INV_X1 U11814 ( .A(n14655), .ZN(n14674) );
  INV_X1 U11815 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U11816 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11126) );
  OAI21_X1 U11817 ( .B1(n14674), .B2(n14350), .A(n11126), .ZN(n9324) );
  AOI21_X1 U11818 ( .B1(n10556), .B2(n14666), .A(n9324), .ZN(n9325) );
  OAI211_X1 U11819 ( .C1(n9327), .C2(n14669), .A(n9326), .B(n9325), .ZN(
        P1_U3252) );
  NAND2_X1 U11820 ( .A1(n6427), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9328) );
  OR2_X1 U11821 ( .A1(n9353), .A2(n9328), .ZN(n14930) );
  NAND2_X1 U11822 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10768) );
  INV_X1 U11823 ( .A(n10768), .ZN(n9351) );
  INV_X1 U11824 ( .A(n6427), .ZN(n9329) );
  NOR2_X1 U11825 ( .A1(n9094), .A2(P2_U3088), .ZN(n13682) );
  NAND2_X1 U11826 ( .A1(n9329), .A2(n13682), .ZN(n9330) );
  OR2_X1 U11827 ( .A1(n9353), .A2(n9330), .ZN(n14853) );
  MUX2_X1 U11828 ( .A(n9331), .B(P2_REG2_REG_2__SCAN_IN), .S(n13159), .Z(
        n13162) );
  AND2_X1 U11829 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9332) );
  OAI21_X1 U11830 ( .B1(n13545), .B2(n13151), .A(n13154), .ZN(n13161) );
  OR2_X1 U11831 ( .A1(n13159), .A2(n9331), .ZN(n13171) );
  NAND2_X1 U11832 ( .A1(n13172), .A2(n13171), .ZN(n9335) );
  MUX2_X1 U11833 ( .A(n9333), .B(P2_REG2_REG_3__SCAN_IN), .S(n13174), .Z(n9334) );
  NAND2_X1 U11834 ( .A1(n9335), .A2(n9334), .ZN(n14801) );
  INV_X1 U11835 ( .A(n13174), .ZN(n13169) );
  NAND2_X1 U11836 ( .A1(n13169), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U11837 ( .A1(n14801), .A2(n14800), .ZN(n9338) );
  MUX2_X1 U11838 ( .A(n9336), .B(P2_REG2_REG_4__SCAN_IN), .S(n14809), .Z(n9337) );
  OR2_X1 U11839 ( .A1(n14809), .A2(n9336), .ZN(n14815) );
  NAND2_X1 U11840 ( .A1(n14816), .A2(n14815), .ZN(n9340) );
  MUX2_X1 U11841 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10402), .S(n14819), .Z(
        n9339) );
  NAND2_X1 U11842 ( .A1(n9340), .A2(n9339), .ZN(n14818) );
  NAND2_X1 U11843 ( .A1(n14819), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U11844 ( .A1(n14818), .A2(n13190), .ZN(n9343) );
  MUX2_X1 U11845 ( .A(n9341), .B(P2_REG2_REG_6__SCAN_IN), .S(n13188), .Z(n9342) );
  NAND2_X1 U11846 ( .A1(n13183), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11847 ( .A1(n13192), .A2(n9348), .ZN(n9346) );
  MUX2_X1 U11848 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9344), .S(n9545), .Z(n9345)
         );
  NAND2_X1 U11849 ( .A1(n9346), .A2(n9345), .ZN(n13200) );
  MUX2_X1 U11850 ( .A(n9344), .B(P2_REG2_REG_7__SCAN_IN), .S(n9545), .Z(n9347)
         );
  NAND3_X1 U11851 ( .A1(n13192), .A2(n9348), .A3(n9347), .ZN(n9349) );
  AND3_X1 U11852 ( .A1(n14917), .A2(n13200), .A3(n9349), .ZN(n9350) );
  AOI211_X1 U11853 ( .C1(n14923), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n9351), .B(
        n9350), .ZN(n9374) );
  NOR2_X1 U11854 ( .A1(n6427), .A2(P2_U3088), .ZN(n13679) );
  NAND2_X1 U11855 ( .A1(n13679), .A2(n9094), .ZN(n9352) );
  OR2_X1 U11856 ( .A1(n9353), .A2(n9352), .ZN(n13246) );
  INV_X1 U11857 ( .A(n13246), .ZN(n14925) );
  INV_X1 U11858 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9354) );
  MUX2_X1 U11859 ( .A(n9354), .B(P2_REG1_REG_2__SCAN_IN), .S(n13159), .Z(
        n13164) );
  INV_X1 U11860 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15067) );
  MUX2_X1 U11861 ( .A(n15067), .B(P2_REG1_REG_1__SCAN_IN), .S(n13151), .Z(
        n13149) );
  AND2_X1 U11862 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13150) );
  NAND2_X1 U11863 ( .A1(n13149), .A2(n13150), .ZN(n13148) );
  OAI21_X1 U11864 ( .B1(n15067), .B2(n13151), .A(n13148), .ZN(n13163) );
  NAND2_X1 U11865 ( .A1(n13164), .A2(n13163), .ZN(n13177) );
  OR2_X1 U11866 ( .A1(n13159), .A2(n9354), .ZN(n13176) );
  NAND2_X1 U11867 ( .A1(n13177), .A2(n13176), .ZN(n9357) );
  INV_X1 U11868 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9355) );
  MUX2_X1 U11869 ( .A(n9355), .B(P2_REG1_REG_3__SCAN_IN), .S(n13174), .Z(n9356) );
  NAND2_X1 U11870 ( .A1(n9357), .A2(n9356), .ZN(n14805) );
  NAND2_X1 U11871 ( .A1(n13169), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n14804) );
  NAND2_X1 U11872 ( .A1(n14805), .A2(n14804), .ZN(n9360) );
  MUX2_X1 U11873 ( .A(n9358), .B(P2_REG1_REG_4__SCAN_IN), .S(n14809), .Z(n9359) );
  NAND2_X1 U11874 ( .A1(n9360), .A2(n9359), .ZN(n14822) );
  OR2_X1 U11875 ( .A1(n14809), .A2(n9358), .ZN(n14821) );
  NAND2_X1 U11876 ( .A1(n14822), .A2(n14821), .ZN(n9363) );
  MUX2_X1 U11877 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9361), .S(n14819), .Z(n9362) );
  NAND2_X1 U11878 ( .A1(n9363), .A2(n9362), .ZN(n14824) );
  NAND2_X1 U11879 ( .A1(n14819), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U11880 ( .A1(n14824), .A2(n13185), .ZN(n9366) );
  MUX2_X1 U11881 ( .A(n9364), .B(P2_REG1_REG_6__SCAN_IN), .S(n13188), .Z(n9365) );
  NAND2_X1 U11882 ( .A1(n9366), .A2(n9365), .ZN(n13187) );
  NAND2_X1 U11883 ( .A1(n13183), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11884 ( .A1(n13187), .A2(n9371), .ZN(n9369) );
  MUX2_X1 U11885 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9367), .S(n9545), .Z(n9368)
         );
  NAND2_X1 U11886 ( .A1(n9369), .A2(n9368), .ZN(n13206) );
  MUX2_X1 U11887 ( .A(n9367), .B(P2_REG1_REG_7__SCAN_IN), .S(n9545), .Z(n9370)
         );
  NAND3_X1 U11888 ( .A1(n13187), .A2(n9371), .A3(n9370), .ZN(n9372) );
  NAND3_X1 U11889 ( .A1(n14925), .A2(n13206), .A3(n9372), .ZN(n9373) );
  OAI211_X1 U11890 ( .C1(n14930), .C2(n9375), .A(n9374), .B(n9373), .ZN(
        P2_U3221) );
  NAND2_X1 U11891 ( .A1(n12521), .A2(P3_DATAO_REG_20__SCAN_IN), .ZN(n9376) );
  OAI21_X1 U11892 ( .B1(n12816), .B2(n12521), .A(n9376), .ZN(P3_U3511) );
  INV_X1 U11893 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U11894 ( .A1(n9378), .A2(n9639), .ZN(n9379) );
  NAND2_X1 U11895 ( .A1(n9379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9467) );
  XNOR2_X1 U11896 ( .A(n9467), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10961) );
  INV_X1 U11897 ( .A(n10961), .ZN(n9701) );
  INV_X1 U11898 ( .A(n10960), .ZN(n9382) );
  OAI222_X1 U11899 ( .A1(P1_U3086), .A2(n9701), .B1(n11530), .B2(n9382), .C1(
        n9380), .C2(n6421), .ZN(P1_U3343) );
  INV_X1 U11900 ( .A(n14861), .ZN(n9381) );
  OAI222_X1 U11901 ( .A1(n11238), .A2(n9383), .B1(n13688), .B2(n9382), .C1(
        n9381), .C2(P2_U3088), .ZN(P2_U3315) );
  NOR2_X1 U11902 ( .A1(n9389), .A2(n9318), .ZN(n9403) );
  INV_X1 U11903 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n14178) );
  MUX2_X1 U11904 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n14178), .S(n10561), .Z(
        n9402) );
  OAI21_X1 U11905 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n9401) );
  NAND2_X1 U11906 ( .A1(n10561), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9386) );
  INV_X1 U11907 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9384) );
  MUX2_X1 U11908 ( .A(n9384), .B(P1_REG2_REG_11__SCAN_IN), .S(n10574), .Z(
        n9385) );
  AOI21_X1 U11909 ( .B1(n9401), .B2(n9386), .A(n9385), .ZN(n9506) );
  NAND3_X1 U11910 ( .A1(n9401), .A2(n9386), .A3(n9385), .ZN(n9387) );
  NAND2_X1 U11911 ( .A1(n9387), .A2(n13914), .ZN(n9398) );
  INV_X1 U11912 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U11913 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11442)
         );
  OAI21_X1 U11914 ( .B1(n14674), .B2(n14355), .A(n11442), .ZN(n9388) );
  AOI21_X1 U11915 ( .B1(n14666), .B2(n10574), .A(n9388), .ZN(n9397) );
  INV_X1 U11916 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14618) );
  MUX2_X1 U11917 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14618), .S(n10574), .Z(
        n9394) );
  NAND2_X1 U11918 ( .A1(n9389), .A2(n15311), .ZN(n9390) );
  NAND2_X1 U11919 ( .A1(n9391), .A2(n9390), .ZN(n9410) );
  INV_X1 U11920 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14770) );
  MUX2_X1 U11921 ( .A(n14770), .B(P1_REG1_REG_10__SCAN_IN), .S(n10561), .Z(
        n9409) );
  OR2_X1 U11922 ( .A1(n9410), .A2(n9409), .ZN(n9407) );
  NAND2_X1 U11923 ( .A1(n10561), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9392) );
  AND2_X1 U11924 ( .A1(n9407), .A2(n9392), .ZN(n9393) );
  NAND2_X1 U11925 ( .A1(n9393), .A2(n9394), .ZN(n9514) );
  OAI21_X1 U11926 ( .B1(n9394), .B2(n9393), .A(n9514), .ZN(n9395) );
  INV_X1 U11927 ( .A(n14669), .ZN(n13908) );
  NAND2_X1 U11928 ( .A1(n9395), .A2(n13908), .ZN(n9396) );
  OAI211_X1 U11929 ( .C1(n9506), .C2(n9398), .A(n9397), .B(n9396), .ZN(
        P1_U3254) );
  INV_X1 U11930 ( .A(n12597), .ZN(n12579) );
  OAI222_X1 U11931 ( .A1(P3_U3151), .A2(n12579), .B1(n12997), .B2(n9400), .C1(
        n14451), .C2(n9399), .ZN(P3_U3280) );
  INV_X1 U11932 ( .A(n9401), .ZN(n9406) );
  NOR3_X1 U11933 ( .A1(n9404), .A2(n9403), .A3(n9402), .ZN(n9405) );
  NOR3_X1 U11934 ( .A1(n9406), .A2(n9405), .A3(n14663), .ZN(n9415) );
  INV_X1 U11935 ( .A(n9407), .ZN(n9408) );
  AOI211_X1 U11936 ( .C1(n9410), .C2(n9409), .A(n14669), .B(n9408), .ZN(n9414)
         );
  INV_X1 U11937 ( .A(n10561), .ZN(n9412) );
  AND2_X1 U11938 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11264) );
  AOI21_X1 U11939 ( .B1(n14655), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11264), 
        .ZN(n9411) );
  OAI21_X1 U11940 ( .B1(n13849), .B2(n9412), .A(n9411), .ZN(n9413) );
  OR3_X1 U11941 ( .A1(n9415), .A2(n9414), .A3(n9413), .ZN(P1_U3253) );
  INV_X1 U11942 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9417) );
  OAI22_X1 U11943 ( .A1(n9417), .A2(n14853), .B1(n13246), .B2(n9416), .ZN(
        n9420) );
  NAND2_X1 U11944 ( .A1(n14917), .A2(n9417), .ZN(n9418) );
  OAI211_X1 U11945 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n13246), .A(n9418), .B(
        n14930), .ZN(n9419) );
  MUX2_X1 U11946 ( .A(n9420), .B(n9419), .S(P2_IR_REG_0__SCAN_IN), .Z(n9421)
         );
  INV_X1 U11947 ( .A(n9421), .ZN(n9423) );
  AOI22_X1 U11948 ( .A1(n14923), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9422) );
  NAND2_X1 U11949 ( .A1(n9423), .A2(n9422), .ZN(P2_U3214) );
  NOR2_X1 U11950 ( .A1(n12986), .A2(n9424), .ZN(n9427) );
  INV_X1 U11951 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9425) );
  NOR2_X1 U11952 ( .A1(n9451), .A2(n9425), .ZN(P3_U3260) );
  INV_X1 U11953 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9426) );
  NOR2_X1 U11954 ( .A1(n9427), .A2(n9426), .ZN(P3_U3258) );
  CLKBUF_X1 U11955 ( .A(n9427), .Z(n9451) );
  INV_X1 U11956 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9428) );
  NOR2_X1 U11957 ( .A1(n9451), .A2(n9428), .ZN(P3_U3261) );
  INV_X1 U11958 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9429) );
  NOR2_X1 U11959 ( .A1(n9427), .A2(n9429), .ZN(P3_U3262) );
  INV_X1 U11960 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9430) );
  NOR2_X1 U11961 ( .A1(n9451), .A2(n9430), .ZN(P3_U3256) );
  INV_X1 U11962 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9431) );
  NOR2_X1 U11963 ( .A1(n9451), .A2(n9431), .ZN(P3_U3255) );
  INV_X1 U11964 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9432) );
  NOR2_X1 U11965 ( .A1(n9451), .A2(n9432), .ZN(P3_U3254) );
  INV_X1 U11966 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9433) );
  NOR2_X1 U11967 ( .A1(n9451), .A2(n9433), .ZN(P3_U3253) );
  INV_X1 U11968 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9434) );
  NOR2_X1 U11969 ( .A1(n9451), .A2(n9434), .ZN(P3_U3263) );
  INV_X1 U11970 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9435) );
  NOR2_X1 U11971 ( .A1(n9451), .A2(n9435), .ZN(P3_U3257) );
  INV_X1 U11972 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9436) );
  NOR2_X1 U11973 ( .A1(n9451), .A2(n9436), .ZN(P3_U3252) );
  INV_X1 U11974 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9437) );
  NOR2_X1 U11975 ( .A1(n9451), .A2(n9437), .ZN(P3_U3251) );
  INV_X1 U11976 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9438) );
  NOR2_X1 U11977 ( .A1(n9451), .A2(n9438), .ZN(P3_U3250) );
  INV_X1 U11978 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U11979 ( .A1(n9451), .A2(n9439), .ZN(P3_U3249) );
  INV_X1 U11980 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9440) );
  NOR2_X1 U11981 ( .A1(n9451), .A2(n9440), .ZN(P3_U3248) );
  INV_X1 U11982 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9441) );
  NOR2_X1 U11983 ( .A1(n9451), .A2(n9441), .ZN(P3_U3247) );
  INV_X1 U11984 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9442) );
  NOR2_X1 U11985 ( .A1(n9451), .A2(n9442), .ZN(P3_U3246) );
  INV_X1 U11986 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n15201) );
  NOR2_X1 U11987 ( .A1(n9427), .A2(n15201), .ZN(P3_U3245) );
  INV_X1 U11988 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15289) );
  NOR2_X1 U11989 ( .A1(n9427), .A2(n15289), .ZN(P3_U3244) );
  INV_X1 U11990 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9443) );
  NOR2_X1 U11991 ( .A1(n9427), .A2(n9443), .ZN(P3_U3243) );
  INV_X1 U11992 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9444) );
  NOR2_X1 U11993 ( .A1(n9427), .A2(n9444), .ZN(P3_U3242) );
  INV_X1 U11994 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15258) );
  NOR2_X1 U11995 ( .A1(n9427), .A2(n15258), .ZN(P3_U3241) );
  INV_X1 U11996 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9445) );
  NOR2_X1 U11997 ( .A1(n9427), .A2(n9445), .ZN(P3_U3240) );
  INV_X1 U11998 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9446) );
  NOR2_X1 U11999 ( .A1(n9427), .A2(n9446), .ZN(P3_U3239) );
  INV_X1 U12000 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9447) );
  NOR2_X1 U12001 ( .A1(n9427), .A2(n9447), .ZN(P3_U3238) );
  INV_X1 U12002 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9448) );
  NOR2_X1 U12003 ( .A1(n9427), .A2(n9448), .ZN(P3_U3237) );
  INV_X1 U12004 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9449) );
  NOR2_X1 U12005 ( .A1(n9451), .A2(n9449), .ZN(P3_U3236) );
  INV_X1 U12006 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9450) );
  NOR2_X1 U12007 ( .A1(n9451), .A2(n9450), .ZN(P3_U3259) );
  INV_X1 U12008 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U12009 ( .A1(n9451), .A2(n9452), .ZN(P3_U3235) );
  INV_X1 U12010 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9453) );
  NOR2_X1 U12011 ( .A1(n9451), .A2(n9453), .ZN(P3_U3234) );
  INV_X1 U12012 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14342) );
  NAND2_X1 U12013 ( .A1(n14666), .A2(n10074), .ZN(n9454) );
  NAND2_X1 U12014 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10518) );
  OAI211_X1 U12015 ( .C1(n14342), .C2(n14674), .A(n9454), .B(n10518), .ZN(
        n9464) );
  INV_X1 U12016 ( .A(n9491), .ZN(n9455) );
  AOI211_X1 U12017 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n14669), .ZN(n9463)
         );
  AND3_X1 U12018 ( .A1(n13903), .A2(n9459), .A3(n9458), .ZN(n9460) );
  NOR3_X1 U12019 ( .A1(n14663), .A2(n9461), .A3(n9460), .ZN(n9462) );
  OR3_X1 U12020 ( .A1(n9464), .A2(n9463), .A3(n9462), .ZN(P1_U3249) );
  INV_X1 U12021 ( .A(n11058), .ZN(n9472) );
  INV_X1 U12022 ( .A(n9976), .ZN(n13228) );
  OAI222_X1 U12023 ( .A1(n11238), .A2(n9465), .B1(n13688), .B2(n9472), .C1(
        n13228), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12024 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U12025 ( .A1(n9467), .A2(n9466), .ZN(n9468) );
  NAND2_X1 U12026 ( .A1(n9468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9470) );
  INV_X1 U12027 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U12028 ( .A1(n9470), .A2(n9469), .ZN(n9677) );
  OR2_X1 U12029 ( .A1(n9470), .A2(n9469), .ZN(n9471) );
  INV_X1 U12030 ( .A(n11061), .ZN(n9749) );
  OAI222_X1 U12031 ( .A1(P1_U3086), .A2(n9749), .B1(n11530), .B2(n9472), .C1(
        n11059), .C2(n6421), .ZN(P1_U3342) );
  INV_X1 U12032 ( .A(n9473), .ZN(n13840) );
  MUX2_X1 U12033 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9309), .S(n9587), .Z(n9476)
         );
  INV_X1 U12034 ( .A(n9474), .ZN(n9475) );
  AOI211_X1 U12035 ( .C1(n13840), .C2(n9476), .A(n9475), .B(n14663), .ZN(n9482) );
  MUX2_X1 U12036 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9289), .S(n9587), .Z(n9477)
         );
  OAI21_X1 U12037 ( .B1(n9478), .B2(n13842), .A(n9477), .ZN(n9479) );
  AND3_X1 U12038 ( .A1(n13908), .A2(n9480), .A3(n9479), .ZN(n9481) );
  NOR2_X1 U12039 ( .A1(n9482), .A2(n9481), .ZN(n9484) );
  AOI22_X1 U12040 ( .A1(n14655), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9483) );
  OAI211_X1 U12041 ( .C1(n9587), .C2(n13849), .A(n9484), .B(n9483), .ZN(
        P1_U3244) );
  INV_X1 U12042 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15203) );
  NAND2_X1 U12043 ( .A1(P3_U3897), .A2(n11202), .ZN(n9485) );
  OAI21_X1 U12044 ( .B1(P3_U3897), .B2(n15203), .A(n9485), .ZN(P3_U3502) );
  INV_X1 U12045 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U12046 ( .A1(P3_U3897), .A2(n12840), .ZN(n9486) );
  OAI21_X1 U12047 ( .B1(P3_U3897), .B2(n15333), .A(n9486), .ZN(P3_U3509) );
  INV_X1 U12048 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15332) );
  NAND2_X1 U12049 ( .A1(P3_U3897), .A2(n10856), .ZN(n9487) );
  OAI21_X1 U12050 ( .B1(P3_U3897), .B2(n15332), .A(n9487), .ZN(P3_U3494) );
  INV_X1 U12051 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U12052 ( .A1(P3_U3897), .A2(n15144), .ZN(n9488) );
  OAI21_X1 U12053 ( .B1(P3_U3897), .B2(n15327), .A(n9488), .ZN(P3_U3493) );
  MUX2_X1 U12054 ( .A(n9298), .B(P1_REG1_REG_7__SCAN_IN), .S(n10079), .Z(n9489) );
  NAND3_X1 U12055 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n9492) );
  NAND3_X1 U12056 ( .A1(n13908), .A2(n9493), .A3(n9492), .ZN(n9500) );
  NAND2_X1 U12057 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10793) );
  AOI211_X1 U12058 ( .C1(n9495), .C2(n9494), .A(n9529), .B(n14663), .ZN(n9496)
         );
  INV_X1 U12059 ( .A(n9496), .ZN(n9497) );
  NAND2_X1 U12060 ( .A1(n10793), .A2(n9497), .ZN(n9498) );
  AOI21_X1 U12061 ( .B1(n14655), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9498), .ZN(
        n9499) );
  OAI211_X1 U12062 ( .C1(n13849), .C2(n9501), .A(n9500), .B(n9499), .ZN(
        P1_U3250) );
  INV_X1 U12063 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U12064 ( .A1(P3_U3897), .A2(n6689), .ZN(n9502) );
  OAI21_X1 U12065 ( .B1(P3_U3897), .B2(n15234), .A(n9502), .ZN(P3_U3492) );
  INV_X1 U12066 ( .A(n12602), .ZN(n12600) );
  OAI222_X1 U12067 ( .A1(P3_U3151), .A2(n12600), .B1(n12997), .B2(n9504), .C1(
        n14451), .C2(n9503), .ZN(P3_U3279) );
  INV_X1 U12068 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9505) );
  MUX2_X1 U12069 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9505), .S(n10961), .Z(
        n9508) );
  AOI21_X1 U12070 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10574), .A(n9506), .ZN(
        n9507) );
  NAND2_X1 U12071 ( .A1(n9507), .A2(n9508), .ZN(n9691) );
  OAI21_X1 U12072 ( .B1(n9508), .B2(n9507), .A(n9691), .ZN(n9520) );
  NAND2_X1 U12073 ( .A1(n9509), .A2(n14618), .ZN(n9512) );
  NAND2_X1 U12074 ( .A1(n9514), .A2(n9512), .ZN(n9510) );
  INV_X1 U12075 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U12076 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9700), .S(n10961), .Z(
        n9511) );
  NAND2_X1 U12077 ( .A1(n9510), .A2(n9511), .ZN(n9703) );
  INV_X1 U12078 ( .A(n9511), .ZN(n9513) );
  NAND3_X1 U12079 ( .A1(n9514), .A2(n9513), .A3(n9512), .ZN(n9515) );
  AOI21_X1 U12080 ( .B1(n9703), .B2(n9515), .A(n14669), .ZN(n9519) );
  INV_X1 U12081 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11486) );
  NOR2_X1 U12082 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11486), .ZN(n9516) );
  AOI21_X1 U12083 ( .B1(n14655), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9516), .ZN(
        n9517) );
  OAI21_X1 U12084 ( .B1(n13849), .B2(n9701), .A(n9517), .ZN(n9518) );
  AOI211_X1 U12085 ( .C1(n9520), .C2(n13914), .A(n9519), .B(n9518), .ZN(n9521)
         );
  INV_X1 U12086 ( .A(n9521), .ZN(P1_U3255) );
  OAI21_X1 U12087 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9534) );
  INV_X1 U12088 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14348) );
  NAND2_X1 U12089 ( .A1(n14666), .A2(n10274), .ZN(n9525) );
  NAND2_X1 U12090 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11012) );
  OAI211_X1 U12091 ( .C1(n14348), .C2(n14674), .A(n9525), .B(n11012), .ZN(
        n9533) );
  INV_X1 U12092 ( .A(n9526), .ZN(n9531) );
  NOR3_X1 U12093 ( .A1(n9529), .A2(n9528), .A3(n9527), .ZN(n9530) );
  NOR3_X1 U12094 ( .A1(n9531), .A2(n9530), .A3(n14663), .ZN(n9532) );
  AOI211_X1 U12095 ( .C1(n13908), .C2(n9534), .A(n9533), .B(n9532), .ZN(n9535)
         );
  INV_X1 U12096 ( .A(n9535), .ZN(P1_U3251) );
  NAND2_X1 U12097 ( .A1(n9545), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U12098 ( .A1(n13200), .A2(n13199), .ZN(n9537) );
  MUX2_X1 U12099 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10748), .S(n13203), .Z(
        n9536) );
  NAND2_X1 U12100 ( .A1(n9537), .A2(n9536), .ZN(n13202) );
  NAND2_X1 U12101 ( .A1(n13203), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12102 ( .A1(n13202), .A2(n9538), .ZN(n14836) );
  MUX2_X1 U12103 ( .A(n10938), .B(P2_REG2_REG_9__SCAN_IN), .S(n9550), .Z(
        n14835) );
  OAI21_X1 U12104 ( .B1(n9550), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14838), .ZN(
        n14854) );
  MUX2_X1 U12105 ( .A(n11044), .B(P2_REG2_REG_10__SCAN_IN), .S(n14848), .Z(
        n14855) );
  NOR2_X1 U12106 ( .A1(n14854), .A2(n14855), .ZN(n14852) );
  MUX2_X1 U12107 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11191), .S(n9975), .Z(
        n9539) );
  NAND2_X1 U12108 ( .A1(n9540), .A2(n9539), .ZN(n9974) );
  OAI21_X1 U12109 ( .B1(n9540), .B2(n9539), .A(n9974), .ZN(n9557) );
  NAND2_X1 U12110 ( .A1(n14923), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n9543) );
  NOR2_X1 U12111 ( .A1(n9541), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11108) );
  INV_X1 U12112 ( .A(n11108), .ZN(n9542) );
  OAI211_X1 U12113 ( .C1(n14930), .C2(n9544), .A(n9543), .B(n9542), .ZN(n9556)
         );
  INV_X1 U12114 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15075) );
  NAND2_X1 U12115 ( .A1(n9545), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U12116 ( .A1(n13206), .A2(n13205), .ZN(n9548) );
  MUX2_X1 U12117 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9546), .S(n13203), .Z(n9547) );
  NAND2_X1 U12118 ( .A1(n9548), .A2(n9547), .ZN(n13208) );
  NAND2_X1 U12119 ( .A1(n13203), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9549) );
  AND2_X1 U12120 ( .A1(n13208), .A2(n9549), .ZN(n14832) );
  MUX2_X1 U12121 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15075), .S(n9550), .Z(
        n14831) );
  AOI21_X1 U12122 ( .B1(n15075), .B2(n14842), .A(n14834), .ZN(n14851) );
  MUX2_X1 U12123 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9551), .S(n14848), .Z(
        n14850) );
  NAND2_X1 U12124 ( .A1(n14851), .A2(n14850), .ZN(n14849) );
  NAND2_X1 U12125 ( .A1(n14848), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9553) );
  INV_X1 U12126 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15079) );
  MUX2_X1 U12127 ( .A(n15079), .B(P2_REG1_REG_11__SCAN_IN), .S(n9975), .Z(
        n9552) );
  AOI21_X1 U12128 ( .B1(n14849), .B2(n9553), .A(n9552), .ZN(n9970) );
  AND3_X1 U12129 ( .A1(n14849), .A2(n9553), .A3(n9552), .ZN(n9554) );
  NOR3_X1 U12130 ( .A1(n9970), .A2(n9554), .A3(n13246), .ZN(n9555) );
  AOI211_X1 U12131 ( .C1(n14917), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9558)
         );
  INV_X1 U12132 ( .A(n9558), .ZN(P2_U3225) );
  NAND3_X1 U12133 ( .A1(n13966), .A2(n9684), .A3(n9559), .ZN(n9575) );
  NOR2_X1 U12134 ( .A1(n9575), .A2(n9576), .ZN(n13805) );
  NAND2_X1 U12135 ( .A1(n13805), .A2(n14575), .ZN(n14551) );
  NAND2_X1 U12136 ( .A1(n10254), .A2(n13838), .ZN(n9566) );
  INV_X1 U12137 ( .A(n9560), .ZN(n9564) );
  NAND2_X1 U12138 ( .A1(n9564), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U12139 ( .A1(n9567), .A2(n9628), .ZN(n9627) );
  OAI21_X1 U12140 ( .B1(n9567), .B2(n9628), .A(n9627), .ZN(n13839) );
  NOR2_X1 U12141 ( .A1(n9575), .A2(n9568), .ZN(n9579) );
  NOR2_X1 U12142 ( .A1(n9569), .A2(n11860), .ZN(n14470) );
  INV_X1 U12143 ( .A(n14470), .ZN(n14580) );
  INV_X1 U12144 ( .A(n9569), .ZN(n9570) );
  NAND2_X1 U12145 ( .A1(n9570), .A2(n14184), .ZN(n9571) );
  NAND2_X1 U12146 ( .A1(n14580), .A2(n9571), .ZN(n14755) );
  NOR2_X1 U12147 ( .A1(n14755), .A2(n9572), .ZN(n9573) );
  NAND2_X1 U12148 ( .A1(n9579), .A2(n9573), .ZN(n14559) );
  NAND2_X1 U12149 ( .A1(n9575), .A2(n9574), .ZN(n10179) );
  INV_X1 U12150 ( .A(n10179), .ZN(n9577) );
  NOR2_X1 U12151 ( .A1(n9577), .A2(n9576), .ZN(n9731) );
  INV_X1 U12152 ( .A(n9731), .ZN(n9578) );
  AOI22_X1 U12153 ( .A1(n13839), .A2(n13810), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n9578), .ZN(n9583) );
  NAND2_X1 U12154 ( .A1(n9579), .A2(n14470), .ZN(n9581) );
  NAND2_X2 U12155 ( .A1(n9580), .A2(n9687), .ZN(n14698) );
  NAND2_X1 U12156 ( .A1(n9581), .A2(n14698), .ZN(n14564) );
  NAND2_X1 U12157 ( .A1(n14564), .A2(n9584), .ZN(n9582) );
  OAI211_X1 U12158 ( .C1(n9732), .C2(n14551), .A(n9583), .B(n9582), .ZN(
        P1_U3232) );
  INV_X1 U12159 ( .A(n11535), .ZN(n9596) );
  INV_X1 U12160 ( .A(n9585), .ZN(n9586) );
  NAND2_X1 U12161 ( .A1(n9925), .A2(n9586), .ZN(n9595) );
  NAND2_X1 U12162 ( .A1(n6412), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9592) );
  INV_X1 U12163 ( .A(n9587), .ZN(n9588) );
  NAND3_X1 U12164 ( .A1(n6424), .A2(n9588), .A3(n6415), .ZN(n9591) );
  INV_X1 U12165 ( .A(n9592), .ZN(n9589) );
  NAND2_X1 U12166 ( .A1(n11914), .A2(n9589), .ZN(n9590) );
  OAI211_X1 U12167 ( .C1(n6424), .C2(n9592), .A(n9591), .B(n9590), .ZN(n9593)
         );
  INV_X1 U12168 ( .A(n9593), .ZN(n9594) );
  AND2_X2 U12169 ( .A1(n9595), .A2(n9594), .ZN(n14717) );
  NAND2_X1 U12170 ( .A1(n13837), .A2(n14717), .ZN(n11546) );
  OR2_X2 U12171 ( .A1(n13837), .A2(n14717), .ZN(n11547) );
  INV_X1 U12172 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9597) );
  INV_X1 U12173 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10051) );
  INV_X1 U12174 ( .A(n9604), .ZN(n9605) );
  NAND2_X1 U12175 ( .A1(n9605), .A2(n9925), .ZN(n9608) );
  AOI22_X1 U12176 ( .A1(n11660), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n11659), 
        .B2(n9606), .ZN(n9607) );
  XNOR2_X1 U12177 ( .A(n9924), .B(n9951), .ZN(n9619) );
  AND2_X2 U12178 ( .A1(n11547), .A2(n11546), .ZN(n11878) );
  INV_X1 U12179 ( .A(n9905), .ZN(n9610) );
  INV_X1 U12180 ( .A(n14717), .ZN(n9609) );
  XNOR2_X1 U12181 ( .A(n9952), .B(n9951), .ZN(n9617) );
  OR2_X1 U12182 ( .A1(n11862), .A2(n6424), .ZN(n14165) );
  NAND2_X1 U12183 ( .A1(n11707), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9615) );
  OR2_X1 U12184 ( .A1(n11818), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9614) );
  OR2_X1 U12185 ( .A1(n11820), .A2(n14699), .ZN(n9613) );
  OAI22_X1 U12186 ( .A1(n9732), .A2(n14165), .B1(n10185), .B2(n11394), .ZN(
        n9616) );
  AOI21_X1 U12187 ( .B1(n9617), .B2(n14762), .A(n9616), .ZN(n9618) );
  OAI21_X1 U12188 ( .B1(n14570), .B2(n9619), .A(n9618), .ZN(n10053) );
  INV_X1 U12189 ( .A(n10053), .ZN(n9620) );
  AND2_X1 U12190 ( .A1(n14717), .A2(n9906), .ZN(n9908) );
  OAI211_X1 U12191 ( .C1(n11552), .C2(n9908), .A(n14707), .B(n14706), .ZN(
        n10052) );
  NAND2_X1 U12192 ( .A1(n9620), .A2(n10052), .ZN(n10058) );
  INV_X1 U12193 ( .A(n10058), .ZN(n9622) );
  NAND2_X1 U12194 ( .A1(n14772), .A2(n14755), .ZN(n14259) );
  INV_X1 U12195 ( .A(n14259), .ZN(n14263) );
  AOI22_X1 U12196 ( .A1(n14263), .A2(n11542), .B1(n6820), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n9621) );
  OAI21_X1 U12197 ( .B1(n9622), .B2(n6820), .A(n9621), .ZN(P1_U3530) );
  XNOR2_X1 U12198 ( .A(n9623), .B(n9724), .ZN(n9624) );
  OAI21_X1 U12199 ( .B1(n12039), .B2(n9628), .A(n9627), .ZN(n9629) );
  OAI21_X1 U12200 ( .B1(n9630), .B2(n9629), .A(n9728), .ZN(n9631) );
  NAND2_X1 U12201 ( .A1(n9631), .A2(n13810), .ZN(n9634) );
  INV_X2 U12202 ( .A(n14165), .ZN(n14572) );
  INV_X1 U12203 ( .A(n13805), .ZN(n13815) );
  NAND2_X1 U12204 ( .A1(n13836), .A2(n14575), .ZN(n9916) );
  OAI22_X1 U12205 ( .A1(n9731), .A2(n9910), .B1(n13815), .B2(n9916), .ZN(n9632) );
  AOI21_X1 U12206 ( .B1(n13794), .B2(n13838), .A(n9632), .ZN(n9633) );
  OAI211_X1 U12207 ( .C1(n14717), .C2(n13821), .A(n9634), .B(n9633), .ZN(
        P1_U3222) );
  INV_X1 U12208 ( .A(n12641), .ZN(n12651) );
  INV_X1 U12209 ( .A(n9635), .ZN(n9637) );
  OAI222_X1 U12210 ( .A1(n12651), .A2(P3_U3151), .B1(n14451), .B2(n9637), .C1(
        n9636), .C2(n12997), .ZN(P3_U3278) );
  INV_X1 U12211 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9638) );
  NAND3_X1 U12212 ( .A1(n15288), .A2(n9639), .A3(n9638), .ZN(n9640) );
  OR2_X1 U12213 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  NOR2_X1 U12214 ( .A1(n9643), .A2(n9642), .ZN(n9714) );
  INV_X1 U12215 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U12216 ( .A1(n9714), .A2(n9715), .ZN(n9717) );
  NAND2_X1 U12217 ( .A1(n9717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9644) );
  MUX2_X1 U12218 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9644), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9645) );
  OR2_X1 U12219 ( .A1(n9717), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n10061) );
  AND2_X1 U12220 ( .A1(n9645), .A2(n10061), .ZN(n13912) );
  INV_X1 U12221 ( .A(n13912), .ZN(n10667) );
  INV_X1 U12222 ( .A(n11375), .ZN(n9647) );
  OAI222_X1 U12223 ( .A1(P1_U3086), .A2(n10667), .B1(n11530), .B2(n9647), .C1(
        n9646), .C2(n6421), .ZN(P1_U3339) );
  INV_X1 U12224 ( .A(n13235), .ZN(n14904) );
  OAI222_X1 U12225 ( .A1(n11238), .A2(n9648), .B1(n13688), .B2(n9647), .C1(
        n14904), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U12226 ( .A(n15059), .ZN(n15013) );
  NAND2_X1 U12227 ( .A1(n10946), .A2(n10674), .ZN(n9753) );
  INV_X1 U12228 ( .A(n9753), .ZN(n9760) );
  AND2_X1 U12229 ( .A1(n13530), .A2(n9760), .ZN(n14934) );
  INV_X1 U12230 ( .A(n10144), .ZN(n9757) );
  AND2_X1 U12231 ( .A1(n6413), .A2(n13254), .ZN(n9772) );
  INV_X1 U12232 ( .A(n9772), .ZN(n9656) );
  NAND2_X1 U12233 ( .A1(n8354), .A2(n9649), .ZN(n9650) );
  NAND2_X1 U12234 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  OR2_X1 U12235 ( .A1(n8951), .A2(n10674), .ZN(n9654) );
  OR2_X1 U12236 ( .A1(n10369), .A2(n10946), .ZN(n9653) );
  OAI21_X1 U12237 ( .B1(n15064), .B2(n15026), .A(n14932), .ZN(n9655) );
  NAND2_X1 U12238 ( .A1(n9656), .A2(n9655), .ZN(n14939) );
  AOI211_X1 U12239 ( .C1(n15013), .C2(n14932), .A(n14934), .B(n14939), .ZN(
        n14980) );
  INV_X1 U12240 ( .A(P2_B_REG_SCAN_IN), .ZN(n13255) );
  XOR2_X1 U12241 ( .A(n11236), .B(n13255), .Z(n9657) );
  INV_X1 U12242 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14975) );
  NAND2_X1 U12243 ( .A1(n14944), .A2(n14975), .ZN(n9659) );
  NAND2_X1 U12244 ( .A1(n13689), .A2(n11236), .ZN(n9658) );
  NAND2_X1 U12245 ( .A1(n10365), .A2(n14979), .ZN(n14974) );
  INV_X1 U12246 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14977) );
  NAND2_X1 U12247 ( .A1(n14944), .A2(n14977), .ZN(n9663) );
  NAND2_X1 U12248 ( .A1(n13689), .A2(n11361), .ZN(n9662) );
  NAND2_X1 U12249 ( .A1(n9663), .A2(n9662), .ZN(n14978) );
  NOR4_X1 U12250 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n9667) );
  NOR4_X1 U12251 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n9666) );
  NOR4_X1 U12252 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n9665) );
  NOR4_X1 U12253 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9664) );
  NAND4_X1 U12254 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n9673)
         );
  NOR2_X1 U12255 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n9671) );
  NOR4_X1 U12256 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9670) );
  NOR4_X1 U12257 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9669) );
  NOR4_X1 U12258 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9668) );
  NAND4_X1 U12259 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n9672)
         );
  OAI21_X1 U12260 ( .B1(n9673), .B2(n9672), .A(n14944), .ZN(n10199) );
  OR2_X1 U12261 ( .A1(n15059), .A2(n9674), .ZN(n9761) );
  NAND2_X1 U12262 ( .A1(n9769), .A2(n9757), .ZN(n10363) );
  AND2_X1 U12263 ( .A1(n9761), .A2(n10363), .ZN(n10198) );
  NAND3_X1 U12264 ( .A1(n14978), .A2(n10199), .A3(n10198), .ZN(n9675) );
  NAND2_X1 U12265 ( .A1(n15078), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9676) );
  OAI21_X1 U12266 ( .B1(n14980), .B2(n15078), .A(n9676), .ZN(P2_U3499) );
  NAND2_X1 U12267 ( .A1(n9677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U12268 ( .A(n9678), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11147) );
  INV_X1 U12269 ( .A(n11147), .ZN(n10658) );
  INV_X1 U12270 ( .A(n11146), .ZN(n9680) );
  OAI222_X1 U12271 ( .A1(P1_U3086), .A2(n10658), .B1(n11530), .B2(n9680), .C1(
        n9679), .C2(n6421), .ZN(P1_U3341) );
  INV_X1 U12272 ( .A(n14876), .ZN(n13219) );
  OAI222_X1 U12273 ( .A1(n11238), .A2(n9681), .B1(n13688), .B2(n9680), .C1(
        n13219), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12274 ( .A(n12668), .ZN(n12644) );
  INV_X1 U12275 ( .A(SI_18_), .ZN(n9683) );
  OAI222_X1 U12276 ( .A1(P3_U3151), .A2(n12644), .B1(n12997), .B2(n9683), .C1(
        n14451), .C2(n9682), .ZN(P3_U3277) );
  INV_X1 U12277 ( .A(n9684), .ZN(n9685) );
  NOR2_X1 U12278 ( .A1(n13966), .A2(n9687), .ZN(n9688) );
  INV_X2 U12279 ( .A(n14763), .ZN(n14764) );
  NAND2_X1 U12280 ( .A1(n14764), .A2(n9689), .ZN(n9690) );
  OAI21_X1 U12281 ( .B1(n14764), .B2(n9285), .A(n9690), .ZN(P1_U3459) );
  OAI21_X1 U12282 ( .B1(n10961), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9691), .ZN(
        n9742) );
  INV_X1 U12283 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9692) );
  MUX2_X1 U12284 ( .A(n9692), .B(P1_REG2_REG_13__SCAN_IN), .S(n11061), .Z(
        n9743) );
  NOR2_X1 U12285 ( .A1(n9742), .A2(n9743), .ZN(n9741) );
  INV_X1 U12286 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U12287 ( .A(n9693), .B(P1_REG2_REG_14__SCAN_IN), .S(n11147), .Z(
        n9695) );
  NAND2_X1 U12288 ( .A1(n11061), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U12289 ( .A1(n9695), .A2(n9696), .ZN(n9694) );
  OAI21_X1 U12290 ( .B1(n9741), .B2(n9694), .A(n13914), .ZN(n9712) );
  INV_X1 U12291 ( .A(n9741), .ZN(n9697) );
  AOI21_X1 U12292 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n10656) );
  INV_X1 U12293 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12294 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14548)
         );
  OAI21_X1 U12295 ( .B1(n14674), .B2(n9698), .A(n14548), .ZN(n9699) );
  AOI21_X1 U12296 ( .B1(n11147), .B2(n14666), .A(n9699), .ZN(n9711) );
  INV_X1 U12297 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14612) );
  MUX2_X1 U12298 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14612), .S(n11147), .Z(
        n9708) );
  NAND2_X1 U12299 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  NAND2_X1 U12300 ( .A1(n9703), .A2(n9702), .ZN(n9737) );
  INV_X1 U12301 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9704) );
  MUX2_X1 U12302 ( .A(n9704), .B(P1_REG1_REG_13__SCAN_IN), .S(n11061), .Z(
        n9705) );
  NAND2_X1 U12303 ( .A1(n11061), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12304 ( .A1(n9707), .A2(n9708), .ZN(n10665) );
  OAI21_X1 U12305 ( .B1(n9708), .B2(n9707), .A(n10665), .ZN(n9709) );
  NAND2_X1 U12306 ( .A1(n9709), .A2(n13908), .ZN(n9710) );
  OAI211_X1 U12307 ( .C1(n9712), .C2(n10656), .A(n9711), .B(n9710), .ZN(
        P1_U3257) );
  INV_X1 U12308 ( .A(n11337), .ZN(n9719) );
  INV_X1 U12309 ( .A(n14884), .ZN(n13231) );
  OAI222_X1 U12310 ( .A1(n11238), .A2(n9713), .B1(n13688), .B2(n9719), .C1(
        P2_U3088), .C2(n13231), .ZN(P2_U3312) );
  OR2_X1 U12311 ( .A1(n9714), .A2(n9159), .ZN(n9716) );
  MUX2_X1 U12312 ( .A(n9716), .B(P1_IR_REG_31__SCAN_IN), .S(n9715), .Z(n9718)
         );
  NAND2_X1 U12313 ( .A1(n9718), .A2(n9717), .ZN(n11339) );
  OAI222_X1 U12314 ( .A1(n11339), .A2(P1_U3086), .B1(n11530), .B2(n9719), .C1(
        n11338), .C2(n6421), .ZN(P1_U3340) );
  NAND2_X1 U12315 ( .A1(n10061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9720) );
  XNOR2_X1 U12316 ( .A(n9720), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11644) );
  INV_X1 U12317 ( .A(n11644), .ZN(n11024) );
  INV_X1 U12318 ( .A(n11643), .ZN(n9723) );
  OAI222_X1 U12319 ( .A1(P1_U3086), .A2(n11024), .B1(n11530), .B2(n9723), .C1(
        n9721), .C2(n6421), .ZN(P1_U3338) );
  INV_X1 U12320 ( .A(n14905), .ZN(n13237) );
  OAI222_X1 U12321 ( .A1(P2_U3088), .A2(n13237), .B1(n13688), .B2(n9723), .C1(
        n9722), .C2(n11238), .ZN(P2_U3310) );
  OAI22_X1 U12322 ( .A1(n10184), .A2(n11556), .B1(n11552), .B2(n12047), .ZN(
        n10186) );
  XOR2_X1 U12323 ( .A(n10186), .B(n10187), .Z(n9730) );
  INV_X1 U12324 ( .A(n9726), .ZN(n9727) );
  OAI21_X1 U12325 ( .B1(n9730), .B2(n9729), .A(n10191), .ZN(n9735) );
  OAI22_X1 U12326 ( .A1(n9731), .A2(n10051), .B1(n14551), .B2(n10185), .ZN(
        n9734) );
  INV_X1 U12327 ( .A(n13794), .ZN(n14554) );
  OAI22_X1 U12328 ( .A1(n11552), .A2(n13821), .B1(n14554), .B2(n9732), .ZN(
        n9733) );
  AOI211_X1 U12329 ( .C1(n9735), .C2(n13810), .A(n9734), .B(n9733), .ZN(n9736)
         );
  INV_X1 U12330 ( .A(n9736), .ZN(P1_U3237) );
  INV_X1 U12331 ( .A(n9737), .ZN(n9740) );
  MUX2_X1 U12332 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9704), .S(n11061), .Z(
        n9739) );
  OAI211_X1 U12333 ( .C1(n9740), .C2(n9739), .A(n13908), .B(n9738), .ZN(n9748)
         );
  NAND2_X1 U12334 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13777)
         );
  AOI211_X1 U12335 ( .C1(n9743), .C2(n9742), .A(n9741), .B(n14663), .ZN(n9744)
         );
  INV_X1 U12336 ( .A(n9744), .ZN(n9745) );
  NAND2_X1 U12337 ( .A1(n13777), .A2(n9745), .ZN(n9746) );
  AOI21_X1 U12338 ( .B1(n14655), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9746), .ZN(
        n9747) );
  OAI211_X1 U12339 ( .C1(n13849), .C2(n9749), .A(n9748), .B(n9747), .ZN(
        P1_U3256) );
  OAI222_X1 U12340 ( .A1(n14451), .A2(n9751), .B1(n12997), .B2(n9750), .C1(
        P3_U3151), .C2(n12499), .ZN(P3_U3276) );
  INV_X1 U12341 ( .A(n10199), .ZN(n9752) );
  OR2_X1 U12342 ( .A1(n10366), .A2(n14974), .ZN(n9756) );
  NOR2_X1 U12343 ( .A1(n8951), .A2(n9753), .ZN(n10370) );
  INV_X1 U12344 ( .A(n10370), .ZN(n9755) );
  INV_X1 U12345 ( .A(n9761), .ZN(n9754) );
  OAI21_X1 U12346 ( .B1(n9756), .B2(n9755), .A(n14938), .ZN(n14794) );
  INV_X1 U12347 ( .A(n14794), .ZN(n13109) );
  INV_X1 U12348 ( .A(n9756), .ZN(n9759) );
  NOR2_X1 U12349 ( .A1(n15053), .A2(n9757), .ZN(n9758) );
  OR2_X1 U12350 ( .A1(n14777), .A2(n13496), .ZN(n13110) );
  INV_X1 U12351 ( .A(n13110), .ZN(n13096) );
  INV_X1 U12352 ( .A(n10365), .ZN(n9762) );
  OAI21_X1 U12353 ( .B1(n9762), .B2(n10366), .A(n9761), .ZN(n9766) );
  INV_X1 U12354 ( .A(n10363), .ZN(n9763) );
  NOR2_X1 U12355 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  NAND2_X1 U12356 ( .A1(n9766), .A2(n9765), .ZN(n10494) );
  OR2_X1 U12357 ( .A1(n10494), .A2(P2_U3088), .ZN(n10349) );
  AOI22_X1 U12358 ( .A1(n13096), .A2(n9767), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10349), .ZN(n9775) );
  AND2_X1 U12359 ( .A1(n13530), .A2(n11136), .ZN(n9768) );
  NOR2_X1 U12360 ( .A1(n13539), .A2(n9768), .ZN(n10307) );
  INV_X1 U12361 ( .A(n10307), .ZN(n9773) );
  INV_X1 U12362 ( .A(n14974), .ZN(n9771) );
  NOR2_X1 U12363 ( .A1(n10366), .A2(n9769), .ZN(n9770) );
  AOI22_X1 U12364 ( .A1(n14788), .A2(n9773), .B1(n9772), .B2(n14534), .ZN(
        n9774) );
  OAI211_X1 U12365 ( .C1(n13109), .C2(n10305), .A(n9775), .B(n9774), .ZN(
        P2_U3204) );
  INV_X1 U12366 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U12367 ( .A1(n10004), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9785) );
  OAI21_X1 U12368 ( .B1(n10004), .B2(P3_REG1_REG_6__SCAN_IN), .A(n9785), .ZN(
        n9993) );
  XNOR2_X1 U12369 ( .A(n10005), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10008) );
  INV_X1 U12370 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9875) );
  OAI21_X1 U12371 ( .B1(n10050), .B2(n9776), .A(n7548), .ZN(n10036) );
  INV_X1 U12372 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15188) );
  INV_X1 U12373 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9777) );
  OR2_X1 U12374 ( .A1(n10005), .A2(n9777), .ZN(n9778) );
  NAND2_X1 U12375 ( .A1(n9779), .A2(n10035), .ZN(n9780) );
  INV_X1 U12376 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15190) );
  INV_X1 U12377 ( .A(n9780), .ZN(n9847) );
  XNOR2_X1 U12378 ( .A(n9860), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n9846) );
  INV_X1 U12379 ( .A(n9860), .ZN(n9830) );
  NAND2_X1 U12380 ( .A1(n9830), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9781) );
  INV_X1 U12381 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12382 ( .A1(n9782), .A2(n10163), .ZN(n9783) );
  INV_X1 U12383 ( .A(n9785), .ZN(n9786) );
  AOI21_X1 U12384 ( .B1(n10322), .B2(n9787), .A(n9877), .ZN(n9843) );
  OR2_X1 U12385 ( .A1(n9790), .A2(P3_U3151), .ZN(n12506) );
  NAND2_X1 U12386 ( .A1(n9788), .A2(n12506), .ZN(n9793) );
  AOI21_X1 U12387 ( .B1(n12487), .B2(n9790), .A(n9789), .ZN(n9792) );
  NAND2_X1 U12388 ( .A1(n9793), .A2(n9792), .ZN(n9838) );
  INV_X1 U12389 ( .A(n9838), .ZN(n9791) );
  MUX2_X1 U12390 ( .A(P3_U3897), .B(n9791), .S(n8139), .Z(n15106) );
  INV_X1 U12391 ( .A(n9792), .ZN(n9794) );
  NAND2_X1 U12392 ( .A1(n15082), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n9825) );
  AND2_X1 U12393 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10433) );
  INV_X1 U12394 ( .A(n10433), .ZN(n9824) );
  OR2_X1 U12395 ( .A1(n12521), .A2(n9795), .ZN(n15110) );
  INV_X1 U12396 ( .A(n15110), .ZN(n15131) );
  MUX2_X1 U12397 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12626), .Z(n9884) );
  XNOR2_X1 U12398 ( .A(n9884), .B(n9894), .ZN(n9821) );
  MUX2_X1 U12399 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12675), .Z(n9797) );
  OR2_X1 U12400 ( .A1(n9797), .A2(n10004), .ZN(n9819) );
  XOR2_X1 U12401 ( .A(n10004), .B(n9797), .Z(n9988) );
  NAND2_X1 U12402 ( .A1(n12626), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9800) );
  INV_X1 U12403 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9798) );
  OR2_X1 U12404 ( .A1(n12675), .A2(n9798), .ZN(n9799) );
  NAND2_X1 U12405 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  OR2_X1 U12406 ( .A1(n10163), .A2(n9801), .ZN(n9818) );
  XNOR2_X1 U12407 ( .A(n9801), .B(n9831), .ZN(n10161) );
  INV_X1 U12408 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9802) );
  OR2_X1 U12409 ( .A1(n6417), .A2(n9802), .ZN(n9804) );
  NAND2_X1 U12410 ( .A1(n6418), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U12411 ( .A1(n9804), .A2(n9803), .ZN(n9807) );
  XNOR2_X1 U12412 ( .A(n9807), .B(n10050), .ZN(n10042) );
  OR2_X1 U12413 ( .A1(n6418), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U12414 ( .A1(n6417), .A2(n9875), .ZN(n9805) );
  NAND2_X1 U12415 ( .A1(n9806), .A2(n9805), .ZN(n15085) );
  OAI22_X1 U12416 ( .A1(n10042), .A2(n15084), .B1(n10050), .B2(n9807), .ZN(
        n10011) );
  MUX2_X1 U12417 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6418), .Z(n9808) );
  XNOR2_X1 U12418 ( .A(n9808), .B(n10005), .ZN(n10012) );
  INV_X1 U12419 ( .A(n9808), .ZN(n9809) );
  AOI22_X1 U12420 ( .A1(n10011), .A2(n10012), .B1(n10005), .B2(n9809), .ZN(
        n10023) );
  INV_X1 U12421 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9810) );
  OR2_X1 U12422 ( .A1(n12626), .A2(n9810), .ZN(n9813) );
  NAND2_X1 U12423 ( .A1(n6417), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U12424 ( .A1(n9813), .A2(n9812), .ZN(n9815) );
  XOR2_X1 U12425 ( .A(n9814), .B(n9815), .Z(n10022) );
  INV_X1 U12426 ( .A(n9845), .ZN(n9817) );
  MUX2_X1 U12427 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12675), .Z(n9816) );
  XOR2_X1 U12428 ( .A(n9860), .B(n9816), .Z(n9844) );
  NAND2_X1 U12429 ( .A1(n10161), .A2(n10162), .ZN(n10160) );
  NAND2_X1 U12430 ( .A1(n9818), .A2(n10160), .ZN(n9987) );
  NAND2_X1 U12431 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  NAND2_X1 U12432 ( .A1(n9819), .A2(n9986), .ZN(n9820) );
  NAND2_X1 U12433 ( .A1(n9821), .A2(n9820), .ZN(n9885) );
  OAI21_X1 U12434 ( .B1(n9821), .B2(n9820), .A(n9885), .ZN(n9822) );
  NAND2_X1 U12435 ( .A1(n15131), .A2(n9822), .ZN(n9823) );
  NAND3_X1 U12436 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9841) );
  INV_X1 U12437 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U12438 ( .A1(n10004), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9834) );
  OAI21_X1 U12439 ( .B1(n10004), .B2(P3_REG2_REG_6__SCAN_IN), .A(n9834), .ZN(
        n9990) );
  AND2_X1 U12440 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n15268), .ZN(n9827) );
  NAND2_X1 U12441 ( .A1(n9828), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9826) );
  OAI21_X1 U12442 ( .B1(n9829), .B2(n10035), .A(n9850), .ZN(n10025) );
  INV_X1 U12443 ( .A(n10024), .ZN(n9852) );
  INV_X1 U12444 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10859) );
  XNOR2_X1 U12445 ( .A(n9860), .B(n10859), .ZN(n9851) );
  AOI21_X1 U12446 ( .B1(n9852), .B2(n9850), .A(n9851), .ZN(n9854) );
  NOR2_X1 U12447 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  AOI21_X1 U12448 ( .B1(n9836), .B2(n9835), .A(n9895), .ZN(n9839) );
  NOR2_X1 U12449 ( .A1(n9839), .A2(n15136), .ZN(n9840) );
  AOI211_X1 U12450 ( .C1(n15106), .C2(n9894), .A(n9841), .B(n9840), .ZN(n9842)
         );
  OAI21_X1 U12451 ( .B1(n9843), .B2(n15125), .A(n9842), .ZN(P3_U3189) );
  XNOR2_X1 U12452 ( .A(n9845), .B(n9844), .ZN(n9862) );
  OR3_X1 U12453 ( .A1(n10026), .A2(n9847), .A3(n9846), .ZN(n9848) );
  AND2_X1 U12454 ( .A1(n9849), .A2(n9848), .ZN(n9858) );
  AND3_X1 U12455 ( .A1(n9852), .A2(n9851), .A3(n9850), .ZN(n9853) );
  INV_X1 U12456 ( .A(n15136), .ZN(n12546) );
  OAI21_X1 U12457 ( .B1(n9854), .B2(n9853), .A(n12546), .ZN(n9857) );
  INV_X1 U12458 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U12459 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9855), .ZN(n10628) );
  AOI21_X1 U12460 ( .B1(n15082), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10628), .ZN(
        n9856) );
  OAI211_X1 U12461 ( .C1(n9858), .C2(n15125), .A(n9857), .B(n9856), .ZN(n9859)
         );
  AOI21_X1 U12462 ( .B1(n9860), .B2(n15106), .A(n9859), .ZN(n9861) );
  OAI21_X1 U12463 ( .B1(n9862), .B2(n15110), .A(n9861), .ZN(P3_U3186) );
  XNOR2_X1 U12464 ( .A(n12339), .B(n9863), .ZN(n9864) );
  NAND2_X1 U12465 ( .A1(n9864), .A2(n12854), .ZN(n9866) );
  AOI22_X1 U12466 ( .A1(n15145), .A2(n10856), .B1(n15143), .B2(n6689), .ZN(
        n9865) );
  NAND2_X1 U12467 ( .A1(n9866), .A2(n9865), .ZN(n10264) );
  AOI21_X1 U12468 ( .B1(n15177), .B2(n10263), .A(n10264), .ZN(n9923) );
  AOI22_X1 U12469 ( .A1(n8256), .A2(n10648), .B1(n15187), .B2(
        P3_REG0_REG_2__SCAN_IN), .ZN(n9867) );
  OAI21_X1 U12470 ( .B1(n15187), .B2(n9923), .A(n9867), .ZN(P3_U3396) );
  NAND2_X1 U12471 ( .A1(n8275), .A2(n10380), .ZN(n9874) );
  NAND2_X1 U12472 ( .A1(n9868), .A2(n15149), .ZN(n9870) );
  OR2_X1 U12473 ( .A1(n9869), .A2(n10380), .ZN(n12333) );
  NAND2_X1 U12474 ( .A1(n12333), .A2(n15140), .ZN(n10379) );
  NAND2_X1 U12475 ( .A1(n9870), .A2(n10379), .ZN(n9872) );
  NAND2_X1 U12476 ( .A1(n15145), .A2(n6689), .ZN(n9871) );
  NAND2_X1 U12477 ( .A1(n9872), .A2(n9871), .ZN(n10237) );
  NAND2_X1 U12478 ( .A1(n15199), .A2(n10237), .ZN(n9873) );
  OAI211_X1 U12479 ( .C1(n15199), .C2(n9875), .A(n9874), .B(n9873), .ZN(
        P3_U3459) );
  NAND2_X1 U12480 ( .A1(n10335), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10327) );
  OAI21_X1 U12481 ( .B1(n10335), .B2(P3_REG1_REG_8__SCAN_IN), .A(n10327), .ZN(
        n9879) );
  INV_X1 U12482 ( .A(n10328), .ZN(n9878) );
  AOI21_X1 U12483 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9904) );
  INV_X1 U12484 ( .A(n10335), .ZN(n9902) );
  NAND2_X1 U12485 ( .A1(n15082), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n9892) );
  INV_X1 U12486 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10763) );
  OR2_X1 U12487 ( .A1(n12626), .A2(n10763), .ZN(n9882) );
  NAND2_X1 U12488 ( .A1(n12675), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U12489 ( .A1(n9882), .A2(n9881), .ZN(n10336) );
  XNOR2_X1 U12490 ( .A(n10336), .B(n9902), .ZN(n9888) );
  OR2_X1 U12491 ( .A1(n9884), .A2(n9883), .ZN(n9886) );
  NAND2_X1 U12492 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  NAND2_X1 U12493 ( .A1(n9888), .A2(n9887), .ZN(n10334) );
  OAI21_X1 U12494 ( .B1(n9888), .B2(n9887), .A(n10334), .ZN(n9890) );
  NOR2_X1 U12495 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9889), .ZN(n10678) );
  AOI21_X1 U12496 ( .B1(n15131), .B2(n9890), .A(n10678), .ZN(n9891) );
  NAND2_X1 U12497 ( .A1(n9892), .A2(n9891), .ZN(n9901) );
  NOR2_X1 U12498 ( .A1(n9894), .A2(n9893), .ZN(n9896) );
  NAND2_X1 U12499 ( .A1(n10335), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10341) );
  OAI21_X1 U12500 ( .B1(n10335), .B2(P3_REG2_REG_8__SCAN_IN), .A(n10341), .ZN(
        n9897) );
  NAND2_X1 U12501 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  AOI21_X1 U12502 ( .B1(n10342), .B2(n9899), .A(n15136), .ZN(n9900) );
  AOI211_X1 U12503 ( .C1(n15106), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9903)
         );
  OAI21_X1 U12504 ( .B1(n9904), .B2(n15125), .A(n9903), .ZN(P3_U3190) );
  XNOR2_X1 U12505 ( .A(n11878), .B(n9905), .ZN(n14715) );
  NAND2_X1 U12506 ( .A1(n13967), .A2(n13966), .ZN(n9909) );
  NAND2_X1 U12507 ( .A1(n14700), .A2(n14762), .ZN(n14114) );
  NOR2_X1 U12508 ( .A1(n14717), .A2(n9906), .ZN(n9907) );
  NOR2_X1 U12509 ( .A1(n9908), .A2(n9907), .ZN(n14716) );
  OR2_X1 U12510 ( .A1(n9909), .A2(n14184), .ZN(n14173) );
  NOR2_X1 U12511 ( .A1(n14173), .A2(n14718), .ZN(n14013) );
  OAI22_X1 U12512 ( .A1(n14700), .A2(n9309), .B1(n9910), .B2(n14698), .ZN(
        n9912) );
  NAND2_X1 U12513 ( .A1(n14700), .A2(n14470), .ZN(n14101) );
  NOR2_X1 U12514 ( .A1(n14101), .A2(n14717), .ZN(n9911) );
  AOI211_X1 U12515 ( .C1(n14716), .C2(n14013), .A(n9912), .B(n9911), .ZN(n9920) );
  XNOR2_X1 U12516 ( .A(n14716), .B(n13837), .ZN(n9915) );
  INV_X1 U12517 ( .A(n11878), .ZN(n9913) );
  NOR2_X1 U12518 ( .A1(n9913), .A2(n14572), .ZN(n9914) );
  MUX2_X1 U12519 ( .A(n9915), .B(n9914), .S(n13838), .Z(n9918) );
  AOI21_X1 U12520 ( .B1(n13838), .B2(n14572), .A(n14751), .ZN(n9917) );
  OAI21_X1 U12521 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n14720) );
  NAND2_X1 U12522 ( .A1(n14700), .A2(n14720), .ZN(n9919) );
  OAI211_X1 U12523 ( .C1(n14715), .C2(n14114), .A(n9920), .B(n9919), .ZN(
        P1_U3292) );
  OAI22_X1 U12524 ( .A1(n12933), .A2(n12349), .B1(n15199), .B2(n9777), .ZN(
        n9921) );
  INV_X1 U12525 ( .A(n9921), .ZN(n9922) );
  OAI21_X1 U12526 ( .B1(n9923), .B2(n15196), .A(n9922), .ZN(P3_U3461) );
  OR2_X1 U12527 ( .A1(n11552), .A2(n13836), .ZN(n11544) );
  OR2_X1 U12528 ( .A1(n9926), .A2(n10072), .ZN(n9928) );
  AOI22_X1 U12529 ( .A1(n6422), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11659), 
        .B2(n13863), .ZN(n9927) );
  NAND2_X1 U12530 ( .A1(n10185), .A2(n14705), .ZN(n11558) );
  INV_X1 U12531 ( .A(n10185), .ZN(n13835) );
  NAND2_X1 U12532 ( .A1(n14695), .A2(n14694), .ZN(n9929) );
  OR2_X1 U12533 ( .A1(n9930), .A2(n10072), .ZN(n9932) );
  AOI22_X1 U12534 ( .A1(n11660), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11659), 
        .B2(n13880), .ZN(n9931) );
  NAND2_X1 U12535 ( .A1(n9932), .A2(n9931), .ZN(n11565) );
  NAND2_X1 U12536 ( .A1(n11707), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9937) );
  XNOR2_X1 U12537 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10256) );
  OR2_X1 U12538 ( .A1(n11818), .A2(n10256), .ZN(n9935) );
  OR2_X1 U12539 ( .A1(n11820), .A2(n9313), .ZN(n9934) );
  NAND4_X2 U12540 ( .A1(n9937), .A2(n9935), .A3(n9934), .A4(n9936), .ZN(n13834) );
  NAND2_X1 U12541 ( .A1(n10112), .A2(n7314), .ZN(n9939) );
  NAND2_X1 U12542 ( .A1(n11565), .A2(n10253), .ZN(n9938) );
  NAND2_X1 U12543 ( .A1(n9940), .A2(n9925), .ZN(n9942) );
  AOI22_X1 U12544 ( .A1(n11660), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11659), 
        .B2(n13892), .ZN(n9941) );
  AOI21_X1 U12545 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U12546 ( .A1(n9943), .A2(n9957), .ZN(n13744) );
  NAND2_X1 U12547 ( .A1(n11706), .A2(n13744), .ZN(n9950) );
  OR2_X1 U12548 ( .A1(n6802), .A2(n9967), .ZN(n9949) );
  INV_X1 U12549 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9945) );
  OR2_X1 U12550 ( .A1(n11797), .A2(n9945), .ZN(n9948) );
  OR2_X1 U12551 ( .A1(n11820), .A2(n9946), .ZN(n9947) );
  XNOR2_X1 U12552 ( .A(n13743), .B(n6845), .ZN(n11881) );
  INV_X1 U12553 ( .A(n11881), .ZN(n10089) );
  XNOR2_X1 U12554 ( .A(n10090), .B(n10089), .ZN(n9965) );
  NAND2_X1 U12555 ( .A1(n9952), .A2(n9951), .ZN(n9954) );
  NAND2_X1 U12556 ( .A1(n11556), .A2(n11552), .ZN(n9953) );
  INV_X1 U12557 ( .A(n14694), .ZN(n14703) );
  NAND2_X1 U12558 ( .A1(n6990), .A2(n10185), .ZN(n9955) );
  INV_X1 U12559 ( .A(n11565), .ZN(n14731) );
  NAND2_X1 U12560 ( .A1(n14731), .A2(n10253), .ZN(n9956) );
  XNOR2_X1 U12561 ( .A(n10069), .B(n10089), .ZN(n9963) );
  NAND2_X1 U12562 ( .A1(n11707), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9961) );
  OR2_X1 U12563 ( .A1(n11820), .A2(n9316), .ZN(n9960) );
  OAI21_X1 U12564 ( .B1(n9957), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10083), .ZN(
        n10517) );
  OR2_X1 U12565 ( .A1(n11818), .A2(n10517), .ZN(n9959) );
  OR2_X1 U12566 ( .A1(n6802), .A2(n10135), .ZN(n9958) );
  NAND4_X1 U12567 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n13832) );
  AOI22_X1 U12568 ( .A1(n14572), .A2(n13834), .B1(n13832), .B2(n14575), .ZN(
        n9962) );
  OAI21_X1 U12569 ( .B1(n9963), .B2(n14609), .A(n9962), .ZN(n9964) );
  AOI21_X1 U12570 ( .B1(n14751), .B2(n9965), .A(n9964), .ZN(n10209) );
  INV_X1 U12571 ( .A(n13743), .ZN(n10065) );
  INV_X1 U12572 ( .A(n10123), .ZN(n9966) );
  OAI211_X1 U12573 ( .C1(n10065), .C2(n10116), .A(n9966), .B(n14707), .ZN(
        n10204) );
  NAND2_X1 U12574 ( .A1(n10209), .A2(n10204), .ZN(n10067) );
  OAI22_X1 U12575 ( .A1(n14259), .A2(n10065), .B1(n14772), .B2(n9967), .ZN(
        n9968) );
  AOI21_X1 U12576 ( .B1(n10067), .B2(n14772), .A(n9968), .ZN(n9969) );
  INV_X1 U12577 ( .A(n9969), .ZN(P1_U3533) );
  AOI21_X1 U12578 ( .B1(n9975), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9970), .ZN(
        n14867) );
  MUX2_X1 U12579 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8612), .S(n14861), .Z(
        n14868) );
  NAND2_X1 U12580 ( .A1(n14867), .A2(n14868), .ZN(n14866) );
  OAI21_X1 U12581 ( .B1(n14861), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14866), 
        .ZN(n9973) );
  INV_X1 U12582 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13229) );
  MUX2_X1 U12583 ( .A(n13229), .B(P2_REG1_REG_13__SCAN_IN), .S(n9976), .Z(
        n9972) );
  INV_X1 U12584 ( .A(n13227), .ZN(n9971) );
  AOI211_X1 U12585 ( .C1(n9973), .C2(n9972), .A(n13246), .B(n9971), .ZN(n9982)
         );
  OAI21_X1 U12586 ( .B1(n9975), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9974), .ZN(
        n14863) );
  MUX2_X1 U12587 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8615), .S(n14861), .Z(
        n14864) );
  NAND2_X1 U12588 ( .A1(n14863), .A2(n14864), .ZN(n14862) );
  OAI21_X1 U12589 ( .B1(n14861), .B2(P2_REG2_REG_12__SCAN_IN), .A(n14862), 
        .ZN(n9978) );
  MUX2_X1 U12590 ( .A(n13217), .B(P2_REG2_REG_13__SCAN_IN), .S(n9976), .Z(
        n9977) );
  NOR2_X1 U12591 ( .A1(n9978), .A2(n9977), .ZN(n13215) );
  AOI211_X1 U12592 ( .C1(n9978), .C2(n9977), .A(n14853), .B(n13215), .ZN(n9981) );
  NAND2_X1 U12593 ( .A1(n14923), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U12594 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14785)
         );
  OAI211_X1 U12595 ( .C1(n14930), .C2(n13228), .A(n9979), .B(n14785), .ZN(
        n9980) );
  OR3_X1 U12596 ( .A1(n9982), .A2(n9981), .A3(n9980), .ZN(P2_U3227) );
  INV_X1 U12597 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12598 ( .A1(n8256), .A2(n10380), .ZN(n9984) );
  NAND2_X1 U12599 ( .A1(n15185), .A2(n10237), .ZN(n9983) );
  OAI211_X1 U12600 ( .C1(n9985), .C2(n15185), .A(n9984), .B(n9983), .ZN(
        P3_U3390) );
  OAI21_X1 U12601 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n10002) );
  AOI21_X1 U12602 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9996) );
  AOI21_X1 U12603 ( .B1(n9994), .B2(n9993), .A(n9992), .ZN(n9995) );
  OAI22_X1 U12604 ( .A1(n9996), .A2(n15136), .B1(n15125), .B2(n9995), .ZN(
        n10001) );
  INV_X1 U12605 ( .A(n15082), .ZN(n15126) );
  INV_X1 U12606 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9999) );
  INV_X1 U12607 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9997) );
  NOR2_X1 U12608 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9997), .ZN(n10467) );
  INV_X1 U12609 ( .A(n10467), .ZN(n9998) );
  OAI21_X1 U12610 ( .B1(n15126), .B2(n9999), .A(n9998), .ZN(n10000) );
  AOI211_X1 U12611 ( .C1(n15131), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10003) );
  OAI21_X1 U12612 ( .B1(n10004), .B2(n15122), .A(n10003), .ZN(P3_U3188) );
  INV_X1 U12613 ( .A(n10005), .ZN(n10021) );
  OAI21_X1 U12614 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10019) );
  AOI21_X1 U12615 ( .B1(n10010), .B2(n10009), .A(n6607), .ZN(n10014) );
  XOR2_X1 U12616 ( .A(n10012), .B(n10011), .Z(n10013) );
  OAI22_X1 U12617 ( .A1(n15136), .A2(n10014), .B1(n10013), .B2(n15110), .ZN(
        n10018) );
  INV_X1 U12618 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10015) );
  OAI22_X1 U12619 ( .A1(n15126), .A2(n10016), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10015), .ZN(n10017) );
  AOI211_X1 U12620 ( .C1(n6983), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10020) );
  OAI21_X1 U12621 ( .B1(n10021), .B2(n15122), .A(n10020), .ZN(P3_U3184) );
  XNOR2_X1 U12622 ( .A(n10023), .B(n10022), .ZN(n10033) );
  AOI21_X1 U12623 ( .B1(n9810), .B2(n10025), .A(n10024), .ZN(n10031) );
  NOR2_X1 U12624 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10532), .ZN(n10527) );
  AOI21_X1 U12625 ( .B1(n15190), .B2(n10027), .A(n10026), .ZN(n10028) );
  NOR2_X1 U12626 ( .A1(n15125), .A2(n10028), .ZN(n10029) );
  AOI211_X1 U12627 ( .C1(n15082), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10527), .B(
        n10029), .ZN(n10030) );
  OAI21_X1 U12628 ( .B1(n10031), .B2(n15136), .A(n10030), .ZN(n10032) );
  AOI21_X1 U12629 ( .B1(n15131), .B2(n10033), .A(n10032), .ZN(n10034) );
  OAI21_X1 U12630 ( .B1(n10035), .B2(n15122), .A(n10034), .ZN(P3_U3185) );
  NAND2_X1 U12631 ( .A1(n10036), .A2(n15188), .ZN(n10037) );
  NAND2_X1 U12632 ( .A1(n10038), .A2(n10037), .ZN(n10048) );
  AOI21_X1 U12633 ( .B1(n9802), .B2(n10040), .A(n10039), .ZN(n10041) );
  NOR2_X1 U12634 ( .A1(n15136), .A2(n10041), .ZN(n10047) );
  INV_X1 U12635 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U12636 ( .A1(n15082), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10045) );
  XNOR2_X1 U12637 ( .A(n10042), .B(n15084), .ZN(n10043) );
  NAND2_X1 U12638 ( .A1(n15131), .A2(n10043), .ZN(n10044) );
  OAI211_X1 U12639 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10815), .A(n10045), .B(
        n10044), .ZN(n10046) );
  AOI211_X1 U12640 ( .C1(n6983), .C2(n10048), .A(n10047), .B(n10046), .ZN(
        n10049) );
  OAI21_X1 U12641 ( .B1(n10050), .B2(n15122), .A(n10049), .ZN(P3_U3183) );
  OAI22_X1 U12642 ( .A1(n14173), .A2(n10052), .B1(n10051), .B2(n14698), .ZN(
        n10055) );
  MUX2_X1 U12643 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10053), .S(n14700), .Z(
        n10054) );
  AOI211_X1 U12644 ( .C1(n14702), .C2(n11542), .A(n10055), .B(n10054), .ZN(
        n10056) );
  INV_X1 U12645 ( .A(n10056), .ZN(P1_U3291) );
  NAND2_X1 U12646 ( .A1(n14764), .A2(n14755), .ZN(n14300) );
  OAI22_X1 U12647 ( .A1(n14300), .A2(n11552), .B1(n14764), .B2(n9597), .ZN(
        n10057) );
  AOI21_X1 U12648 ( .B1(n14764), .B2(n10058), .A(n10057), .ZN(n10059) );
  INV_X1 U12649 ( .A(n10059), .ZN(P1_U3465) );
  INV_X1 U12650 ( .A(n11631), .ZN(n10064) );
  INV_X1 U12651 ( .A(n13239), .ZN(n14929) );
  OAI222_X1 U12652 ( .A1(n11238), .A2(n10060), .B1(n13688), .B2(n10064), .C1(
        n14929), .C2(P2_U3088), .ZN(P2_U3309) );
  OAI21_X1 U12653 ( .B1(n10061), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10062) );
  XNOR2_X1 U12654 ( .A(n10062), .B(P1_IR_REG_18__SCAN_IN), .ZN(n11632) );
  INV_X1 U12655 ( .A(n11632), .ZN(n11030) );
  OAI222_X1 U12656 ( .A1(P1_U3086), .A2(n11030), .B1(n11530), .B2(n10064), 
        .C1(n10063), .C2(n6421), .ZN(P1_U3337) );
  OAI22_X1 U12657 ( .A1(n14300), .A2(n10065), .B1(n14764), .B2(n9945), .ZN(
        n10066) );
  AOI21_X1 U12658 ( .B1(n10067), .B2(n14764), .A(n10066), .ZN(n10068) );
  INV_X1 U12659 ( .A(n10068), .ZN(P1_U3474) );
  NAND2_X1 U12660 ( .A1(n10069), .A2(n11881), .ZN(n10071) );
  OR2_X1 U12661 ( .A1(n13743), .A2(n13833), .ZN(n10070) );
  INV_X2 U12662 ( .A(n10072), .ZN(n11791) );
  AOI22_X1 U12663 ( .A1(n11660), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11659), 
        .B2(n10074), .ZN(n10075) );
  INV_X1 U12664 ( .A(n13832), .ZN(n13741) );
  XNOR2_X1 U12665 ( .A(n11578), .B(n13741), .ZN(n11882) );
  NAND2_X1 U12666 ( .A1(n10125), .A2(n11882), .ZN(n10077) );
  OR2_X1 U12667 ( .A1(n11578), .A2(n13832), .ZN(n10076) );
  AOI22_X1 U12668 ( .A1(n11660), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11659), 
        .B2(n10079), .ZN(n10080) );
  NAND2_X1 U12669 ( .A1(n11817), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10088) );
  INV_X1 U12670 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10081) );
  OR2_X1 U12671 ( .A1(n11797), .A2(n10081), .ZN(n10087) );
  AND2_X1 U12672 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  OR2_X1 U12673 ( .A1(n10084), .A2(n10095), .ZN(n10792) );
  OR2_X1 U12674 ( .A1(n11818), .A2(n10792), .ZN(n10086) );
  OR2_X1 U12675 ( .A1(n11820), .A2(n9317), .ZN(n10085) );
  NAND4_X1 U12676 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n13831) );
  XNOR2_X1 U12677 ( .A(n10271), .B(n11883), .ZN(n10105) );
  NAND2_X1 U12678 ( .A1(n13743), .A2(n6845), .ZN(n10091) );
  INV_X1 U12679 ( .A(n11882), .ZN(n10124) );
  NAND2_X1 U12680 ( .A1(n11578), .A2(n13741), .ZN(n10092) );
  XNOR2_X1 U12681 ( .A(n10279), .B(n11883), .ZN(n10103) );
  NAND2_X1 U12682 ( .A1(n11707), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10101) );
  INV_X1 U12683 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10094) );
  OR2_X1 U12684 ( .A1(n6802), .A2(n10094), .ZN(n10100) );
  NAND2_X1 U12685 ( .A1(n10095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10284) );
  OR2_X1 U12686 ( .A1(n10095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12687 ( .A1(n10284), .A2(n10096), .ZN(n11013) );
  OR2_X1 U12688 ( .A1(n11818), .A2(n11013), .ZN(n10099) );
  OR2_X1 U12689 ( .A1(n11820), .A2(n10097), .ZN(n10098) );
  NAND4_X1 U12690 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n13830) );
  INV_X1 U12691 ( .A(n13830), .ZN(n10795) );
  OAI22_X1 U12692 ( .A1(n10795), .A2(n11394), .B1(n13741), .B2(n14165), .ZN(
        n10102) );
  AOI21_X1 U12693 ( .B1(n10103), .B2(n14751), .A(n10102), .ZN(n10104) );
  OAI21_X1 U12694 ( .B1(n10105), .B2(n14609), .A(n10104), .ZN(n10298) );
  INV_X1 U12695 ( .A(n11578), .ZN(n10138) );
  AOI211_X1 U12696 ( .C1(n11587), .C2(n10122), .A(n14718), .B(n10277), .ZN(
        n10301) );
  NOR2_X1 U12697 ( .A1(n10298), .A2(n10301), .ZN(n10110) );
  INV_X1 U12698 ( .A(n11587), .ZN(n10297) );
  OAI22_X1 U12699 ( .A1(n14259), .A2(n10297), .B1(n14772), .B2(n9298), .ZN(
        n10106) );
  INV_X1 U12700 ( .A(n10106), .ZN(n10107) );
  OAI21_X1 U12701 ( .B1(n10110), .B2(n6820), .A(n10107), .ZN(P1_U3535) );
  OAI22_X1 U12702 ( .A1(n14300), .A2(n10297), .B1(n14764), .B2(n10081), .ZN(
        n10108) );
  INV_X1 U12703 ( .A(n10108), .ZN(n10109) );
  OAI21_X1 U12704 ( .B1(n10110), .B2(n14763), .A(n10109), .ZN(P1_U3480) );
  XNOR2_X1 U12705 ( .A(n11880), .B(n10111), .ZN(n14734) );
  INV_X1 U12706 ( .A(n14114), .ZN(n14712) );
  AOI22_X1 U12707 ( .A1(n14734), .A2(n14712), .B1(n14702), .B2(n11565), .ZN(
        n10121) );
  XNOR2_X1 U12708 ( .A(n10112), .B(n7314), .ZN(n10113) );
  NAND2_X1 U12709 ( .A1(n10113), .A2(n14751), .ZN(n10115) );
  AOI22_X1 U12710 ( .A1(n13835), .A2(n14572), .B1(n14575), .B2(n13833), .ZN(
        n10114) );
  NAND2_X1 U12711 ( .A1(n10115), .A2(n10114), .ZN(n14732) );
  INV_X1 U12712 ( .A(n10116), .ZN(n10117) );
  OAI211_X1 U12713 ( .C1(n14731), .C2(n14710), .A(n10117), .B(n14707), .ZN(
        n14730) );
  OAI22_X1 U12714 ( .A1(n14730), .A2(n14184), .B1(n14698), .B2(n10256), .ZN(
        n10118) );
  NOR2_X1 U12715 ( .A1(n14732), .A2(n10118), .ZN(n10119) );
  MUX2_X1 U12716 ( .A(n9313), .B(n10119), .S(n14700), .Z(n10120) );
  NAND2_X1 U12717 ( .A1(n10121), .A2(n10120), .ZN(P1_U3289) );
  OAI211_X1 U12718 ( .C1(n10138), .C2(n10123), .A(n14707), .B(n10122), .ZN(
        n10133) );
  XNOR2_X1 U12719 ( .A(n10125), .B(n10124), .ZN(n10127) );
  AOI22_X1 U12720 ( .A1(n14572), .A2(n13833), .B1(n13831), .B2(n14575), .ZN(
        n10126) );
  OAI21_X1 U12721 ( .B1(n10127), .B2(n14609), .A(n10126), .ZN(n10128) );
  AOI21_X1 U12722 ( .B1(n14751), .B2(n10129), .A(n10128), .ZN(n10134) );
  MUX2_X1 U12723 ( .A(n9316), .B(n10134), .S(n14700), .Z(n10132) );
  INV_X1 U12724 ( .A(n10517), .ZN(n10130) );
  INV_X1 U12725 ( .A(n14698), .ZN(n14683) );
  AOI22_X1 U12726 ( .A1(n14702), .A2(n11578), .B1(n10130), .B2(n14683), .ZN(
        n10131) );
  OAI211_X1 U12727 ( .C1(n14173), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        P1_U3287) );
  NAND2_X1 U12728 ( .A1(n10134), .A2(n10133), .ZN(n10140) );
  OAI22_X1 U12729 ( .A1(n14259), .A2(n10138), .B1(n14772), .B2(n10135), .ZN(
        n10136) );
  AOI21_X1 U12730 ( .B1(n10140), .B2(n14772), .A(n10136), .ZN(n10137) );
  INV_X1 U12731 ( .A(n10137), .ZN(P1_U3534) );
  INV_X1 U12732 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15310) );
  OAI22_X1 U12733 ( .A1(n14300), .A2(n10138), .B1(n14764), .B2(n15310), .ZN(
        n10139) );
  AOI21_X1 U12734 ( .B1(n10140), .B2(n14764), .A(n10139), .ZN(n10141) );
  INV_X1 U12735 ( .A(n10141), .ZN(P1_U3477) );
  INV_X2 U12736 ( .A(n15078), .ZN(n15081) );
  NAND2_X1 U12737 ( .A1(n13146), .A2(n13530), .ZN(n13537) );
  NAND2_X1 U12738 ( .A1(n13538), .A2(n13537), .ZN(n13536) );
  INV_X1 U12739 ( .A(n6413), .ZN(n10147) );
  INV_X1 U12740 ( .A(n9053), .ZN(n13532) );
  NAND2_X1 U12741 ( .A1(n10147), .A2(n13532), .ZN(n10142) );
  NAND2_X1 U12742 ( .A1(n13536), .A2(n10142), .ZN(n10605) );
  NAND2_X1 U12743 ( .A1(n10605), .A2(n10604), .ZN(n10607) );
  INV_X1 U12744 ( .A(n13144), .ZN(n10150) );
  NAND2_X1 U12745 ( .A1(n10150), .A2(n9052), .ZN(n10143) );
  NAND2_X1 U12746 ( .A1(n10607), .A2(n10143), .ZN(n10384) );
  XNOR2_X1 U12747 ( .A(n10384), .B(n10383), .ZN(n10377) );
  NAND2_X1 U12748 ( .A1(n10377), .A2(n14999), .ZN(n10158) );
  NAND2_X1 U12749 ( .A1(n13142), .A2(n13254), .ZN(n10146) );
  OR2_X1 U12750 ( .A1(n10144), .A2(n6427), .ZN(n13508) );
  NAND2_X1 U12751 ( .A1(n13144), .A2(n13116), .ZN(n10145) );
  NAND2_X1 U12752 ( .A1(n10146), .A2(n10145), .ZN(n14774) );
  AOI21_X1 U12753 ( .B1(n15053), .B2(n14783), .A(n14774), .ZN(n10157) );
  NAND2_X1 U12754 ( .A1(n13540), .A2(n13539), .ZN(n10149) );
  NAND2_X1 U12755 ( .A1(n10147), .A2(n9053), .ZN(n10148) );
  NAND2_X1 U12756 ( .A1(n10149), .A2(n10148), .ZN(n10610) );
  NAND2_X1 U12757 ( .A1(n10150), .A2(n10621), .ZN(n10151) );
  OR2_X1 U12758 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NAND2_X1 U12759 ( .A1(n10545), .A2(n10154), .ZN(n10155) );
  NAND2_X1 U12760 ( .A1(n10155), .A2(n15026), .ZN(n10373) );
  INV_X1 U12761 ( .A(n14783), .ZN(n10385) );
  INV_X1 U12762 ( .A(n10538), .ZN(n10156) );
  OAI211_X1 U12763 ( .C1(n10385), .C2(n10616), .A(n10156), .B(n13496), .ZN(
        n10371) );
  NAND4_X1 U12764 ( .A1(n10158), .A2(n10157), .A3(n10373), .A4(n10371), .ZN(
        n10202) );
  NAND2_X1 U12765 ( .A1(n10202), .A2(n15081), .ZN(n10159) );
  OAI21_X1 U12766 ( .B1(n15081), .B2(n9355), .A(n10159), .ZN(P2_U3502) );
  OAI21_X1 U12767 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10173) );
  NOR2_X1 U12768 ( .A1(n15122), .A2(n10163), .ZN(n10172) );
  AOI21_X1 U12769 ( .B1(n10165), .B2(n10221), .A(n10164), .ZN(n10170) );
  OAI21_X1 U12770 ( .B1(n10167), .B2(n10166), .A(n12546), .ZN(n10169) );
  AND2_X1 U12771 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10637) );
  AOI21_X1 U12772 ( .B1(n15082), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10637), .ZN(
        n10168) );
  OAI211_X1 U12773 ( .C1(n10170), .C2(n15125), .A(n10169), .B(n10168), .ZN(
        n10171) );
  AOI211_X1 U12774 ( .C1(n15131), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10174) );
  INV_X1 U12775 ( .A(n10174), .ZN(P3_U3187) );
  AND2_X1 U12776 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U12777 ( .A1(n9560), .A2(n10177), .ZN(n11916) );
  INV_X1 U12778 ( .A(n11916), .ZN(n10178) );
  NAND2_X1 U12779 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  NAND2_X1 U12780 ( .A1(n10180), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14568) );
  INV_X1 U12781 ( .A(n14568), .ZN(n13817) );
  INV_X1 U12782 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13857) );
  NAND2_X1 U12783 ( .A1(n13836), .A2(n14572), .ZN(n10182) );
  NAND2_X1 U12784 ( .A1(n13834), .A2(n14575), .ZN(n10181) );
  NAND2_X1 U12785 ( .A1(n10182), .A2(n10181), .ZN(n14696) );
  AOI22_X1 U12786 ( .A1(n13805), .A2(n14696), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10183) );
  OAI21_X1 U12787 ( .B1(n13821), .B2(n6990), .A(n10183), .ZN(n10196) );
  OAI22_X1 U12788 ( .A1(n10184), .A2(n10185), .B1(n6990), .B2(n12047), .ZN(
        n10251) );
  XNOR2_X1 U12789 ( .A(n10250), .B(n10251), .ZN(n10194) );
  AOI211_X1 U12790 ( .C1(n10194), .C2(n10193), .A(n14559), .B(n10192), .ZN(
        n10195) );
  AOI211_X1 U12791 ( .C1(n13817), .C2(n13857), .A(n10196), .B(n10195), .ZN(
        n10197) );
  INV_X1 U12792 ( .A(n10197), .ZN(P1_U3218) );
  NAND3_X1 U12793 ( .A1(n14979), .A2(n10199), .A3(n10198), .ZN(n10200) );
  NOR2_X1 U12794 ( .A1(n10365), .A2(n10200), .ZN(n10201) );
  AND2_X2 U12795 ( .A1(n10201), .A2(n14978), .ZN(n15066) );
  NAND2_X1 U12796 ( .A1(n10202), .A2(n15066), .ZN(n10203) );
  OAI21_X1 U12797 ( .B1(n15066), .B2(n8390), .A(n10203), .ZN(P2_U3439) );
  INV_X2 U12798 ( .A(n14700), .ZN(n14684) );
  NOR2_X1 U12799 ( .A1(n14173), .A2(n10204), .ZN(n10207) );
  INV_X1 U12800 ( .A(n13744), .ZN(n10205) );
  OAI22_X1 U12801 ( .A1(n14700), .A2(n9946), .B1(n10205), .B2(n14698), .ZN(
        n10206) );
  AOI211_X1 U12802 ( .C1(n14702), .C2(n13743), .A(n10207), .B(n10206), .ZN(
        n10208) );
  OAI21_X1 U12803 ( .B1(n10209), .B2(n14684), .A(n10208), .ZN(P1_U3288) );
  INV_X1 U12804 ( .A(n11658), .ZN(n10211) );
  OAI222_X1 U12805 ( .A1(n11238), .A2(n15215), .B1(n13688), .B2(n10211), .C1(
        n10369), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U12806 ( .A1(P1_U3086), .A2(n14471), .B1(n11530), .B2(n10211), 
        .C1(n10210), .C2(n6421), .ZN(P1_U3336) );
  OAI21_X1 U12807 ( .B1(n10213), .B2(n12366), .A(n10212), .ZN(n10464) );
  INV_X1 U12808 ( .A(n10214), .ZN(n10215) );
  AOI21_X1 U12809 ( .B1(n12366), .B2(n10216), .A(n10215), .ZN(n10217) );
  OAI222_X1 U12810 ( .A1(n12873), .A2(n10437), .B1(n12875), .B2(n10641), .C1(
        n15149), .C2(n10217), .ZN(n10461) );
  AOI21_X1 U12811 ( .B1(n15177), .B2(n10464), .A(n10461), .ZN(n10225) );
  INV_X1 U12812 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10218) );
  OAI22_X1 U12813 ( .A1(n10222), .A2(n12981), .B1(n15185), .B2(n10218), .ZN(
        n10219) );
  INV_X1 U12814 ( .A(n10219), .ZN(n10220) );
  OAI21_X1 U12815 ( .B1(n10225), .B2(n15187), .A(n10220), .ZN(P3_U3405) );
  OAI22_X1 U12816 ( .A1(n12933), .A2(n10222), .B1(n15199), .B2(n10221), .ZN(
        n10223) );
  INV_X1 U12817 ( .A(n10223), .ZN(n10224) );
  OAI21_X1 U12818 ( .B1(n10225), .B2(n15196), .A(n10224), .ZN(P3_U3464) );
  OAI21_X1 U12819 ( .B1(n14013), .B2(n14702), .A(n9584), .ZN(n10230) );
  INV_X1 U12820 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10226) );
  OAI22_X1 U12821 ( .A1(n14684), .A2(n10227), .B1(n10226), .B2(n14698), .ZN(
        n10228) );
  INV_X1 U12822 ( .A(n10228), .ZN(n10229) );
  OAI211_X1 U12823 ( .C1(n9284), .C2(n14700), .A(n10230), .B(n10229), .ZN(
        P1_U3293) );
  NAND2_X1 U12824 ( .A1(n10232), .A2(n10231), .ZN(n10235) );
  NAND2_X1 U12825 ( .A1(n10233), .A2(n12985), .ZN(n10234) );
  NAND3_X1 U12826 ( .A1(n10236), .A2(n10235), .A3(n10234), .ZN(n10239) );
  INV_X2 U12827 ( .A(n15154), .ZN(n15156) );
  AOI21_X1 U12828 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15151), .A(n10237), .ZN(
        n10241) );
  NAND2_X1 U12829 ( .A1(n15184), .A2(n15150), .ZN(n10238) );
  INV_X1 U12830 ( .A(n12883), .ZN(n12741) );
  AOI22_X1 U12831 ( .A1(n15156), .A2(P3_REG2_REG_0__SCAN_IN), .B1(n12741), 
        .B2(n10380), .ZN(n10240) );
  OAI21_X1 U12832 ( .B1(n15156), .B2(n10241), .A(n10240), .ZN(P3_U3233) );
  INV_X1 U12833 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U12834 ( .A1(n6457), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U12835 ( .A1(n8215), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U12836 ( .A1(n8216), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10242) );
  AND3_X1 U12837 ( .A1(n10244), .A2(n10243), .A3(n10242), .ZN(n10245) );
  AND2_X1 U12838 ( .A1(n10246), .A2(n10245), .ZN(n12690) );
  NAND2_X1 U12839 ( .A1(n6738), .A2(P3_U3897), .ZN(n10247) );
  OAI21_X1 U12840 ( .B1(P3_U3897), .B2(n15297), .A(n10247), .ZN(P3_U3522) );
  OAI222_X1 U12841 ( .A1(n14451), .A2(n10249), .B1(n12997), .B2(n10248), .C1(
        P3_U3151), .C2(n8101), .ZN(P3_U3274) );
  OAI22_X1 U12842 ( .A1(n10184), .A2(n10253), .B1(n14731), .B2(n12047), .ZN(
        n10503) );
  AOI22_X1 U12843 ( .A1(n12122), .A2(n13834), .B1(n12129), .B2(n11565), .ZN(
        n10255) );
  XOR2_X1 U12844 ( .A(n12130), .B(n10255), .Z(n10504) );
  XNOR2_X1 U12845 ( .A(n10505), .B(n10504), .ZN(n10260) );
  NAND2_X1 U12846 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13871) );
  OAI21_X1 U12847 ( .B1(n14551), .B2(n6845), .A(n13871), .ZN(n10258) );
  OAI22_X1 U12848 ( .A1(n13821), .A2(n14731), .B1(n14568), .B2(n10256), .ZN(
        n10257) );
  AOI211_X1 U12849 ( .C1(n13794), .C2(n13835), .A(n10258), .B(n10257), .ZN(
        n10259) );
  OAI21_X1 U12850 ( .B1(n10260), .B2(n14559), .A(n10259), .ZN(P1_U3230) );
  NOR2_X1 U12851 ( .A1(n8101), .A2(n15150), .ZN(n10261) );
  NAND2_X1 U12852 ( .A1(n15154), .A2(n10261), .ZN(n10414) );
  INV_X1 U12853 ( .A(n12771), .ZN(n15141) );
  NAND2_X1 U12854 ( .A1(n15154), .A2(n15141), .ZN(n10262) );
  INV_X1 U12855 ( .A(n12885), .ZN(n12806) );
  INV_X1 U12856 ( .A(n10263), .ZN(n10269) );
  NOR3_X1 U12857 ( .A1(n15173), .A2(n12493), .A3(n12349), .ZN(n10265) );
  AOI211_X1 U12858 ( .C1(n15151), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10265), .B(
        n10264), .ZN(n10266) );
  MUX2_X1 U12859 ( .A(n10267), .B(n10266), .S(n15154), .Z(n10268) );
  OAI21_X1 U12860 ( .B1(n12806), .B2(n10269), .A(n10268), .ZN(P3_U3231) );
  OR2_X1 U12861 ( .A1(n11587), .A2(n13831), .ZN(n10272) );
  NAND2_X1 U12862 ( .A1(n10273), .A2(n11791), .ZN(n10276) );
  AOI22_X1 U12863 ( .A1(n6422), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10274), 
        .B2(n11659), .ZN(n10275) );
  NAND2_X1 U12864 ( .A1(n10276), .A2(n10275), .ZN(n14737) );
  XNOR2_X1 U12865 ( .A(n14737), .B(n13830), .ZN(n11884) );
  XNOR2_X1 U12866 ( .A(n10594), .B(n10593), .ZN(n14742) );
  INV_X1 U12867 ( .A(n14737), .ZN(n10278) );
  OAI211_X1 U12868 ( .C1(n10278), .C2(n10277), .A(n14707), .B(n14687), .ZN(
        n14738) );
  OAI22_X1 U12869 ( .A1(n14738), .A2(n14173), .B1(n14101), .B2(n10278), .ZN(
        n10295) );
  INV_X1 U12870 ( .A(n13831), .ZN(n10787) );
  NAND2_X1 U12871 ( .A1(n11587), .A2(n10787), .ZN(n10280) );
  AOI21_X1 U12872 ( .B1(n10281), .B2(n10593), .A(n14570), .ZN(n10282) );
  NAND2_X1 U12873 ( .A1(n10282), .A2(n10554), .ZN(n14740) );
  NAND2_X1 U12874 ( .A1(n13831), .A2(n14572), .ZN(n10291) );
  NAND2_X1 U12875 ( .A1(n11707), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10289) );
  OR2_X1 U12876 ( .A1(n6802), .A2(n15311), .ZN(n10288) );
  INV_X1 U12877 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12878 ( .A1(n10284), .A2(n10283), .ZN(n10285) );
  NAND2_X1 U12879 ( .A1(n10566), .A2(n10285), .ZN(n14681) );
  OR2_X1 U12880 ( .A1(n11818), .A2(n14681), .ZN(n10287) );
  OR2_X1 U12881 ( .A1(n11820), .A2(n9318), .ZN(n10286) );
  NAND4_X1 U12882 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n13829) );
  NAND2_X1 U12883 ( .A1(n13829), .A2(n14575), .ZN(n10290) );
  NAND2_X1 U12884 ( .A1(n10291), .A2(n10290), .ZN(n14736) );
  INV_X1 U12885 ( .A(n14736), .ZN(n10292) );
  OAI211_X1 U12886 ( .C1(n14698), .C2(n11013), .A(n14740), .B(n10292), .ZN(
        n10293) );
  MUX2_X1 U12887 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10293), .S(n14700), .Z(
        n10294) );
  AOI211_X1 U12888 ( .C1(n14712), .C2(n14742), .A(n10295), .B(n10294), .ZN(
        n10296) );
  INV_X1 U12889 ( .A(n10296), .ZN(P1_U3285) );
  INV_X1 U12890 ( .A(n14173), .ZN(n14711) );
  OAI22_X1 U12891 ( .A1(n14101), .A2(n10297), .B1(n10792), .B2(n14698), .ZN(
        n10300) );
  MUX2_X1 U12892 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10298), .S(n14700), .Z(
        n10299) );
  AOI211_X1 U12893 ( .C1(n14711), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10302) );
  INV_X1 U12894 ( .A(n10302), .ZN(P1_U3286) );
  XNOR2_X1 U12895 ( .A(n11976), .B(n9052), .ZN(n10481) );
  INV_X1 U12896 ( .A(n10303), .ZN(n11136) );
  NAND2_X1 U12897 ( .A1(n13144), .A2(n13529), .ZN(n10480) );
  XNOR2_X1 U12898 ( .A(n10481), .B(n10480), .ZN(n10484) );
  INV_X1 U12899 ( .A(n10304), .ZN(n10309) );
  NAND2_X1 U12900 ( .A1(n6413), .A2(n10303), .ZN(n10308) );
  XNOR2_X1 U12901 ( .A(n10304), .B(n10308), .ZN(n10353) );
  NAND2_X1 U12902 ( .A1(n11976), .A2(n10305), .ZN(n10306) );
  NAND2_X1 U12903 ( .A1(n10307), .A2(n10306), .ZN(n10352) );
  AND2_X1 U12904 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  XOR2_X1 U12905 ( .A(n10484), .B(n10485), .Z(n10314) );
  NAND2_X1 U12906 ( .A1(n13143), .A2(n13254), .ZN(n10311) );
  NAND2_X1 U12907 ( .A1(n6413), .A2(n13116), .ZN(n10310) );
  NAND2_X1 U12908 ( .A1(n10311), .A2(n10310), .ZN(n10611) );
  AOI22_X1 U12909 ( .A1(n14782), .A2(n10621), .B1(n14534), .B2(n10611), .ZN(
        n10313) );
  NAND2_X1 U12910 ( .A1(n10349), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10312) );
  OAI211_X1 U12911 ( .C1(n10314), .C2(n14777), .A(n10313), .B(n10312), .ZN(
        P2_U3209) );
  OAI21_X1 U12912 ( .B1(n10316), .B2(n12373), .A(n10315), .ZN(n10693) );
  OAI211_X1 U12913 ( .C1(n10319), .C2(n10318), .A(n10317), .B(n12854), .ZN(
        n10321) );
  AOI22_X1 U12914 ( .A1(n15145), .A2(n12516), .B1(n15143), .B2(n12518), .ZN(
        n10320) );
  NAND2_X1 U12915 ( .A1(n10321), .A2(n10320), .ZN(n10690) );
  AOI21_X1 U12916 ( .B1(n15177), .B2(n10693), .A(n10690), .ZN(n10326) );
  OAI22_X1 U12917 ( .A1(n12933), .A2(n10689), .B1(n15199), .B2(n10322), .ZN(
        n10323) );
  INV_X1 U12918 ( .A(n10323), .ZN(n10324) );
  OAI21_X1 U12919 ( .B1(n10326), .B2(n15196), .A(n10324), .ZN(P3_U3466) );
  AOI22_X1 U12920 ( .A1(n8256), .A2(n10434), .B1(n15187), .B2(
        P3_REG0_REG_7__SCAN_IN), .ZN(n10325) );
  OAI21_X1 U12921 ( .B1(n10326), .B2(n15187), .A(n10325), .ZN(P3_U3411) );
  INV_X1 U12922 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10882) );
  AOI21_X1 U12923 ( .B1(n10882), .B2(n10329), .A(n10911), .ZN(n10348) );
  NAND2_X1 U12924 ( .A1(n15082), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n10340) );
  OR2_X1 U12925 ( .A1(n12626), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U12926 ( .A1(n12626), .A2(n10882), .ZN(n10330) );
  AND2_X1 U12927 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  NAND2_X1 U12928 ( .A1(n10332), .A2(n14443), .ZN(n10901) );
  INV_X1 U12929 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U12930 ( .A1(n10333), .A2(n10910), .ZN(n10899) );
  AND2_X1 U12931 ( .A1(n10901), .A2(n10899), .ZN(n10337) );
  XNOR2_X1 U12932 ( .A(n10337), .B(n10902), .ZN(n10338) );
  AND2_X1 U12933 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n10999) );
  AOI21_X1 U12934 ( .B1(n15131), .B2(n10338), .A(n10999), .ZN(n10339) );
  NAND2_X1 U12935 ( .A1(n10340), .A2(n10339), .ZN(n10346) );
  INV_X1 U12936 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10846) );
  AOI21_X1 U12937 ( .B1(n10846), .B2(n10343), .A(n10888), .ZN(n10344) );
  NOR2_X1 U12938 ( .A1(n10344), .A2(n15136), .ZN(n10345) );
  AOI211_X1 U12939 ( .C1(n15106), .C2(n10910), .A(n10346), .B(n10345), .ZN(
        n10347) );
  OAI21_X1 U12940 ( .B1(n10348), .B2(n15125), .A(n10347), .ZN(P3_U3191) );
  INV_X1 U12941 ( .A(n10349), .ZN(n10358) );
  NOR2_X1 U12942 ( .A1(n10350), .A2(n13508), .ZN(n10351) );
  AOI21_X1 U12943 ( .B1(n13144), .B2(n13254), .A(n10351), .ZN(n13544) );
  INV_X1 U12944 ( .A(n13544), .ZN(n14982) );
  AOI22_X1 U12945 ( .A1(n14782), .A2(n9053), .B1(n14534), .B2(n14982), .ZN(
        n10357) );
  NOR2_X1 U12946 ( .A1(n10353), .A2(n10352), .ZN(n10354) );
  OAI21_X1 U12947 ( .B1(n10355), .B2(n10354), .A(n14788), .ZN(n10356) );
  OAI211_X1 U12948 ( .C1(n10358), .C2(n13531), .A(n10357), .B(n10356), .ZN(
        P2_U3194) );
  NOR2_X1 U12949 ( .A1(n12997), .A2(SI_22_), .ZN(n10359) );
  AOI21_X1 U12950 ( .B1(n12331), .B2(P3_STATE_REG_SCAN_IN), .A(n10359), .ZN(
        n10360) );
  OAI21_X1 U12951 ( .B1(n10361), .B2(n14451), .A(n10360), .ZN(n10362) );
  INV_X1 U12952 ( .A(n10362), .ZN(P3_U3273) );
  NAND2_X1 U12953 ( .A1(n14979), .A2(n10363), .ZN(n10364) );
  OR2_X1 U12954 ( .A1(n10365), .A2(n10364), .ZN(n10367) );
  OAI21_X2 U12955 ( .B1(n10367), .B2(n10366), .A(n14938), .ZN(n13543) );
  NOR2_X1 U12956 ( .A1(n8354), .A2(n10369), .ZN(n14931) );
  NAND2_X1 U12957 ( .A1(n14941), .A2(n14931), .ZN(n10615) );
  NAND2_X1 U12958 ( .A1(n14941), .A2(n15064), .ZN(n10368) );
  NAND2_X1 U12959 ( .A1(n10615), .A2(n10368), .ZN(n13542) );
  NAND2_X1 U12960 ( .A1(n14941), .A2(n10370), .ZN(n13533) );
  OAI22_X1 U12961 ( .A1(n13500), .A2(n10371), .B1(n10385), .B2(n13533), .ZN(
        n10376) );
  INV_X1 U12962 ( .A(n14938), .ZN(n13493) );
  AOI21_X1 U12963 ( .B1(n13493), .B2(n8409), .A(n14774), .ZN(n10372) );
  NAND2_X1 U12964 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  INV_X2 U12965 ( .A(n13543), .ZN(n14943) );
  MUX2_X1 U12966 ( .A(n10374), .B(P2_REG2_REG_3__SCAN_IN), .S(n14943), .Z(
        n10375) );
  AOI211_X1 U12967 ( .C1(n10377), .C2(n13542), .A(n10376), .B(n10375), .ZN(
        n10378) );
  INV_X1 U12968 ( .A(n10378), .ZN(P2_U3262) );
  INV_X1 U12969 ( .A(n10379), .ZN(n12306) );
  INV_X1 U12970 ( .A(n12281), .ZN(n12226) );
  NAND2_X1 U12971 ( .A1(n12226), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10800) );
  NAND2_X1 U12972 ( .A1(n10800), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U12973 ( .A1(n12282), .A2(n6689), .B1(n12287), .B2(n10380), .ZN(
        n10381) );
  OAI211_X1 U12974 ( .C1(n12306), .C2(n12289), .A(n10382), .B(n10381), .ZN(
        P3_U3172) );
  INV_X1 U12975 ( .A(n11680), .ZN(n10685) );
  OAI222_X1 U12976 ( .A1(n11860), .A2(P1_U3086), .B1(n11530), .B2(n10685), 
        .C1(n11681), .C2(n6421), .ZN(P1_U3335) );
  NAND2_X1 U12977 ( .A1(n10384), .A2(n10383), .ZN(n10387) );
  INV_X1 U12978 ( .A(n13143), .ZN(n10489) );
  NAND2_X1 U12979 ( .A1(n10489), .A2(n10385), .ZN(n10386) );
  INV_X1 U12980 ( .A(n13142), .ZN(n10391) );
  NAND2_X1 U12981 ( .A1(n10391), .A2(n14995), .ZN(n10388) );
  XNOR2_X1 U12982 ( .A(n10441), .B(n10395), .ZN(n15005) );
  INV_X1 U12983 ( .A(n15005), .ZN(n10408) );
  NAND2_X1 U12984 ( .A1(n10489), .A2(n14783), .ZN(n10543) );
  INV_X1 U12985 ( .A(n10544), .ZN(n10389) );
  NAND2_X1 U12986 ( .A1(n10390), .A2(n10389), .ZN(n10393) );
  NAND2_X1 U12987 ( .A1(n10391), .A2(n10541), .ZN(n10394) );
  INV_X1 U12988 ( .A(n10395), .ZN(n10392) );
  NAND3_X1 U12989 ( .A1(n10393), .A2(n10395), .A3(n10394), .ZN(n10396) );
  NAND2_X1 U12990 ( .A1(n10725), .A2(n10396), .ZN(n10397) );
  NAND2_X1 U12991 ( .A1(n10397), .A2(n15026), .ZN(n10400) );
  NAND2_X1 U12992 ( .A1(n13140), .A2(n13254), .ZN(n10399) );
  NAND2_X1 U12993 ( .A1(n13142), .A2(n13116), .ZN(n10398) );
  AND2_X1 U12994 ( .A1(n10399), .A2(n10398), .ZN(n11989) );
  NAND2_X1 U12995 ( .A1(n10400), .A2(n11989), .ZN(n10401) );
  AOI21_X1 U12996 ( .B1(n15005), .B2(n15064), .A(n10401), .ZN(n15007) );
  MUX2_X1 U12997 ( .A(n10402), .B(n15007), .S(n14941), .Z(n10407) );
  NAND2_X1 U12998 ( .A1(n10537), .A2(n15001), .ZN(n10403) );
  NAND2_X1 U12999 ( .A1(n10403), .A2(n13496), .ZN(n10404) );
  NOR2_X1 U13000 ( .A1(n10717), .A2(n10404), .ZN(n15003) );
  OAI22_X1 U13001 ( .A1(n13533), .A2(n7032), .B1(n14938), .B2(n11987), .ZN(
        n10405) );
  AOI21_X1 U13002 ( .B1(n13535), .B2(n15003), .A(n10405), .ZN(n10406) );
  OAI211_X1 U13003 ( .C1(n10408), .C2(n10615), .A(n10407), .B(n10406), .ZN(
        P2_U3260) );
  XNOR2_X1 U13004 ( .A(n10409), .B(n8225), .ZN(n10413) );
  AOI22_X1 U13005 ( .A1(n15145), .A2(n12520), .B1(n15143), .B2(n15144), .ZN(
        n10412) );
  OAI211_X1 U13006 ( .C1(n7558), .C2(n8225), .A(n12854), .B(n10410), .ZN(
        n10411) );
  OAI211_X1 U13007 ( .C1(n10413), .C2(n12771), .A(n10412), .B(n10411), .ZN(
        n15162) );
  INV_X1 U13008 ( .A(n15162), .ZN(n10418) );
  INV_X1 U13009 ( .A(n10413), .ZN(n15165) );
  INV_X1 U13010 ( .A(n10414), .ZN(n15152) );
  NOR2_X1 U13011 ( .A1(n15154), .A2(n9810), .ZN(n10416) );
  OAI22_X1 U13012 ( .A1(n12883), .A2(n15161), .B1(n11405), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n10415) );
  AOI211_X1 U13013 ( .C1(n15165), .C2(n15152), .A(n10416), .B(n10415), .ZN(
        n10417) );
  OAI21_X1 U13014 ( .B1(n15156), .B2(n10418), .A(n10417), .ZN(P3_U3230) );
  OAI21_X1 U13015 ( .B1(n10420), .B2(n12305), .A(n10419), .ZN(n15176) );
  INV_X1 U13016 ( .A(n10478), .ZN(n10421) );
  OAI22_X1 U13017 ( .A1(n12883), .A2(n15172), .B1(n11405), .B2(n10421), .ZN(
        n10428) );
  OAI211_X1 U13018 ( .C1(n10424), .C2(n10423), .A(n10422), .B(n12854), .ZN(
        n10426) );
  AOI22_X1 U13019 ( .A1(n15145), .A2(n12517), .B1(n15143), .B2(n12519), .ZN(
        n10425) );
  NAND2_X1 U13020 ( .A1(n10426), .A2(n10425), .ZN(n15174) );
  MUX2_X1 U13021 ( .A(n15174), .B(P3_REG2_REG_6__SCAN_IN), .S(n15156), .Z(
        n10427) );
  AOI211_X1 U13022 ( .C1(n12885), .C2(n15176), .A(n10428), .B(n10427), .ZN(
        n10429) );
  INV_X1 U13023 ( .A(n10429), .ZN(P3_U3227) );
  OAI211_X1 U13024 ( .C1(n10432), .C2(n10431), .A(n10430), .B(n12272), .ZN(
        n10440) );
  AOI21_X1 U13025 ( .B1(n12282), .B2(n12516), .A(n10433), .ZN(n10436) );
  NAND2_X1 U13026 ( .A1(n12287), .A2(n10434), .ZN(n10435) );
  OAI211_X1 U13027 ( .C1(n12285), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        n10438) );
  AOI21_X1 U13028 ( .B1(n10687), .B2(n12281), .A(n10438), .ZN(n10439) );
  NAND2_X1 U13029 ( .A1(n10440), .A2(n10439), .ZN(P3_U3153) );
  NAND2_X1 U13030 ( .A1(n10442), .A2(n7032), .ZN(n10443) );
  OR2_X1 U13031 ( .A1(n10444), .A2(n10722), .ZN(n10715) );
  NAND2_X1 U13032 ( .A1(n13140), .A2(n10720), .ZN(n10445) );
  NAND2_X1 U13033 ( .A1(n10715), .A2(n10445), .ZN(n10448) );
  INV_X1 U13034 ( .A(n10458), .ZN(n10447) );
  INV_X1 U13035 ( .A(n10444), .ZN(n10446) );
  OAI21_X1 U13036 ( .B1(n10448), .B2(n10447), .A(n10742), .ZN(n15023) );
  INV_X1 U13037 ( .A(n10720), .ZN(n15011) );
  INV_X1 U13038 ( .A(n10746), .ZN(n10449) );
  AOI211_X1 U13039 ( .C1(n15020), .C2(n10716), .A(n13529), .B(n10449), .ZN(
        n15018) );
  INV_X1 U13040 ( .A(n10769), .ZN(n10453) );
  NAND2_X1 U13041 ( .A1(n13138), .A2(n13254), .ZN(n10451) );
  NAND2_X1 U13042 ( .A1(n13140), .A2(n13116), .ZN(n10450) );
  NAND2_X1 U13043 ( .A1(n10451), .A2(n10450), .ZN(n15019) );
  MUX2_X1 U13044 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15019), .S(n14941), .Z(
        n10452) );
  AOI21_X1 U13045 ( .B1(n13493), .B2(n10453), .A(n10452), .ZN(n10454) );
  OAI21_X1 U13046 ( .B1(n7033), .B2(n13533), .A(n10454), .ZN(n10455) );
  AOI21_X1 U13047 ( .B1(n15018), .B2(n13535), .A(n10455), .ZN(n10460) );
  INV_X1 U13048 ( .A(n13140), .ZN(n10456) );
  NAND2_X1 U13049 ( .A1(n10456), .A2(n10720), .ZN(n10457) );
  NAND2_X1 U13050 ( .A1(n10727), .A2(n10457), .ZN(n10735) );
  XNOR2_X1 U13051 ( .A(n10735), .B(n10458), .ZN(n15025) );
  NAND2_X1 U13052 ( .A1(n13543), .A2(n15026), .ZN(n13473) );
  INV_X1 U13053 ( .A(n13473), .ZN(n13541) );
  NAND2_X1 U13054 ( .A1(n15025), .A2(n13541), .ZN(n10459) );
  OAI211_X1 U13055 ( .C1(n15023), .C2(n13524), .A(n10460), .B(n10459), .ZN(
        P2_U3258) );
  INV_X1 U13056 ( .A(n10461), .ZN(n10466) );
  AOI22_X1 U13057 ( .A1(n12741), .A2(n10638), .B1(n15151), .B2(n10643), .ZN(
        n10462) );
  OAI21_X1 U13058 ( .B1(n9798), .B2(n15154), .A(n10462), .ZN(n10463) );
  AOI21_X1 U13059 ( .B1(n12885), .B2(n10464), .A(n10463), .ZN(n10465) );
  OAI21_X1 U13060 ( .B1(n10466), .B2(n15156), .A(n10465), .ZN(P3_U3228) );
  AOI21_X1 U13061 ( .B1(n12282), .B2(n12517), .A(n10467), .ZN(n10470) );
  NAND2_X1 U13062 ( .A1(n12287), .A2(n10468), .ZN(n10469) );
  OAI211_X1 U13063 ( .C1(n12285), .C2(n10471), .A(n10470), .B(n10469), .ZN(
        n10477) );
  INV_X1 U13064 ( .A(n10473), .ZN(n10474) );
  AOI211_X1 U13065 ( .C1(n10475), .C2(n10472), .A(n12289), .B(n10474), .ZN(
        n10476) );
  AOI211_X1 U13066 ( .C1(n10478), .C2(n12281), .A(n10477), .B(n10476), .ZN(
        n10479) );
  INV_X1 U13067 ( .A(n10479), .ZN(P3_U3179) );
  INV_X1 U13068 ( .A(n10480), .ZN(n10483) );
  INV_X1 U13069 ( .A(n10481), .ZN(n10482) );
  XNOR2_X1 U13070 ( .A(n14783), .B(n11976), .ZN(n10487) );
  AND2_X1 U13071 ( .A1(n13143), .A2(n13529), .ZN(n10486) );
  NAND2_X1 U13072 ( .A1(n10487), .A2(n10486), .ZN(n10491) );
  OAI21_X1 U13073 ( .B1(n10487), .B2(n10486), .A(n10491), .ZN(n14778) );
  INV_X1 U13074 ( .A(n10487), .ZN(n10488) );
  NOR3_X1 U13075 ( .A1(n13110), .A2(n10489), .A3(n10488), .ZN(n10490) );
  AOI21_X1 U13076 ( .B1(n14776), .B2(n14788), .A(n10490), .ZN(n10502) );
  XNOR2_X1 U13077 ( .A(n11976), .B(n14995), .ZN(n10700) );
  NAND2_X1 U13078 ( .A1(n13142), .A2(n13529), .ZN(n10701) );
  XNOR2_X1 U13079 ( .A(n10700), .B(n10701), .ZN(n10492) );
  INV_X1 U13080 ( .A(n10492), .ZN(n10501) );
  INV_X1 U13081 ( .A(n10491), .ZN(n10493) );
  NAND2_X1 U13082 ( .A1(n10494), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14797) );
  NOR2_X1 U13083 ( .A1(n14797), .A2(n10539), .ZN(n10499) );
  INV_X1 U13084 ( .A(n14534), .ZN(n14787) );
  NAND2_X1 U13085 ( .A1(n13141), .A2(n13254), .ZN(n10496) );
  NAND2_X1 U13086 ( .A1(n13143), .A2(n13116), .ZN(n10495) );
  AND2_X1 U13087 ( .A1(n10496), .A2(n10495), .ZN(n10548) );
  NAND2_X1 U13088 ( .A1(n14782), .A2(n10541), .ZN(n10497) );
  NAND2_X1 U13089 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14811) );
  OAI211_X1 U13090 ( .C1(n14787), .C2(n10548), .A(n10497), .B(n14811), .ZN(
        n10498) );
  AOI211_X1 U13091 ( .C1(n11993), .C2(n14788), .A(n10499), .B(n10498), .ZN(
        n10500) );
  OAI21_X1 U13092 ( .B1(n10502), .B2(n10501), .A(n10500), .ZN(P2_U3202) );
  NAND2_X1 U13093 ( .A1(n12122), .A2(n13833), .ZN(n10507) );
  NAND2_X1 U13094 ( .A1(n12129), .A2(n13743), .ZN(n10506) );
  NAND2_X1 U13095 ( .A1(n10507), .A2(n10506), .ZN(n10508) );
  INV_X2 U13096 ( .A(n12039), .ZN(n12130) );
  XNOR2_X1 U13097 ( .A(n10508), .B(n12130), .ZN(n10511) );
  NAND2_X1 U13098 ( .A1(n12122), .A2(n13743), .ZN(n10509) );
  OAI21_X1 U13099 ( .B1(n10184), .B2(n6845), .A(n10509), .ZN(n10510) );
  NOR2_X1 U13100 ( .A1(n10511), .A2(n10510), .ZN(n13736) );
  NAND2_X1 U13101 ( .A1(n10511), .A2(n10510), .ZN(n13734) );
  NAND2_X1 U13102 ( .A1(n11578), .A2(n12129), .ZN(n10513) );
  NAND2_X1 U13103 ( .A1(n12122), .A2(n13832), .ZN(n10512) );
  NAND2_X1 U13104 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  XNOR2_X1 U13105 ( .A(n10514), .B(n12130), .ZN(n10784) );
  AOI22_X1 U13106 ( .A1(n9562), .A2(n13832), .B1(n11578), .B2(n12122), .ZN(
        n10786) );
  XNOR2_X1 U13107 ( .A(n10784), .B(n10786), .ZN(n10515) );
  OAI211_X1 U13108 ( .C1(n10516), .C2(n10515), .A(n10785), .B(n13810), .ZN(
        n10523) );
  NOR2_X1 U13109 ( .A1(n14568), .A2(n10517), .ZN(n10521) );
  NAND2_X1 U13110 ( .A1(n13794), .A2(n13833), .ZN(n10519) );
  OAI211_X1 U13111 ( .C1(n10787), .C2(n14551), .A(n10519), .B(n10518), .ZN(
        n10520) );
  AOI211_X1 U13112 ( .C1(n11578), .C2(n14564), .A(n10521), .B(n10520), .ZN(
        n10522) );
  NAND2_X1 U13113 ( .A1(n10523), .A2(n10522), .ZN(P1_U3239) );
  OAI211_X1 U13114 ( .C1(n10526), .C2(n10525), .A(n10524), .B(n12272), .ZN(
        n10534) );
  AOI21_X1 U13115 ( .B1(n12282), .B2(n12520), .A(n10527), .ZN(n10530) );
  NAND2_X1 U13116 ( .A1(n12287), .A2(n10528), .ZN(n10529) );
  OAI211_X1 U13117 ( .C1(n12285), .C2(n10802), .A(n10530), .B(n10529), .ZN(
        n10531) );
  AOI21_X1 U13118 ( .B1(n10532), .B2(n12281), .A(n10531), .ZN(n10533) );
  NAND2_X1 U13119 ( .A1(n10534), .A2(n10533), .ZN(P3_U3158) );
  OAI21_X1 U13120 ( .B1(n10536), .B2(n10544), .A(n10535), .ZN(n14998) );
  OAI211_X1 U13121 ( .C1(n10538), .C2(n14995), .A(n13496), .B(n10537), .ZN(
        n14994) );
  INV_X1 U13122 ( .A(n10539), .ZN(n10540) );
  AOI22_X1 U13123 ( .A1(n13518), .A2(n10541), .B1(n10540), .B2(n13493), .ZN(
        n10542) );
  OAI21_X1 U13124 ( .B1(n13500), .B2(n14994), .A(n10542), .ZN(n10551) );
  NAND3_X1 U13125 ( .A1(n10545), .A2(n10544), .A3(n10543), .ZN(n10546) );
  NAND2_X1 U13126 ( .A1(n10393), .A2(n10546), .ZN(n10547) );
  NAND2_X1 U13127 ( .A1(n10547), .A2(n15026), .ZN(n10549) );
  NAND2_X1 U13128 ( .A1(n10549), .A2(n10548), .ZN(n14996) );
  MUX2_X1 U13129 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n14996), .S(n13543), .Z(
        n10550) );
  AOI211_X1 U13130 ( .C1(n13542), .C2(n14998), .A(n10551), .B(n10550), .ZN(
        n10552) );
  INV_X1 U13131 ( .A(n10552), .ZN(P2_U3261) );
  OR2_X1 U13132 ( .A1(n14737), .A2(n10795), .ZN(n10553) );
  NAND2_X1 U13133 ( .A1(n10555), .A2(n11791), .ZN(n10558) );
  AOI22_X1 U13134 ( .A1(n10556), .A2(n11659), .B1(n11660), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n10557) );
  XNOR2_X1 U13135 ( .A(n14688), .B(n13829), .ZN(n14677) );
  INV_X1 U13136 ( .A(n14677), .ZN(n14685) );
  INV_X1 U13137 ( .A(n13829), .ZN(n11119) );
  NAND2_X1 U13138 ( .A1(n14688), .A2(n11119), .ZN(n10559) );
  NAND2_X1 U13139 ( .A1(n10560), .A2(n11791), .ZN(n10563) );
  AOI22_X1 U13140 ( .A1(n10561), .A2(n11659), .B1(n6422), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10562) );
  NAND2_X1 U13141 ( .A1(n11817), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10571) );
  INV_X1 U13142 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10564) );
  OR2_X1 U13143 ( .A1(n11797), .A2(n10564), .ZN(n10570) );
  INV_X1 U13144 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U13145 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13146 ( .A1(n10578), .A2(n10567), .ZN(n14177) );
  OR2_X1 U13147 ( .A1(n11818), .A2(n14177), .ZN(n10569) );
  OR2_X1 U13148 ( .A1(n11820), .A2(n14178), .ZN(n10568) );
  NAND4_X1 U13149 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n13828) );
  INV_X1 U13150 ( .A(n13828), .ZN(n11258) );
  OR2_X1 U13151 ( .A1(n14756), .A2(n11258), .ZN(n10572) );
  NAND2_X1 U13152 ( .A1(n10573), .A2(n11791), .ZN(n10576) );
  AOI22_X1 U13153 ( .A1(n10574), .A2(n11659), .B1(n11660), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U13154 ( .A1(n11707), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10583) );
  OR2_X1 U13155 ( .A1(n6802), .A2(n14618), .ZN(n10582) );
  INV_X1 U13156 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10577) );
  AND2_X1 U13157 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  OR2_X1 U13158 ( .A1(n10579), .A2(n10585), .ZN(n11445) );
  OR2_X1 U13159 ( .A1(n11818), .A2(n11445), .ZN(n10581) );
  OR2_X1 U13160 ( .A1(n11820), .A2(n9384), .ZN(n10580) );
  NAND4_X1 U13161 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(
        n13827) );
  OR2_X1 U13162 ( .A1(n11609), .A2(n13827), .ZN(n10964) );
  NAND2_X1 U13163 ( .A1(n11609), .A2(n13827), .ZN(n10967) );
  AND2_X1 U13164 ( .A1(n10964), .A2(n10967), .ZN(n11887) );
  XNOR2_X1 U13165 ( .A(n10976), .B(n11887), .ZN(n10584) );
  NAND2_X1 U13166 ( .A1(n10584), .A2(n14751), .ZN(n10592) );
  NAND2_X1 U13167 ( .A1(n11707), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10590) );
  OR2_X1 U13168 ( .A1(n6802), .A2(n9700), .ZN(n10589) );
  NAND2_X1 U13169 ( .A1(n10585), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10969) );
  OR2_X1 U13170 ( .A1(n10585), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13171 ( .A1(n10969), .A2(n10586), .ZN(n11485) );
  OR2_X1 U13172 ( .A1(n11818), .A2(n11485), .ZN(n10588) );
  OR2_X1 U13173 ( .A1(n11820), .A2(n9505), .ZN(n10587) );
  NAND4_X1 U13174 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n13826) );
  AOI22_X1 U13175 ( .A1(n14572), .A2(n13828), .B1(n13826), .B2(n14575), .ZN(
        n10591) );
  NAND2_X1 U13176 ( .A1(n10592), .A2(n10591), .ZN(n14615) );
  INV_X1 U13177 ( .A(n14615), .ZN(n10603) );
  OR2_X1 U13178 ( .A1(n14688), .A2(n13829), .ZN(n10595) );
  OR2_X1 U13179 ( .A1(n14756), .A2(n13828), .ZN(n10596) );
  XNOR2_X1 U13180 ( .A(n10966), .B(n11887), .ZN(n14617) );
  INV_X1 U13181 ( .A(n11609), .ZN(n14614) );
  INV_X1 U13182 ( .A(n14183), .ZN(n10598) );
  INV_X1 U13183 ( .A(n10982), .ZN(n10984) );
  OAI211_X1 U13184 ( .C1(n14614), .C2(n10598), .A(n10984), .B(n14707), .ZN(
        n14613) );
  OAI22_X1 U13185 ( .A1(n14700), .A2(n9384), .B1(n11445), .B2(n14698), .ZN(
        n10599) );
  AOI21_X1 U13186 ( .B1(n11609), .B2(n14702), .A(n10599), .ZN(n10600) );
  OAI21_X1 U13187 ( .B1(n14613), .B2(n14173), .A(n10600), .ZN(n10601) );
  AOI21_X1 U13188 ( .B1(n14617), .B2(n14712), .A(n10601), .ZN(n10602) );
  OAI21_X1 U13189 ( .B1(n10603), .B2(n14684), .A(n10602), .ZN(P1_U3282) );
  OR2_X1 U13190 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  NAND2_X1 U13191 ( .A1(n10607), .A2(n10606), .ZN(n14991) );
  NAND2_X1 U13192 ( .A1(n14991), .A2(n15064), .ZN(n10614) );
  OAI21_X1 U13193 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(n10612) );
  AOI21_X1 U13194 ( .B1(n10612), .B2(n15026), .A(n10611), .ZN(n10613) );
  AND2_X1 U13195 ( .A1(n10614), .A2(n10613), .ZN(n14993) );
  INV_X1 U13196 ( .A(n10615), .ZN(n10624) );
  INV_X1 U13197 ( .A(n10616), .ZN(n10618) );
  AOI21_X1 U13198 ( .B1(n13527), .B2(n10621), .A(n13529), .ZN(n10617) );
  NAND2_X1 U13199 ( .A1(n10618), .A2(n10617), .ZN(n14989) );
  OAI22_X1 U13200 ( .A1(n13543), .A2(n9331), .B1(n10619), .B2(n14938), .ZN(
        n10620) );
  AOI21_X1 U13201 ( .B1(n13518), .B2(n10621), .A(n10620), .ZN(n10622) );
  OAI21_X1 U13202 ( .B1(n13500), .B2(n14989), .A(n10622), .ZN(n10623) );
  AOI21_X1 U13203 ( .B1(n10624), .B2(n14991), .A(n10623), .ZN(n10625) );
  OAI21_X1 U13204 ( .B1(n14943), .B2(n14993), .A(n10625), .ZN(P2_U3263) );
  AOI21_X1 U13205 ( .B1(n10627), .B2(n10626), .A(n6603), .ZN(n10634) );
  AOI21_X1 U13206 ( .B1(n12282), .B2(n12519), .A(n10628), .ZN(n10630) );
  NAND2_X1 U13207 ( .A1(n12287), .A2(n15167), .ZN(n10629) );
  OAI211_X1 U13208 ( .C1(n12285), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10632) );
  AOI21_X1 U13209 ( .B1(n10860), .B2(n12281), .A(n10632), .ZN(n10633) );
  OAI21_X1 U13210 ( .B1(n10634), .B2(n12289), .A(n10633), .ZN(P3_U3170) );
  XOR2_X1 U13211 ( .A(n10635), .B(n10636), .Z(n10645) );
  AOI21_X1 U13212 ( .B1(n12282), .B2(n12518), .A(n10637), .ZN(n10640) );
  NAND2_X1 U13213 ( .A1(n12287), .A2(n10638), .ZN(n10639) );
  OAI211_X1 U13214 ( .C1(n12285), .C2(n10641), .A(n10640), .B(n10639), .ZN(
        n10642) );
  AOI21_X1 U13215 ( .B1(n10643), .B2(n12281), .A(n10642), .ZN(n10644) );
  OAI21_X1 U13216 ( .B1(n10645), .B2(n12289), .A(n10644), .ZN(P3_U3167) );
  XOR2_X1 U13217 ( .A(n10647), .B(n10646), .Z(n10653) );
  AOI22_X1 U13218 ( .A1(n12282), .A2(n10856), .B1(n12287), .B2(n10648), .ZN(
        n10649) );
  OAI21_X1 U13219 ( .B1(n10650), .B2(n12285), .A(n10649), .ZN(n10651) );
  AOI21_X1 U13220 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10800), .A(n10651), .ZN(
        n10652) );
  OAI21_X1 U13221 ( .B1(n10653), .B2(n12289), .A(n10652), .ZN(P3_U3177) );
  INV_X1 U13222 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10654) );
  MUX2_X1 U13223 ( .A(n10654), .B(P1_REG2_REG_17__SCAN_IN), .S(n11644), .Z(
        n10655) );
  INV_X1 U13224 ( .A(n10655), .ZN(n10663) );
  INV_X1 U13225 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10661) );
  MUX2_X1 U13226 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n10661), .S(n13912), .Z(
        n13915) );
  INV_X1 U13227 ( .A(n11339), .ZN(n14665) );
  INV_X1 U13228 ( .A(n10656), .ZN(n10657) );
  OAI21_X1 U13229 ( .B1(n9693), .B2(n10658), .A(n10657), .ZN(n10659) );
  NOR2_X1 U13230 ( .A1(n14665), .A2(n10659), .ZN(n10660) );
  XNOR2_X1 U13231 ( .A(n10659), .B(n14665), .ZN(n14662) );
  NOR2_X1 U13232 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14662), .ZN(n14661) );
  NOR2_X1 U13233 ( .A1(n10660), .A2(n14661), .ZN(n13916) );
  NAND2_X1 U13234 ( .A1(n13915), .A2(n13916), .ZN(n13913) );
  OAI21_X1 U13235 ( .B1(n10667), .B2(n10661), .A(n13913), .ZN(n10662) );
  NAND2_X1 U13236 ( .A1(n10663), .A2(n10662), .ZN(n11020) );
  OAI211_X1 U13237 ( .C1(n10663), .C2(n10662), .A(n13914), .B(n11020), .ZN(
        n10673) );
  NAND2_X1 U13238 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13754)
         );
  INV_X1 U13239 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14603) );
  MUX2_X1 U13240 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14603), .S(n13912), .Z(
        n13909) );
  OR2_X1 U13241 ( .A1(n11147), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U13242 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  XNOR2_X1 U13243 ( .A(n10666), .B(n11339), .ZN(n14660) );
  NOR2_X1 U13244 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14660), .ZN(n14659) );
  AOI21_X1 U13245 ( .B1(n10666), .B2(n11339), .A(n14659), .ZN(n13910) );
  NAND2_X1 U13246 ( .A1(n13909), .A2(n13910), .ZN(n13907) );
  OAI21_X1 U13247 ( .B1(n14603), .B2(n10667), .A(n13907), .ZN(n10669) );
  INV_X1 U13248 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11390) );
  MUX2_X1 U13249 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n11390), .S(n11644), .Z(
        n10668) );
  NAND2_X1 U13250 ( .A1(n10668), .A2(n10669), .ZN(n11023) );
  OAI211_X1 U13251 ( .C1(n10669), .C2(n10668), .A(n11023), .B(n13908), .ZN(
        n10670) );
  NAND2_X1 U13252 ( .A1(n13754), .A2(n10670), .ZN(n10671) );
  AOI21_X1 U13253 ( .B1(n14655), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10671), 
        .ZN(n10672) );
  OAI211_X1 U13254 ( .C1(n13849), .C2(n11024), .A(n10673), .B(n10672), .ZN(
        P1_U3260) );
  INV_X1 U13255 ( .A(n11695), .ZN(n10675) );
  OAI222_X1 U13256 ( .A1(n11238), .A2(n15225), .B1(n13688), .B2(n10675), .C1(
        n10674), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13257 ( .A1(P1_U3086), .A2(n11870), .B1(n11530), .B2(n10675), 
        .C1(n11696), .C2(n6421), .ZN(P1_U3334) );
  OAI21_X1 U13258 ( .B1(n10677), .B2(n10676), .A(n12272), .ZN(n10684) );
  AOI21_X1 U13259 ( .B1(n12282), .B2(n12515), .A(n10678), .ZN(n10680) );
  NAND2_X1 U13260 ( .A1(n12287), .A2(n12384), .ZN(n10679) );
  OAI211_X1 U13261 ( .C1(n12285), .C2(n10758), .A(n10680), .B(n10679), .ZN(
        n10681) );
  AOI21_X1 U13262 ( .B1(n10761), .B2(n12281), .A(n10681), .ZN(n10682) );
  OAI21_X1 U13263 ( .B1(n10684), .B2(n10683), .A(n10682), .ZN(P3_U3161) );
  OAI222_X1 U13264 ( .A1(n11238), .A2(n10686), .B1(P2_U3088), .B2(n8951), .C1(
        n13688), .C2(n10685), .ZN(P2_U3307) );
  INV_X1 U13265 ( .A(n10687), .ZN(n10688) );
  OAI22_X1 U13266 ( .A1(n12883), .A2(n10689), .B1(n11405), .B2(n10688), .ZN(
        n10692) );
  MUX2_X1 U13267 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n10690), .S(n15154), .Z(
        n10691) );
  AOI211_X1 U13268 ( .C1(n12885), .C2(n10693), .A(n10692), .B(n10691), .ZN(
        n10694) );
  INV_X1 U13269 ( .A(n10694), .ZN(P3_U3226) );
  NAND2_X1 U13270 ( .A1(n13139), .A2(n13254), .ZN(n10696) );
  NAND2_X1 U13271 ( .A1(n13141), .A2(n13116), .ZN(n10695) );
  AND2_X1 U13272 ( .A1(n10696), .A2(n10695), .ZN(n10729) );
  INV_X1 U13273 ( .A(n10729), .ZN(n10697) );
  AOI22_X1 U13274 ( .A1(n14534), .A2(n10697), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10698) );
  OAI21_X1 U13275 ( .B1(n14797), .B2(n10718), .A(n10698), .ZN(n10709) );
  XNOR2_X1 U13276 ( .A(n10720), .B(n11976), .ZN(n10770) );
  AND2_X1 U13277 ( .A1(n13140), .A2(n13529), .ZN(n10699) );
  NAND2_X1 U13278 ( .A1(n10770), .A2(n10699), .ZN(n10775) );
  OAI21_X1 U13279 ( .B1(n10770), .B2(n10699), .A(n10775), .ZN(n10707) );
  NAND2_X1 U13280 ( .A1(n13141), .A2(n13529), .ZN(n10703) );
  INV_X1 U13281 ( .A(n10703), .ZN(n10705) );
  XNOR2_X1 U13282 ( .A(n11976), .B(n15001), .ZN(n10704) );
  INV_X1 U13283 ( .A(n10700), .ZN(n11990) );
  INV_X1 U13284 ( .A(n10701), .ZN(n10702) );
  XNOR2_X1 U13285 ( .A(n10704), .B(n10703), .ZN(n11991) );
  NOR2_X2 U13286 ( .A1(n10706), .A2(n10707), .ZN(n10778) );
  AOI211_X1 U13287 ( .C1(n10707), .C2(n10706), .A(n14777), .B(n10778), .ZN(
        n10708) );
  AOI211_X1 U13288 ( .C1(n10720), .C2(n14782), .A(n10709), .B(n10708), .ZN(
        n10710) );
  INV_X1 U13289 ( .A(n10710), .ZN(P2_U3211) );
  NAND2_X1 U13290 ( .A1(n10711), .A2(n14446), .ZN(n10712) );
  OAI211_X1 U13291 ( .C1(n10713), .C2(n12997), .A(n10712), .B(n12506), .ZN(
        P3_U3272) );
  NAND2_X1 U13292 ( .A1(n10444), .A2(n10722), .ZN(n10714) );
  AND2_X1 U13293 ( .A1(n10715), .A2(n10714), .ZN(n15014) );
  OAI211_X1 U13294 ( .C1(n10717), .C2(n15011), .A(n13496), .B(n10716), .ZN(
        n15010) );
  INV_X1 U13295 ( .A(n10718), .ZN(n10719) );
  AOI22_X1 U13296 ( .A1(n13518), .A2(n10720), .B1(n13493), .B2(n10719), .ZN(
        n10721) );
  OAI21_X1 U13297 ( .B1(n13500), .B2(n15010), .A(n10721), .ZN(n10732) );
  INV_X1 U13298 ( .A(n10722), .ZN(n10724) );
  NAND3_X1 U13299 ( .A1(n10725), .A2(n10724), .A3(n10723), .ZN(n10726) );
  NAND2_X1 U13300 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  NAND2_X1 U13301 ( .A1(n10728), .A2(n15026), .ZN(n10730) );
  NAND2_X1 U13302 ( .A1(n10730), .A2(n10729), .ZN(n15009) );
  MUX2_X1 U13303 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n15009), .S(n14941), .Z(
        n10731) );
  AOI211_X1 U13304 ( .C1(n15014), .C2(n13542), .A(n10732), .B(n10731), .ZN(
        n10733) );
  INV_X1 U13305 ( .A(n10733), .ZN(P2_U3259) );
  INV_X1 U13306 ( .A(n13139), .ZN(n10865) );
  OR2_X1 U13307 ( .A1(n10865), .A2(n15020), .ZN(n10734) );
  NAND2_X1 U13308 ( .A1(n10735), .A2(n10734), .ZN(n10737) );
  NAND2_X1 U13309 ( .A1(n15020), .A2(n10865), .ZN(n10736) );
  NAND2_X1 U13310 ( .A1(n10737), .A2(n10736), .ZN(n10922) );
  XNOR2_X1 U13311 ( .A(n10922), .B(n10921), .ZN(n10740) );
  NAND2_X1 U13312 ( .A1(n13137), .A2(n13254), .ZN(n10739) );
  NAND2_X1 U13313 ( .A1(n13139), .A2(n13116), .ZN(n10738) );
  NAND2_X1 U13314 ( .A1(n10739), .A2(n10738), .ZN(n10868) );
  AOI21_X1 U13315 ( .B1(n10740), .B2(n15026), .A(n10868), .ZN(n15033) );
  NAND2_X1 U13316 ( .A1(n15020), .A2(n13139), .ZN(n10741) );
  INV_X1 U13317 ( .A(n10921), .ZN(n10743) );
  OR2_X1 U13318 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  NAND2_X1 U13319 ( .A1(n10930), .A2(n10745), .ZN(n15028) );
  INV_X1 U13320 ( .A(n15028), .ZN(n10752) );
  AOI21_X1 U13321 ( .B1(n10746), .B2(n15029), .A(n13529), .ZN(n10747) );
  NAND2_X1 U13322 ( .A1(n10747), .A2(n10935), .ZN(n15031) );
  OAI22_X1 U13323 ( .A1(n13543), .A2(n10748), .B1(n10870), .B2(n14938), .ZN(
        n10749) );
  AOI21_X1 U13324 ( .B1(n13518), .B2(n15029), .A(n10749), .ZN(n10750) );
  OAI21_X1 U13325 ( .B1(n15031), .B2(n13500), .A(n10750), .ZN(n10751) );
  AOI21_X1 U13326 ( .B1(n10752), .B2(n13542), .A(n10751), .ZN(n10753) );
  OAI21_X1 U13327 ( .B1(n14943), .B2(n15033), .A(n10753), .ZN(P2_U3257) );
  INV_X1 U13328 ( .A(n10754), .ZN(n10755) );
  AOI21_X1 U13329 ( .B1(n12378), .B2(n10756), .A(n10755), .ZN(n10757) );
  OAI222_X1 U13330 ( .A1(n12873), .A2(n11205), .B1(n12875), .B2(n10758), .C1(
        n15149), .C2(n10757), .ZN(n10831) );
  INV_X1 U13331 ( .A(n10831), .ZN(n10766) );
  OAI21_X1 U13332 ( .B1(n10760), .B2(n12378), .A(n10759), .ZN(n10832) );
  AOI22_X1 U13333 ( .A1(n12741), .A2(n12384), .B1(n15151), .B2(n10761), .ZN(
        n10762) );
  OAI21_X1 U13334 ( .B1(n10763), .B2(n15154), .A(n10762), .ZN(n10764) );
  AOI21_X1 U13335 ( .B1(n10832), .B2(n12885), .A(n10764), .ZN(n10765) );
  OAI21_X1 U13336 ( .B1(n10766), .B2(n15156), .A(n10765), .ZN(P3_U3225) );
  NAND2_X1 U13337 ( .A1(n14534), .A2(n15019), .ZN(n10767) );
  OAI211_X1 U13338 ( .C1(n14797), .C2(n10769), .A(n10768), .B(n10767), .ZN(
        n10782) );
  NAND3_X1 U13339 ( .A1(n13096), .A2(n13140), .A3(n10770), .ZN(n10780) );
  XNOR2_X1 U13340 ( .A(n15020), .B(n11976), .ZN(n10771) );
  AND2_X1 U13341 ( .A1(n13139), .A2(n13529), .ZN(n10772) );
  NAND2_X1 U13342 ( .A1(n10771), .A2(n10772), .ZN(n10817) );
  INV_X1 U13343 ( .A(n10771), .ZN(n10864) );
  INV_X1 U13344 ( .A(n10772), .ZN(n10773) );
  NAND2_X1 U13345 ( .A1(n10864), .A2(n10773), .ZN(n10774) );
  AND2_X1 U13346 ( .A1(n10817), .A2(n10774), .ZN(n10776) );
  OAI21_X1 U13347 ( .B1(n10778), .B2(n10776), .A(n14788), .ZN(n10779) );
  INV_X1 U13348 ( .A(n10775), .ZN(n10777) );
  OAI21_X2 U13349 ( .B1(n10778), .B2(n10777), .A(n10776), .ZN(n10818) );
  INV_X1 U13350 ( .A(n10818), .ZN(n10867) );
  AOI21_X1 U13351 ( .B1(n10780), .B2(n10779), .A(n10867), .ZN(n10781) );
  AOI211_X1 U13352 ( .C1(n15020), .C2(n14782), .A(n10782), .B(n10781), .ZN(
        n10783) );
  INV_X1 U13353 ( .A(n10783), .ZN(P2_U3185) );
  NOR2_X1 U13354 ( .A1(n10184), .A2(n10787), .ZN(n10788) );
  AOI21_X1 U13355 ( .B1(n11587), .B2(n12122), .A(n10788), .ZN(n11008) );
  AOI22_X1 U13356 ( .A1(n11587), .A2(n12129), .B1(n12122), .B2(n13831), .ZN(
        n10789) );
  XNOR2_X1 U13357 ( .A(n10789), .B(n12130), .ZN(n11007) );
  XOR2_X1 U13358 ( .A(n11008), .B(n11007), .Z(n10790) );
  OAI211_X1 U13359 ( .C1(n10791), .C2(n10790), .A(n11006), .B(n13810), .ZN(
        n10799) );
  NOR2_X1 U13360 ( .A1(n14568), .A2(n10792), .ZN(n10797) );
  NAND2_X1 U13361 ( .A1(n13794), .A2(n13832), .ZN(n10794) );
  OAI211_X1 U13362 ( .C1(n10795), .C2(n14551), .A(n10794), .B(n10793), .ZN(
        n10796) );
  AOI211_X1 U13363 ( .C1(n11587), .C2(n14564), .A(n10797), .B(n10796), .ZN(
        n10798) );
  NAND2_X1 U13364 ( .A1(n10799), .A2(n10798), .ZN(P1_U3213) );
  INV_X1 U13365 ( .A(n10800), .ZN(n10816) );
  INV_X1 U13366 ( .A(n12285), .ZN(n12224) );
  INV_X1 U13367 ( .A(n12282), .ZN(n12191) );
  OAI22_X1 U13368 ( .A1(n10802), .A2(n12191), .B1(n12278), .B2(n10801), .ZN(
        n10803) );
  AOI21_X1 U13369 ( .B1(n12224), .B2(n15142), .A(n10803), .ZN(n10814) );
  INV_X1 U13370 ( .A(n10804), .ZN(n15138) );
  OAI21_X1 U13371 ( .B1(n15138), .B2(n10806), .A(n10805), .ZN(n10812) );
  NAND3_X1 U13372 ( .A1(n10808), .A2(n10807), .A3(n6689), .ZN(n10809) );
  AOI21_X1 U13373 ( .B1(n10810), .B2(n10809), .A(n15139), .ZN(n10811) );
  OAI21_X1 U13374 ( .B1(n10812), .B2(n10811), .A(n12272), .ZN(n10813) );
  OAI211_X1 U13375 ( .C1(n10816), .C2(n10815), .A(n10814), .B(n10813), .ZN(
        P3_U3162) );
  XNOR2_X1 U13376 ( .A(n15029), .B(n11972), .ZN(n10819) );
  NAND2_X1 U13377 ( .A1(n13138), .A2(n10303), .ZN(n10820) );
  XNOR2_X1 U13378 ( .A(n10819), .B(n10820), .ZN(n10875) );
  INV_X1 U13379 ( .A(n10819), .ZN(n10826) );
  NAND2_X1 U13380 ( .A1(n13137), .A2(n13529), .ZN(n11096) );
  XNOR2_X1 U13381 ( .A(n15038), .B(n11972), .ZN(n11095) );
  XOR2_X1 U13382 ( .A(n11096), .B(n11095), .Z(n10828) );
  NAND2_X1 U13383 ( .A1(n13136), .A2(n13254), .ZN(n10822) );
  NAND2_X1 U13384 ( .A1(n13138), .A2(n13116), .ZN(n10821) );
  AND2_X1 U13385 ( .A1(n10822), .A2(n10821), .ZN(n10927) );
  INV_X1 U13386 ( .A(n10927), .ZN(n10823) );
  AOI22_X1 U13387 ( .A1(n14534), .A2(n10823), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10824) );
  OAI21_X1 U13388 ( .B1(n14797), .B2(n10937), .A(n10824), .ZN(n10825) );
  AOI21_X1 U13389 ( .B1(n15038), .B2(n14794), .A(n10825), .ZN(n10830) );
  OAI22_X1 U13390 ( .A1(n13110), .A2(n10923), .B1(n10826), .B2(n14777), .ZN(
        n10827) );
  NAND3_X1 U13391 ( .A1(n10871), .A2(n10828), .A3(n10827), .ZN(n10829) );
  OAI211_X1 U13392 ( .C1(n6595), .C2(n14777), .A(n10830), .B(n10829), .ZN(
        P2_U3203) );
  AOI21_X1 U13393 ( .B1(n15177), .B2(n10832), .A(n10831), .ZN(n10839) );
  INV_X1 U13394 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n10833) );
  OAI22_X1 U13395 ( .A1(n12383), .A2(n12981), .B1(n15185), .B2(n10833), .ZN(
        n10834) );
  INV_X1 U13396 ( .A(n10834), .ZN(n10835) );
  OAI21_X1 U13397 ( .B1(n10839), .B2(n15187), .A(n10835), .ZN(P3_U3414) );
  INV_X1 U13398 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10836) );
  OAI22_X1 U13399 ( .A1(n12933), .A2(n12383), .B1(n15199), .B2(n10836), .ZN(
        n10837) );
  INV_X1 U13400 ( .A(n10837), .ZN(n10838) );
  OAI21_X1 U13401 ( .B1(n10839), .B2(n15196), .A(n10838), .ZN(P3_U3467) );
  INV_X1 U13402 ( .A(n10842), .ZN(n12388) );
  XNOR2_X1 U13403 ( .A(n10840), .B(n12388), .ZN(n10878) );
  INV_X1 U13404 ( .A(n10878), .ZN(n10851) );
  OAI211_X1 U13405 ( .C1(n10843), .C2(n10842), .A(n10841), .B(n12854), .ZN(
        n10845) );
  AOI22_X1 U13406 ( .A1(n15145), .A2(n12514), .B1(n15143), .B2(n12516), .ZN(
        n10844) );
  NAND2_X1 U13407 ( .A1(n10845), .A2(n10844), .ZN(n10877) );
  NOR2_X1 U13408 ( .A1(n15154), .A2(n10846), .ZN(n10849) );
  INV_X1 U13409 ( .A(n10847), .ZN(n11004) );
  OAI22_X1 U13410 ( .A1(n12883), .A2(n12391), .B1(n11405), .B2(n11004), .ZN(
        n10848) );
  AOI211_X1 U13411 ( .C1(n10877), .C2(n15154), .A(n10849), .B(n10848), .ZN(
        n10850) );
  OAI21_X1 U13412 ( .B1(n12806), .B2(n10851), .A(n10850), .ZN(P3_U3224) );
  OAI21_X1 U13413 ( .B1(n10853), .B2(n12307), .A(n10852), .ZN(n15168) );
  INV_X1 U13414 ( .A(n15168), .ZN(n10863) );
  OAI211_X1 U13415 ( .C1(n10855), .C2(n12356), .A(n10854), .B(n12854), .ZN(
        n10858) );
  AOI22_X1 U13416 ( .A1(n15145), .A2(n12519), .B1(n15143), .B2(n10856), .ZN(
        n10857) );
  AND2_X1 U13417 ( .A1(n10858), .A2(n10857), .ZN(n15169) );
  MUX2_X1 U13418 ( .A(n15169), .B(n10859), .S(n15156), .Z(n10862) );
  AOI22_X1 U13419 ( .A1(n12741), .A2(n15167), .B1(n15151), .B2(n10860), .ZN(
        n10861) );
  OAI211_X1 U13420 ( .C1(n12806), .C2(n10863), .A(n10862), .B(n10861), .ZN(
        P3_U3229) );
  NOR3_X1 U13421 ( .A1(n13110), .A2(n10865), .A3(n10864), .ZN(n10866) );
  AOI21_X1 U13422 ( .B1(n10867), .B2(n14788), .A(n10866), .ZN(n10876) );
  AND2_X1 U13423 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13197) );
  AOI21_X1 U13424 ( .B1(n14534), .B2(n10868), .A(n13197), .ZN(n10869) );
  OAI21_X1 U13425 ( .B1(n14797), .B2(n10870), .A(n10869), .ZN(n10873) );
  NOR2_X1 U13426 ( .A1(n10871), .A2(n14777), .ZN(n10872) );
  AOI211_X1 U13427 ( .C1(n15029), .C2(n14794), .A(n10873), .B(n10872), .ZN(
        n10874) );
  OAI21_X1 U13428 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(P2_U3193) );
  AOI21_X1 U13429 ( .B1(n10878), .B2(n15177), .A(n10877), .ZN(n10885) );
  INV_X1 U13430 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n10879) );
  OAI22_X1 U13431 ( .A1(n12391), .A2(n12981), .B1(n15185), .B2(n10879), .ZN(
        n10880) );
  INV_X1 U13432 ( .A(n10880), .ZN(n10881) );
  OAI21_X1 U13433 ( .B1(n10885), .B2(n15187), .A(n10881), .ZN(P3_U3417) );
  OAI22_X1 U13434 ( .A1(n12933), .A2(n12391), .B1(n15199), .B2(n10882), .ZN(
        n10883) );
  INV_X1 U13435 ( .A(n10883), .ZN(n10884) );
  OAI21_X1 U13436 ( .B1(n10885), .B2(n15196), .A(n10884), .ZN(P3_U3468) );
  INV_X1 U13437 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10894) );
  INV_X1 U13438 ( .A(n14449), .ZN(n11324) );
  NAND2_X1 U13439 ( .A1(n15095), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10892) );
  OR2_X1 U13440 ( .A1(n15095), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10889) );
  NAND2_X1 U13441 ( .A1(n10892), .A2(n10889), .ZN(n15093) );
  AOI21_X1 U13442 ( .B1(n10894), .B2(n10893), .A(n11305), .ZN(n10920) );
  OR2_X1 U13443 ( .A1(n12675), .A2(n10894), .ZN(n10896) );
  NAND2_X1 U13444 ( .A1(n12626), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n10895) );
  NAND2_X1 U13445 ( .A1(n10896), .A2(n10895), .ZN(n11314) );
  XNOR2_X1 U13446 ( .A(n14449), .B(n11314), .ZN(n10905) );
  MUX2_X1 U13447 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12626), .Z(n10897) );
  NOR2_X1 U13448 ( .A1(n10897), .A2(n15095), .ZN(n10903) );
  AOI21_X1 U13449 ( .B1(n15095), .B2(n10897), .A(n10903), .ZN(n10898) );
  INV_X1 U13450 ( .A(n10898), .ZN(n15108) );
  INV_X1 U13451 ( .A(n10899), .ZN(n10900) );
  NOR2_X1 U13452 ( .A1(n15108), .A2(n15109), .ZN(n15107) );
  NOR2_X1 U13453 ( .A1(n10903), .A2(n15107), .ZN(n10904) );
  AOI21_X1 U13454 ( .B1(n10905), .B2(n10904), .A(n11315), .ZN(n10908) );
  NAND2_X1 U13455 ( .A1(n15082), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n10907) );
  AND2_X1 U13456 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11452) );
  INV_X1 U13457 ( .A(n11452), .ZN(n10906) );
  OAI211_X1 U13458 ( .C1(n10908), .C2(n15110), .A(n10907), .B(n10906), .ZN(
        n10918) );
  INV_X1 U13459 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U13460 ( .A1(n10910), .A2(n10909), .ZN(n10912) );
  NAND2_X1 U13461 ( .A1(n15095), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n10914) );
  OR2_X1 U13462 ( .A1(n15095), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n10913) );
  NAND2_X1 U13463 ( .A1(n10914), .A2(n10913), .ZN(n15099) );
  AND2_X2 U13464 ( .A1(n15102), .A2(n10914), .ZN(n11323) );
  AOI21_X1 U13465 ( .B1(n15343), .B2(n10915), .A(n11325), .ZN(n10916) );
  NOR2_X1 U13466 ( .A1(n10916), .A2(n15125), .ZN(n10917) );
  AOI211_X1 U13467 ( .C1(n15106), .C2(n11324), .A(n10918), .B(n10917), .ZN(
        n10919) );
  OAI21_X1 U13468 ( .B1(n10920), .B2(n15136), .A(n10919), .ZN(P3_U3193) );
  NAND2_X1 U13469 ( .A1(n10922), .A2(n10921), .ZN(n10925) );
  NAND2_X1 U13470 ( .A1(n15029), .A2(n10923), .ZN(n10924) );
  INV_X1 U13471 ( .A(n10931), .ZN(n11031) );
  XNOR2_X1 U13472 ( .A(n11032), .B(n11031), .ZN(n10926) );
  NAND2_X1 U13473 ( .A1(n10926), .A2(n15026), .ZN(n10928) );
  NAND2_X1 U13474 ( .A1(n10928), .A2(n10927), .ZN(n15042) );
  INV_X1 U13475 ( .A(n15042), .ZN(n10944) );
  NAND2_X1 U13476 ( .A1(n15029), .A2(n13138), .ZN(n10929) );
  OR2_X1 U13477 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  NAND2_X1 U13478 ( .A1(n11039), .A2(n10933), .ZN(n15037) );
  INV_X1 U13479 ( .A(n15037), .ZN(n10942) );
  NAND2_X1 U13480 ( .A1(n10935), .A2(n15038), .ZN(n10934) );
  NAND2_X1 U13481 ( .A1(n10934), .A2(n13496), .ZN(n10936) );
  OR2_X1 U13482 ( .A1(n10936), .A2(n11043), .ZN(n15039) );
  OAI22_X1 U13483 ( .A1(n13543), .A2(n10938), .B1(n10937), .B2(n14938), .ZN(
        n10939) );
  AOI21_X1 U13484 ( .B1(n13518), .B2(n15038), .A(n10939), .ZN(n10940) );
  OAI21_X1 U13485 ( .B1(n15039), .B2(n13500), .A(n10940), .ZN(n10941) );
  AOI21_X1 U13486 ( .B1(n10942), .B2(n13542), .A(n10941), .ZN(n10943) );
  OAI21_X1 U13487 ( .B1(n14943), .B2(n10944), .A(n10943), .ZN(P2_U3256) );
  INV_X1 U13488 ( .A(n10945), .ZN(n10947) );
  OAI222_X1 U13489 ( .A1(n11238), .A2(n10948), .B1(n13688), .B2(n10947), .C1(
        P2_U3088), .C2(n10946), .ZN(P2_U3305) );
  OAI211_X1 U13490 ( .C1(n10950), .C2(n12310), .A(n10949), .B(n12854), .ZN(
        n10952) );
  AOI22_X1 U13491 ( .A1(n15145), .A2(n11202), .B1(n15143), .B2(n12515), .ZN(
        n10951) );
  NAND2_X1 U13492 ( .A1(n10952), .A2(n10951), .ZN(n15181) );
  INV_X1 U13493 ( .A(n15181), .ZN(n10959) );
  INV_X1 U13494 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10954) );
  INV_X1 U13495 ( .A(n11200), .ZN(n10953) );
  OAI22_X1 U13496 ( .A1(n15154), .A2(n10954), .B1(n10953), .B2(n11405), .ZN(
        n10957) );
  AND2_X1 U13497 ( .A1(n10955), .A2(n12310), .ZN(n15180) );
  NOR3_X1 U13498 ( .A1(n6589), .A2(n15180), .A3(n12806), .ZN(n10956) );
  AOI211_X1 U13499 ( .C1(n12741), .C2(n15183), .A(n10957), .B(n10956), .ZN(
        n10958) );
  OAI21_X1 U13500 ( .B1(n15156), .B2(n10959), .A(n10958), .ZN(P3_U3223) );
  NAND2_X1 U13501 ( .A1(n10960), .A2(n11791), .ZN(n10963) );
  AOI22_X1 U13502 ( .A1(n10961), .A2(n11659), .B1(n6422), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10962) );
  XNOR2_X1 U13503 ( .A(n11613), .B(n13826), .ZN(n11888) );
  INV_X1 U13504 ( .A(n10964), .ZN(n10965) );
  XOR2_X1 U13505 ( .A(n11065), .B(n11888), .Z(n10981) );
  INV_X1 U13506 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13507 ( .A1(n10969), .A2(n10968), .ZN(n10970) );
  NAND2_X1 U13508 ( .A1(n11072), .A2(n10970), .ZN(n14477) );
  OR2_X1 U13509 ( .A1(n14477), .A2(n11818), .ZN(n10974) );
  NAND2_X1 U13510 ( .A1(n11707), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10973) );
  OR2_X1 U13511 ( .A1(n11820), .A2(n9692), .ZN(n10972) );
  OR2_X1 U13512 ( .A1(n6802), .A2(n9704), .ZN(n10971) );
  NAND4_X1 U13513 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n13825) );
  AOI22_X1 U13514 ( .A1(n14575), .A2(n13825), .B1(n13827), .B2(n14572), .ZN(
        n10980) );
  INV_X1 U13515 ( .A(n13827), .ZN(n10977) );
  NOR2_X1 U13516 ( .A1(n11609), .A2(n10977), .ZN(n10975) );
  NAND2_X1 U13517 ( .A1(n10978), .A2(n11888), .ZN(n11057) );
  OAI211_X1 U13518 ( .C1(n10978), .C2(n11888), .A(n11057), .B(n14751), .ZN(
        n10979) );
  OAI211_X1 U13519 ( .C1(n10981), .C2(n14609), .A(n10980), .B(n10979), .ZN(
        n10990) );
  INV_X1 U13520 ( .A(n11613), .ZN(n11491) );
  NAND2_X1 U13521 ( .A1(n11491), .A2(n10982), .ZN(n11150) );
  INV_X1 U13522 ( .A(n11150), .ZN(n10983) );
  AOI211_X1 U13523 ( .C1(n11613), .C2(n10984), .A(n14718), .B(n10983), .ZN(
        n10991) );
  NOR2_X1 U13524 ( .A1(n10990), .A2(n10991), .ZN(n10989) );
  INV_X1 U13525 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10985) );
  OAI22_X1 U13526 ( .A1(n11491), .A2(n14300), .B1(n14764), .B2(n10985), .ZN(
        n10986) );
  INV_X1 U13527 ( .A(n10986), .ZN(n10987) );
  OAI21_X1 U13528 ( .B1(n10989), .B2(n14763), .A(n10987), .ZN(P1_U3495) );
  AOI22_X1 U13529 ( .A1(n11613), .A2(n14263), .B1(n6820), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n10988) );
  OAI21_X1 U13530 ( .B1(n10989), .B2(n6820), .A(n10988), .ZN(P1_U3540) );
  AOI21_X1 U13531 ( .B1(n10991), .B2(n14471), .A(n10990), .ZN(n10994) );
  OAI22_X1 U13532 ( .A1(n14700), .A2(n9505), .B1(n11485), .B2(n14698), .ZN(
        n10992) );
  AOI21_X1 U13533 ( .B1(n11613), .B2(n14702), .A(n10992), .ZN(n10993) );
  OAI21_X1 U13534 ( .B1(n10994), .B2(n14684), .A(n10993), .ZN(P1_U3281) );
  OAI21_X1 U13535 ( .B1(n10997), .B2(n10996), .A(n10995), .ZN(n10998) );
  NAND2_X1 U13536 ( .A1(n10998), .A2(n12272), .ZN(n11003) );
  AOI21_X1 U13537 ( .B1(n12282), .B2(n12514), .A(n10999), .ZN(n11000) );
  OAI21_X1 U13538 ( .B1(n12278), .B2(n12391), .A(n11000), .ZN(n11001) );
  AOI21_X1 U13539 ( .B1(n12224), .B2(n12516), .A(n11001), .ZN(n11002) );
  OAI211_X1 U13540 ( .C1(n11004), .C2(n12226), .A(n11003), .B(n11002), .ZN(
        P3_U3171) );
  AOI22_X1 U13541 ( .A1(n14737), .A2(n12129), .B1(n12122), .B2(n13830), .ZN(
        n11005) );
  XNOR2_X1 U13542 ( .A(n11005), .B(n12130), .ZN(n11114) );
  AOI22_X1 U13543 ( .A1(n14737), .A2(n12122), .B1(n9562), .B2(n13830), .ZN(
        n11115) );
  XNOR2_X1 U13544 ( .A(n11114), .B(n11115), .ZN(n11010) );
  AOI21_X1 U13545 ( .B1(n11010), .B2(n11009), .A(n6592), .ZN(n11016) );
  NAND2_X1 U13546 ( .A1(n13805), .A2(n14736), .ZN(n11011) );
  OAI211_X1 U13547 ( .C1(n14568), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11014) );
  AOI21_X1 U13548 ( .B1(n14737), .B2(n14564), .A(n11014), .ZN(n11015) );
  OAI21_X1 U13549 ( .B1(n11016), .B2(n14559), .A(n11015), .ZN(P1_U3221) );
  INV_X1 U13550 ( .A(n11017), .ZN(n11018) );
  OAI222_X1 U13551 ( .A1(P3_U3151), .A2(n11019), .B1(n14451), .B2(n11018), 
        .C1(n7376), .C2(n12997), .ZN(P3_U3271) );
  NAND2_X1 U13552 ( .A1(n11644), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U13553 ( .A1(n11021), .A2(n11020), .ZN(n11212) );
  XOR2_X1 U13554 ( .A(n11632), .B(n11212), .Z(n11022) );
  NAND2_X1 U13555 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11022), .ZN(n11214) );
  OAI211_X1 U13556 ( .C1(n11022), .C2(P1_REG2_REG_18__SCAN_IN), .A(n13914), 
        .B(n11214), .ZN(n11029) );
  NAND2_X1 U13557 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13795)
         );
  OAI21_X1 U13558 ( .B1(n11390), .B2(n11024), .A(n11023), .ZN(n11216) );
  XNOR2_X1 U13559 ( .A(n11216), .B(n11030), .ZN(n11025) );
  NAND2_X1 U13560 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11025), .ZN(n11218) );
  OAI211_X1 U13561 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11025), .A(n13908), 
        .B(n11218), .ZN(n11026) );
  NAND2_X1 U13562 ( .A1(n13795), .A2(n11026), .ZN(n11027) );
  AOI21_X1 U13563 ( .B1(n14655), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11027), 
        .ZN(n11028) );
  OAI211_X1 U13564 ( .C1(n13849), .C2(n11030), .A(n11029), .B(n11028), .ZN(
        P1_U3261) );
  NAND2_X1 U13565 ( .A1(n15038), .A2(n11033), .ZN(n11034) );
  INV_X1 U13566 ( .A(n11040), .ZN(n11170) );
  XNOR2_X1 U13567 ( .A(n11171), .B(n11170), .ZN(n11035) );
  NAND2_X1 U13568 ( .A1(n11035), .A2(n15026), .ZN(n11038) );
  NAND2_X1 U13569 ( .A1(n13135), .A2(n13254), .ZN(n11037) );
  NAND2_X1 U13570 ( .A1(n13137), .A2(n13116), .ZN(n11036) );
  AND2_X1 U13571 ( .A1(n11037), .A2(n11036), .ZN(n13022) );
  NAND2_X1 U13572 ( .A1(n11038), .A2(n13022), .ZN(n15049) );
  INV_X1 U13573 ( .A(n15049), .ZN(n11050) );
  NAND2_X1 U13574 ( .A1(n11041), .A2(n11040), .ZN(n11166) );
  OR2_X1 U13575 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  NAND2_X1 U13576 ( .A1(n11166), .A2(n11042), .ZN(n15044) );
  INV_X1 U13577 ( .A(n15044), .ZN(n11048) );
  OAI211_X1 U13578 ( .C1(n11043), .C2(n15047), .A(n13496), .B(n11192), .ZN(
        n15045) );
  OAI22_X1 U13579 ( .A1(n13543), .A2(n11044), .B1(n13025), .B2(n14938), .ZN(
        n11045) );
  AOI21_X1 U13580 ( .B1(n13518), .B2(n13024), .A(n11045), .ZN(n11046) );
  OAI21_X1 U13581 ( .B1(n15045), .B2(n13500), .A(n11046), .ZN(n11047) );
  AOI21_X1 U13582 ( .B1(n11048), .B2(n13542), .A(n11047), .ZN(n11049) );
  OAI21_X1 U13583 ( .B1(n14943), .B2(n11050), .A(n11049), .ZN(P2_U3255) );
  NAND2_X1 U13584 ( .A1(n11725), .A2(n14310), .ZN(n11051) );
  OAI211_X1 U13585 ( .C1(n11726), .C2(n6421), .A(n11051), .B(n11918), .ZN(
        P1_U3332) );
  NAND2_X1 U13586 ( .A1(n11725), .A2(n11052), .ZN(n11054) );
  OAI211_X1 U13587 ( .C1(n11055), .C2(n13686), .A(n11054), .B(n11053), .ZN(
        P2_U3304) );
  INV_X1 U13588 ( .A(n13826), .ZN(n11482) );
  OR2_X1 U13589 ( .A1(n11613), .A2(n11482), .ZN(n11056) );
  NAND2_X1 U13590 ( .A1(n11057), .A2(n11056), .ZN(n11064) );
  NAND2_X1 U13591 ( .A1(n11058), .A2(n11791), .ZN(n11063) );
  NOR2_X1 U13592 ( .A1(n11857), .A2(n11059), .ZN(n11060) );
  AOI21_X1 U13593 ( .B1(n11061), .B2(n11659), .A(n11060), .ZN(n11062) );
  XNOR2_X1 U13594 ( .A(n14469), .B(n13825), .ZN(n11889) );
  OAI211_X1 U13595 ( .C1(n11064), .C2(n11889), .A(n11160), .B(n14751), .ZN(
        n11079) );
  INV_X1 U13596 ( .A(n11889), .ZN(n11069) );
  OR2_X1 U13597 ( .A1(n11613), .A2(n13826), .ZN(n11066) );
  OAI21_X1 U13598 ( .B1(n11069), .B2(n11068), .A(n11158), .ZN(n11070) );
  NAND2_X1 U13599 ( .A1(n11070), .A2(n14762), .ZN(n11078) );
  INV_X1 U13600 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11071) );
  AND2_X1 U13601 ( .A1(n11072), .A2(n11071), .ZN(n11073) );
  OR2_X1 U13602 ( .A1(n11073), .A2(n11153), .ZN(n14550) );
  OR2_X1 U13603 ( .A1(n11820), .A2(n9693), .ZN(n11075) );
  OR2_X1 U13604 ( .A1(n6802), .A2(n14612), .ZN(n11074) );
  AND2_X1 U13605 ( .A1(n11075), .A2(n11074), .ZN(n11077) );
  NAND2_X1 U13606 ( .A1(n11707), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11076) );
  OAI211_X1 U13607 ( .C1(n14550), .C2(n11818), .A(n11077), .B(n11076), .ZN(
        n13824) );
  AOI22_X1 U13608 ( .A1(n13824), .A2(n14575), .B1(n14572), .B2(n13826), .ZN(
        n13778) );
  NAND3_X1 U13609 ( .A1(n11079), .A2(n11078), .A3(n13778), .ZN(n14468) );
  XNOR2_X1 U13610 ( .A(n11150), .B(n14469), .ZN(n11080) );
  NOR2_X1 U13611 ( .A1(n11080), .A2(n14718), .ZN(n14472) );
  NOR2_X1 U13612 ( .A1(n14468), .A2(n14472), .ZN(n11085) );
  INV_X1 U13613 ( .A(n14469), .ZN(n13783) );
  INV_X1 U13614 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11081) );
  OAI22_X1 U13615 ( .A1(n13783), .A2(n14300), .B1(n14764), .B2(n11081), .ZN(
        n11082) );
  INV_X1 U13616 ( .A(n11082), .ZN(n11083) );
  OAI21_X1 U13617 ( .B1(n11085), .B2(n14763), .A(n11083), .ZN(P1_U3498) );
  AOI22_X1 U13618 ( .A1(n14469), .A2(n14263), .B1(n6820), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11084) );
  OAI21_X1 U13619 ( .B1(n11085), .B2(n6820), .A(n11084), .ZN(P1_U3541) );
  XNOR2_X1 U13620 ( .A(n11086), .B(n12399), .ZN(n11087) );
  OAI222_X1 U13621 ( .A1(n12873), .A2(n12246), .B1(n12875), .B2(n11455), .C1(
        n11087), .C2(n15149), .ZN(n14514) );
  INV_X1 U13622 ( .A(n14514), .ZN(n11094) );
  OAI21_X1 U13623 ( .B1(n6589), .B2(n11088), .A(n12399), .ZN(n11090) );
  NAND2_X1 U13624 ( .A1(n11090), .A2(n11089), .ZN(n14516) );
  AOI22_X1 U13625 ( .A1(n15156), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15151), 
        .B2(n11451), .ZN(n11091) );
  OAI21_X1 U13626 ( .B1(n14513), .B2(n12883), .A(n11091), .ZN(n11092) );
  AOI21_X1 U13627 ( .B1(n14516), .B2(n12885), .A(n11092), .ZN(n11093) );
  OAI21_X1 U13628 ( .B1(n11094), .B2(n15156), .A(n11093), .ZN(P3_U3222) );
  XNOR2_X1 U13629 ( .A(n13024), .B(n11976), .ZN(n11098) );
  INV_X1 U13630 ( .A(n11098), .ZN(n11100) );
  NAND2_X1 U13631 ( .A1(n13136), .A2(n13529), .ZN(n11099) );
  INV_X1 U13632 ( .A(n11095), .ZN(n11097) );
  XNOR2_X1 U13633 ( .A(n11098), .B(n11099), .ZN(n13020) );
  XNOR2_X1 U13634 ( .A(n15054), .B(n11101), .ZN(n11103) );
  NAND2_X1 U13635 ( .A1(n13135), .A2(n10303), .ZN(n11102) );
  NOR2_X1 U13636 ( .A1(n11103), .A2(n11102), .ZN(n11133) );
  INV_X1 U13637 ( .A(n11133), .ZN(n11104) );
  NAND2_X1 U13638 ( .A1(n11103), .A2(n11102), .ZN(n11134) );
  NAND2_X1 U13639 ( .A1(n11104), .A2(n11134), .ZN(n11105) );
  XNOR2_X1 U13640 ( .A(n11135), .B(n11105), .ZN(n11112) );
  NAND2_X1 U13641 ( .A1(n15054), .A2(n14782), .ZN(n11110) );
  NAND2_X1 U13642 ( .A1(n13134), .A2(n13254), .ZN(n11107) );
  NAND2_X1 U13643 ( .A1(n13136), .A2(n13116), .ZN(n11106) );
  NAND2_X1 U13644 ( .A1(n11107), .A2(n11106), .ZN(n15052) );
  AOI21_X1 U13645 ( .B1(n14534), .B2(n15052), .A(n11108), .ZN(n11109) );
  OAI211_X1 U13646 ( .C1(n14797), .C2(n11188), .A(n11110), .B(n11109), .ZN(
        n11111) );
  AOI21_X1 U13647 ( .B1(n11112), .B2(n14788), .A(n11111), .ZN(n11113) );
  INV_X1 U13648 ( .A(n11113), .ZN(P2_U3208) );
  NAND2_X1 U13649 ( .A1(n14688), .A2(n12129), .ZN(n11117) );
  NAND2_X1 U13650 ( .A1(n12122), .A2(n13829), .ZN(n11116) );
  NAND2_X1 U13651 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  XNOR2_X1 U13652 ( .A(n11118), .B(n12130), .ZN(n11254) );
  NOR2_X1 U13653 ( .A1(n10184), .A2(n11119), .ZN(n11120) );
  AOI21_X1 U13654 ( .B1(n14688), .B2(n12122), .A(n11120), .ZN(n11255) );
  XNOR2_X1 U13655 ( .A(n11254), .B(n11255), .ZN(n11121) );
  OAI211_X1 U13656 ( .C1(n11122), .C2(n11121), .A(n11257), .B(n13810), .ZN(
        n11129) );
  NAND2_X1 U13657 ( .A1(n13830), .A2(n14572), .ZN(n11124) );
  NAND2_X1 U13658 ( .A1(n13828), .A2(n14575), .ZN(n11123) );
  NAND2_X1 U13659 ( .A1(n11124), .A2(n11123), .ZN(n14679) );
  NAND2_X1 U13660 ( .A1(n13805), .A2(n14679), .ZN(n11125) );
  OAI211_X1 U13661 ( .C1(n14568), .C2(n14681), .A(n11126), .B(n11125), .ZN(
        n11127) );
  AOI21_X1 U13662 ( .B1(n14688), .B2(n14564), .A(n11127), .ZN(n11128) );
  NAND2_X1 U13663 ( .A1(n11129), .A2(n11128), .ZN(P1_U3231) );
  INV_X1 U13664 ( .A(n11130), .ZN(n11132) );
  OAI222_X1 U13665 ( .A1(n14451), .A2(n11132), .B1(n12997), .B2(n15313), .C1(
        P3_U3151), .C2(n11131), .ZN(P3_U3270) );
  AOI21_X2 U13666 ( .B1(n11135), .B2(n11134), .A(n11133), .ZN(n11288) );
  XNOR2_X1 U13667 ( .A(n11243), .B(n11972), .ZN(n11138) );
  AND2_X1 U13668 ( .A1(n13134), .A2(n13529), .ZN(n11137) );
  NOR2_X1 U13669 ( .A1(n11138), .A2(n11137), .ZN(n11287) );
  INV_X1 U13670 ( .A(n11287), .ZN(n11139) );
  NAND2_X1 U13671 ( .A1(n11138), .A2(n11137), .ZN(n11286) );
  NAND2_X1 U13672 ( .A1(n11139), .A2(n11286), .ZN(n11140) );
  XNOR2_X1 U13673 ( .A(n11288), .B(n11140), .ZN(n11145) );
  AOI22_X1 U13674 ( .A1(n13116), .A2(n13135), .B1(n13133), .B2(n13254), .ZN(
        n11267) );
  INV_X1 U13675 ( .A(n11267), .ZN(n11141) );
  AOI22_X1 U13676 ( .A1(n14534), .A2(n11141), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11142) );
  OAI21_X1 U13677 ( .B1(n14797), .B2(n11179), .A(n11142), .ZN(n11143) );
  AOI21_X1 U13678 ( .B1(n11243), .B2(n14794), .A(n11143), .ZN(n11144) );
  OAI21_X1 U13679 ( .B1(n11145), .B2(n14777), .A(n11144), .ZN(P2_U3196) );
  NAND2_X1 U13680 ( .A1(n11146), .A2(n11791), .ZN(n11149) );
  AOI22_X1 U13681 ( .A1(n11147), .A2(n11659), .B1(n11660), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11148) );
  INV_X1 U13682 ( .A(n11352), .ZN(n11151) );
  AOI211_X1 U13683 ( .C1(n14606), .C2(n11152), .A(n14718), .B(n11151), .ZN(
        n14604) );
  NOR2_X1 U13684 ( .A1(n14698), .A2(n14550), .ZN(n11157) );
  NOR2_X1 U13685 ( .A1(n11153), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11154) );
  OR2_X1 U13686 ( .A1(n11346), .A2(n11154), .ZN(n13813) );
  AOI22_X1 U13687 ( .A1(n11817), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n11707), 
        .B2(P1_REG0_REG_15__SCAN_IN), .ZN(n11156) );
  INV_X1 U13688 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11354) );
  OR2_X1 U13689 ( .A1(n11820), .A2(n11354), .ZN(n11155) );
  OAI211_X1 U13690 ( .C1(n13813), .C2(n11818), .A(n11156), .B(n11155), .ZN(
        n13823) );
  INV_X1 U13691 ( .A(n13823), .ZN(n14553) );
  INV_X1 U13692 ( .A(n13825), .ZN(n14539) );
  OAI22_X1 U13693 ( .A1(n14553), .A2(n11394), .B1(n14539), .B2(n14165), .ZN(
        n14605) );
  AOI211_X1 U13694 ( .C1(n14604), .C2(n14471), .A(n11157), .B(n14605), .ZN(
        n11165) );
  INV_X1 U13695 ( .A(n13824), .ZN(n12026) );
  OR2_X1 U13696 ( .A1(n14606), .A2(n12026), .ZN(n11622) );
  NAND2_X1 U13697 ( .A1(n14606), .A2(n12026), .ZN(n11624) );
  NAND2_X1 U13698 ( .A1(n11622), .A2(n11624), .ZN(n11891) );
  INV_X1 U13699 ( .A(n11891), .ZN(n11161) );
  OAI21_X1 U13700 ( .B1(n6576), .B2(n11891), .A(n11336), .ZN(n14608) );
  INV_X1 U13701 ( .A(n14608), .ZN(n11162) );
  OR2_X1 U13702 ( .A1(n14469), .A2(n14539), .ZN(n11159) );
  OAI21_X1 U13703 ( .B1(n6452), .B2(n11161), .A(n7177), .ZN(n14611) );
  NOR2_X1 U13704 ( .A1(n14684), .A2(n14570), .ZN(n14181) );
  AOI22_X1 U13705 ( .A1(n14712), .A2(n11162), .B1(n14611), .B2(n14181), .ZN(
        n11164) );
  AOI22_X1 U13706 ( .A1(n14606), .A2(n14702), .B1(n14684), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n11163) );
  OAI211_X1 U13707 ( .C1(n14684), .C2(n11165), .A(n11164), .B(n11163), .ZN(
        P1_U3279) );
  NAND2_X1 U13708 ( .A1(n11166), .A2(n7539), .ZN(n11186) );
  INV_X1 U13709 ( .A(n15054), .ZN(n11167) );
  NAND2_X1 U13710 ( .A1(n11167), .A2(n11176), .ZN(n11169) );
  XOR2_X1 U13711 ( .A(n11239), .B(n11178), .Z(n11273) );
  NAND2_X1 U13712 ( .A1(n13024), .A2(n11172), .ZN(n11173) );
  NAND2_X1 U13713 ( .A1(n11174), .A2(n11173), .ZN(n11185) );
  INV_X1 U13714 ( .A(n11187), .ZN(n11175) );
  NAND2_X1 U13715 ( .A1(n15054), .A2(n11176), .ZN(n11177) );
  XOR2_X1 U13716 ( .A(n11241), .B(n11178), .Z(n11271) );
  INV_X1 U13717 ( .A(n11243), .ZN(n11268) );
  AOI211_X1 U13718 ( .C1(n11243), .C2(n6590), .A(n13529), .B(n11248), .ZN(
        n11270) );
  NAND2_X1 U13719 ( .A1(n11270), .A2(n13535), .ZN(n11182) );
  OAI22_X1 U13720 ( .A1(n14943), .A2(n11267), .B1(n11179), .B2(n14938), .ZN(
        n11180) );
  AOI21_X1 U13721 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n14943), .A(n11180), 
        .ZN(n11181) );
  OAI211_X1 U13722 ( .C1(n11268), .C2(n13533), .A(n11182), .B(n11181), .ZN(
        n11183) );
  AOI21_X1 U13723 ( .B1(n11271), .B2(n13541), .A(n11183), .ZN(n11184) );
  OAI21_X1 U13724 ( .B1(n11273), .B2(n13524), .A(n11184), .ZN(P2_U3253) );
  XNOR2_X1 U13725 ( .A(n11185), .B(n11187), .ZN(n15058) );
  XNOR2_X1 U13726 ( .A(n11186), .B(n11187), .ZN(n15060) );
  INV_X1 U13727 ( .A(n15060), .ZN(n15063) );
  NAND2_X1 U13728 ( .A1(n15063), .A2(n13542), .ZN(n11197) );
  INV_X1 U13729 ( .A(n11188), .ZN(n11189) );
  AOI22_X1 U13730 ( .A1(n14941), .A2(n15052), .B1(n11189), .B2(n13493), .ZN(
        n11190) );
  OAI21_X1 U13731 ( .B1(n11191), .B2(n13543), .A(n11190), .ZN(n11195) );
  AOI21_X1 U13732 ( .B1(n11192), .B2(n15054), .A(n13529), .ZN(n11193) );
  NAND2_X1 U13733 ( .A1(n11193), .A2(n6590), .ZN(n15055) );
  NOR2_X1 U13734 ( .A1(n15055), .A2(n13500), .ZN(n11194) );
  AOI211_X1 U13735 ( .C1(n13518), .C2(n15054), .A(n11195), .B(n11194), .ZN(
        n11196) );
  OAI211_X1 U13736 ( .C1(n15058), .C2(n13473), .A(n11197), .B(n11196), .ZN(
        P2_U3254) );
  OAI222_X1 U13737 ( .A1(P3_U3151), .A2(n6848), .B1(n14451), .B2(n11199), .C1(
        n11198), .C2(n12997), .ZN(P3_U3269) );
  NAND2_X1 U13738 ( .A1(n12281), .A2(n11200), .ZN(n11204) );
  INV_X1 U13739 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11201) );
  NOR2_X1 U13740 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11201), .ZN(n15096) );
  AOI21_X1 U13741 ( .B1(n12282), .B2(n11202), .A(n15096), .ZN(n11203) );
  OAI211_X1 U13742 ( .C1(n11205), .C2(n12285), .A(n11204), .B(n11203), .ZN(
        n11210) );
  AOI211_X1 U13743 ( .C1(n11208), .C2(n11207), .A(n12289), .B(n11206), .ZN(
        n11209) );
  AOI211_X1 U13744 ( .C1(n15183), .C2(n12287), .A(n11210), .B(n11209), .ZN(
        n11211) );
  INV_X1 U13745 ( .A(n11211), .ZN(P3_U3157) );
  INV_X1 U13746 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U13747 ( .A1(n11632), .A2(n11212), .ZN(n11213) );
  NAND2_X1 U13748 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  XNOR2_X1 U13749 ( .A(n11215), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n11222) );
  AOI21_X1 U13750 ( .B1(n11222), .B2(n13914), .A(n14666), .ZN(n11221) );
  NAND2_X1 U13751 ( .A1(n11632), .A2(n11216), .ZN(n11217) );
  NAND2_X1 U13752 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  XNOR2_X1 U13753 ( .A(n11219), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U13754 ( .A1(n11223), .A2(n13908), .ZN(n11220) );
  NAND2_X1 U13755 ( .A1(n11221), .A2(n11220), .ZN(n11225) );
  OAI22_X1 U13756 ( .A1(n11223), .A2(n14669), .B1(n11222), .B2(n14663), .ZN(
        n11224) );
  MUX2_X1 U13757 ( .A(n11225), .B(n11224), .S(n14471), .Z(n11226) );
  INV_X1 U13758 ( .A(n11226), .ZN(n11227) );
  NAND2_X1 U13759 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13710)
         );
  OAI211_X1 U13760 ( .C1(n11228), .C2(n14674), .A(n11227), .B(n13710), .ZN(
        P1_U3262) );
  XNOR2_X1 U13761 ( .A(n11229), .B(n12314), .ZN(n14509) );
  XNOR2_X1 U13762 ( .A(n11230), .B(n12314), .ZN(n11231) );
  OAI222_X1 U13763 ( .A1(n12875), .A2(n12181), .B1(n12873), .B2(n11468), .C1(
        n11231), .C2(n15149), .ZN(n14510) );
  NAND2_X1 U13764 ( .A1(n14510), .A2(n15154), .ZN(n11235) );
  INV_X1 U13765 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11311) );
  INV_X1 U13766 ( .A(n12177), .ZN(n11232) );
  OAI22_X1 U13767 ( .A1(n15154), .A2(n11311), .B1(n11232), .B2(n11405), .ZN(
        n11233) );
  AOI21_X1 U13768 ( .B1(n12741), .B2(n14512), .A(n11233), .ZN(n11234) );
  OAI211_X1 U13769 ( .C1(n12806), .C2(n14509), .A(n11235), .B(n11234), .ZN(
        P3_U3221) );
  INV_X1 U13770 ( .A(n11741), .ZN(n11364) );
  OAI222_X1 U13771 ( .A1(n11238), .A2(n11237), .B1(n13688), .B2(n11364), .C1(
        n11236), .C2(P2_U3088), .ZN(P2_U3303) );
  OAI21_X1 U13772 ( .B1(n11268), .B2(n11242), .A(n11239), .ZN(n11240) );
  OAI21_X1 U13773 ( .B1(n13134), .B2(n11243), .A(n11240), .ZN(n11412) );
  XOR2_X1 U13774 ( .A(n11412), .B(n11246), .Z(n11431) );
  OR2_X1 U13775 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  XNOR2_X1 U13776 ( .A(n11417), .B(n11246), .ZN(n11429) );
  INV_X1 U13777 ( .A(n11418), .ZN(n11247) );
  OAI211_X1 U13778 ( .C1(n11427), .C2(n11248), .A(n11247), .B(n13496), .ZN(
        n11426) );
  AOI22_X1 U13779 ( .A1(n13116), .A2(n13134), .B1(n13132), .B2(n13254), .ZN(
        n14786) );
  OAI22_X1 U13780 ( .A1(n14943), .A2(n14786), .B1(n14798), .B2(n14938), .ZN(
        n11250) );
  NOR2_X1 U13781 ( .A1(n11427), .A2(n13533), .ZN(n11249) );
  AOI211_X1 U13782 ( .C1(n14943), .C2(P2_REG2_REG_13__SCAN_IN), .A(n11250), 
        .B(n11249), .ZN(n11251) );
  OAI21_X1 U13783 ( .B1(n11426), .B2(n13500), .A(n11251), .ZN(n11252) );
  AOI21_X1 U13784 ( .B1(n11429), .B2(n13541), .A(n11252), .ZN(n11253) );
  OAI21_X1 U13785 ( .B1(n11431), .B2(n13524), .A(n11253), .ZN(P2_U3252) );
  INV_X1 U13786 ( .A(n11254), .ZN(n11256) );
  NOR2_X1 U13787 ( .A1(n10184), .A2(n11258), .ZN(n11259) );
  AOI21_X1 U13788 ( .B1(n14756), .B2(n12122), .A(n11259), .ZN(n11435) );
  AOI22_X1 U13789 ( .A1(n14756), .A2(n12129), .B1(n12122), .B2(n13828), .ZN(
        n11260) );
  XNOR2_X1 U13790 ( .A(n11260), .B(n12130), .ZN(n11434) );
  XOR2_X1 U13791 ( .A(n11435), .B(n11434), .Z(n11261) );
  OAI211_X1 U13792 ( .C1(n11262), .C2(n11261), .A(n11439), .B(n13810), .ZN(
        n11266) );
  NAND2_X1 U13793 ( .A1(n13829), .A2(n14572), .ZN(n14186) );
  NAND2_X1 U13794 ( .A1(n13827), .A2(n14575), .ZN(n14185) );
  NAND2_X1 U13795 ( .A1(n14186), .A2(n14185), .ZN(n14754) );
  NOR2_X1 U13796 ( .A1(n14568), .A2(n14177), .ZN(n11263) );
  AOI211_X1 U13797 ( .C1(n13805), .C2(n14754), .A(n11264), .B(n11263), .ZN(
        n11265) );
  OAI211_X1 U13798 ( .C1(n6993), .C2(n13821), .A(n11266), .B(n11265), .ZN(
        P1_U3217) );
  INV_X1 U13799 ( .A(n15053), .ZN(n15046) );
  OAI21_X1 U13800 ( .B1(n11268), .B2(n15046), .A(n11267), .ZN(n11269) );
  AOI211_X1 U13801 ( .C1(n11271), .C2(n15026), .A(n11270), .B(n11269), .ZN(
        n11272) );
  OAI21_X1 U13802 ( .B1(n11273), .B2(n15022), .A(n11272), .ZN(n11275) );
  NAND2_X1 U13803 ( .A1(n11275), .A2(n15081), .ZN(n11274) );
  OAI21_X1 U13804 ( .B1(n15081), .B2(n8612), .A(n11274), .ZN(P2_U3511) );
  INV_X1 U13805 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11277) );
  NAND2_X1 U13806 ( .A1(n11275), .A2(n15066), .ZN(n11276) );
  OAI21_X1 U13807 ( .B1(n15066), .B2(n11277), .A(n11276), .ZN(P2_U3466) );
  XNOR2_X1 U13808 ( .A(n11278), .B(n12406), .ZN(n14505) );
  XNOR2_X1 U13809 ( .A(n11279), .B(n12406), .ZN(n11280) );
  OAI222_X1 U13810 ( .A1(n12875), .A2(n12246), .B1(n12873), .B2(n12874), .C1(
        n11280), .C2(n15149), .ZN(n14507) );
  NAND2_X1 U13811 ( .A1(n14507), .A2(n15154), .ZN(n11285) );
  INV_X1 U13812 ( .A(n14504), .ZN(n11283) );
  INV_X1 U13813 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11308) );
  INV_X1 U13814 ( .A(n12242), .ZN(n11281) );
  OAI22_X1 U13815 ( .A1(n15154), .A2(n11308), .B1(n11281), .B2(n11405), .ZN(
        n11282) );
  AOI21_X1 U13816 ( .B1(n11283), .B2(n12741), .A(n11282), .ZN(n11284) );
  OAI211_X1 U13817 ( .C1(n12806), .C2(n14505), .A(n11285), .B(n11284), .ZN(
        P3_U3220) );
  XNOR2_X1 U13818 ( .A(n14795), .B(n11101), .ZN(n11295) );
  NAND2_X1 U13819 ( .A1(n13133), .A2(n10303), .ZN(n11289) );
  NOR2_X1 U13820 ( .A1(n11295), .A2(n11289), .ZN(n11290) );
  AOI21_X1 U13821 ( .B1(n11295), .B2(n11289), .A(n11290), .ZN(n14789) );
  NAND2_X1 U13822 ( .A1(n14790), .A2(n14789), .ZN(n11293) );
  XNOR2_X1 U13823 ( .A(n11512), .B(n11976), .ZN(n11494) );
  NAND2_X1 U13824 ( .A1(n13132), .A2(n10303), .ZN(n11492) );
  XNOR2_X1 U13825 ( .A(n11494), .B(n11492), .ZN(n11296) );
  INV_X1 U13826 ( .A(n11290), .ZN(n11291) );
  NAND2_X1 U13827 ( .A1(n11293), .A2(n11292), .ZN(n11496) );
  NAND2_X1 U13828 ( .A1(n13096), .A2(n13133), .ZN(n11294) );
  OAI22_X1 U13829 ( .A1(n11293), .A2(n14777), .B1(n11295), .B2(n11294), .ZN(
        n11298) );
  INV_X1 U13830 ( .A(n11296), .ZN(n11297) );
  NAND2_X1 U13831 ( .A1(n11298), .A2(n11297), .ZN(n11303) );
  NOR2_X1 U13832 ( .A1(n14797), .A2(n11420), .ZN(n11301) );
  AOI22_X1 U13833 ( .A1(n13116), .A2(n13133), .B1(n13131), .B2(n13254), .ZN(
        n13644) );
  OAI22_X1 U13834 ( .A1(n14787), .A2(n13644), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11299), .ZN(n11300) );
  AOI211_X1 U13835 ( .C1(n11512), .C2(n14782), .A(n11301), .B(n11300), .ZN(
        n11302) );
  OAI211_X1 U13836 ( .C1(n11496), .C2(n14777), .A(n11303), .B(n11302), .ZN(
        P2_U3187) );
  INV_X1 U13837 ( .A(n14455), .ZN(n12532) );
  NOR2_X1 U13838 ( .A1(n11324), .A2(n11304), .ZN(n11306) );
  MUX2_X1 U13839 ( .A(n11311), .B(P3_REG2_REG_12__SCAN_IN), .S(n15123), .Z(
        n15116) );
  AOI21_X1 U13840 ( .B1(n11308), .B2(n11307), .A(n12527), .ZN(n11334) );
  OR2_X1 U13841 ( .A1(n12626), .A2(n11308), .ZN(n11310) );
  NAND2_X1 U13842 ( .A1(n12626), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n11309) );
  AND2_X1 U13843 ( .A1(n11310), .A2(n11309), .ZN(n12533) );
  XNOR2_X1 U13844 ( .A(n12533), .B(n12532), .ZN(n11319) );
  INV_X1 U13845 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11327) );
  MUX2_X1 U13846 ( .A(n11311), .B(n11327), .S(n12675), .Z(n11313) );
  OR2_X1 U13847 ( .A1(n11312), .A2(n11313), .ZN(n11317) );
  XNOR2_X1 U13848 ( .A(n11313), .B(n15123), .ZN(n15133) );
  INV_X1 U13849 ( .A(n11314), .ZN(n11316) );
  AOI21_X1 U13850 ( .B1(n11324), .B2(n11316), .A(n11315), .ZN(n15132) );
  NAND2_X1 U13851 ( .A1(n15133), .A2(n15132), .ZN(n15130) );
  NAND2_X1 U13852 ( .A1(n11317), .A2(n15130), .ZN(n11318) );
  AOI21_X1 U13853 ( .B1(n11319), .B2(n11318), .A(n12534), .ZN(n11322) );
  NAND2_X1 U13854 ( .A1(n15082), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n11321) );
  AND2_X1 U13855 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12243) );
  INV_X1 U13856 ( .A(n12243), .ZN(n11320) );
  OAI211_X1 U13857 ( .C1(n11322), .C2(n15110), .A(n11321), .B(n11320), .ZN(
        n11332) );
  INV_X1 U13858 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14508) );
  NOR2_X1 U13859 ( .A1(n11324), .A2(n11323), .ZN(n11326) );
  MUX2_X1 U13860 ( .A(n11327), .B(P3_REG1_REG_12__SCAN_IN), .S(n15123), .Z(
        n15120) );
  NAND2_X1 U13861 ( .A1(n15123), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11328) );
  AOI21_X1 U13862 ( .B1(n14508), .B2(n11329), .A(n12523), .ZN(n11330) );
  NOR2_X1 U13863 ( .A1(n11330), .A2(n15125), .ZN(n11331) );
  AOI211_X1 U13864 ( .C1(n15106), .C2(n12532), .A(n11332), .B(n11331), .ZN(
        n11333) );
  OAI21_X1 U13865 ( .B1(n11334), .B2(n15136), .A(n11333), .ZN(P3_U3195) );
  NAND2_X1 U13866 ( .A1(n14606), .A2(n13824), .ZN(n11335) );
  NAND2_X1 U13867 ( .A1(n11336), .A2(n11335), .ZN(n11381) );
  NAND2_X1 U13868 ( .A1(n11337), .A2(n11791), .ZN(n11342) );
  OAI22_X1 U13869 ( .A1(n11339), .A2(n11715), .B1(n11857), .B2(n11338), .ZN(
        n11340) );
  INV_X1 U13870 ( .A(n11340), .ZN(n11341) );
  NAND2_X1 U13871 ( .A1(n12036), .A2(n14553), .ZN(n11626) );
  NAND2_X1 U13872 ( .A1(n11629), .A2(n11626), .ZN(n11893) );
  XNOR2_X1 U13873 ( .A(n11381), .B(n11893), .ZN(n11367) );
  OAI211_X1 U13874 ( .C1(n11345), .C2(n11380), .A(n11374), .B(n14751), .ZN(
        n11351) );
  OR2_X1 U13875 ( .A1(n11346), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U13876 ( .A1(n11386), .A2(n11347), .ZN(n14567) );
  INV_X1 U13877 ( .A(n11820), .ZN(n11830) );
  AOI22_X1 U13878 ( .A1(n11830), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11707), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U13879 ( .A1(n11817), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11348) );
  OAI211_X1 U13880 ( .C1(n14567), .C2(n11818), .A(n11349), .B(n11348), .ZN(
        n14573) );
  AND2_X1 U13881 ( .A1(n13824), .A2(n14572), .ZN(n11350) );
  AOI21_X1 U13882 ( .B1(n14573), .B2(n14575), .A(n11350), .ZN(n13814) );
  AND2_X1 U13883 ( .A1(n11351), .A2(n13814), .ZN(n11366) );
  INV_X1 U13884 ( .A(n11366), .ZN(n11358) );
  NAND2_X1 U13885 ( .A1(n12036), .A2(n11352), .ZN(n11353) );
  NAND3_X1 U13886 ( .A1(n11384), .A2(n14707), .A3(n11353), .ZN(n11365) );
  OAI22_X1 U13887 ( .A1(n14700), .A2(n11354), .B1(n13813), .B2(n14698), .ZN(
        n11355) );
  AOI21_X1 U13888 ( .B1(n12036), .B2(n14702), .A(n11355), .ZN(n11356) );
  OAI21_X1 U13889 ( .B1(n11365), .B2(n14173), .A(n11356), .ZN(n11357) );
  AOI21_X1 U13890 ( .B1(n11358), .B2(n14700), .A(n11357), .ZN(n11359) );
  OAI21_X1 U13891 ( .B1(n14114), .B2(n11367), .A(n11359), .ZN(P1_U3278) );
  INV_X1 U13892 ( .A(n11754), .ZN(n11362) );
  OAI222_X1 U13893 ( .A1(P1_U3086), .A2(n11360), .B1(n11530), .B2(n11362), 
        .C1(n11755), .C2(n6421), .ZN(P1_U3330) );
  OAI222_X1 U13894 ( .A1(n13686), .A2(n11363), .B1(n13688), .B2(n11362), .C1(
        n11361), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U13895 ( .A1(P1_U3086), .A2(n11532), .B1(n11530), .B2(n11364), 
        .C1(n11742), .C2(n6421), .ZN(P1_U3331) );
  OAI211_X1 U13896 ( .C1(n11367), .C2(n14609), .A(n11366), .B(n11365), .ZN(
        n11372) );
  INV_X1 U13897 ( .A(n12036), .ZN(n13822) );
  INV_X1 U13898 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11368) );
  OAI22_X1 U13899 ( .A1(n13822), .A2(n14259), .B1(n14772), .B2(n11368), .ZN(
        n11369) );
  AOI21_X1 U13900 ( .B1(n11372), .B2(n14772), .A(n11369), .ZN(n11370) );
  INV_X1 U13901 ( .A(n11370), .ZN(P1_U3543) );
  INV_X1 U13902 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15216) );
  OAI22_X1 U13903 ( .A1(n13822), .A2(n14300), .B1(n14764), .B2(n15216), .ZN(
        n11371) );
  AOI21_X1 U13904 ( .B1(n11372), .B2(n14764), .A(n11371), .ZN(n11373) );
  INV_X1 U13905 ( .A(n11373), .ZN(P1_U3504) );
  NAND2_X1 U13906 ( .A1(n11375), .A2(n11791), .ZN(n11377) );
  AOI22_X1 U13907 ( .A1(n13912), .A2(n11659), .B1(n11660), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n11376) );
  INV_X1 U13908 ( .A(n14573), .ZN(n13972) );
  XNOR2_X1 U13909 ( .A(n14598), .B(n13972), .ZN(n11892) );
  INV_X1 U13910 ( .A(n11892), .ZN(n11378) );
  OAI21_X1 U13911 ( .B1(n11379), .B2(n11378), .A(n13934), .ZN(n14602) );
  INV_X1 U13912 ( .A(n14602), .ZN(n11400) );
  INV_X1 U13913 ( .A(n14181), .ZN(n14107) );
  OR2_X1 U13914 ( .A1(n12036), .A2(n13823), .ZN(n11382) );
  OAI21_X1 U13915 ( .B1(n11383), .B2(n11892), .A(n13975), .ZN(n14595) );
  AOI211_X1 U13916 ( .C1(n14598), .C2(n11384), .A(n14718), .B(n14585), .ZN(
        n14596) );
  NOR2_X1 U13917 ( .A1(n14698), .A2(n14567), .ZN(n11395) );
  INV_X1 U13918 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U13919 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  AND2_X1 U13920 ( .A1(n11636), .A2(n11387), .ZN(n14578) );
  NAND2_X1 U13921 ( .A1(n14578), .A2(n11706), .ZN(n11393) );
  NAND2_X1 U13922 ( .A1(n11707), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13923 ( .A1(n11830), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11388) );
  OAI211_X1 U13924 ( .C1(n6802), .C2(n11390), .A(n11389), .B(n11388), .ZN(
        n11391) );
  INV_X1 U13925 ( .A(n11391), .ZN(n11392) );
  NAND2_X1 U13926 ( .A1(n11393), .A2(n11392), .ZN(n13935) );
  INV_X1 U13927 ( .A(n13935), .ZN(n14552) );
  OAI22_X1 U13928 ( .A1(n14552), .A2(n11394), .B1(n14553), .B2(n14165), .ZN(
        n14597) );
  AOI211_X1 U13929 ( .C1(n14596), .C2(n14471), .A(n11395), .B(n14597), .ZN(
        n11397) );
  AOI22_X1 U13930 ( .A1(n14598), .A2(n14702), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14684), .ZN(n11396) );
  OAI21_X1 U13931 ( .B1(n11397), .B2(n14684), .A(n11396), .ZN(n11398) );
  AOI21_X1 U13932 ( .B1(n14712), .B2(n14595), .A(n11398), .ZN(n11399) );
  OAI21_X1 U13933 ( .B1(n11400), .B2(n14107), .A(n11399), .ZN(P1_U3277) );
  XNOR2_X1 U13934 ( .A(n11401), .B(n7423), .ZN(n14500) );
  XNOR2_X1 U13935 ( .A(n11403), .B(n11402), .ZN(n11404) );
  OAI222_X1 U13936 ( .A1(n12875), .A2(n11468), .B1(n12873), .B2(n12206), .C1(
        n11404), .C2(n15149), .ZN(n14502) );
  NAND2_X1 U13937 ( .A1(n14502), .A2(n15154), .ZN(n11411) );
  INV_X1 U13938 ( .A(n14499), .ZN(n11409) );
  INV_X1 U13939 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11407) );
  INV_X1 U13940 ( .A(n11471), .ZN(n11406) );
  OAI22_X1 U13941 ( .A1(n15154), .A2(n11407), .B1(n11406), .B2(n11405), .ZN(
        n11408) );
  AOI21_X1 U13942 ( .B1(n11409), .B2(n12741), .A(n11408), .ZN(n11410) );
  OAI211_X1 U13943 ( .C1(n12806), .C2(n14500), .A(n11411), .B(n11410), .ZN(
        P3_U3219) );
  XNOR2_X1 U13944 ( .A(n11504), .B(n11509), .ZN(n13650) );
  INV_X1 U13945 ( .A(n11414), .ZN(n11415) );
  XNOR2_X1 U13946 ( .A(n11510), .B(n11509), .ZN(n13648) );
  INV_X1 U13947 ( .A(n11512), .ZN(n13646) );
  OAI211_X1 U13948 ( .C1(n13646), .C2(n11418), .A(n13496), .B(n11506), .ZN(
        n13645) );
  NOR2_X1 U13949 ( .A1(n13543), .A2(n11419), .ZN(n11422) );
  OAI22_X1 U13950 ( .A1(n14943), .A2(n13644), .B1(n11420), .B2(n14938), .ZN(
        n11421) );
  AOI211_X1 U13951 ( .C1(n11512), .C2(n13518), .A(n11422), .B(n11421), .ZN(
        n11423) );
  OAI21_X1 U13952 ( .B1(n13645), .B2(n13500), .A(n11423), .ZN(n11424) );
  AOI21_X1 U13953 ( .B1(n13648), .B2(n13541), .A(n11424), .ZN(n11425) );
  OAI21_X1 U13954 ( .B1(n13650), .B2(n13524), .A(n11425), .ZN(P2_U3251) );
  OAI211_X1 U13955 ( .C1(n11427), .C2(n15046), .A(n11426), .B(n14786), .ZN(
        n11428) );
  AOI21_X1 U13956 ( .B1(n11429), .B2(n15026), .A(n11428), .ZN(n11430) );
  OAI21_X1 U13957 ( .B1(n11431), .B2(n15022), .A(n11430), .ZN(n11449) );
  NAND2_X1 U13958 ( .A1(n11449), .A2(n15081), .ZN(n11432) );
  OAI21_X1 U13959 ( .B1(n15081), .B2(n13229), .A(n11432), .ZN(P2_U3512) );
  AOI22_X1 U13960 ( .A1(n11609), .A2(n12129), .B1(n12122), .B2(n13827), .ZN(
        n11433) );
  XNOR2_X1 U13961 ( .A(n11433), .B(n12130), .ZN(n11474) );
  AOI22_X1 U13962 ( .A1(n11609), .A2(n12122), .B1(n9562), .B2(n13827), .ZN(
        n11475) );
  XNOR2_X1 U13963 ( .A(n11474), .B(n11475), .ZN(n11441) );
  INV_X1 U13964 ( .A(n11435), .ZN(n11436) );
  AOI21_X1 U13965 ( .B1(n11441), .B2(n11440), .A(n11478), .ZN(n11448) );
  OAI21_X1 U13966 ( .B1(n14551), .B2(n11482), .A(n11442), .ZN(n11443) );
  AOI21_X1 U13967 ( .B1(n13794), .B2(n13828), .A(n11443), .ZN(n11444) );
  OAI21_X1 U13968 ( .B1(n11445), .B2(n14568), .A(n11444), .ZN(n11446) );
  AOI21_X1 U13969 ( .B1(n11609), .B2(n14564), .A(n11446), .ZN(n11447) );
  OAI21_X1 U13970 ( .B1(n11448), .B2(n14559), .A(n11447), .ZN(P1_U3236) );
  NAND2_X1 U13971 ( .A1(n11449), .A2(n15066), .ZN(n11450) );
  OAI21_X1 U13972 ( .B1(n15066), .B2(n8634), .A(n11450), .ZN(P2_U3469) );
  NAND2_X1 U13973 ( .A1(n12281), .A2(n11451), .ZN(n11454) );
  AOI21_X1 U13974 ( .B1(n12282), .B2(n12513), .A(n11452), .ZN(n11453) );
  OAI211_X1 U13975 ( .C1(n11455), .C2(n12285), .A(n11454), .B(n11453), .ZN(
        n11461) );
  NAND2_X1 U13976 ( .A1(n11457), .A2(n11456), .ZN(n11458) );
  XNOR2_X1 U13977 ( .A(n11458), .B(n12181), .ZN(n11459) );
  NOR2_X1 U13978 ( .A1(n11459), .A2(n12289), .ZN(n11460) );
  AOI211_X1 U13979 ( .C1(n11462), .C2(n12287), .A(n11461), .B(n11460), .ZN(
        n11463) );
  INV_X1 U13980 ( .A(n11463), .ZN(P3_U3176) );
  XNOR2_X1 U13981 ( .A(n11464), .B(n11465), .ZN(n11473) );
  INV_X1 U13982 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11466) );
  NOR2_X1 U13983 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11466), .ZN(n12531) );
  AOI21_X1 U13984 ( .B1(n12282), .B2(n12855), .A(n12531), .ZN(n11467) );
  OAI21_X1 U13985 ( .B1(n12285), .B2(n11468), .A(n11467), .ZN(n11470) );
  NOR2_X1 U13986 ( .A1(n14499), .A2(n12278), .ZN(n11469) );
  AOI211_X1 U13987 ( .C1(n11471), .C2(n12281), .A(n11470), .B(n11469), .ZN(
        n11472) );
  OAI21_X1 U13988 ( .B1(n11473), .B2(n12289), .A(n11472), .ZN(P3_U3155) );
  INV_X1 U13989 ( .A(n11474), .ZN(n11477) );
  INV_X1 U13990 ( .A(n11475), .ZN(n11476) );
  NAND2_X1 U13991 ( .A1(n11613), .A2(n12129), .ZN(n11480) );
  NAND2_X1 U13992 ( .A1(n12122), .A2(n13826), .ZN(n11479) );
  NAND2_X1 U13993 ( .A1(n11480), .A2(n11479), .ZN(n11481) );
  XNOR2_X1 U13994 ( .A(n11481), .B(n12130), .ZN(n12017) );
  NOR2_X1 U13995 ( .A1(n10184), .A2(n11482), .ZN(n11483) );
  AOI21_X1 U13996 ( .B1(n11613), .B2(n12122), .A(n11483), .ZN(n12018) );
  XNOR2_X1 U13997 ( .A(n12017), .B(n12018), .ZN(n11484) );
  OAI211_X1 U13998 ( .C1(n6588), .C2(n11484), .A(n12020), .B(n13810), .ZN(
        n11490) );
  NOR2_X1 U13999 ( .A1(n14568), .A2(n11485), .ZN(n11488) );
  OAI22_X1 U14000 ( .A1(n14551), .A2(n14539), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11486), .ZN(n11487) );
  AOI211_X1 U14001 ( .C1(n13794), .C2(n13827), .A(n11488), .B(n11487), .ZN(
        n11489) );
  OAI211_X1 U14002 ( .C1(n11491), .C2(n13821), .A(n11490), .B(n11489), .ZN(
        P1_U3224) );
  INV_X1 U14003 ( .A(n11492), .ZN(n11493) );
  NAND2_X1 U14004 ( .A1(n11496), .A2(n11495), .ZN(n11921) );
  XNOR2_X1 U14005 ( .A(n13640), .B(n11972), .ZN(n11919) );
  XNOR2_X1 U14006 ( .A(n11921), .B(n11919), .ZN(n11498) );
  NAND2_X1 U14007 ( .A1(n11498), .A2(n11497), .ZN(n11923) );
  INV_X1 U14008 ( .A(n11923), .ZN(n11503) );
  AOI22_X1 U14009 ( .A1(n11498), .A2(n14788), .B1(n13096), .B2(n13131), .ZN(
        n11502) );
  INV_X1 U14010 ( .A(n13254), .ZN(n13510) );
  INV_X1 U14011 ( .A(n13132), .ZN(n11511) );
  OAI22_X1 U14012 ( .A1(n13300), .A2(n13510), .B1(n11511), .B2(n13508), .ZN(
        n11514) );
  AOI22_X1 U14013 ( .A1(n14534), .A2(n11514), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11499) );
  OAI21_X1 U14014 ( .B1(n14797), .B2(n11516), .A(n11499), .ZN(n11500) );
  AOI21_X1 U14015 ( .B1(n13640), .B2(n14794), .A(n11500), .ZN(n11501) );
  OAI21_X1 U14016 ( .B1(n11503), .B2(n11502), .A(n11501), .ZN(P2_U3213) );
  XNOR2_X1 U14017 ( .A(n13298), .B(n13295), .ZN(n13643) );
  OR2_X2 U14018 ( .A1(n11506), .A2(n13640), .ZN(n13519) );
  INV_X1 U14019 ( .A(n13519), .ZN(n11505) );
  AOI211_X1 U14020 ( .C1(n13640), .C2(n11506), .A(n13529), .B(n11505), .ZN(
        n13639) );
  INV_X1 U14021 ( .A(n13640), .ZN(n13296) );
  OAI22_X1 U14022 ( .A1(n13296), .A2(n13533), .B1(n14941), .B2(n11507), .ZN(
        n11508) );
  AOI21_X1 U14023 ( .B1(n13639), .B2(n13535), .A(n11508), .ZN(n11519) );
  NAND2_X1 U14024 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  XNOR2_X1 U14025 ( .A(n13264), .B(n13295), .ZN(n11515) );
  AOI21_X1 U14026 ( .B1(n11515), .B2(n15026), .A(n11514), .ZN(n13642) );
  OAI21_X1 U14027 ( .B1(n11516), .B2(n14938), .A(n13642), .ZN(n11517) );
  NAND2_X1 U14028 ( .A1(n11517), .A2(n14941), .ZN(n11518) );
  OAI211_X1 U14029 ( .C1(n13643), .C2(n13524), .A(n11519), .B(n11518), .ZN(
        P2_U3250) );
  NAND2_X1 U14030 ( .A1(n14312), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14031 ( .A1(n12000), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12291) );
  INV_X1 U14032 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U14033 ( .A1(n11835), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11523) );
  AND2_X1 U14034 ( .A1(n12291), .A2(n11523), .ZN(n11525) );
  INV_X1 U14035 ( .A(n11524), .ZN(n11526) );
  NAND2_X1 U14036 ( .A1(n11526), .A2(n6729), .ZN(n11527) );
  NAND2_X1 U14037 ( .A1(n12292), .A2(n11527), .ZN(n12297) );
  INV_X1 U14038 ( .A(n12297), .ZN(n11528) );
  INV_X1 U14039 ( .A(SI_30_), .ZN(n12298) );
  OAI222_X1 U14040 ( .A1(P3_U3151), .A2(n11529), .B1(n14451), .B2(n11528), 
        .C1(n12298), .C2(n12997), .ZN(P3_U3265) );
  INV_X1 U14041 ( .A(n11834), .ZN(n11999) );
  OAI222_X1 U14042 ( .A1(P1_U3086), .A2(n11531), .B1(n11530), .B2(n11999), 
        .C1(n11835), .C2(n6421), .ZN(P1_U3325) );
  INV_X1 U14043 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14044 ( .A1(n6405), .A2(n11534), .B1(n11533), .B2(n11532), .ZN(
        P1_U3445) );
  NAND2_X1 U14045 ( .A1(n11547), .A2(n11535), .ZN(n11539) );
  NAND2_X1 U14046 ( .A1(n11537), .A2(n11870), .ZN(n11839) );
  NAND2_X1 U14047 ( .A1(n11537), .A2(n11869), .ZN(n11538) );
  AND2_X1 U14048 ( .A1(n11876), .A2(n11541), .ZN(n11550) );
  INV_X1 U14049 ( .A(n11555), .ZN(n11553) );
  NAND2_X1 U14050 ( .A1(n11574), .A2(n11542), .ZN(n11554) );
  NAND2_X1 U14051 ( .A1(n11574), .A2(n13836), .ZN(n11543) );
  NAND4_X1 U14052 ( .A1(n11558), .A2(n11555), .A3(n11544), .A4(n11543), .ZN(
        n11545) );
  OAI21_X1 U14053 ( .B1(n11553), .B2(n11554), .A(n11545), .ZN(n11549) );
  MUX2_X1 U14054 ( .A(n11547), .B(n11546), .S(n11574), .Z(n11548) );
  OAI211_X1 U14055 ( .C1(n11551), .C2(n11550), .A(n11549), .B(n11548), .ZN(
        n11564) );
  NAND4_X1 U14056 ( .A1(n14694), .A2(n11552), .A3(n11844), .A4(n13836), .ZN(
        n11563) );
  NAND2_X1 U14057 ( .A1(n11553), .A2(n11844), .ZN(n11562) );
  INV_X1 U14058 ( .A(n11554), .ZN(n11557) );
  NAND3_X1 U14059 ( .A1(n11557), .A2(n11556), .A3(n11555), .ZN(n11561) );
  INV_X1 U14060 ( .A(n11558), .ZN(n11559) );
  NAND2_X1 U14061 ( .A1(n11559), .A2(n11574), .ZN(n11560) );
  MUX2_X1 U14062 ( .A(n13834), .B(n11565), .S(n11574), .Z(n11569) );
  NAND2_X1 U14063 ( .A1(n11568), .A2(n11569), .ZN(n11567) );
  MUX2_X1 U14064 ( .A(n11565), .B(n13834), .S(n11574), .Z(n11566) );
  NAND2_X1 U14065 ( .A1(n11567), .A2(n11566), .ZN(n11573) );
  INV_X1 U14066 ( .A(n11568), .ZN(n11571) );
  INV_X1 U14067 ( .A(n11569), .ZN(n11570) );
  NAND2_X1 U14068 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  MUX2_X1 U14069 ( .A(n13833), .B(n13743), .S(n11574), .Z(n11575) );
  MUX2_X1 U14070 ( .A(n13832), .B(n11578), .S(n11574), .Z(n11582) );
  NAND2_X1 U14071 ( .A1(n11581), .A2(n11582), .ZN(n11580) );
  MUX2_X1 U14072 ( .A(n13832), .B(n11578), .S(n11844), .Z(n11579) );
  NAND2_X1 U14073 ( .A1(n11580), .A2(n11579), .ZN(n11586) );
  INV_X1 U14074 ( .A(n11581), .ZN(n11584) );
  INV_X1 U14075 ( .A(n11582), .ZN(n11583) );
  NAND2_X1 U14076 ( .A1(n11584), .A2(n11583), .ZN(n11585) );
  MUX2_X1 U14077 ( .A(n13831), .B(n11587), .S(n11844), .Z(n11589) );
  MUX2_X1 U14078 ( .A(n13831), .B(n11587), .S(n11867), .Z(n11588) );
  MUX2_X1 U14079 ( .A(n13830), .B(n14737), .S(n11867), .Z(n11593) );
  NAND2_X1 U14080 ( .A1(n11592), .A2(n11593), .ZN(n11591) );
  MUX2_X1 U14081 ( .A(n13830), .B(n14737), .S(n11844), .Z(n11590) );
  NAND2_X1 U14082 ( .A1(n11591), .A2(n11590), .ZN(n11597) );
  INV_X1 U14083 ( .A(n11592), .ZN(n11595) );
  INV_X1 U14084 ( .A(n11593), .ZN(n11594) );
  NAND2_X1 U14085 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  MUX2_X1 U14086 ( .A(n13829), .B(n14688), .S(n11844), .Z(n11599) );
  MUX2_X1 U14087 ( .A(n13829), .B(n14688), .S(n11867), .Z(n11598) );
  INV_X1 U14088 ( .A(n11599), .ZN(n11600) );
  MUX2_X1 U14089 ( .A(n13828), .B(n14756), .S(n11867), .Z(n11604) );
  NAND2_X1 U14090 ( .A1(n11603), .A2(n11604), .ZN(n11602) );
  MUX2_X1 U14091 ( .A(n13828), .B(n14756), .S(n11844), .Z(n11601) );
  NAND2_X1 U14092 ( .A1(n11602), .A2(n11601), .ZN(n11608) );
  INV_X1 U14093 ( .A(n11603), .ZN(n11606) );
  INV_X1 U14094 ( .A(n11604), .ZN(n11605) );
  NAND2_X1 U14095 ( .A1(n11606), .A2(n11605), .ZN(n11607) );
  MUX2_X1 U14096 ( .A(n13827), .B(n11609), .S(n11844), .Z(n11611) );
  MUX2_X1 U14097 ( .A(n13827), .B(n11609), .S(n11867), .Z(n11610) );
  INV_X1 U14098 ( .A(n11611), .ZN(n11612) );
  MUX2_X1 U14099 ( .A(n13826), .B(n11613), .S(n11867), .Z(n11617) );
  NAND2_X1 U14100 ( .A1(n11616), .A2(n11617), .ZN(n11615) );
  MUX2_X1 U14101 ( .A(n13826), .B(n11613), .S(n11844), .Z(n11614) );
  INV_X1 U14102 ( .A(n11616), .ZN(n11619) );
  INV_X1 U14103 ( .A(n11617), .ZN(n11618) );
  MUX2_X1 U14104 ( .A(n13825), .B(n14469), .S(n11844), .Z(n11621) );
  MUX2_X1 U14105 ( .A(n14539), .B(n13783), .S(n11867), .Z(n11620) );
  AOI21_X1 U14106 ( .B1(n11629), .B2(n11622), .A(n11844), .ZN(n11623) );
  AOI21_X1 U14107 ( .B1(n11626), .B2(n11624), .A(n11867), .ZN(n11625) );
  AOI21_X1 U14108 ( .B1(n11627), .B2(n11626), .A(n11625), .ZN(n11628) );
  MUX2_X1 U14109 ( .A(n13972), .B(n13973), .S(n11844), .Z(n11648) );
  MUX2_X1 U14110 ( .A(n14573), .B(n14598), .S(n11867), .Z(n11630) );
  NAND2_X1 U14111 ( .A1(n11631), .A2(n11791), .ZN(n11634) );
  AOI22_X1 U14112 ( .A1(n11632), .A2(n11659), .B1(n11660), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n11633) );
  XNOR2_X1 U14113 ( .A(n14303), .B(n11844), .ZN(n11649) );
  INV_X1 U14114 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11635) );
  AND2_X1 U14115 ( .A1(n11636), .A2(n11635), .ZN(n11637) );
  OR2_X1 U14116 ( .A1(n11637), .A2(n11663), .ZN(n14168) );
  INV_X1 U14117 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14118 ( .A1(n11707), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11639) );
  INV_X1 U14119 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14169) );
  OR2_X1 U14120 ( .A1(n11820), .A2(n14169), .ZN(n11638) );
  OAI211_X1 U14121 ( .C1(n6802), .C2(n11640), .A(n11639), .B(n11638), .ZN(
        n11641) );
  INV_X1 U14122 ( .A(n11641), .ZN(n11642) );
  OAI21_X1 U14123 ( .B1(n14168), .B2(n11818), .A(n11642), .ZN(n14576) );
  XNOR2_X1 U14124 ( .A(n14576), .B(n11867), .ZN(n11650) );
  NAND2_X1 U14125 ( .A1(n11643), .A2(n11791), .ZN(n11646) );
  AOI22_X1 U14126 ( .A1(n11644), .A2(n11659), .B1(n6422), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n11645) );
  NOR2_X1 U14127 ( .A1(n13749), .A2(n13935), .ZN(n13976) );
  MUX2_X1 U14128 ( .A(n13935), .B(n13749), .S(n11844), .Z(n11651) );
  OAI22_X1 U14129 ( .A1(n11649), .A2(n11650), .B1(n13976), .B2(n11651), .ZN(
        n11647) );
  INV_X1 U14130 ( .A(n11649), .ZN(n11654) );
  NAND2_X1 U14131 ( .A1(n13749), .A2(n13935), .ZN(n13977) );
  AOI21_X1 U14132 ( .B1(n11651), .B2(n13977), .A(n11650), .ZN(n11653) );
  NAND3_X1 U14133 ( .A1(n11651), .A2(n13977), .A3(n11650), .ZN(n11652) );
  INV_X1 U14134 ( .A(n11655), .ZN(n11656) );
  NAND2_X1 U14135 ( .A1(n11657), .A2(n11656), .ZN(n11669) );
  NAND2_X1 U14136 ( .A1(n11658), .A2(n11791), .ZN(n11662) );
  AOI22_X1 U14137 ( .A1(n6422), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14184), 
        .B2(n11659), .ZN(n11661) );
  NOR2_X1 U14138 ( .A1(n11663), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11664) );
  OR2_X1 U14139 ( .A1(n11674), .A2(n11664), .ZN(n14141) );
  INV_X1 U14140 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U14141 ( .A1(n11817), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14142 ( .A1(n11830), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11665) );
  OAI211_X1 U14143 ( .C1(n11797), .C2(n15312), .A(n11666), .B(n11665), .ZN(
        n11667) );
  INV_X1 U14144 ( .A(n11667), .ZN(n11668) );
  OAI21_X1 U14145 ( .B1(n14141), .B2(n11818), .A(n11668), .ZN(n14163) );
  XNOR2_X1 U14146 ( .A(n14153), .B(n14163), .ZN(n14146) );
  NAND2_X1 U14147 ( .A1(n11669), .A2(n14146), .ZN(n11673) );
  NAND2_X1 U14148 ( .A1(n14163), .A2(n11867), .ZN(n11671) );
  OR2_X1 U14149 ( .A1(n14163), .A2(n11867), .ZN(n11670) );
  MUX2_X1 U14150 ( .A(n11671), .B(n11670), .S(n14153), .Z(n11672) );
  NAND2_X1 U14151 ( .A1(n11673), .A2(n11672), .ZN(n11685) );
  NOR2_X1 U14152 ( .A1(n11674), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11675) );
  OR2_X1 U14153 ( .A1(n11688), .A2(n11675), .ZN(n13769) );
  INV_X1 U14154 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U14155 ( .A1(n11830), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11677) );
  NAND2_X1 U14156 ( .A1(n11707), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11676) );
  OAI211_X1 U14157 ( .C1(n6802), .C2(n14253), .A(n11677), .B(n11676), .ZN(
        n11678) );
  INV_X1 U14158 ( .A(n11678), .ZN(n11679) );
  OAI21_X1 U14159 ( .B1(n13769), .B2(n11818), .A(n11679), .ZN(n14149) );
  NAND2_X1 U14160 ( .A1(n11680), .A2(n11791), .ZN(n11683) );
  OR2_X1 U14161 ( .A1(n11857), .A2(n11681), .ZN(n11682) );
  MUX2_X1 U14162 ( .A(n14149), .B(n14132), .S(n11844), .Z(n11686) );
  MUX2_X1 U14163 ( .A(n14149), .B(n14132), .S(n11867), .Z(n11684) );
  INV_X1 U14164 ( .A(n11686), .ZN(n11687) );
  NOR2_X1 U14165 ( .A1(n11688), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11689) );
  OR2_X1 U14166 ( .A1(n11704), .A2(n11689), .ZN(n14111) );
  INV_X1 U14167 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14168 ( .A1(n11830), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14169 ( .A1(n11707), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11690) );
  OAI211_X1 U14170 ( .C1(n6802), .C2(n11692), .A(n11691), .B(n11690), .ZN(
        n11693) );
  INV_X1 U14171 ( .A(n11693), .ZN(n11694) );
  OAI21_X1 U14172 ( .B1(n14111), .B2(n11818), .A(n11694), .ZN(n13983) );
  NAND2_X1 U14173 ( .A1(n11695), .A2(n11791), .ZN(n11698) );
  OR2_X1 U14174 ( .A1(n11857), .A2(n11696), .ZN(n11697) );
  MUX2_X1 U14175 ( .A(n13983), .B(n14292), .S(n11867), .Z(n11702) );
  MUX2_X1 U14176 ( .A(n13983), .B(n14292), .S(n11844), .Z(n11699) );
  NAND2_X1 U14177 ( .A1(n11700), .A2(n11699), .ZN(n11703) );
  OR2_X1 U14178 ( .A1(n11704), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11705) );
  NAND2_X1 U14179 ( .A1(n11704), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11719) );
  AND2_X1 U14180 ( .A1(n11705), .A2(n11719), .ZN(n14099) );
  NAND2_X1 U14181 ( .A1(n14099), .A2(n11706), .ZN(n11712) );
  INV_X1 U14182 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15314) );
  NAND2_X1 U14183 ( .A1(n11707), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14184 ( .A1(n11830), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11708) );
  OAI211_X1 U14185 ( .C1(n6802), .C2(n15314), .A(n11709), .B(n11708), .ZN(
        n11710) );
  INV_X1 U14186 ( .A(n11710), .ZN(n11711) );
  NAND2_X1 U14187 ( .A1(n11712), .A2(n11711), .ZN(n13985) );
  XNOR2_X1 U14188 ( .A(n11714), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U14189 ( .A1(n11817), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11724) );
  INV_X1 U14190 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11718) );
  OR2_X1 U14191 ( .A1(n11797), .A2(n11718), .ZN(n11723) );
  OAI21_X1 U14192 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11720), .A(n11735), 
        .ZN(n14085) );
  OR2_X1 U14193 ( .A1(n11818), .A2(n14085), .ZN(n11722) );
  INV_X1 U14194 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14086) );
  OR2_X1 U14195 ( .A1(n11820), .A2(n14086), .ZN(n11721) );
  NAND4_X1 U14196 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n14063) );
  NAND2_X1 U14197 ( .A1(n11725), .A2(n11791), .ZN(n11728) );
  OR2_X1 U14198 ( .A1(n11857), .A2(n11726), .ZN(n11727) );
  MUX2_X1 U14199 ( .A(n14063), .B(n14232), .S(n11867), .Z(n11732) );
  NAND2_X1 U14200 ( .A1(n11731), .A2(n11732), .ZN(n11730) );
  MUX2_X1 U14201 ( .A(n14063), .B(n14232), .S(n11844), .Z(n11729) );
  INV_X1 U14202 ( .A(n11731), .ZN(n11734) );
  INV_X1 U14203 ( .A(n11732), .ZN(n11733) );
  NAND2_X1 U14204 ( .A1(n11817), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11740) );
  INV_X1 U14205 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14286) );
  OR2_X1 U14206 ( .A1(n11797), .A2(n14286), .ZN(n11739) );
  OAI21_X1 U14207 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11736), .A(n11748), 
        .ZN(n14071) );
  OR2_X1 U14208 ( .A1(n11818), .A2(n14071), .ZN(n11738) );
  INV_X1 U14209 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14072) );
  OR2_X1 U14210 ( .A1(n11820), .A2(n14072), .ZN(n11737) );
  NAND4_X1 U14211 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n13988) );
  OR2_X1 U14212 ( .A1(n11857), .A2(n11742), .ZN(n11743) );
  MUX2_X1 U14213 ( .A(n13988), .B(n14073), .S(n11844), .Z(n11745) );
  NAND2_X1 U14214 ( .A1(n11817), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11753) );
  INV_X1 U14215 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n14282) );
  OR2_X1 U14216 ( .A1(n11797), .A2(n14282), .ZN(n11752) );
  INV_X1 U14217 ( .A(n11748), .ZN(n11746) );
  NAND2_X1 U14218 ( .A1(n11746), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11769) );
  INV_X1 U14219 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14220 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND2_X1 U14221 ( .A1(n11769), .A2(n11749), .ZN(n14055) );
  OR2_X1 U14222 ( .A1(n11818), .A2(n14055), .ZN(n11751) );
  INV_X1 U14223 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14056) );
  OR2_X1 U14224 ( .A1(n11820), .A2(n14056), .ZN(n11750) );
  NAND4_X1 U14225 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n14062) );
  NAND2_X1 U14226 ( .A1(n11754), .A2(n11791), .ZN(n11757) );
  OR2_X1 U14227 ( .A1(n11857), .A2(n11755), .ZN(n11756) );
  MUX2_X1 U14228 ( .A(n14062), .B(n14220), .S(n11867), .Z(n11761) );
  NAND2_X1 U14229 ( .A1(n11760), .A2(n11761), .ZN(n11759) );
  MUX2_X1 U14230 ( .A(n14062), .B(n14220), .S(n11844), .Z(n11758) );
  NAND2_X1 U14231 ( .A1(n11759), .A2(n11758), .ZN(n11765) );
  INV_X1 U14232 ( .A(n11760), .ZN(n11763) );
  INV_X1 U14233 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U14234 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  NAND2_X1 U14235 ( .A1(n11817), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11774) );
  INV_X1 U14236 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11766) );
  OR2_X1 U14237 ( .A1(n11797), .A2(n11766), .ZN(n11773) );
  INV_X1 U14238 ( .A(n11769), .ZN(n11767) );
  NAND2_X1 U14239 ( .A1(n11767), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11785) );
  INV_X1 U14240 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U14241 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  NAND2_X1 U14242 ( .A1(n11785), .A2(n11770), .ZN(n14031) );
  OR2_X1 U14243 ( .A1(n11818), .A2(n14031), .ZN(n11772) );
  INV_X1 U14244 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14034) );
  OR2_X1 U14245 ( .A1(n11820), .A2(n14034), .ZN(n11771) );
  NAND4_X1 U14246 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n14020) );
  NAND2_X1 U14247 ( .A1(n13685), .A2(n11791), .ZN(n11776) );
  OR2_X1 U14248 ( .A1(n11857), .A2(n14321), .ZN(n11775) );
  MUX2_X1 U14249 ( .A(n14020), .B(n14038), .S(n11844), .Z(n11779) );
  MUX2_X1 U14250 ( .A(n14020), .B(n14038), .S(n11867), .Z(n11777) );
  INV_X1 U14251 ( .A(n11778), .ZN(n11781) );
  INV_X1 U14252 ( .A(n11779), .ZN(n11780) );
  NAND2_X1 U14253 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  NAND2_X1 U14254 ( .A1(n11817), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11790) );
  INV_X1 U14255 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14275) );
  OR2_X1 U14256 ( .A1(n11797), .A2(n14275), .ZN(n11789) );
  INV_X1 U14257 ( .A(n11785), .ZN(n11783) );
  NAND2_X1 U14258 ( .A1(n11783), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11800) );
  INV_X1 U14259 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U14260 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  NAND2_X1 U14261 ( .A1(n11800), .A2(n11786), .ZN(n14023) );
  OR2_X1 U14262 ( .A1(n11818), .A2(n14023), .ZN(n11788) );
  INV_X1 U14263 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14024) );
  OR2_X1 U14264 ( .A1(n11820), .A2(n14024), .ZN(n11787) );
  NAND4_X1 U14265 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n13999) );
  OR2_X1 U14266 ( .A1(n11857), .A2(n14318), .ZN(n11792) );
  MUX2_X1 U14267 ( .A(n13999), .B(n14026), .S(n11867), .Z(n11795) );
  MUX2_X1 U14268 ( .A(n13999), .B(n14026), .S(n11844), .Z(n11794) );
  NAND2_X1 U14269 ( .A1(n11817), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11806) );
  INV_X1 U14270 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n11796) );
  OR2_X1 U14271 ( .A1(n11797), .A2(n11796), .ZN(n11805) );
  INV_X1 U14272 ( .A(n11800), .ZN(n11798) );
  NAND2_X1 U14273 ( .A1(n11798), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13969) );
  INV_X1 U14274 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14275 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  NAND2_X1 U14276 ( .A1(n13969), .A2(n11801), .ZN(n14005) );
  OR2_X1 U14277 ( .A1(n11818), .A2(n14005), .ZN(n11804) );
  INV_X1 U14278 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11802) );
  OR2_X1 U14279 ( .A1(n11820), .A2(n11802), .ZN(n11803) );
  NAND4_X1 U14280 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n14019) );
  OR2_X1 U14281 ( .A1(n11857), .A2(n14315), .ZN(n11807) );
  MUX2_X1 U14282 ( .A(n14019), .B(n14205), .S(n11844), .Z(n11812) );
  NAND2_X1 U14283 ( .A1(n11811), .A2(n11812), .ZN(n11810) );
  MUX2_X1 U14284 ( .A(n14019), .B(n14205), .S(n11867), .Z(n11809) );
  NAND2_X1 U14285 ( .A1(n11810), .A2(n11809), .ZN(n11816) );
  INV_X1 U14286 ( .A(n11811), .ZN(n11814) );
  INV_X1 U14287 ( .A(n11812), .ZN(n11813) );
  NAND2_X1 U14288 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  NAND2_X1 U14289 ( .A1(n11707), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14290 ( .A1(n11817), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11823) );
  OR2_X1 U14291 ( .A1(n11818), .A2(n13969), .ZN(n11822) );
  INV_X1 U14292 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n11819) );
  OR2_X1 U14293 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  NAND4_X1 U14294 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n13998) );
  NAND2_X1 U14295 ( .A1(n13675), .A2(n11791), .ZN(n11826) );
  OR2_X1 U14296 ( .A1(n11857), .A2(n14312), .ZN(n11825) );
  MUX2_X1 U14297 ( .A(n13998), .B(n14202), .S(n11867), .Z(n11846) );
  INV_X1 U14298 ( .A(n11827), .ZN(n11833) );
  INV_X1 U14299 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U14300 ( .A1(n11830), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11829) );
  NAND2_X1 U14301 ( .A1(n11707), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11828) );
  OAI211_X1 U14302 ( .C1(n6802), .C2(n14194), .A(n11829), .B(n11828), .ZN(
        n13925) );
  INV_X1 U14303 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14198) );
  NAND2_X1 U14304 ( .A1(n11830), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14305 ( .A1(n11707), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11831) );
  OAI211_X1 U14306 ( .C1(n6802), .C2(n14198), .A(n11832), .B(n11831), .ZN(
        n13963) );
  OAI21_X1 U14307 ( .B1(n11833), .B2(n13925), .A(n13963), .ZN(n11838) );
  NAND2_X1 U14308 ( .A1(n11834), .A2(n11791), .ZN(n11837) );
  OR2_X1 U14309 ( .A1(n11857), .A2(n11835), .ZN(n11836) );
  MUX2_X1 U14310 ( .A(n11838), .B(n14272), .S(n11844), .Z(n11852) );
  NAND2_X1 U14311 ( .A1(n11899), .A2(n11867), .ZN(n11842) );
  INV_X1 U14312 ( .A(n13925), .ZN(n11868) );
  OAI21_X1 U14313 ( .B1(n11867), .B2(n11868), .A(n11839), .ZN(n11840) );
  NAND2_X1 U14314 ( .A1(n11840), .A2(n13963), .ZN(n11841) );
  NAND2_X1 U14315 ( .A1(n11842), .A2(n11841), .ZN(n11851) );
  INV_X1 U14316 ( .A(n11843), .ZN(n11850) );
  INV_X1 U14317 ( .A(n13998), .ZN(n12137) );
  MUX2_X1 U14318 ( .A(n12137), .B(n6419), .S(n11844), .Z(n11845) );
  AOI21_X1 U14319 ( .B1(n11847), .B2(n11846), .A(n11845), .ZN(n11848) );
  INV_X1 U14320 ( .A(n11848), .ZN(n11849) );
  NAND2_X1 U14321 ( .A1(n11850), .A2(n11849), .ZN(n11856) );
  INV_X1 U14322 ( .A(n11851), .ZN(n11854) );
  INV_X1 U14323 ( .A(n11852), .ZN(n11853) );
  NAND2_X1 U14324 ( .A1(n13669), .A2(n11791), .ZN(n11859) );
  INV_X1 U14325 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14307) );
  OR2_X1 U14326 ( .A1(n11857), .A2(n14307), .ZN(n11858) );
  XNOR2_X1 U14327 ( .A(n13922), .B(n11868), .ZN(n11872) );
  NAND2_X1 U14328 ( .A1(n7533), .A2(n11860), .ZN(n11861) );
  NAND2_X1 U14329 ( .A1(n11862), .A2(n11861), .ZN(n11865) );
  OR2_X1 U14330 ( .A1(n11863), .A2(n14471), .ZN(n11864) );
  NAND2_X1 U14331 ( .A1(n11865), .A2(n11864), .ZN(n11905) );
  NAND2_X1 U14332 ( .A1(n11870), .A2(n11869), .ZN(n11903) );
  NAND2_X1 U14333 ( .A1(n11905), .A2(n11903), .ZN(n11906) );
  INV_X1 U14334 ( .A(n11872), .ZN(n11907) );
  INV_X1 U14335 ( .A(n13999), .ZN(n11873) );
  INV_X1 U14336 ( .A(n14020), .ZN(n13958) );
  XNOR2_X1 U14337 ( .A(n14038), .B(n13958), .ZN(n14039) );
  XNOR2_X1 U14338 ( .A(n14220), .B(n14062), .ZN(n13955) );
  XNOR2_X1 U14339 ( .A(n14238), .B(n13985), .ZN(n14095) );
  INV_X1 U14340 ( .A(n13983), .ZN(n13946) );
  XNOR2_X1 U14341 ( .A(n14292), .B(n13946), .ZN(n14112) );
  INV_X1 U14342 ( .A(n14149), .ZN(n13711) );
  OR2_X1 U14343 ( .A1(n14132), .A2(n13711), .ZN(n13945) );
  NAND2_X1 U14344 ( .A1(n14132), .A2(n13711), .ZN(n11874) );
  NAND2_X1 U14345 ( .A1(n13945), .A2(n11874), .ZN(n13944) );
  INV_X1 U14346 ( .A(n13976), .ZN(n11875) );
  NAND2_X1 U14347 ( .A1(n11875), .A2(n13977), .ZN(n14583) );
  NAND4_X1 U14348 ( .A1(n14694), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11879) );
  NOR4_X1 U14349 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11885) );
  NAND4_X1 U14350 ( .A1(n14677), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11886) );
  NOR3_X1 U14351 ( .A1(n11887), .A2(n7146), .A3(n11886), .ZN(n11890) );
  NAND4_X1 U14352 ( .A1(n14583), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11894) );
  NOR4_X1 U14353 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11895) );
  XNOR2_X1 U14354 ( .A(n14303), .B(n14576), .ZN(n14160) );
  NAND3_X1 U14355 ( .A1(n14146), .A2(n11895), .A3(n14160), .ZN(n11896) );
  NOR4_X1 U14356 ( .A1(n14095), .A2(n14112), .A3(n13944), .A4(n11896), .ZN(
        n11897) );
  XNOR2_X1 U14357 ( .A(n14073), .B(n13988), .ZN(n14065) );
  XNOR2_X1 U14358 ( .A(n14232), .B(n14063), .ZN(n14081) );
  NAND4_X1 U14359 ( .A1(n13955), .A2(n11897), .A3(n14065), .A4(n14081), .ZN(
        n11898) );
  NOR4_X1 U14360 ( .A1(n14009), .A2(n14018), .A3(n14039), .A4(n11898), .ZN(
        n11901) );
  XNOR2_X1 U14361 ( .A(n11899), .B(n13963), .ZN(n11900) );
  NAND4_X1 U14362 ( .A1(n11907), .A2(n11901), .A3(n11900), .A4(n13992), .ZN(
        n11902) );
  XNOR2_X1 U14363 ( .A(n11902), .B(n14471), .ZN(n11904) );
  NOR2_X1 U14364 ( .A1(n11904), .A2(n11903), .ZN(n11912) );
  INV_X1 U14365 ( .A(n11905), .ZN(n11910) );
  NOR2_X1 U14366 ( .A1(n11907), .A2(n11906), .ZN(n11909) );
  NAND2_X1 U14367 ( .A1(n11914), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11915) );
  OAI21_X1 U14368 ( .B1(n11918), .B2(n6831), .A(P1_B_REG_SCAN_IN), .ZN(n11917)
         );
  INV_X1 U14369 ( .A(n11919), .ZN(n11920) );
  NAND2_X1 U14370 ( .A1(n11923), .A2(n11922), .ZN(n14530) );
  INV_X1 U14371 ( .A(n14530), .ZN(n11925) );
  INV_X1 U14372 ( .A(n14536), .ZN(n13299) );
  XNOR2_X1 U14373 ( .A(n13299), .B(n11972), .ZN(n13066) );
  NAND2_X1 U14374 ( .A1(n13130), .A2(n13529), .ZN(n11926) );
  XNOR2_X1 U14375 ( .A(n13066), .B(n11926), .ZN(n14529) );
  NAND2_X1 U14376 ( .A1(n13066), .A2(n11926), .ZN(n11927) );
  XNOR2_X1 U14377 ( .A(n13628), .B(n11101), .ZN(n11928) );
  NAND2_X1 U14378 ( .A1(n13129), .A2(n13529), .ZN(n11929) );
  XNOR2_X1 U14379 ( .A(n11928), .B(n11929), .ZN(n13068) );
  INV_X1 U14380 ( .A(n11928), .ZN(n11931) );
  INV_X1 U14381 ( .A(n11929), .ZN(n11930) );
  XNOR2_X1 U14382 ( .A(n13623), .B(n11101), .ZN(n13031) );
  NAND2_X1 U14383 ( .A1(n13128), .A2(n13529), .ZN(n11932) );
  NOR2_X1 U14384 ( .A1(n13031), .A2(n11932), .ZN(n11933) );
  AOI21_X1 U14385 ( .B1(n13031), .B2(n11932), .A(n11933), .ZN(n13103) );
  XNOR2_X1 U14386 ( .A(n13618), .B(n11972), .ZN(n13087) );
  NAND2_X1 U14387 ( .A1(n13127), .A2(n13529), .ZN(n11936) );
  XNOR2_X1 U14388 ( .A(n13087), .B(n11936), .ZN(n13038) );
  INV_X1 U14389 ( .A(n11933), .ZN(n11934) );
  INV_X1 U14390 ( .A(n11936), .ZN(n11937) );
  XNOR2_X1 U14391 ( .A(n13449), .B(n11972), .ZN(n11942) );
  NAND2_X1 U14392 ( .A1(n13309), .A2(n13529), .ZN(n11940) );
  XNOR2_X1 U14393 ( .A(n11942), .B(n11940), .ZN(n13088) );
  INV_X1 U14394 ( .A(n11940), .ZN(n11941) );
  XNOR2_X1 U14395 ( .A(n13604), .B(n11972), .ZN(n11945) );
  NAND2_X1 U14396 ( .A1(n13126), .A2(n13529), .ZN(n11946) );
  XNOR2_X1 U14397 ( .A(n11945), .B(n11946), .ZN(n13045) );
  INV_X1 U14398 ( .A(n13045), .ZN(n11944) );
  INV_X1 U14399 ( .A(n11945), .ZN(n11948) );
  INV_X1 U14400 ( .A(n11946), .ZN(n11947) );
  NAND2_X1 U14401 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  NAND2_X1 U14402 ( .A1(n13042), .A2(n11949), .ZN(n11951) );
  XNOR2_X1 U14403 ( .A(n13598), .B(n11972), .ZN(n11950) );
  NAND2_X1 U14404 ( .A1(n11951), .A2(n11950), .ZN(n11953) );
  OR2_X1 U14405 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  NAND2_X1 U14406 ( .A1(n11953), .A2(n11952), .ZN(n13095) );
  XNOR2_X1 U14407 ( .A(n13410), .B(n11101), .ZN(n11954) );
  NAND2_X1 U14408 ( .A1(n13281), .A2(n13529), .ZN(n13010) );
  INV_X1 U14409 ( .A(n11954), .ZN(n11955) );
  XNOR2_X1 U14410 ( .A(n13587), .B(n11972), .ZN(n11956) );
  AND2_X1 U14411 ( .A1(n13314), .A2(n13529), .ZN(n11957) );
  NAND2_X1 U14412 ( .A1(n11956), .A2(n11957), .ZN(n11960) );
  INV_X1 U14413 ( .A(n11956), .ZN(n13052) );
  INV_X1 U14414 ( .A(n11957), .ZN(n11958) );
  NAND2_X1 U14415 ( .A1(n13052), .A2(n11958), .ZN(n11959) );
  NAND2_X1 U14416 ( .A1(n13049), .A2(n11960), .ZN(n11965) );
  XNOR2_X1 U14417 ( .A(n6879), .B(n11972), .ZN(n11961) );
  AND2_X1 U14418 ( .A1(n13316), .A2(n13529), .ZN(n11962) );
  NAND2_X1 U14419 ( .A1(n11961), .A2(n11962), .ZN(n11966) );
  INV_X1 U14420 ( .A(n11961), .ZN(n13111) );
  INV_X1 U14421 ( .A(n11962), .ZN(n11963) );
  NAND2_X1 U14422 ( .A1(n13111), .A2(n11963), .ZN(n11964) );
  NAND2_X1 U14423 ( .A1(n11965), .A2(n13050), .ZN(n13053) );
  XNOR2_X1 U14424 ( .A(n13373), .B(n11972), .ZN(n11970) );
  NAND2_X1 U14425 ( .A1(n13318), .A2(n13529), .ZN(n11968) );
  XNOR2_X1 U14426 ( .A(n11970), .B(n11968), .ZN(n13112) );
  INV_X1 U14427 ( .A(n11968), .ZN(n11969) );
  XNOR2_X1 U14428 ( .A(n13568), .B(n11972), .ZN(n11974) );
  AND2_X1 U14429 ( .A1(n13286), .A2(n13529), .ZN(n11973) );
  NAND2_X1 U14430 ( .A1(n11974), .A2(n11973), .ZN(n11975) );
  OAI21_X1 U14431 ( .B1(n11974), .B2(n11973), .A(n11975), .ZN(n13001) );
  NAND2_X1 U14432 ( .A1(n13006), .A2(n11975), .ZN(n11980) );
  NAND2_X1 U14433 ( .A1(n13124), .A2(n13529), .ZN(n11977) );
  XNOR2_X1 U14434 ( .A(n11977), .B(n11976), .ZN(n11978) );
  XNOR2_X1 U14435 ( .A(n13558), .B(n11978), .ZN(n11979) );
  XNOR2_X1 U14436 ( .A(n11980), .B(n11979), .ZN(n11986) );
  NAND2_X1 U14437 ( .A1(n13123), .A2(n13254), .ZN(n11982) );
  NAND2_X1 U14438 ( .A1(n13286), .A2(n13116), .ZN(n11981) );
  NAND2_X1 U14439 ( .A1(n11982), .A2(n11981), .ZN(n13337) );
  AOI22_X1 U14440 ( .A1(n14534), .A2(n13337), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11983) );
  OAI21_X1 U14441 ( .B1(n14797), .B2(n13345), .A(n11983), .ZN(n11984) );
  AOI21_X1 U14442 ( .B1(n13558), .B2(n14782), .A(n11984), .ZN(n11985) );
  OAI21_X1 U14443 ( .B1(n11986), .B2(n14777), .A(n11985), .ZN(P2_U3192) );
  INV_X1 U14444 ( .A(n14797), .ZN(n13058) );
  INV_X1 U14445 ( .A(n11987), .ZN(n11996) );
  NAND2_X1 U14446 ( .A1(n14782), .A2(n15001), .ZN(n11988) );
  NAND2_X1 U14447 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14829) );
  OAI211_X1 U14448 ( .C1(n14787), .C2(n11989), .A(n11988), .B(n14829), .ZN(
        n11995) );
  AOI22_X1 U14449 ( .A1(n13096), .A2(n13142), .B1(n14788), .B2(n11990), .ZN(
        n11992) );
  NOR3_X1 U14450 ( .A1(n11993), .A2(n11992), .A3(n11991), .ZN(n11994) );
  AOI211_X1 U14451 ( .C1(n13058), .C2(n11996), .A(n11995), .B(n11994), .ZN(
        n11997) );
  OAI21_X1 U14452 ( .B1(n11998), .B2(n14777), .A(n11997), .ZN(P2_U3199) );
  INV_X1 U14453 ( .A(n12001), .ZN(n12003) );
  OAI222_X1 U14454 ( .A1(n14451), .A2(n12003), .B1(n12997), .B2(n12002), .C1(
        P3_U3151), .C2(n12675), .ZN(P3_U3268) );
  XNOR2_X1 U14455 ( .A(n12703), .B(n12006), .ZN(n12007) );
  AOI22_X1 U14456 ( .A1(n12705), .A2(n12281), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12009) );
  NAND2_X1 U14457 ( .A1(n12698), .A2(n12282), .ZN(n12008) );
  OAI211_X1 U14458 ( .C1(n12726), .C2(n12285), .A(n12009), .B(n12008), .ZN(
        n12010) );
  AOI21_X1 U14459 ( .B1(n12011), .B2(n12287), .A(n12010), .ZN(n12012) );
  OAI21_X1 U14460 ( .B1(n12013), .B2(n12289), .A(n12012), .ZN(P3_U3160) );
  OAI222_X1 U14461 ( .A1(n14451), .A2(n12016), .B1(n12997), .B2(n12015), .C1(
        P3_U3151), .C2(n12014), .ZN(P3_U3275) );
  INV_X1 U14462 ( .A(n12017), .ZN(n12019) );
  OAI22_X1 U14463 ( .A1(n13783), .A2(n9563), .B1(n14539), .B2(n12047), .ZN(
        n12021) );
  XNOR2_X1 U14464 ( .A(n12021), .B(n12130), .ZN(n12028) );
  NOR2_X1 U14465 ( .A1(n10184), .A2(n14539), .ZN(n12022) );
  AOI21_X1 U14466 ( .B1(n14469), .B2(n12122), .A(n12022), .ZN(n12029) );
  XNOR2_X1 U14467 ( .A(n12028), .B(n12029), .ZN(n13775) );
  NAND2_X1 U14468 ( .A1(n14606), .A2(n12129), .ZN(n12024) );
  NAND2_X1 U14469 ( .A1(n12122), .A2(n13824), .ZN(n12023) );
  NAND2_X1 U14470 ( .A1(n12024), .A2(n12023), .ZN(n12025) );
  XNOR2_X1 U14471 ( .A(n12025), .B(n12130), .ZN(n12032) );
  NOR2_X1 U14472 ( .A1(n10184), .A2(n12026), .ZN(n12027) );
  AOI21_X1 U14473 ( .B1(n14606), .B2(n12122), .A(n12027), .ZN(n12033) );
  XNOR2_X1 U14474 ( .A(n12032), .B(n12033), .ZN(n14540) );
  INV_X1 U14475 ( .A(n12028), .ZN(n12030) );
  OR2_X1 U14476 ( .A1(n12030), .A2(n12029), .ZN(n14541) );
  INV_X1 U14477 ( .A(n12032), .ZN(n12034) );
  NAND2_X1 U14478 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  NAND2_X1 U14479 ( .A1(n12036), .A2(n12129), .ZN(n12038) );
  NAND2_X1 U14480 ( .A1(n12122), .A2(n13823), .ZN(n12037) );
  NAND2_X1 U14481 ( .A1(n12038), .A2(n12037), .ZN(n12040) );
  XNOR2_X1 U14482 ( .A(n12040), .B(n12039), .ZN(n12044) );
  NOR2_X1 U14483 ( .A1(n12046), .A2(n12044), .ZN(n14557) );
  OAI22_X1 U14484 ( .A1(n13973), .A2(n9563), .B1(n13972), .B2(n12047), .ZN(
        n12041) );
  XNOR2_X1 U14485 ( .A(n12041), .B(n12130), .ZN(n12049) );
  OR2_X1 U14486 ( .A1(n13973), .A2(n12047), .ZN(n12043) );
  NAND2_X1 U14487 ( .A1(n9562), .A2(n14573), .ZN(n12042) );
  NAND2_X1 U14488 ( .A1(n12043), .A2(n12042), .ZN(n12050) );
  XNOR2_X1 U14489 ( .A(n12049), .B(n12050), .ZN(n14556) );
  NOR2_X1 U14490 ( .A1(n14557), .A2(n14556), .ZN(n12048) );
  INV_X1 U14491 ( .A(n12044), .ZN(n12045) );
  OAI22_X1 U14492 ( .A1(n13822), .A2(n12047), .B1(n14553), .B2(n10184), .ZN(
        n13811) );
  INV_X1 U14493 ( .A(n12049), .ZN(n12052) );
  INV_X1 U14494 ( .A(n12050), .ZN(n12051) );
  NAND2_X1 U14495 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  NAND2_X1 U14496 ( .A1(n13749), .A2(n12129), .ZN(n12055) );
  NAND2_X1 U14497 ( .A1(n13935), .A2(n12122), .ZN(n12054) );
  NAND2_X1 U14498 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  XNOR2_X1 U14499 ( .A(n12056), .B(n12130), .ZN(n12057) );
  AOI22_X1 U14500 ( .A1(n13749), .A2(n12122), .B1(n9562), .B2(n13935), .ZN(
        n12058) );
  XNOR2_X1 U14501 ( .A(n12057), .B(n12058), .ZN(n13752) );
  INV_X1 U14502 ( .A(n12057), .ZN(n12059) );
  NAND2_X1 U14503 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  NAND2_X1 U14504 ( .A1(n14303), .A2(n12129), .ZN(n12062) );
  NAND2_X1 U14505 ( .A1(n14576), .A2(n12122), .ZN(n12061) );
  NAND2_X1 U14506 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  XNOR2_X1 U14507 ( .A(n12063), .B(n12130), .ZN(n12064) );
  AOI22_X1 U14508 ( .A1(n14303), .A2(n12122), .B1(n9562), .B2(n14576), .ZN(
        n12065) );
  XNOR2_X1 U14509 ( .A(n12064), .B(n12065), .ZN(n13792) );
  INV_X1 U14510 ( .A(n12064), .ZN(n12066) );
  AND2_X1 U14511 ( .A1(n14163), .A2(n9562), .ZN(n12067) );
  AOI21_X1 U14512 ( .B1(n14153), .B2(n12122), .A(n12067), .ZN(n12071) );
  NAND2_X1 U14513 ( .A1(n14153), .A2(n12129), .ZN(n12069) );
  NAND2_X1 U14514 ( .A1(n14163), .A2(n12122), .ZN(n12068) );
  NAND2_X1 U14515 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  XNOR2_X1 U14516 ( .A(n12070), .B(n12130), .ZN(n12073) );
  XOR2_X1 U14517 ( .A(n12071), .B(n12073), .Z(n13706) );
  INV_X1 U14518 ( .A(n12071), .ZN(n12072) );
  NAND2_X1 U14519 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  AND2_X1 U14520 ( .A1(n14149), .A2(n9562), .ZN(n12075) );
  AOI21_X1 U14521 ( .B1(n14132), .B2(n12122), .A(n12075), .ZN(n12078) );
  AOI22_X1 U14522 ( .A1(n14132), .A2(n12129), .B1(n12122), .B2(n14149), .ZN(
        n12076) );
  XNOR2_X1 U14523 ( .A(n12076), .B(n12130), .ZN(n12077) );
  XOR2_X1 U14524 ( .A(n12078), .B(n12077), .Z(n13767) );
  INV_X1 U14525 ( .A(n12077), .ZN(n12080) );
  INV_X1 U14526 ( .A(n12078), .ZN(n12079) );
  NAND2_X1 U14527 ( .A1(n12080), .A2(n12079), .ZN(n12081) );
  AOI22_X1 U14528 ( .A1(n14292), .A2(n12129), .B1(n12122), .B2(n13983), .ZN(
        n12082) );
  XNOR2_X1 U14529 ( .A(n12082), .B(n12130), .ZN(n12085) );
  AOI22_X1 U14530 ( .A1(n14292), .A2(n12122), .B1(n9562), .B2(n13983), .ZN(
        n12084) );
  XNOR2_X1 U14531 ( .A(n12085), .B(n12084), .ZN(n13719) );
  NAND2_X1 U14532 ( .A1(n12085), .A2(n12084), .ZN(n12086) );
  NAND2_X1 U14533 ( .A1(n13986), .A2(n12129), .ZN(n12088) );
  NAND2_X1 U14534 ( .A1(n13985), .A2(n12122), .ZN(n12087) );
  NAND2_X1 U14535 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  XNOR2_X1 U14536 ( .A(n12089), .B(n12130), .ZN(n12090) );
  AOI22_X1 U14537 ( .A1(n13986), .A2(n12122), .B1(n9562), .B2(n13985), .ZN(
        n12091) );
  XNOR2_X1 U14538 ( .A(n12090), .B(n12091), .ZN(n13786) );
  INV_X1 U14539 ( .A(n12090), .ZN(n12092) );
  NAND2_X1 U14540 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  NAND2_X1 U14541 ( .A1(n14232), .A2(n12129), .ZN(n12095) );
  NAND2_X1 U14542 ( .A1(n12122), .A2(n14063), .ZN(n12094) );
  NAND2_X1 U14543 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  XNOR2_X1 U14544 ( .A(n12096), .B(n12130), .ZN(n12097) );
  AOI22_X1 U14545 ( .A1(n14232), .A2(n12122), .B1(n9562), .B2(n14063), .ZN(
        n12098) );
  XNOR2_X1 U14546 ( .A(n12097), .B(n12098), .ZN(n13699) );
  INV_X1 U14547 ( .A(n12097), .ZN(n12099) );
  NAND2_X1 U14548 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U14549 ( .A1(n14073), .A2(n12129), .ZN(n12103) );
  NAND2_X1 U14550 ( .A1(n12122), .A2(n13988), .ZN(n12102) );
  NAND2_X1 U14551 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  XNOR2_X1 U14552 ( .A(n12104), .B(n12130), .ZN(n12105) );
  AOI22_X1 U14553 ( .A1(n14073), .A2(n12122), .B1(n9562), .B2(n13988), .ZN(
        n12106) );
  XNOR2_X1 U14554 ( .A(n12105), .B(n12106), .ZN(n13760) );
  INV_X1 U14555 ( .A(n12105), .ZN(n12107) );
  NAND2_X1 U14556 ( .A1(n12107), .A2(n12106), .ZN(n12108) );
  NAND2_X1 U14557 ( .A1(n14220), .A2(n12129), .ZN(n12110) );
  NAND2_X1 U14558 ( .A1(n12122), .A2(n14062), .ZN(n12109) );
  NAND2_X1 U14559 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  XNOR2_X1 U14560 ( .A(n12111), .B(n12130), .ZN(n12112) );
  AOI22_X1 U14561 ( .A1(n14220), .A2(n12122), .B1(n9562), .B2(n14062), .ZN(
        n12113) );
  XNOR2_X1 U14562 ( .A(n12112), .B(n12113), .ZN(n13727) );
  INV_X1 U14563 ( .A(n12112), .ZN(n12114) );
  NAND2_X1 U14564 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U14565 ( .A1(n14038), .A2(n12129), .ZN(n12117) );
  NAND2_X1 U14566 ( .A1(n12122), .A2(n14020), .ZN(n12116) );
  NAND2_X1 U14567 ( .A1(n12117), .A2(n12116), .ZN(n12118) );
  XNOR2_X1 U14568 ( .A(n12118), .B(n12130), .ZN(n12119) );
  AOI22_X1 U14569 ( .A1(n14038), .A2(n12122), .B1(n9562), .B2(n14020), .ZN(
        n12120) );
  XNOR2_X1 U14570 ( .A(n12119), .B(n12120), .ZN(n13802) );
  INV_X1 U14571 ( .A(n12119), .ZN(n12121) );
  NAND2_X1 U14572 ( .A1(n14026), .A2(n12129), .ZN(n12124) );
  NAND2_X1 U14573 ( .A1(n12122), .A2(n13999), .ZN(n12123) );
  NAND2_X1 U14574 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  XNOR2_X1 U14575 ( .A(n12125), .B(n12130), .ZN(n12126) );
  AOI22_X1 U14576 ( .A1(n14026), .A2(n12122), .B1(n9562), .B2(n13999), .ZN(
        n12127) );
  XNOR2_X1 U14577 ( .A(n12126), .B(n12127), .ZN(n13692) );
  INV_X1 U14578 ( .A(n12126), .ZN(n12128) );
  AOI22_X1 U14579 ( .A1(n14205), .A2(n12129), .B1(n12122), .B2(n14019), .ZN(
        n12133) );
  AOI22_X1 U14580 ( .A1(n14205), .A2(n12122), .B1(n9562), .B2(n14019), .ZN(
        n12131) );
  XNOR2_X1 U14581 ( .A(n12131), .B(n12130), .ZN(n12132) );
  XOR2_X1 U14582 ( .A(n12133), .B(n12132), .Z(n12134) );
  XNOR2_X1 U14583 ( .A(n12135), .B(n12134), .ZN(n12141) );
  NOR2_X1 U14584 ( .A1(n14568), .A2(n14005), .ZN(n12139) );
  AOI22_X1 U14585 ( .A1(n13794), .A2(n13999), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12136) );
  OAI21_X1 U14586 ( .B1(n12137), .B2(n14551), .A(n12136), .ZN(n12138) );
  AOI211_X1 U14587 ( .C1(n14205), .C2(n14564), .A(n12139), .B(n12138), .ZN(
        n12140) );
  OAI21_X1 U14588 ( .B1(n12141), .B2(n14559), .A(n12140), .ZN(P1_U3220) );
  INV_X1 U14589 ( .A(n12142), .ZN(n12146) );
  AOI22_X1 U14590 ( .A1(n12688), .A2(n12881), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15156), .ZN(n12143) );
  OAI21_X1 U14591 ( .B1(n12144), .B2(n12883), .A(n12143), .ZN(n12145) );
  AOI21_X1 U14592 ( .B1(n12146), .B2(n12885), .A(n12145), .ZN(n12147) );
  OAI21_X1 U14593 ( .B1(n12148), .B2(n15156), .A(n12147), .ZN(P3_U3204) );
  AOI21_X1 U14594 ( .B1(n12510), .B2(n12149), .A(n6432), .ZN(n12156) );
  INV_X1 U14595 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12150) );
  OAI22_X1 U14596 ( .A1(n8007), .A2(n12285), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12150), .ZN(n12154) );
  INV_X1 U14597 ( .A(n12773), .ZN(n12151) );
  OAI22_X1 U14598 ( .A1(n12152), .A2(n12191), .B1(n12151), .B2(n12226), .ZN(
        n12153) );
  AOI211_X1 U14599 ( .C1(n12330), .C2(n12287), .A(n12154), .B(n12153), .ZN(
        n12155) );
  OAI21_X1 U14600 ( .B1(n12156), .B2(n12289), .A(n12155), .ZN(P3_U3156) );
  XNOR2_X1 U14601 ( .A(n12159), .B(n12158), .ZN(n12164) );
  NAND2_X1 U14602 ( .A1(n12224), .A2(n12840), .ZN(n12160) );
  NAND2_X1 U14603 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12678)
         );
  OAI211_X1 U14604 ( .C1(n12816), .C2(n12191), .A(n12160), .B(n12678), .ZN(
        n12162) );
  NOR2_X1 U14605 ( .A1(n12977), .A2(n12278), .ZN(n12161) );
  AOI211_X1 U14606 ( .C1(n12819), .C2(n12281), .A(n12162), .B(n12161), .ZN(
        n12163) );
  OAI21_X1 U14607 ( .B1(n12164), .B2(n12289), .A(n12163), .ZN(P3_U3159) );
  INV_X1 U14608 ( .A(n12453), .ZN(n12969) );
  INV_X1 U14609 ( .A(n12166), .ZN(n12232) );
  INV_X1 U14610 ( .A(n12167), .ZN(n12169) );
  NOR3_X1 U14611 ( .A1(n12232), .A2(n12169), .A3(n12168), .ZN(n12172) );
  INV_X1 U14612 ( .A(n12170), .ZN(n12171) );
  OAI21_X1 U14613 ( .B1(n12172), .B2(n12171), .A(n12272), .ZN(n12176) );
  AOI22_X1 U14614 ( .A1(n12768), .A2(n12282), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12173) );
  OAI21_X1 U14615 ( .B1(n12816), .B2(n12285), .A(n12173), .ZN(n12174) );
  AOI21_X1 U14616 ( .B1(n12793), .B2(n12281), .A(n12174), .ZN(n12175) );
  OAI211_X1 U14617 ( .C1(n12969), .C2(n12278), .A(n12176), .B(n12175), .ZN(
        P3_U3163) );
  NAND2_X1 U14618 ( .A1(n12281), .A2(n12177), .ZN(n12180) );
  INV_X1 U14619 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12178) );
  NOR2_X1 U14620 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12178), .ZN(n15129) );
  AOI21_X1 U14621 ( .B1(n12282), .B2(n12512), .A(n15129), .ZN(n12179) );
  OAI211_X1 U14622 ( .C1(n12181), .C2(n12285), .A(n12180), .B(n12179), .ZN(
        n12187) );
  XNOR2_X1 U14623 ( .A(n12182), .B(n12513), .ZN(n12183) );
  XNOR2_X1 U14624 ( .A(n12184), .B(n12183), .ZN(n12185) );
  NOR2_X1 U14625 ( .A1(n12185), .A2(n12289), .ZN(n12186) );
  AOI211_X1 U14626 ( .C1(n14512), .C2(n12287), .A(n12187), .B(n12186), .ZN(
        n12188) );
  INV_X1 U14627 ( .A(n12188), .ZN(P3_U3164) );
  AOI22_X1 U14628 ( .A1(n8195), .A2(n12224), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12190) );
  NAND2_X1 U14629 ( .A1(n12742), .A2(n12281), .ZN(n12189) );
  OAI211_X1 U14630 ( .C1(n12714), .C2(n12191), .A(n12190), .B(n12189), .ZN(
        n12199) );
  INV_X1 U14631 ( .A(n12193), .ZN(n12194) );
  NAND3_X1 U14632 ( .A1(n12192), .A2(n12195), .A3(n12194), .ZN(n12196) );
  AOI21_X1 U14633 ( .B1(n12197), .B2(n12196), .A(n12289), .ZN(n12198) );
  AOI211_X1 U14634 ( .C1(n12900), .C2(n12287), .A(n12199), .B(n12198), .ZN(
        n12200) );
  INV_X1 U14635 ( .A(n12200), .ZN(P3_U3165) );
  XNOR2_X1 U14636 ( .A(n12201), .B(n12202), .ZN(n12209) );
  NAND2_X1 U14637 ( .A1(n12281), .A2(n12864), .ZN(n12205) );
  NOR2_X1 U14638 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12203), .ZN(n12594) );
  AOI21_X1 U14639 ( .B1(n12282), .B2(n12856), .A(n12594), .ZN(n12204) );
  OAI211_X1 U14640 ( .C1(n12206), .C2(n12285), .A(n12205), .B(n12204), .ZN(
        n12207) );
  AOI21_X1 U14641 ( .B1(n12938), .B2(n12287), .A(n12207), .ZN(n12208) );
  OAI21_X1 U14642 ( .B1(n12209), .B2(n12289), .A(n12208), .ZN(P3_U3166) );
  INV_X1 U14643 ( .A(n12211), .ZN(n12212) );
  AOI21_X1 U14644 ( .B1(n12213), .B2(n12210), .A(n12212), .ZN(n12218) );
  NAND2_X1 U14645 ( .A1(n12281), .A2(n12846), .ZN(n12215) );
  AND2_X1 U14646 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12620) );
  AOI21_X1 U14647 ( .B1(n12282), .B2(n12840), .A(n12620), .ZN(n12214) );
  OAI211_X1 U14648 ( .C1(n12872), .C2(n12285), .A(n12215), .B(n12214), .ZN(
        n12216) );
  AOI21_X1 U14649 ( .B1(n12934), .B2(n12287), .A(n12216), .ZN(n12217) );
  OAI21_X1 U14650 ( .B1(n12218), .B2(n12289), .A(n12217), .ZN(P3_U3168) );
  INV_X1 U14651 ( .A(n12219), .ZN(n12221) );
  NOR3_X1 U14652 ( .A1(n6432), .A2(n12221), .A3(n12220), .ZN(n12223) );
  INV_X1 U14653 ( .A(n12192), .ZN(n12222) );
  OAI21_X1 U14654 ( .B1(n12223), .B2(n12222), .A(n12272), .ZN(n12230) );
  INV_X1 U14655 ( .A(n12757), .ZN(n12227) );
  AOI22_X1 U14656 ( .A1(n12510), .A2(n12224), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12225) );
  OAI21_X1 U14657 ( .B1(n12227), .B2(n12226), .A(n12225), .ZN(n12228) );
  AOI21_X1 U14658 ( .B1(n12509), .B2(n12282), .A(n12228), .ZN(n12229) );
  OAI211_X1 U14659 ( .C1(n12759), .C2(n12278), .A(n12230), .B(n12229), .ZN(
        P3_U3169) );
  AOI21_X1 U14660 ( .B1(n12233), .B2(n12231), .A(n12232), .ZN(n12239) );
  NAND2_X1 U14661 ( .A1(n12281), .A2(n12808), .ZN(n12235) );
  AOI22_X1 U14662 ( .A1(n12282), .A2(n12801), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12234) );
  OAI211_X1 U14663 ( .C1(n12828), .C2(n12285), .A(n12235), .B(n12234), .ZN(
        n12236) );
  AOI21_X1 U14664 ( .B1(n12237), .B2(n12287), .A(n12236), .ZN(n12238) );
  OAI21_X1 U14665 ( .B1(n12239), .B2(n12289), .A(n12238), .ZN(P3_U3173) );
  XOR2_X1 U14666 ( .A(n12241), .B(n12240), .Z(n12249) );
  NOR2_X1 U14667 ( .A1(n12278), .A2(n14504), .ZN(n12248) );
  NAND2_X1 U14668 ( .A1(n12281), .A2(n12242), .ZN(n12245) );
  AOI21_X1 U14669 ( .B1(n12282), .B2(n12511), .A(n12243), .ZN(n12244) );
  OAI211_X1 U14670 ( .C1(n12246), .C2(n12285), .A(n12245), .B(n12244), .ZN(
        n12247) );
  AOI211_X1 U14671 ( .C1(n12249), .C2(n12272), .A(n12248), .B(n12247), .ZN(
        n12250) );
  INV_X1 U14672 ( .A(n12250), .ZN(P3_U3174) );
  INV_X1 U14673 ( .A(n12251), .ZN(n12252) );
  AOI21_X1 U14674 ( .B1(n12768), .B2(n12253), .A(n12252), .ZN(n12259) );
  AOI22_X1 U14675 ( .A1(n12510), .A2(n12282), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12255) );
  NAND2_X1 U14676 ( .A1(n12281), .A2(n12784), .ZN(n12254) );
  OAI211_X1 U14677 ( .C1(n12781), .C2(n12285), .A(n12255), .B(n12254), .ZN(
        n12256) );
  AOI21_X1 U14678 ( .B1(n12257), .B2(n12287), .A(n12256), .ZN(n12258) );
  OAI21_X1 U14679 ( .B1(n12259), .B2(n12289), .A(n12258), .ZN(P3_U3175) );
  AOI21_X1 U14680 ( .B1(n12261), .B2(n12260), .A(n12289), .ZN(n12263) );
  NAND2_X1 U14681 ( .A1(n12263), .A2(n12262), .ZN(n12268) );
  INV_X1 U14682 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n12264) );
  NOR2_X1 U14683 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12264), .ZN(n12657) );
  AOI21_X1 U14684 ( .B1(n12282), .B2(n12800), .A(n12657), .ZN(n12265) );
  OAI21_X1 U14685 ( .B1(n12285), .B2(n12829), .A(n12265), .ZN(n12266) );
  AOI21_X1 U14686 ( .B1(n12831), .B2(n12281), .A(n12266), .ZN(n12267) );
  OAI211_X1 U14687 ( .C1(n12982), .C2(n12278), .A(n12268), .B(n12267), .ZN(
        P3_U3178) );
  OAI21_X1 U14688 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12273) );
  NAND2_X1 U14689 ( .A1(n12273), .A2(n12272), .ZN(n12277) );
  AOI22_X1 U14690 ( .A1(n12729), .A2(n12281), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12274) );
  OAI21_X1 U14691 ( .B1(n12749), .B2(n12285), .A(n12274), .ZN(n12275) );
  AOI21_X1 U14692 ( .B1(n12697), .B2(n12282), .A(n12275), .ZN(n12276) );
  OAI211_X1 U14693 ( .C1(n12955), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        P3_U3180) );
  XNOR2_X1 U14694 ( .A(n12279), .B(n12280), .ZN(n12290) );
  NAND2_X1 U14695 ( .A1(n12281), .A2(n12880), .ZN(n12284) );
  AND2_X1 U14696 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12552) );
  AOI21_X1 U14697 ( .B1(n12282), .B2(n12839), .A(n12552), .ZN(n12283) );
  OAI211_X1 U14698 ( .C1(n12874), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12286) );
  AOI21_X1 U14699 ( .B1(n12879), .B2(n12287), .A(n12286), .ZN(n12288) );
  OAI21_X1 U14700 ( .B1(n12290), .B2(n12289), .A(n12288), .ZN(P3_U3181) );
  XNOR2_X1 U14701 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12293) );
  INV_X1 U14702 ( .A(SI_31_), .ZN(n12993) );
  OR2_X1 U14703 ( .A1(n12299), .A2(n12993), .ZN(n12295) );
  OR2_X1 U14704 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  INV_X1 U14705 ( .A(n12301), .ZN(n12507) );
  NAND2_X1 U14706 ( .A1(n12302), .A2(n12301), .ZN(n12303) );
  NAND2_X1 U14707 ( .A1(n12460), .A2(n12461), .ZN(n12782) );
  INV_X1 U14708 ( .A(n12782), .ZN(n12778) );
  INV_X1 U14709 ( .A(n12804), .ZN(n12320) );
  NAND4_X1 U14710 ( .A1(n12306), .A2(n12305), .A3(n12345), .A4(n12304), .ZN(
        n12309) );
  NAND4_X1 U14711 ( .A1(n15138), .A2(n12307), .A3(n12373), .A4(n12366), .ZN(
        n12308) );
  NOR3_X1 U14712 ( .A1(n12309), .A2(n12308), .A3(n8175), .ZN(n12312) );
  INV_X1 U14713 ( .A(n12399), .ZN(n12311) );
  NAND4_X1 U14714 ( .A1(n12312), .A2(n7276), .A3(n12311), .A4(n12388), .ZN(
        n12313) );
  NOR3_X1 U14715 ( .A1(n12406), .A2(n12314), .A3(n12313), .ZN(n12315) );
  NAND4_X1 U14716 ( .A1(n12859), .A2(n7423), .A3(n12877), .A4(n12315), .ZN(
        n12316) );
  NOR4_X1 U14717 ( .A1(n12817), .A2(n7434), .A3(n12837), .A4(n12316), .ZN(
        n12319) );
  INV_X1 U14718 ( .A(n12454), .ZN(n12318) );
  NAND2_X1 U14719 ( .A1(n12318), .A2(n12317), .ZN(n12792) );
  NAND4_X1 U14720 ( .A1(n12778), .A2(n12320), .A3(n12319), .A4(n12792), .ZN(
        n12321) );
  NOR4_X1 U14721 ( .A1(n12739), .A2(n12465), .A3(n12767), .A4(n12321), .ZN(
        n12322) );
  INV_X1 U14722 ( .A(n12324), .ZN(n12325) );
  INV_X1 U14723 ( .A(n12465), .ZN(n12755) );
  XNOR2_X1 U14724 ( .A(n12327), .B(n12487), .ZN(n12328) );
  AOI21_X1 U14725 ( .B1(n12755), .B2(n12329), .A(n12328), .ZN(n12469) );
  NAND3_X1 U14726 ( .A1(n12330), .A2(n8026), .A3(n12487), .ZN(n12467) );
  NAND2_X1 U14727 ( .A1(n12333), .A2(n12331), .ZN(n12332) );
  MUX2_X1 U14728 ( .A(n12332), .B(n15140), .S(n8101), .Z(n12337) );
  INV_X1 U14729 ( .A(n12333), .ZN(n12335) );
  NAND2_X1 U14730 ( .A1(n12483), .A2(n12344), .ZN(n12334) );
  OAI21_X1 U14731 ( .B1(n12335), .B2(n10804), .A(n12334), .ZN(n12336) );
  NAND2_X1 U14732 ( .A1(n12337), .A2(n12336), .ZN(n12346) );
  NOR2_X1 U14733 ( .A1(n12339), .A2(n12338), .ZN(n12343) );
  NAND2_X1 U14734 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  AOI21_X1 U14735 ( .B1(n12346), .B2(n12343), .A(n12342), .ZN(n12348) );
  NAND3_X1 U14736 ( .A1(n12346), .A2(n12345), .A3(n12344), .ZN(n12347) );
  MUX2_X1 U14737 ( .A(n12348), .B(n12347), .S(n12487), .Z(n12355) );
  INV_X1 U14738 ( .A(n12351), .ZN(n12354) );
  NAND2_X1 U14739 ( .A1(n15144), .A2(n12349), .ZN(n12350) );
  NAND2_X1 U14740 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  NAND2_X1 U14741 ( .A1(n12487), .A2(n12352), .ZN(n12353) );
  OAI21_X1 U14742 ( .B1(n12355), .B2(n12354), .A(n12353), .ZN(n12359) );
  AOI21_X1 U14743 ( .B1(n12487), .B2(n12357), .A(n12356), .ZN(n12358) );
  NAND2_X1 U14744 ( .A1(n12359), .A2(n12358), .ZN(n12367) );
  NAND3_X1 U14745 ( .A1(n12367), .A2(n12366), .A3(n12360), .ZN(n12364) );
  AND2_X1 U14746 ( .A1(n12374), .A2(n12361), .ZN(n12363) );
  INV_X1 U14747 ( .A(n12369), .ZN(n12362) );
  AOI21_X1 U14748 ( .B1(n12364), .B2(n12363), .A(n12362), .ZN(n12372) );
  NAND3_X1 U14749 ( .A1(n12367), .A2(n12366), .A3(n12365), .ZN(n12370) );
  NAND3_X1 U14750 ( .A1(n12370), .A2(n12369), .A3(n12368), .ZN(n12371) );
  MUX2_X1 U14751 ( .A(n12372), .B(n12371), .S(n12487), .Z(n12382) );
  OAI21_X1 U14752 ( .B1(n12483), .B2(n12374), .A(n12373), .ZN(n12375) );
  INV_X1 U14753 ( .A(n12375), .ZN(n12381) );
  MUX2_X1 U14754 ( .A(n12377), .B(n12376), .S(n12483), .Z(n12379) );
  NAND2_X1 U14755 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  AOI21_X1 U14756 ( .B1(n12382), .B2(n12381), .A(n12380), .ZN(n12396) );
  NAND2_X1 U14757 ( .A1(n12487), .A2(n12383), .ZN(n12387) );
  NAND2_X1 U14758 ( .A1(n12483), .A2(n12384), .ZN(n12386) );
  MUX2_X1 U14759 ( .A(n12387), .B(n12386), .S(n12385), .Z(n12389) );
  NAND2_X1 U14760 ( .A1(n12389), .A2(n12388), .ZN(n12395) );
  NAND2_X1 U14761 ( .A1(n12487), .A2(n12390), .ZN(n12393) );
  NAND2_X1 U14762 ( .A1(n12483), .A2(n12391), .ZN(n12392) );
  MUX2_X1 U14763 ( .A(n12393), .B(n12392), .S(n12515), .Z(n12394) );
  OAI211_X1 U14764 ( .C1(n12396), .C2(n12395), .A(n7276), .B(n12394), .ZN(
        n12401) );
  MUX2_X1 U14765 ( .A(n12398), .B(n12397), .S(n12483), .Z(n12400) );
  AOI21_X1 U14766 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12412) );
  NAND2_X1 U14767 ( .A1(n12408), .A2(n12402), .ZN(n12405) );
  NAND2_X1 U14768 ( .A1(n12407), .A2(n12403), .ZN(n12404) );
  MUX2_X1 U14769 ( .A(n12405), .B(n12404), .S(n12487), .Z(n12411) );
  INV_X1 U14770 ( .A(n12406), .ZN(n12410) );
  MUX2_X1 U14771 ( .A(n12408), .B(n12407), .S(n12483), .Z(n12409) );
  OAI211_X1 U14772 ( .C1(n12412), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        n12416) );
  MUX2_X1 U14773 ( .A(n12414), .B(n12413), .S(n12487), .Z(n12415) );
  NAND3_X1 U14774 ( .A1(n12416), .A2(n7423), .A3(n12415), .ZN(n12417) );
  OAI21_X1 U14775 ( .B1(n12418), .B2(n12483), .A(n12417), .ZN(n12419) );
  NAND2_X1 U14776 ( .A1(n12419), .A2(n12877), .ZN(n12428) );
  INV_X1 U14777 ( .A(n12420), .ZN(n12421) );
  NAND2_X1 U14778 ( .A1(n12877), .A2(n12421), .ZN(n12424) );
  NAND3_X1 U14779 ( .A1(n12424), .A2(n12423), .A3(n12422), .ZN(n12425) );
  NAND2_X1 U14780 ( .A1(n12425), .A2(n12483), .ZN(n12427) );
  INV_X1 U14781 ( .A(n12429), .ZN(n12426) );
  AOI21_X1 U14782 ( .B1(n12428), .B2(n12427), .A(n12426), .ZN(n12432) );
  AOI21_X1 U14783 ( .B1(n12429), .B2(n12861), .A(n12483), .ZN(n12431) );
  NAND2_X1 U14784 ( .A1(n12487), .A2(n12839), .ZN(n12430) );
  OAI22_X1 U14785 ( .A1(n12432), .A2(n12431), .B1(n12938), .B2(n12430), .ZN(
        n12439) );
  INV_X1 U14786 ( .A(n12433), .ZN(n12438) );
  INV_X1 U14787 ( .A(n12434), .ZN(n12435) );
  NAND2_X1 U14788 ( .A1(n12440), .A2(n12435), .ZN(n12436) );
  NAND4_X1 U14789 ( .A1(n12446), .A2(n12487), .A3(n12437), .A4(n12436), .ZN(
        n12442) );
  AOI22_X1 U14790 ( .A1(n12439), .A2(n12844), .B1(n12438), .B2(n12442), .ZN(
        n12444) );
  NAND3_X1 U14791 ( .A1(n12445), .A2(n12483), .A3(n12440), .ZN(n12441) );
  NAND2_X1 U14792 ( .A1(n12442), .A2(n12441), .ZN(n12443) );
  OAI21_X1 U14793 ( .B1(n12444), .B2(n7434), .A(n12443), .ZN(n12448) );
  MUX2_X1 U14794 ( .A(n12446), .B(n12445), .S(n12487), .Z(n12447) );
  AOI21_X1 U14795 ( .B1(n12448), .B2(n12447), .A(n12804), .ZN(n12459) );
  MUX2_X1 U14796 ( .A(n12450), .B(n12449), .S(n12487), .Z(n12451) );
  NAND2_X1 U14797 ( .A1(n12792), .A2(n12451), .ZN(n12458) );
  OR2_X1 U14798 ( .A1(n12801), .A2(n12483), .ZN(n12452) );
  OAI21_X1 U14799 ( .B1(n12453), .B2(n12487), .A(n12452), .ZN(n12455) );
  NOR2_X1 U14800 ( .A1(n12455), .A2(n12454), .ZN(n12456) );
  NOR2_X1 U14801 ( .A1(n12782), .A2(n12456), .ZN(n12457) );
  OAI21_X1 U14802 ( .B1(n12459), .B2(n12458), .A(n12457), .ZN(n12463) );
  MUX2_X1 U14803 ( .A(n12461), .B(n12460), .S(n12483), .Z(n12462) );
  NAND2_X1 U14804 ( .A1(n12463), .A2(n12462), .ZN(n12464) );
  NAND2_X1 U14805 ( .A1(n12464), .A2(n12762), .ZN(n12466) );
  AOI21_X1 U14806 ( .B1(n12467), .B2(n12466), .A(n12465), .ZN(n12468) );
  NAND3_X1 U14807 ( .A1(n12727), .A2(n12470), .A3(n12473), .ZN(n12472) );
  NAND2_X1 U14808 ( .A1(n12475), .A2(n6473), .ZN(n12476) );
  NAND2_X1 U14809 ( .A1(n12477), .A2(n12713), .ZN(n12480) );
  OR2_X1 U14810 ( .A1(n12478), .A2(n12487), .ZN(n12479) );
  NAND2_X1 U14811 ( .A1(n12480), .A2(n12479), .ZN(n12481) );
  NAND2_X1 U14812 ( .A1(n12481), .A2(n7416), .ZN(n12488) );
  OAI21_X1 U14813 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n12485) );
  NAND2_X1 U14814 ( .A1(n12488), .A2(n12485), .ZN(n12486) );
  OAI211_X1 U14815 ( .C1(n12488), .C2(n12487), .A(n12486), .B(n12494), .ZN(
        n12490) );
  INV_X1 U14816 ( .A(n12494), .ZN(n12495) );
  NOR2_X1 U14817 ( .A1(n12502), .A2(n8139), .ZN(n12505) );
  OAI21_X1 U14818 ( .B1(n12506), .B2(n12503), .A(P3_B_REG_SCAN_IN), .ZN(n12504) );
  MUX2_X1 U14819 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12507), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14820 ( .A(n12698), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12521), .Z(
        P3_U3520) );
  MUX2_X1 U14821 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12508), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14822 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12697), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14823 ( .A(n12736), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12521), .Z(
        P3_U3517) );
  MUX2_X1 U14824 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12509), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14825 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n8195), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14826 ( .A(n12510), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12521), .Z(
        P3_U3514) );
  MUX2_X1 U14827 ( .A(n12768), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12521), .Z(
        P3_U3513) );
  MUX2_X1 U14828 ( .A(n12801), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12521), .Z(
        P3_U3512) );
  MUX2_X1 U14829 ( .A(n12800), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12521), .Z(
        P3_U3510) );
  MUX2_X1 U14830 ( .A(n12856), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12521), .Z(
        P3_U3508) );
  MUX2_X1 U14831 ( .A(n12839), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12521), .Z(
        P3_U3507) );
  MUX2_X1 U14832 ( .A(n12855), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12521), .Z(
        P3_U3506) );
  MUX2_X1 U14833 ( .A(n12511), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12521), .Z(
        P3_U3505) );
  MUX2_X1 U14834 ( .A(n12512), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12521), .Z(
        P3_U3504) );
  MUX2_X1 U14835 ( .A(n12513), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12521), .Z(
        P3_U3503) );
  MUX2_X1 U14836 ( .A(n12514), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12521), .Z(
        P3_U3501) );
  MUX2_X1 U14837 ( .A(n12515), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12521), .Z(
        P3_U3500) );
  MUX2_X1 U14838 ( .A(n12516), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12521), .Z(
        P3_U3499) );
  MUX2_X1 U14839 ( .A(n12517), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12521), .Z(
        P3_U3498) );
  MUX2_X1 U14840 ( .A(n12518), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12521), .Z(
        P3_U3497) );
  MUX2_X1 U14841 ( .A(n12519), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12521), .Z(
        P3_U3496) );
  MUX2_X1 U14842 ( .A(n12520), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12521), .Z(
        P3_U3495) );
  MUX2_X1 U14843 ( .A(n15142), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12521), .Z(
        P3_U3491) );
  NOR2_X1 U14844 ( .A1(n12532), .A2(n12522), .ZN(n12524) );
  NAND2_X1 U14845 ( .A1(n12530), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12553) );
  OR2_X1 U14846 ( .A1(n12530), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12525) );
  NAND2_X1 U14847 ( .A1(n12553), .A2(n12525), .ZN(n12540) );
  AOI21_X1 U14848 ( .B1(n12526), .B2(n12540), .A(n12550), .ZN(n12549) );
  NOR2_X1 U14849 ( .A1(n12532), .A2(n6552), .ZN(n12528) );
  AND2_X1 U14850 ( .A1(n12530), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12570) );
  NOR2_X1 U14851 ( .A1(n12530), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12529) );
  OR2_X1 U14852 ( .A1(n12570), .A2(n12529), .ZN(n12567) );
  XNOR2_X1 U14853 ( .A(n12568), .B(n12567), .ZN(n12547) );
  NOR2_X1 U14854 ( .A1(n15122), .A2(n12530), .ZN(n12545) );
  INV_X1 U14855 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15295) );
  INV_X1 U14856 ( .A(n12531), .ZN(n12543) );
  NAND2_X1 U14857 ( .A1(n12533), .A2(n12532), .ZN(n12536) );
  INV_X1 U14858 ( .A(n12567), .ZN(n12537) );
  INV_X1 U14859 ( .A(n12534), .ZN(n12535) );
  NAND2_X1 U14860 ( .A1(n12536), .A2(n12535), .ZN(n12539) );
  NAND2_X1 U14861 ( .A1(n9796), .A2(n12537), .ZN(n12538) );
  OAI211_X1 U14862 ( .C1(n9796), .C2(n12540), .A(n12539), .B(n12538), .ZN(
        n12541) );
  NAND3_X1 U14863 ( .A1(n15131), .A2(n12556), .A3(n12541), .ZN(n12542) );
  OAI211_X1 U14864 ( .C1(n15126), .C2(n15295), .A(n12543), .B(n12542), .ZN(
        n12544) );
  AOI211_X1 U14865 ( .C1(n12547), .C2(n12546), .A(n12545), .B(n12544), .ZN(
        n12548) );
  OAI21_X1 U14866 ( .B1(n12549), .B2(n15125), .A(n12548), .ZN(P3_U3196) );
  INV_X1 U14867 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14498) );
  XNOR2_X1 U14868 ( .A(n12579), .B(n12578), .ZN(n12551) );
  AOI21_X1 U14869 ( .B1(n14498), .B2(n12551), .A(n12580), .ZN(n12577) );
  NAND2_X1 U14870 ( .A1(n15082), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12566) );
  INV_X1 U14871 ( .A(n12552), .ZN(n12565) );
  INV_X1 U14872 ( .A(n12570), .ZN(n12554) );
  MUX2_X1 U14873 ( .A(n12554), .B(n12553), .S(n12626), .Z(n12555) );
  NAND2_X1 U14874 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  AND2_X1 U14875 ( .A1(n12557), .A2(n12579), .ZN(n12558) );
  NOR2_X1 U14876 ( .A1(n12557), .A2(n12579), .ZN(n12587) );
  OR2_X1 U14877 ( .A1(n12558), .A2(n12587), .ZN(n12562) );
  OR2_X1 U14878 ( .A1(n12675), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U14879 ( .A1(n12626), .A2(n14498), .ZN(n12559) );
  AND2_X1 U14880 ( .A1(n12560), .A2(n12559), .ZN(n12561) );
  NOR2_X1 U14881 ( .A1(n12562), .A2(n12561), .ZN(n12586) );
  AND2_X1 U14882 ( .A1(n12562), .A2(n12561), .ZN(n12563) );
  OAI21_X1 U14883 ( .B1(n12586), .B2(n12563), .A(n15131), .ZN(n12564) );
  NAND3_X1 U14884 ( .A1(n12566), .A2(n12565), .A3(n12564), .ZN(n12575) );
  INV_X1 U14885 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12572) );
  NOR2_X1 U14886 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  NOR2_X2 U14887 ( .A1(n12570), .A2(n12569), .ZN(n12596) );
  AOI21_X1 U14888 ( .B1(n12572), .B2(n12571), .A(n12598), .ZN(n12573) );
  NOR2_X1 U14889 ( .A1(n12573), .A2(n15136), .ZN(n12574) );
  AOI211_X1 U14890 ( .C1(n15106), .C2(n12597), .A(n12575), .B(n12574), .ZN(
        n12576) );
  OAI21_X1 U14891 ( .B1(n12577), .B2(n15125), .A(n12576), .ZN(P3_U3197) );
  AND2_X1 U14892 ( .A1(n12579), .A2(n12578), .ZN(n12581) );
  NAND2_X1 U14893 ( .A1(n12600), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U14894 ( .A1(n12602), .A2(n12589), .ZN(n12582) );
  NAND2_X1 U14895 ( .A1(n12612), .A2(n12582), .ZN(n12584) );
  INV_X1 U14896 ( .A(n12613), .ZN(n12583) );
  AOI21_X1 U14897 ( .B1(n12585), .B2(n12584), .A(n12583), .ZN(n12611) );
  NOR2_X1 U14898 ( .A1(n12587), .A2(n12586), .ZN(n12624) );
  INV_X1 U14899 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12601) );
  AOI21_X1 U14900 ( .B1(n12675), .B2(P3_REG1_REG_16__SCAN_IN), .A(n12600), 
        .ZN(n12588) );
  OAI21_X1 U14901 ( .B1(n12675), .B2(n12601), .A(n12588), .ZN(n12623) );
  OR2_X1 U14902 ( .A1(n12675), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U14903 ( .A1(n12675), .A2(n12589), .ZN(n12590) );
  AND3_X1 U14904 ( .A1(n12591), .A2(n12590), .A3(n12600), .ZN(n12625) );
  INV_X1 U14905 ( .A(n12625), .ZN(n12592) );
  NAND2_X1 U14906 ( .A1(n12623), .A2(n12592), .ZN(n12593) );
  XNOR2_X1 U14907 ( .A(n12624), .B(n12593), .ZN(n12609) );
  AOI21_X1 U14908 ( .B1(n15082), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12594), 
        .ZN(n12595) );
  OAI21_X1 U14909 ( .B1(n15122), .B2(n12600), .A(n12595), .ZN(n12608) );
  NOR2_X1 U14910 ( .A1(n12597), .A2(n12596), .ZN(n12599) );
  NAND2_X1 U14911 ( .A1(n12600), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U14912 ( .A1(n12602), .A2(n12601), .ZN(n12603) );
  NAND2_X1 U14913 ( .A1(n12616), .A2(n12603), .ZN(n12604) );
  NAND2_X1 U14914 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  AOI21_X1 U14915 ( .B1(n12617), .B2(n12606), .A(n15136), .ZN(n12607) );
  AOI211_X1 U14916 ( .C1(n15131), .C2(n12609), .A(n12608), .B(n12607), .ZN(
        n12610) );
  OAI21_X1 U14917 ( .B1(n12611), .B2(n15125), .A(n12610), .ZN(P3_U3198) );
  AOI21_X1 U14918 ( .B1(n12615), .B2(n12614), .A(n12636), .ZN(n12634) );
  INV_X1 U14919 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12618) );
  AOI21_X1 U14920 ( .B1(n12619), .B2(n12618), .A(n12642), .ZN(n12622) );
  AOI21_X1 U14921 ( .B1(n15082), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12620), 
        .ZN(n12621) );
  OAI21_X1 U14922 ( .B1(n12622), .B2(n15136), .A(n12621), .ZN(n12632) );
  OAI21_X1 U14923 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n12630) );
  OR2_X1 U14924 ( .A1(n12675), .A2(n12618), .ZN(n12628) );
  NAND2_X1 U14925 ( .A1(n12626), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n12627) );
  NAND2_X1 U14926 ( .A1(n12628), .A2(n12627), .ZN(n12650) );
  XNOR2_X1 U14927 ( .A(n12651), .B(n12650), .ZN(n12629) );
  NOR2_X1 U14928 ( .A1(n12630), .A2(n12629), .ZN(n12652) );
  AOI211_X1 U14929 ( .C1(n12630), .C2(n12629), .A(n12652), .B(n15110), .ZN(
        n12631) );
  OAI21_X1 U14930 ( .B1(n12634), .B2(n15125), .A(n12633), .ZN(P3_U3199) );
  NOR2_X1 U14931 ( .A1(n12641), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U14932 ( .A1(n12644), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12665) );
  OAI21_X1 U14933 ( .B1(n12644), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12665), 
        .ZN(n12638) );
  NOR2_X1 U14934 ( .A1(n12641), .A2(n12640), .ZN(n12643) );
  NAND2_X1 U14935 ( .A1(n12644), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12681) );
  OAI21_X1 U14936 ( .B1(n12644), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12681), 
        .ZN(n12645) );
  AOI21_X1 U14937 ( .B1(n6493), .B2(n12645), .A(n12683), .ZN(n12646) );
  NOR2_X1 U14938 ( .A1(n12646), .A2(n15136), .ZN(n12662) );
  INV_X1 U14939 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U14940 ( .A1(n15106), .A2(n12668), .ZN(n12660) );
  INV_X1 U14941 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12647) );
  OR2_X1 U14942 ( .A1(n12675), .A2(n12647), .ZN(n12649) );
  NAND2_X1 U14943 ( .A1(n12675), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12648) );
  AND2_X1 U14944 ( .A1(n12649), .A2(n12648), .ZN(n12656) );
  NAND2_X1 U14945 ( .A1(n12651), .A2(n12650), .ZN(n12654) );
  INV_X1 U14946 ( .A(n12652), .ZN(n12653) );
  NAND2_X1 U14947 ( .A1(n12654), .A2(n12653), .ZN(n12667) );
  XNOR2_X1 U14948 ( .A(n12667), .B(n12668), .ZN(n12655) );
  NAND2_X1 U14949 ( .A1(n12655), .A2(n12656), .ZN(n12671) );
  OAI21_X1 U14950 ( .B1(n12656), .B2(n12655), .A(n12671), .ZN(n12658) );
  AOI21_X1 U14951 ( .B1(n15131), .B2(n12658), .A(n12657), .ZN(n12659) );
  OAI211_X1 U14952 ( .C1(n14483), .C2(n15126), .A(n12660), .B(n12659), .ZN(
        n12661) );
  NOR2_X1 U14953 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  OAI21_X1 U14954 ( .B1(n12664), .B2(n15125), .A(n12663), .ZN(P3_U3200) );
  XNOR2_X1 U14955 ( .A(n12687), .B(n12928), .ZN(n12673) );
  INV_X1 U14956 ( .A(n12673), .ZN(n12666) );
  INV_X1 U14957 ( .A(n12667), .ZN(n12669) );
  NAND2_X1 U14958 ( .A1(n12669), .A2(n12668), .ZN(n12670) );
  NAND2_X1 U14959 ( .A1(n12671), .A2(n12670), .ZN(n12677) );
  INV_X1 U14960 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12672) );
  MUX2_X1 U14961 ( .A(n12672), .B(P3_REG2_REG_19__SCAN_IN), .S(n12687), .Z(
        n12684) );
  NAND2_X1 U14962 ( .A1(n12673), .A2(n12675), .ZN(n12674) );
  OAI21_X1 U14963 ( .B1(n12684), .B2(n12675), .A(n12674), .ZN(n12676) );
  XNOR2_X1 U14964 ( .A(n12677), .B(n12676), .ZN(n12680) );
  NAND2_X1 U14965 ( .A1(n15082), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12679) );
  OAI211_X1 U14966 ( .C1(n12680), .C2(n15110), .A(n12679), .B(n12678), .ZN(
        n12686) );
  INV_X1 U14967 ( .A(n12681), .ZN(n12682) );
  NAND2_X1 U14968 ( .A1(n12688), .A2(n15151), .ZN(n12691) );
  OR2_X1 U14969 ( .A1(n12690), .A2(n12689), .ZN(n14491) );
  AOI21_X1 U14970 ( .B1(n12691), .B2(n14491), .A(n15156), .ZN(n12693) );
  AOI21_X1 U14971 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15156), .A(n12693), 
        .ZN(n12692) );
  OAI21_X1 U14972 ( .B1(n12945), .B2(n12883), .A(n12692), .ZN(P3_U3202) );
  AOI21_X1 U14973 ( .B1(n15156), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12693), 
        .ZN(n12694) );
  OAI21_X1 U14974 ( .B1(n14492), .B2(n12883), .A(n12694), .ZN(P3_U3203) );
  OAI211_X1 U14975 ( .C1(n12696), .C2(n12703), .A(n12695), .B(n12854), .ZN(
        n12700) );
  AOI22_X1 U14976 ( .A1(n12698), .A2(n15145), .B1(n15143), .B2(n12697), .ZN(
        n12699) );
  NAND2_X1 U14977 ( .A1(n12700), .A2(n12699), .ZN(n12890) );
  INV_X1 U14978 ( .A(n12890), .ZN(n12709) );
  INV_X1 U14979 ( .A(n12701), .ZN(n12702) );
  NOR2_X1 U14980 ( .A1(n12711), .A2(n12702), .ZN(n12704) );
  XNOR2_X1 U14981 ( .A(n12703), .B(n12704), .ZN(n12891) );
  AOI22_X1 U14982 ( .A1(n12705), .A2(n12881), .B1(n15156), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12706) );
  OAI21_X1 U14983 ( .B1(n12948), .B2(n12883), .A(n12706), .ZN(n12707) );
  AOI21_X1 U14984 ( .B1(n12891), .B2(n12885), .A(n12707), .ZN(n12708) );
  OAI21_X1 U14985 ( .B1(n12709), .B2(n15156), .A(n12708), .ZN(P3_U3205) );
  INV_X1 U14986 ( .A(n12711), .ZN(n12712) );
  OAI22_X1 U14987 ( .A1(n12715), .A2(n12873), .B1(n12714), .B2(n12875), .ZN(
        n12716) );
  INV_X1 U14988 ( .A(n12894), .ZN(n12723) );
  AOI22_X1 U14989 ( .A1(n12719), .A2(n12881), .B1(n15156), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12720) );
  OAI21_X1 U14990 ( .B1(n12951), .B2(n12883), .A(n12720), .ZN(n12721) );
  AOI21_X1 U14991 ( .B1(n12895), .B2(n15152), .A(n12721), .ZN(n12722) );
  OAI21_X1 U14992 ( .B1(n12723), .B2(n15156), .A(n12722), .ZN(P3_U3206) );
  XOR2_X1 U14993 ( .A(n12724), .B(n12727), .Z(n12725) );
  OAI222_X1 U14994 ( .A1(n12873), .A2(n12726), .B1(n12875), .B2(n12749), .C1(
        n12725), .C2(n15149), .ZN(n12897) );
  INV_X1 U14995 ( .A(n12897), .ZN(n12733) );
  XNOR2_X1 U14996 ( .A(n12728), .B(n12727), .ZN(n12898) );
  AOI22_X1 U14997 ( .A1(n12729), .A2(n12881), .B1(n15156), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12730) );
  OAI21_X1 U14998 ( .B1(n12955), .B2(n12883), .A(n12730), .ZN(n12731) );
  AOI21_X1 U14999 ( .B1(n12898), .B2(n12885), .A(n12731), .ZN(n12732) );
  OAI21_X1 U15000 ( .B1(n12733), .B2(n15156), .A(n12732), .ZN(P3_U3207) );
  OAI211_X1 U15001 ( .C1(n12735), .C2(n12739), .A(n12734), .B(n12854), .ZN(
        n12738) );
  AOI22_X1 U15002 ( .A1(n12736), .A2(n15145), .B1(n8195), .B2(n15143), .ZN(
        n12737) );
  AND2_X1 U15003 ( .A1(n12738), .A2(n12737), .ZN(n12903) );
  XNOR2_X1 U15004 ( .A(n12740), .B(n12739), .ZN(n12901) );
  NAND2_X1 U15005 ( .A1(n12900), .A2(n12741), .ZN(n12744) );
  AOI22_X1 U15006 ( .A1(n12742), .A2(n15151), .B1(n15156), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15007 ( .A1(n12744), .A2(n12743), .ZN(n12745) );
  AOI21_X1 U15008 ( .B1(n12901), .B2(n12885), .A(n12745), .ZN(n12746) );
  OAI21_X1 U15009 ( .B1(n12903), .B2(n15156), .A(n12746), .ZN(P3_U3208) );
  INV_X1 U15010 ( .A(n12747), .ZN(n12748) );
  AOI21_X1 U15011 ( .B1(n12748), .B2(n12755), .A(n15149), .ZN(n12752) );
  OAI22_X1 U15012 ( .A1(n12749), .A2(n12873), .B1(n8026), .B2(n12875), .ZN(
        n12750) );
  AOI21_X1 U15013 ( .B1(n12752), .B2(n12751), .A(n12750), .ZN(n12907) );
  INV_X1 U15014 ( .A(n12753), .ZN(n12756) );
  OAI21_X1 U15015 ( .B1(n12756), .B2(n12755), .A(n12754), .ZN(n12905) );
  AOI22_X1 U15016 ( .A1(n15151), .A2(n12757), .B1(n15156), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12758) );
  OAI21_X1 U15017 ( .B1(n12759), .B2(n12883), .A(n12758), .ZN(n12760) );
  AOI21_X1 U15018 ( .B1(n12905), .B2(n12885), .A(n12760), .ZN(n12761) );
  OAI21_X1 U15019 ( .B1(n12907), .B2(n15156), .A(n12761), .ZN(P3_U3209) );
  OR2_X1 U15020 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  NAND2_X1 U15021 ( .A1(n12765), .A2(n12764), .ZN(n12772) );
  OAI211_X1 U15022 ( .C1(n6563), .C2(n12767), .A(n12766), .B(n12854), .ZN(
        n12770) );
  AOI22_X1 U15023 ( .A1(n8195), .A2(n15145), .B1(n15143), .B2(n12768), .ZN(
        n12769) );
  OAI211_X1 U15024 ( .C1(n12771), .C2(n12772), .A(n12770), .B(n12769), .ZN(
        n12908) );
  INV_X1 U15025 ( .A(n12908), .ZN(n12777) );
  INV_X1 U15026 ( .A(n12772), .ZN(n12909) );
  AOI22_X1 U15027 ( .A1(n15156), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15151), 
        .B2(n12773), .ZN(n12774) );
  OAI21_X1 U15028 ( .B1(n12961), .B2(n12883), .A(n12774), .ZN(n12775) );
  AOI21_X1 U15029 ( .B1(n12909), .B2(n15152), .A(n12775), .ZN(n12776) );
  OAI21_X1 U15030 ( .B1(n12777), .B2(n15156), .A(n12776), .ZN(P3_U3210) );
  XNOR2_X1 U15031 ( .A(n12779), .B(n12778), .ZN(n12780) );
  OAI222_X1 U15032 ( .A1(n12875), .A2(n12781), .B1(n12873), .B2(n8026), .C1(
        n15149), .C2(n12780), .ZN(n12912) );
  INV_X1 U15033 ( .A(n12912), .ZN(n12788) );
  XNOR2_X1 U15034 ( .A(n12783), .B(n12782), .ZN(n12913) );
  AOI22_X1 U15035 ( .A1(n15156), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15151), 
        .B2(n12784), .ZN(n12785) );
  OAI21_X1 U15036 ( .B1(n12965), .B2(n12883), .A(n12785), .ZN(n12786) );
  AOI21_X1 U15037 ( .B1(n12913), .B2(n12885), .A(n12786), .ZN(n12787) );
  OAI21_X1 U15038 ( .B1(n12788), .B2(n15156), .A(n12787), .ZN(P3_U3211) );
  XOR2_X1 U15039 ( .A(n12792), .B(n12789), .Z(n12790) );
  OAI222_X1 U15040 ( .A1(n12875), .A2(n12816), .B1(n12873), .B2(n8007), .C1(
        n15149), .C2(n12790), .ZN(n12916) );
  INV_X1 U15041 ( .A(n12916), .ZN(n12797) );
  XOR2_X1 U15042 ( .A(n12792), .B(n12791), .Z(n12917) );
  AOI22_X1 U15043 ( .A1(n15156), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12881), 
        .B2(n12793), .ZN(n12794) );
  OAI21_X1 U15044 ( .B1(n12969), .B2(n12883), .A(n12794), .ZN(n12795) );
  AOI21_X1 U15045 ( .B1(n12917), .B2(n12885), .A(n12795), .ZN(n12796) );
  OAI21_X1 U15046 ( .B1(n12797), .B2(n15156), .A(n12796), .ZN(P3_U3212) );
  OAI211_X1 U15047 ( .C1(n12799), .C2(n12804), .A(n12798), .B(n12854), .ZN(
        n12803) );
  AOI22_X1 U15048 ( .A1(n12801), .A2(n15145), .B1(n15143), .B2(n12800), .ZN(
        n12802) );
  NAND2_X1 U15049 ( .A1(n12803), .A2(n12802), .ZN(n12921) );
  INV_X1 U15050 ( .A(n12922), .ZN(n12807) );
  AND2_X1 U15051 ( .A1(n12805), .A2(n12804), .ZN(n12920) );
  NOR3_X1 U15052 ( .A1(n12807), .A2(n12920), .A3(n12806), .ZN(n12811) );
  AOI22_X1 U15053 ( .A1(n15156), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15151), 
        .B2(n12808), .ZN(n12809) );
  OAI21_X1 U15054 ( .B1(n12973), .B2(n12883), .A(n12809), .ZN(n12810) );
  AOI211_X1 U15055 ( .C1(n12921), .C2(n15154), .A(n12811), .B(n12810), .ZN(
        n12812) );
  INV_X1 U15056 ( .A(n12812), .ZN(P3_U3213) );
  OAI211_X1 U15057 ( .C1(n6585), .C2(n12817), .A(n12813), .B(n12854), .ZN(
        n12815) );
  NAND2_X1 U15058 ( .A1(n12840), .A2(n15143), .ZN(n12814) );
  OAI211_X1 U15059 ( .C1(n12816), .C2(n12873), .A(n12815), .B(n12814), .ZN(
        n12926) );
  INV_X1 U15060 ( .A(n12926), .ZN(n12823) );
  XNOR2_X1 U15061 ( .A(n12818), .B(n12817), .ZN(n12927) );
  AOI22_X1 U15062 ( .A1(n15156), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12881), 
        .B2(n12819), .ZN(n12820) );
  OAI21_X1 U15063 ( .B1(n12977), .B2(n12883), .A(n12820), .ZN(n12821) );
  AOI21_X1 U15064 ( .B1(n12927), .B2(n12885), .A(n12821), .ZN(n12822) );
  OAI21_X1 U15065 ( .B1(n12823), .B2(n15156), .A(n12822), .ZN(P3_U3214) );
  AOI21_X1 U15066 ( .B1(n12826), .B2(n12825), .A(n12824), .ZN(n12827) );
  OAI222_X1 U15067 ( .A1(n12875), .A2(n12829), .B1(n12873), .B2(n12828), .C1(
        n15149), .C2(n12827), .ZN(n12930) );
  INV_X1 U15068 ( .A(n12930), .ZN(n12835) );
  AOI21_X1 U15069 ( .B1(n7434), .B2(n12830), .A(n6578), .ZN(n12931) );
  AOI22_X1 U15070 ( .A1(n15156), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12881), 
        .B2(n12831), .ZN(n12832) );
  OAI21_X1 U15071 ( .B1(n12982), .B2(n12883), .A(n12832), .ZN(n12833) );
  AOI21_X1 U15072 ( .B1(n12931), .B2(n12885), .A(n12833), .ZN(n12834) );
  OAI21_X1 U15073 ( .B1(n12835), .B2(n15156), .A(n12834), .ZN(P3_U3215) );
  OAI211_X1 U15074 ( .C1(n12838), .C2(n12837), .A(n12836), .B(n12854), .ZN(
        n12842) );
  AOI22_X1 U15075 ( .A1(n15145), .A2(n12840), .B1(n15143), .B2(n12839), .ZN(
        n12841) );
  AND2_X1 U15076 ( .A1(n12842), .A2(n12841), .ZN(n12937) );
  OAI21_X1 U15077 ( .B1(n12845), .B2(n12844), .A(n12843), .ZN(n12935) );
  AOI22_X1 U15078 ( .A1(n15156), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12881), 
        .B2(n12846), .ZN(n12847) );
  OAI21_X1 U15079 ( .B1(n12848), .B2(n12883), .A(n12847), .ZN(n12849) );
  AOI21_X1 U15080 ( .B1(n12935), .B2(n12885), .A(n12849), .ZN(n12850) );
  OAI21_X1 U15081 ( .B1(n12937), .B2(n15156), .A(n12850), .ZN(P3_U3216) );
  NAND2_X1 U15082 ( .A1(n12852), .A2(n12859), .ZN(n12853) );
  NAND3_X1 U15083 ( .A1(n12851), .A2(n12854), .A3(n12853), .ZN(n12858) );
  AOI22_X1 U15084 ( .A1(n15145), .A2(n12856), .B1(n15143), .B2(n12855), .ZN(
        n12857) );
  NAND2_X1 U15085 ( .A1(n12858), .A2(n12857), .ZN(n12942) );
  INV_X1 U15086 ( .A(n12942), .ZN(n12869) );
  INV_X1 U15087 ( .A(n12859), .ZN(n12860) );
  NAND3_X1 U15088 ( .A1(n12876), .A2(n12861), .A3(n12860), .ZN(n12862) );
  NAND2_X1 U15089 ( .A1(n12863), .A2(n12862), .ZN(n12939) );
  AOI22_X1 U15090 ( .A1(n15156), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12881), 
        .B2(n12864), .ZN(n12865) );
  OAI21_X1 U15091 ( .B1(n12866), .B2(n12883), .A(n12865), .ZN(n12867) );
  AOI21_X1 U15092 ( .B1(n12939), .B2(n12885), .A(n12867), .ZN(n12868) );
  OAI21_X1 U15093 ( .B1(n12869), .B2(n15156), .A(n12868), .ZN(P3_U3217) );
  XOR2_X1 U15094 ( .A(n12870), .B(n12877), .Z(n12871) );
  OAI222_X1 U15095 ( .A1(n12875), .A2(n12874), .B1(n12873), .B2(n12872), .C1(
        n12871), .C2(n15149), .ZN(n14497) );
  INV_X1 U15096 ( .A(n14497), .ZN(n12887) );
  OAI21_X1 U15097 ( .B1(n12878), .B2(n12877), .A(n12876), .ZN(n14494) );
  AOI22_X1 U15098 ( .A1(n15156), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12881), 
        .B2(n12880), .ZN(n12882) );
  OAI21_X1 U15099 ( .B1(n7420), .B2(n12883), .A(n12882), .ZN(n12884) );
  AOI21_X1 U15100 ( .B1(n14494), .B2(n12885), .A(n12884), .ZN(n12886) );
  OAI21_X1 U15101 ( .B1(n12887), .B2(n15156), .A(n12886), .ZN(P3_U3218) );
  INV_X1 U15102 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12888) );
  MUX2_X1 U15103 ( .A(n14491), .B(n12888), .S(n15196), .Z(n12889) );
  OAI21_X1 U15104 ( .B1(n12945), .B2(n12933), .A(n12889), .ZN(P3_U3490) );
  INV_X1 U15105 ( .A(n12893), .ZN(n15164) );
  AOI21_X1 U15106 ( .B1(n12898), .B2(n15177), .A(n12897), .ZN(n12952) );
  MUX2_X1 U15107 ( .A(n15227), .B(n12952), .S(n15199), .Z(n12899) );
  OAI21_X1 U15108 ( .B1(n12955), .B2(n12933), .A(n12899), .ZN(P3_U3485) );
  AOI22_X1 U15109 ( .A1(n12901), .A2(n15177), .B1(n15184), .B2(n12900), .ZN(
        n12902) );
  NAND2_X1 U15110 ( .A1(n12903), .A2(n12902), .ZN(n12956) );
  MUX2_X1 U15111 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12956), .S(n15199), .Z(
        P3_U3484) );
  AOI22_X1 U15112 ( .A1(n12905), .A2(n15177), .B1(n15184), .B2(n12904), .ZN(
        n12906) );
  NAND2_X1 U15113 ( .A1(n12907), .A2(n12906), .ZN(n12957) );
  MUX2_X1 U15114 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12957), .S(n15199), .Z(
        P3_U3483) );
  AOI21_X1 U15115 ( .B1(n15164), .B2(n12909), .A(n12908), .ZN(n12958) );
  MUX2_X1 U15116 ( .A(n12910), .B(n12958), .S(n15199), .Z(n12911) );
  OAI21_X1 U15117 ( .B1(n12961), .B2(n12933), .A(n12911), .ZN(P3_U3482) );
  AOI21_X1 U15118 ( .B1(n15177), .B2(n12913), .A(n12912), .ZN(n12962) );
  MUX2_X1 U15119 ( .A(n12914), .B(n12962), .S(n15199), .Z(n12915) );
  OAI21_X1 U15120 ( .B1(n12965), .B2(n12933), .A(n12915), .ZN(P3_U3481) );
  AOI21_X1 U15121 ( .B1(n12917), .B2(n15177), .A(n12916), .ZN(n12966) );
  MUX2_X1 U15122 ( .A(n12918), .B(n12966), .S(n15199), .Z(n12919) );
  OAI21_X1 U15123 ( .B1(n12969), .B2(n12933), .A(n12919), .ZN(P3_U3480) );
  NOR2_X1 U15124 ( .A1(n12920), .A2(n15179), .ZN(n12923) );
  AOI21_X1 U15125 ( .B1(n12923), .B2(n12922), .A(n12921), .ZN(n12970) );
  MUX2_X1 U15126 ( .A(n12924), .B(n12970), .S(n15199), .Z(n12925) );
  OAI21_X1 U15127 ( .B1(n12973), .B2(n12933), .A(n12925), .ZN(P3_U3479) );
  AOI21_X1 U15128 ( .B1(n15177), .B2(n12927), .A(n12926), .ZN(n12974) );
  MUX2_X1 U15129 ( .A(n12928), .B(n12974), .S(n15199), .Z(n12929) );
  OAI21_X1 U15130 ( .B1(n12933), .B2(n12977), .A(n12929), .ZN(P3_U3478) );
  AOI21_X1 U15131 ( .B1(n12931), .B2(n15177), .A(n12930), .ZN(n12978) );
  MUX2_X1 U15132 ( .A(n15280), .B(n12978), .S(n15199), .Z(n12932) );
  OAI21_X1 U15133 ( .B1(n12982), .B2(n12933), .A(n12932), .ZN(P3_U3477) );
  AOI22_X1 U15134 ( .A1(n12935), .A2(n15177), .B1(n15184), .B2(n12934), .ZN(
        n12936) );
  NAND2_X1 U15135 ( .A1(n12937), .A2(n12936), .ZN(n12983) );
  MUX2_X1 U15136 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12983), .S(n15199), .Z(
        P3_U3476) );
  AND2_X1 U15137 ( .A1(n12938), .A2(n15184), .ZN(n12941) );
  AND2_X1 U15138 ( .A1(n12939), .A2(n15177), .ZN(n12940) );
  MUX2_X1 U15139 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12984), .S(n15199), .Z(
        P3_U3475) );
  INV_X1 U15140 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12943) );
  MUX2_X1 U15141 ( .A(n14491), .B(n12943), .S(n15187), .Z(n12944) );
  OAI21_X1 U15142 ( .B1(n12945), .B2(n12981), .A(n12944), .ZN(P3_U3458) );
  INV_X1 U15143 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12947) );
  INV_X1 U15144 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12950) );
  INV_X1 U15145 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12953) );
  MUX2_X1 U15146 ( .A(n12953), .B(n12952), .S(n15185), .Z(n12954) );
  OAI21_X1 U15147 ( .B1(n12955), .B2(n12981), .A(n12954), .ZN(P3_U3453) );
  MUX2_X1 U15148 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12956), .S(n15185), .Z(
        P3_U3452) );
  MUX2_X1 U15149 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12957), .S(n15185), .Z(
        P3_U3451) );
  INV_X1 U15150 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12959) );
  MUX2_X1 U15151 ( .A(n12959), .B(n12958), .S(n15185), .Z(n12960) );
  OAI21_X1 U15152 ( .B1(n12961), .B2(n12981), .A(n12960), .ZN(P3_U3450) );
  INV_X1 U15153 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12963) );
  MUX2_X1 U15154 ( .A(n12963), .B(n12962), .S(n15185), .Z(n12964) );
  OAI21_X1 U15155 ( .B1(n12965), .B2(n12981), .A(n12964), .ZN(P3_U3449) );
  INV_X1 U15156 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12967) );
  MUX2_X1 U15157 ( .A(n12967), .B(n12966), .S(n15185), .Z(n12968) );
  OAI21_X1 U15158 ( .B1(n12969), .B2(n12981), .A(n12968), .ZN(P3_U3448) );
  INV_X1 U15159 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12971) );
  MUX2_X1 U15160 ( .A(n12971), .B(n12970), .S(n15185), .Z(n12972) );
  OAI21_X1 U15161 ( .B1(n12973), .B2(n12981), .A(n12972), .ZN(P3_U3447) );
  INV_X1 U15162 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12975) );
  MUX2_X1 U15163 ( .A(n12975), .B(n12974), .S(n15185), .Z(n12976) );
  OAI21_X1 U15164 ( .B1(n12981), .B2(n12977), .A(n12976), .ZN(P3_U3446) );
  INV_X1 U15165 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12979) );
  MUX2_X1 U15166 ( .A(n12979), .B(n12978), .S(n15185), .Z(n12980) );
  OAI21_X1 U15167 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(P3_U3444) );
  MUX2_X1 U15168 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12983), .S(n15185), .Z(
        P3_U3441) );
  MUX2_X1 U15169 ( .A(n12984), .B(P3_REG0_REG_16__SCAN_IN), .S(n15187), .Z(
        P3_U3438) );
  MUX2_X1 U15170 ( .A(n12985), .B(P3_D_REG_1__SCAN_IN), .S(n12986), .Z(
        P3_U3377) );
  MUX2_X1 U15171 ( .A(n12987), .B(P3_D_REG_0__SCAN_IN), .S(n12986), .Z(
        P3_U3376) );
  NAND2_X1 U15172 ( .A1(n12988), .A2(n14446), .ZN(n12992) );
  OR4_X1 U15173 ( .A1(n12989), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12990), .A4(
        P3_U3151), .ZN(n12991) );
  OAI211_X1 U15174 ( .C1(n12993), .C2(n12997), .A(n12992), .B(n12991), .ZN(
        P3_U3264) );
  INV_X1 U15175 ( .A(n12994), .ZN(n12995) );
  INV_X1 U15176 ( .A(n12998), .ZN(n12999) );
  OAI222_X1 U15177 ( .A1(n12997), .A2(n13000), .B1(n14451), .B2(n12999), .C1(
        n8139), .C2(P3_U3151), .ZN(P3_U3267) );
  AOI21_X1 U15178 ( .B1(n13002), .B2(n13001), .A(n14777), .ZN(n13007) );
  NAND2_X1 U15179 ( .A1(n13568), .A2(n14782), .ZN(n13004) );
  INV_X1 U15180 ( .A(n13318), .ZN(n13319) );
  INV_X1 U15181 ( .A(n13124), .ZN(n13289) );
  OAI22_X1 U15182 ( .A1(n13319), .A2(n13508), .B1(n13289), .B2(n13510), .ZN(
        n13567) );
  AOI22_X1 U15183 ( .A1(n14534), .A2(n13567), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13003) );
  OAI211_X1 U15184 ( .C1(n14797), .C2(n13357), .A(n13004), .B(n13003), .ZN(
        n13005) );
  AOI21_X1 U15185 ( .B1(n13007), .B2(n13006), .A(n13005), .ZN(n13008) );
  INV_X1 U15186 ( .A(n13008), .ZN(P2_U3186) );
  INV_X1 U15187 ( .A(n13074), .ZN(n13009) );
  NOR2_X1 U15188 ( .A1(n13009), .A2(n13071), .ZN(n13018) );
  NOR2_X1 U15189 ( .A1(n7203), .A2(n13110), .ZN(n13077) );
  INV_X1 U15190 ( .A(n13077), .ZN(n13017) );
  NAND3_X1 U15191 ( .A1(n13018), .A2(n14788), .A3(n13010), .ZN(n13016) );
  AND2_X1 U15192 ( .A1(n13314), .A2(n13254), .ZN(n13011) );
  AOI21_X1 U15193 ( .B1(n13125), .B2(n13116), .A(n13011), .ZN(n13413) );
  INV_X1 U15194 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13012) );
  OAI22_X1 U15195 ( .A1(n13413), .A2(n14787), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13012), .ZN(n13014) );
  INV_X1 U15196 ( .A(n13410), .ZN(n13593) );
  NOR2_X1 U15197 ( .A1(n13593), .A2(n13109), .ZN(n13013) );
  AOI211_X1 U15198 ( .C1(n13058), .C2(n13415), .A(n13014), .B(n13013), .ZN(
        n13015) );
  OAI211_X1 U15199 ( .C1(n13018), .C2(n13017), .A(n13016), .B(n13015), .ZN(
        P2_U3188) );
  OAI211_X1 U15200 ( .C1(n13021), .C2(n13020), .A(n13019), .B(n14788), .ZN(
        n13029) );
  INV_X1 U15201 ( .A(n13022), .ZN(n13023) );
  AOI22_X1 U15202 ( .A1(n14534), .A2(n13023), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13028) );
  NAND2_X1 U15203 ( .A1(n14782), .A2(n13024), .ZN(n13027) );
  OR2_X1 U15204 ( .A1(n14797), .A2(n13025), .ZN(n13026) );
  NAND4_X1 U15205 ( .A1(n13029), .A2(n13028), .A3(n13027), .A4(n13026), .ZN(
        P2_U3189) );
  INV_X1 U15206 ( .A(n13030), .ZN(n13033) );
  NOR3_X1 U15207 ( .A1(n13031), .A2(n13303), .A3(n13110), .ZN(n13032) );
  AOI21_X1 U15208 ( .B1(n13033), .B2(n14788), .A(n13032), .ZN(n13039) );
  OAI22_X1 U15209 ( .A1(n13307), .A2(n13510), .B1(n13303), .B2(n13508), .ZN(
        n13617) );
  NAND2_X1 U15210 ( .A1(n13617), .A2(n14534), .ZN(n13034) );
  NAND2_X1 U15211 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13250)
         );
  OAI211_X1 U15212 ( .C1(n14797), .C2(n13465), .A(n13034), .B(n13250), .ZN(
        n13036) );
  NOR2_X1 U15213 ( .A1(n13086), .A2(n14777), .ZN(n13035) );
  AOI211_X1 U15214 ( .C1(n13618), .C2(n14794), .A(n13036), .B(n13035), .ZN(
        n13037) );
  OAI21_X1 U15215 ( .B1(n13039), .B2(n13038), .A(n13037), .ZN(P2_U3191) );
  AOI22_X1 U15216 ( .A1(n13125), .A2(n13254), .B1(n13116), .B2(n13309), .ZN(
        n13602) );
  INV_X1 U15217 ( .A(n13602), .ZN(n13040) );
  AOI22_X1 U15218 ( .A1(n13040), .A2(n14534), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13041) );
  OAI21_X1 U15219 ( .B1(n13442), .B2(n14797), .A(n13041), .ZN(n13047) );
  INV_X1 U15220 ( .A(n13042), .ZN(n13043) );
  AOI211_X1 U15221 ( .C1(n13045), .C2(n13044), .A(n14777), .B(n13043), .ZN(
        n13046) );
  AOI211_X1 U15222 ( .C1(n13439), .C2(n14782), .A(n13047), .B(n13046), .ZN(
        n13048) );
  INV_X1 U15223 ( .A(n13048), .ZN(P2_U3195) );
  INV_X1 U15224 ( .A(n6879), .ZN(n13389) );
  INV_X1 U15225 ( .A(n13050), .ZN(n13051) );
  AOI21_X1 U15226 ( .B1(n13049), .B2(n13051), .A(n14777), .ZN(n13055) );
  NOR3_X1 U15227 ( .A1(n13052), .A2(n13056), .A3(n13110), .ZN(n13054) );
  OAI21_X1 U15228 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13061) );
  INV_X1 U15229 ( .A(n13384), .ZN(n13059) );
  OAI22_X1 U15230 ( .A1(n13056), .A2(n13508), .B1(n13319), .B2(n13510), .ZN(
        n13581) );
  INV_X1 U15231 ( .A(n13581), .ZN(n13385) );
  INV_X1 U15232 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15213) );
  OAI22_X1 U15233 ( .A1(n14787), .A2(n13385), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15213), .ZN(n13057) );
  AOI21_X1 U15234 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n13060) );
  OAI211_X1 U15235 ( .C1(n13389), .C2(n13109), .A(n13061), .B(n13060), .ZN(
        P2_U3197) );
  NAND2_X1 U15236 ( .A1(n13128), .A2(n13254), .ZN(n13063) );
  NAND2_X1 U15237 ( .A1(n13130), .A2(n13116), .ZN(n13062) );
  NAND2_X1 U15238 ( .A1(n13063), .A2(n13062), .ZN(n13627) );
  AOI22_X1 U15239 ( .A1(n14534), .A2(n13627), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13064) );
  OAI21_X1 U15240 ( .B1(n14797), .B2(n13492), .A(n13064), .ZN(n13065) );
  AOI21_X1 U15241 ( .B1(n13628), .B2(n14794), .A(n13065), .ZN(n13070) );
  OAI22_X1 U15242 ( .A1(n13066), .A2(n14777), .B1(n13300), .B2(n13110), .ZN(
        n13067) );
  NAND3_X1 U15243 ( .A1(n14532), .A2(n13068), .A3(n13067), .ZN(n13069) );
  OAI211_X1 U15244 ( .C1(n6579), .C2(n14777), .A(n13070), .B(n13069), .ZN(
        P2_U3200) );
  INV_X1 U15245 ( .A(n13049), .ZN(n13082) );
  INV_X1 U15246 ( .A(n13071), .ZN(n13076) );
  INV_X1 U15247 ( .A(n13072), .ZN(n13073) );
  AOI21_X1 U15248 ( .B1(n13074), .B2(n13073), .A(n14777), .ZN(n13075) );
  AOI21_X1 U15249 ( .B1(n13077), .B2(n13076), .A(n13075), .ZN(n13081) );
  OAI22_X1 U15250 ( .A1(n7203), .A2(n13508), .B1(n13284), .B2(n13510), .ZN(
        n13393) );
  AOI22_X1 U15251 ( .A1(n13393), .A2(n14534), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13078) );
  OAI21_X1 U15252 ( .B1(n13397), .B2(n14797), .A(n13078), .ZN(n13079) );
  AOI21_X1 U15253 ( .B1(n13587), .B2(n14782), .A(n13079), .ZN(n13080) );
  OAI21_X1 U15254 ( .B1(n13082), .B2(n13081), .A(n13080), .ZN(P2_U3201) );
  INV_X1 U15255 ( .A(n13083), .ZN(n13452) );
  AOI22_X1 U15256 ( .A1(n13126), .A2(n13254), .B1(n13116), .B2(n13127), .ZN(
        n13609) );
  INV_X1 U15257 ( .A(n13609), .ZN(n13084) );
  AOI22_X1 U15258 ( .A1(n13084), .A2(n14534), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13085) );
  OAI21_X1 U15259 ( .B1(n13452), .B2(n14797), .A(n13085), .ZN(n13092) );
  INV_X1 U15260 ( .A(n13086), .ZN(n13090) );
  AOI22_X1 U15261 ( .A1(n13087), .A2(n14788), .B1(n13096), .B2(n13127), .ZN(
        n13089) );
  NOR3_X1 U15262 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(n13091) );
  AOI211_X1 U15263 ( .C1(n13449), .C2(n14794), .A(n13092), .B(n13091), .ZN(
        n13093) );
  OAI21_X1 U15264 ( .B1(n13094), .B2(n14777), .A(n13093), .ZN(P2_U3205) );
  AOI22_X1 U15265 ( .A1(n7125), .A2(n14788), .B1(n13096), .B2(n13125), .ZN(
        n13102) );
  INV_X1 U15266 ( .A(n13097), .ZN(n13101) );
  OAI22_X1 U15267 ( .A1(n7203), .A2(n13510), .B1(n13310), .B2(n13508), .ZN(
        n13422) );
  AOI22_X1 U15268 ( .A1(n13422), .A2(n14534), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13098) );
  OAI21_X1 U15269 ( .B1(n13427), .B2(n14797), .A(n13098), .ZN(n13099) );
  AOI21_X1 U15270 ( .B1(n13598), .B2(n14782), .A(n13099), .ZN(n13100) );
  OAI21_X1 U15271 ( .B1(n13102), .B2(n13101), .A(n13100), .ZN(P2_U3207) );
  INV_X1 U15272 ( .A(n13623), .ZN(n13483) );
  OAI211_X1 U15273 ( .C1(n13104), .C2(n13103), .A(n13030), .B(n14788), .ZN(
        n13108) );
  INV_X1 U15274 ( .A(n13127), .ZN(n13274) );
  OAI22_X1 U15275 ( .A1(n13274), .A2(n13510), .B1(n13511), .B2(n13508), .ZN(
        n13475) );
  NAND2_X1 U15276 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14921)
         );
  INV_X1 U15277 ( .A(n14921), .ZN(n13106) );
  NOR2_X1 U15278 ( .A1(n14797), .A2(n13480), .ZN(n13105) );
  AOI211_X1 U15279 ( .C1(n14534), .C2(n13475), .A(n13106), .B(n13105), .ZN(
        n13107) );
  OAI211_X1 U15280 ( .C1(n13483), .C2(n13109), .A(n13108), .B(n13107), .ZN(
        P2_U3210) );
  NOR2_X1 U15281 ( .A1(n13053), .A2(n14777), .ZN(n13115) );
  NOR3_X1 U15282 ( .A1(n13111), .A2(n13284), .A3(n13110), .ZN(n13114) );
  INV_X1 U15283 ( .A(n13112), .ZN(n13113) );
  OAI21_X1 U15284 ( .B1(n13115), .B2(n13114), .A(n13113), .ZN(n13121) );
  AOI22_X1 U15285 ( .A1(n13116), .A2(n13316), .B1(n13286), .B2(n13254), .ZN(
        n13572) );
  INV_X1 U15286 ( .A(n13572), .ZN(n13117) );
  AOI22_X1 U15287 ( .A1(n14534), .A2(n13117), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13118) );
  OAI21_X1 U15288 ( .B1(n14797), .B2(n13370), .A(n13118), .ZN(n13119) );
  AOI21_X1 U15289 ( .B1(n13373), .B2(n14794), .A(n13119), .ZN(n13120) );
  OAI211_X1 U15290 ( .C1(n14777), .C2(n13122), .A(n13121), .B(n13120), .ZN(
        P2_U3212) );
  CLKBUF_X2 U15291 ( .A(P2_U3947), .Z(n14773) );
  MUX2_X1 U15292 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13257), .S(n14773), .Z(
        P2_U3562) );
  MUX2_X1 U15293 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13290), .S(n14773), .Z(
        P2_U3561) );
  MUX2_X1 U15294 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13123), .S(n14773), .Z(
        P2_U3560) );
  MUX2_X1 U15295 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13124), .S(n14773), .Z(
        P2_U3559) );
  MUX2_X1 U15296 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13286), .S(n14773), .Z(
        P2_U3558) );
  MUX2_X1 U15297 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13318), .S(n14773), .Z(
        P2_U3557) );
  MUX2_X1 U15298 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13316), .S(n14773), .Z(
        P2_U3556) );
  MUX2_X1 U15299 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13314), .S(n14773), .Z(
        P2_U3555) );
  MUX2_X1 U15300 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13281), .S(n14773), .Z(
        P2_U3554) );
  MUX2_X1 U15301 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13125), .S(n14773), .Z(
        P2_U3553) );
  MUX2_X1 U15302 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13126), .S(n14773), .Z(
        P2_U3552) );
  MUX2_X1 U15303 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13309), .S(n14773), .Z(
        P2_U3551) );
  MUX2_X1 U15304 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13127), .S(n14773), .Z(
        P2_U3550) );
  MUX2_X1 U15305 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13128), .S(n14773), .Z(
        P2_U3549) );
  MUX2_X1 U15306 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13129), .S(n14773), .Z(
        P2_U3548) );
  MUX2_X1 U15307 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13130), .S(n14773), .Z(
        P2_U3547) );
  MUX2_X1 U15308 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13131), .S(n14773), .Z(
        P2_U3546) );
  MUX2_X1 U15309 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13132), .S(n14773), .Z(
        P2_U3545) );
  MUX2_X1 U15310 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13133), .S(n14773), .Z(
        P2_U3544) );
  MUX2_X1 U15311 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13134), .S(n14773), .Z(
        P2_U3543) );
  MUX2_X1 U15312 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13135), .S(n14773), .Z(
        P2_U3542) );
  MUX2_X1 U15313 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13136), .S(n14773), .Z(
        P2_U3541) );
  MUX2_X1 U15314 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13137), .S(n14773), .Z(
        P2_U3540) );
  MUX2_X1 U15315 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13138), .S(n14773), .Z(
        P2_U3539) );
  MUX2_X1 U15316 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13139), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15317 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13140), .S(n14773), .Z(
        P2_U3537) );
  MUX2_X1 U15318 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13141), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U15319 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13142), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15320 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13143), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15321 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13144), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U15322 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6413), .S(n14773), .Z(
        P2_U3532) );
  MUX2_X1 U15323 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13146), .S(n14773), .Z(
        P2_U3531) );
  INV_X1 U15324 ( .A(n14930), .ZN(n14906) );
  INV_X1 U15325 ( .A(n13151), .ZN(n13147) );
  AOI22_X1 U15326 ( .A1(n14906), .A2(n13147), .B1(n14923), .B2(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U15327 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(P2_U3088), .ZN(n13157) );
  OAI211_X1 U15328 ( .C1(n13150), .C2(n13149), .A(n14925), .B(n13148), .ZN(
        n13156) );
  MUX2_X1 U15329 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n13545), .S(n13151), .Z(
        n13152) );
  OAI21_X1 U15330 ( .B1(n9417), .B2(n6659), .A(n13152), .ZN(n13153) );
  NAND3_X1 U15331 ( .A1(n14917), .A2(n13154), .A3(n13153), .ZN(n13155) );
  NAND4_X1 U15332 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        P2_U3215) );
  INV_X1 U15333 ( .A(n13159), .ZN(n13160) );
  AOI22_X1 U15334 ( .A1(n14906), .A2(n13160), .B1(n14923), .B2(
        P2_ADDR_REG_2__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U15335 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n13167) );
  OAI211_X1 U15336 ( .C1(n13162), .C2(n13161), .A(n14917), .B(n13172), .ZN(
        n13166) );
  OAI211_X1 U15337 ( .C1(n13164), .C2(n13163), .A(n14925), .B(n13177), .ZN(
        n13165) );
  NAND4_X1 U15338 ( .A1(n13168), .A2(n13167), .A3(n13166), .A4(n13165), .ZN(
        P2_U3216) );
  AOI22_X1 U15339 ( .A1(n14906), .A2(n13169), .B1(n14923), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U15340 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13181) );
  MUX2_X1 U15341 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9333), .S(n13174), .Z(
        n13170) );
  NAND3_X1 U15342 ( .A1(n13172), .A2(n13171), .A3(n13170), .ZN(n13173) );
  NAND3_X1 U15343 ( .A1(n14917), .A2(n14801), .A3(n13173), .ZN(n13180) );
  MUX2_X1 U15344 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9355), .S(n13174), .Z(
        n13175) );
  NAND3_X1 U15345 ( .A1(n13177), .A2(n13176), .A3(n13175), .ZN(n13178) );
  NAND3_X1 U15346 ( .A1(n14925), .A2(n14805), .A3(n13178), .ZN(n13179) );
  NAND4_X1 U15347 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        P2_U3217) );
  AOI22_X1 U15348 ( .A1(n14906), .A2(n13183), .B1(n14923), .B2(
        P2_ADDR_REG_6__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U15349 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13195) );
  MUX2_X1 U15350 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9364), .S(n13188), .Z(
        n13184) );
  NAND3_X1 U15351 ( .A1(n14824), .A2(n13185), .A3(n13184), .ZN(n13186) );
  NAND3_X1 U15352 ( .A1(n14925), .A2(n13187), .A3(n13186), .ZN(n13194) );
  MUX2_X1 U15353 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9341), .S(n13188), .Z(
        n13189) );
  NAND3_X1 U15354 ( .A1(n14818), .A2(n13190), .A3(n13189), .ZN(n13191) );
  NAND3_X1 U15355 ( .A1(n14917), .A2(n13192), .A3(n13191), .ZN(n13193) );
  NAND4_X1 U15356 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n13193), .ZN(
        P2_U3220) );
  AOI21_X1 U15357 ( .B1(n14923), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n13197), .ZN(
        n13212) );
  MUX2_X1 U15358 ( .A(n10748), .B(P2_REG2_REG_8__SCAN_IN), .S(n13203), .Z(
        n13198) );
  NAND3_X1 U15359 ( .A1(n13200), .A2(n13199), .A3(n13198), .ZN(n13201) );
  NAND3_X1 U15360 ( .A1(n14917), .A2(n13202), .A3(n13201), .ZN(n13211) );
  NAND2_X1 U15361 ( .A1(n14906), .A2(n13203), .ZN(n13210) );
  MUX2_X1 U15362 ( .A(n9546), .B(P2_REG1_REG_8__SCAN_IN), .S(n13203), .Z(
        n13204) );
  NAND3_X1 U15363 ( .A1(n13206), .A2(n13205), .A3(n13204), .ZN(n13207) );
  NAND3_X1 U15364 ( .A1(n14925), .A2(n13208), .A3(n13207), .ZN(n13209) );
  NAND4_X1 U15365 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        P2_U3222) );
  INV_X1 U15366 ( .A(n14923), .ZN(n14846) );
  NAND2_X1 U15367 ( .A1(n14905), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13223) );
  INV_X1 U15368 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13214) );
  INV_X1 U15369 ( .A(n13223), .ZN(n13213) );
  AOI21_X1 U15370 ( .B1(n13214), .B2(n13237), .A(n13213), .ZN(n14912) );
  AOI22_X1 U15371 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n13235), .B1(n14904), 
        .B2(n13516), .ZN(n14901) );
  INV_X1 U15372 ( .A(n13215), .ZN(n13216) );
  OAI21_X1 U15373 ( .B1(n13217), .B2(n13228), .A(n13216), .ZN(n13218) );
  NAND2_X1 U15374 ( .A1(n14876), .A2(n13218), .ZN(n13220) );
  NAND2_X1 U15375 ( .A1(n13220), .A2(n14874), .ZN(n13221) );
  NAND2_X1 U15376 ( .A1(n13221), .A2(n14884), .ZN(n13222) );
  NAND2_X1 U15377 ( .A1(n13222), .A2(n14885), .ZN(n14900) );
  NAND2_X1 U15378 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  OAI21_X1 U15379 ( .B1(n14904), .B2(n13516), .A(n14899), .ZN(n14911) );
  NAND2_X1 U15380 ( .A1(n14912), .A2(n14911), .ZN(n14910) );
  NAND2_X1 U15381 ( .A1(n13223), .A2(n14910), .ZN(n13224) );
  NOR2_X1 U15382 ( .A1(n13239), .A2(n13224), .ZN(n13225) );
  XOR2_X1 U15383 ( .A(n14929), .B(n13224), .Z(n14918) );
  NOR2_X1 U15384 ( .A1(n13225), .A2(n14919), .ZN(n13226) );
  XOR2_X1 U15385 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13226), .Z(n13243) );
  XNOR2_X1 U15386 ( .A(n14905), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14907) );
  XNOR2_X1 U15387 ( .A(n14904), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14894) );
  OAI21_X1 U15388 ( .B1(n13229), .B2(n13228), .A(n13227), .ZN(n14877) );
  INV_X1 U15389 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13230) );
  XNOR2_X1 U15390 ( .A(n14876), .B(n13230), .ZN(n14878) );
  AOI22_X1 U15391 ( .A1(n14877), .A2(n14878), .B1(n14876), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n13232) );
  XNOR2_X1 U15392 ( .A(n13232), .B(n13231), .ZN(n14887) );
  OAI22_X1 U15393 ( .A1(n14887), .A2(n13233), .B1(n13232), .B2(n13231), .ZN(
        n14895) );
  NAND2_X1 U15394 ( .A1(n14894), .A2(n14895), .ZN(n14893) );
  INV_X1 U15395 ( .A(n14893), .ZN(n13234) );
  AOI21_X1 U15396 ( .B1(n13235), .B2(P2_REG1_REG_16__SCAN_IN), .A(n13234), 
        .ZN(n14908) );
  OAI22_X1 U15397 ( .A1(n14907), .A2(n14908), .B1(n13237), .B2(n13236), .ZN(
        n13238) );
  XNOR2_X1 U15398 ( .A(n13238), .B(n14929), .ZN(n14926) );
  NAND2_X1 U15399 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14926), .ZN(n14924) );
  NAND2_X1 U15400 ( .A1(n13239), .A2(n13238), .ZN(n13240) );
  NAND2_X1 U15401 ( .A1(n14924), .A2(n13240), .ZN(n13242) );
  INV_X1 U15402 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13241) );
  XNOR2_X1 U15403 ( .A(n13242), .B(n13241), .ZN(n13247) );
  AOI22_X1 U15404 ( .A1(n13243), .A2(n14917), .B1(n14925), .B2(n13247), .ZN(
        n13249) );
  INV_X1 U15405 ( .A(n13243), .ZN(n13244) );
  NAND2_X1 U15406 ( .A1(n14917), .A2(n13244), .ZN(n13245) );
  MUX2_X1 U15407 ( .A(n13249), .B(n13248), .S(n8318), .Z(n13251) );
  OAI211_X1 U15408 ( .C1(n14846), .C2(n13252), .A(n13251), .B(n13250), .ZN(
        P2_U3233) );
  OR2_X2 U15409 ( .A1(n13519), .A2(n14536), .ZN(n13520) );
  NAND2_X1 U15410 ( .A1(n13498), .A2(n13483), .ZN(n13485) );
  NOR2_X2 U15411 ( .A1(n6879), .A2(n13400), .ZN(n13383) );
  NAND2_X1 U15412 ( .A1(n13574), .A2(n13383), .ZN(n13368) );
  OAI21_X1 U15413 ( .B1(n9094), .B2(n13255), .A(n13254), .ZN(n13291) );
  INV_X1 U15414 ( .A(n13291), .ZN(n13256) );
  NAND2_X1 U15415 ( .A1(n13257), .A2(n13256), .ZN(n13550) );
  NOR2_X1 U15416 ( .A1(n14943), .A2(n13550), .ZN(n13262) );
  NOR2_X1 U15417 ( .A1(n6769), .A2(n13533), .ZN(n13258) );
  AOI211_X1 U15418 ( .C1(n14943), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13262), 
        .B(n13258), .ZN(n13259) );
  OAI21_X1 U15419 ( .B1(n13549), .B2(n13500), .A(n13259), .ZN(P2_U3234) );
  OAI211_X1 U15420 ( .C1(n13552), .C2(n13328), .A(n13496), .B(n13260), .ZN(
        n13551) );
  NOR2_X1 U15421 ( .A1(n13552), .A2(n13533), .ZN(n13261) );
  AOI211_X1 U15422 ( .C1(n14943), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13262), 
        .B(n13261), .ZN(n13263) );
  OAI21_X1 U15423 ( .B1(n13500), .B2(n13551), .A(n13263), .ZN(P2_U3235) );
  OR2_X1 U15424 ( .A1(n13640), .A2(n13509), .ZN(n13265) );
  NAND2_X1 U15425 ( .A1(n13266), .A2(n13265), .ZN(n13507) );
  INV_X1 U15426 ( .A(n13514), .ZN(n13267) );
  NAND2_X1 U15427 ( .A1(n13507), .A2(n13267), .ZN(n13269) );
  OR2_X1 U15428 ( .A1(n14536), .A2(n13300), .ZN(n13268) );
  NAND2_X1 U15429 ( .A1(n13269), .A2(n13268), .ZN(n13504) );
  NOR2_X1 U15430 ( .A1(n13628), .A2(n13511), .ZN(n13271) );
  NAND2_X1 U15431 ( .A1(n13628), .A2(n13511), .ZN(n13270) );
  AND2_X1 U15432 ( .A1(n13623), .A2(n13303), .ZN(n13272) );
  OR2_X1 U15433 ( .A1(n13623), .A2(n13303), .ZN(n13273) );
  NOR2_X1 U15434 ( .A1(n13618), .A2(n13274), .ZN(n13275) );
  NAND2_X1 U15435 ( .A1(n13458), .A2(n13457), .ZN(n13278) );
  NAND2_X1 U15436 ( .A1(n13449), .A2(n13307), .ZN(n13277) );
  NAND2_X1 U15437 ( .A1(n13278), .A2(n13277), .ZN(n13436) );
  AND2_X1 U15438 ( .A1(n13439), .A2(n13310), .ZN(n13279) );
  INV_X1 U15439 ( .A(n13425), .ZN(n13280) );
  AOI21_X1 U15440 ( .B1(n7203), .B2(n13410), .A(n13282), .ZN(n13392) );
  INV_X1 U15441 ( .A(n13587), .ZN(n13283) );
  INV_X1 U15442 ( .A(n13379), .ZN(n13285) );
  INV_X1 U15443 ( .A(n13286), .ZN(n13322) );
  INV_X1 U15444 ( .A(n15057), .ZN(n13288) );
  INV_X1 U15445 ( .A(n13290), .ZN(n13292) );
  AOI21_X1 U15446 ( .B1(n13124), .B2(n13116), .A(n13293), .ZN(n13294) );
  INV_X1 U15447 ( .A(n13568), .ZN(n13361) );
  INV_X1 U15448 ( .A(n13295), .ZN(n13297) );
  NAND2_X1 U15449 ( .A1(n13515), .A2(n13514), .ZN(n13513) );
  INV_X1 U15450 ( .A(n13628), .ZN(n13301) );
  INV_X1 U15451 ( .A(n13304), .ZN(n13306) );
  NAND2_X1 U15452 ( .A1(n13426), .A2(n13425), .ZN(n13424) );
  NAND2_X1 U15453 ( .A1(n13389), .A2(n13284), .ZN(n13317) );
  NAND2_X1 U15454 ( .A1(n13373), .A2(n13318), .ZN(n13320) );
  NAND2_X1 U15455 ( .A1(n13340), .A2(n13324), .ZN(n13327) );
  XNOR2_X1 U15456 ( .A(n13327), .B(n13326), .ZN(n13553) );
  INV_X1 U15457 ( .A(n13555), .ZN(n13333) );
  AOI211_X1 U15458 ( .C1(n13555), .C2(n13343), .A(n13529), .B(n13328), .ZN(
        n13554) );
  NAND2_X1 U15459 ( .A1(n13554), .A2(n13535), .ZN(n13332) );
  INV_X1 U15460 ( .A(n13329), .ZN(n13330) );
  AOI22_X1 U15461 ( .A1(n14943), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13330), 
        .B2(n13493), .ZN(n13331) );
  OAI211_X1 U15462 ( .C1(n13333), .C2(n13533), .A(n13332), .B(n13331), .ZN(
        n13334) );
  AOI21_X1 U15463 ( .B1(n13553), .B2(n13542), .A(n13334), .ZN(n13335) );
  OAI21_X1 U15464 ( .B1(n6406), .B2(n14943), .A(n13335), .ZN(P2_U3236) );
  AOI21_X1 U15465 ( .B1(n7208), .B2(n13341), .A(n15057), .ZN(n13339) );
  AOI21_X1 U15466 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n13562) );
  OAI21_X1 U15467 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n13557) );
  INV_X1 U15468 ( .A(n13557), .ZN(n13350) );
  AOI21_X1 U15469 ( .B1(n13558), .B2(n13355), .A(n10303), .ZN(n13344) );
  NAND2_X1 U15470 ( .A1(n13344), .A2(n13343), .ZN(n13560) );
  OAI22_X1 U15471 ( .A1(n13543), .A2(n13346), .B1(n13345), .B2(n14938), .ZN(
        n13347) );
  AOI21_X1 U15472 ( .B1(n13558), .B2(n13518), .A(n13347), .ZN(n13348) );
  OAI21_X1 U15473 ( .B1(n13560), .B2(n13500), .A(n13348), .ZN(n13349) );
  AOI21_X1 U15474 ( .B1(n13350), .B2(n13542), .A(n13349), .ZN(n13351) );
  OAI21_X1 U15475 ( .B1(n14943), .B2(n13562), .A(n13351), .ZN(P2_U3237) );
  XNOR2_X1 U15476 ( .A(n13352), .B(n13353), .ZN(n13571) );
  OR2_X1 U15477 ( .A1(n13354), .A2(n13353), .ZN(n13565) );
  NAND3_X1 U15478 ( .A1(n13565), .A2(n13564), .A3(n13542), .ZN(n13364) );
  AOI21_X1 U15479 ( .B1(n13568), .B2(n13368), .A(n10303), .ZN(n13356) );
  INV_X1 U15480 ( .A(n13567), .ZN(n13358) );
  OAI22_X1 U15481 ( .A1(n14943), .A2(n13358), .B1(n13357), .B2(n14938), .ZN(
        n13359) );
  AOI21_X1 U15482 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(n14943), .A(n13359), 
        .ZN(n13360) );
  OAI21_X1 U15483 ( .B1(n13361), .B2(n13533), .A(n13360), .ZN(n13362) );
  AOI21_X1 U15484 ( .B1(n13535), .B2(n13566), .A(n13362), .ZN(n13363) );
  OAI211_X1 U15485 ( .C1(n13571), .C2(n13473), .A(n13364), .B(n13363), .ZN(
        P2_U3238) );
  XNOR2_X1 U15486 ( .A(n13365), .B(n7216), .ZN(n13578) );
  XNOR2_X1 U15487 ( .A(n13367), .B(n13366), .ZN(n13576) );
  OAI211_X1 U15488 ( .C1(n13574), .C2(n13383), .A(n13496), .B(n13368), .ZN(
        n13573) );
  NOR2_X1 U15489 ( .A1(n13543), .A2(n13369), .ZN(n13372) );
  OAI22_X1 U15490 ( .A1(n14943), .A2(n13572), .B1(n13370), .B2(n14938), .ZN(
        n13371) );
  AOI211_X1 U15491 ( .C1(n13373), .C2(n13518), .A(n13372), .B(n13371), .ZN(
        n13374) );
  OAI21_X1 U15492 ( .B1(n13573), .B2(n13500), .A(n13374), .ZN(n13375) );
  AOI21_X1 U15493 ( .B1(n13576), .B2(n13541), .A(n13375), .ZN(n13376) );
  OAI21_X1 U15494 ( .B1(n13578), .B2(n13524), .A(n13376), .ZN(P2_U3239) );
  XNOR2_X1 U15495 ( .A(n13377), .B(n13379), .ZN(n13585) );
  OAI21_X1 U15496 ( .B1(n13380), .B2(n13379), .A(n13378), .ZN(n13579) );
  NAND2_X1 U15497 ( .A1(n6879), .A2(n13400), .ZN(n13381) );
  NAND2_X1 U15498 ( .A1(n13381), .A2(n13496), .ZN(n13382) );
  NOR2_X1 U15499 ( .A1(n13383), .A2(n13382), .ZN(n13580) );
  NAND2_X1 U15500 ( .A1(n13580), .A2(n13535), .ZN(n13388) );
  OAI22_X1 U15501 ( .A1(n14943), .A2(n13385), .B1(n13384), .B2(n14938), .ZN(
        n13386) );
  AOI21_X1 U15502 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(n14943), .A(n13386), 
        .ZN(n13387) );
  OAI211_X1 U15503 ( .C1(n13389), .C2(n13533), .A(n13388), .B(n13387), .ZN(
        n13390) );
  AOI21_X1 U15504 ( .B1(n13579), .B2(n13542), .A(n13390), .ZN(n13391) );
  OAI21_X1 U15505 ( .B1(n13585), .B2(n13473), .A(n13391), .ZN(P2_U3240) );
  XNOR2_X1 U15506 ( .A(n13392), .B(n13395), .ZN(n13394) );
  AOI21_X1 U15507 ( .B1(n13394), .B2(n15026), .A(n13393), .ZN(n13589) );
  XNOR2_X1 U15508 ( .A(n13396), .B(n13395), .ZN(n13590) );
  OAI22_X1 U15509 ( .A1(n14941), .A2(n13398), .B1(n13397), .B2(n14938), .ZN(
        n13399) );
  AOI21_X1 U15510 ( .B1(n13587), .B2(n13518), .A(n13399), .ZN(n13403) );
  AOI21_X1 U15511 ( .B1(n13587), .B2(n13412), .A(n10303), .ZN(n13401) );
  AND2_X1 U15512 ( .A1(n13401), .A2(n13400), .ZN(n13586) );
  NAND2_X1 U15513 ( .A1(n13586), .A2(n13535), .ZN(n13402) );
  OAI211_X1 U15514 ( .C1(n13590), .C2(n13524), .A(n13403), .B(n13402), .ZN(
        n13404) );
  INV_X1 U15515 ( .A(n13404), .ZN(n13405) );
  OAI21_X1 U15516 ( .B1(n14943), .B2(n13589), .A(n13405), .ZN(P2_U3241) );
  XNOR2_X1 U15517 ( .A(n13406), .B(n13408), .ZN(n13407) );
  NAND2_X1 U15518 ( .A1(n13407), .A2(n15026), .ZN(n13592) );
  XOR2_X1 U15519 ( .A(n13409), .B(n13408), .Z(n13595) );
  NAND2_X1 U15520 ( .A1(n13595), .A2(n13542), .ZN(n13420) );
  NAND2_X1 U15521 ( .A1(n13410), .A2(n13430), .ZN(n13411) );
  NAND3_X1 U15522 ( .A1(n13412), .A2(n13496), .A3(n13411), .ZN(n13414) );
  AND2_X1 U15523 ( .A1(n13414), .A2(n13413), .ZN(n13591) );
  INV_X1 U15524 ( .A(n13591), .ZN(n13418) );
  AOI22_X1 U15525 ( .A1(n14943), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13415), 
        .B2(n13493), .ZN(n13416) );
  OAI21_X1 U15526 ( .B1(n13593), .B2(n13533), .A(n13416), .ZN(n13417) );
  AOI21_X1 U15527 ( .B1(n13418), .B2(n13535), .A(n13417), .ZN(n13419) );
  OAI211_X1 U15528 ( .C1(n14943), .C2(n13592), .A(n13420), .B(n13419), .ZN(
        P2_U3242) );
  XNOR2_X1 U15529 ( .A(n13421), .B(n13425), .ZN(n13423) );
  AOI21_X1 U15530 ( .B1(n13423), .B2(n15026), .A(n13422), .ZN(n13600) );
  OAI21_X1 U15531 ( .B1(n13426), .B2(n13425), .A(n13424), .ZN(n13601) );
  INV_X1 U15532 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13428) );
  OAI22_X1 U15533 ( .A1(n13543), .A2(n13428), .B1(n13427), .B2(n14938), .ZN(
        n13429) );
  AOI21_X1 U15534 ( .B1(n13598), .B2(n13518), .A(n13429), .ZN(n13433) );
  AOI21_X1 U15535 ( .B1(n13598), .B2(n13440), .A(n10303), .ZN(n13431) );
  AND2_X1 U15536 ( .A1(n13431), .A2(n13430), .ZN(n13597) );
  NAND2_X1 U15537 ( .A1(n13597), .A2(n13535), .ZN(n13432) );
  OAI211_X1 U15538 ( .C1(n13601), .C2(n13524), .A(n13433), .B(n13432), .ZN(
        n13434) );
  INV_X1 U15539 ( .A(n13434), .ZN(n13435) );
  OAI21_X1 U15540 ( .B1(n14943), .B2(n13600), .A(n13435), .ZN(P2_U3243) );
  XNOR2_X1 U15541 ( .A(n13436), .B(n13437), .ZN(n13608) );
  XNOR2_X1 U15542 ( .A(n13438), .B(n13437), .ZN(n13606) );
  AOI21_X1 U15543 ( .B1(n13439), .B2(n13450), .A(n10303), .ZN(n13441) );
  NAND2_X1 U15544 ( .A1(n13441), .A2(n13440), .ZN(n13603) );
  OAI22_X1 U15545 ( .A1(n13602), .A2(n14943), .B1(n13442), .B2(n14938), .ZN(
        n13444) );
  NOR2_X1 U15546 ( .A1(n13604), .A2(n13533), .ZN(n13443) );
  AOI211_X1 U15547 ( .C1(n14943), .C2(P2_REG2_REG_21__SCAN_IN), .A(n13444), 
        .B(n13443), .ZN(n13445) );
  OAI21_X1 U15548 ( .B1(n13500), .B2(n13603), .A(n13445), .ZN(n13446) );
  AOI21_X1 U15549 ( .B1(n13606), .B2(n13542), .A(n13446), .ZN(n13447) );
  OAI21_X1 U15550 ( .B1(n13608), .B2(n13473), .A(n13447), .ZN(P2_U3244) );
  XNOR2_X1 U15551 ( .A(n13448), .B(n13457), .ZN(n13614) );
  AOI21_X1 U15552 ( .B1(n13449), .B2(n13464), .A(n10303), .ZN(n13451) );
  NAND2_X1 U15553 ( .A1(n13451), .A2(n13450), .ZN(n13610) );
  INV_X1 U15554 ( .A(n13610), .ZN(n13456) );
  OAI22_X1 U15555 ( .A1(n13609), .A2(n14943), .B1(n13452), .B2(n14938), .ZN(
        n13453) );
  AOI21_X1 U15556 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(n14943), .A(n13453), 
        .ZN(n13454) );
  OAI21_X1 U15557 ( .B1(n6770), .B2(n13533), .A(n13454), .ZN(n13455) );
  AOI21_X1 U15558 ( .B1(n13456), .B2(n13535), .A(n13455), .ZN(n13460) );
  XNOR2_X1 U15559 ( .A(n13458), .B(n13457), .ZN(n13612) );
  NAND2_X1 U15560 ( .A1(n13612), .A2(n13541), .ZN(n13459) );
  OAI211_X1 U15561 ( .C1(n13614), .C2(n13524), .A(n13460), .B(n13459), .ZN(
        P2_U3245) );
  XNOR2_X1 U15562 ( .A(n13461), .B(n13462), .ZN(n13621) );
  XNOR2_X1 U15563 ( .A(n13463), .B(n13462), .ZN(n13615) );
  NAND2_X1 U15564 ( .A1(n13615), .A2(n13542), .ZN(n13472) );
  AOI211_X1 U15565 ( .C1(n13618), .C2(n13485), .A(n13529), .B(n6771), .ZN(
        n13616) );
  NAND2_X1 U15566 ( .A1(n13618), .A2(n13518), .ZN(n13468) );
  INV_X1 U15567 ( .A(n13465), .ZN(n13466) );
  AOI22_X1 U15568 ( .A1(n13617), .A2(n13543), .B1(n13466), .B2(n13493), .ZN(
        n13467) );
  OAI211_X1 U15569 ( .C1(n14941), .C2(n13469), .A(n13468), .B(n13467), .ZN(
        n13470) );
  AOI21_X1 U15570 ( .B1(n13616), .B2(n13535), .A(n13470), .ZN(n13471) );
  OAI211_X1 U15571 ( .C1(n13621), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        P2_U3246) );
  XNOR2_X1 U15572 ( .A(n13474), .B(n13479), .ZN(n13476) );
  AOI21_X1 U15573 ( .B1(n13476), .B2(n15026), .A(n13475), .ZN(n13625) );
  AOI21_X1 U15574 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n13626) );
  OAI22_X1 U15575 ( .A1(n14941), .A2(n13481), .B1(n13480), .B2(n14938), .ZN(
        n13482) );
  AOI21_X1 U15576 ( .B1(n13623), .B2(n13518), .A(n13482), .ZN(n13487) );
  OR2_X1 U15577 ( .A1(n13498), .A2(n13483), .ZN(n13484) );
  AND3_X1 U15578 ( .A1(n13485), .A2(n13496), .A3(n13484), .ZN(n13622) );
  NAND2_X1 U15579 ( .A1(n13622), .A2(n13535), .ZN(n13486) );
  OAI211_X1 U15580 ( .C1(n13626), .C2(n13524), .A(n13487), .B(n13486), .ZN(
        n13488) );
  INV_X1 U15581 ( .A(n13488), .ZN(n13489) );
  OAI21_X1 U15582 ( .B1(n14943), .B2(n13625), .A(n13489), .ZN(P2_U3247) );
  OAI21_X1 U15583 ( .B1(n13491), .B2(n13503), .A(n13490), .ZN(n13631) );
  INV_X1 U15584 ( .A(n13492), .ZN(n13494) );
  AOI22_X1 U15585 ( .A1(n13543), .A2(n13627), .B1(n13494), .B2(n13493), .ZN(
        n13495) );
  OAI21_X1 U15586 ( .B1(n13214), .B2(n14941), .A(n13495), .ZN(n13502) );
  NAND2_X1 U15587 ( .A1(n13520), .A2(n13628), .ZN(n13497) );
  NAND2_X1 U15588 ( .A1(n13497), .A2(n13496), .ZN(n13499) );
  OR2_X1 U15589 ( .A1(n13499), .A2(n13498), .ZN(n13629) );
  NOR2_X1 U15590 ( .A1(n13629), .A2(n13500), .ZN(n13501) );
  AOI211_X1 U15591 ( .C1(n13518), .C2(n13628), .A(n13502), .B(n13501), .ZN(
        n13506) );
  XNOR2_X1 U15592 ( .A(n13504), .B(n13503), .ZN(n13633) );
  NAND2_X1 U15593 ( .A1(n13633), .A2(n13541), .ZN(n13505) );
  OAI211_X1 U15594 ( .C1(n13631), .C2(n13524), .A(n13506), .B(n13505), .ZN(
        P2_U3248) );
  XNOR2_X1 U15595 ( .A(n13507), .B(n13514), .ZN(n13512) );
  OAI22_X1 U15596 ( .A1(n13511), .A2(n13510), .B1(n13509), .B2(n13508), .ZN(
        n14535) );
  AOI21_X1 U15597 ( .B1(n13512), .B2(n15026), .A(n14535), .ZN(n13637) );
  OAI21_X1 U15598 ( .B1(n13515), .B2(n13514), .A(n13513), .ZN(n13638) );
  OAI22_X1 U15599 ( .A1(n13543), .A2(n13516), .B1(n14538), .B2(n14938), .ZN(
        n13517) );
  AOI21_X1 U15600 ( .B1(n14536), .B2(n13518), .A(n13517), .ZN(n13523) );
  AOI21_X1 U15601 ( .B1(n13519), .B2(n14536), .A(n10303), .ZN(n13521) );
  AND2_X1 U15602 ( .A1(n13521), .A2(n13520), .ZN(n13635) );
  NAND2_X1 U15603 ( .A1(n13635), .A2(n13535), .ZN(n13522) );
  OAI211_X1 U15604 ( .C1(n13638), .C2(n13524), .A(n13523), .B(n13522), .ZN(
        n13525) );
  INV_X1 U15605 ( .A(n13525), .ZN(n13526) );
  OAI21_X1 U15606 ( .B1(n14943), .B2(n13637), .A(n13526), .ZN(P2_U3249) );
  INV_X1 U15607 ( .A(n13527), .ZN(n13528) );
  AOI211_X1 U15608 ( .C1(n13530), .C2(n9053), .A(n13529), .B(n13528), .ZN(
        n14981) );
  OAI22_X1 U15609 ( .A1(n13533), .A2(n13532), .B1(n14938), .B2(n13531), .ZN(
        n13534) );
  AOI21_X1 U15610 ( .B1(n13535), .B2(n14981), .A(n13534), .ZN(n13548) );
  OAI21_X1 U15611 ( .B1(n13538), .B2(n13537), .A(n13536), .ZN(n14983) );
  XNOR2_X1 U15612 ( .A(n13540), .B(n13539), .ZN(n14988) );
  AOI22_X1 U15613 ( .A1(n13542), .A2(n14983), .B1(n13541), .B2(n14988), .ZN(
        n13547) );
  MUX2_X1 U15614 ( .A(n13545), .B(n13544), .S(n13543), .Z(n13546) );
  NAND3_X1 U15615 ( .A1(n13548), .A2(n13547), .A3(n13546), .ZN(P2_U3264) );
  OAI211_X1 U15616 ( .C1(n6769), .C2(n15046), .A(n13549), .B(n13550), .ZN(
        n13651) );
  MUX2_X1 U15617 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13651), .S(n15081), .Z(
        P2_U3530) );
  OAI211_X1 U15618 ( .C1(n13552), .C2(n15046), .A(n13551), .B(n13550), .ZN(
        n13652) );
  MUX2_X1 U15619 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13652), .S(n15081), .Z(
        P2_U3529) );
  NAND2_X1 U15620 ( .A1(n13553), .A2(n14999), .ZN(n13556) );
  MUX2_X1 U15621 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13653), .S(n15081), .Z(
        P2_U3528) );
  NAND2_X1 U15622 ( .A1(n13558), .A2(n15053), .ZN(n13559) );
  MUX2_X1 U15623 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13654), .S(n15081), .Z(
        P2_U3527) );
  NAND3_X1 U15624 ( .A1(n13565), .A2(n13564), .A3(n14999), .ZN(n13570) );
  AOI211_X1 U15625 ( .C1(n15053), .C2(n13568), .A(n13567), .B(n13566), .ZN(
        n13569) );
  OAI211_X1 U15626 ( .C1(n15057), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        n13655) );
  MUX2_X1 U15627 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13655), .S(n15081), .Z(
        P2_U3526) );
  OAI211_X1 U15628 ( .C1(n13574), .C2(n15046), .A(n13573), .B(n13572), .ZN(
        n13575) );
  AOI21_X1 U15629 ( .B1(n13576), .B2(n15026), .A(n13575), .ZN(n13577) );
  OAI21_X1 U15630 ( .B1(n13578), .B2(n15022), .A(n13577), .ZN(n13656) );
  MUX2_X1 U15631 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13656), .S(n15081), .Z(
        P2_U3525) );
  NAND2_X1 U15632 ( .A1(n13579), .A2(n14999), .ZN(n13584) );
  AOI211_X1 U15633 ( .C1(n15053), .C2(n6879), .A(n13581), .B(n13580), .ZN(
        n13583) );
  OAI211_X1 U15634 ( .C1(n15057), .C2(n13585), .A(n13584), .B(n13583), .ZN(
        n13657) );
  MUX2_X1 U15635 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13657), .S(n15081), .Z(
        P2_U3524) );
  AOI21_X1 U15636 ( .B1(n15053), .B2(n13587), .A(n13586), .ZN(n13588) );
  OAI211_X1 U15637 ( .C1(n13590), .C2(n15022), .A(n13589), .B(n13588), .ZN(
        n13658) );
  MUX2_X1 U15638 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13658), .S(n15081), .Z(
        P2_U3523) );
  OAI211_X1 U15639 ( .C1(n13593), .C2(n15046), .A(n13592), .B(n13591), .ZN(
        n13594) );
  AOI21_X1 U15640 ( .B1(n13595), .B2(n14999), .A(n13594), .ZN(n13596) );
  INV_X1 U15641 ( .A(n13596), .ZN(n13659) );
  MUX2_X1 U15642 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13659), .S(n15081), .Z(
        P2_U3522) );
  AOI21_X1 U15643 ( .B1(n15053), .B2(n13598), .A(n13597), .ZN(n13599) );
  OAI211_X1 U15644 ( .C1(n13601), .C2(n15022), .A(n13600), .B(n13599), .ZN(
        n13660) );
  MUX2_X1 U15645 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13660), .S(n15081), .Z(
        P2_U3521) );
  OAI211_X1 U15646 ( .C1(n13604), .C2(n15046), .A(n13603), .B(n13602), .ZN(
        n13605) );
  AOI21_X1 U15647 ( .B1(n13606), .B2(n14999), .A(n13605), .ZN(n13607) );
  OAI21_X1 U15648 ( .B1(n15057), .B2(n13608), .A(n13607), .ZN(n13661) );
  MUX2_X1 U15649 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13661), .S(n15081), .Z(
        P2_U3520) );
  OAI211_X1 U15650 ( .C1(n6770), .C2(n15046), .A(n13610), .B(n13609), .ZN(
        n13611) );
  AOI21_X1 U15651 ( .B1(n13612), .B2(n15026), .A(n13611), .ZN(n13613) );
  OAI21_X1 U15652 ( .B1(n13614), .B2(n15022), .A(n13613), .ZN(n13662) );
  MUX2_X1 U15653 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13662), .S(n15081), .Z(
        P2_U3519) );
  NAND2_X1 U15654 ( .A1(n13615), .A2(n14999), .ZN(n13620) );
  AOI211_X1 U15655 ( .C1(n15053), .C2(n13618), .A(n13617), .B(n13616), .ZN(
        n13619) );
  OAI211_X1 U15656 ( .C1(n15057), .C2(n13621), .A(n13620), .B(n13619), .ZN(
        n13663) );
  MUX2_X1 U15657 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13663), .S(n15081), .Z(
        P2_U3518) );
  AOI21_X1 U15658 ( .B1(n15053), .B2(n13623), .A(n13622), .ZN(n13624) );
  OAI211_X1 U15659 ( .C1(n13626), .C2(n15022), .A(n13625), .B(n13624), .ZN(
        n13664) );
  MUX2_X1 U15660 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13664), .S(n15081), .Z(
        P2_U3517) );
  AOI21_X1 U15661 ( .B1(n13628), .B2(n15053), .A(n13627), .ZN(n13630) );
  OAI211_X1 U15662 ( .C1(n13631), .C2(n15022), .A(n13630), .B(n13629), .ZN(
        n13632) );
  AOI21_X1 U15663 ( .B1(n13633), .B2(n15026), .A(n13632), .ZN(n13634) );
  INV_X1 U15664 ( .A(n13634), .ZN(n13665) );
  MUX2_X1 U15665 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13665), .S(n15081), .Z(
        P2_U3516) );
  AOI21_X1 U15666 ( .B1(n15053), .B2(n14536), .A(n13635), .ZN(n13636) );
  OAI211_X1 U15667 ( .C1(n13638), .C2(n15022), .A(n13637), .B(n13636), .ZN(
        n13666) );
  MUX2_X1 U15668 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13666), .S(n15081), .Z(
        P2_U3515) );
  AOI21_X1 U15669 ( .B1(n15053), .B2(n13640), .A(n13639), .ZN(n13641) );
  OAI211_X1 U15670 ( .C1(n13643), .C2(n15022), .A(n13642), .B(n13641), .ZN(
        n13667) );
  MUX2_X1 U15671 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13667), .S(n15081), .Z(
        P2_U3514) );
  OAI211_X1 U15672 ( .C1(n13646), .C2(n15046), .A(n13645), .B(n13644), .ZN(
        n13647) );
  AOI21_X1 U15673 ( .B1(n13648), .B2(n15026), .A(n13647), .ZN(n13649) );
  OAI21_X1 U15674 ( .B1(n13650), .B2(n15022), .A(n13649), .ZN(n13668) );
  MUX2_X1 U15675 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13668), .S(n15081), .Z(
        P2_U3513) );
  MUX2_X1 U15676 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13651), .S(n15066), .Z(
        P2_U3498) );
  MUX2_X1 U15677 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13652), .S(n15066), .Z(
        P2_U3497) );
  MUX2_X1 U15678 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13653), .S(n15066), .Z(
        P2_U3496) );
  MUX2_X1 U15679 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13654), .S(n15066), .Z(
        P2_U3495) );
  MUX2_X1 U15680 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13655), .S(n15066), .Z(
        P2_U3494) );
  MUX2_X1 U15681 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13656), .S(n15066), .Z(
        P2_U3493) );
  MUX2_X1 U15682 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13657), .S(n15066), .Z(
        P2_U3492) );
  MUX2_X1 U15683 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13658), .S(n15066), .Z(
        P2_U3491) );
  MUX2_X1 U15684 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13659), .S(n15066), .Z(
        P2_U3490) );
  MUX2_X1 U15685 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13660), .S(n15066), .Z(
        P2_U3489) );
  MUX2_X1 U15686 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13661), .S(n15066), .Z(
        P2_U3488) );
  MUX2_X1 U15687 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13662), .S(n15066), .Z(
        P2_U3487) );
  MUX2_X1 U15688 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13663), .S(n15066), .Z(
        P2_U3486) );
  MUX2_X1 U15689 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13664), .S(n15066), .Z(
        P2_U3484) );
  MUX2_X1 U15690 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13665), .S(n15066), .Z(
        P2_U3481) );
  MUX2_X1 U15691 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13666), .S(n15066), .Z(
        P2_U3478) );
  MUX2_X1 U15692 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13667), .S(n15066), .Z(
        P2_U3475) );
  MUX2_X1 U15693 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13668), .S(n15066), .Z(
        P2_U3472) );
  INV_X1 U15694 ( .A(n13669), .ZN(n13674) );
  NOR4_X1 U15695 ( .A1(n13670), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13671), .A4(
        P2_U3088), .ZN(n13672) );
  AOI21_X1 U15696 ( .B1(n13683), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13672), 
        .ZN(n13673) );
  OAI21_X1 U15697 ( .B1(n13674), .B2(n13688), .A(n13673), .ZN(P2_U3296) );
  INV_X1 U15698 ( .A(n13675), .ZN(n14313) );
  OAI222_X1 U15699 ( .A1(n13686), .A2(n13677), .B1(P2_U3088), .B2(n13676), 
        .C1(n13688), .C2(n14313), .ZN(P2_U3298) );
  INV_X1 U15700 ( .A(n13678), .ZN(n14316) );
  AOI21_X1 U15701 ( .B1(n13683), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13679), 
        .ZN(n13680) );
  OAI21_X1 U15702 ( .B1(n14316), .B2(n13688), .A(n13680), .ZN(P2_U3299) );
  INV_X1 U15703 ( .A(n13681), .ZN(n14319) );
  AOI21_X1 U15704 ( .B1(n13683), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n13682), 
        .ZN(n13684) );
  OAI21_X1 U15705 ( .B1(n14319), .B2(n13688), .A(n13684), .ZN(P2_U3300) );
  INV_X1 U15706 ( .A(n13685), .ZN(n14322) );
  OAI222_X1 U15707 ( .A1(n13689), .A2(P2_U3088), .B1(n13688), .B2(n14322), 
        .C1(n13687), .C2(n13686), .ZN(P2_U3301) );
  MUX2_X1 U15708 ( .A(n13690), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15709 ( .A(n13692), .B(n13691), .Z(n13697) );
  NOR2_X1 U15710 ( .A1(n14568), .A2(n14023), .ZN(n13695) );
  AOI22_X1 U15711 ( .A1(n13794), .A2(n14020), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13693) );
  OAI21_X1 U15712 ( .B1(n13960), .B2(n14551), .A(n13693), .ZN(n13694) );
  AOI211_X1 U15713 ( .C1(n14026), .C2(n14564), .A(n13695), .B(n13694), .ZN(
        n13696) );
  OAI21_X1 U15714 ( .B1(n13697), .B2(n14559), .A(n13696), .ZN(P1_U3214) );
  XOR2_X1 U15715 ( .A(n13699), .B(n13698), .Z(n13705) );
  NAND2_X1 U15716 ( .A1(n13985), .A2(n14572), .ZN(n13701) );
  NAND2_X1 U15717 ( .A1(n13988), .A2(n14575), .ZN(n13700) );
  NAND2_X1 U15718 ( .A1(n13701), .A2(n13700), .ZN(n14231) );
  AOI22_X1 U15719 ( .A1(n14231), .A2(n13805), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13702) );
  OAI21_X1 U15720 ( .B1(n14085), .B2(n14568), .A(n13702), .ZN(n13703) );
  AOI21_X1 U15721 ( .B1(n14232), .B2(n14564), .A(n13703), .ZN(n13704) );
  OAI21_X1 U15722 ( .B1(n13705), .B2(n14559), .A(n13704), .ZN(P1_U3216) );
  AOI21_X1 U15723 ( .B1(n13707), .B2(n13706), .A(n14559), .ZN(n13709) );
  NAND2_X1 U15724 ( .A1(n13709), .A2(n13708), .ZN(n13715) );
  NOR2_X1 U15725 ( .A1(n14568), .A2(n14141), .ZN(n13713) );
  OAI21_X1 U15726 ( .B1(n13711), .B2(n14551), .A(n13710), .ZN(n13712) );
  AOI211_X1 U15727 ( .C1(n13794), .C2(n14576), .A(n13713), .B(n13712), .ZN(
        n13714) );
  OAI211_X1 U15728 ( .C1(n13920), .C2(n13821), .A(n13715), .B(n13714), .ZN(
        P1_U3219) );
  INV_X1 U15729 ( .A(n13716), .ZN(n13717) );
  AOI21_X1 U15730 ( .B1(n13719), .B2(n13718), .A(n13717), .ZN(n13725) );
  NAND2_X1 U15731 ( .A1(n13985), .A2(n14575), .ZN(n13721) );
  NAND2_X1 U15732 ( .A1(n14149), .A2(n14572), .ZN(n13720) );
  NAND2_X1 U15733 ( .A1(n13721), .A2(n13720), .ZN(n14110) );
  AOI22_X1 U15734 ( .A1(n14110), .A2(n13805), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13722) );
  OAI21_X1 U15735 ( .B1(n14111), .B2(n14568), .A(n13722), .ZN(n13723) );
  AOI21_X1 U15736 ( .B1(n14292), .B2(n14564), .A(n13723), .ZN(n13724) );
  OAI21_X1 U15737 ( .B1(n13725), .B2(n14559), .A(n13724), .ZN(P1_U3223) );
  XOR2_X1 U15738 ( .A(n13727), .B(n13726), .Z(n13733) );
  NAND2_X1 U15739 ( .A1(n13988), .A2(n14572), .ZN(n13729) );
  NAND2_X1 U15740 ( .A1(n14020), .A2(n14575), .ZN(n13728) );
  NAND2_X1 U15741 ( .A1(n13729), .A2(n13728), .ZN(n14046) );
  AOI22_X1 U15742 ( .A1(n13805), .A2(n14046), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13730) );
  OAI21_X1 U15743 ( .B1(n14055), .B2(n14568), .A(n13730), .ZN(n13731) );
  AOI21_X1 U15744 ( .B1(n14220), .B2(n14564), .A(n13731), .ZN(n13732) );
  OAI21_X1 U15745 ( .B1(n13733), .B2(n14559), .A(n13732), .ZN(P1_U3225) );
  INV_X1 U15746 ( .A(n13734), .ZN(n13735) );
  NOR2_X1 U15747 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  XNOR2_X1 U15748 ( .A(n13738), .B(n13737), .ZN(n13739) );
  NAND2_X1 U15749 ( .A1(n13739), .A2(n13810), .ZN(n13748) );
  NAND2_X1 U15750 ( .A1(n13794), .A2(n13834), .ZN(n13740) );
  NAND2_X1 U15751 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13890) );
  OAI211_X1 U15752 ( .C1(n13741), .C2(n14551), .A(n13740), .B(n13890), .ZN(
        n13742) );
  INV_X1 U15753 ( .A(n13742), .ZN(n13747) );
  NAND2_X1 U15754 ( .A1(n14564), .A2(n13743), .ZN(n13746) );
  NAND2_X1 U15755 ( .A1(n13817), .A2(n13744), .ZN(n13745) );
  NAND4_X1 U15756 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        P1_U3227) );
  OAI21_X1 U15757 ( .B1(n13752), .B2(n13751), .A(n13750), .ZN(n13753) );
  NAND2_X1 U15758 ( .A1(n13753), .A2(n13810), .ZN(n13758) );
  INV_X1 U15759 ( .A(n14576), .ZN(n13940) );
  NAND2_X1 U15760 ( .A1(n13794), .A2(n14573), .ZN(n13755) );
  OAI211_X1 U15761 ( .C1(n13940), .C2(n14551), .A(n13755), .B(n13754), .ZN(
        n13756) );
  AOI21_X1 U15762 ( .B1(n14578), .B2(n13817), .A(n13756), .ZN(n13757) );
  OAI211_X1 U15763 ( .C1(n14591), .C2(n13821), .A(n13758), .B(n13757), .ZN(
        P1_U3228) );
  XOR2_X1 U15764 ( .A(n13760), .B(n13759), .Z(n13765) );
  NOR2_X1 U15765 ( .A1(n14568), .A2(n14071), .ZN(n13763) );
  INV_X1 U15766 ( .A(n14062), .ZN(n13956) );
  AOI22_X1 U15767 ( .A1(n13794), .A2(n14063), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13761) );
  OAI21_X1 U15768 ( .B1(n13956), .B2(n14551), .A(n13761), .ZN(n13762) );
  AOI211_X1 U15769 ( .C1(n14073), .C2(n14564), .A(n13763), .B(n13762), .ZN(
        n13764) );
  OAI21_X1 U15770 ( .B1(n13765), .B2(n14559), .A(n13764), .ZN(P1_U3229) );
  INV_X1 U15771 ( .A(n14132), .ZN(n14297) );
  OAI211_X1 U15772 ( .C1(n13768), .C2(n13767), .A(n13766), .B(n13810), .ZN(
        n13774) );
  INV_X1 U15773 ( .A(n13769), .ZN(n14125) );
  AND2_X1 U15774 ( .A1(n14163), .A2(n14572), .ZN(n13770) );
  AOI21_X1 U15775 ( .B1(n13983), .B2(n14575), .A(n13770), .ZN(n14123) );
  INV_X1 U15776 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13771) );
  OAI22_X1 U15777 ( .A1(n14123), .A2(n13815), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13771), .ZN(n13772) );
  AOI21_X1 U15778 ( .B1(n14125), .B2(n13817), .A(n13772), .ZN(n13773) );
  OAI211_X1 U15779 ( .C1(n14297), .C2(n13821), .A(n13774), .B(n13773), .ZN(
        P1_U3233) );
  OAI211_X1 U15780 ( .C1(n13776), .C2(n13775), .A(n14542), .B(n13810), .ZN(
        n13782) );
  INV_X1 U15781 ( .A(n14477), .ZN(n13780) );
  OAI21_X1 U15782 ( .B1(n13815), .B2(n13778), .A(n13777), .ZN(n13779) );
  AOI21_X1 U15783 ( .B1(n13780), .B2(n13817), .A(n13779), .ZN(n13781) );
  OAI211_X1 U15784 ( .C1(n13783), .C2(n13821), .A(n13782), .B(n13781), .ZN(
        P1_U3234) );
  OAI21_X1 U15785 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(n13787) );
  NAND2_X1 U15786 ( .A1(n13787), .A2(n13810), .ZN(n13791) );
  AOI22_X1 U15787 ( .A1(n13983), .A2(n14572), .B1(n14575), .B2(n14063), .ZN(
        n14236) );
  INV_X1 U15788 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13788) );
  OAI22_X1 U15789 ( .A1(n14236), .A2(n13815), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13788), .ZN(n13789) );
  AOI21_X1 U15790 ( .B1(n14099), .B2(n13817), .A(n13789), .ZN(n13790) );
  OAI211_X1 U15791 ( .C1(n13821), .C2(n14238), .A(n13791), .B(n13790), .ZN(
        P1_U3235) );
  XOR2_X1 U15792 ( .A(n13793), .B(n13792), .Z(n13800) );
  NOR2_X1 U15793 ( .A1(n14568), .A2(n14168), .ZN(n13798) );
  INV_X1 U15794 ( .A(n14163), .ZN(n13943) );
  NAND2_X1 U15795 ( .A1(n13794), .A2(n13935), .ZN(n13796) );
  OAI211_X1 U15796 ( .C1(n13943), .C2(n14551), .A(n13796), .B(n13795), .ZN(
        n13797) );
  AOI211_X1 U15797 ( .C1(n14303), .C2(n14564), .A(n13798), .B(n13797), .ZN(
        n13799) );
  OAI21_X1 U15798 ( .B1(n13800), .B2(n14559), .A(n13799), .ZN(P1_U3238) );
  XOR2_X1 U15799 ( .A(n13802), .B(n13801), .Z(n13809) );
  NAND2_X1 U15800 ( .A1(n14062), .A2(n14572), .ZN(n13804) );
  NAND2_X1 U15801 ( .A1(n13999), .A2(n14575), .ZN(n13803) );
  NAND2_X1 U15802 ( .A1(n13804), .A2(n13803), .ZN(n14213) );
  AOI22_X1 U15803 ( .A1(n13805), .A2(n14213), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13806) );
  OAI21_X1 U15804 ( .B1(n14031), .B2(n14568), .A(n13806), .ZN(n13807) );
  AOI21_X1 U15805 ( .B1(n14038), .B2(n14564), .A(n13807), .ZN(n13808) );
  OAI21_X1 U15806 ( .B1(n13809), .B2(n14559), .A(n13808), .ZN(P1_U3240) );
  OAI211_X1 U15807 ( .C1(n13812), .C2(n13811), .A(n14555), .B(n13810), .ZN(
        n13820) );
  INV_X1 U15808 ( .A(n13813), .ZN(n13818) );
  NAND2_X1 U15809 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14672)
         );
  OAI21_X1 U15810 ( .B1(n13815), .B2(n13814), .A(n14672), .ZN(n13816) );
  AOI21_X1 U15811 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(n13819) );
  OAI211_X1 U15812 ( .C1(n13822), .C2(n13821), .A(n13820), .B(n13819), .ZN(
        P1_U3241) );
  MUX2_X1 U15813 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13925), .S(n13844), .Z(
        P1_U3591) );
  MUX2_X1 U15814 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13963), .S(n13844), .Z(
        P1_U3590) );
  MUX2_X1 U15815 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13998), .S(n13844), .Z(
        P1_U3589) );
  MUX2_X1 U15816 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14019), .S(n13844), .Z(
        P1_U3588) );
  MUX2_X1 U15817 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13999), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15818 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14020), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15819 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14062), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15820 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13988), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15821 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14063), .S(n13844), .Z(
        P1_U3583) );
  MUX2_X1 U15822 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13985), .S(n13844), .Z(
        P1_U3582) );
  MUX2_X1 U15823 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13983), .S(n13844), .Z(
        P1_U3581) );
  MUX2_X1 U15824 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14149), .S(n13844), .Z(
        P1_U3580) );
  MUX2_X1 U15825 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14163), .S(n13844), .Z(
        P1_U3579) );
  MUX2_X1 U15826 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14576), .S(n13844), .Z(
        P1_U3578) );
  MUX2_X1 U15827 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13935), .S(n13844), .Z(
        P1_U3577) );
  MUX2_X1 U15828 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14573), .S(n13844), .Z(
        P1_U3576) );
  MUX2_X1 U15829 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13823), .S(n13844), .Z(
        P1_U3575) );
  MUX2_X1 U15830 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13824), .S(n13844), .Z(
        P1_U3574) );
  MUX2_X1 U15831 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13825), .S(n13844), .Z(
        P1_U3573) );
  MUX2_X1 U15832 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13826), .S(n13844), .Z(
        P1_U3572) );
  MUX2_X1 U15833 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13827), .S(n13844), .Z(
        P1_U3571) );
  MUX2_X1 U15834 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13828), .S(n13844), .Z(
        P1_U3570) );
  MUX2_X1 U15835 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13829), .S(n13844), .Z(
        P1_U3569) );
  MUX2_X1 U15836 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13830), .S(n13844), .Z(
        P1_U3568) );
  MUX2_X1 U15837 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13831), .S(n13844), .Z(
        P1_U3567) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13832), .S(n13844), .Z(
        P1_U3566) );
  MUX2_X1 U15839 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13833), .S(n13844), .Z(
        P1_U3565) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13834), .S(n13844), .Z(
        P1_U3564) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13835), .S(n13844), .Z(
        P1_U3563) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13836), .S(n13844), .Z(
        P1_U3562) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13837), .S(n13844), .Z(
        P1_U3561) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13838), .S(n13844), .Z(
        P1_U3560) );
  MUX2_X1 U15845 ( .A(n13840), .B(n13839), .S(n6415), .Z(n13845) );
  OAI21_X1 U15846 ( .B1(n6415), .B2(P1_REG2_REG_0__SCAN_IN), .A(n13841), .ZN(
        n14652) );
  NAND2_X1 U15847 ( .A1(n14652), .A2(n13842), .ZN(n13843) );
  OAI211_X1 U15848 ( .C1(n13845), .C2(n6424), .A(n13844), .B(n13843), .ZN(
        n13889) );
  AOI22_X1 U15849 ( .A1(n14655), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13856) );
  OAI21_X1 U15850 ( .B1(n13847), .B2(n13846), .A(n13866), .ZN(n13848) );
  OAI22_X1 U15851 ( .A1(n13850), .A2(n13849), .B1(n14669), .B2(n13848), .ZN(
        n13851) );
  INV_X1 U15852 ( .A(n13851), .ZN(n13855) );
  OAI211_X1 U15853 ( .C1(n13853), .C2(n13852), .A(n13914), .B(n13861), .ZN(
        n13854) );
  NAND4_X1 U15854 ( .A1(n13889), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        P1_U3245) );
  INV_X1 U15855 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14332) );
  OAI22_X1 U15856 ( .A1(n14674), .A2(n14332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13857), .ZN(n13858) );
  AOI21_X1 U15857 ( .B1(n13863), .B2(n14666), .A(n13858), .ZN(n13870) );
  MUX2_X1 U15858 ( .A(n14699), .B(P1_REG2_REG_3__SCAN_IN), .S(n13863), .Z(
        n13859) );
  NAND3_X1 U15859 ( .A1(n13861), .A2(n13860), .A3(n13859), .ZN(n13862) );
  NAND3_X1 U15860 ( .A1(n13914), .A2(n13876), .A3(n13862), .ZN(n13869) );
  MUX2_X1 U15861 ( .A(n9611), .B(P1_REG1_REG_3__SCAN_IN), .S(n13863), .Z(
        n13864) );
  NAND3_X1 U15862 ( .A1(n13866), .A2(n13865), .A3(n13864), .ZN(n13867) );
  NAND3_X1 U15863 ( .A1(n13908), .A2(n13883), .A3(n13867), .ZN(n13868) );
  NAND3_X1 U15864 ( .A1(n13870), .A2(n13869), .A3(n13868), .ZN(P1_U3246) );
  INV_X1 U15865 ( .A(n13871), .ZN(n13872) );
  AOI21_X1 U15866 ( .B1(n14655), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n13872), .ZN(
        n13888) );
  INV_X1 U15867 ( .A(n13873), .ZN(n13901) );
  NAND3_X1 U15868 ( .A1(n13876), .A2(n13875), .A3(n13874), .ZN(n13877) );
  NAND3_X1 U15869 ( .A1(n13914), .A2(n13901), .A3(n13877), .ZN(n13879) );
  NAND2_X1 U15870 ( .A1(n14666), .A2(n13880), .ZN(n13878) );
  AND2_X1 U15871 ( .A1(n13879), .A2(n13878), .ZN(n13887) );
  MUX2_X1 U15872 ( .A(n9933), .B(P1_REG1_REG_4__SCAN_IN), .S(n13880), .Z(
        n13881) );
  NAND3_X1 U15873 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n13884) );
  NAND3_X1 U15874 ( .A1(n13908), .A2(n13885), .A3(n13884), .ZN(n13886) );
  NAND4_X1 U15875 ( .A1(n13889), .A2(n13888), .A3(n13887), .A4(n13886), .ZN(
        P1_U3247) );
  INV_X1 U15876 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15233) );
  OAI21_X1 U15877 ( .B1(n14674), .B2(n15233), .A(n13890), .ZN(n13891) );
  AOI21_X1 U15878 ( .B1(n13892), .B2(n14666), .A(n13891), .ZN(n13906) );
  OAI21_X1 U15879 ( .B1(n13895), .B2(n13894), .A(n13893), .ZN(n13896) );
  NAND2_X1 U15880 ( .A1(n13908), .A2(n13896), .ZN(n13905) );
  INV_X1 U15881 ( .A(n13897), .ZN(n13900) );
  MUX2_X1 U15882 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9946), .S(n13898), .Z(
        n13899) );
  NAND3_X1 U15883 ( .A1(n13901), .A2(n13900), .A3(n13899), .ZN(n13902) );
  NAND3_X1 U15884 ( .A1(n13914), .A2(n13903), .A3(n13902), .ZN(n13904) );
  NAND3_X1 U15885 ( .A1(n13906), .A2(n13905), .A3(n13904), .ZN(P1_U3248) );
  NAND2_X1 U15886 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14565)
         );
  OAI211_X1 U15887 ( .C1(n13910), .C2(n13909), .A(n13908), .B(n13907), .ZN(
        n13911) );
  AND2_X1 U15888 ( .A1(n14565), .A2(n13911), .ZN(n13919) );
  AOI22_X1 U15889 ( .A1(n14666), .A2(n13912), .B1(n14655), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n13918) );
  OAI211_X1 U15890 ( .C1(n13916), .C2(n13915), .A(n13914), .B(n13913), .ZN(
        n13917) );
  NAND3_X1 U15891 ( .A1(n13919), .A2(n13918), .A3(n13917), .ZN(P1_U3259) );
  NOR2_X2 U15892 ( .A1(n14220), .A2(n14045), .ZN(n14044) );
  OR2_X1 U15893 ( .A1(n6415), .A2(n13923), .ZN(n13924) );
  NAND2_X1 U15894 ( .A1(n14575), .A2(n13924), .ZN(n13964) );
  INV_X1 U15895 ( .A(n13964), .ZN(n13926) );
  NAND2_X1 U15896 ( .A1(n13926), .A2(n13925), .ZN(n14196) );
  NOR2_X1 U15897 ( .A1(n14684), .A2(n14196), .ZN(n13931) );
  NOR2_X1 U15898 ( .A1(n14268), .A2(n14101), .ZN(n13927) );
  AOI211_X1 U15899 ( .C1(n14684), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13931), 
        .B(n13927), .ZN(n13928) );
  OAI21_X1 U15900 ( .B1(n14193), .B2(n14173), .A(n13928), .ZN(P1_U3263) );
  OAI211_X1 U15901 ( .C1(n14272), .C2(n13962), .A(n14707), .B(n13929), .ZN(
        n14197) );
  NOR2_X1 U15902 ( .A1(n14272), .A2(n14101), .ZN(n13930) );
  AOI211_X1 U15903 ( .C1(n14684), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13931), 
        .B(n13930), .ZN(n13932) );
  OAI21_X1 U15904 ( .B1(n14173), .B2(n14197), .A(n13932), .ZN(P1_U3264) );
  OR2_X1 U15905 ( .A1(n13973), .A2(n14573), .ZN(n13933) );
  NAND2_X1 U15906 ( .A1(n14569), .A2(n13935), .ZN(n13939) );
  NAND2_X1 U15907 ( .A1(n13936), .A2(n14552), .ZN(n13937) );
  NAND2_X1 U15908 ( .A1(n13937), .A2(n14591), .ZN(n13938) );
  OR2_X1 U15909 ( .A1(n14303), .A2(n13940), .ZN(n13941) );
  INV_X1 U15910 ( .A(n14112), .ZN(n13984) );
  NAND2_X1 U15911 ( .A1(n14108), .A2(n13984), .ZN(n13948) );
  OR2_X1 U15912 ( .A1(n14292), .A2(n13946), .ZN(n13947) );
  INV_X1 U15913 ( .A(n13985), .ZN(n13949) );
  NAND2_X1 U15914 ( .A1(n13986), .A2(n13949), .ZN(n13950) );
  NAND2_X1 U15915 ( .A1(n14082), .A2(n14081), .ZN(n14080) );
  INV_X1 U15916 ( .A(n14063), .ZN(n13951) );
  NAND2_X1 U15917 ( .A1(n14232), .A2(n13951), .ZN(n13952) );
  INV_X1 U15918 ( .A(n13988), .ZN(n13953) );
  OR2_X1 U15919 ( .A1(n14073), .A2(n13953), .ZN(n13954) );
  NAND2_X1 U15920 ( .A1(n14220), .A2(n13956), .ZN(n13957) );
  NAND2_X1 U15921 ( .A1(n14280), .A2(n14020), .ZN(n13959) );
  INV_X1 U15922 ( .A(n14026), .ZN(n14276) );
  AOI211_X1 U15923 ( .C1(n14202), .C2(n14003), .A(n14718), .B(n13962), .ZN(
        n14200) );
  INV_X1 U15924 ( .A(n13963), .ZN(n13965) );
  NOR2_X1 U15925 ( .A1(n13965), .A2(n13964), .ZN(n14201) );
  NAND3_X1 U15926 ( .A1(n13967), .A2(n14201), .A3(n13966), .ZN(n13968) );
  OAI21_X1 U15927 ( .B1(n14698), .B2(n13969), .A(n13968), .ZN(n13970) );
  AOI21_X1 U15928 ( .B1(n14684), .B2(P1_REG2_REG_29__SCAN_IN), .A(n13970), 
        .ZN(n13971) );
  OAI21_X1 U15929 ( .B1(n6419), .B2(n14101), .A(n13971), .ZN(n13995) );
  NAND2_X1 U15930 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  OR2_X1 U15931 ( .A1(n14303), .A2(n14576), .ZN(n13978) );
  NAND2_X1 U15932 ( .A1(n14158), .A2(n13978), .ZN(n13980) );
  NAND2_X1 U15933 ( .A1(n14303), .A2(n14576), .ZN(n13979) );
  OR2_X1 U15934 ( .A1(n14153), .A2(n14163), .ZN(n13981) );
  NAND2_X1 U15935 ( .A1(n14132), .A2(n14149), .ZN(n13982) );
  NAND2_X1 U15936 ( .A1(n14232), .A2(n14063), .ZN(n13987) );
  NAND2_X1 U15937 ( .A1(n14078), .A2(n13987), .ZN(n14061) );
  NAND2_X1 U15938 ( .A1(n14220), .A2(n14062), .ZN(n13989) );
  AND2_X1 U15939 ( .A1(n14038), .A2(n14020), .ZN(n13990) );
  NOR2_X1 U15940 ( .A1(n14026), .A2(n13999), .ZN(n13991) );
  INV_X1 U15941 ( .A(n13992), .ZN(n13993) );
  NOR2_X1 U15942 ( .A1(n14203), .A2(n14114), .ZN(n13994) );
  OAI21_X1 U15943 ( .B1(n14204), .B2(n14684), .A(n13996), .ZN(P1_U3356) );
  NAND2_X1 U15944 ( .A1(n13999), .A2(n14572), .ZN(n14000) );
  INV_X1 U15945 ( .A(n14003), .ZN(n14004) );
  AOI21_X1 U15946 ( .B1(n14205), .B2(n6468), .A(n14004), .ZN(n14206) );
  INV_X1 U15947 ( .A(n14005), .ZN(n14006) );
  AOI22_X1 U15948 ( .A1(n14684), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14006), 
        .B2(n14683), .ZN(n14007) );
  OAI21_X1 U15949 ( .B1(n13921), .B2(n14101), .A(n14007), .ZN(n14012) );
  OAI21_X1 U15950 ( .B1(n14010), .B2(n14009), .A(n14008), .ZN(n14209) );
  NOR2_X1 U15951 ( .A1(n14209), .A2(n14114), .ZN(n14011) );
  AOI211_X1 U15952 ( .C1(n14206), .C2(n14013), .A(n14012), .B(n14011), .ZN(
        n14014) );
  OAI21_X1 U15953 ( .B1(n14208), .B2(n14684), .A(n14014), .ZN(P1_U3265) );
  AOI21_X1 U15954 ( .B1(n14026), .B2(n14035), .A(n14718), .ZN(n14015) );
  AND2_X1 U15955 ( .A1(n14015), .A2(n6468), .ZN(n14210) );
  INV_X1 U15956 ( .A(n14210), .ZN(n14029) );
  INV_X1 U15957 ( .A(n14017), .ZN(n14016) );
  AOI22_X1 U15958 ( .A1(n14572), .A2(n14020), .B1(n14019), .B2(n14575), .ZN(
        n14021) );
  NAND2_X1 U15959 ( .A1(n14022), .A2(n14021), .ZN(n14211) );
  NAND2_X1 U15960 ( .A1(n14211), .A2(n14700), .ZN(n14028) );
  OAI22_X1 U15961 ( .A1(n14700), .A2(n14024), .B1(n14023), .B2(n14698), .ZN(
        n14025) );
  AOI21_X1 U15962 ( .B1(n14026), .B2(n14702), .A(n14025), .ZN(n14027) );
  OAI211_X1 U15963 ( .C1(n14173), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        P1_U3266) );
  XNOR2_X1 U15964 ( .A(n14030), .B(n14039), .ZN(n14217) );
  INV_X1 U15965 ( .A(n14031), .ZN(n14032) );
  AOI22_X1 U15966 ( .A1(n14700), .A2(n14213), .B1(n14032), .B2(n14683), .ZN(
        n14033) );
  OAI21_X1 U15967 ( .B1(n14034), .B2(n14700), .A(n14033), .ZN(n14037) );
  OAI211_X1 U15968 ( .C1(n14280), .C2(n14044), .A(n14707), .B(n14035), .ZN(
        n14215) );
  NOR2_X1 U15969 ( .A1(n14215), .A2(n14173), .ZN(n14036) );
  AOI211_X1 U15970 ( .C1(n14702), .C2(n14038), .A(n14037), .B(n14036), .ZN(
        n14043) );
  INV_X1 U15971 ( .A(n14039), .ZN(n14040) );
  XNOR2_X1 U15972 ( .A(n14041), .B(n14040), .ZN(n14212) );
  NAND2_X1 U15973 ( .A1(n14212), .A2(n14181), .ZN(n14042) );
  OAI211_X1 U15974 ( .C1(n14217), .C2(n14114), .A(n14043), .B(n14042), .ZN(
        P1_U3267) );
  AOI211_X1 U15975 ( .C1(n14220), .C2(n14045), .A(n14718), .B(n14044), .ZN(
        n14047) );
  OR2_X1 U15976 ( .A1(n14047), .A2(n14046), .ZN(n14221) );
  INV_X1 U15977 ( .A(n14048), .ZN(n14049) );
  AOI21_X1 U15978 ( .B1(n14052), .B2(n14050), .A(n14049), .ZN(n14054) );
  OAI211_X1 U15979 ( .C1(n14052), .C2(n6531), .A(n14051), .B(n14762), .ZN(
        n14053) );
  OAI21_X1 U15980 ( .B1(n14054), .B2(n14570), .A(n14053), .ZN(n14222) );
  AOI21_X1 U15981 ( .B1(n14471), .B2(n14221), .A(n14222), .ZN(n14059) );
  OAI22_X1 U15982 ( .A1(n14700), .A2(n14056), .B1(n14055), .B2(n14698), .ZN(
        n14057) );
  AOI21_X1 U15983 ( .B1(n14220), .B2(n14702), .A(n14057), .ZN(n14058) );
  OAI21_X1 U15984 ( .B1(n14059), .B2(n14684), .A(n14058), .ZN(P1_U3268) );
  AOI21_X1 U15985 ( .B1(n14065), .B2(n14061), .A(n14060), .ZN(n14069) );
  AOI22_X1 U15986 ( .A1(n14572), .A2(n14063), .B1(n14062), .B2(n14575), .ZN(
        n14068) );
  OAI211_X1 U15987 ( .C1(n14066), .C2(n14065), .A(n14064), .B(n14751), .ZN(
        n14067) );
  OAI211_X1 U15988 ( .C1(n14069), .C2(n14609), .A(n14068), .B(n14067), .ZN(
        n14226) );
  INV_X1 U15989 ( .A(n14226), .ZN(n14077) );
  XNOR2_X1 U15990 ( .A(n14073), .B(n14083), .ZN(n14070) );
  NOR2_X1 U15991 ( .A1(n14070), .A2(n14718), .ZN(n14225) );
  OAI22_X1 U15992 ( .A1(n14700), .A2(n14072), .B1(n14071), .B2(n14698), .ZN(
        n14075) );
  NOR2_X1 U15993 ( .A1(n6991), .A2(n14101), .ZN(n14074) );
  AOI211_X1 U15994 ( .C1(n14225), .C2(n14711), .A(n14075), .B(n14074), .ZN(
        n14076) );
  OAI21_X1 U15995 ( .B1(n14077), .B2(n14684), .A(n14076), .ZN(P1_U3269) );
  INV_X1 U15996 ( .A(n14081), .ZN(n14079) );
  OAI21_X1 U15997 ( .B1(n6494), .B2(n14079), .A(n14078), .ZN(n14235) );
  OAI21_X1 U15998 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14229) );
  INV_X1 U15999 ( .A(n14232), .ZN(n14090) );
  AOI21_X1 U16000 ( .B1(n14232), .B2(n14098), .A(n14718), .ZN(n14084) );
  AND2_X1 U16001 ( .A1(n14084), .A2(n14083), .ZN(n14230) );
  NAND2_X1 U16002 ( .A1(n14230), .A2(n14711), .ZN(n14089) );
  OAI22_X1 U16003 ( .A1(n14700), .A2(n14086), .B1(n14085), .B2(n14698), .ZN(
        n14087) );
  AOI21_X1 U16004 ( .B1(n14231), .B2(n14700), .A(n14087), .ZN(n14088) );
  OAI211_X1 U16005 ( .C1(n14090), .C2(n14101), .A(n14089), .B(n14088), .ZN(
        n14091) );
  AOI21_X1 U16006 ( .B1(n14229), .B2(n14181), .A(n14091), .ZN(n14092) );
  OAI21_X1 U16007 ( .B1(n14114), .B2(n14235), .A(n14092), .ZN(P1_U3270) );
  XOR2_X1 U16008 ( .A(n14093), .B(n14095), .Z(n14242) );
  OAI21_X1 U16009 ( .B1(n14096), .B2(n14095), .A(n14094), .ZN(n14240) );
  OAI211_X1 U16010 ( .C1(n14238), .C2(n14097), .A(n14707), .B(n14098), .ZN(
        n14237) );
  INV_X1 U16011 ( .A(n14099), .ZN(n14100) );
  OAI22_X1 U16012 ( .A1(n14236), .A2(n14684), .B1(n14100), .B2(n14698), .ZN(
        n14103) );
  NOR2_X1 U16013 ( .A1(n14238), .A2(n14101), .ZN(n14102) );
  AOI211_X1 U16014 ( .C1(n14684), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14103), 
        .B(n14102), .ZN(n14104) );
  OAI21_X1 U16015 ( .B1(n14173), .B2(n14237), .A(n14104), .ZN(n14105) );
  AOI21_X1 U16016 ( .B1(n14712), .B2(n14240), .A(n14105), .ZN(n14106) );
  OAI21_X1 U16017 ( .B1(n14242), .B2(n14107), .A(n14106), .ZN(P1_U3271) );
  XNOR2_X1 U16018 ( .A(n14108), .B(n14112), .ZN(n14109) );
  NAND2_X1 U16019 ( .A1(n14109), .A2(n14751), .ZN(n14246) );
  INV_X1 U16020 ( .A(n14110), .ZN(n14243) );
  OAI211_X1 U16021 ( .C1(n14698), .C2(n14111), .A(n14246), .B(n14243), .ZN(
        n14120) );
  XNOR2_X1 U16022 ( .A(n14113), .B(n14112), .ZN(n14247) );
  NOR2_X1 U16023 ( .A1(n14247), .A2(n14114), .ZN(n14119) );
  AOI21_X1 U16024 ( .B1(n14292), .B2(n14130), .A(n14718), .ZN(n14116) );
  NAND2_X1 U16025 ( .A1(n14116), .A2(n14115), .ZN(n14244) );
  AOI22_X1 U16026 ( .A1(n14292), .A2(n14702), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14684), .ZN(n14117) );
  OAI21_X1 U16027 ( .B1(n14244), .B2(n14173), .A(n14117), .ZN(n14118) );
  AOI211_X1 U16028 ( .C1(n14120), .C2(n14700), .A(n14119), .B(n14118), .ZN(
        n14121) );
  INV_X1 U16029 ( .A(n14121), .ZN(P1_U3272) );
  OAI211_X1 U16030 ( .C1(n6567), .C2(n14126), .A(n14122), .B(n14751), .ZN(
        n14124) );
  NAND2_X1 U16031 ( .A1(n14124), .A2(n14123), .ZN(n14250) );
  AOI21_X1 U16032 ( .B1(n14125), .B2(n14683), .A(n14250), .ZN(n14137) );
  NAND2_X1 U16033 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  AND2_X1 U16034 ( .A1(n14129), .A2(n14128), .ZN(n14252) );
  INV_X1 U16035 ( .A(n14130), .ZN(n14131) );
  AOI211_X1 U16036 ( .C1(n14132), .C2(n14140), .A(n14718), .B(n14131), .ZN(
        n14251) );
  INV_X1 U16037 ( .A(n14251), .ZN(n14134) );
  AOI22_X1 U16038 ( .A1(n14132), .A2(n14702), .B1(n14684), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14133) );
  OAI21_X1 U16039 ( .B1(n14134), .B2(n14173), .A(n14133), .ZN(n14135) );
  AOI21_X1 U16040 ( .B1(n14712), .B2(n14252), .A(n14135), .ZN(n14136) );
  OAI21_X1 U16041 ( .B1(n14137), .B2(n14684), .A(n14136), .ZN(P1_U3273) );
  INV_X1 U16042 ( .A(n14138), .ZN(n14171) );
  NAND2_X1 U16043 ( .A1(n14153), .A2(n14171), .ZN(n14139) );
  AND3_X1 U16044 ( .A1(n14140), .A2(n14707), .A3(n14139), .ZN(n14255) );
  NOR2_X1 U16045 ( .A1(n14141), .A2(n14698), .ZN(n14152) );
  INV_X1 U16046 ( .A(n14144), .ZN(n14143) );
  AOI22_X1 U16047 ( .A1(n14142), .A2(n14751), .B1(n14143), .B2(n14762), .ZN(
        n14148) );
  INV_X1 U16048 ( .A(n14142), .ZN(n14145) );
  AOI22_X1 U16049 ( .A1(n14145), .A2(n14751), .B1(n14762), .B2(n14144), .ZN(
        n14147) );
  MUX2_X1 U16050 ( .A(n14148), .B(n14147), .S(n14146), .Z(n14151) );
  AOI22_X1 U16051 ( .A1(n14149), .A2(n14575), .B1(n14572), .B2(n14576), .ZN(
        n14150) );
  NAND2_X1 U16052 ( .A1(n14151), .A2(n14150), .ZN(n14256) );
  AOI211_X1 U16053 ( .C1(n14255), .C2(n14471), .A(n14152), .B(n14256), .ZN(
        n14155) );
  AOI22_X1 U16054 ( .A1(n14153), .A2(n14702), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n14684), .ZN(n14154) );
  OAI21_X1 U16055 ( .B1(n14155), .B2(n14684), .A(n14154), .ZN(P1_U3274) );
  NAND2_X1 U16056 ( .A1(n14156), .A2(n14751), .ZN(n14157) );
  OAI21_X1 U16057 ( .B1(n14609), .B2(n14158), .A(n14157), .ZN(n14162) );
  INV_X1 U16058 ( .A(n14158), .ZN(n14159) );
  OAI22_X1 U16059 ( .A1(n14156), .A2(n14570), .B1(n14159), .B2(n14609), .ZN(
        n14161) );
  MUX2_X1 U16060 ( .A(n14162), .B(n14161), .S(n14160), .Z(n14167) );
  NAND2_X1 U16061 ( .A1(n14163), .A2(n14575), .ZN(n14164) );
  OAI21_X1 U16062 ( .B1(n14552), .B2(n14165), .A(n14164), .ZN(n14166) );
  NOR2_X1 U16063 ( .A1(n14167), .A2(n14166), .ZN(n14261) );
  OAI22_X1 U16064 ( .A1(n14700), .A2(n14169), .B1(n14168), .B2(n14698), .ZN(
        n14170) );
  AOI21_X1 U16065 ( .B1(n14303), .B2(n14702), .A(n14170), .ZN(n14175) );
  AOI21_X1 U16066 ( .B1(n14584), .B2(n14303), .A(n14718), .ZN(n14172) );
  NAND2_X1 U16067 ( .A1(n14172), .A2(n14171), .ZN(n14260) );
  OR2_X1 U16068 ( .A1(n14260), .A2(n14173), .ZN(n14174) );
  OAI211_X1 U16069 ( .C1(n14261), .C2(n14684), .A(n14175), .B(n14174), .ZN(
        P1_U3275) );
  XNOR2_X1 U16070 ( .A(n14176), .B(n7146), .ZN(n14761) );
  NAND2_X1 U16071 ( .A1(n14761), .A2(n14712), .ZN(n14192) );
  OAI22_X1 U16072 ( .A1(n14700), .A2(n14178), .B1(n14177), .B2(n14698), .ZN(
        n14179) );
  AOI21_X1 U16073 ( .B1(n14702), .B2(n14756), .A(n14179), .ZN(n14191) );
  NAND2_X1 U16074 ( .A1(n14180), .A2(n7146), .ZN(n14752) );
  NAND3_X1 U16075 ( .A1(n14753), .A2(n14752), .A3(n14181), .ZN(n14190) );
  NAND2_X1 U16076 ( .A1(n14756), .A2(n14689), .ZN(n14182) );
  NAND3_X1 U16077 ( .A1(n14183), .A2(n14707), .A3(n14182), .ZN(n14757) );
  AOI21_X1 U16078 ( .B1(n14757), .B2(n14185), .A(n14184), .ZN(n14188) );
  INV_X1 U16079 ( .A(n14186), .ZN(n14187) );
  OAI21_X1 U16080 ( .B1(n14188), .B2(n14187), .A(n14700), .ZN(n14189) );
  NAND4_X1 U16081 ( .A1(n14192), .A2(n14191), .A3(n14190), .A4(n14189), .ZN(
        P1_U3283) );
  MUX2_X1 U16082 ( .A(n14194), .B(n14265), .S(n14772), .Z(n14195) );
  AND2_X1 U16083 ( .A1(n14197), .A2(n14196), .ZN(n14269) );
  MUX2_X1 U16084 ( .A(n14198), .B(n14269), .S(n14772), .Z(n14199) );
  OAI21_X1 U16085 ( .B1(n14272), .B2(n14259), .A(n14199), .ZN(P1_U3558) );
  AOI22_X1 U16086 ( .A1(n14206), .A2(n14707), .B1(n14205), .B2(n14755), .ZN(
        n14207) );
  MUX2_X1 U16087 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14273), .S(n14772), .Z(
        P1_U3556) );
  INV_X1 U16088 ( .A(n14213), .ZN(n14214) );
  AND2_X1 U16089 ( .A1(n14215), .A2(n14214), .ZN(n14216) );
  MUX2_X1 U16090 ( .A(n14277), .B(P1_REG1_REG_26__SCAN_IN), .S(n6820), .Z(
        n14218) );
  INV_X1 U16091 ( .A(n14218), .ZN(n14219) );
  INV_X1 U16092 ( .A(n14220), .ZN(n14284) );
  INV_X1 U16093 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n14223) );
  NOR2_X1 U16094 ( .A1(n14222), .A2(n14221), .ZN(n14281) );
  MUX2_X1 U16095 ( .A(n14223), .B(n14281), .S(n14772), .Z(n14224) );
  OAI21_X1 U16096 ( .B1(n14284), .B2(n14259), .A(n14224), .ZN(P1_U3553) );
  INV_X1 U16097 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14227) );
  NOR2_X1 U16098 ( .A1(n14226), .A2(n14225), .ZN(n14285) );
  MUX2_X1 U16099 ( .A(n14227), .B(n14285), .S(n14772), .Z(n14228) );
  OAI21_X1 U16100 ( .B1(n6991), .B2(n14259), .A(n14228), .ZN(P1_U3552) );
  NAND2_X1 U16101 ( .A1(n14229), .A2(n14751), .ZN(n14234) );
  AOI211_X1 U16102 ( .C1(n14232), .C2(n14755), .A(n14231), .B(n14230), .ZN(
        n14233) );
  OAI211_X1 U16103 ( .C1(n14235), .C2(n14609), .A(n14234), .B(n14233), .ZN(
        n14288) );
  MUX2_X1 U16104 ( .A(n14288), .B(P1_REG1_REG_23__SCAN_IN), .S(n6820), .Z(
        P1_U3551) );
  INV_X1 U16105 ( .A(n14755), .ZN(n14746) );
  OAI211_X1 U16106 ( .C1(n14746), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14239) );
  AOI21_X1 U16107 ( .B1(n14240), .B2(n14762), .A(n14239), .ZN(n14241) );
  OAI21_X1 U16108 ( .B1(n14242), .B2(n14570), .A(n14241), .ZN(n14289) );
  MUX2_X1 U16109 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14289), .S(n14772), .Z(
        P1_U3550) );
  AND2_X1 U16110 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  OAI211_X1 U16111 ( .C1(n14247), .C2(n14609), .A(n14246), .B(n14245), .ZN(
        n14290) );
  MUX2_X1 U16112 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14290), .S(n14772), .Z(
        n14248) );
  AOI21_X1 U16113 ( .B1(n14263), .B2(n14292), .A(n14248), .ZN(n14249) );
  INV_X1 U16114 ( .A(n14249), .ZN(P1_U3549) );
  AOI211_X1 U16115 ( .C1(n14762), .C2(n14252), .A(n14251), .B(n14250), .ZN(
        n14294) );
  MUX2_X1 U16116 ( .A(n14253), .B(n14294), .S(n14772), .Z(n14254) );
  OAI21_X1 U16117 ( .B1(n14297), .B2(n14259), .A(n14254), .ZN(P1_U3548) );
  INV_X1 U16118 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14257) );
  NOR2_X1 U16119 ( .A1(n14256), .A2(n14255), .ZN(n14298) );
  MUX2_X1 U16120 ( .A(n14257), .B(n14298), .S(n14772), .Z(n14258) );
  OAI21_X1 U16121 ( .B1(n13920), .B2(n14259), .A(n14258), .ZN(P1_U3547) );
  NAND2_X1 U16122 ( .A1(n14261), .A2(n14260), .ZN(n14301) );
  MUX2_X1 U16123 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14301), .S(n14772), .Z(
        n14262) );
  AOI21_X1 U16124 ( .B1(n14263), .B2(n14303), .A(n14262), .ZN(n14264) );
  INV_X1 U16125 ( .A(n14264), .ZN(P1_U3546) );
  INV_X1 U16126 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14266) );
  MUX2_X1 U16127 ( .A(n14266), .B(n14265), .S(n14764), .Z(n14267) );
  INV_X1 U16128 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14270) );
  MUX2_X1 U16129 ( .A(n14270), .B(n14269), .S(n14764), .Z(n14271) );
  OAI21_X1 U16130 ( .B1(n14272), .B2(n14300), .A(n14271), .ZN(P1_U3526) );
  MUX2_X1 U16131 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14273), .S(n14764), .Z(
        P1_U3524) );
  MUX2_X1 U16132 ( .A(n14277), .B(P1_REG0_REG_26__SCAN_IN), .S(n14763), .Z(
        n14278) );
  INV_X1 U16133 ( .A(n14278), .ZN(n14279) );
  MUX2_X1 U16134 ( .A(n14282), .B(n14281), .S(n14764), .Z(n14283) );
  OAI21_X1 U16135 ( .B1(n14284), .B2(n14300), .A(n14283), .ZN(P1_U3521) );
  MUX2_X1 U16136 ( .A(n14286), .B(n14285), .S(n14764), .Z(n14287) );
  OAI21_X1 U16137 ( .B1(n6991), .B2(n14300), .A(n14287), .ZN(P1_U3520) );
  MUX2_X1 U16138 ( .A(n14288), .B(P1_REG0_REG_23__SCAN_IN), .S(n14763), .Z(
        P1_U3519) );
  MUX2_X1 U16139 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14289), .S(n14764), .Z(
        P1_U3518) );
  MUX2_X1 U16140 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14290), .S(n14764), .Z(
        n14291) );
  AOI21_X1 U16141 ( .B1(n6824), .B2(n14292), .A(n14291), .ZN(n14293) );
  INV_X1 U16142 ( .A(n14293), .ZN(P1_U3517) );
  INV_X1 U16143 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14295) );
  MUX2_X1 U16144 ( .A(n14295), .B(n14294), .S(n14764), .Z(n14296) );
  OAI21_X1 U16145 ( .B1(n14297), .B2(n14300), .A(n14296), .ZN(P1_U3516) );
  MUX2_X1 U16146 ( .A(n15312), .B(n14298), .S(n14764), .Z(n14299) );
  OAI21_X1 U16147 ( .B1(n13920), .B2(n14300), .A(n14299), .ZN(P1_U3515) );
  MUX2_X1 U16148 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14301), .S(n14764), .Z(
        n14302) );
  AOI21_X1 U16149 ( .B1(n6824), .B2(n14303), .A(n14302), .ZN(n14304) );
  INV_X1 U16150 ( .A(n14304), .ZN(P1_U3513) );
  INV_X1 U16151 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14306) );
  NAND3_X1 U16152 ( .A1(n14306), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14308) );
  OAI22_X1 U16153 ( .A1(n14305), .A2(n14308), .B1(n14307), .B2(n6421), .ZN(
        n14309) );
  AOI21_X1 U16154 ( .B1(n13669), .B2(n14310), .A(n14309), .ZN(n14311) );
  INV_X1 U16155 ( .A(n14311), .ZN(P1_U3324) );
  OAI222_X1 U16156 ( .A1(P1_U3086), .A2(n14314), .B1(n11530), .B2(n14313), 
        .C1(n14312), .C2(n6421), .ZN(P1_U3326) );
  OAI222_X1 U16157 ( .A1(P1_U3086), .A2(n6424), .B1(n11530), .B2(n14316), .C1(
        n14315), .C2(n6421), .ZN(P1_U3327) );
  OAI222_X1 U16158 ( .A1(P1_U3086), .A2(n6415), .B1(n11530), .B2(n14319), .C1(
        n14318), .C2(n6421), .ZN(P1_U3328) );
  INV_X1 U16159 ( .A(n14320), .ZN(n14324) );
  OAI222_X1 U16160 ( .A1(n14324), .A2(P1_U3086), .B1(n11530), .B2(n14322), 
        .C1(n14321), .C2(n6421), .ZN(P1_U3329) );
  MUX2_X1 U16161 ( .A(n6831), .B(n14325), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16162 ( .A(n14327), .ZN(n14328) );
  MUX2_X1 U16163 ( .A(n14328), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16164 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14364) );
  OR2_X1 U16165 ( .A1(n14364), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14362) );
  INV_X1 U16166 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14675) );
  INV_X1 U16167 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14329) );
  NOR2_X1 U16168 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14329), .ZN(n14361) );
  XOR2_X1 U16169 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14418) );
  INV_X1 U16170 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14359) );
  INV_X1 U16171 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14357) );
  XOR2_X1 U16172 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14369) );
  XNOR2_X1 U16173 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14350), .ZN(n14374) );
  XNOR2_X1 U16174 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14402) );
  XNOR2_X1 U16175 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14377) );
  NAND2_X1 U16176 ( .A1(n14380), .A2(n14379), .ZN(n14330) );
  NAND2_X1 U16177 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14331), .ZN(n14334) );
  NAND2_X1 U16178 ( .A1(n14376), .A2(n14332), .ZN(n14333) );
  NAND2_X1 U16179 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14335), .ZN(n14337) );
  INV_X1 U16180 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14336) );
  NAND2_X1 U16181 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14338), .ZN(n14340) );
  NAND2_X1 U16182 ( .A1(n14389), .A2(n15233), .ZN(n14339) );
  OR2_X1 U16183 ( .A1(n14342), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14341) );
  INV_X1 U16184 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U16185 ( .A1(n14344), .A2(n14343), .ZN(n14346) );
  XNOR2_X1 U16186 ( .A(n14344), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U16187 ( .A1(n14397), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14345) );
  NOR2_X1 U16188 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14351), .ZN(n14409) );
  NAND2_X1 U16189 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14351), .ZN(n14411) );
  INV_X1 U16190 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14353) );
  XNOR2_X1 U16191 ( .A(n14353), .B(n14355), .ZN(n14371) );
  NAND2_X1 U16192 ( .A1(n14372), .A2(n14371), .ZN(n14354) );
  AND2_X1 U16193 ( .A1(n14359), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14358) );
  OAI22_X1 U16194 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14359), .B1(n14415), 
        .B2(n14358), .ZN(n14417) );
  NOR2_X1 U16195 ( .A1(n14418), .A2(n14417), .ZN(n14360) );
  AOI21_X1 U16196 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15295), .A(n14360), 
        .ZN(n14368) );
  OAI22_X1 U16197 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14675), .B1(n14361), 
        .B2(n14368), .ZN(n14366) );
  AOI22_X1 U16198 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14364), .B1(n14362), 
        .B2(n14366), .ZN(n14426) );
  XOR2_X1 U16199 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14426), .Z(n14428) );
  XNOR2_X1 U16200 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14428), .ZN(n14423) );
  NAND2_X1 U16201 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14364), .ZN(n14363) );
  OAI21_X1 U16202 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14364), .A(n14363), 
        .ZN(n14365) );
  XOR2_X1 U16203 ( .A(n14366), .B(n14365), .Z(n14649) );
  XOR2_X1 U16204 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14367) );
  XOR2_X1 U16205 ( .A(n14368), .B(n14367), .Z(n14421) );
  XOR2_X1 U16206 ( .A(n14370), .B(n14369), .Z(n14632) );
  XNOR2_X1 U16207 ( .A(n14372), .B(n14371), .ZN(n14628) );
  XOR2_X1 U16208 ( .A(n14374), .B(n14373), .Z(n14407) );
  INV_X1 U16209 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14813) );
  NOR2_X1 U16210 ( .A1(n14387), .A2(n14813), .ZN(n14388) );
  XNOR2_X1 U16211 ( .A(n14376), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15367) );
  XOR2_X1 U16212 ( .A(n14378), .B(n14377), .Z(n14438) );
  INV_X1 U16213 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14383) );
  NOR2_X1 U16214 ( .A1(n14382), .A2(n14383), .ZN(n14384) );
  AOI21_X1 U16215 ( .B1(n15090), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14380), .ZN(
        n15361) );
  INV_X1 U16216 ( .A(n15361), .ZN(n14381) );
  NAND2_X1 U16217 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n14381), .ZN(n15371) );
  NOR2_X1 U16218 ( .A1(n14438), .A2(n14437), .ZN(n14385) );
  NAND2_X1 U16219 ( .A1(n14438), .A2(n14437), .ZN(n14436) );
  NAND2_X1 U16220 ( .A1(n15367), .A2(n15366), .ZN(n14386) );
  NOR2_X1 U16221 ( .A1(n15367), .A2(n15366), .ZN(n15365) );
  XNOR2_X1 U16222 ( .A(n14813), .B(n14387), .ZN(n15356) );
  NOR2_X1 U16223 ( .A1(n15357), .A2(n15356), .ZN(n15355) );
  NAND2_X1 U16224 ( .A1(n14390), .A2(n14391), .ZN(n14392) );
  INV_X1 U16225 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15359) );
  INV_X1 U16226 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15278) );
  NOR2_X1 U16227 ( .A1(n14393), .A2(n15278), .ZN(n14396) );
  XNOR2_X1 U16228 ( .A(n14393), .B(n15278), .ZN(n14458) );
  XOR2_X1 U16229 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n14394) );
  XNOR2_X1 U16230 ( .A(n14395), .B(n14394), .ZN(n14457) );
  INV_X1 U16231 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14399) );
  NOR2_X1 U16232 ( .A1(n14398), .A2(n14399), .ZN(n14400) );
  XNOR2_X1 U16233 ( .A(n14397), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15364) );
  XNOR2_X1 U16234 ( .A(n14402), .B(n14401), .ZN(n14404) );
  NAND2_X1 U16235 ( .A1(n14403), .A2(n14404), .ZN(n14405) );
  INV_X1 U16236 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14460) );
  NOR2_X1 U16237 ( .A1(n14407), .A2(n14406), .ZN(n14408) );
  INV_X1 U16238 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14847) );
  INV_X1 U16239 ( .A(n14409), .ZN(n14410) );
  NAND2_X1 U16240 ( .A1(n14411), .A2(n14410), .ZN(n14412) );
  XNOR2_X1 U16241 ( .A(n14412), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U16242 ( .A1(n14632), .A2(n14631), .ZN(n14413) );
  XOR2_X1 U16243 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14414) );
  XOR2_X1 U16244 ( .A(n14415), .B(n14414), .Z(n14635) );
  NAND2_X1 U16245 ( .A1(n14636), .A2(n14635), .ZN(n14416) );
  XOR2_X1 U16246 ( .A(n14418), .B(n14417), .Z(n14420) );
  INV_X1 U16247 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14642) );
  INV_X1 U16248 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14647) );
  NAND2_X1 U16249 ( .A1(n14423), .A2(n14424), .ZN(n14425) );
  INV_X1 U16250 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15294) );
  INV_X1 U16251 ( .A(n14426), .ZN(n14427) );
  NOR2_X1 U16252 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14427), .ZN(n14431) );
  INV_X1 U16253 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14429) );
  NOR2_X1 U16254 ( .A1(n14429), .A2(n14428), .ZN(n14430) );
  OR2_X1 U16255 ( .A1(n14431), .A2(n14430), .ZN(n14480) );
  NAND2_X1 U16256 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14483), .ZN(n14432) );
  OAI21_X1 U16257 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14483), .A(n14432), 
        .ZN(n14481) );
  XNOR2_X1 U16258 ( .A(n14480), .B(n14481), .ZN(n14484) );
  XNOR2_X1 U16259 ( .A(n14433), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16260 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14434) );
  OAI21_X1 U16261 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14434), 
        .ZN(U28) );
  AOI21_X1 U16262 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14435) );
  OAI21_X1 U16263 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14435), 
        .ZN(U29) );
  OAI21_X1 U16264 ( .B1(n14438), .B2(n14437), .A(n14436), .ZN(n14439) );
  XNOR2_X1 U16265 ( .A(n14439), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  INV_X1 U16266 ( .A(n14440), .ZN(n14441) );
  AOI22_X1 U16267 ( .A1(n14441), .A2(n14446), .B1(SI_9_), .B2(n14445), .ZN(
        n14442) );
  OAI21_X1 U16268 ( .B1(P3_U3151), .B2(n14443), .A(n14442), .ZN(P3_U3286) );
  INV_X1 U16269 ( .A(n14444), .ZN(n14447) );
  AOI22_X1 U16270 ( .A1(n14447), .A2(n14446), .B1(SI_11_), .B2(n14445), .ZN(
        n14448) );
  OAI21_X1 U16271 ( .B1(P3_U3151), .B2(n14449), .A(n14448), .ZN(P3_U3284) );
  OAI22_X1 U16272 ( .A1(n14452), .A2(n14451), .B1(n14450), .B2(n12997), .ZN(
        n14453) );
  INV_X1 U16273 ( .A(n14453), .ZN(n14454) );
  OAI21_X1 U16274 ( .B1(P3_U3151), .B2(n14455), .A(n14454), .ZN(P3_U3282) );
  AOI21_X1 U16275 ( .B1(n14458), .B2(n14457), .A(n14456), .ZN(SUB_1596_U57) );
  OAI21_X1 U16276 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(SUB_1596_U55) );
  AOI21_X1 U16277 ( .B1(n14847), .B2(n14463), .A(n14462), .ZN(SUB_1596_U54) );
  OAI21_X1 U16278 ( .B1(n14466), .B2(n14465), .A(n14464), .ZN(n14467) );
  XNOR2_X1 U16279 ( .A(n14467), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U16280 ( .A(n14468), .ZN(n14474) );
  AOI22_X1 U16281 ( .A1(n14472), .A2(n14471), .B1(n14470), .B2(n14469), .ZN(
        n14473) );
  NAND2_X1 U16282 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  AOI22_X1 U16283 ( .A1(n14684), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n14475), 
        .B2(n14700), .ZN(n14476) );
  OAI21_X1 U16284 ( .B1(n14698), .B2(n14477), .A(n14476), .ZN(P1_U3280) );
  OAI21_X1 U16285 ( .B1(n14479), .B2(n15294), .A(n14478), .ZN(SUB_1596_U63) );
  NOR2_X1 U16286 ( .A1(n14481), .A2(n14480), .ZN(n14482) );
  AOI21_X1 U16287 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14483), .A(n14482), 
        .ZN(n14490) );
  XNOR2_X1 U16288 ( .A(n14487), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14488) );
  XNOR2_X1 U16289 ( .A(n14488), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14489) );
  OAI21_X1 U16290 ( .B1(n14492), .B2(n15173), .A(n14491), .ZN(n14517) );
  OAI22_X1 U16291 ( .A1(n15196), .A2(n14517), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15199), .ZN(n14493) );
  INV_X1 U16292 ( .A(n14493), .ZN(P3_U3489) );
  INV_X1 U16293 ( .A(n14494), .ZN(n14495) );
  OAI22_X1 U16294 ( .A1(n14495), .A2(n15179), .B1(n7420), .B2(n15173), .ZN(
        n14496) );
  NOR2_X1 U16295 ( .A1(n14497), .A2(n14496), .ZN(n14519) );
  AOI22_X1 U16296 ( .A1(n15199), .A2(n14519), .B1(n14498), .B2(n15196), .ZN(
        P3_U3474) );
  OAI22_X1 U16297 ( .A1(n14500), .A2(n15179), .B1(n14499), .B2(n15173), .ZN(
        n14501) );
  NOR2_X1 U16298 ( .A1(n14502), .A2(n14501), .ZN(n14521) );
  INV_X1 U16299 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U16300 ( .A1(n15199), .A2(n14521), .B1(n14503), .B2(n15196), .ZN(
        P3_U3473) );
  OAI22_X1 U16301 ( .A1(n14505), .A2(n15179), .B1(n14504), .B2(n15173), .ZN(
        n14506) );
  NOR2_X1 U16302 ( .A1(n14507), .A2(n14506), .ZN(n14523) );
  AOI22_X1 U16303 ( .A1(n15199), .A2(n14523), .B1(n14508), .B2(n15196), .ZN(
        P3_U3472) );
  NOR2_X1 U16304 ( .A1(n14509), .A2(n15179), .ZN(n14511) );
  AOI211_X1 U16305 ( .C1(n15184), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14525) );
  AOI22_X1 U16306 ( .A1(n15199), .A2(n14525), .B1(n11327), .B2(n15196), .ZN(
        P3_U3471) );
  NOR2_X1 U16307 ( .A1(n15173), .A2(n14513), .ZN(n14515) );
  AOI211_X1 U16308 ( .C1(n15177), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        n14527) );
  AOI22_X1 U16309 ( .A1(n15199), .A2(n14527), .B1(n15343), .B2(n15196), .ZN(
        P3_U3470) );
  OAI22_X1 U16310 ( .A1(n15185), .A2(P3_REG0_REG_30__SCAN_IN), .B1(n14517), 
        .B2(n15187), .ZN(n14518) );
  INV_X1 U16311 ( .A(n14518), .ZN(P3_U3457) );
  INV_X1 U16312 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14520) );
  AOI22_X1 U16313 ( .A1(n15187), .A2(n14520), .B1(n14519), .B2(n15185), .ZN(
        P3_U3435) );
  INV_X1 U16314 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14522) );
  AOI22_X1 U16315 ( .A1(n15187), .A2(n14522), .B1(n14521), .B2(n15185), .ZN(
        P3_U3432) );
  INV_X1 U16316 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U16317 ( .A1(n15187), .A2(n14524), .B1(n14523), .B2(n15185), .ZN(
        P3_U3429) );
  INV_X1 U16318 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U16319 ( .A1(n15187), .A2(n14526), .B1(n14525), .B2(n15185), .ZN(
        P3_U3426) );
  INV_X1 U16320 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U16321 ( .A1(n15187), .A2(n14528), .B1(n14527), .B2(n15185), .ZN(
        P3_U3423) );
  NAND2_X1 U16322 ( .A1(n14530), .A2(n14529), .ZN(n14531) );
  NAND2_X1 U16323 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  AOI222_X1 U16324 ( .A1(n14782), .A2(n14536), .B1(n14535), .B2(n14534), .C1(
        n14533), .C2(n14788), .ZN(n14537) );
  NAND2_X1 U16325 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14897)
         );
  OAI211_X1 U16326 ( .C1(n14797), .C2(n14538), .A(n14537), .B(n14897), .ZN(
        P2_U3198) );
  OAI22_X1 U16327 ( .A1(n14554), .A2(n14539), .B1(n14553), .B2(n14551), .ZN(
        n14547) );
  AOI21_X1 U16328 ( .B1(n14542), .B2(n14541), .A(n14540), .ZN(n14543) );
  INV_X1 U16329 ( .A(n14543), .ZN(n14545) );
  AOI21_X1 U16330 ( .B1(n14545), .B2(n14544), .A(n14559), .ZN(n14546) );
  AOI211_X1 U16331 ( .C1(n14606), .C2(n14564), .A(n14547), .B(n14546), .ZN(
        n14549) );
  OAI211_X1 U16332 ( .C1(n14568), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        P1_U3215) );
  OAI22_X1 U16333 ( .A1(n14554), .A2(n14553), .B1(n14552), .B2(n14551), .ZN(
        n14563) );
  INV_X1 U16334 ( .A(n14555), .ZN(n14558) );
  OAI21_X1 U16335 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14561) );
  AOI21_X1 U16336 ( .B1(n14561), .B2(n14560), .A(n14559), .ZN(n14562) );
  AOI211_X1 U16337 ( .C1(n14598), .C2(n14564), .A(n14563), .B(n14562), .ZN(
        n14566) );
  OAI211_X1 U16338 ( .C1(n14568), .C2(n14567), .A(n14566), .B(n14565), .ZN(
        P1_U3226) );
  XNOR2_X1 U16339 ( .A(n14569), .B(n14583), .ZN(n14571) );
  NOR2_X1 U16340 ( .A1(n14571), .A2(n14570), .ZN(n14592) );
  AND2_X1 U16341 ( .A1(n14573), .A2(n14572), .ZN(n14574) );
  AOI21_X1 U16342 ( .B1(n14576), .B2(n14575), .A(n14574), .ZN(n14589) );
  INV_X1 U16343 ( .A(n14589), .ZN(n14577) );
  AOI211_X1 U16344 ( .C1(n14683), .C2(n14578), .A(n14577), .B(n14684), .ZN(
        n14579) );
  OAI21_X1 U16345 ( .B1(n14591), .B2(n14580), .A(n14579), .ZN(n14581) );
  OAI22_X1 U16346 ( .A1(n14592), .A2(n14581), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n14700), .ZN(n14588) );
  XOR2_X1 U16347 ( .A(n14582), .B(n14583), .Z(n14594) );
  OAI211_X1 U16348 ( .C1(n14585), .C2(n14591), .A(n14584), .B(n14707), .ZN(
        n14590) );
  INV_X1 U16349 ( .A(n14590), .ZN(n14586) );
  AOI22_X1 U16350 ( .A1(n14594), .A2(n14712), .B1(n14711), .B2(n14586), .ZN(
        n14587) );
  NAND2_X1 U16351 ( .A1(n14588), .A2(n14587), .ZN(P1_U3276) );
  OAI211_X1 U16352 ( .C1(n14591), .C2(n14746), .A(n14590), .B(n14589), .ZN(
        n14593) );
  AOI211_X1 U16353 ( .C1(n14594), .C2(n14762), .A(n14593), .B(n14592), .ZN(
        n14620) );
  AOI22_X1 U16354 ( .A1(n14772), .A2(n14620), .B1(n11390), .B2(n6820), .ZN(
        P1_U3545) );
  INV_X1 U16355 ( .A(n14595), .ZN(n14600) );
  AOI211_X1 U16356 ( .C1(n14598), .C2(n14755), .A(n14597), .B(n14596), .ZN(
        n14599) );
  OAI21_X1 U16357 ( .B1(n14600), .B2(n14609), .A(n14599), .ZN(n14601) );
  AOI21_X1 U16358 ( .B1(n14751), .B2(n14602), .A(n14601), .ZN(n14622) );
  AOI22_X1 U16359 ( .A1(n14772), .A2(n14622), .B1(n14603), .B2(n6820), .ZN(
        P1_U3544) );
  AOI211_X1 U16360 ( .C1(n14606), .C2(n14755), .A(n14605), .B(n14604), .ZN(
        n14607) );
  OAI21_X1 U16361 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14610) );
  AOI21_X1 U16362 ( .B1(n14751), .B2(n14611), .A(n14610), .ZN(n14623) );
  AOI22_X1 U16363 ( .A1(n14772), .A2(n14623), .B1(n14612), .B2(n6820), .ZN(
        P1_U3542) );
  OAI21_X1 U16364 ( .B1(n14614), .B2(n14746), .A(n14613), .ZN(n14616) );
  AOI211_X1 U16365 ( .C1(n14762), .C2(n14617), .A(n14616), .B(n14615), .ZN(
        n14625) );
  AOI22_X1 U16366 ( .A1(n14772), .A2(n14625), .B1(n14618), .B2(n6820), .ZN(
        P1_U3539) );
  INV_X1 U16367 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14619) );
  AOI22_X1 U16368 ( .A1(n14764), .A2(n14620), .B1(n14619), .B2(n14763), .ZN(
        P1_U3510) );
  INV_X1 U16369 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U16370 ( .A1(n14764), .A2(n14622), .B1(n14621), .B2(n14763), .ZN(
        P1_U3507) );
  INV_X1 U16371 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U16372 ( .A1(n14764), .A2(n14623), .B1(n15239), .B2(n14763), .ZN(
        P1_U3501) );
  INV_X1 U16373 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U16374 ( .A1(n14764), .A2(n14625), .B1(n14624), .B2(n14763), .ZN(
        P1_U3492) );
  OAI21_X1 U16375 ( .B1(n14628), .B2(n14627), .A(n14626), .ZN(n14629) );
  XNOR2_X1 U16376 ( .A(n14629), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  AOI21_X1 U16377 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14633) );
  XOR2_X1 U16378 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14633), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16379 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  XOR2_X1 U16380 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14637), .Z(SUB_1596_U67)
         );
  OAI222_X1 U16381 ( .A1(n14642), .A2(n14641), .B1(n14642), .B2(n14640), .C1(
        n14639), .C2(n14638), .ZN(SUB_1596_U66) );
  OAI222_X1 U16382 ( .A1(n14647), .A2(n14646), .B1(n14647), .B2(n14645), .C1(
        n14644), .C2(n14643), .ZN(SUB_1596_U65) );
  OAI21_X1 U16383 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(n14651) );
  XNOR2_X1 U16384 ( .A(n14651), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AOI21_X1 U16385 ( .B1(n6415), .B2(n9478), .A(n14652), .ZN(n14654) );
  XNOR2_X1 U16386 ( .A(n14654), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16387 ( .A1(n14655), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14656) );
  OAI21_X1 U16388 ( .B1(n14658), .B2(n14657), .A(n14656), .ZN(P1_U3243) );
  AOI21_X1 U16389 ( .B1(n14660), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14659), 
        .ZN(n14670) );
  AOI21_X1 U16390 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14662), .A(n14661), 
        .ZN(n14664) );
  OR2_X1 U16391 ( .A1(n14664), .A2(n14663), .ZN(n14668) );
  NAND2_X1 U16392 ( .A1(n14666), .A2(n14665), .ZN(n14667) );
  OAI211_X1 U16393 ( .C1(n14670), .C2(n14669), .A(n14668), .B(n14667), .ZN(
        n14671) );
  INV_X1 U16394 ( .A(n14671), .ZN(n14673) );
  OAI211_X1 U16395 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        P1_U3258) );
  OAI21_X1 U16396 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(n14680) );
  AOI21_X1 U16397 ( .B1(n14680), .B2(n14751), .A(n14679), .ZN(n14745) );
  INV_X1 U16398 ( .A(n14681), .ZN(n14682) );
  AOI222_X1 U16399 ( .A1(n14688), .A2(n14702), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n14684), .C1(n14683), .C2(n14682), .ZN(n14693) );
  XNOR2_X1 U16400 ( .A(n14686), .B(n14685), .ZN(n14749) );
  INV_X1 U16401 ( .A(n14687), .ZN(n14690) );
  INV_X1 U16402 ( .A(n14688), .ZN(n14747) );
  OAI211_X1 U16403 ( .C1(n14690), .C2(n14747), .A(n14707), .B(n14689), .ZN(
        n14744) );
  INV_X1 U16404 ( .A(n14744), .ZN(n14691) );
  AOI22_X1 U16405 ( .A1(n14749), .A2(n14712), .B1(n14711), .B2(n14691), .ZN(
        n14692) );
  OAI211_X1 U16406 ( .C1(n14684), .C2(n14745), .A(n14693), .B(n14692), .ZN(
        P1_U3284) );
  XNOR2_X1 U16407 ( .A(n14695), .B(n14694), .ZN(n14697) );
  AOI21_X1 U16408 ( .B1(n14697), .B2(n14751), .A(n14696), .ZN(n14725) );
  OAI22_X1 U16409 ( .A1(n14700), .A2(n14699), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14698), .ZN(n14701) );
  AOI21_X1 U16410 ( .B1(n14702), .B2(n14705), .A(n14701), .ZN(n14714) );
  XNOR2_X1 U16411 ( .A(n14704), .B(n14703), .ZN(n14728) );
  NAND2_X1 U16412 ( .A1(n14706), .A2(n14705), .ZN(n14708) );
  NAND2_X1 U16413 ( .A1(n14708), .A2(n14707), .ZN(n14709) );
  NOR2_X1 U16414 ( .A1(n14710), .A2(n14709), .ZN(n14723) );
  AOI22_X1 U16415 ( .A1(n14712), .A2(n14728), .B1(n14711), .B2(n14723), .ZN(
        n14713) );
  OAI211_X1 U16416 ( .C1(n14684), .C2(n14725), .A(n14714), .B(n14713), .ZN(
        P1_U3290) );
  AND2_X1 U16417 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n6405), .ZN(P1_U3294) );
  AND2_X1 U16418 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n6405), .ZN(P1_U3295) );
  AND2_X1 U16419 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n6405), .ZN(P1_U3296) );
  AND2_X1 U16420 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n6405), .ZN(P1_U3297) );
  AND2_X1 U16421 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n6405), .ZN(P1_U3298) );
  AND2_X1 U16422 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n6405), .ZN(P1_U3299) );
  AND2_X1 U16423 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n6405), .ZN(P1_U3300) );
  AND2_X1 U16424 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n6405), .ZN(P1_U3301) );
  AND2_X1 U16425 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n6405), .ZN(P1_U3302) );
  AND2_X1 U16426 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n6405), .ZN(P1_U3303) );
  AND2_X1 U16427 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n6405), .ZN(P1_U3304) );
  AND2_X1 U16428 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n6405), .ZN(P1_U3305) );
  AND2_X1 U16429 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n6405), .ZN(P1_U3306) );
  AND2_X1 U16430 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n6405), .ZN(P1_U3307) );
  AND2_X1 U16431 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n6405), .ZN(P1_U3308) );
  AND2_X1 U16432 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n6405), .ZN(P1_U3309) );
  AND2_X1 U16433 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n6405), .ZN(P1_U3310) );
  AND2_X1 U16434 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n6405), .ZN(P1_U3311) );
  AND2_X1 U16435 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n6405), .ZN(P1_U3312) );
  AND2_X1 U16436 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n6405), .ZN(P1_U3313) );
  AND2_X1 U16437 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n6405), .ZN(P1_U3314) );
  AND2_X1 U16438 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n6405), .ZN(P1_U3315) );
  AND2_X1 U16439 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n6405), .ZN(P1_U3316) );
  AND2_X1 U16440 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n6405), .ZN(P1_U3318) );
  AND2_X1 U16441 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n6405), .ZN(P1_U3319) );
  AND2_X1 U16442 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n6405), .ZN(P1_U3320) );
  AND2_X1 U16443 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n6405), .ZN(P1_U3321) );
  AND2_X1 U16444 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n6405), .ZN(P1_U3322) );
  AND2_X1 U16445 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n6405), .ZN(P1_U3323) );
  INV_X1 U16446 ( .A(n14715), .ZN(n14722) );
  INV_X1 U16447 ( .A(n14716), .ZN(n14719) );
  OAI22_X1 U16448 ( .A1(n14719), .A2(n14718), .B1(n14717), .B2(n14746), .ZN(
        n14721) );
  AOI211_X1 U16449 ( .C1(n14762), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        n14765) );
  AOI22_X1 U16450 ( .A1(n14764), .A2(n14765), .B1(n9274), .B2(n14763), .ZN(
        P1_U3462) );
  INV_X1 U16451 ( .A(n14723), .ZN(n14724) );
  OAI21_X1 U16452 ( .B1(n6990), .B2(n14746), .A(n14724), .ZN(n14727) );
  INV_X1 U16453 ( .A(n14725), .ZN(n14726) );
  AOI211_X1 U16454 ( .C1(n14762), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14766) );
  INV_X1 U16455 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14729) );
  AOI22_X1 U16456 ( .A1(n14764), .A2(n14766), .B1(n14729), .B2(n14763), .ZN(
        P1_U3468) );
  OAI21_X1 U16457 ( .B1(n14731), .B2(n14746), .A(n14730), .ZN(n14733) );
  AOI211_X1 U16458 ( .C1(n14762), .C2(n14734), .A(n14733), .B(n14732), .ZN(
        n14767) );
  INV_X1 U16459 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U16460 ( .A1(n14764), .A2(n14767), .B1(n14735), .B2(n14763), .ZN(
        P1_U3471) );
  AOI21_X1 U16461 ( .B1(n14737), .B2(n14755), .A(n14736), .ZN(n14739) );
  NAND3_X1 U16462 ( .A1(n14740), .A2(n14739), .A3(n14738), .ZN(n14741) );
  AOI21_X1 U16463 ( .B1(n14762), .B2(n14742), .A(n14741), .ZN(n14768) );
  INV_X1 U16464 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14743) );
  AOI22_X1 U16465 ( .A1(n14764), .A2(n14768), .B1(n14743), .B2(n14763), .ZN(
        P1_U3483) );
  OAI211_X1 U16466 ( .C1(n14747), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14748) );
  AOI21_X1 U16467 ( .B1(n14762), .B2(n14749), .A(n14748), .ZN(n14769) );
  INV_X1 U16468 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U16469 ( .A1(n14764), .A2(n14769), .B1(n14750), .B2(n14763), .ZN(
        P1_U3486) );
  NAND3_X1 U16470 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(n14759) );
  AOI21_X1 U16471 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14758) );
  NAND3_X1 U16472 ( .A1(n14759), .A2(n14758), .A3(n14757), .ZN(n14760) );
  AOI21_X1 U16473 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14771) );
  AOI22_X1 U16474 ( .A1(n14764), .A2(n14771), .B1(n10564), .B2(n14763), .ZN(
        P1_U3489) );
  AOI22_X1 U16475 ( .A1(n14772), .A2(n14765), .B1(n9289), .B2(n6820), .ZN(
        P1_U3529) );
  AOI22_X1 U16476 ( .A1(n14772), .A2(n14766), .B1(n9611), .B2(n6820), .ZN(
        P1_U3531) );
  AOI22_X1 U16477 ( .A1(n14772), .A2(n14767), .B1(n9933), .B2(n6820), .ZN(
        P1_U3532) );
  AOI22_X1 U16478 ( .A1(n14772), .A2(n14768), .B1(n10094), .B2(n6820), .ZN(
        P1_U3536) );
  AOI22_X1 U16479 ( .A1(n14772), .A2(n14769), .B1(n15311), .B2(n6820), .ZN(
        P1_U3537) );
  AOI22_X1 U16480 ( .A1(n14772), .A2(n14771), .B1(n14770), .B2(n6820), .ZN(
        P1_U3538) );
  NOR2_X1 U16481 ( .A1(n14923), .A2(n14773), .ZN(P2_U3087) );
  INV_X1 U16482 ( .A(n14774), .ZN(n14775) );
  OAI22_X1 U16483 ( .A1(n14787), .A2(n14775), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8409), .ZN(n14781) );
  AOI211_X1 U16484 ( .C1(n14779), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        n14780) );
  AOI211_X1 U16485 ( .C1(n14783), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        n14784) );
  OAI21_X1 U16486 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14797), .A(n14784), .ZN(
        P2_U3190) );
  OAI21_X1 U16487 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14793) );
  OAI211_X1 U16488 ( .C1(n14790), .C2(n14789), .A(n11293), .B(n14788), .ZN(
        n14791) );
  INV_X1 U16489 ( .A(n14791), .ZN(n14792) );
  AOI211_X1 U16490 ( .C1(n14795), .C2(n14794), .A(n14793), .B(n14792), .ZN(
        n14796) );
  OAI21_X1 U16491 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(P2_U3206) );
  MUX2_X1 U16492 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9336), .S(n14809), .Z(
        n14799) );
  NAND3_X1 U16493 ( .A1(n14801), .A2(n14800), .A3(n14799), .ZN(n14802) );
  NAND3_X1 U16494 ( .A1(n14917), .A2(n14816), .A3(n14802), .ZN(n14808) );
  MUX2_X1 U16495 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9358), .S(n14809), .Z(
        n14803) );
  NAND3_X1 U16496 ( .A1(n14805), .A2(n14804), .A3(n14803), .ZN(n14806) );
  NAND3_X1 U16497 ( .A1(n14925), .A2(n14822), .A3(n14806), .ZN(n14807) );
  OAI211_X1 U16498 ( .C1(n14930), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        n14810) );
  INV_X1 U16499 ( .A(n14810), .ZN(n14812) );
  OAI211_X1 U16500 ( .C1(n14846), .C2(n14813), .A(n14812), .B(n14811), .ZN(
        P2_U3218) );
  MUX2_X1 U16501 ( .A(n10402), .B(P2_REG2_REG_5__SCAN_IN), .S(n14819), .Z(
        n14814) );
  NAND3_X1 U16502 ( .A1(n14816), .A2(n14815), .A3(n14814), .ZN(n14817) );
  NAND3_X1 U16503 ( .A1(n14917), .A2(n14818), .A3(n14817), .ZN(n14826) );
  MUX2_X1 U16504 ( .A(n9361), .B(P2_REG1_REG_5__SCAN_IN), .S(n14819), .Z(
        n14820) );
  NAND3_X1 U16505 ( .A1(n14822), .A2(n14821), .A3(n14820), .ZN(n14823) );
  NAND3_X1 U16506 ( .A1(n14925), .A2(n14824), .A3(n14823), .ZN(n14825) );
  OAI211_X1 U16507 ( .C1(n14930), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        n14828) );
  INV_X1 U16508 ( .A(n14828), .ZN(n14830) );
  OAI211_X1 U16509 ( .C1(n14846), .C2(n15359), .A(n14830), .B(n14829), .ZN(
        P2_U3219) );
  NOR2_X1 U16510 ( .A1(n14832), .A2(n14831), .ZN(n14833) );
  OAI21_X1 U16511 ( .B1(n14834), .B2(n14833), .A(n14925), .ZN(n14841) );
  NAND2_X1 U16512 ( .A1(n14836), .A2(n14835), .ZN(n14837) );
  NAND2_X1 U16513 ( .A1(n14838), .A2(n14837), .ZN(n14839) );
  NAND2_X1 U16514 ( .A1(n14917), .A2(n14839), .ZN(n14840) );
  OAI211_X1 U16515 ( .C1(n14930), .C2(n14842), .A(n14841), .B(n14840), .ZN(
        n14843) );
  INV_X1 U16516 ( .A(n14843), .ZN(n14845) );
  NAND2_X1 U16517 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14844) );
  OAI211_X1 U16518 ( .C1(n14847), .C2(n14846), .A(n14845), .B(n14844), .ZN(
        P2_U3223) );
  AOI22_X1 U16519 ( .A1(n14906), .A2(n14848), .B1(n14923), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U16520 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14859)
         );
  OAI211_X1 U16521 ( .C1(n14851), .C2(n14850), .A(n14849), .B(n14925), .ZN(
        n14858) );
  AOI211_X1 U16522 ( .C1(n14855), .C2(n14854), .A(n14853), .B(n14852), .ZN(
        n14856) );
  INV_X1 U16523 ( .A(n14856), .ZN(n14857) );
  NAND4_X1 U16524 ( .A1(n14860), .A2(n14859), .A3(n14858), .A4(n14857), .ZN(
        P2_U3224) );
  AOI22_X1 U16525 ( .A1(n14906), .A2(n14861), .B1(n14923), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n14873) );
  NAND2_X1 U16526 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14872)
         );
  OAI21_X1 U16527 ( .B1(n14864), .B2(n14863), .A(n14862), .ZN(n14865) );
  NAND2_X1 U16528 ( .A1(n14865), .A2(n14917), .ZN(n14871) );
  OAI21_X1 U16529 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14869) );
  NAND2_X1 U16530 ( .A1(n14869), .A2(n14925), .ZN(n14870) );
  NAND4_X1 U16531 ( .A1(n14873), .A2(n14872), .A3(n14871), .A4(n14870), .ZN(
        P2_U3226) );
  AOI22_X1 U16532 ( .A1(n14923), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14883) );
  OAI211_X1 U16533 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n14875), .A(n14917), 
        .B(n14874), .ZN(n14882) );
  NAND2_X1 U16534 ( .A1(n14876), .A2(n14906), .ZN(n14881) );
  XOR2_X1 U16535 ( .A(n14878), .B(n14877), .Z(n14879) );
  NAND2_X1 U16536 ( .A1(n14879), .A2(n14925), .ZN(n14880) );
  NAND4_X1 U16537 ( .A1(n14883), .A2(n14882), .A3(n14881), .A4(n14880), .ZN(
        P2_U3228) );
  AOI22_X1 U16538 ( .A1(n14923), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14892) );
  NAND2_X1 U16539 ( .A1(n14906), .A2(n14884), .ZN(n14891) );
  OAI211_X1 U16540 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14886), .A(n14917), 
        .B(n14885), .ZN(n14890) );
  XNOR2_X1 U16541 ( .A(n14887), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n14888) );
  NAND2_X1 U16542 ( .A1(n14888), .A2(n14925), .ZN(n14889) );
  NAND4_X1 U16543 ( .A1(n14892), .A2(n14891), .A3(n14890), .A4(n14889), .ZN(
        P2_U3229) );
  OAI211_X1 U16544 ( .C1(n14895), .C2(n14894), .A(n14925), .B(n14893), .ZN(
        n14896) );
  NAND2_X1 U16545 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  AOI21_X1 U16546 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n14923), .A(n14898), 
        .ZN(n14903) );
  OAI211_X1 U16547 ( .C1(n14901), .C2(n14900), .A(n14917), .B(n14899), .ZN(
        n14902) );
  OAI211_X1 U16548 ( .C1(n14930), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        P2_U3230) );
  AOI22_X1 U16549 ( .A1(n14923), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14916) );
  NAND2_X1 U16550 ( .A1(n14906), .A2(n14905), .ZN(n14915) );
  XOR2_X1 U16551 ( .A(n14908), .B(n14907), .Z(n14909) );
  NAND2_X1 U16552 ( .A1(n14925), .A2(n14909), .ZN(n14914) );
  OAI211_X1 U16553 ( .C1(n14912), .C2(n14911), .A(n14917), .B(n14910), .ZN(
        n14913) );
  NAND4_X1 U16554 ( .A1(n14916), .A2(n14915), .A3(n14914), .A4(n14913), .ZN(
        P2_U3231) );
  OAI221_X1 U16555 ( .B1(n14919), .B2(P2_REG2_REG_18__SCAN_IN), .C1(n14919), 
        .C2(n14918), .A(n14917), .ZN(n14920) );
  NAND2_X1 U16556 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  AOI21_X1 U16557 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n14923), .A(n14922), 
        .ZN(n14928) );
  OAI211_X1 U16558 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14926), .A(n14925), 
        .B(n14924), .ZN(n14927) );
  OAI211_X1 U16559 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        P2_U3232) );
  INV_X1 U16560 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U16561 ( .A1(n14932), .A2(n14931), .ZN(n14936) );
  NAND2_X1 U16562 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  OAI211_X1 U16563 ( .C1(n14938), .C2(n14937), .A(n14936), .B(n14935), .ZN(
        n14940) );
  NOR2_X1 U16564 ( .A1(n14940), .A2(n14939), .ZN(n14942) );
  AOI22_X1 U16565 ( .A1(n14943), .A2(n9417), .B1(n14942), .B2(n14941), .ZN(
        P2_U3265) );
  INV_X1 U16566 ( .A(n14979), .ZN(n14976) );
  INV_X1 U16567 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16568 ( .A1(n14973), .A2(n15337), .ZN(P2_U3266) );
  INV_X1 U16569 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15319) );
  NOR2_X1 U16570 ( .A1(n14973), .A2(n15319), .ZN(P2_U3267) );
  INV_X1 U16571 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14945) );
  NOR2_X1 U16572 ( .A1(n14973), .A2(n14945), .ZN(P2_U3268) );
  INV_X1 U16573 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U16574 ( .A1(n14969), .A2(n14946), .ZN(P2_U3269) );
  INV_X1 U16575 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14947) );
  NOR2_X1 U16576 ( .A1(n14969), .A2(n14947), .ZN(P2_U3270) );
  INV_X1 U16577 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14948) );
  NOR2_X1 U16578 ( .A1(n14969), .A2(n14948), .ZN(P2_U3271) );
  INV_X1 U16579 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14949) );
  NOR2_X1 U16580 ( .A1(n14969), .A2(n14949), .ZN(P2_U3272) );
  INV_X1 U16581 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14950) );
  NOR2_X1 U16582 ( .A1(n14969), .A2(n14950), .ZN(P2_U3273) );
  INV_X1 U16583 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U16584 ( .A1(n14969), .A2(n15338), .ZN(P2_U3274) );
  INV_X1 U16585 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14951) );
  NOR2_X1 U16586 ( .A1(n14969), .A2(n14951), .ZN(P2_U3275) );
  INV_X1 U16587 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14952) );
  NOR2_X1 U16588 ( .A1(n14969), .A2(n14952), .ZN(P2_U3276) );
  INV_X1 U16589 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14953) );
  NOR2_X1 U16590 ( .A1(n14969), .A2(n14953), .ZN(P2_U3277) );
  INV_X1 U16591 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14954) );
  NOR2_X1 U16592 ( .A1(n14973), .A2(n14954), .ZN(P2_U3278) );
  INV_X1 U16593 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14955) );
  NOR2_X1 U16594 ( .A1(n14973), .A2(n14955), .ZN(P2_U3279) );
  INV_X1 U16595 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14956) );
  NOR2_X1 U16596 ( .A1(n14973), .A2(n14956), .ZN(P2_U3280) );
  INV_X1 U16597 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14957) );
  NOR2_X1 U16598 ( .A1(n14973), .A2(n14957), .ZN(P2_U3281) );
  INV_X1 U16599 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14958) );
  NOR2_X1 U16600 ( .A1(n14973), .A2(n14958), .ZN(P2_U3282) );
  INV_X1 U16601 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14959) );
  NOR2_X1 U16602 ( .A1(n14973), .A2(n14959), .ZN(P2_U3283) );
  INV_X1 U16603 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14960) );
  NOR2_X1 U16604 ( .A1(n14973), .A2(n14960), .ZN(P2_U3284) );
  INV_X1 U16605 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14961) );
  NOR2_X1 U16606 ( .A1(n14973), .A2(n14961), .ZN(P2_U3285) );
  INV_X1 U16607 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14962) );
  NOR2_X1 U16608 ( .A1(n14973), .A2(n14962), .ZN(P2_U3286) );
  INV_X1 U16609 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14963) );
  NOR2_X1 U16610 ( .A1(n14973), .A2(n14963), .ZN(P2_U3287) );
  INV_X1 U16611 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14964) );
  NOR2_X1 U16612 ( .A1(n14973), .A2(n14964), .ZN(P2_U3288) );
  INV_X1 U16613 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14965) );
  NOR2_X1 U16614 ( .A1(n14973), .A2(n14965), .ZN(P2_U3289) );
  INV_X1 U16615 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14966) );
  NOR2_X1 U16616 ( .A1(n14969), .A2(n14966), .ZN(P2_U3290) );
  INV_X1 U16617 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14967) );
  NOR2_X1 U16618 ( .A1(n14973), .A2(n14967), .ZN(P2_U3291) );
  INV_X1 U16619 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14968) );
  NOR2_X1 U16620 ( .A1(n14969), .A2(n14968), .ZN(P2_U3292) );
  INV_X1 U16621 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14970) );
  NOR2_X1 U16622 ( .A1(n14973), .A2(n14970), .ZN(P2_U3293) );
  INV_X1 U16623 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14971) );
  NOR2_X1 U16624 ( .A1(n14973), .A2(n14971), .ZN(P2_U3294) );
  INV_X1 U16625 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14972) );
  NOR2_X1 U16626 ( .A1(n14973), .A2(n14972), .ZN(P2_U3295) );
  OAI21_X1 U16627 ( .B1(n14979), .B2(n14975), .A(n14974), .ZN(P2_U3416) );
  AOI22_X1 U16628 ( .A1(n14979), .A2(n14978), .B1(n14977), .B2(n14976), .ZN(
        P2_U3417) );
  AOI22_X1 U16629 ( .A1(n15066), .A2(n14980), .B1(n8338), .B2(n15065), .ZN(
        P2_U3430) );
  INV_X1 U16630 ( .A(n14983), .ZN(n14986) );
  AOI211_X1 U16631 ( .C1(n15053), .C2(n9053), .A(n14982), .B(n14981), .ZN(
        n14985) );
  NAND2_X1 U16632 ( .A1(n14983), .A2(n15064), .ZN(n14984) );
  OAI211_X1 U16633 ( .C1(n14986), .C2(n15059), .A(n14985), .B(n14984), .ZN(
        n14987) );
  AOI21_X1 U16634 ( .B1(n14988), .B2(n15026), .A(n14987), .ZN(n15068) );
  AOI22_X1 U16635 ( .A1(n15066), .A2(n15068), .B1(n8300), .B2(n15065), .ZN(
        P2_U3433) );
  OAI21_X1 U16636 ( .B1(n9052), .B2(n15046), .A(n14989), .ZN(n14990) );
  AOI21_X1 U16637 ( .B1(n14991), .B2(n15013), .A(n14990), .ZN(n14992) );
  AND2_X1 U16638 ( .A1(n14993), .A2(n14992), .ZN(n15069) );
  AOI22_X1 U16639 ( .A1(n15066), .A2(n15069), .B1(n8362), .B2(n15065), .ZN(
        P2_U3436) );
  OAI21_X1 U16640 ( .B1(n14995), .B2(n15046), .A(n14994), .ZN(n14997) );
  AOI211_X1 U16641 ( .C1(n14999), .C2(n14998), .A(n14997), .B(n14996), .ZN(
        n15070) );
  INV_X1 U16642 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U16643 ( .A1(n15066), .A2(n15070), .B1(n15000), .B2(n15065), .ZN(
        P2_U3442) );
  AND2_X1 U16644 ( .A1(n15001), .A2(n15053), .ZN(n15002) );
  OR2_X1 U16645 ( .A1(n15003), .A2(n15002), .ZN(n15004) );
  AOI21_X1 U16646 ( .B1(n15005), .B2(n15013), .A(n15004), .ZN(n15006) );
  AND2_X1 U16647 ( .A1(n15007), .A2(n15006), .ZN(n15071) );
  INV_X1 U16648 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16649 ( .A1(n15066), .A2(n15071), .B1(n15008), .B2(n15065), .ZN(
        P2_U3445) );
  AOI21_X1 U16650 ( .B1(n15014), .B2(n15064), .A(n15009), .ZN(n15016) );
  OAI21_X1 U16651 ( .B1(n15011), .B2(n15046), .A(n15010), .ZN(n15012) );
  AOI21_X1 U16652 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15015) );
  AND2_X1 U16653 ( .A1(n15016), .A2(n15015), .ZN(n15072) );
  INV_X1 U16654 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15017) );
  AOI22_X1 U16655 ( .A1(n15066), .A2(n15072), .B1(n15017), .B2(n15065), .ZN(
        P2_U3448) );
  AOI211_X1 U16656 ( .C1(n15053), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15021) );
  OAI21_X1 U16657 ( .B1(n15023), .B2(n15022), .A(n15021), .ZN(n15024) );
  AOI21_X1 U16658 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15073) );
  INV_X1 U16659 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15027) );
  AOI22_X1 U16660 ( .A1(n15066), .A2(n15073), .B1(n15027), .B2(n15065), .ZN(
        P2_U3451) );
  OR2_X1 U16661 ( .A1(n15028), .A2(n15059), .ZN(n15035) );
  NAND2_X1 U16662 ( .A1(n15029), .A2(n15053), .ZN(n15030) );
  AND2_X1 U16663 ( .A1(n15031), .A2(n15030), .ZN(n15032) );
  INV_X1 U16664 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U16665 ( .A1(n15066), .A2(n15074), .B1(n15036), .B2(n15065), .ZN(
        P2_U3454) );
  NOR2_X1 U16666 ( .A1(n15037), .A2(n15059), .ZN(n15043) );
  INV_X1 U16667 ( .A(n15038), .ZN(n15040) );
  OAI21_X1 U16668 ( .B1(n15040), .B2(n15046), .A(n15039), .ZN(n15041) );
  NOR4_X1 U16669 ( .A1(n15043), .A2(n7106), .A3(n15042), .A4(n15041), .ZN(
        n15076) );
  AOI22_X1 U16670 ( .A1(n15066), .A2(n15076), .B1(n8542), .B2(n15065), .ZN(
        P2_U3457) );
  NOR2_X1 U16671 ( .A1(n15044), .A2(n15059), .ZN(n15050) );
  OAI21_X1 U16672 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15048) );
  NOR4_X1 U16673 ( .A1(n15050), .A2(n7107), .A3(n15049), .A4(n15048), .ZN(
        n15077) );
  INV_X1 U16674 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U16675 ( .A1(n15066), .A2(n15077), .B1(n15051), .B2(n15065), .ZN(
        P2_U3460) );
  AOI21_X1 U16676 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15056) );
  OAI211_X1 U16677 ( .C1(n15058), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15062) );
  NOR2_X1 U16678 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  AOI211_X1 U16679 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15080) );
  AOI22_X1 U16680 ( .A1(n15066), .A2(n15080), .B1(n8590), .B2(n15065), .ZN(
        P2_U3463) );
  AOI22_X1 U16681 ( .A1(n15081), .A2(n15068), .B1(n15067), .B2(n15078), .ZN(
        P2_U3500) );
  AOI22_X1 U16682 ( .A1(n15081), .A2(n15069), .B1(n9354), .B2(n15078), .ZN(
        P2_U3501) );
  AOI22_X1 U16683 ( .A1(n15081), .A2(n15070), .B1(n9358), .B2(n15078), .ZN(
        P2_U3503) );
  AOI22_X1 U16684 ( .A1(n15081), .A2(n15071), .B1(n9361), .B2(n15078), .ZN(
        P2_U3504) );
  AOI22_X1 U16685 ( .A1(n15081), .A2(n15072), .B1(n9364), .B2(n15078), .ZN(
        P2_U3505) );
  AOI22_X1 U16686 ( .A1(n15081), .A2(n15073), .B1(n9367), .B2(n15078), .ZN(
        P2_U3506) );
  AOI22_X1 U16687 ( .A1(n15081), .A2(n15074), .B1(n9546), .B2(n15078), .ZN(
        P2_U3507) );
  AOI22_X1 U16688 ( .A1(n15081), .A2(n15076), .B1(n15075), .B2(n15078), .ZN(
        P2_U3508) );
  AOI22_X1 U16689 ( .A1(n15081), .A2(n15077), .B1(n9551), .B2(n15078), .ZN(
        P2_U3509) );
  AOI22_X1 U16690 ( .A1(n15081), .A2(n15080), .B1(n15079), .B2(n15078), .ZN(
        P2_U3510) );
  NOR2_X1 U16691 ( .A1(P3_U3897), .A2(n15082), .ZN(P3_U3150) );
  NAND3_X1 U16692 ( .A1(n15136), .A2(n15125), .A3(n15110), .ZN(n15087) );
  NAND2_X1 U16693 ( .A1(n15087), .A2(n15086), .ZN(n15088) );
  OAI211_X1 U16694 ( .C1(n15090), .C2(n15126), .A(n15089), .B(n15088), .ZN(
        P3_U3182) );
  INV_X1 U16695 ( .A(n15091), .ZN(n15092) );
  AOI21_X1 U16696 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15114) );
  INV_X1 U16697 ( .A(n15095), .ZN(n15105) );
  INV_X1 U16698 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15098) );
  INV_X1 U16699 ( .A(n15096), .ZN(n15097) );
  OAI21_X1 U16700 ( .B1(n15126), .B2(n15098), .A(n15097), .ZN(n15104) );
  NAND2_X1 U16701 ( .A1(n15100), .A2(n15099), .ZN(n15101) );
  AOI21_X1 U16702 ( .B1(n15102), .B2(n15101), .A(n15125), .ZN(n15103) );
  AOI211_X1 U16703 ( .C1(n15106), .C2(n15105), .A(n15104), .B(n15103), .ZN(
        n15113) );
  AOI21_X1 U16704 ( .B1(n15109), .B2(n15108), .A(n15107), .ZN(n15111) );
  OR2_X1 U16705 ( .A1(n15111), .A2(n15110), .ZN(n15112) );
  OAI211_X1 U16706 ( .C1(n15114), .C2(n15136), .A(n15113), .B(n15112), .ZN(
        P3_U3192) );
  AOI21_X1 U16707 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15137) );
  INV_X1 U16708 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15127) );
  INV_X1 U16709 ( .A(n15118), .ZN(n15119) );
  AOI21_X1 U16710 ( .B1(n15121), .B2(n15120), .A(n15119), .ZN(n15124) );
  OAI222_X1 U16711 ( .A1(n15127), .A2(n15126), .B1(n15125), .B2(n15124), .C1(
        n15123), .C2(n15122), .ZN(n15128) );
  NOR2_X1 U16712 ( .A1(n15129), .A2(n15128), .ZN(n15135) );
  OAI211_X1 U16713 ( .C1(n15133), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15134) );
  OAI211_X1 U16714 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        P3_U3194) );
  NOR2_X1 U16715 ( .A1(n15173), .A2(n10801), .ZN(n15158) );
  XNOR2_X1 U16716 ( .A(n15139), .B(n15138), .ZN(n15148) );
  XNOR2_X1 U16717 ( .A(n10804), .B(n15140), .ZN(n15159) );
  NAND2_X1 U16718 ( .A1(n15141), .A2(n15159), .ZN(n15147) );
  AOI22_X1 U16719 ( .A1(n15145), .A2(n15144), .B1(n15143), .B2(n15142), .ZN(
        n15146) );
  OAI211_X1 U16720 ( .C1(n15149), .C2(n15148), .A(n15147), .B(n15146), .ZN(
        n15157) );
  AOI21_X1 U16721 ( .B1(n15158), .B2(n15150), .A(n15157), .ZN(n15155) );
  AOI22_X1 U16722 ( .A1(n15152), .A2(n15159), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15151), .ZN(n15153) );
  OAI221_X1 U16723 ( .B1(n15156), .B2(n15155), .C1(n15154), .C2(n9802), .A(
        n15153), .ZN(P3_U3232) );
  AOI211_X1 U16724 ( .C1(n15164), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15189) );
  AOI22_X1 U16725 ( .A1(n15187), .A2(n15160), .B1(n15189), .B2(n15185), .ZN(
        P3_U3393) );
  INV_X1 U16726 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15166) );
  NOR2_X1 U16727 ( .A1(n15173), .A2(n15161), .ZN(n15163) );
  AOI211_X1 U16728 ( .C1(n15165), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15191) );
  AOI22_X1 U16729 ( .A1(n15187), .A2(n15166), .B1(n15191), .B2(n15185), .ZN(
        P3_U3399) );
  INV_X1 U16730 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U16731 ( .A1(n15177), .A2(n15168), .B1(n15167), .B2(n15184), .ZN(
        n15170) );
  AND2_X1 U16732 ( .A1(n15170), .A2(n15169), .ZN(n15193) );
  AOI22_X1 U16733 ( .A1(n15187), .A2(n15171), .B1(n15193), .B2(n15185), .ZN(
        P3_U3402) );
  INV_X1 U16734 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15178) );
  NOR2_X1 U16735 ( .A1(n15173), .A2(n15172), .ZN(n15175) );
  AOI211_X1 U16736 ( .C1(n15177), .C2(n15176), .A(n15175), .B(n15174), .ZN(
        n15195) );
  AOI22_X1 U16737 ( .A1(n15187), .A2(n15178), .B1(n15195), .B2(n15185), .ZN(
        P3_U3408) );
  INV_X1 U16738 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15186) );
  NOR3_X1 U16739 ( .A1(n6589), .A2(n15180), .A3(n15179), .ZN(n15182) );
  AOI211_X1 U16740 ( .C1(n15184), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        n15198) );
  AOI22_X1 U16741 ( .A1(n15187), .A2(n15186), .B1(n15198), .B2(n15185), .ZN(
        P3_U3420) );
  AOI22_X1 U16742 ( .A1(n15199), .A2(n15189), .B1(n15188), .B2(n15196), .ZN(
        P3_U3460) );
  AOI22_X1 U16743 ( .A1(n15199), .A2(n15191), .B1(n15190), .B2(n15196), .ZN(
        P3_U3462) );
  INV_X1 U16744 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U16745 ( .A1(n15199), .A2(n15193), .B1(n15192), .B2(n15196), .ZN(
        P3_U3463) );
  INV_X1 U16746 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U16747 ( .A1(n15199), .A2(n15195), .B1(n15194), .B2(n15196), .ZN(
        P3_U3465) );
  INV_X1 U16748 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15197) );
  AOI22_X1 U16749 ( .A1(n15199), .A2(n15198), .B1(n15197), .B2(n15196), .ZN(
        P3_U3469) );
  AOI22_X1 U16750 ( .A1(n15201), .A2(keyinput18), .B1(keyinput48), .B2(n10097), 
        .ZN(n15200) );
  OAI221_X1 U16751 ( .B1(n15201), .B2(keyinput18), .C1(n10097), .C2(keyinput48), .A(n15200), .ZN(n15210) );
  AOI22_X1 U16752 ( .A1(n15203), .A2(keyinput61), .B1(n15319), .B2(keyinput28), 
        .ZN(n15202) );
  OAI221_X1 U16753 ( .B1(n15203), .B2(keyinput61), .C1(n15319), .C2(keyinput28), .A(n15202), .ZN(n15209) );
  AOI22_X1 U16754 ( .A1(n15311), .A2(keyinput14), .B1(n7560), .B2(keyinput53), 
        .ZN(n15204) );
  OAI221_X1 U16755 ( .B1(n15311), .B2(keyinput14), .C1(n7560), .C2(keyinput53), 
        .A(n15204), .ZN(n15208) );
  XOR2_X1 U16756 ( .A(n10016), .B(keyinput58), .Z(n15206) );
  XNOR2_X1 U16757 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput38), .ZN(n15205) );
  NAND2_X1 U16758 ( .A1(n15206), .A2(n15205), .ZN(n15207) );
  NOR4_X1 U16759 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        n15252) );
  AOI22_X1 U16760 ( .A1(n15312), .A2(keyinput41), .B1(n15337), .B2(keyinput39), 
        .ZN(n15211) );
  OAI221_X1 U16761 ( .B1(n15312), .B2(keyinput41), .C1(n15337), .C2(keyinput39), .A(n15211), .ZN(n15222) );
  AOI22_X1 U16762 ( .A1(n10938), .A2(keyinput60), .B1(n15213), .B2(keyinput27), 
        .ZN(n15212) );
  OAI221_X1 U16763 ( .B1(n10938), .B2(keyinput60), .C1(n15213), .C2(keyinput27), .A(n15212), .ZN(n15221) );
  AOI22_X1 U16764 ( .A1(n15333), .A2(keyinput55), .B1(n15215), .B2(keyinput37), 
        .ZN(n15214) );
  OAI221_X1 U16765 ( .B1(n15333), .B2(keyinput55), .C1(n15215), .C2(keyinput37), .A(n15214), .ZN(n15220) );
  XOR2_X1 U16766 ( .A(n15216), .B(keyinput54), .Z(n15218) );
  XNOR2_X1 U16767 ( .A(SI_0_), .B(keyinput26), .ZN(n15217) );
  NAND2_X1 U16768 ( .A1(n15218), .A2(n15217), .ZN(n15219) );
  NOR4_X1 U16769 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15251) );
  AOI22_X1 U16770 ( .A1(n15225), .A2(keyinput3), .B1(keyinput59), .B2(n15224), 
        .ZN(n15223) );
  OAI221_X1 U16771 ( .B1(n15225), .B2(keyinput3), .C1(n15224), .C2(keyinput59), 
        .A(n15223), .ZN(n15231) );
  AOI22_X1 U16772 ( .A1(n15228), .A2(keyinput45), .B1(n15227), .B2(keyinput40), 
        .ZN(n15226) );
  OAI221_X1 U16773 ( .B1(n15228), .B2(keyinput45), .C1(n15227), .C2(keyinput40), .A(n15226), .ZN(n15230) );
  XOR2_X1 U16774 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput47), .Z(n15229) );
  OR3_X1 U16775 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n15237) );
  AOI22_X1 U16776 ( .A1(n15233), .A2(keyinput35), .B1(n15343), .B2(keyinput12), 
        .ZN(n15232) );
  OAI221_X1 U16777 ( .B1(n15233), .B2(keyinput35), .C1(n15343), .C2(keyinput12), .A(n15232), .ZN(n15236) );
  XNOR2_X1 U16778 ( .A(n15234), .B(keyinput21), .ZN(n15235) );
  NOR3_X1 U16779 ( .A1(n15237), .A2(n15236), .A3(n15235), .ZN(n15250) );
  AOI22_X1 U16780 ( .A1(n15239), .A2(keyinput7), .B1(n15325), .B2(keyinput52), 
        .ZN(n15238) );
  OAI221_X1 U16781 ( .B1(n15239), .B2(keyinput7), .C1(n15325), .C2(keyinput52), 
        .A(n15238), .ZN(n15248) );
  INV_X1 U16782 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U16783 ( .A1(n15327), .A2(keyinput32), .B1(n15342), .B2(keyinput15), 
        .ZN(n15240) );
  OAI221_X1 U16784 ( .B1(n15327), .B2(keyinput32), .C1(n15342), .C2(keyinput15), .A(n15240), .ZN(n15247) );
  AOI22_X1 U16785 ( .A1(n15341), .A2(keyinput19), .B1(keyinput22), .B2(n15310), 
        .ZN(n15241) );
  OAI221_X1 U16786 ( .B1(n15341), .B2(keyinput19), .C1(n15310), .C2(keyinput22), .A(n15241), .ZN(n15246) );
  INV_X1 U16787 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15244) );
  INV_X1 U16788 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U16789 ( .A1(n15244), .A2(keyinput56), .B1(n15243), .B2(keyinput44), 
        .ZN(n15242) );
  OAI221_X1 U16790 ( .B1(n15244), .B2(keyinput56), .C1(n15243), .C2(keyinput44), .A(n15242), .ZN(n15245) );
  NOR4_X1 U16791 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        n15249) );
  NAND4_X1 U16792 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        n15306) );
  INV_X1 U16793 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n15254) );
  AOI22_X1 U16794 ( .A1(n15332), .A2(keyinput10), .B1(n15254), .B2(keyinput24), 
        .ZN(n15253) );
  OAI221_X1 U16795 ( .B1(n15332), .B2(keyinput10), .C1(n15254), .C2(keyinput24), .A(n15253), .ZN(n15264) );
  INV_X1 U16796 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U16797 ( .A1(n15313), .A2(keyinput31), .B1(keyinput16), .B2(n15256), 
        .ZN(n15255) );
  OAI221_X1 U16798 ( .B1(n15313), .B2(keyinput31), .C1(n15256), .C2(keyinput16), .A(n15255), .ZN(n15263) );
  AOI22_X1 U16799 ( .A1(n15258), .A2(keyinput9), .B1(keyinput4), .B2(n15314), 
        .ZN(n15257) );
  OAI221_X1 U16800 ( .B1(n15258), .B2(keyinput9), .C1(n15314), .C2(keyinput4), 
        .A(n15257), .ZN(n15262) );
  XNOR2_X1 U16801 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput33), .ZN(n15260)
         );
  XNOR2_X1 U16802 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput20), .ZN(n15259) );
  NAND2_X1 U16803 ( .A1(n15260), .A2(n15259), .ZN(n15261) );
  NOR4_X1 U16804 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15304) );
  INV_X1 U16805 ( .A(P1_WR_REG_SCAN_IN), .ZN(n15266) );
  AOI22_X1 U16806 ( .A1(n15266), .A2(keyinput49), .B1(n9344), .B2(keyinput34), 
        .ZN(n15265) );
  OAI221_X1 U16807 ( .B1(n15266), .B2(keyinput49), .C1(n9344), .C2(keyinput34), 
        .A(n15265), .ZN(n15275) );
  AOI22_X1 U16808 ( .A1(n15268), .A2(keyinput63), .B1(keyinput5), .B2(n15345), 
        .ZN(n15267) );
  OAI221_X1 U16809 ( .B1(n15268), .B2(keyinput63), .C1(n15345), .C2(keyinput5), 
        .A(n15267), .ZN(n15274) );
  XOR2_X1 U16810 ( .A(n9798), .B(keyinput0), .Z(n15272) );
  XNOR2_X1 U16811 ( .A(keyinput36), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n15271) );
  XNOR2_X1 U16812 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput50), .ZN(n15270) );
  XNOR2_X1 U16813 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput13), .ZN(n15269) );
  NAND4_X1 U16814 ( .A1(n15272), .A2(n15271), .A3(n15270), .A4(n15269), .ZN(
        n15273) );
  NOR3_X1 U16815 ( .A1(n15275), .A2(n15274), .A3(n15273), .ZN(n15303) );
  AOI22_X1 U16816 ( .A1(n11407), .A2(keyinput42), .B1(keyinput25), .B2(n9331), 
        .ZN(n15276) );
  OAI221_X1 U16817 ( .B1(n11407), .B2(keyinput42), .C1(n9331), .C2(keyinput25), 
        .A(n15276), .ZN(n15286) );
  AOI22_X1 U16818 ( .A1(n15344), .A2(keyinput62), .B1(keyinput29), .B2(n15278), 
        .ZN(n15277) );
  OAI221_X1 U16819 ( .B1(n15344), .B2(keyinput62), .C1(n15278), .C2(keyinput29), .A(n15277), .ZN(n15285) );
  AOI22_X1 U16820 ( .A1(n15280), .A2(keyinput17), .B1(keyinput30), .B2(n8542), 
        .ZN(n15279) );
  OAI221_X1 U16821 ( .B1(n15280), .B2(keyinput17), .C1(n8542), .C2(keyinput30), 
        .A(n15279), .ZN(n15284) );
  XNOR2_X1 U16822 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput8), .ZN(n15282) );
  XNOR2_X1 U16823 ( .A(SI_7_), .B(keyinput46), .ZN(n15281) );
  NAND2_X1 U16824 ( .A1(n15282), .A2(n15281), .ZN(n15283) );
  NOR4_X1 U16825 ( .A1(n15286), .A2(n15285), .A3(n15284), .A4(n15283), .ZN(
        n15302) );
  INV_X1 U16826 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n15288) );
  AOI22_X1 U16827 ( .A1(n15338), .A2(keyinput57), .B1(keyinput1), .B2(n15288), 
        .ZN(n15287) );
  OAI221_X1 U16828 ( .B1(n15338), .B2(keyinput57), .C1(n15288), .C2(keyinput1), 
        .A(n15287), .ZN(n15292) );
  XNOR2_X1 U16829 ( .A(n15324), .B(keyinput23), .ZN(n15291) );
  XNOR2_X1 U16830 ( .A(n15289), .B(keyinput11), .ZN(n15290) );
  OR3_X1 U16831 ( .A1(n15292), .A2(n15291), .A3(n15290), .ZN(n15300) );
  AOI22_X1 U16832 ( .A1(n15295), .A2(keyinput43), .B1(keyinput6), .B2(n15294), 
        .ZN(n15293) );
  OAI221_X1 U16833 ( .B1(n15295), .B2(keyinput43), .C1(n15294), .C2(keyinput6), 
        .A(n15293), .ZN(n15299) );
  AOI22_X1 U16834 ( .A1(n13469), .A2(keyinput51), .B1(keyinput2), .B2(n15297), 
        .ZN(n15296) );
  OAI221_X1 U16835 ( .B1(n13469), .B2(keyinput51), .C1(n15297), .C2(keyinput2), 
        .A(n15296), .ZN(n15298) );
  NOR3_X1 U16836 ( .A1(n15300), .A2(n15299), .A3(n15298), .ZN(n15301) );
  NAND4_X1 U16837 ( .A1(n15304), .A2(n15303), .A3(n15302), .A4(n15301), .ZN(
        n15305) );
  NOR2_X1 U16838 ( .A1(n15306), .A2(n15305), .ZN(n15309) );
  NAND2_X1 U16839 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n6405), .ZN(n15308) );
  XNOR2_X1 U16840 ( .A(n15309), .B(n15308), .ZN(n15354) );
  NOR4_X1 U16841 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_REG1_REG_26__SCAN_IN), .A4(P3_REG0_REG_2__SCAN_IN), .ZN(n15352) );
  NAND4_X1 U16842 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15316) );
  NAND4_X1 U16843 ( .A1(n9344), .A2(n9355), .A3(n9331), .A4(n15314), .ZN(
        n15315) );
  INV_X1 U16844 ( .A(SI_7_), .ZN(n15317) );
  AND3_X1 U16845 ( .A1(n15319), .A2(n15318), .A3(n15317), .ZN(n15351) );
  NAND4_X1 U16846 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(P2_REG0_REG_9__SCAN_IN), .A4(P1_IR_REG_27__SCAN_IN), .ZN(n15323)
         );
  NAND4_X1 U16847 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(P1_REG2_REG_8__SCAN_IN), 
        .A3(P3_ADDR_REG_14__SCAN_IN), .A4(P2_ADDR_REG_12__SCAN_IN), .ZN(n15322) );
  NAND4_X1 U16848 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), .A3(P2_REG0_REG_16__SCAN_IN), .A4(P1_REG0_REG_15__SCAN_IN), .ZN(n15321) );
  NAND4_X1 U16849 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P3_REG1_REG_18__SCAN_IN), .A3(P3_REG2_REG_31__SCAN_IN), .A4(P1_WR_REG_SCAN_IN), .ZN(n15320) );
  NOR4_X1 U16850 ( .A1(n15323), .A2(n15322), .A3(n15321), .A4(n15320), .ZN(
        n15350) );
  NOR4_X1 U16851 ( .A1(n15326), .A2(n15325), .A3(n15324), .A4(
        P1_IR_REG_25__SCAN_IN), .ZN(n15331) );
  INV_X1 U16852 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n15329) );
  NAND4_X1 U16853 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .A3(
        P1_IR_REG_10__SCAN_IN), .A4(n15327), .ZN(n15328) );
  NOR3_X1 U16854 ( .A1(n15329), .A2(n15278), .A3(n15328), .ZN(n15330) );
  NAND4_X1 U16855 ( .A1(n15331), .A2(P2_REG0_REG_22__SCAN_IN), .A3(
        P1_ADDR_REG_5__SCAN_IN), .A4(n15330), .ZN(n15334) );
  OR3_X1 U16856 ( .A1(n15334), .A2(n15333), .A3(n15332), .ZN(n15340) );
  NOR4_X1 U16857 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_DATAO_REG_11__SCAN_IN), 
        .A3(P3_DATAO_REG_1__SCAN_IN), .A4(P3_DATAO_REG_31__SCAN_IN), .ZN(
        n15335) );
  NAND4_X1 U16858 ( .A1(n15336), .A2(P3_ADDR_REG_2__SCAN_IN), .A3(
        P3_ADDR_REG_1__SCAN_IN), .A4(n15335), .ZN(n15339) );
  NOR4_X1 U16859 ( .A1(n15340), .A2(n15339), .A3(n15338), .A4(n15337), .ZN(
        n15348) );
  NOR4_X1 U16860 ( .A1(n15344), .A2(n15343), .A3(n15342), .A4(n15341), .ZN(
        n15347) );
  NOR4_X1 U16861 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(P3_REG2_REG_14__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(n15345), .ZN(n15346) );
  AND3_X1 U16862 ( .A1(n15348), .A2(n15347), .A3(n15346), .ZN(n15349) );
  NAND4_X1 U16863 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15353) );
  XNOR2_X1 U16864 ( .A(n15354), .B(n15353), .ZN(P1_U3317) );
  AOI21_X1 U16865 ( .B1(n15357), .B2(n15356), .A(n15355), .ZN(SUB_1596_U59) );
  OAI21_X1 U16866 ( .B1(n15360), .B2(n15359), .A(n15358), .ZN(SUB_1596_U58) );
  XNOR2_X1 U16867 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15361), .ZN(SUB_1596_U53)
         );
  AOI21_X1 U16868 ( .B1(n15364), .B2(n15363), .A(n15362), .ZN(SUB_1596_U56) );
  AOI21_X1 U16869 ( .B1(n15367), .B2(n15366), .A(n15365), .ZN(n15368) );
  XOR2_X1 U16870 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15368), .Z(SUB_1596_U60) );
  AOI21_X1 U16871 ( .B1(n15371), .B2(n15370), .A(n15369), .ZN(SUB_1596_U5) );
  BUF_X1 U7275 ( .A(n8371), .Z(n8455) );
  OR2_X2 U7239 ( .A1(n12331), .A2(n8101), .ZN(n12483) );
  INV_X2 U7161 ( .A(n12483), .ZN(n12487) );
  NAND2_X1 U9571 ( .A1(n7304), .A2(n7306), .ZN(n14030) );
  NAND2_X1 U7442 ( .A1(n7561), .A2(n7560), .ZN(n7591) );
  CLKBUF_X2 U7166 ( .A(n9811), .Z(n6416) );
  CLKBUF_X1 U7170 ( .A(n7657), .Z(n8216) );
  CLKBUF_X1 U7179 ( .A(n9093), .Z(n6427) );
  NAND2_X1 U7188 ( .A1(n14317), .A2(n14653), .ZN(n11715) );
  CLKBUF_X1 U7213 ( .A(n9944), .Z(n11797) );
  NAND2_X1 U7215 ( .A1(n6966), .A2(n13944), .ZN(n14129) );
  INV_X1 U7225 ( .A(n14705), .ZN(n6990) );
  NAND2_X1 U7228 ( .A1(n9607), .A2(n9608), .ZN(n11542) );
  NAND2_X1 U7477 ( .A1(n8303), .A2(n13676), .ZN(n8411) );
  AND2_X1 U8838 ( .A1(n9580), .A2(n9261), .ZN(n15375) );
endmodule

