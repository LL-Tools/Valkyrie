

module b15_C_gen_AntiSAT_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785;

  INV_X2 U3434 ( .A(n3512), .ZN(n5857) );
  BUF_X2 U3435 ( .A(n3857), .Z(n2988) );
  CLKBUF_X1 U3436 ( .A(n3273), .Z(n4245) );
  CLKBUF_X2 U3437 ( .A(n3138), .Z(n3002) );
  CLKBUF_X2 U3438 ( .A(n3211), .Z(n4128) );
  CLKBUF_X2 U3439 ( .A(n3210), .Z(n4244) );
  CLKBUF_X2 U3440 ( .A(n3219), .Z(n4337) );
  NAND2_X1 U3441 ( .A1(n3614), .A2(n4343), .ZN(n3297) );
  CLKBUF_X2 U3442 ( .A(n3272), .Z(n2991) );
  INV_X1 U3443 ( .A(n3227), .ZN(n3240) );
  AND2_X2 U3444 ( .A1(n5762), .A2(n4408), .ZN(n3353) );
  AND2_X1 U34450 ( .A1(n3117), .A2(n5762), .ZN(n3398) );
  AND2_X1 U34460 ( .A1(n4409), .A2(n4503), .ZN(n3210) );
  AND2_X1 U34470 ( .A1(n3117), .A2(n3119), .ZN(n3138) );
  INV_X1 U3449 ( .A(n6785), .ZN(n2987) );
  AND2_X2 U34510 ( .A1(n4503), .A2(n4408), .ZN(n4243) );
  AND2_X1 U34520 ( .A1(n4337), .A2(n3236), .ZN(n3549) );
  AND2_X1 U34530 ( .A1(n3244), .A2(n3236), .ZN(n3638) );
  INV_X1 U3454 ( .A(n6032), .ZN(n6029) );
  XNOR2_X1 U34560 ( .A(n3322), .B(n3372), .ZN(n3857) );
  OAI22_X2 U3458 ( .A1(n5575), .A2(n5557), .B1(n5564), .B2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5558) );
  NAND2_X2 U34590 ( .A1(n3178), .A2(n3109), .ZN(n4343) );
  AND2_X2 U34600 ( .A1(n4503), .A2(n4408), .ZN(n2989) );
  AND2_X2 U34610 ( .A1(n5762), .A2(n4408), .ZN(n2990) );
  AND2_X2 U34620 ( .A1(n4069), .A2(n3020), .ZN(n5452) );
  OAI222_X1 U34630 ( .A1(n3873), .A2(n6328), .B1(n6322), .B2(n5756), .C1(n6371), .C2(n5755), .ZN(n5757) );
  NAND2_X1 U34640 ( .A1(n4480), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U34650 ( .A1(n3746), .A2(n3624), .ZN(n6201) );
  NAND2_X1 U3466 ( .A1(n5489), .A2(n4444), .ZN(n5843) );
  NAND2_X1 U3467 ( .A1(n3052), .A2(n3050), .ZN(n3332) );
  XNOR2_X1 U34680 ( .A(n3341), .B(n3320), .ZN(n4318) );
  NAND2_X2 U34690 ( .A1(n3251), .A2(n3250), .ZN(n3341) );
  CLKBUF_X1 U34700 ( .A(n3343), .Z(n2994) );
  AND3_X1 U34710 ( .A1(n3244), .A2(n3240), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3577) );
  NAND2_X2 U34720 ( .A1(n3202), .A2(n3201), .ZN(n3236) );
  BUF_X2 U34730 ( .A(n3179), .Z(n4238) );
  AND2_X2 U34740 ( .A1(n6441), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5762) );
  AND2_X1 U3475 ( .A1(n3111), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3119)
         );
  INV_X1 U3476 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6441) );
  AND2_X1 U3477 ( .A1(n3767), .A2(n3031), .ZN(n3030) );
  OR2_X1 U3478 ( .A1(n4309), .A2(n6201), .ZN(n3767) );
  OR2_X1 U3479 ( .A1(n4309), .A2(n6124), .ZN(n4310) );
  AND2_X1 U3480 ( .A1(n3013), .A2(n4235), .ZN(n3076) );
  NOR2_X1 U3481 ( .A1(n5528), .A2(n5641), .ZN(n5508) );
  CLKBUF_X1 U3482 ( .A(n5420), .Z(n5421) );
  NAND2_X1 U3483 ( .A1(n5162), .A2(n5163), .ZN(n6105) );
  NAND2_X2 U3484 ( .A1(n5172), .A2(n4005), .ZN(n5230) );
  OR2_X1 U3485 ( .A1(n3992), .A2(n3991), .ZN(n4005) );
  NAND2_X1 U3486 ( .A1(n4713), .A2(n3490), .ZN(n4878) );
  NAND2_X1 U3487 ( .A1(n4526), .A2(n3438), .ZN(n4542) );
  INV_X1 U3488 ( .A(n4924), .ZN(n4925) );
  NOR2_X1 U3489 ( .A1(n4672), .A2(n3091), .ZN(n4924) );
  NAND2_X1 U3490 ( .A1(n4524), .A2(n4523), .ZN(n4526) );
  OR2_X1 U3491 ( .A1(n4544), .A2(n3049), .ZN(n3048) );
  XNOR2_X1 U3492 ( .A(n3511), .B(n6177), .ZN(n4966) );
  XNOR2_X1 U3493 ( .A(n3494), .B(n3493), .ZN(n3891) );
  NAND2_X1 U3494 ( .A1(n3340), .A2(n3339), .ZN(n6130) );
  NAND2_X1 U3495 ( .A1(n3479), .A2(n3478), .ZN(n3494) );
  NAND2_X1 U3496 ( .A1(n3411), .A2(n4313), .ZN(n3412) );
  NOR2_X1 U3497 ( .A1(n6069), .A2(n6571), .ZN(n6099) );
  NOR2_X1 U3498 ( .A1(n4634), .A2(n5188), .ZN(n6408) );
  NOR2_X1 U3499 ( .A1(n6719), .A2(n5188), .ZN(n6402) );
  NOR2_X1 U3500 ( .A1(n6738), .A2(n5188), .ZN(n6396) );
  NOR2_X1 U3501 ( .A1(n6683), .A2(n5188), .ZN(n6390) );
  AND2_X1 U3502 ( .A1(n3374), .A2(n3373), .ZN(n3407) );
  CLKBUF_X1 U3503 ( .A(n4351), .Z(n4760) );
  OR2_X1 U3504 ( .A1(n5485), .A2(n5410), .ZN(n5473) );
  NAND2_X1 U3505 ( .A1(n3332), .A2(n3331), .ZN(n4314) );
  NAND2_X1 U3506 ( .A1(n3332), .A2(n3284), .ZN(n3370) );
  OR2_X2 U3507 ( .A1(n4737), .A2(n4385), .ZN(n4446) );
  OAI21_X2 U3508 ( .B1(n4318), .B2(STATE2_REG_0__SCAN_IN), .A(n3321), .ZN(
        n3372) );
  NAND2_X1 U3509 ( .A1(n3344), .A2(n2994), .ZN(n3382) );
  AND2_X1 U3510 ( .A1(n3343), .A2(n3319), .ZN(n3342) );
  OR2_X1 U3511 ( .A1(n3247), .A2(n3503), .ZN(n3741) );
  NAND3_X1 U3512 ( .A1(n3191), .A2(n3239), .A3(n3304), .ZN(n3303) );
  NAND2_X1 U3513 ( .A1(n3169), .A2(n3219), .ZN(n3228) );
  OR2_X1 U3514 ( .A1(n3265), .A2(n3264), .ZN(n3504) );
  NAND2_X1 U3515 ( .A1(n3169), .A2(n3227), .ZN(n3077) );
  INV_X2 U3516 ( .A(n3244), .ZN(n3307) );
  AND4_X2 U3517 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3227)
         );
  INV_X2 U3518 ( .A(n3236), .ZN(n3612) );
  OR2_X2 U3519 ( .A1(n3217), .A2(n3216), .ZN(n3244) );
  AND3_X1 U3520 ( .A1(n3162), .A2(n3161), .A3(n3160), .ZN(n3167) );
  AND4_X1 U3521 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3201)
         );
  AND4_X1 U3522 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3152)
         );
  AND4_X1 U3523 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3154)
         );
  AND4_X1 U3524 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3178)
         );
  AND4_X1 U3525 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3155)
         );
  AND4_X1 U3526 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3124)
         );
  AND4_X1 U3527 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3202)
         );
  AND4_X1 U3528 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3125)
         );
  BUF_X2 U3529 ( .A(n3398), .Z(n3258) );
  CLKBUF_X1 U3530 ( .A(n3204), .Z(n4109) );
  BUF_X2 U3531 ( .A(n3259), .Z(n3267) );
  AND2_X2 U3532 ( .A1(n3117), .A2(n4503), .ZN(n3393) );
  AND2_X2 U3533 ( .A1(n3119), .A2(n4408), .ZN(n3157) );
  AND2_X2 U3534 ( .A1(n3047), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3117)
         );
  CLKBUF_X1 U3535 ( .A(n6441), .Z(n2996) );
  AND2_X2 U3536 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4503) );
  NOR2_X2 U3537 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5760) );
  INV_X1 U3538 ( .A(n3169), .ZN(n2992) );
  NAND2_X1 U3539 ( .A1(n3597), .A2(n3612), .ZN(n2993) );
  OR2_X2 U3540 ( .A1(n2997), .A2(n2998), .ZN(n3241) );
  NAND2_X1 U3541 ( .A1(n3597), .A2(n3612), .ZN(n3622) );
  NOR2_X2 U3542 ( .A1(n3303), .A2(n3302), .ZN(n3597) );
  NAND2_X2 U3543 ( .A1(n3252), .A2(n3341), .ZN(n3862) );
  OAI211_X1 U3544 ( .C1(n3314), .C2(n3112), .A(n3315), .B(n3316), .ZN(n3343)
         );
  AND2_X2 U3545 ( .A1(n3118), .A2(n5760), .ZN(n3003) );
  CLKBUF_X1 U3546 ( .A(n4526), .Z(n2995) );
  INV_X2 U3547 ( .A(n3241), .ZN(n3169) );
  NOR2_X1 U3548 ( .A1(n3234), .A2(n3297), .ZN(n3593) );
  NAND2_X2 U3549 ( .A1(n3167), .A2(n3015), .ZN(n3192) );
  NAND4_X1 U3550 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n2997)
         );
  NAND4_X1 U3551 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n2998)
         );
  AND2_X2 U3553 ( .A1(n3611), .A2(n3244), .ZN(n4280) );
  AND2_X2 U3554 ( .A1(n3323), .A2(n3299), .ZN(n3611) );
  AND2_X1 U3555 ( .A1(n3117), .A2(n4503), .ZN(n3000) );
  AND2_X2 U3556 ( .A1(n3117), .A2(n4503), .ZN(n3001) );
  AND2_X4 U3557 ( .A1(n5760), .A2(n4409), .ZN(n3180) );
  NOR2_X4 U3558 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4409) );
  NAND2_X2 U3559 ( .A1(n5553), .A2(n5552), .ZN(n5563) );
  NOR2_X1 U3560 ( .A1(n3460), .A2(n3439), .ZN(n3452) );
  NAND2_X2 U3561 ( .A1(n3406), .A2(n3405), .ZN(n3410) );
  NAND2_X2 U3562 ( .A1(n4878), .A2(n4880), .ZN(n4879) );
  NAND2_X2 U3563 ( .A1(n3412), .A2(n3460), .ZN(n3873) );
  OAI21_X2 U3564 ( .B1(n6105), .B2(n3014), .A(n3517), .ZN(n5236) );
  AND2_X1 U3565 ( .A1(n3119), .A2(n4409), .ZN(n3272) );
  AND2_X4 U3566 ( .A1(n3118), .A2(n5760), .ZN(n3004) );
  AND2_X1 U3567 ( .A1(n3118), .A2(n5760), .ZN(n3838) );
  OR2_X1 U3568 ( .A1(n3217), .A2(n3216), .ZN(n3005) );
  OR2_X1 U3569 ( .A1(n3217), .A2(n3216), .ZN(n3006) );
  AND2_X4 U3570 ( .A1(n3118), .A2(n4503), .ZN(n3204) );
  OAI21_X1 U3571 ( .B1(n3303), .B2(n3218), .A(n3307), .ZN(n3247) );
  OAI21_X1 U3572 ( .B1(n3556), .B2(n3169), .A(n3192), .ZN(n3203) );
  OR2_X1 U3573 ( .A1(n3244), .A2(n6466), .ZN(n3392) );
  AOI21_X1 U3574 ( .B1(n6446), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3546), 
        .ZN(n3582) );
  INV_X1 U3575 ( .A(n4203), .ZN(n4258) );
  NOR2_X1 U3576 ( .A1(n5296), .A2(n6466), .ZN(n4203) );
  NAND2_X1 U3577 ( .A1(n3092), .A2(n4926), .ZN(n3091) );
  INV_X1 U3578 ( .A(n3094), .ZN(n3092) );
  INV_X1 U3579 ( .A(n4673), .ZN(n3925) );
  INV_X1 U3580 ( .A(n3892), .ZN(n4261) );
  NAND2_X1 U3581 ( .A1(n6374), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3988) );
  CLKBUF_X1 U3582 ( .A(n3892), .Z(n4208) );
  NOR2_X2 U3583 ( .A1(n2992), .A2(n6374), .ZN(n4018) );
  OR2_X1 U3584 ( .A1(n3240), .A2(n6466), .ZN(n3391) );
  NAND2_X1 U3585 ( .A1(n4367), .A2(n4283), .ZN(n5269) );
  INV_X1 U3586 ( .A(n6477), .ZN(n4431) );
  INV_X1 U3587 ( .A(n3988), .ZN(n4277) );
  INV_X1 U3588 ( .A(n3638), .ZN(n4368) );
  INV_X1 U3589 ( .A(n2988), .ZN(n4511) );
  OR2_X1 U3590 ( .A1(n3619), .A2(n3556), .ZN(n6455) );
  AND2_X1 U3591 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  AND2_X1 U3592 ( .A1(n3451), .A2(n3450), .ZN(n3461) );
  NAND2_X1 U3593 ( .A1(n3431), .A2(n3430), .ZN(n3463) );
  NAND2_X1 U3594 ( .A1(n3522), .A2(n3016), .ZN(n3059) );
  OR2_X1 U3595 ( .A1(n3228), .A2(n3240), .ZN(n3230) );
  NOR2_X1 U3596 ( .A1(n3101), .A2(n3099), .ZN(n3098) );
  INV_X1 U3597 ( .A(n5361), .ZN(n3101) );
  NAND2_X1 U3598 ( .A1(n3100), .A2(n4191), .ZN(n3099) );
  INV_X1 U3599 ( .A(n5375), .ZN(n3100) );
  INV_X1 U3600 ( .A(n5422), .ZN(n4191) );
  OR2_X1 U3601 ( .A1(n5446), .A2(n5439), .ZN(n3104) );
  INV_X1 U3602 ( .A(n5459), .ZN(n3082) );
  AND2_X1 U3603 ( .A1(n4091), .A2(n4068), .ZN(n3083) );
  INV_X1 U3604 ( .A(n5470), .ZN(n4091) );
  NAND2_X1 U3605 ( .A1(n4424), .A2(n4425), .ZN(n3078) );
  NAND2_X1 U3606 ( .A1(n3045), .A2(n5377), .ZN(n3044) );
  INV_X1 U3607 ( .A(n5430), .ZN(n3045) );
  NAND2_X1 U3608 ( .A1(n5447), .A2(n3042), .ZN(n3041) );
  INV_X1 U3609 ( .A(n5464), .ZN(n3042) );
  NAND2_X1 U3610 ( .A1(n3053), .A2(n3008), .ZN(n5549) );
  INV_X1 U3611 ( .A(n4709), .ZN(n3659) );
  NOR2_X1 U3612 ( .A1(n3034), .A2(n4517), .ZN(n3033) );
  INV_X1 U3613 ( .A(n4552), .ZN(n3034) );
  AND2_X1 U3614 ( .A1(n5461), .A2(n3638), .ZN(n3695) );
  INV_X1 U3615 ( .A(n3695), .ZN(n3727) );
  AND2_X1 U3616 ( .A1(n5771), .A2(n3245), .ZN(n3070) );
  OR2_X1 U3617 ( .A1(n3279), .A2(n3278), .ZN(n3376) );
  OR2_X1 U3618 ( .A1(n3363), .A2(n3362), .ZN(n3413) );
  NAND2_X1 U3619 ( .A1(n3168), .A2(n3614), .ZN(n3191) );
  OR2_X1 U3620 ( .A1(n4317), .A2(n4561), .ZN(n6321) );
  NAND2_X1 U3621 ( .A1(n5269), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4827) );
  AND2_X1 U3622 ( .A1(n4127), .A2(n4126), .ZN(n5453) );
  NAND2_X1 U3623 ( .A1(n4211), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4237)
         );
  AND2_X1 U3624 ( .A1(n5571), .A2(n3892), .ZN(n4170) );
  AND2_X1 U3625 ( .A1(n3982), .A2(n3981), .ZN(n5048) );
  AND4_X1 U3626 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n4673)
         );
  NAND2_X1 U3627 ( .A1(n3895), .A2(n3894), .ZN(n4707) );
  INV_X1 U3628 ( .A(n4516), .ZN(n3889) );
  INV_X1 U3629 ( .A(n3870), .ZN(n3875) );
  NAND2_X1 U3630 ( .A1(n3875), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3874)
         );
  OAI211_X1 U3631 ( .C1(n3878), .C2(n2996), .A(n3872), .B(n3871), .ZN(n4482)
         );
  INV_X1 U3632 ( .A(n3626), .ZN(n5461) );
  NOR3_X1 U3633 ( .A1(n5431), .A2(n3046), .A3(n5430), .ZN(n5426) );
  OR2_X1 U3634 ( .A1(n3018), .A2(n5390), .ZN(n5431) );
  NAND2_X1 U3635 ( .A1(n5901), .A2(n3010), .ZN(n5485) );
  NOR2_X1 U3636 ( .A1(n3523), .A2(n3061), .ZN(n3060) );
  AND2_X1 U3637 ( .A1(n3512), .A2(n5613), .ZN(n3523) );
  INV_X1 U3638 ( .A(n3520), .ZN(n3061) );
  NOR2_X1 U3639 ( .A1(n5980), .A2(n5050), .ZN(n5901) );
  NOR2_X1 U3640 ( .A1(n3744), .A2(n3743), .ZN(n5315) );
  NAND2_X1 U3641 ( .A1(n3618), .A2(n3617), .ZN(n3746) );
  OR2_X1 U3642 ( .A1(n4737), .A2(n3616), .ZN(n3617) );
  AND2_X1 U3643 ( .A1(n4842), .A2(n4315), .ZN(n6369) );
  INV_X1 U3644 ( .A(n4562), .ZN(n6370) );
  CLKBUF_X1 U3645 ( .A(n3855), .Z(n4312) );
  NAND2_X1 U3646 ( .A1(n3588), .A2(n3587), .ZN(n5314) );
  NAND2_X1 U3647 ( .A1(n3600), .A2(n3586), .ZN(n3587) );
  NAND2_X1 U3648 ( .A1(n3585), .A2(n3584), .ZN(n3588) );
  AND2_X1 U3649 ( .A1(n5269), .A2(n4286), .ZN(n6026) );
  AND2_X1 U3650 ( .A1(n5489), .A2(n4274), .ZN(n6066) );
  INV_X1 U3651 ( .A(n5489), .ZN(n6065) );
  AND2_X1 U3652 ( .A1(n5489), .A2(n4445), .ZN(n5279) );
  NAND2_X1 U3653 ( .A1(n4222), .A2(n4262), .ZN(n5302) );
  OR2_X1 U3654 ( .A1(n4220), .A2(n4221), .ZN(n4222) );
  INV_X1 U3655 ( .A(n6139), .ZN(n6109) );
  NAND2_X1 U3656 ( .A1(n6124), .A2(n4230), .ZN(n5616) );
  OR2_X1 U3657 ( .A1(n3073), .A2(n3534), .ZN(n3105) );
  XNOR2_X1 U3658 ( .A(n3731), .B(n3730), .ZN(n5414) );
  XNOR2_X1 U3659 ( .A(n4228), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5638)
         );
  XNOR2_X1 U3660 ( .A(n3370), .B(n3371), .ZN(n3322) );
  INV_X1 U3661 ( .A(n4315), .ZN(n6322) );
  AND2_X1 U3662 ( .A1(n3313), .A2(n3312), .ZN(n3316) );
  AND2_X1 U3663 ( .A1(n3477), .A2(n3476), .ZN(n3481) );
  OR2_X1 U3664 ( .A1(n3449), .A2(n3448), .ZN(n3482) );
  OR2_X1 U3665 ( .A1(n3429), .A2(n3428), .ZN(n3483) );
  AND2_X2 U3666 ( .A1(n3112), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3118)
         );
  OR2_X1 U3667 ( .A1(n3404), .A2(n3403), .ZN(n3432) );
  NAND2_X1 U3668 ( .A1(n3577), .A2(n3549), .ZN(n3578) );
  OR2_X1 U3669 ( .A1(n3548), .A2(n3547), .ZN(n3579) );
  NAND2_X1 U3670 ( .A1(n5230), .A2(n3086), .ZN(n5397) );
  NOR2_X1 U3671 ( .A1(n3090), .A2(n3087), .ZN(n3086) );
  INV_X1 U3672 ( .A(n5482), .ZN(n3090) );
  INV_X1 U3673 ( .A(n3088), .ZN(n3087) );
  NOR2_X1 U3674 ( .A1(n5259), .A2(n3089), .ZN(n3088) );
  INV_X1 U3675 ( .A(n5232), .ZN(n3089) );
  AOI21_X1 U3676 ( .B1(n3863), .B2(EAX_REG_13__SCAN_IN), .A(n3990), .ZN(n3991)
         );
  NAND2_X1 U3677 ( .A1(n3095), .A2(n3925), .ZN(n3094) );
  INV_X1 U3678 ( .A(n4756), .ZN(n3095) );
  INV_X1 U3679 ( .A(n5261), .ZN(n3039) );
  INV_X1 U3680 ( .A(n3058), .ZN(n3057) );
  OAI21_X1 U3681 ( .B1(n3059), .B2(n3060), .A(n3524), .ZN(n3058) );
  NAND2_X1 U3682 ( .A1(n3055), .A2(n3054), .ZN(n3053) );
  INV_X1 U3683 ( .A(n3059), .ZN(n3054) );
  NOR2_X1 U3684 ( .A1(n3011), .A2(n3068), .ZN(n3067) );
  NOR2_X1 U3685 ( .A1(n3663), .A2(n4710), .ZN(n3038) );
  NOR2_X1 U3686 ( .A1(n3147), .A2(n3146), .ZN(n3153) );
  AND2_X1 U3687 ( .A1(n2989), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U3688 ( .A1(n3638), .A2(n5454), .ZN(n3723) );
  NAND2_X1 U3689 ( .A1(n3304), .A2(n3240), .ZN(n3589) );
  INV_X1 U3690 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U3691 ( .A1(n3138), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3188) );
  AOI21_X1 U3692 ( .B1(n2990), .B2(INSTQUEUE_REG_11__0__SCAN_IN), .A(n3209), 
        .ZN(n3215) );
  AND2_X1 U3693 ( .A1(n3004), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U3694 ( .A1(n3179), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U3695 ( .A1(n3211), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3162) );
  AOI21_X1 U3696 ( .B1(n6483), .B2(n4741), .A(n6470), .ZN(n4324) );
  NAND2_X1 U3697 ( .A1(n3392), .A2(n3391), .ZN(n3586) );
  INV_X1 U3698 ( .A(n3578), .ZN(n3583) );
  NOR2_X1 U3699 ( .A1(n6533), .A2(n5404), .ZN(n5935) );
  INV_X1 U3700 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U3701 ( .A1(n5901), .A2(n3019), .ZN(n5262) );
  AND2_X1 U3702 ( .A1(n5901), .A2(n5900), .ZN(n5903) );
  AND2_X1 U3703 ( .A1(n4740), .A2(n4739), .ZN(n6069) );
  NAND2_X1 U3704 ( .A1(n4446), .A2(n4738), .ZN(n4740) );
  OR2_X1 U3705 ( .A1(n4237), .A2(n4236), .ZN(n4284) );
  AOI22_X1 U3706 ( .A1(n3854), .A2(n3853), .B1(n3892), .B2(n5339), .ZN(n4220)
         );
  AND2_X1 U3707 ( .A1(n3852), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4211)
         );
  INV_X1 U3708 ( .A(n5348), .ZN(n3096) );
  AOI22_X1 U3709 ( .A1(n4210), .A2(n4209), .B1(n4208), .B2(n5534), .ZN(n5361)
         );
  AND2_X1 U3710 ( .A1(n4188), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4193)
         );
  INV_X1 U3711 ( .A(n3099), .ZN(n3097) );
  NAND2_X1 U3712 ( .A1(n3103), .A2(n5387), .ZN(n3102) );
  INV_X1 U3713 ( .A(n3104), .ZN(n3103) );
  AND2_X1 U3714 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3851), .ZN(n4162)
         );
  NAND2_X1 U3715 ( .A1(n4162), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4169)
         );
  AND2_X1 U3716 ( .A1(n4106), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4125)
         );
  NOR2_X1 U3717 ( .A1(n4050), .A2(n5405), .ZN(n4084) );
  OR2_X1 U3718 ( .A1(n5942), .A2(n4261), .ZN(n4089) );
  NAND2_X1 U3719 ( .A1(n4037), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4050)
         );
  CLKBUF_X1 U3720 ( .A(n5397), .Z(n5398) );
  NOR2_X1 U3721 ( .A1(n4021), .A2(n5271), .ZN(n4037) );
  INV_X1 U3722 ( .A(n3985), .ZN(n4006) );
  AND2_X1 U3723 ( .A1(n3968), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3986)
         );
  NAND2_X1 U3724 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3985)
         );
  NAND2_X1 U3725 ( .A1(n3941), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3954)
         );
  INV_X1 U3726 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5983) );
  NOR2_X1 U3727 ( .A1(n3926), .A2(n6006), .ZN(n3941) );
  AND2_X1 U3728 ( .A1(n3902), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3920)
         );
  INV_X1 U3729 ( .A(n4672), .ZN(n3093) );
  NAND2_X1 U3730 ( .A1(n3896), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3901)
         );
  INV_X1 U3731 ( .A(n3874), .ZN(n3883) );
  OAI21_X1 U3732 ( .B1(n3873), .B2(n4035), .A(n3880), .ZN(n4489) );
  NAND2_X1 U3733 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3870) );
  NAND2_X1 U3734 ( .A1(n3856), .A2(n3988), .ZN(n3081) );
  NOR2_X1 U3735 ( .A1(n5351), .A2(n5307), .ZN(n5326) );
  NAND2_X1 U3736 ( .A1(n5364), .A2(n5349), .ZN(n5351) );
  NOR3_X1 U3737 ( .A1(n5431), .A2(n3044), .A3(n3043), .ZN(n5364) );
  OR2_X1 U3738 ( .A1(n3046), .A2(n5362), .ZN(n3043) );
  AND2_X1 U3739 ( .A1(n3075), .A2(n3530), .ZN(n3074) );
  INV_X1 U3740 ( .A(n5543), .ZN(n3075) );
  AND2_X1 U3741 ( .A1(n3715), .A2(n3714), .ZN(n5430) );
  NOR2_X1 U3742 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  OR2_X1 U3743 ( .A1(n3041), .A2(n5440), .ZN(n3040) );
  AND2_X1 U3745 ( .A1(n3677), .A2(n3676), .ZN(n5050) );
  OR2_X1 U3746 ( .A1(n5976), .A2(n3674), .ZN(n5980) );
  NAND2_X1 U3747 ( .A1(n3659), .A2(n3035), .ZN(n5976) );
  NOR2_X1 U3748 ( .A1(n3037), .A2(n3036), .ZN(n3035) );
  INV_X1 U3749 ( .A(n4809), .ZN(n3036) );
  INV_X1 U3750 ( .A(n3038), .ZN(n3037) );
  INV_X1 U3751 ( .A(n3502), .ZN(n3068) );
  AND2_X1 U3752 ( .A1(n3659), .A2(n3038), .ZN(n4810) );
  NAND2_X1 U3753 ( .A1(n3032), .A2(n3007), .ZN(n4709) );
  NAND2_X1 U3754 ( .A1(n3032), .A2(n3033), .ZN(n4663) );
  NOR2_X1 U3755 ( .A1(n4518), .A2(n4517), .ZN(n4553) );
  NOR2_X1 U3756 ( .A1(n4548), .A2(n6227), .ZN(n4545) );
  AND2_X1 U3757 ( .A1(n5743), .A2(n5906), .ZN(n4548) );
  NAND2_X1 U3758 ( .A1(n3857), .A2(n3549), .ZN(n3327) );
  NAND2_X1 U3759 ( .A1(n3639), .A2(n5454), .ZN(n4418) );
  AND2_X1 U3760 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3084) );
  AND3_X1 U3761 ( .A1(n3072), .A2(n3246), .A3(n3070), .ZN(n3069) );
  AND2_X1 U3762 ( .A1(n3051), .A2(n3329), .ZN(n3050) );
  OAI211_X1 U3763 ( .C1(n3504), .C2(n3391), .A(n3296), .B(n3295), .ZN(n3371)
         );
  NAND2_X1 U3764 ( .A1(n3366), .A2(n3365), .ZN(n3369) );
  NAND2_X1 U3765 ( .A1(n3364), .A2(n3413), .ZN(n3365) );
  OR2_X1 U3766 ( .A1(n3228), .A2(n3589), .ZN(n5296) );
  CLKBUF_X1 U3767 ( .A(n3157), .Z(n5764) );
  NAND2_X1 U3768 ( .A1(n3384), .A2(n3383), .ZN(n4379) );
  INV_X1 U3769 ( .A(n6439), .ZN(n6443) );
  AND2_X1 U3770 ( .A1(n4350), .A2(n6237), .ZN(n4559) );
  NOR2_X1 U3771 ( .A1(n6366), .A2(n2988), .ZN(n4677) );
  AND2_X1 U3772 ( .A1(n2988), .A2(n4314), .ZN(n4840) );
  NOR2_X1 U3773 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4324), .ZN(n4765) );
  AND2_X1 U3774 ( .A1(n4312), .A2(n4533), .ZN(n4538) );
  AOI22_X1 U3775 ( .A1(n3398), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3132) );
  NOR2_X1 U3776 ( .A1(n6558), .A2(n4324), .ZN(n4574) );
  INV_X1 U3777 ( .A(n6569), .ZN(n4367) );
  NAND2_X1 U3778 ( .A1(n4386), .A2(n4364), .ZN(n6569) );
  INV_X1 U3779 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6758) );
  INV_X1 U3780 ( .A(n6026), .ZN(n6009) );
  INV_X1 U3781 ( .A(n6031), .ZN(n6005) );
  OR2_X1 U3782 ( .A1(n4827), .A2(n4290), .ZN(n5267) );
  INV_X1 U3783 ( .A(n6016), .ZN(n6034) );
  OR2_X1 U3784 ( .A1(n4821), .A2(n6026), .ZN(n5070) );
  INV_X1 U3785 ( .A(n5469), .ZN(n6052) );
  AND2_X1 U3786 ( .A1(n6055), .A2(n5488), .ZN(n6051) );
  AND2_X2 U3787 ( .A1(n4432), .A2(n4431), .ZN(n6055) );
  INV_X1 U3788 ( .A(n6051), .ZN(n6045) );
  INV_X1 U3789 ( .A(n6052), .ZN(n5487) );
  INV_X1 U3790 ( .A(n5843), .ZN(n6063) );
  NAND2_X1 U3791 ( .A1(n4271), .A2(n4478), .ZN(n5489) );
  INV_X1 U3792 ( .A(n5279), .ZN(n4668) );
  INV_X2 U3795 ( .A(n4476), .ZN(n4473) );
  OR2_X1 U3796 ( .A1(n4737), .A2(n4270), .ZN(n4478) );
  OR2_X1 U3797 ( .A1(n4269), .A2(READY_N), .ZN(n4270) );
  AOI21_X1 U3798 ( .B1(n6573), .B2(READY_N), .A(n4386), .ZN(n4476) );
  XNOR2_X1 U3799 ( .A(n4285), .B(n4296), .ZN(n4831) );
  OR2_X1 U3800 ( .A1(n4284), .A2(n5331), .ZN(n4285) );
  INV_X1 U3801 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5567) );
  CLKBUF_X1 U3802 ( .A(n4991), .Z(n4992) );
  INV_X1 U3803 ( .A(n5616), .ZN(n6129) );
  INV_X2 U3804 ( .A(n6122), .ZN(n6133) );
  OR2_X1 U3805 ( .A1(n5701), .A2(n3761), .ZN(n5686) );
  NOR3_X1 U3806 ( .A1(n5473), .A2(n3706), .A3(n5464), .ZN(n5448) );
  AND2_X1 U3807 ( .A1(n5475), .A2(n5474), .ZN(n5939) );
  NAND2_X1 U3808 ( .A1(n3521), .A2(n3060), .ZN(n3056) );
  NAND2_X1 U3809 ( .A1(n4879), .A2(n3502), .ZN(n4967) );
  NAND2_X1 U3810 ( .A1(n4543), .A2(n3459), .ZN(n4715) );
  NAND2_X1 U3811 ( .A1(n3746), .A2(n5315), .ZN(n5717) );
  INV_X1 U3812 ( .A(n5717), .ZN(n6214) );
  INV_X1 U3813 ( .A(n6201), .ZN(n6229) );
  INV_X1 U3814 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5184) );
  CLKBUF_X1 U3815 ( .A(n4318), .Z(n4319) );
  INV_X1 U3816 ( .A(n4312), .ZN(n6237) );
  CLKBUF_X1 U3817 ( .A(n4316), .Z(n4317) );
  INV_X1 U3818 ( .A(n6365), .ZN(n6371) );
  INV_X1 U3819 ( .A(n5782), .ZN(n5299) );
  INV_X1 U3821 ( .A(n6274), .ZN(n6264) );
  OR2_X1 U3822 ( .A1(n4602), .A2(n4760), .ZN(n5047) );
  INV_X1 U3823 ( .A(n6311), .ZN(n6313) );
  OR2_X1 U3824 ( .A1(n6333), .A2(n6332), .ZN(n6357) );
  NOR2_X2 U3825 ( .A1(n4682), .A2(n4760), .ZN(n6356) );
  OAI211_X1 U3826 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6374), .A(n4848), .B(n4847), .ZN(n4871) );
  INV_X1 U3827 ( .A(n5199), .ZN(n6362) );
  INV_X1 U3828 ( .A(n5219), .ZN(n6388) );
  INV_X1 U3829 ( .A(n5215), .ZN(n6394) );
  INV_X1 U3830 ( .A(n5203), .ZN(n6400) );
  INV_X1 U3831 ( .A(n5207), .ZN(n6406) );
  INV_X1 U3832 ( .A(n5197), .ZN(n5223) );
  AND2_X1 U3833 ( .A1(DATAI_6_), .A2(n4765), .ZN(n6415) );
  AND2_X1 U3834 ( .A1(n4538), .A2(n4760), .ZN(n5089) );
  OAI21_X1 U3835 ( .B1(n4890), .B2(n4889), .A(n4888), .ZN(n4921) );
  AND2_X1 U3836 ( .A1(n4761), .A2(n4312), .ZN(n4920) );
  INV_X1 U3837 ( .A(n5105), .ZN(n6421) );
  NOR2_X1 U3838 ( .A1(n5314), .A2(n6560), .ZN(n6470) );
  NAND2_X1 U3839 ( .A1(n3609), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U3840 ( .B1(n5638), .B2(n6124), .A(n3076), .ZN(U2957) );
  INV_X1 U3841 ( .A(n3766), .ZN(n3031) );
  OR2_X1 U3842 ( .A1(n5444), .A2(n5446), .ZN(n5438) );
  NAND2_X1 U3843 ( .A1(n4192), .A2(n4191), .ZN(n5374) );
  NAND2_X1 U3844 ( .A1(n3093), .A2(n3925), .ZN(n4671) );
  AND2_X1 U3845 ( .A1(n3073), .A2(n3021), .ZN(n4224) );
  AND2_X1 U3846 ( .A1(n3033), .A2(n3656), .ZN(n3007) );
  OR2_X1 U3847 ( .A1(n3556), .A2(n3626), .ZN(n3245) );
  AND2_X1 U3848 ( .A1(n3057), .A2(n3025), .ZN(n3008) );
  INV_X1 U3849 ( .A(n3863), .ZN(n3905) );
  AND2_X1 U3850 ( .A1(n3019), .A2(n3039), .ZN(n3009) );
  AND2_X1 U3851 ( .A1(n3009), .A2(n5483), .ZN(n3010) );
  NAND2_X1 U3852 ( .A1(n3053), .A2(n3057), .ZN(n5599) );
  NOR2_X1 U3853 ( .A1(n5444), .A2(n3104), .ZN(n5386) );
  AND2_X1 U3854 ( .A1(n3511), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3011)
         );
  NAND2_X1 U3855 ( .A1(n3531), .A2(n3530), .ZN(n5517) );
  AND2_X1 U3856 ( .A1(n5230), .A2(n3088), .ZN(n3012) );
  NAND2_X1 U3857 ( .A1(n3056), .A2(n3522), .ZN(n5605) );
  OR2_X1 U3858 ( .A1(n5302), .A2(n6122), .ZN(n3013) );
  AND2_X1 U3859 ( .A1(n3512), .A2(n3515), .ZN(n3014) );
  AND4_X1 U3860 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3015)
         );
  OR2_X1 U3861 ( .A1(n3512), .A2(n5898), .ZN(n3016) );
  XNOR2_X1 U3862 ( .A(n3369), .B(n3368), .ZN(n3408) );
  AND2_X1 U3863 ( .A1(n3220), .A2(n3304), .ZN(n3229) );
  INV_X1 U3864 ( .A(n3073), .ZN(n5542) );
  NAND2_X1 U3865 ( .A1(n3531), .A2(n3074), .ZN(n3073) );
  OR2_X1 U3866 ( .A1(n6130), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3017)
         );
  NAND2_X1 U3867 ( .A1(n3352), .A2(n3351), .ZN(n3383) );
  NAND2_X1 U3868 ( .A1(n3230), .A2(n3229), .ZN(n3234) );
  XNOR2_X1 U3869 ( .A(n3382), .B(n3383), .ZN(n4316) );
  OR3_X1 U3870 ( .A1(n5473), .A2(n3706), .A3(n3040), .ZN(n3018) );
  INV_X1 U3871 ( .A(n3410), .ZN(n4313) );
  NAND2_X1 U3872 ( .A1(n3227), .A2(n3219), .ZN(n3556) );
  NAND2_X1 U3873 ( .A1(n4069), .A2(n4068), .ZN(n5399) );
  AND2_X1 U3874 ( .A1(n5900), .A2(n5234), .ZN(n3019) );
  AND2_X1 U3875 ( .A1(n3083), .A2(n3082), .ZN(n3020) );
  NOR2_X1 U3876 ( .A1(n4672), .A2(n3094), .ZN(n4757) );
  NAND2_X1 U3877 ( .A1(n5230), .A2(n5232), .ZN(n5231) );
  NAND2_X1 U3878 ( .A1(n3521), .A2(n3520), .ZN(n5612) );
  NAND2_X1 U3879 ( .A1(n3512), .A2(n5670), .ZN(n3021) );
  INV_X1 U3880 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3047) );
  OR3_X1 U3881 ( .A1(n5473), .A2(n3706), .A3(n3041), .ZN(n3022) );
  OR3_X1 U3882 ( .A1(n5431), .A2(n3044), .A3(n3046), .ZN(n3023) );
  OR2_X1 U3883 ( .A1(n5473), .A2(n5464), .ZN(n3024) );
  NAND2_X1 U3884 ( .A1(n3512), .A2(n3525), .ZN(n3025) );
  INV_X1 U3885 ( .A(n4710), .ZN(n3658) );
  AND2_X1 U3886 ( .A1(n3993), .A2(n4005), .ZN(n5168) );
  INV_X1 U3887 ( .A(n4662), .ZN(n3656) );
  AND2_X1 U3888 ( .A1(n3098), .A2(n3096), .ZN(n3026) );
  AND2_X1 U3889 ( .A1(n3021), .A2(n3532), .ZN(n3027) );
  NAND2_X1 U3890 ( .A1(n3746), .A2(n3733), .ZN(n6193) );
  AND2_X1 U3891 ( .A1(n3659), .A2(n3658), .ZN(n3028) );
  NAND2_X1 U3892 ( .A1(n3080), .A2(n3079), .ZN(n4480) );
  AOI21_X1 U3893 ( .B1(n3900), .B2(n4018), .A(n3899), .ZN(n4617) );
  AND2_X1 U3894 ( .A1(n3338), .A2(n3339), .ZN(n4496) );
  AND2_X1 U3895 ( .A1(n5901), .A2(n3009), .ZN(n3029) );
  INV_X1 U3896 ( .A(n3078), .ZN(n4423) );
  INV_X1 U3897 ( .A(n3192), .ZN(n3614) );
  NOR2_X1 U3898 ( .A1(n3308), .A2(n4267), .ZN(n3620) );
  OR2_X1 U3899 ( .A1(n4484), .A2(n3644), .ZN(n4518) );
  INV_X1 U3900 ( .A(n4518), .ZN(n3032) );
  OR2_X2 U3901 ( .A1(n4737), .A2(n6455), .ZN(n6124) );
  AND2_X1 U3902 ( .A1(n5777), .A2(n6486), .ZN(n6199) );
  OAI21_X1 U3903 ( .B1(n5414), .B2(n6193), .A(n3030), .ZN(U2987) );
  INV_X1 U3904 ( .A(n5424), .ZN(n3046) );
  OAI211_X2 U3905 ( .C1(n4542), .C2(n3049), .A(n3048), .B(n4714), .ZN(n4713)
         );
  INV_X1 U3906 ( .A(n3459), .ZN(n3049) );
  NAND2_X1 U3907 ( .A1(n4542), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U3908 ( .A1(n3328), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3909 ( .A1(n3862), .A2(n3328), .ZN(n3052) );
  INV_X1 U3910 ( .A(n3521), .ZN(n3055) );
  OAI21_X1 U3911 ( .B1(n4879), .B2(n3063), .A(n3062), .ZN(n5137) );
  AOI21_X1 U3912 ( .B1(n4966), .B2(n3068), .A(n3011), .ZN(n3062) );
  INV_X1 U3913 ( .A(n4966), .ZN(n3063) );
  NAND2_X1 U3914 ( .A1(n3066), .A2(n3064), .ZN(n3513) );
  INV_X1 U3915 ( .A(n3065), .ZN(n3064) );
  OAI21_X1 U3916 ( .B1(n4966), .B2(n3011), .A(n5138), .ZN(n3065) );
  NAND2_X1 U3917 ( .A1(n4879), .A2(n3067), .ZN(n3066) );
  NAND2_X1 U3918 ( .A1(n4967), .A2(n4966), .ZN(n4965) );
  NAND3_X1 U3919 ( .A1(n3069), .A2(n3741), .A3(n3071), .ZN(n3250) );
  OAI21_X1 U3920 ( .B1(n3222), .B2(n3239), .A(n3238), .ZN(n3071) );
  OAI21_X1 U3921 ( .B1(n3234), .B2(n3237), .A(n3236), .ZN(n3072) );
  NAND2_X1 U3922 ( .A1(n3073), .A2(n3027), .ZN(n5528) );
  OAI21_X2 U3923 ( .B1(n5236), .B2(n5237), .A(n5238), .ZN(n5871) );
  NAND2_X1 U3924 ( .A1(n3077), .A2(n3156), .ZN(n3168) );
  NOR2_X1 U3925 ( .A1(n4272), .A2(n3077), .ZN(n3299) );
  NAND3_X1 U3926 ( .A1(n3078), .A2(n3856), .A3(n3988), .ZN(n4481) );
  NAND2_X1 U3927 ( .A1(n3081), .A2(n4423), .ZN(n3079) );
  NAND2_X1 U3928 ( .A1(n4481), .A2(n4482), .ZN(n3080) );
  NAND2_X1 U3929 ( .A1(n4069), .A2(n3083), .ZN(n5458) );
  NAND2_X1 U3930 ( .A1(n3085), .A2(n3084), .ZN(n3233) );
  INV_X1 U3931 ( .A(n3314), .ZN(n3345) );
  NAND2_X1 U3932 ( .A1(n3085), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U3933 ( .A1(n3231), .A2(n3593), .A3(n3596), .A4(n3247), .ZN(n3085)
         );
  NAND2_X1 U3934 ( .A1(n4192), .A2(n3098), .ZN(n5347) );
  AND2_X1 U3935 ( .A1(n4192), .A2(n3097), .ZN(n5360) );
  AND2_X2 U3936 ( .A1(n4192), .A2(n3026), .ZN(n4221) );
  NOR2_X1 U3937 ( .A1(n5444), .A2(n3102), .ZN(n5385) );
  NAND2_X1 U3938 ( .A1(n5452), .A2(n5453), .ZN(n5444) );
  AOI22_X1 U3939 ( .A1(n3204), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3208) );
  AND2_X1 U3940 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3106) );
  OR2_X1 U3941 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3107)
         );
  OR2_X1 U3942 ( .A1(n3317), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3108)
         );
  AND4_X1 U3943 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3109)
         );
  INV_X1 U3944 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6006) );
  AND2_X1 U3945 ( .A1(n4276), .A2(n4275), .ZN(n3110) );
  NOR2_X1 U3946 ( .A1(n3594), .A2(n3307), .ZN(n3221) );
  NAND2_X1 U3947 ( .A1(n3219), .A2(n3241), .ZN(n3156) );
  INV_X1 U3948 ( .A(n3461), .ZN(n3462) );
  AND2_X1 U3949 ( .A1(n5184), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3554)
         );
  INV_X1 U3950 ( .A(n5401), .ZN(n4068) );
  AND2_X1 U3951 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  INV_X1 U3952 ( .A(n3481), .ZN(n3478) );
  OR2_X1 U3953 ( .A1(n3294), .A2(n3293), .ZN(n3375) );
  NAND2_X1 U3954 ( .A1(n3318), .A2(n3108), .ZN(n3319) );
  NOR2_X1 U3955 ( .A1(n3169), .A2(n3556), .ZN(n3301) );
  INV_X1 U3956 ( .A(n3391), .ZN(n3364) );
  AOI22_X1 U3957 ( .A1(n3138), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U3958 ( .A1(n3138), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3129) );
  INV_X1 U3959 ( .A(n3579), .ZN(n3601) );
  OR2_X1 U3960 ( .A1(n3475), .A2(n3474), .ZN(n3496) );
  AOI22_X1 U3961 ( .A1(n3398), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3185) );
  AND2_X1 U3962 ( .A1(n3305), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3881) );
  INV_X1 U3963 ( .A(n4144), .ZN(n3851) );
  NOR2_X1 U3964 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  NOR2_X1 U3965 ( .A1(n4169), .A2(n5567), .ZN(n4175) );
  INV_X1 U3966 ( .A(n5267), .ZN(n5061) );
  NAND2_X1 U3967 ( .A1(n3236), .A2(n4343), .ZN(n3626) );
  INV_X1 U3968 ( .A(n3905), .ZN(n4206) );
  OR2_X1 U3969 ( .A1(n4737), .A2(n6433), .ZN(n4738) );
  NAND2_X1 U3970 ( .A1(n4006), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4021)
         );
  INV_X1 U3971 ( .A(n5586), .ZN(n5552) );
  NAND2_X1 U3972 ( .A1(n3307), .A2(n3612), .ZN(n4267) );
  NAND2_X1 U3973 ( .A1(n3390), .A2(n3389), .ZN(n4596) );
  OAI21_X1 U3974 ( .B1(n5022), .B2(n6560), .A(n5018), .ZN(n5041) );
  INV_X1 U3975 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6437) );
  OR3_X1 U3976 ( .A1(n4376), .A2(n4375), .A3(n4374), .ZN(n6439) );
  AND2_X1 U3977 ( .A1(n4175), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4188)
         );
  NAND2_X1 U3978 ( .A1(n4125), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4144)
         );
  INV_X1 U3979 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U3980 ( .A1(n4831), .A2(n6465), .ZN(n4286) );
  AND2_X1 U3981 ( .A1(n4831), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4832) );
  OR2_X1 U3982 ( .A1(n4827), .A2(n5413), .ZN(n4295) );
  AND2_X1 U3983 ( .A1(n3710), .A2(n3709), .ZN(n5440) );
  AND2_X1 U3984 ( .A1(n3681), .A2(n3680), .ZN(n5900) );
  NAND2_X1 U3985 ( .A1(n4193), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4207)
         );
  AND2_X1 U3986 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4084), .ZN(n4106)
         );
  NOR2_X1 U3987 ( .A1(n3954), .A2(n5983), .ZN(n3968) );
  NAND2_X1 U3988 ( .A1(n3920), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3926)
         );
  INV_X1 U3989 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3904) );
  AND2_X1 U3990 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3883), .ZN(n3896)
         );
  AND2_X1 U3991 ( .A1(n6242), .A2(n6241), .ZN(n6246) );
  INV_X1 U3992 ( .A(n4677), .ZN(n4682) );
  OR2_X1 U3993 ( .A1(n3873), .A2(n4312), .ZN(n6366) );
  INV_X1 U3994 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6446) );
  INV_X1 U3995 ( .A(n4765), .ZN(n5188) );
  INV_X1 U3996 ( .A(n4280), .ZN(n5310) );
  OAI21_X1 U3997 ( .B1(n5414), .B2(n6024), .A(n4302), .ZN(n4303) );
  NOR2_X1 U3998 ( .A1(n6703), .A2(n5824), .ZN(n5811) );
  AND2_X1 U3999 ( .A1(n5269), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6031) );
  INV_X1 U4000 ( .A(n5994), .ZN(n6021) );
  AND2_X1 U4001 ( .A1(n5269), .A2(n4832), .ZN(n6032) );
  NOR2_X2 U4002 ( .A1(n4295), .A2(n4288), .ZN(n6041) );
  INV_X1 U4003 ( .A(n6055), .ZN(n5479) );
  AND2_X1 U4004 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  INV_X1 U4005 ( .A(n4478), .ZN(n4459) );
  AND2_X1 U4006 ( .A1(n5458), .A2(n5471), .ZN(n6056) );
  AND2_X1 U4007 ( .A1(n5173), .A2(n5172), .ZN(n6048) );
  NOR2_X1 U4008 ( .A1(n3901), .A2(n3904), .ZN(n3902) );
  INV_X1 U4009 ( .A(n6124), .ZN(n6135) );
  OR2_X1 U4010 ( .A1(n5314), .A2(n6477), .ZN(n4737) );
  OR2_X1 U4011 ( .A1(n5689), .A2(n3756), .ZN(n5676) );
  AND2_X1 U4012 ( .A1(n6147), .A2(n6146), .ZN(n6182) );
  INV_X1 U4013 ( .A(n6191), .ZN(n6213) );
  INV_X1 U4014 ( .A(n6193), .ZN(n6223) );
  NOR2_X1 U4015 ( .A1(n4511), .A2(n6758), .ZN(n6364) );
  NOR2_X1 U4016 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5777) );
  INV_X1 U4017 ( .A(n4964), .ZN(n4586) );
  AND2_X1 U4018 ( .A1(n4359), .A2(n4358), .ZN(n4959) );
  OAI221_X1 U4019 ( .B1(n4357), .B2(n6560), .C1(n4357), .C2(n4354), .A(n4848), 
        .ZN(n4958) );
  INV_X1 U4020 ( .A(n6267), .ZN(n6268) );
  INV_X1 U4021 ( .A(n5047), .ZN(n4626) );
  OR2_X1 U4022 ( .A1(n6282), .A2(n2988), .ZN(n4602) );
  INV_X1 U4023 ( .A(n4629), .ZN(n6277) );
  INV_X1 U4024 ( .A(n4840), .ZN(n4892) );
  NAND2_X1 U4025 ( .A1(n4312), .A2(n4313), .ZN(n6282) );
  INV_X1 U4026 ( .A(n4849), .ZN(n4874) );
  INV_X1 U4027 ( .A(n5226), .ZN(n6382) );
  INV_X1 U4028 ( .A(n5211), .ZN(n6412) );
  INV_X1 U4029 ( .A(n6366), .ZN(n5177) );
  AND2_X1 U4030 ( .A1(n4538), .A2(n4314), .ZN(n5228) );
  OAI211_X1 U4031 ( .C1(n5095), .C2(n6560), .A(n5092), .B(n5091), .ZN(n5126)
         );
  AND2_X1 U4032 ( .A1(n6465), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3609) );
  INV_X1 U4033 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6465) );
  OR2_X1 U4034 ( .A1(n4737), .A2(n5310), .ZN(n4386) );
  INV_X1 U4035 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6466) );
  INV_X1 U4036 ( .A(n4303), .ZN(n4304) );
  OR2_X1 U4037 ( .A1(n4827), .A2(n4825), .ZN(n6016) );
  INV_X1 U4038 ( .A(n6041), .ZN(n6024) );
  INV_X1 U4039 ( .A(n5070), .ZN(n6038) );
  NAND2_X1 U4040 ( .A1(n3304), .A2(n6055), .ZN(n5469) );
  INV_X1 U4041 ( .A(n5256), .ZN(n5135) );
  NAND2_X1 U4042 ( .A1(n4223), .A2(n6365), .ZN(n6122) );
  NAND2_X1 U4043 ( .A1(n5616), .A2(n4233), .ZN(n6139) );
  INV_X1 U4044 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4384) );
  NAND2_X1 U4045 ( .A1(n4559), .A2(n4314), .ZN(n4820) );
  NAND2_X1 U4046 ( .A1(n4559), .A2(n4760), .ZN(n4964) );
  NAND2_X1 U4047 ( .A1(n5010), .A2(n6237), .ZN(n6274) );
  OR2_X1 U4048 ( .A1(n4602), .A2(n4314), .ZN(n4629) );
  INV_X1 U4049 ( .A(n6278), .ZN(n4736) );
  OR2_X1 U4050 ( .A1(n6282), .A2(n4892), .ZN(n6311) );
  OR2_X1 U4051 ( .A1(n6282), .A2(n6281), .ZN(n6360) );
  NAND2_X1 U4052 ( .A1(n4677), .A2(n4760), .ZN(n4849) );
  NAND2_X1 U4053 ( .A1(n5177), .A2(n4840), .ZN(n6429) );
  NAND2_X1 U4054 ( .A1(n5177), .A2(n5176), .ZN(n6418) );
  INV_X1 U4055 ( .A(n5089), .ZN(n5134) );
  INV_X1 U4057 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6560) );
  INV_X1 U4058 ( .A(n6556), .ZN(n6487) );
  AND2_X1 U4059 ( .A1(n6498), .A2(STATE_REG_1__SCAN_IN), .ZN(n6581) );
  INV_X1 U4060 ( .A(n6550), .ZN(n6547) );
  INV_X1 U4061 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3111) );
  AND2_X2 U4062 ( .A1(n3117), .A2(n5760), .ZN(n3179) );
  INV_X1 U4063 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3112) );
  AND2_X2 U4064 ( .A1(n3118), .A2(n5762), .ZN(n3266) );
  AOI22_X1 U4065 ( .A1(n3266), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4066 ( .A1(n3272), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3114) );
  AND2_X4 U4067 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4408) );
  AND2_X2 U4068 ( .A1(n5760), .A2(n4408), .ZN(n3259) );
  AOI22_X1 U4069 ( .A1(n3398), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3113) );
  AND2_X2 U4070 ( .A1(n5762), .A2(n4409), .ZN(n3273) );
  AOI22_X1 U4071 ( .A1(n3273), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4072 ( .A1(n3204), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3122) );
  AOI22_X1 U4073 ( .A1(n3157), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3121) );
  AND2_X2 U4074 ( .A1(n3119), .A2(n3118), .ZN(n3211) );
  AOI22_X1 U4075 ( .A1(n3211), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3120) );
  NAND2_X2 U4076 ( .A1(n3125), .A2(n3124), .ZN(n3219) );
  AOI22_X1 U4077 ( .A1(n3272), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4078 ( .A1(n3204), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4079 ( .A1(n3211), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4080 ( .A1(n3273), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4081 ( .A1(n3157), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4082 ( .A1(n3266), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4083 ( .A1(n3004), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U4084 ( .A1(n3157), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4085 ( .A1(n3211), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U4086 ( .A1(n3353), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3134)
         );
  NAND2_X1 U4087 ( .A1(n3138), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4088 ( .A1(n3266), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4089 ( .A1(n3179), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U4090 ( .A1(n3210), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3139)
         );
  NAND2_X1 U4091 ( .A1(n3273), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U4092 ( .A1(n3393), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3144)
         );
  NAND2_X1 U4093 ( .A1(n3204), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3143)
         );
  NAND3_X1 U4094 ( .A1(n3145), .A2(n3144), .A3(n3143), .ZN(n3146) );
  NAND2_X1 U4095 ( .A1(n3398), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3151)
         );
  NAND2_X1 U4096 ( .A1(n3272), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4097 ( .A1(n3259), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4098 ( .A1(n3180), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4099 ( .A1(n3266), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4100 ( .A1(n3157), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4101 ( .A1(n3398), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3158) );
  AND2_X1 U4102 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  AOI22_X1 U4103 ( .A1(n3273), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4104 ( .A1(n3272), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4105 ( .A1(n3179), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4106 ( .A1(n2990), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4107 ( .A1(n3272), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4108 ( .A1(n3138), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4109 ( .A1(n3398), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4110 ( .A1(n3266), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4111 ( .A1(n3157), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4112 ( .A1(n3211), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4113 ( .A1(n3273), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4114 ( .A1(n3204), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U4115 ( .A1(n3228), .A2(n4343), .ZN(n3239) );
  AOI22_X1 U4116 ( .A1(n3204), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4117 ( .A1(n3273), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4118 ( .A1(n3272), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4119 ( .A1(n3157), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3181) );
  NAND4_X1 U4120 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3190)
         );
  AOI22_X1 U4121 ( .A1(n3266), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4122 ( .A1(n3211), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3186) );
  NAND4_X1 U4123 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3189)
         );
  OR2_X2 U4124 ( .A1(n3190), .A2(n3189), .ZN(n3304) );
  AOI22_X1 U4125 ( .A1(n3273), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4126 ( .A1(n3138), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4127 ( .A1(n3179), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4128 ( .A1(n3157), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4129 ( .A1(n3266), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4130 ( .A1(n3004), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4131 ( .A1(n3211), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4132 ( .A1(n3272), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4133 ( .A1(n3203), .A2(n3612), .ZN(n3218) );
  AOI22_X1 U4134 ( .A1(n3138), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3398), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4135 ( .A1(n3273), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4136 ( .A1(n3272), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3205) );
  NAND4_X1 U4137 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3217)
         );
  AOI22_X1 U4138 ( .A1(n3266), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4139 ( .A1(n3211), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3212) );
  NAND4_X1 U4140 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3216)
         );
  INV_X1 U4141 ( .A(n3219), .ZN(n3298) );
  NAND2_X1 U4142 ( .A1(n3298), .A2(n3241), .ZN(n3220) );
  NAND2_X1 U4143 ( .A1(n3229), .A2(n3227), .ZN(n3222) );
  INV_X1 U4144 ( .A(n3228), .ZN(n3594) );
  NAND2_X1 U4145 ( .A1(n3222), .A2(n3221), .ZN(n3596) );
  AND2_X2 U4146 ( .A1(n3005), .A2(n3612), .ZN(n3238) );
  NAND2_X1 U4147 ( .A1(n3238), .A2(n3222), .ZN(n3224) );
  NAND2_X1 U4148 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6490) );
  OAI21_X1 U4149 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6490), .ZN(n3599) );
  NAND2_X1 U4150 ( .A1(n3612), .A2(n3599), .ZN(n3300) );
  NAND2_X1 U4151 ( .A1(n3300), .A2(n3298), .ZN(n3223) );
  NAND2_X1 U4152 ( .A1(n3224), .A2(n3223), .ZN(n3226) );
  INV_X1 U4153 ( .A(n3245), .ZN(n3225) );
  NOR2_X1 U4154 ( .A1(n3226), .A2(n3225), .ZN(n3231) );
  NAND2_X1 U4155 ( .A1(n5777), .A2(n6466), .ZN(n4229) );
  MUX2_X1 U4156 ( .A(n3609), .B(n4229), .S(n5184), .Z(n3232) );
  NAND2_X1 U4157 ( .A1(n3233), .A2(n3232), .ZN(n3251) );
  INV_X1 U4158 ( .A(n3251), .ZN(n3249) );
  NAND2_X1 U4159 ( .A1(n3228), .A2(n3240), .ZN(n3235) );
  NAND2_X1 U4160 ( .A1(n3235), .A2(n4343), .ZN(n3237) );
  NOR2_X1 U4161 ( .A1(n3192), .A2(n3006), .ZN(n3734) );
  INV_X1 U4162 ( .A(n3589), .ZN(n3243) );
  NOR2_X1 U4163 ( .A1(n3241), .A2(n4343), .ZN(n3242) );
  NAND3_X1 U4164 ( .A1(n3734), .A2(n3243), .A3(n3242), .ZN(n5771) );
  NAND2_X1 U4165 ( .A1(n5777), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6478) );
  AOI21_X1 U4166 ( .B1(n3192), .B2(n3244), .A(n6478), .ZN(n3246) );
  AND2_X1 U4167 ( .A1(n3549), .A2(n3227), .ZN(n3503) );
  INV_X1 U4168 ( .A(n3250), .ZN(n3248) );
  NAND2_X1 U4169 ( .A1(n3249), .A2(n3248), .ZN(n3252) );
  AOI22_X1 U4170 ( .A1(n3004), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4171 ( .A1(n4109), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4172 ( .A1(n3138), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3255) );
  INV_X1 U4173 ( .A(n3266), .ZN(n3253) );
  INV_X2 U4174 ( .A(n3253), .ZN(n4147) );
  AOI22_X1 U4175 ( .A1(n4147), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4176 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3265)
         );
  AOI22_X1 U4177 ( .A1(n4128), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4178 ( .A1(n3258), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4179 ( .A1(n3273), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4180 ( .A1(n2991), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3260) );
  NAND4_X1 U4181 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3264)
         );
  INV_X1 U4182 ( .A(n3504), .ZN(n3508) );
  AOI22_X1 U4183 ( .A1(n3157), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4184 ( .A1(n3353), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4185 ( .A1(n4147), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4186 ( .A1(n3180), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3268) );
  NAND4_X1 U4187 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3279)
         );
  AOI22_X1 U4188 ( .A1(n3002), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4189 ( .A1(n3273), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4190 ( .A1(n4128), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4191 ( .A1(n4238), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4192 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  XNOR2_X1 U4193 ( .A(n3508), .B(n3376), .ZN(n3280) );
  NAND2_X1 U4194 ( .A1(n3280), .A2(n3364), .ZN(n3328) );
  INV_X1 U4195 ( .A(n3376), .ZN(n3283) );
  NAND2_X1 U4196 ( .A1(n3577), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3282) );
  AOI21_X1 U4197 ( .B1(n3227), .B2(n3504), .A(n6466), .ZN(n3281) );
  OAI211_X1 U4198 ( .C1(n3283), .C2(n3006), .A(n3282), .B(n3281), .ZN(n3329)
         );
  NAND2_X1 U4199 ( .A1(n3364), .A2(n3504), .ZN(n3284) );
  NAND2_X1 U4200 ( .A1(n3577), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3296) );
  INV_X1 U4201 ( .A(n3392), .ZN(n3367) );
  AOI22_X1 U4202 ( .A1(n3157), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4203 ( .A1(n3266), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4204 ( .A1(n3258), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4205 ( .A1(n3002), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4206 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3294)
         );
  AOI22_X1 U4207 ( .A1(n4128), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4208 ( .A1(n3393), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4209 ( .A1(n4109), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4210 ( .A1(n3180), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3289) );
  NAND4_X1 U4211 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3293)
         );
  NAND2_X1 U4212 ( .A1(n3367), .A2(n3375), .ZN(n3295) );
  INV_X1 U4213 ( .A(n3297), .ZN(n3323) );
  NAND2_X1 U4214 ( .A1(n3298), .A2(n3304), .ZN(n4272) );
  NAND2_X1 U4215 ( .A1(n4280), .A2(n3300), .ZN(n3310) );
  NAND2_X1 U4216 ( .A1(n3307), .A2(n3301), .ZN(n3302) );
  INV_X1 U4217 ( .A(n4343), .ZN(n3625) );
  NAND3_X1 U4218 ( .A1(n3625), .A2(n3614), .A3(n3298), .ZN(n4405) );
  INV_X1 U4219 ( .A(n4405), .ZN(n3306) );
  NAND2_X1 U4220 ( .A1(n3241), .A2(n3304), .ZN(n4273) );
  INV_X1 U4221 ( .A(n4273), .ZN(n3305) );
  NAND2_X1 U4222 ( .A1(n3306), .A2(n3305), .ZN(n3308) );
  INV_X1 U4223 ( .A(n3620), .ZN(n3309) );
  NAND3_X1 U4224 ( .A1(n3310), .A2(n3622), .A3(n3309), .ZN(n3311) );
  NAND2_X1 U4225 ( .A1(n3311), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3315) );
  INV_X1 U4226 ( .A(n4229), .ZN(n3350) );
  XNOR2_X1 U4227 ( .A(n5184), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5180)
         );
  NAND2_X1 U4228 ( .A1(n3350), .A2(n5180), .ZN(n3313) );
  INV_X1 U4229 ( .A(n3609), .ZN(n3349) );
  NAND2_X1 U4230 ( .A1(n3349), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3312) );
  INV_X1 U4231 ( .A(n3315), .ZN(n3318) );
  INV_X1 U4232 ( .A(n3316), .ZN(n3317) );
  INV_X1 U4233 ( .A(n3342), .ZN(n3320) );
  NAND2_X1 U4234 ( .A1(n3364), .A2(n3375), .ZN(n3321) );
  XNOR2_X1 U4235 ( .A(n3376), .B(n3375), .ZN(n3324) );
  INV_X1 U4236 ( .A(n3238), .ZN(n6573) );
  OAI211_X1 U4237 ( .C1(n3324), .C2(n6573), .A(n3323), .B(n4337), .ZN(n3325)
         );
  INV_X1 U4238 ( .A(n3325), .ZN(n3326) );
  NAND2_X1 U4239 ( .A1(n3327), .A2(n3326), .ZN(n4497) );
  INV_X1 U4240 ( .A(n3328), .ZN(n3330) );
  OR2_X1 U4241 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  INV_X1 U4242 ( .A(n4314), .ZN(n4351) );
  NAND2_X1 U4243 ( .A1(n4351), .A2(n3549), .ZN(n3335) );
  NAND2_X1 U4244 ( .A1(n3307), .A2(n4343), .ZN(n3377) );
  OAI21_X1 U4245 ( .B1(n6573), .B2(n3376), .A(n3377), .ZN(n3333) );
  INV_X1 U4246 ( .A(n3333), .ZN(n3334) );
  NAND2_X1 U4247 ( .A1(n3335), .A2(n3334), .ZN(n4417) );
  NAND2_X1 U4248 ( .A1(n4417), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3336)
         );
  INV_X1 U4249 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U4250 ( .A1(n3336), .A2(n6234), .ZN(n3338) );
  AND2_X1 U4251 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4252 ( .A1(n4417), .A2(n3337), .ZN(n3339) );
  NAND2_X1 U4253 ( .A1(n4497), .A2(n4496), .ZN(n3340) );
  NAND2_X1 U4254 ( .A1(n6130), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3380)
         );
  NAND2_X1 U4255 ( .A1(n3342), .A2(n3341), .ZN(n3344) );
  NAND2_X1 U4256 ( .A1(n3345), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3352) );
  AND2_X1 U4257 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3346) );
  NAND2_X1 U4258 ( .A1(n3346), .A2(n4844), .ZN(n6361) );
  INV_X1 U4259 ( .A(n3346), .ZN(n3347) );
  NAND2_X1 U4260 ( .A1(n3347), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4261 ( .A1(n6361), .A2(n3348), .ZN(n4325) );
  AOI22_X1 U4262 ( .A1(n3350), .A2(n4325), .B1(n3349), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4263 ( .A1(n4316), .A2(n6466), .ZN(n3366) );
  AOI22_X1 U4264 ( .A1(n3157), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4265 ( .A1(n4128), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4266 ( .A1(n4245), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4267 ( .A1(n4109), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3354) );
  NAND4_X1 U4268 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3363)
         );
  AOI22_X1 U4269 ( .A1(n3002), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4270 ( .A1(n4147), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4271 ( .A1(n2991), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4272 ( .A1(n3258), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U4273 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3362)
         );
  AOI22_X1 U4274 ( .A1(n3577), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3367), 
        .B2(n3413), .ZN(n3368) );
  OAI21_X1 U4275 ( .B1(n3372), .B2(n3371), .A(n3370), .ZN(n3374) );
  NAND2_X1 U4276 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  XNOR2_X1 U4277 ( .A(n3408), .B(n3407), .ZN(n3855) );
  NAND2_X1 U4278 ( .A1(n3376), .A2(n3375), .ZN(n3415) );
  XNOR2_X1 U4279 ( .A(n3415), .B(n3413), .ZN(n3378) );
  OAI21_X1 U4280 ( .B1(n3378), .B2(n6573), .A(n3377), .ZN(n3379) );
  AOI21_X1 U4281 ( .B1(n3855), .B2(n3549), .A(n3379), .ZN(n6131) );
  NAND2_X1 U4282 ( .A1(n3380), .A2(n6131), .ZN(n3381) );
  AND2_X1 U4283 ( .A1(n3381), .A2(n3017), .ZN(n6121) );
  INV_X1 U4284 ( .A(n3382), .ZN(n3384) );
  NAND2_X1 U4285 ( .A1(n3345), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3390) );
  NAND3_X1 U4286 ( .A1(n6446), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6290) );
  INV_X1 U4287 ( .A(n6290), .ZN(n3385) );
  NAND2_X1 U4288 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3385), .ZN(n6283) );
  NAND2_X1 U4289 ( .A1(n6446), .A2(n6283), .ZN(n3387) );
  NAND3_X1 U4290 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5086) );
  INV_X1 U4291 ( .A(n5086), .ZN(n3386) );
  NAND2_X1 U4292 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3386), .ZN(n4917) );
  NAND2_X1 U4293 ( .A1(n3387), .A2(n4917), .ZN(n5179) );
  OAI22_X1 U4294 ( .A1(n4229), .A2(n5179), .B1(n3609), .B2(n6446), .ZN(n3388)
         );
  INV_X1 U4295 ( .A(n3388), .ZN(n3389) );
  XNOR2_X2 U4296 ( .A(n4379), .B(n4596), .ZN(n4315) );
  NAND2_X1 U4297 ( .A1(n4315), .A2(n6466), .ZN(n3406) );
  AOI22_X1 U4298 ( .A1(n5764), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4299 ( .A1(n4128), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4300 ( .A1(n4245), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4301 ( .A1(n3204), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3394) );
  NAND4_X1 U4302 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3404)
         );
  AOI22_X1 U4303 ( .A1(n3002), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4304 ( .A1(n4147), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4305 ( .A1(n2991), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4306 ( .A1(n3258), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3399) );
  NAND4_X1 U4307 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3403)
         );
  AOI22_X1 U4308 ( .A1(n3586), .A2(n3432), .B1(n3577), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3405) );
  INV_X1 U4309 ( .A(n3407), .ZN(n3409) );
  NAND3_X2 U4310 ( .A1(n3408), .A2(n3410), .A3(n3409), .ZN(n3460) );
  NAND2_X1 U4311 ( .A1(n3408), .A2(n3409), .ZN(n3411) );
  INV_X1 U4312 ( .A(n3549), .ZN(n3417) );
  INV_X1 U4313 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4314 ( .A1(n3415), .A2(n3414), .ZN(n3433) );
  XNOR2_X1 U4315 ( .A(n3433), .B(n3432), .ZN(n3416) );
  OAI22_X2 U4316 ( .A1(n3873), .A2(n3417), .B1(n6573), .B2(n3416), .ZN(n3418)
         );
  INV_X1 U4317 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6207) );
  XNOR2_X1 U4318 ( .A(n3418), .B(n6207), .ZN(n6119) );
  NAND2_X1 U4319 ( .A1(n6121), .A2(n6119), .ZN(n6120) );
  NAND2_X1 U4320 ( .A1(n3418), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3419)
         );
  NAND2_X1 U4321 ( .A1(n6120), .A2(n3419), .ZN(n4524) );
  AOI22_X1 U4322 ( .A1(n4128), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4323 ( .A1(n4147), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4324 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3258), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4325 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n2991), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3420) );
  NAND4_X1 U4326 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3429)
         );
  AOI22_X1 U4327 ( .A1(n5764), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4328 ( .A1(n4245), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4329 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3002), .B1(n3180), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4330 ( .A1(n3353), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4331 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3428)
         );
  NAND2_X1 U4332 ( .A1(n3586), .A2(n3483), .ZN(n3431) );
  NAND2_X1 U4333 ( .A1(n3577), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3430) );
  XNOR2_X1 U4334 ( .A(n3460), .B(n3463), .ZN(n3888) );
  NAND2_X1 U4335 ( .A1(n3888), .A2(n3549), .ZN(n3436) );
  NAND2_X1 U4336 ( .A1(n3433), .A2(n3432), .ZN(n3485) );
  XNOR2_X1 U4337 ( .A(n3485), .B(n3483), .ZN(n3434) );
  NAND2_X1 U4338 ( .A1(n3434), .A2(n3238), .ZN(n3435) );
  NAND2_X1 U4339 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  INV_X1 U4340 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6198) );
  XNOR2_X1 U4341 ( .A(n3437), .B(n6198), .ZN(n4523) );
  NAND2_X1 U4342 ( .A1(n3437), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3438)
         );
  INV_X1 U4343 ( .A(n3463), .ZN(n3439) );
  AOI22_X1 U4344 ( .A1(n5764), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4345 ( .A1(n4128), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4346 ( .A1(n4245), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4347 ( .A1(n3204), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4348 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3449)
         );
  AOI22_X1 U4349 ( .A1(n3002), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4350 ( .A1(n4147), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4351 ( .A1(n2991), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4352 ( .A1(n3258), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4353 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3448)
         );
  NAND2_X1 U4354 ( .A1(n3586), .A2(n3482), .ZN(n3451) );
  NAND2_X1 U4355 ( .A1(n3577), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3450) );
  XNOR2_X1 U4356 ( .A(n3452), .B(n3461), .ZN(n3900) );
  NAND2_X1 U4357 ( .A1(n3900), .A2(n3549), .ZN(n3457) );
  INV_X1 U4358 ( .A(n3483), .ZN(n3453) );
  OR2_X1 U4359 ( .A1(n3485), .A2(n3453), .ZN(n3454) );
  XNOR2_X1 U4360 ( .A(n3454), .B(n3482), .ZN(n3455) );
  NAND2_X1 U4361 ( .A1(n3455), .A2(n3238), .ZN(n3456) );
  NAND2_X1 U4362 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  INV_X1 U4363 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4550) );
  XNOR2_X1 U4364 ( .A(n3458), .B(n4550), .ZN(n4544) );
  NAND2_X1 U4365 ( .A1(n3458), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3459)
         );
  INV_X1 U4366 ( .A(n3460), .ZN(n3465) );
  NAND2_X1 U4367 ( .A1(n3465), .A2(n3464), .ZN(n3480) );
  INV_X1 U4368 ( .A(n3480), .ZN(n3479) );
  AOI22_X1 U4369 ( .A1(n5764), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4370 ( .A1(n4128), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4371 ( .A1(n4245), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4372 ( .A1(n3204), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4373 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3475)
         );
  AOI22_X1 U4374 ( .A1(n3002), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4375 ( .A1(n4147), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4376 ( .A1(n2991), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4377 ( .A1(n3258), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4378 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3474)
         );
  NAND2_X1 U4379 ( .A1(n3586), .A2(n3496), .ZN(n3477) );
  NAND2_X1 U4380 ( .A1(n3577), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U4381 ( .A1(n3480), .A2(n3481), .ZN(n3908) );
  NAND3_X1 U4382 ( .A1(n3494), .A2(n3908), .A3(n3549), .ZN(n3488) );
  NAND2_X1 U4383 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  OR2_X1 U4384 ( .A1(n3485), .A2(n3484), .ZN(n3495) );
  XNOR2_X1 U4385 ( .A(n3495), .B(n3496), .ZN(n3486) );
  NAND2_X1 U4386 ( .A1(n3486), .A2(n3238), .ZN(n3487) );
  NAND2_X1 U4387 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  INV_X1 U4388 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3745) );
  XNOR2_X1 U4389 ( .A(n3489), .B(n3745), .ZN(n4714) );
  NAND2_X1 U4390 ( .A1(n3489), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3490)
         );
  NAND2_X1 U4391 ( .A1(n3586), .A2(n3504), .ZN(n3492) );
  NAND2_X1 U4392 ( .A1(n3577), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U4393 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  NAND2_X1 U4394 ( .A1(n3891), .A2(n3549), .ZN(n3500) );
  INV_X1 U4395 ( .A(n3495), .ZN(n3497) );
  NAND2_X1 U4396 ( .A1(n3497), .A2(n3496), .ZN(n3509) );
  XNOR2_X1 U4397 ( .A(n3509), .B(n3504), .ZN(n3498) );
  NAND2_X1 U4398 ( .A1(n3498), .A2(n3238), .ZN(n3499) );
  NAND2_X1 U4399 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  INV_X1 U4400 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6186) );
  XNOR2_X1 U4401 ( .A(n3501), .B(n6186), .ZN(n4880) );
  NAND2_X1 U4402 ( .A1(n3501), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3502)
         );
  INV_X1 U4403 ( .A(n3503), .ZN(n3506) );
  NAND2_X1 U4404 ( .A1(n3504), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3505) );
  NAND2_X4 U4405 ( .A1(n3494), .A2(n3507), .ZN(n3512) );
  OR3_X1 U4406 ( .A1(n3509), .A2(n3508), .A3(n6573), .ZN(n3510) );
  NAND2_X1 U4407 ( .A1(n3512), .A2(n3510), .ZN(n3511) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6177) );
  INV_X1 U4409 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U4410 ( .A1(n3512), .A2(n6148), .ZN(n5138) );
  NAND2_X1 U4411 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5139)
         );
  NAND2_X1 U4412 ( .A1(n3513), .A2(n5139), .ZN(n5162) );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4414 ( .A1(n3512), .A2(n3514), .ZN(n5163) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4416 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U4417 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3516) );
  AND2_X1 U4418 ( .A1(n6104), .A2(n3516), .ZN(n3517) );
  INV_X1 U4419 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3518) );
  NOR2_X1 U4420 ( .A1(n3512), .A2(n3518), .ZN(n5237) );
  NAND2_X1 U4421 ( .A1(n3512), .A2(n3518), .ZN(n5238) );
  XNOR2_X1 U4422 ( .A(n3512), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5870)
         );
  NAND2_X1 U4423 ( .A1(n5871), .A2(n5870), .ZN(n3521) );
  INV_X1 U4424 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4425 ( .A1(n3512), .A2(n3519), .ZN(n3520) );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U4427 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3522) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U4429 ( .A1(n3512), .A2(n5898), .ZN(n3524) );
  AND2_X1 U4430 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4431 ( .A1(n3760), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3525) );
  INV_X1 U4432 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5856) );
  INV_X1 U4433 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5859) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5874) );
  NAND3_X1 U4435 ( .A1(n5856), .A2(n5859), .A3(n5874), .ZN(n3526) );
  NAND2_X1 U4436 ( .A1(n5857), .A2(n3526), .ZN(n3527) );
  NAND2_X1 U4437 ( .A1(n5549), .A2(n3527), .ZN(n5548) );
  NAND2_X1 U4438 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3762) );
  AND2_X1 U4439 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5695) );
  AND2_X1 U4440 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U4441 ( .A1(n5695), .A2(n5707), .ZN(n5565) );
  OAI21_X1 U4442 ( .B1(n3762), .B2(n5565), .A(n3512), .ZN(n3528) );
  NAND2_X1 U4443 ( .A1(n5548), .A2(n3528), .ZN(n3531) );
  NOR2_X1 U4444 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5675) );
  NOR2_X1 U4445 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5694) );
  NOR2_X1 U4446 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5708) );
  NAND3_X1 U4447 ( .A1(n5675), .A2(n5694), .A3(n5708), .ZN(n3529) );
  NAND2_X1 U4448 ( .A1(n5857), .A2(n3529), .ZN(n3530) );
  XOR2_X1 U4449 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n3512), .Z(n5543) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5670) );
  AND2_X1 U4451 ( .A1(n3512), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3532)
         );
  NAND2_X1 U4452 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U4453 ( .A1(n5508), .A2(n3106), .ZN(n3535) );
  NOR2_X1 U4454 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5643) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U4456 ( .A1(n5643), .A2(n5519), .ZN(n3533) );
  NOR2_X1 U4457 ( .A1(n3512), .A2(n3533), .ZN(n4225) );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5624) );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5632) );
  NAND3_X1 U4460 ( .A1(n4225), .A2(n5624), .A3(n5632), .ZN(n3534) );
  NAND2_X1 U4461 ( .A1(n3535), .A2(n3105), .ZN(n3536) );
  XNOR2_X1 U4462 ( .A(n3536), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4309)
         );
  XNOR2_X1 U4463 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4464 ( .A1(n3554), .A2(n3550), .ZN(n3538) );
  NAND2_X1 U4465 ( .A1(n6437), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4466 ( .A1(n3538), .A2(n3537), .ZN(n3567) );
  XNOR2_X1 U4467 ( .A(n4844), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3566)
         );
  INV_X1 U4468 ( .A(n3566), .ZN(n3539) );
  NAND2_X1 U4469 ( .A1(n3567), .A2(n3539), .ZN(n3541) );
  NAND2_X1 U4470 ( .A1(n4844), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U4471 ( .A1(n3541), .A2(n3540), .ZN(n3544) );
  XNOR2_X1 U4472 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U4473 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3582), .ZN(n3542) );
  NOR2_X1 U4474 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3542), .ZN(n3548)
         );
  NOR2_X1 U4475 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  OR2_X1 U4476 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  INV_X1 U4477 ( .A(n3550), .ZN(n3551) );
  XNOR2_X1 U4478 ( .A(n3551), .B(n3554), .ZN(n3603) );
  NAND2_X1 U4479 ( .A1(n3586), .A2(n3236), .ZN(n3552) );
  NAND2_X1 U4480 ( .A1(n3552), .A2(n4337), .ZN(n3563) );
  AND2_X1 U4481 ( .A1(n3047), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3553)
         );
  NOR2_X1 U4482 ( .A1(n3554), .A2(n3553), .ZN(n3557) );
  NAND2_X1 U4483 ( .A1(n3586), .A2(n3557), .ZN(n3555) );
  NAND2_X1 U4484 ( .A1(n3578), .A2(n3555), .ZN(n3562) );
  NAND2_X1 U4485 ( .A1(n3556), .A2(n3557), .ZN(n3558) );
  NAND2_X1 U4486 ( .A1(n3558), .A2(n3006), .ZN(n3560) );
  NAND2_X1 U4487 ( .A1(n3298), .A2(n3244), .ZN(n3559) );
  NAND2_X1 U4488 ( .A1(n3559), .A2(n3612), .ZN(n3572) );
  NAND2_X1 U4489 ( .A1(n3560), .A2(n3572), .ZN(n3561) );
  OAI211_X1 U4490 ( .C1(n3563), .C2(n3603), .A(n3562), .B(n3561), .ZN(n3565)
         );
  NAND3_X1 U4491 ( .A1(n3563), .A2(STATE2_REG_0__SCAN_IN), .A3(n3603), .ZN(
        n3564) );
  OAI211_X1 U4492 ( .C1(n3578), .C2(n3603), .A(n3565), .B(n3564), .ZN(n3571)
         );
  XNOR2_X1 U4493 ( .A(n3567), .B(n3566), .ZN(n3602) );
  INV_X1 U4494 ( .A(n3577), .ZN(n3569) );
  NAND2_X1 U4495 ( .A1(n3586), .A2(n3602), .ZN(n3568) );
  OAI211_X1 U4496 ( .C1(n3602), .C2(n3569), .A(n3568), .B(n3572), .ZN(n3570)
         );
  NAND2_X1 U4497 ( .A1(n3571), .A2(n3570), .ZN(n3575) );
  INV_X1 U4498 ( .A(n3572), .ZN(n3573) );
  NAND3_X1 U4499 ( .A1(n3573), .A2(n3602), .A3(n3586), .ZN(n3574) );
  NAND2_X1 U4500 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  OAI21_X1 U4501 ( .B1(n3577), .B2(n3601), .A(n3576), .ZN(n3581) );
  AOI22_X1 U4502 ( .A1(n3579), .A2(n3583), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6466), .ZN(n3580) );
  NAND2_X1 U4503 ( .A1(n3581), .A2(n3580), .ZN(n3585) );
  OAI222_X1 U4504 ( .A1(n4384), .A2(n3582), .B1(n4384), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3582), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4505 ( .A1(n3600), .A2(n3583), .ZN(n3584) );
  INV_X1 U4506 ( .A(n5296), .ZN(n3590) );
  NAND2_X1 U4507 ( .A1(n3590), .A2(n3236), .ZN(n3743) );
  INV_X1 U4508 ( .A(n3743), .ZN(n3591) );
  NAND2_X1 U4509 ( .A1(n5314), .A2(n3591), .ZN(n3608) );
  NAND2_X1 U4510 ( .A1(n5296), .A2(n3307), .ZN(n3592) );
  NAND2_X1 U4511 ( .A1(n3593), .A2(n3592), .ZN(n3619) );
  NAND2_X1 U4512 ( .A1(n3594), .A2(n3238), .ZN(n3595) );
  NAND2_X1 U4513 ( .A1(n3596), .A2(n3595), .ZN(n3739) );
  OR2_X1 U4514 ( .A1(n3619), .A2(n3739), .ZN(n3598) );
  INV_X1 U4515 ( .A(n3597), .ZN(n4281) );
  NAND2_X1 U4516 ( .A1(n3598), .A2(n4281), .ZN(n4371) );
  OR2_X1 U4517 ( .A1(n3599), .A2(STATE_REG_0__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U4518 ( .A1(n3236), .A2(n6495), .ZN(n3606) );
  INV_X1 U4519 ( .A(n3600), .ZN(n3605) );
  NAND3_X1 U4520 ( .A1(n3603), .A2(n3602), .A3(n3601), .ZN(n3604) );
  NAND2_X1 U4521 ( .A1(n3605), .A2(n3604), .ZN(n5312) );
  NOR2_X1 U4522 ( .A1(READY_N), .A2(n5312), .ZN(n4264) );
  NAND3_X1 U4523 ( .A1(n3606), .A2(n4264), .A3(n3192), .ZN(n3607) );
  NAND3_X1 U4524 ( .A1(n3608), .A2(n4371), .A3(n3607), .ZN(n3610) );
  NAND2_X1 U4525 ( .A1(n3610), .A2(n4431), .ZN(n3618) );
  NAND2_X1 U4526 ( .A1(n3612), .A2(n6495), .ZN(n4289) );
  NAND3_X1 U4527 ( .A1(n3611), .A2(n4287), .A3(n4289), .ZN(n3613) );
  NAND3_X1 U4528 ( .A1(n3613), .A2(n3244), .A3(n4273), .ZN(n3615) );
  NAND2_X1 U4529 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  OR2_X1 U4530 ( .A1(n3619), .A2(n4267), .ZN(n5311) );
  NAND2_X1 U4531 ( .A1(n3620), .A2(n3240), .ZN(n3621) );
  NAND2_X1 U4532 ( .A1(n3611), .A2(n3638), .ZN(n4269) );
  AND2_X1 U4533 ( .A1(n3621), .A2(n4269), .ZN(n3623) );
  NAND4_X1 U4534 ( .A1(n5311), .A2(n6455), .A3(n3623), .A4(n2993), .ZN(n3624)
         );
  INV_X1 U4535 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U4536 ( .A1(n3695), .A2(n4828), .ZN(n3630) );
  NAND2_X1 U4537 ( .A1(n3625), .A2(n3244), .ZN(n3639) );
  NAND2_X1 U4538 ( .A1(n3639), .A2(n6234), .ZN(n3628) );
  NAND2_X1 U4539 ( .A1(n3638), .A2(n4828), .ZN(n3627) );
  NAND3_X1 U4540 ( .A1(n3628), .A2(n5454), .A3(n3627), .ZN(n3629) );
  NAND2_X1 U4541 ( .A1(n3630), .A2(n3629), .ZN(n3634) );
  NAND2_X1 U4542 ( .A1(n3639), .A2(EBX_REG_0__SCAN_IN), .ZN(n3632) );
  INV_X1 U4543 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U4544 ( .A1(n5454), .A2(n4972), .ZN(n3631) );
  NAND2_X1 U4545 ( .A1(n3632), .A2(n3631), .ZN(n4419) );
  XNOR2_X1 U4546 ( .A(n3634), .B(n4419), .ZN(n4830) );
  NAND2_X1 U4547 ( .A1(n4830), .A2(n3638), .ZN(n4433) );
  INV_X1 U4548 ( .A(n4419), .ZN(n3633) );
  OR2_X1 U4549 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  NAND2_X1 U4550 ( .A1(n4433), .A2(n3635), .ZN(n4484) );
  MUX2_X1 U4551 ( .A(n3723), .B(n5454), .S(EBX_REG_3__SCAN_IN), .Z(n3636) );
  OAI21_X1 U4552 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4418), .A(n3636), 
        .ZN(n3637) );
  INV_X1 U4553 ( .A(n3637), .ZN(n4491) );
  MUX2_X1 U4554 ( .A(n3727), .B(n3639), .S(EBX_REG_2__SCAN_IN), .Z(n3643) );
  INV_X1 U4555 ( .A(n3639), .ZN(n3640) );
  NAND2_X1 U4556 ( .A1(n4368), .A2(n3640), .ZN(n3689) );
  NAND3_X1 U4557 ( .A1(n4368), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n5454), 
        .ZN(n3641) );
  AND2_X1 U4558 ( .A1(n3689), .A2(n3641), .ZN(n3642) );
  NAND2_X1 U4559 ( .A1(n3643), .A2(n3642), .ZN(n4492) );
  NAND2_X1 U4560 ( .A1(n4491), .A2(n4492), .ZN(n3644) );
  INV_X1 U4561 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U4562 ( .A1(n3695), .A2(n4520), .ZN(n3648) );
  NAND2_X1 U4563 ( .A1(n3639), .A2(n6198), .ZN(n3646) );
  NAND2_X1 U4564 ( .A1(n3638), .A2(n4520), .ZN(n3645) );
  NAND3_X1 U4565 ( .A1(n3646), .A2(n5454), .A3(n3645), .ZN(n3647) );
  AND2_X1 U4566 ( .A1(n3648), .A2(n3647), .ZN(n4517) );
  MUX2_X1 U4567 ( .A(n3723), .B(n5454), .S(EBX_REG_5__SCAN_IN), .Z(n3649) );
  INV_X1 U4568 ( .A(n3649), .ZN(n3651) );
  NOR2_X1 U4569 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3650)
         );
  NOR2_X1 U4570 ( .A1(n3651), .A2(n3650), .ZN(n4552) );
  INV_X1 U4571 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U4572 ( .A1(n3695), .A2(n6017), .ZN(n3655) );
  NAND2_X1 U4573 ( .A1(n3639), .A2(n3745), .ZN(n3653) );
  NAND2_X1 U4574 ( .A1(n3638), .A2(n6017), .ZN(n3652) );
  NAND3_X1 U4575 ( .A1(n3653), .A2(n5454), .A3(n3652), .ZN(n3654) );
  AND2_X1 U4576 ( .A1(n3655), .A2(n3654), .ZN(n4662) );
  MUX2_X1 U4577 ( .A(n3723), .B(n5454), .S(EBX_REG_7__SCAN_IN), .Z(n3657) );
  NAND2_X1 U4578 ( .A1(n3107), .A2(n3657), .ZN(n4710) );
  MUX2_X1 U4579 ( .A(n3727), .B(n3639), .S(EBX_REG_8__SCAN_IN), .Z(n3662) );
  NAND2_X1 U4580 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n4368), .ZN(n3660)
         );
  AND2_X1 U4581 ( .A1(n3689), .A2(n3660), .ZN(n3661) );
  NAND2_X1 U4582 ( .A1(n3662), .A2(n3661), .ZN(n4696) );
  INV_X1 U4583 ( .A(n4696), .ZN(n3663) );
  MUX2_X1 U4584 ( .A(n3723), .B(n5454), .S(EBX_REG_9__SCAN_IN), .Z(n3664) );
  INV_X1 U4585 ( .A(n3664), .ZN(n3666) );
  NOR2_X1 U4586 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3665)
         );
  NOR2_X1 U4587 ( .A1(n3666), .A2(n3665), .ZN(n4809) );
  MUX2_X1 U4588 ( .A(n3727), .B(n3639), .S(EBX_REG_10__SCAN_IN), .Z(n3669) );
  NAND2_X1 U4589 ( .A1(n4368), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3667) );
  AND2_X1 U4590 ( .A1(n3689), .A2(n3667), .ZN(n3668) );
  NAND2_X1 U4591 ( .A1(n3669), .A2(n3668), .ZN(n5978) );
  INV_X1 U4592 ( .A(n3723), .ZN(n3716) );
  INV_X1 U4593 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U4594 ( .A1(n3716), .A2(n6054), .ZN(n3673) );
  NAND2_X1 U4595 ( .A1(n3638), .A2(n6054), .ZN(n3671) );
  NAND2_X1 U4596 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3670) );
  NAND3_X1 U4597 ( .A1(n3671), .A2(n3639), .A3(n3670), .ZN(n3672) );
  AND2_X1 U4598 ( .A1(n3673), .A2(n3672), .ZN(n5977) );
  NAND2_X1 U4599 ( .A1(n5978), .A2(n5977), .ZN(n3674) );
  MUX2_X1 U4600 ( .A(n3727), .B(n3639), .S(EBX_REG_12__SCAN_IN), .Z(n3677) );
  NAND2_X1 U4601 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4368), .ZN(n3675) );
  AND2_X1 U4602 ( .A1(n3689), .A2(n3675), .ZN(n3676) );
  INV_X1 U4603 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U4604 ( .A1(n3716), .A2(n6050), .ZN(n3681) );
  NAND2_X1 U4605 ( .A1(n3638), .A2(n6050), .ZN(n3679) );
  NAND2_X1 U4606 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3678) );
  NAND3_X1 U4607 ( .A1(n3679), .A2(n3639), .A3(n3678), .ZN(n3680) );
  MUX2_X1 U4608 ( .A(n3727), .B(n3639), .S(EBX_REG_14__SCAN_IN), .Z(n3684) );
  NAND2_X1 U4609 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4368), .ZN(n3682) );
  AND2_X1 U4610 ( .A1(n3689), .A2(n3682), .ZN(n3683) );
  NAND2_X1 U4611 ( .A1(n3684), .A2(n3683), .ZN(n5234) );
  INV_X1 U4612 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U4613 ( .A1(n3638), .A2(n5275), .ZN(n3686) );
  NAND2_X1 U4614 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3685) );
  NAND3_X1 U4615 ( .A1(n3686), .A2(n3639), .A3(n3685), .ZN(n3687) );
  OAI21_X1 U4616 ( .B1(n3723), .B2(EBX_REG_15__SCAN_IN), .A(n3687), .ZN(n5261)
         );
  MUX2_X1 U4617 ( .A(n3727), .B(n3639), .S(EBX_REG_16__SCAN_IN), .Z(n3691) );
  NAND2_X1 U4618 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4368), .ZN(n3688) );
  AND2_X1 U4619 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  NAND2_X1 U4620 ( .A1(n3691), .A2(n3690), .ZN(n5483) );
  INV_X1 U4621 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U4622 ( .A1(n3638), .A2(n5406), .ZN(n3693) );
  NAND2_X1 U4623 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3692) );
  NAND3_X1 U4624 ( .A1(n3693), .A2(n3639), .A3(n3692), .ZN(n3694) );
  OAI21_X1 U4625 ( .B1(n3723), .B2(EBX_REG_17__SCAN_IN), .A(n3694), .ZN(n5410)
         );
  INV_X1 U4626 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U4627 ( .A1(n3695), .A2(n5842), .ZN(n3699) );
  INV_X1 U4628 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U4629 ( .A1(n3639), .A2(n5721), .ZN(n3697) );
  NAND2_X1 U4630 ( .A1(n3638), .A2(n5842), .ZN(n3696) );
  NAND3_X1 U4631 ( .A1(n3697), .A2(n5454), .A3(n3696), .ZN(n3698) );
  AND2_X1 U4632 ( .A1(n3699), .A2(n3698), .ZN(n5464) );
  OR2_X1 U4633 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3702)
         );
  INV_X1 U4634 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4635 ( .A1(n3638), .A2(n3700), .ZN(n3701) );
  AND2_X1 U4636 ( .A1(n3702), .A2(n3701), .ZN(n5455) );
  OR2_X1 U4637 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3703)
         );
  INV_X1 U4638 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U4639 ( .A1(n3638), .A2(n5477), .ZN(n5462) );
  NAND2_X1 U4640 ( .A1(n3703), .A2(n5462), .ZN(n5463) );
  NAND2_X1 U4641 ( .A1(n5461), .A2(EBX_REG_20__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4642 ( .A1(n5463), .A2(n5454), .ZN(n3704) );
  OAI211_X1 U4643 ( .C1(n5455), .C2(n5463), .A(n3705), .B(n3704), .ZN(n3706)
         );
  MUX2_X1 U4644 ( .A(n3723), .B(n5454), .S(EBX_REG_21__SCAN_IN), .Z(n3707) );
  OAI21_X1 U4645 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4418), .A(n3707), 
        .ZN(n3708) );
  INV_X1 U4646 ( .A(n3708), .ZN(n5447) );
  MUX2_X1 U4647 ( .A(n3727), .B(n3639), .S(EBX_REG_22__SCAN_IN), .Z(n3710) );
  NAND2_X1 U4648 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n4368), .ZN(n3709) );
  INV_X1 U4649 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U4650 ( .A1(n3638), .A2(n5435), .ZN(n3712) );
  NAND2_X1 U4651 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3711) );
  NAND3_X1 U4652 ( .A1(n3712), .A2(n3639), .A3(n3711), .ZN(n3713) );
  OAI21_X1 U4653 ( .B1(n3723), .B2(EBX_REG_23__SCAN_IN), .A(n3713), .ZN(n5390)
         );
  MUX2_X1 U4654 ( .A(n3727), .B(n3639), .S(EBX_REG_24__SCAN_IN), .Z(n3715) );
  NAND2_X1 U4655 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4368), .ZN(n3714) );
  INV_X1 U4656 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U4657 ( .A1(n3716), .A2(n5427), .ZN(n3720) );
  NAND2_X1 U4658 ( .A1(n3638), .A2(n5427), .ZN(n3718) );
  NAND2_X1 U4659 ( .A1(n5454), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3717) );
  NAND3_X1 U4660 ( .A1(n3718), .A2(n3639), .A3(n3717), .ZN(n3719) );
  AND2_X1 U4661 ( .A1(n3720), .A2(n3719), .ZN(n5424) );
  MUX2_X1 U4662 ( .A(n3727), .B(n3639), .S(EBX_REG_26__SCAN_IN), .Z(n3722) );
  NAND2_X1 U4663 ( .A1(n4368), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U4664 ( .A1(n3722), .A2(n3721), .ZN(n5377) );
  MUX2_X1 U4665 ( .A(n3723), .B(n5454), .S(EBX_REG_27__SCAN_IN), .Z(n3724) );
  OAI21_X1 U4666 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4418), .A(n3724), 
        .ZN(n5362) );
  MUX2_X1 U4667 ( .A(n3727), .B(n3639), .S(EBX_REG_28__SCAN_IN), .Z(n3726) );
  NAND2_X1 U4668 ( .A1(n4368), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4669 ( .A1(n3726), .A2(n3725), .ZN(n5349) );
  OAI22_X1 U4670 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n4368), .B2(EBX_REG_29__SCAN_IN), .ZN(n5307) );
  NOR2_X1 U4671 ( .A1(n3727), .A2(EBX_REG_29__SCAN_IN), .ZN(n5305) );
  INV_X1 U4672 ( .A(n5351), .ZN(n5324) );
  AOI22_X1 U4673 ( .A1(n5326), .A2(n5454), .B1(n5305), .B2(n5324), .ZN(n5309)
         );
  NAND2_X1 U4674 ( .A1(n4418), .A2(EBX_REG_30__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4675 ( .A1(n4368), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4676 ( .A1(n3729), .A2(n3728), .ZN(n5327) );
  INV_X1 U4677 ( .A(n5326), .ZN(n5325) );
  NAND2_X1 U4678 ( .A1(n5325), .A2(n5454), .ZN(n5329) );
  OAI21_X1 U4679 ( .B1(n5309), .B2(n5327), .A(n5329), .ZN(n3731) );
  OAI22_X1 U4680 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4368), .B2(EBX_REG_31__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4681 ( .A1(n3620), .A2(n3227), .ZN(n3732) );
  NAND2_X1 U4682 ( .A1(n3611), .A2(n3238), .ZN(n4385) );
  NAND2_X1 U4683 ( .A1(n3732), .A2(n4385), .ZN(n3733) );
  AND2_X1 U4684 ( .A1(n3734), .A2(n3236), .ZN(n4370) );
  OAI21_X1 U4685 ( .B1(n4370), .B2(n4418), .A(n3297), .ZN(n3737) );
  OAI21_X1 U4686 ( .B1(n4273), .B2(n3244), .A(n3192), .ZN(n3736) );
  NAND2_X1 U4687 ( .A1(n3234), .A2(n5461), .ZN(n3735) );
  NAND3_X1 U4688 ( .A1(n3737), .A2(n3736), .A3(n3735), .ZN(n3738) );
  NOR2_X1 U4689 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  NAND2_X1 U4690 ( .A1(n3741), .A2(n3740), .ZN(n3744) );
  INV_X1 U4691 ( .A(n3744), .ZN(n4407) );
  OAI211_X1 U4692 ( .C1(n3245), .C2(n3006), .A(n4407), .B(n5771), .ZN(n3742)
         );
  NAND2_X1 U4693 ( .A1(n3746), .A2(n3742), .ZN(n5743) );
  AND2_X1 U4694 ( .A1(n3597), .A2(n3236), .ZN(n5769) );
  NAND2_X1 U4695 ( .A1(n3746), .A2(n5769), .ZN(n5906) );
  NAND2_X1 U4696 ( .A1(n4548), .A2(n5717), .ZN(n6221) );
  INV_X1 U4697 ( .A(n6221), .ZN(n6157) );
  NAND2_X1 U4698 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U4699 ( .A1(n3519), .A2(n5904), .ZN(n5742) );
  NAND2_X1 U4700 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5742), .ZN(n5892) );
  NAND2_X1 U4701 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5733) );
  NOR2_X1 U4702 ( .A1(n5892), .A2(n5733), .ZN(n3759) );
  INV_X1 U4703 ( .A(n4548), .ZN(n6156) );
  NOR2_X1 U4704 ( .A1(n6207), .A2(n6198), .ZN(n6189) );
  NAND2_X1 U4705 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6189), .ZN(n4718)
         );
  NOR2_X1 U4706 ( .A1(n3745), .A2(n4718), .ZN(n6147) );
  NAND3_X1 U4707 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6147), .ZN(n6155) );
  NAND2_X1 U4708 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6174) );
  INV_X1 U4709 ( .A(n6174), .ZN(n6158) );
  NAND3_X1 U4710 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6158), .ZN(n3748) );
  NOR2_X1 U4711 ( .A1(n6155), .A2(n3748), .ZN(n5744) );
  INV_X1 U4712 ( .A(n5744), .ZN(n5905) );
  INV_X1 U4713 ( .A(n3746), .ZN(n3747) );
  NAND2_X1 U4714 ( .A1(n6466), .A2(n6374), .ZN(n6476) );
  INV_X1 U4715 ( .A(n6476), .ZN(n6486) );
  INV_X1 U4716 ( .A(n6199), .ZN(n6191) );
  NAND2_X1 U4717 ( .A1(n3747), .A2(n6191), .ZN(n6233) );
  OAI21_X1 U4718 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5743), .A(n6233), 
        .ZN(n6153) );
  AOI21_X1 U4719 ( .B1(n6156), .B2(n5905), .A(n6153), .ZN(n5242) );
  OAI21_X1 U4720 ( .B1(n4548), .B2(n3759), .A(n5242), .ZN(n5714) );
  INV_X1 U4721 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U4722 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U4723 ( .A1(n6211), .A2(n6210), .ZN(n6209) );
  NAND2_X1 U4724 ( .A1(n6147), .A2(n6209), .ZN(n6152) );
  NOR2_X1 U4725 ( .A1(n3748), .A2(n6152), .ZN(n5241) );
  NAND2_X1 U4726 ( .A1(n5241), .A2(n3759), .ZN(n5711) );
  INV_X1 U4727 ( .A(n5711), .ZN(n3749) );
  NAND3_X1 U4728 ( .A1(n3749), .A2(n5707), .A3(n3760), .ZN(n3750) );
  AND2_X1 U4729 ( .A1(n6221), .A2(n3750), .ZN(n3751) );
  NOR2_X1 U4730 ( .A1(n5714), .A2(n3751), .ZN(n5692) );
  INV_X1 U4731 ( .A(n5695), .ZN(n3761) );
  NAND2_X1 U4732 ( .A1(n6221), .A2(n3761), .ZN(n3752) );
  NAND2_X1 U4733 ( .A1(n5692), .A2(n3752), .ZN(n5689) );
  INV_X1 U4734 ( .A(n5906), .ZN(n3753) );
  NOR2_X1 U4735 ( .A1(n3753), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6227)
         );
  INV_X1 U4736 ( .A(n4545), .ZN(n3755) );
  INV_X1 U4737 ( .A(n3762), .ZN(n3754) );
  AOI21_X1 U4738 ( .B1(n5717), .B2(n3755), .A(n3754), .ZN(n3756) );
  INV_X1 U4739 ( .A(n5676), .ZN(n3758) );
  NAND2_X1 U4740 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4741 ( .A1(n6221), .A2(n3763), .ZN(n3757) );
  NAND2_X1 U4742 ( .A1(n3758), .A2(n3757), .ZN(n5655) );
  AOI21_X1 U4743 ( .B1(n6221), .B2(n5641), .A(n5655), .ZN(n5633) );
  OAI21_X1 U4744 ( .B1(n6157), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5633), 
        .ZN(n5620) );
  AOI21_X1 U4745 ( .B1(n6221), .B2(n5624), .A(n5620), .ZN(n3765) );
  INV_X1 U4746 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U4747 ( .A1(n6213), .A2(REIP_REG_31__SCAN_IN), .ZN(n4307) );
  NAND2_X1 U4748 ( .A1(n4545), .A2(n5744), .ZN(n5875) );
  NAND2_X1 U4749 ( .A1(n6214), .A2(n5241), .ZN(n5747) );
  NAND2_X1 U4750 ( .A1(n5875), .A2(n5747), .ZN(n6141) );
  NAND2_X1 U4751 ( .A1(n6141), .A2(n3759), .ZN(n5885) );
  INV_X1 U4752 ( .A(n3760), .ZN(n5715) );
  NOR2_X1 U4753 ( .A1(n5885), .A2(n5715), .ZN(n5722) );
  NAND2_X1 U4754 ( .A1(n5722), .A2(n5707), .ZN(n5701) );
  NOR2_X1 U4755 ( .A1(n5686), .A2(n3762), .ZN(n5671) );
  INV_X1 U4756 ( .A(n3763), .ZN(n5659) );
  NAND2_X1 U4757 ( .A1(n5671), .A2(n5659), .ZN(n5650) );
  NOR3_X1 U4758 ( .A1(n5650), .A2(n5632), .A3(n5641), .ZN(n5621) );
  NAND3_X1 U4759 ( .A1(n5621), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4412), .ZN(n3764) );
  OAI211_X1 U4760 ( .C1(n3765), .C2(n4412), .A(n4307), .B(n3764), .ZN(n3766)
         );
  AOI22_X1 U4761 ( .A1(n3157), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4762 ( .A1(n4245), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4763 ( .A1(n4147), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4764 ( .A1(n3180), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4765 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3777)
         );
  AOI22_X1 U4766 ( .A1(n3211), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4767 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n2991), .B1(n3258), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4768 ( .A1(n3002), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4769 ( .A1(n4109), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4770 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3776)
         );
  NOR2_X1 U4771 ( .A1(n3777), .A2(n3776), .ZN(n4201) );
  AOI22_X1 U4772 ( .A1(n5764), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4773 ( .A1(n4128), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4109), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4774 ( .A1(n4147), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4775 ( .A1(n3002), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4776 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3787)
         );
  AOI22_X1 U4777 ( .A1(n4245), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4778 ( .A1(n2991), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4779 ( .A1(n3258), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4780 ( .A1(n2990), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4781 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3786)
         );
  NOR2_X1 U4782 ( .A1(n3787), .A2(n3786), .ZN(n4180) );
  AOI22_X1 U4783 ( .A1(n5764), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4784 ( .A1(n4128), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4785 ( .A1(n3273), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4786 ( .A1(n3204), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4787 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4788 ( .A1(n3002), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4789 ( .A1(n4147), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4790 ( .A1(n2991), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4791 ( .A1(n3258), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4792 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  NOR2_X1 U4793 ( .A1(n3797), .A2(n3796), .ZN(n4166) );
  AOI22_X1 U4794 ( .A1(n3838), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4795 ( .A1(n3002), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4796 ( .A1(n4109), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4797 ( .A1(n2991), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3798) );
  NAND4_X1 U4798 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3807)
         );
  AOI22_X1 U4799 ( .A1(n4128), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5764), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4800 ( .A1(n4147), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4801 ( .A1(n3393), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4802 ( .A1(n4114), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4803 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3806)
         );
  NOR2_X1 U4804 ( .A1(n3807), .A2(n3806), .ZN(n4165) );
  OR2_X1 U4805 ( .A1(n4166), .A2(n4165), .ZN(n4174) );
  AOI22_X1 U4806 ( .A1(n3004), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4807 ( .A1(n5764), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4808 ( .A1(n3002), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4809 ( .A1(n4147), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4810 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3817)
         );
  AOI22_X1 U4811 ( .A1(n4128), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4812 ( .A1(n4109), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4813 ( .A1(n4244), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4814 ( .A1(n4238), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4815 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3816)
         );
  NOR2_X1 U4816 ( .A1(n3817), .A2(n3816), .ZN(n4173) );
  OR2_X1 U4817 ( .A1(n4174), .A2(n4173), .ZN(n4181) );
  NOR2_X1 U4818 ( .A1(n4180), .A2(n4181), .ZN(n4196) );
  AOI22_X1 U4819 ( .A1(n3157), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4820 ( .A1(n4128), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4821 ( .A1(n4245), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4822 ( .A1(n4109), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4823 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3827)
         );
  AOI22_X1 U4824 ( .A1(n3002), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4825 ( .A1(n4147), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4826 ( .A1(n2991), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4827 ( .A1(n3258), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3822) );
  NAND4_X1 U4828 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3826)
         );
  OR2_X1 U4829 ( .A1(n3827), .A2(n3826), .ZN(n4195) );
  NAND2_X1 U4830 ( .A1(n4196), .A2(n4195), .ZN(n4202) );
  NOR2_X1 U4831 ( .A1(n4201), .A2(n4202), .ZN(n4215) );
  AOI22_X1 U4832 ( .A1(n3157), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4833 ( .A1(n3211), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4834 ( .A1(n3273), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4835 ( .A1(n4109), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4836 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3837)
         );
  AOI22_X1 U4837 ( .A1(n3002), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4838 ( .A1(n4147), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4839 ( .A1(n2991), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4840 ( .A1(n3258), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4841 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  OR2_X1 U4842 ( .A1(n3837), .A2(n3836), .ZN(n4214) );
  NAND2_X1 U4843 ( .A1(n4215), .A2(n4214), .ZN(n4252) );
  AOI22_X1 U4844 ( .A1(n3211), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4845 ( .A1(n3273), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4846 ( .A1(n3000), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4847 ( .A1(n2991), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4848 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4849 ( .A1(n3157), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4850 ( .A1(n4147), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4851 ( .A1(n4238), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4852 ( .A1(n3002), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4853 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4854 ( .A1(n3848), .A2(n3847), .ZN(n4253) );
  XOR2_X1 U4855 ( .A(n4252), .B(n4253), .Z(n3849) );
  NAND2_X1 U4856 ( .A1(n3849), .A2(n4203), .ZN(n3854) );
  INV_X2 U4857 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6374) );
  NOR2_X2 U4858 ( .A1(n3304), .A2(n6374), .ZN(n3863) );
  INV_X1 U4859 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4236) );
  AOI21_X1 U4860 ( .B1(n4236), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3850) );
  AOI21_X1 U4861 ( .B1(n4206), .B2(EAX_REG_29__SCAN_IN), .A(n3850), .ZN(n3853)
         );
  NOR2_X2 U4862 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3892) );
  INV_X1 U4863 ( .A(n4207), .ZN(n3852) );
  XNOR2_X1 U4864 ( .A(n4237), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5339)
         );
  NAND2_X1 U4865 ( .A1(n3855), .A2(n4018), .ZN(n3856) );
  NAND2_X1 U4866 ( .A1(n2988), .A2(n4018), .ZN(n3861) );
  AOI22_X1 U4867 ( .A1(n4206), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6374), .ZN(n3859) );
  NAND2_X1 U4868 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3858) );
  AND2_X1 U4869 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  NAND2_X1 U4870 ( .A1(n3861), .A2(n3860), .ZN(n4424) );
  AOI21_X1 U4871 ( .B1(n4314), .B2(n3169), .A(n6374), .ZN(n4438) );
  INV_X1 U4872 ( .A(n3862), .ZN(n6368) );
  NAND2_X1 U4873 ( .A1(n6368), .A2(n4018), .ZN(n3867) );
  AOI22_X1 U4874 ( .A1(n3863), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6374), .ZN(n3865) );
  NAND2_X1 U4875 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3864) );
  AND2_X1 U4876 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  NAND2_X1 U4877 ( .A1(n3867), .A2(n3866), .ZN(n4437) );
  NAND2_X1 U4878 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  INV_X1 U4879 ( .A(n4437), .ZN(n3868) );
  NAND2_X1 U4880 ( .A1(n3868), .A2(n4208), .ZN(n3869) );
  NAND2_X1 U4881 ( .A1(n4436), .A2(n3869), .ZN(n4425) );
  INV_X1 U4882 ( .A(n3881), .ZN(n3878) );
  OAI21_X1 U4883 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3870), .ZN(n6138) );
  AOI22_X1 U4884 ( .A1(n4277), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4208), 
        .B2(n6138), .ZN(n3872) );
  NAND2_X1 U4885 ( .A1(n4206), .A2(EAX_REG_2__SCAN_IN), .ZN(n3871) );
  INV_X1 U4886 ( .A(n4018), .ZN(n4035) );
  OAI21_X1 U4887 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3875), .A(n3874), 
        .ZN(n6128) );
  AOI22_X1 U4888 ( .A1(n3892), .A2(n6128), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3877) );
  NAND2_X1 U4889 ( .A1(n4206), .A2(EAX_REG_3__SCAN_IN), .ZN(n3876) );
  OAI211_X1 U4890 ( .C1(n3878), .C2(n3111), .A(n3877), .B(n3876), .ZN(n3879)
         );
  INV_X1 U4891 ( .A(n3879), .ZN(n3880) );
  INV_X1 U4892 ( .A(n4488), .ZN(n3890) );
  NAND2_X1 U4893 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3886) );
  INV_X1 U4894 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5076) );
  AOI21_X1 U4895 ( .B1(n5076), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3882) );
  AOI21_X1 U4896 ( .B1(n4206), .B2(EAX_REG_4__SCAN_IN), .A(n3882), .ZN(n3885)
         );
  NOR2_X1 U4897 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3883), .ZN(n3884)
         );
  NOR2_X1 U4898 ( .A1(n3896), .A2(n3884), .ZN(n5073) );
  AOI22_X1 U4899 ( .A1(n3886), .A2(n3885), .B1(n3892), .B2(n5073), .ZN(n3887)
         );
  AOI21_X1 U4900 ( .B1(n3888), .B2(n4018), .A(n3887), .ZN(n4516) );
  NAND2_X1 U4901 ( .A1(n3890), .A2(n3889), .ZN(n4515) );
  INV_X1 U4902 ( .A(n4515), .ZN(n3909) );
  NAND2_X1 U4903 ( .A1(n3891), .A2(n4018), .ZN(n3895) );
  INV_X1 U4904 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4997) );
  XNOR2_X1 U4905 ( .A(n3902), .B(n4997), .ZN(n4998) );
  OAI22_X1 U4906 ( .A1(n4998), .A2(n4261), .B1(n3988), .B2(n4997), .ZN(n3893)
         );
  AOI21_X1 U4907 ( .B1(n4206), .B2(EAX_REG_7__SCAN_IN), .A(n3893), .ZN(n3894)
         );
  INV_X1 U4908 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3898) );
  XNOR2_X1 U4909 ( .A(n3896), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U4910 ( .A1(n5062), .A2(n3892), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3897) );
  OAI21_X1 U4911 ( .B1(n3905), .B2(n3898), .A(n3897), .ZN(n3899) );
  AND2_X1 U4912 ( .A1(n3901), .A2(n3904), .ZN(n3903) );
  OR2_X1 U4913 ( .A1(n3903), .A2(n3902), .ZN(n6118) );
  INV_X1 U4914 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4669) );
  OAI22_X1 U4915 ( .A1(n3905), .A2(n4669), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3904), .ZN(n3906) );
  MUX2_X1 U4916 ( .A(n6118), .B(n3906), .S(n4261), .Z(n3907) );
  AOI21_X1 U4917 ( .B1(n3908), .B2(n4018), .A(n3907), .ZN(n4661) );
  NOR2_X1 U4918 ( .A1(n4617), .A2(n4661), .ZN(n4659) );
  NAND3_X1 U4919 ( .A1(n3909), .A2(n4707), .A3(n4659), .ZN(n4672) );
  AOI22_X1 U4920 ( .A1(n5764), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4921 ( .A1(n3258), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4922 ( .A1(n2991), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4923 ( .A1(n4128), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4924 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4925 ( .A1(n4147), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4926 ( .A1(n3204), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4927 ( .A1(n3838), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4928 ( .A1(n3002), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4929 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  OAI21_X1 U4930 ( .B1(n3919), .B2(n3918), .A(n4018), .ZN(n3924) );
  NAND2_X1 U4931 ( .A1(n4206), .A2(EAX_REG_8__SCAN_IN), .ZN(n3923) );
  XNOR2_X1 U4932 ( .A(n3920), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U4933 ( .A1(n4985), .A2(n3892), .ZN(n3922) );
  NAND2_X1 U4934 ( .A1(n4277), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3921)
         );
  XOR2_X1 U4935 ( .A(n6006), .B(n3926), .Z(n5142) );
  INV_X1 U4936 ( .A(n5142), .ZN(n6008) );
  AOI22_X1 U4937 ( .A1(n3004), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4938 ( .A1(n4147), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4939 ( .A1(n3258), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4940 ( .A1(n3002), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4941 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3936)
         );
  AOI22_X1 U4942 ( .A1(n5764), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4943 ( .A1(n3393), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4944 ( .A1(n3180), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4945 ( .A1(n4128), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4946 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3935)
         );
  NOR2_X1 U4947 ( .A1(n3936), .A2(n3935), .ZN(n3939) );
  NAND2_X1 U4948 ( .A1(n4206), .A2(EAX_REG_9__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U4949 ( .A1(n4277), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3937)
         );
  OAI211_X1 U4950 ( .C1(n4035), .C2(n3939), .A(n3938), .B(n3937), .ZN(n3940)
         );
  AOI21_X1 U4951 ( .B1(n6008), .B2(n4208), .A(n3940), .ZN(n4756) );
  INV_X1 U4952 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U4953 ( .A(n3941), .B(n5996), .ZN(n6001) );
  AOI22_X1 U4954 ( .A1(n4206), .A2(EAX_REG_10__SCAN_IN), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4955 ( .A1(n4147), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4956 ( .A1(n3204), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4957 ( .A1(n3002), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4958 ( .A1(n2991), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4959 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3951)
         );
  AOI22_X1 U4960 ( .A1(n5764), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4961 ( .A1(n4128), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4962 ( .A1(n4238), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4963 ( .A1(n3258), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4964 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  OAI21_X1 U4965 ( .B1(n3951), .B2(n3950), .A(n4018), .ZN(n3952) );
  OAI211_X1 U4966 ( .C1(n6001), .C2(n4261), .A(n3953), .B(n3952), .ZN(n4926)
         );
  XOR2_X1 U4967 ( .A(n5983), .B(n3954), .Z(n6108) );
  AOI22_X1 U4968 ( .A1(n5764), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4969 ( .A1(n4128), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4970 ( .A1(n3258), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4971 ( .A1(n3000), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4972 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3964)
         );
  AOI22_X1 U4973 ( .A1(n4147), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4974 ( .A1(n3002), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4975 ( .A1(n3180), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4976 ( .A1(n3353), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4977 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  OR2_X1 U4978 ( .A1(n3964), .A2(n3963), .ZN(n3965) );
  AOI22_X1 U4979 ( .A1(n4018), .A2(n3965), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3967) );
  NAND2_X1 U4980 ( .A1(n4206), .A2(EAX_REG_11__SCAN_IN), .ZN(n3966) );
  OAI211_X1 U4981 ( .C1(n6108), .C2(n4261), .A(n3967), .B(n3966), .ZN(n4990)
         );
  NAND2_X1 U4982 ( .A1(n4924), .A2(n4990), .ZN(n4991) );
  INV_X1 U4983 ( .A(n4991), .ZN(n3984) );
  XNOR2_X1 U4984 ( .A(n3968), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5254)
         );
  INV_X1 U4985 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5054) );
  AOI21_X1 U4986 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5054), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3970) );
  AND2_X1 U4987 ( .A1(n4206), .A2(EAX_REG_12__SCAN_IN), .ZN(n3969) );
  OAI22_X1 U4988 ( .A1(n5254), .A2(n4261), .B1(n3970), .B2(n3969), .ZN(n3982)
         );
  AOI22_X1 U4989 ( .A1(n4245), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4990 ( .A1(n3204), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4991 ( .A1(n3004), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4992 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n2991), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4993 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4994 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4128), .B1(n4147), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4995 ( .A1(n5764), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4996 ( .A1(n4238), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4997 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3258), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4998 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  OAI21_X1 U4999 ( .B1(n3980), .B2(n3979), .A(n4018), .ZN(n3981) );
  INV_X1 U5000 ( .A(n5048), .ZN(n3983) );
  NAND2_X1 U5001 ( .A1(n3984), .A2(n3983), .ZN(n3992) );
  INV_X1 U5002 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3989) );
  OAI21_X1 U5003 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3986), .A(n3985), 
        .ZN(n5975) );
  NAND2_X1 U5004 ( .A1(n5975), .A2(n3892), .ZN(n3987) );
  OAI21_X1 U5005 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n3990) );
  NAND2_X1 U5006 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  AOI22_X1 U5007 ( .A1(n5764), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5008 ( .A1(n4147), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5009 ( .A1(n4128), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5010 ( .A1(n2991), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U5011 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4003)
         );
  AOI22_X1 U5012 ( .A1(n3204), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5013 ( .A1(n4238), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U5014 ( .A1(n3002), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5015 ( .A1(n3838), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U5016 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4002)
         );
  OR2_X1 U5017 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  AND2_X1 U5018 ( .A1(n4018), .A2(n4004), .ZN(n5169) );
  NAND2_X1 U5019 ( .A1(n5168), .A2(n5169), .ZN(n5172) );
  XOR2_X1 U5020 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4006), .Z(n5959) );
  AOI22_X1 U5021 ( .A1(n3004), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5022 ( .A1(n4128), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5023 ( .A1(n3258), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5024 ( .A1(n4245), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U5025 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4016)
         );
  AOI22_X1 U5026 ( .A1(n4147), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5027 ( .A1(n3002), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5028 ( .A1(n2991), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U5029 ( .A1(n5764), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U5030 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  OR2_X1 U5031 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  AOI22_X1 U5032 ( .A1(n4018), .A2(n4017), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U5033 ( .A1(n4206), .A2(EAX_REG_14__SCAN_IN), .ZN(n4019) );
  OAI211_X1 U5034 ( .C1(n5959), .C2(n4261), .A(n4020), .B(n4019), .ZN(n5232)
         );
  XNOR2_X1 U5035 ( .A(n4021), .B(n5271), .ZN(n5607) );
  AOI22_X1 U5036 ( .A1(n4128), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5037 ( .A1(n3204), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5038 ( .A1(n4147), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5039 ( .A1(n4238), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U5040 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4031)
         );
  AOI22_X1 U5041 ( .A1(n5764), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5042 ( .A1(n3002), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5043 ( .A1(n3000), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5044 ( .A1(n2991), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U5045 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4030)
         );
  NOR2_X1 U5046 ( .A1(n4031), .A2(n4030), .ZN(n4034) );
  NAND2_X1 U5047 ( .A1(n4206), .A2(EAX_REG_15__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U5048 ( .A1(n4277), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4032)
         );
  OAI211_X1 U5049 ( .C1(n4035), .C2(n4034), .A(n4033), .B(n4032), .ZN(n4036)
         );
  AOI21_X1 U5050 ( .B1(n5607), .B2(n3892), .A(n4036), .ZN(n5259) );
  XOR2_X1 U5051 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4037), .Z(n5950) );
  AOI22_X1 U5052 ( .A1(n3863), .A2(EAX_REG_16__SCAN_IN), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5053 ( .A1(n4128), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5764), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5054 ( .A1(n4147), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5055 ( .A1(n3258), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5056 ( .A1(n4114), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5057 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U5058 ( .A1(n3004), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5059 ( .A1(n3002), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5060 ( .A1(n3204), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5061 ( .A1(n4245), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5062 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  OAI21_X1 U5063 ( .B1(n4047), .B2(n4046), .A(n4203), .ZN(n4048) );
  OAI211_X1 U5064 ( .C1(n5950), .C2(n4261), .A(n4049), .B(n4048), .ZN(n5482)
         );
  INV_X1 U5065 ( .A(n5397), .ZN(n4069) );
  XNOR2_X1 U5066 ( .A(n4050), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5867)
         );
  NAND2_X1 U5067 ( .A1(n5867), .A2(n3892), .ZN(n4067) );
  AOI22_X1 U5068 ( .A1(n4147), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5069 ( .A1(n4128), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5070 ( .A1(n4114), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5071 ( .A1(n3258), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U5072 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4062)
         );
  AOI22_X1 U5073 ( .A1(n3204), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U5074 ( .A1(n2991), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4056) );
  NAND2_X1 U5075 ( .A1(n5764), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4055)
         );
  AND3_X1 U5076 ( .A1(n4056), .A2(n4055), .A3(n4261), .ZN(n4059) );
  AOI22_X1 U5077 ( .A1(n2990), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5078 ( .A1(n4245), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4057) );
  NAND4_X1 U5079 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4061)
         );
  NAND2_X1 U5080 ( .A1(n4258), .A2(n4261), .ZN(n4139) );
  OAI21_X1 U5081 ( .B1(n4062), .B2(n4061), .A(n4139), .ZN(n4065) );
  NOR2_X1 U5082 ( .A1(n5405), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4063) );
  AOI21_X1 U5083 ( .B1(n4206), .B2(EAX_REG_17__SCAN_IN), .A(n4063), .ZN(n4064)
         );
  NAND2_X1 U5084 ( .A1(n4065), .A2(n4064), .ZN(n4066) );
  NAND2_X1 U5085 ( .A1(n4067), .A2(n4066), .ZN(n5401) );
  AOI22_X1 U5086 ( .A1(n5764), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5087 ( .A1(n4147), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5088 ( .A1(n3258), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5089 ( .A1(n3002), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U5090 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4079)
         );
  AOI22_X1 U5091 ( .A1(n4128), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5092 ( .A1(n3393), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5093 ( .A1(n4109), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5094 ( .A1(n3180), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5095 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4078)
         );
  NOR2_X1 U5096 ( .A1(n4079), .A2(n4078), .ZN(n4083) );
  NAND2_X1 U5097 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4080)
         );
  NAND2_X1 U5098 ( .A1(n4261), .A2(n4080), .ZN(n4081) );
  AOI21_X1 U5099 ( .B1(n3863), .B2(EAX_REG_18__SCAN_IN), .A(n4081), .ZN(n4082)
         );
  OAI21_X1 U5100 ( .B1(n4258), .B2(n4083), .A(n4082), .ZN(n4090) );
  INV_X1 U5101 ( .A(n4106), .ZN(n4088) );
  INV_X1 U5102 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4086) );
  INV_X1 U5103 ( .A(n4084), .ZN(n4085) );
  NAND2_X1 U5104 ( .A1(n4086), .A2(n4085), .ZN(n4087) );
  NAND2_X1 U5105 ( .A1(n4088), .A2(n4087), .ZN(n5942) );
  NAND2_X1 U5106 ( .A1(n4090), .A2(n4089), .ZN(n5470) );
  AOI22_X1 U5107 ( .A1(n5764), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5108 ( .A1(n4238), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5109 ( .A1(n4128), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5110 ( .A1(n3002), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4092) );
  NAND4_X1 U5111 ( .A1(n4095), .A2(n4094), .A3(n4093), .A4(n4092), .ZN(n4103)
         );
  AOI22_X1 U5112 ( .A1(n3004), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5113 ( .A1(n4147), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U5114 ( .A1(n2991), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U5115 ( .A1(n2990), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4096)
         );
  AND3_X1 U5116 ( .A1(n4097), .A2(n4096), .A3(n4261), .ZN(n4099) );
  AOI22_X1 U5117 ( .A1(n4109), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4098) );
  NAND4_X1 U5118 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(n4102)
         );
  OAI21_X1 U5119 ( .B1(n4103), .B2(n4102), .A(n4139), .ZN(n4105) );
  AOI22_X1 U5120 ( .A1(n3863), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6374), .ZN(n4104) );
  NAND2_X1 U5121 ( .A1(n4105), .A2(n4104), .ZN(n4108) );
  INV_X1 U5122 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5834) );
  XNOR2_X1 U5123 ( .A(n4106), .B(n5834), .ZN(n5839) );
  NAND2_X1 U5124 ( .A1(n5839), .A2(n3892), .ZN(n4107) );
  NAND2_X1 U5125 ( .A1(n4108), .A2(n4107), .ZN(n5459) );
  AOI22_X1 U5126 ( .A1(n5764), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5127 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4147), .B1(n4109), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5128 ( .A1(n2990), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5129 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3002), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U5130 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4120)
         );
  AOI22_X1 U5131 ( .A1(n4128), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5132 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3258), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5133 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n2991), .B1(n4114), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5134 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3273), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U5135 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4119)
         );
  NOR2_X1 U5136 ( .A1(n4120), .A2(n4119), .ZN(n4124) );
  NAND2_X1 U5137 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4121)
         );
  NAND2_X1 U5138 ( .A1(n4261), .A2(n4121), .ZN(n4122) );
  AOI21_X1 U5139 ( .B1(n3863), .B2(EAX_REG_20__SCAN_IN), .A(n4122), .ZN(n4123)
         );
  OAI21_X1 U5140 ( .B1(n4258), .B2(n4124), .A(n4123), .ZN(n4127) );
  OAI21_X1 U5141 ( .B1(n4125), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4144), 
        .ZN(n5825) );
  OR2_X1 U5142 ( .A1(n5825), .A2(n4261), .ZN(n4126) );
  AOI22_X1 U5143 ( .A1(n3003), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5144 ( .A1(n4128), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5145 ( .A1(n4238), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5146 ( .A1(n4244), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U5147 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4141)
         );
  AOI22_X1 U5148 ( .A1(n2990), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5149 ( .A1(n4147), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5150 ( .A1(n3002), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U5151 ( .A1(n5764), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4134)
         );
  NAND2_X1 U5152 ( .A1(n3180), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4133) );
  AND3_X1 U5153 ( .A1(n4134), .A2(n4261), .A3(n4133), .ZN(n4135) );
  NAND4_X1 U5154 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4140)
         );
  OAI21_X1 U5155 ( .B1(n4141), .B2(n4140), .A(n4139), .ZN(n4143) );
  AOI22_X1 U5156 ( .A1(n3863), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6374), .ZN(n4142) );
  NAND2_X1 U5157 ( .A1(n4143), .A2(n4142), .ZN(n4146) );
  XNOR2_X1 U5158 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4144), .ZN(n5817)
         );
  NAND2_X1 U5159 ( .A1(n5817), .A2(n3892), .ZN(n4145) );
  NAND2_X1 U5160 ( .A1(n4146), .A2(n4145), .ZN(n5446) );
  AOI22_X1 U5161 ( .A1(n5764), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5162 ( .A1(n3353), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5163 ( .A1(n4147), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5164 ( .A1(n4245), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U5165 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4157)
         );
  AOI22_X1 U5166 ( .A1(n3002), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5167 ( .A1(n4238), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5168 ( .A1(n3180), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5169 ( .A1(n4128), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5170 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  NOR2_X1 U5171 ( .A1(n4157), .A2(n4156), .ZN(n4161) );
  NAND2_X1 U5172 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4158)
         );
  NAND2_X1 U5173 ( .A1(n4261), .A2(n4158), .ZN(n4159) );
  AOI21_X1 U5174 ( .B1(n3863), .B2(EAX_REG_22__SCAN_IN), .A(n4159), .ZN(n4160)
         );
  OAI21_X1 U5175 ( .B1(n4258), .B2(n4161), .A(n4160), .ZN(n4164) );
  OAI21_X1 U5176 ( .B1(n4162), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4169), 
        .ZN(n5804) );
  OR2_X1 U5177 ( .A1(n5804), .A2(n4261), .ZN(n4163) );
  NAND2_X1 U5178 ( .A1(n4164), .A2(n4163), .ZN(n5439) );
  XOR2_X1 U5179 ( .A(n4166), .B(n4165), .Z(n4167) );
  NAND2_X1 U5180 ( .A1(n4167), .A2(n4203), .ZN(n4172) );
  OAI21_X1 U5181 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5567), .A(n4261), .ZN(
        n4168) );
  AOI21_X1 U5182 ( .B1(n3863), .B2(EAX_REG_23__SCAN_IN), .A(n4168), .ZN(n4171)
         );
  XNOR2_X1 U5183 ( .A(n4169), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5571)
         );
  AOI21_X1 U5184 ( .B1(n4172), .B2(n4171), .A(n4170), .ZN(n5387) );
  XNOR2_X1 U5185 ( .A(n4174), .B(n4173), .ZN(n4179) );
  NOR2_X1 U5186 ( .A1(n4175), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4176)
         );
  OR2_X1 U5187 ( .A1(n4188), .A2(n4176), .ZN(n5795) );
  AOI22_X1 U5188 ( .A1(n5795), .A2(n4208), .B1(PHYADDRPOINTER_REG_24__SCAN_IN), 
        .B2(n4277), .ZN(n4178) );
  NAND2_X1 U5189 ( .A1(n3863), .A2(EAX_REG_24__SCAN_IN), .ZN(n4177) );
  OAI211_X1 U5190 ( .C1(n4179), .C2(n4258), .A(n4178), .B(n4177), .ZN(n5429)
         );
  NAND2_X1 U5191 ( .A1(n5385), .A2(n5429), .ZN(n5420) );
  INV_X1 U5192 ( .A(n5420), .ZN(n4192) );
  XOR2_X1 U5193 ( .A(n4181), .B(n4180), .Z(n4182) );
  NAND2_X1 U5194 ( .A1(n4182), .A2(n4203), .ZN(n4186) );
  NAND2_X1 U5195 ( .A1(n6374), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4183)
         );
  NAND2_X1 U5196 ( .A1(n4261), .A2(n4183), .ZN(n4184) );
  AOI21_X1 U5197 ( .B1(n3863), .B2(EAX_REG_25__SCAN_IN), .A(n4184), .ZN(n4185)
         );
  NAND2_X1 U5198 ( .A1(n4186), .A2(n4185), .ZN(n4190) );
  INV_X1 U5199 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4187) );
  XNOR2_X1 U5200 ( .A(n4188), .B(n4187), .ZN(n5785) );
  NAND2_X1 U5201 ( .A1(n5785), .A2(n4208), .ZN(n4189) );
  NAND2_X1 U5202 ( .A1(n4190), .A2(n4189), .ZN(n5422) );
  OR2_X1 U5203 ( .A1(n4193), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4194)
         );
  NAND2_X1 U5204 ( .A1(n4207), .A2(n4194), .ZN(n5538) );
  XNOR2_X1 U5205 ( .A(n4196), .B(n4195), .ZN(n4199) );
  AOI21_X1 U5206 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6374), .A(n4208), 
        .ZN(n4198) );
  NAND2_X1 U5207 ( .A1(n3863), .A2(EAX_REG_26__SCAN_IN), .ZN(n4197) );
  OAI211_X1 U5208 ( .C1(n4199), .C2(n4258), .A(n4198), .B(n4197), .ZN(n4200)
         );
  OAI21_X1 U5209 ( .B1(n4261), .B2(n5538), .A(n4200), .ZN(n5375) );
  XOR2_X1 U5210 ( .A(n4202), .B(n4201), .Z(n4204) );
  NAND2_X1 U5211 ( .A1(n4204), .A2(n4203), .ZN(n4210) );
  INV_X1 U5212 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5530) );
  NOR2_X1 U5213 ( .A1(n5530), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4205) );
  AOI211_X1 U5214 ( .C1(n4206), .C2(EAX_REG_27__SCAN_IN), .A(n3892), .B(n4205), 
        .ZN(n4209) );
  XNOR2_X1 U5215 ( .A(n4207), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5534)
         );
  INV_X1 U5216 ( .A(n4211), .ZN(n4212) );
  INV_X1 U5217 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U5218 ( .A1(n4212), .A2(n5352), .ZN(n4213) );
  NAND2_X1 U5219 ( .A1(n4237), .A2(n4213), .ZN(n5523) );
  XNOR2_X1 U5220 ( .A(n4215), .B(n4214), .ZN(n4218) );
  AOI21_X1 U5221 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6374), .A(n3892), 
        .ZN(n4217) );
  NAND2_X1 U5222 ( .A1(n3863), .A2(EAX_REG_28__SCAN_IN), .ZN(n4216) );
  OAI211_X1 U5223 ( .C1(n4218), .C2(n4258), .A(n4217), .B(n4216), .ZN(n4219)
         );
  OAI21_X1 U5224 ( .B1(n4261), .B2(n5523), .A(n4219), .ZN(n5348) );
  NAND2_X1 U5225 ( .A1(n4221), .A2(n4220), .ZN(n4262) );
  NAND3_X1 U5226 ( .A1(n6466), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6484) );
  INV_X1 U5227 ( .A(n6484), .ZN(n4223) );
  NOR2_X2 U5228 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6365) );
  INV_X1 U5229 ( .A(n5508), .ZN(n4227) );
  INV_X1 U5230 ( .A(n4224), .ZN(n4226) );
  NAND2_X1 U5231 ( .A1(n4226), .A2(n4225), .ZN(n5510) );
  NAND2_X1 U5232 ( .A1(n4227), .A2(n5510), .ZN(n4228) );
  NAND2_X1 U5233 ( .A1(n6371), .A2(n4229), .ZN(n6570) );
  NAND2_X1 U5234 ( .A1(n6570), .A2(n6466), .ZN(n4230) );
  NAND2_X1 U5235 ( .A1(n6466), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4232) );
  NAND2_X1 U5236 ( .A1(n6758), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4231) );
  AND2_X1 U5237 ( .A1(n4232), .A2(n4231), .ZN(n4435) );
  INV_X1 U5238 ( .A(n4435), .ZN(n4233) );
  NAND2_X1 U5239 ( .A1(n6213), .A2(REIP_REG_29__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U5240 ( .B1(n5616), .B2(n4236), .A(n5631), .ZN(n4234) );
  AOI21_X1 U5241 ( .B1(n6109), .B2(n5339), .A(n4234), .ZN(n4235) );
  INV_X1 U5242 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5331) );
  XNOR2_X1 U5243 ( .A(n4284), .B(n5331), .ZN(n5513) );
  AOI22_X1 U5244 ( .A1(n3157), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5245 ( .A1(n3266), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5246 ( .A1(n4238), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5247 ( .A1(n2991), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4239) );
  NAND4_X1 U5248 ( .A1(n4242), .A2(n4241), .A3(n4240), .A4(n4239), .ZN(n4251)
         );
  AOI22_X1 U5249 ( .A1(n4128), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U5250 ( .A1(n3002), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U5251 ( .A1(n3000), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4243), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U5252 ( .A1(n4245), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4246) );
  NAND4_X1 U5253 ( .A1(n4249), .A2(n4248), .A3(n4247), .A4(n4246), .ZN(n4250)
         );
  NOR2_X1 U5254 ( .A1(n4251), .A2(n4250), .ZN(n4255) );
  NOR2_X1 U5255 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  XOR2_X1 U5256 ( .A(n4255), .B(n4254), .Z(n4259) );
  AOI21_X1 U5257 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6374), .A(n3892), 
        .ZN(n4257) );
  NAND2_X1 U5258 ( .A1(n3863), .A2(EAX_REG_30__SCAN_IN), .ZN(n4256) );
  OAI211_X1 U5259 ( .C1(n4259), .C2(n4258), .A(n4257), .B(n4256), .ZN(n4260)
         );
  OAI21_X1 U5260 ( .B1(n4261), .B2(n5513), .A(n4260), .ZN(n4263) );
  NOR2_X2 U5261 ( .A1(n4262), .A2(n4263), .ZN(n4279) );
  AOI21_X1 U5262 ( .B1(n4262), .B2(n4263), .A(n4279), .ZN(n5515) );
  INV_X1 U5263 ( .A(n5515), .ZN(n5416) );
  INV_X1 U5264 ( .A(n4264), .ZN(n4265) );
  OAI22_X1 U5265 ( .A1(n5314), .A2(n5311), .B1(n2993), .B2(n4265), .ZN(n4376)
         );
  INV_X1 U5266 ( .A(n3304), .ZN(n5488) );
  NAND3_X1 U5267 ( .A1(n5488), .A2(n3227), .A3(n2992), .ZN(n4266) );
  OR2_X1 U5268 ( .A1(n4405), .A2(n4266), .ZN(n4427) );
  NOR2_X1 U5269 ( .A1(n4427), .A2(n4267), .ZN(n4268) );
  OAI21_X1 U5270 ( .B1(n4376), .B2(n4268), .A(n4431), .ZN(n4271) );
  AND2_X1 U5271 ( .A1(n4273), .A2(n4272), .ZN(n4444) );
  AND2_X1 U5272 ( .A1(n5489), .A2(n3305), .ZN(n6062) );
  AOI22_X1 U5273 ( .A1(n6062), .A2(DATAI_30_), .B1(n6065), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4276) );
  INV_X1 U5274 ( .A(n4272), .ZN(n4274) );
  NAND2_X1 U5275 ( .A1(n6066), .A2(DATAI_14_), .ZN(n4275) );
  OAI21_X1 U5276 ( .B1(n5416), .B2(n5843), .A(n3110), .ZN(U2861) );
  AOI22_X1 U5277 ( .A1(n3863), .A2(EAX_REG_31__SCAN_IN), .B1(n4277), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4278) );
  XNOR2_X1 U5278 ( .A(n4279), .B(n4278), .ZN(n5491) );
  NOR2_X1 U5279 ( .A1(n5312), .A2(n4281), .ZN(n5318) );
  NAND2_X1 U5280 ( .A1(n5318), .A2(n4431), .ZN(n4364) );
  NOR2_X1 U5281 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6574) );
  INV_X1 U5282 ( .A(n6574), .ZN(n6483) );
  NOR3_X1 U5283 ( .A1(n6466), .A2(n6560), .A3(n6483), .ZN(n6467) );
  NOR3_X1 U5284 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6476), .A3(n6465), .ZN(
        n6479) );
  OR2_X1 U5285 ( .A1(n6199), .A2(n6479), .ZN(n4282) );
  NOR2_X1 U5286 ( .A1(n6467), .A2(n4282), .ZN(n4283) );
  INV_X1 U5287 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U5288 ( .A1(n5491), .A2(n6026), .ZN(n4305) );
  INV_X1 U5289 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5413) );
  INV_X1 U5290 ( .A(READY_N), .ZN(n4287) );
  NAND2_X1 U5291 ( .A1(n6758), .A2(n4287), .ZN(n4822) );
  NAND2_X1 U5292 ( .A1(n3638), .A2(n4822), .ZN(n4288) );
  INV_X1 U5293 ( .A(n4822), .ZN(n4294) );
  NAND3_X1 U5294 ( .A1(n4289), .A2(n4294), .A3(n3244), .ZN(n4290) );
  INV_X1 U5295 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U5296 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4292) );
  NAND3_X1 U5297 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4291) );
  INV_X1 U5298 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6531) );
  INV_X1 U5299 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6528) );
  INV_X1 U5300 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6517) );
  INV_X1 U5301 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6515) );
  INV_X1 U5302 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6511) );
  NAND3_X1 U5303 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5074) );
  NOR2_X1 U5304 ( .A1(n6511), .A2(n5074), .ZN(n5060) );
  NAND2_X1 U5305 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5060), .ZN(n4999) );
  NOR2_X1 U5306 ( .A1(n6515), .A2(n4999), .ZN(n5001) );
  NAND2_X1 U5307 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5001), .ZN(n4982) );
  NOR2_X1 U5308 ( .A1(n6517), .A2(n4982), .ZN(n4983) );
  NAND4_X1 U5309 ( .A1(REIP_REG_11__SCAN_IN), .A2(n4983), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5310 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5968) );
  NOR2_X1 U5311 ( .A1(n5049), .A2(n5968), .ZN(n5957) );
  NAND2_X1 U5312 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5957), .ZN(n5265) );
  NOR3_X1 U5313 ( .A1(n6531), .A2(n6528), .A3(n5265), .ZN(n4297) );
  AND3_X1 U5314 ( .A1(n5269), .A2(REIP_REG_17__SCAN_IN), .A3(n4297), .ZN(n5402) );
  NAND4_X1 U5315 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5402), .ZN(n5803) );
  NOR2_X1 U5316 ( .A1(n4291), .A2(n5803), .ZN(n5389) );
  AND3_X1 U5317 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U5318 ( .A1(n5267), .A2(n5269), .ZN(n5992) );
  INV_X1 U5319 ( .A(n5992), .ZN(n5403) );
  AOI21_X1 U5320 ( .B1(n5389), .B2(n5367), .A(n5403), .ZN(n5373) );
  AOI21_X1 U5321 ( .B1(n5061), .B2(n4292), .A(n5373), .ZN(n4293) );
  INV_X1 U5322 ( .A(n4293), .ZN(n5354) );
  AOI21_X1 U5323 ( .B1(n5061), .B2(n6549), .A(n5354), .ZN(n5334) );
  OAI21_X1 U5324 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5267), .A(n5334), .ZN(n4301) );
  INV_X1 U5325 ( .A(n6495), .ZN(n4739) );
  NAND2_X1 U5326 ( .A1(n4739), .A2(n4294), .ZN(n6461) );
  NAND2_X1 U5327 ( .A1(n3238), .A2(n6461), .ZN(n4824) );
  OAI22_X1 U5328 ( .A1(n6005), .A2(n4296), .B1(n4295), .B2(n4824), .ZN(n4300)
         );
  INV_X1 U5329 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6703) );
  INV_X1 U5330 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U5331 ( .A1(n5061), .A2(n4297), .ZN(n5404) );
  NAND3_X1 U5332 ( .A1(n5935), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5824) );
  NAND4_X1 U5333 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5811), .ZN(n5788) );
  NAND2_X1 U5334 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5367), .ZN(n4298) );
  NOR2_X1 U5335 ( .A1(n5788), .A2(n4298), .ZN(n5358) );
  NAND2_X1 U5336 ( .A1(n5358), .A2(REIP_REG_28__SCAN_IN), .ZN(n5346) );
  INV_X1 U5337 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6587) );
  NOR4_X1 U5338 ( .A1(n5346), .A2(REIP_REG_31__SCAN_IN), .A3(n6587), .A4(n6549), .ZN(n4299) );
  AOI211_X1 U5339 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4301), .A(n4300), .B(n4299), .ZN(n4302) );
  NAND2_X1 U5340 ( .A1(n4305), .A2(n4304), .ZN(U2796) );
  NAND2_X1 U5341 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4306)
         );
  OAI211_X1 U5342 ( .C1(n6139), .C2(n4831), .A(n4307), .B(n4306), .ZN(n4308)
         );
  AOI21_X1 U5343 ( .B1(n5491), .B2(n6133), .A(n4308), .ZN(n4311) );
  NAND2_X1 U5344 ( .A1(n4311), .A2(n4310), .ZN(U2955) );
  OAI21_X1 U5345 ( .B1(n6277), .B2(n6313), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4320) );
  INV_X1 U5346 ( .A(n4319), .ZN(n4561) );
  NAND2_X1 U5347 ( .A1(n4317), .A2(n4561), .ZN(n5093) );
  OR2_X1 U5348 ( .A1(n4315), .A2(n5093), .ZN(n6285) );
  NAND3_X1 U5349 ( .A1(n4320), .A2(n6365), .A3(n6285), .ZN(n4322) );
  NOR2_X1 U5350 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6290), .ZN(n6276)
         );
  INV_X1 U5351 ( .A(n6276), .ZN(n4345) );
  NOR2_X1 U5352 ( .A1(n4325), .A2(n6374), .ZN(n5087) );
  NAND2_X1 U5353 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4741) );
  OAI21_X1 U5354 ( .B1(n5180), .B2(n6374), .A(n4765), .ZN(n5088) );
  AOI211_X1 U5355 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4345), .A(n5087), .B(
        n5088), .ZN(n4321) );
  NAND3_X1 U5356 ( .A1(n6446), .A2(n4322), .A3(n4321), .ZN(n6278) );
  INV_X1 U5357 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4323) );
  NOR2_X1 U5358 ( .A1(n4736), .A2(n4323), .ZN(n4330) );
  NAND2_X1 U5359 ( .A1(n6133), .A2(DATAI_28_), .ZN(n6347) );
  NOR2_X1 U5360 ( .A1(n4629), .A2(n6347), .ZN(n4329) );
  NAND2_X1 U5361 ( .A1(n6133), .A2(DATAI_20_), .ZN(n6405) );
  NOR2_X1 U5362 ( .A1(n6311), .A2(n6405), .ZN(n4328) );
  NAND2_X1 U5363 ( .A1(n6466), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U5364 ( .A1(n4574), .A2(n3240), .ZN(n5203) );
  AND2_X1 U5365 ( .A1(n4325), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5182) );
  NAND3_X1 U5366 ( .A1(n5182), .A2(n5180), .A3(n6446), .ZN(n4326) );
  OAI21_X1 U5367 ( .B1(n6285), .B2(n6371), .A(n4326), .ZN(n6275) );
  INV_X1 U5368 ( .A(n6275), .ZN(n4344) );
  INV_X1 U5369 ( .A(DATAI_4_), .ZN(n6719) );
  INV_X1 U5370 ( .A(n6402), .ZN(n5122) );
  OAI22_X1 U5371 ( .A1(n5203), .A2(n4345), .B1(n4344), .B2(n5122), .ZN(n4327)
         );
  OR4_X1 U5372 ( .A1(n4330), .A2(n4329), .A3(n4328), .A4(n4327), .ZN(U3072) );
  INV_X1 U5373 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4331) );
  NOR2_X1 U5374 ( .A1(n4736), .A2(n4331), .ZN(n4335) );
  NAND2_X1 U5375 ( .A1(n6133), .A2(DATAI_26_), .ZN(n6393) );
  NOR2_X1 U5376 ( .A1(n4629), .A2(n6393), .ZN(n4334) );
  NAND2_X1 U5377 ( .A1(n6133), .A2(DATAI_18_), .ZN(n6301) );
  NOR2_X1 U5378 ( .A1(n6311), .A2(n6301), .ZN(n4333) );
  NAND2_X1 U5379 ( .A1(n4574), .A2(n3192), .ZN(n5219) );
  INV_X1 U5380 ( .A(DATAI_2_), .ZN(n6683) );
  INV_X1 U5381 ( .A(n6390), .ZN(n5128) );
  OAI22_X1 U5382 ( .A1(n5219), .A2(n4345), .B1(n4344), .B2(n5128), .ZN(n4332)
         );
  OR4_X1 U5383 ( .A1(n4335), .A2(n4334), .A3(n4333), .A4(n4332), .ZN(U3070) );
  INV_X1 U5384 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4336) );
  NOR2_X1 U5385 ( .A1(n4736), .A2(n4336), .ZN(n4341) );
  NAND2_X1 U5386 ( .A1(n6133), .A2(DATAI_29_), .ZN(n6411) );
  NOR2_X1 U5387 ( .A1(n4629), .A2(n6411), .ZN(n4340) );
  NAND2_X1 U5388 ( .A1(n6133), .A2(DATAI_21_), .ZN(n6263) );
  NOR2_X1 U5389 ( .A1(n6311), .A2(n6263), .ZN(n4339) );
  NAND2_X1 U5390 ( .A1(n4574), .A2(n4337), .ZN(n5207) );
  INV_X1 U5391 ( .A(DATAI_5_), .ZN(n4634) );
  INV_X1 U5392 ( .A(n6408), .ZN(n5100) );
  OAI22_X1 U5393 ( .A1(n5207), .A2(n4345), .B1(n4344), .B2(n5100), .ZN(n4338)
         );
  OR4_X1 U5394 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(U3073) );
  INV_X1 U5395 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4342) );
  NOR2_X1 U5396 ( .A1(n4736), .A2(n4342), .ZN(n4349) );
  NAND2_X1 U5397 ( .A1(n6133), .A2(DATAI_27_), .ZN(n6399) );
  NOR2_X1 U5398 ( .A1(n4629), .A2(n6399), .ZN(n4348) );
  NAND2_X1 U5399 ( .A1(n6133), .A2(DATAI_19_), .ZN(n6257) );
  NOR2_X1 U5400 ( .A1(n6311), .A2(n6257), .ZN(n4347) );
  NAND2_X1 U5401 ( .A1(n4574), .A2(n4343), .ZN(n5215) );
  INV_X1 U5402 ( .A(DATAI_3_), .ZN(n6738) );
  INV_X1 U5403 ( .A(n6396), .ZN(n5110) );
  OAI22_X1 U5404 ( .A1(n5215), .A2(n4345), .B1(n4344), .B2(n5110), .ZN(n4346)
         );
  OR4_X1 U5405 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(U3071) );
  NAND3_X1 U5406 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6446), .A3(n4844), .ZN(n6245) );
  NOR2_X1 U5407 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6245), .ZN(n4357)
         );
  AND2_X1 U5408 ( .A1(n3873), .A2(n4511), .ZN(n4350) );
  AND2_X1 U5409 ( .A1(n3873), .A2(n4840), .ZN(n4352) );
  NAND2_X1 U5410 ( .A1(n4352), .A2(n6237), .ZN(n6267) );
  NAND2_X1 U5411 ( .A1(n6365), .A2(n6758), .ZN(n6328) );
  OAI21_X1 U5412 ( .B1(n4586), .B2(n6268), .A(n6328), .ZN(n4353) );
  NOR2_X1 U5413 ( .A1(n4317), .A2(n4319), .ZN(n4842) );
  NAND2_X1 U5414 ( .A1(n6322), .A2(n4842), .ZN(n6240) );
  NAND2_X1 U5415 ( .A1(n4353), .A2(n6240), .ZN(n4354) );
  NOR2_X1 U5416 ( .A1(n5182), .A2(n5088), .ZN(n4848) );
  INV_X1 U5417 ( .A(n4958), .ZN(n4356) );
  INV_X1 U5418 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4355) );
  NOR2_X1 U5419 ( .A1(n4356), .A2(n4355), .ZN(n4363) );
  NAND2_X1 U5420 ( .A1(n6133), .A2(DATAI_24_), .ZN(n6381) );
  NOR2_X1 U5421 ( .A1(n4964), .A2(n6381), .ZN(n4362) );
  NAND2_X1 U5422 ( .A1(n6133), .A2(DATAI_16_), .ZN(n6295) );
  NOR2_X1 U5423 ( .A1(n6267), .A2(n6295), .ZN(n4361) );
  NAND2_X1 U5424 ( .A1(n4574), .A2(n3244), .ZN(n5199) );
  INV_X1 U5425 ( .A(n4357), .ZN(n4960) );
  OR2_X1 U5426 ( .A1(n6240), .A2(n6371), .ZN(n4359) );
  NAND3_X1 U5427 ( .A1(n5087), .A2(n5180), .A3(n6446), .ZN(n4358) );
  INV_X1 U5428 ( .A(DATAI_0_), .ZN(n6760) );
  NOR2_X2 U5429 ( .A1(n6760), .A2(n5188), .ZN(n6378) );
  INV_X1 U5430 ( .A(n6378), .ZN(n5096) );
  OAI22_X1 U5431 ( .A1(n5199), .A2(n4960), .B1(n4959), .B2(n5096), .ZN(n4360)
         );
  OR4_X1 U5432 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(U3036) );
  INV_X1 U5433 ( .A(n4364), .ZN(n4365) );
  INV_X1 U5434 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6579) );
  NAND2_X1 U5435 ( .A1(n6365), .A2(n6465), .ZN(n5917) );
  OAI211_X1 U5436 ( .C1(n4365), .C2(n6579), .A(n4386), .B(n5917), .ZN(U2788)
         );
  INV_X1 U5437 ( .A(n4267), .ZN(n5319) );
  NOR2_X1 U5438 ( .A1(n5319), .A2(n3638), .ZN(n5321) );
  INV_X1 U5439 ( .A(n5917), .ZN(n4980) );
  OAI21_X1 U5440 ( .B1(n4980), .B2(READREQUEST_REG_SCAN_IN), .A(n4367), .ZN(
        n4366) );
  OAI21_X1 U5441 ( .B1(n4367), .B2(n5321), .A(n4366), .ZN(U3474) );
  NAND2_X1 U5442 ( .A1(n5314), .A2(n5315), .ZN(n4430) );
  INV_X1 U5443 ( .A(n4430), .ZN(n4375) );
  AOI21_X1 U5444 ( .B1(n4368), .B2(n6495), .A(READY_N), .ZN(n4369) );
  OAI21_X1 U5445 ( .B1(n5769), .B2(n3611), .A(n4369), .ZN(n4373) );
  INV_X1 U5446 ( .A(n4370), .ZN(n4372) );
  OAI211_X1 U5447 ( .C1(n5314), .C2(n4373), .A(n4372), .B(n4371), .ZN(n4374)
         );
  INV_X1 U5448 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6594) );
  OR2_X1 U5449 ( .A1(n6466), .A2(n4741), .ZN(n6557) );
  OAI22_X1 U5450 ( .A1(n6443), .A2(n6477), .B1(n6594), .B2(n6557), .ZN(n4381)
         );
  INV_X1 U5451 ( .A(n4381), .ZN(n4377) );
  NAND2_X1 U5452 ( .A1(n6558), .A2(n4377), .ZN(n5782) );
  INV_X1 U5453 ( .A(n4596), .ZN(n4378) );
  NOR2_X1 U5454 ( .A1(n4379), .A2(n4378), .ZN(n4380) );
  XNOR2_X1 U5455 ( .A(n4380), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5077)
         );
  INV_X1 U5456 ( .A(n2993), .ZN(n4382) );
  NAND3_X1 U5457 ( .A1(n4382), .A2(n5777), .A3(n4381), .ZN(n4383) );
  OAI22_X1 U5458 ( .A1(n5782), .A2(n4384), .B1(n5077), .B2(n4383), .ZN(U3455)
         );
  INV_X1 U5459 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U5460 ( .A1(n4473), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U5461 ( .A1(n4459), .A2(DATAI_11_), .ZN(n4465) );
  OAI211_X1 U5462 ( .C1(n6079), .C2(n4446), .A(n4387), .B(n4465), .ZN(U2950)
         );
  INV_X1 U5463 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U5464 ( .A1(n4473), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5465 ( .A1(n4459), .A2(DATAI_12_), .ZN(n4463) );
  OAI211_X1 U5466 ( .C1(n6077), .C2(n4446), .A(n4388), .B(n4463), .ZN(U2951)
         );
  INV_X1 U5467 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U5468 ( .A1(n4473), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U5469 ( .A1(n4459), .A2(DATAI_9_), .ZN(n4396) );
  OAI211_X1 U5470 ( .C1(n4753), .C2(n4446), .A(n4389), .B(n4396), .ZN(U2933)
         );
  INV_X1 U5471 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U5472 ( .A1(n4473), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5473 ( .A1(n4459), .A2(DATAI_10_), .ZN(n4393) );
  OAI211_X1 U5474 ( .C1(n6081), .C2(n4446), .A(n4390), .B(n4393), .ZN(U2949)
         );
  NAND2_X1 U5475 ( .A1(n4473), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5476 ( .A1(n4459), .A2(DATAI_6_), .ZN(n4400) );
  OAI211_X1 U5477 ( .C1(n4669), .C2(n4446), .A(n4391), .B(n4400), .ZN(U2945)
         );
  NAND2_X1 U5478 ( .A1(n4473), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U5479 ( .A1(n4459), .A2(DATAI_5_), .ZN(n4454) );
  OAI211_X1 U5480 ( .C1(n3898), .C2(n4446), .A(n4392), .B(n4454), .ZN(U2944)
         );
  INV_X1 U5481 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U5482 ( .A1(n4473), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4394) );
  OAI211_X1 U5483 ( .C1(n4747), .C2(n4446), .A(n4394), .B(n4393), .ZN(U2934)
         );
  INV_X1 U5484 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U5485 ( .A1(n4473), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5486 ( .A1(n4459), .A2(DATAI_8_), .ZN(n4398) );
  OAI211_X1 U5487 ( .C1(n4755), .C2(n4446), .A(n4395), .B(n4398), .ZN(U2932)
         );
  INV_X1 U5488 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U5489 ( .A1(n4473), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U5490 ( .C1(n6083), .C2(n4446), .A(n4397), .B(n4396), .ZN(U2948)
         );
  INV_X1 U5491 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5492 ( .A1(n4473), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4399) );
  OAI211_X1 U5493 ( .C1(n6085), .C2(n4446), .A(n4399), .B(n4398), .ZN(U2947)
         );
  INV_X1 U5494 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U5495 ( .A1(n4473), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4401) );
  OAI211_X1 U5496 ( .C1(n5158), .C2(n4446), .A(n4401), .B(n4400), .ZN(U2930)
         );
  INV_X1 U5497 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U5498 ( .A1(n4473), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U5499 ( .A1(n4459), .A2(DATAI_14_), .ZN(n4449) );
  OAI211_X1 U5500 ( .C1(n6073), .C2(n4446), .A(n4402), .B(n4449), .ZN(U2953)
         );
  INV_X1 U5501 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U5502 ( .A1(n4473), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U5503 ( .A1(n4459), .A2(DATAI_13_), .ZN(n4447) );
  OAI211_X1 U5504 ( .C1(n6075), .C2(n4446), .A(n4403), .B(n4447), .ZN(U2952)
         );
  INV_X1 U5505 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U5506 ( .A1(n4473), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5507 ( .A1(n4459), .A2(DATAI_7_), .ZN(n4457) );
  OAI211_X1 U5508 ( .C1(n5161), .C2(n4446), .A(n4404), .B(n4457), .ZN(U2931)
         );
  INV_X1 U5509 ( .A(n3611), .ZN(n6462) );
  AND4_X1 U5510 ( .A1(n3245), .A2(n2993), .A3(n6462), .A4(n4405), .ZN(n4406)
         );
  NAND2_X1 U5511 ( .A1(n4407), .A2(n4406), .ZN(n5758) );
  INV_X1 U5512 ( .A(n5758), .ZN(n5297) );
  NOR3_X1 U5513 ( .A1(n5296), .A2(n4408), .A3(n4409), .ZN(n4410) );
  AOI21_X1 U5514 ( .B1(n5769), .B2(n3112), .A(n4410), .ZN(n4411) );
  OAI21_X1 U5515 ( .B1(n4319), .B2(n5297), .A(n4411), .ZN(n6434) );
  INV_X1 U5516 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5288) );
  NOR2_X1 U5517 ( .A1(n6465), .A2(n5288), .ZN(n4414) );
  AOI22_X1 U5518 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4412), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6234), .ZN(n5287) );
  INV_X1 U5519 ( .A(n4409), .ZN(n4413) );
  INV_X1 U5520 ( .A(n6470), .ZN(n5778) );
  NOR2_X1 U5521 ( .A1(n5778), .A2(n4408), .ZN(n5293) );
  AOI222_X1 U5522 ( .A1(n6434), .A2(n5777), .B1(n4414), .B2(n5287), .C1(n4413), 
        .C2(n5293), .ZN(n4416) );
  NAND2_X1 U5523 ( .A1(n5299), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4415) );
  OAI21_X1 U5524 ( .B1(n5299), .B2(n4416), .A(n4415), .ZN(U3460) );
  XNOR2_X1 U5525 ( .A(n4417), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4443)
         );
  NAND2_X1 U5526 ( .A1(n5743), .A2(n5717), .ZN(n5740) );
  NAND2_X1 U5527 ( .A1(n5288), .A2(n5740), .ZN(n6232) );
  OR2_X1 U5528 ( .A1(n4418), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4420)
         );
  AND2_X1 U5529 ( .A1(n4420), .A2(n4419), .ZN(n4487) );
  AND2_X1 U5530 ( .A1(n6199), .A2(REIP_REG_0__SCAN_IN), .ZN(n4440) );
  AOI21_X1 U5531 ( .B1(n6233), .B2(n5906), .A(n5288), .ZN(n4421) );
  AOI211_X1 U5532 ( .C1(n6223), .C2(n4487), .A(n4440), .B(n4421), .ZN(n4422)
         );
  OAI211_X1 U5533 ( .C1(n4443), .C2(n6201), .A(n6232), .B(n4422), .ZN(U3018)
         );
  NOR2_X1 U5534 ( .A1(n4424), .A2(n4425), .ZN(n4426) );
  NOR2_X1 U5535 ( .A1(n4423), .A2(n4426), .ZN(n4500) );
  INV_X1 U5536 ( .A(n4500), .ZN(n4839) );
  INV_X1 U5537 ( .A(n4427), .ZN(n4428) );
  NAND2_X1 U5538 ( .A1(n4428), .A2(n3638), .ZN(n4429) );
  NAND2_X1 U5539 ( .A1(n4430), .A2(n4429), .ZN(n4432) );
  OAI21_X1 U5540 ( .B1(n4830), .B2(n3638), .A(n4433), .ZN(n6222) );
  AOI22_X1 U5541 ( .A1(n6051), .A2(n6222), .B1(n5479), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4434) );
  OAI21_X1 U5542 ( .B1(n4839), .B2(n5469), .A(n4434), .ZN(U2858) );
  NAND2_X1 U5543 ( .A1(n4435), .A2(n5616), .ZN(n4441) );
  OAI21_X1 U5544 ( .B1(n4438), .B2(n4437), .A(n4436), .ZN(n4979) );
  NOR2_X1 U5545 ( .A1(n4979), .A2(n6122), .ZN(n4439) );
  AOI211_X1 U5546 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4441), .A(n4440), 
        .B(n4439), .ZN(n4442) );
  OAI21_X1 U5547 ( .B1(n4443), .B2(n6124), .A(n4442), .ZN(U2986) );
  INV_X1 U5548 ( .A(n4444), .ZN(n4445) );
  INV_X1 U5549 ( .A(DATAI_1_), .ZN(n4573) );
  INV_X1 U5550 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6098) );
  OAI222_X1 U5551 ( .A1(n4839), .A2(n5843), .B1(n4668), .B2(n4573), .C1(n5489), 
        .C2(n6098), .ZN(U2890) );
  INV_X1 U5552 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5553 ( .A1(n4473), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4448) );
  OAI211_X1 U5554 ( .C1(n4749), .C2(n4446), .A(n4448), .B(n4447), .ZN(U2937)
         );
  INV_X1 U5555 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5556 ( .A1(n4473), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4450) );
  OAI211_X1 U5557 ( .C1(n4743), .C2(n4446), .A(n4450), .B(n4449), .ZN(U2938)
         );
  INV_X1 U5558 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5559 ( .A1(n4473), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4451) );
  NAND2_X1 U5560 ( .A1(n4459), .A2(DATAI_2_), .ZN(n4474) );
  OAI211_X1 U5561 ( .C1(n5152), .C2(n4446), .A(n4451), .B(n4474), .ZN(U2926)
         );
  INV_X1 U5562 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U5563 ( .A1(n4473), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5564 ( .A1(n4459), .A2(DATAI_3_), .ZN(n4467) );
  OAI211_X1 U5565 ( .C1(n5154), .C2(n4446), .A(n4452), .B(n4467), .ZN(U2927)
         );
  INV_X1 U5566 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U5567 ( .A1(n4473), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5568 ( .A1(n4459), .A2(DATAI_4_), .ZN(n4469) );
  OAI211_X1 U5569 ( .C1(n5156), .C2(n4446), .A(n4453), .B(n4469), .ZN(U2928)
         );
  INV_X1 U5570 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U5571 ( .A1(n4473), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4455) );
  OAI211_X1 U5572 ( .C1(n5150), .C2(n4446), .A(n4455), .B(n4454), .ZN(U2929)
         );
  INV_X1 U5573 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U5574 ( .A1(n4473), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U5575 ( .A1(n4459), .A2(DATAI_0_), .ZN(n4461) );
  OAI211_X1 U5576 ( .C1(n5146), .C2(n4446), .A(n4456), .B(n4461), .ZN(U2924)
         );
  INV_X1 U5577 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U5578 ( .A1(n4473), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4458) );
  OAI211_X1 U5579 ( .C1(n6087), .C2(n4446), .A(n4458), .B(n4457), .ZN(U2946)
         );
  NAND2_X1 U5580 ( .A1(n4473), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5581 ( .A1(n4459), .A2(DATAI_1_), .ZN(n4471) );
  OAI211_X1 U5582 ( .C1(n6098), .C2(n4446), .A(n4460), .B(n4471), .ZN(U2940)
         );
  INV_X1 U5583 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5584 ( .A1(n4473), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4462) );
  OAI211_X1 U5585 ( .C1(n6103), .C2(n4446), .A(n4462), .B(n4461), .ZN(U2939)
         );
  INV_X1 U5586 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5587 ( .A1(n4473), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4464) );
  OAI211_X1 U5588 ( .C1(n4751), .C2(n4446), .A(n4464), .B(n4463), .ZN(U2936)
         );
  INV_X1 U5589 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U5590 ( .A1(n4473), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4466) );
  OAI211_X1 U5591 ( .C1(n4745), .C2(n4446), .A(n4466), .B(n4465), .ZN(U2935)
         );
  INV_X1 U5592 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U5593 ( .A1(n4473), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4468) );
  OAI211_X1 U5594 ( .C1(n6094), .C2(n4446), .A(n4468), .B(n4467), .ZN(U2942)
         );
  INV_X1 U5595 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U5596 ( .A1(n4473), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4470) );
  OAI211_X1 U5597 ( .C1(n6092), .C2(n4446), .A(n4470), .B(n4469), .ZN(U2943)
         );
  INV_X1 U5598 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U5599 ( .A1(n4473), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4472) );
  OAI211_X1 U5600 ( .C1(n5148), .C2(n4446), .A(n4472), .B(n4471), .ZN(U2925)
         );
  INV_X1 U5601 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U5602 ( .A1(n4473), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4475) );
  OAI211_X1 U5603 ( .C1(n6096), .C2(n4446), .A(n4475), .B(n4474), .ZN(U2941)
         );
  INV_X1 U5604 ( .A(DATAI_15_), .ZN(n4479) );
  INV_X1 U5605 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4477) );
  INV_X1 U5606 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6071) );
  OAI222_X1 U5607 ( .A1(n4479), .A2(n4478), .B1(n4477), .B2(n4476), .C1(n4446), 
        .C2(n6071), .ZN(U2954) );
  NOR2_X1 U5608 ( .A1(n4481), .A2(n4482), .ZN(n4483) );
  NOR2_X1 U5609 ( .A1(n4480), .A2(n4483), .ZN(n6134) );
  INV_X1 U5610 ( .A(n6134), .ZN(n4486) );
  XNOR2_X1 U5611 ( .A(n4484), .B(n4492), .ZN(n6212) );
  AOI22_X1 U5612 ( .A1(n6051), .A2(n6212), .B1(n5479), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4485) );
  OAI21_X1 U5613 ( .B1(n4486), .B2(n5469), .A(n4485), .ZN(U2857) );
  OAI222_X1 U5614 ( .A1(n4486), .A2(n5843), .B1(n4668), .B2(n6683), .C1(n5489), 
        .C2(n6096), .ZN(U2889) );
  INV_X1 U5615 ( .A(n4487), .ZN(n4974) );
  OAI222_X1 U5616 ( .A1(n4979), .A2(n5487), .B1(n4972), .B2(n6055), .C1(n6045), 
        .C2(n4974), .ZN(U2859) );
  OR2_X1 U5617 ( .A1(n4480), .A2(n4489), .ZN(n4490) );
  NAND2_X1 U5618 ( .A1(n4488), .A2(n4490), .ZN(n6123) );
  INV_X1 U5619 ( .A(n4484), .ZN(n4493) );
  AOI21_X1 U5620 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(n4494) );
  NOR2_X1 U5621 ( .A1(n4494), .A2(n3032), .ZN(n6200) );
  AOI22_X1 U5622 ( .A1(n6051), .A2(n6200), .B1(n5479), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4495) );
  OAI21_X1 U5623 ( .B1(n6123), .B2(n5469), .A(n4495), .ZN(U2856) );
  XOR2_X1 U5624 ( .A(n4497), .B(n4496), .Z(n6230) );
  INV_X1 U5625 ( .A(n6230), .ZN(n4502) );
  NAND2_X1 U5626 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4498)
         );
  NAND2_X1 U5627 ( .A1(n6213), .A2(REIP_REG_1__SCAN_IN), .ZN(n6224) );
  OAI211_X1 U5628 ( .C1(n6139), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4498), 
        .B(n6224), .ZN(n4499) );
  AOI21_X1 U5629 ( .B1(n4500), .B2(n6133), .A(n4499), .ZN(n4501) );
  OAI21_X1 U5630 ( .B1(n4502), .B2(n6124), .A(n4501), .ZN(U2985) );
  OAI222_X1 U5631 ( .A1(n4979), .A2(n5843), .B1(n4668), .B2(n6760), .C1(n5489), 
        .C2(n6103), .ZN(U2891) );
  OAI222_X1 U5632 ( .A1(n6123), .A2(n5843), .B1(n4668), .B2(n6738), .C1(n5489), 
        .C2(n6094), .ZN(U2888) );
  NAND2_X1 U5633 ( .A1(n4503), .A2(n6594), .ZN(n4504) );
  NOR2_X1 U5634 ( .A1(n4504), .A2(n4409), .ZN(n4509) );
  OR2_X1 U5635 ( .A1(n2993), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4505) );
  OR2_X1 U5636 ( .A1(n5077), .A2(n4505), .ZN(n4508) );
  MUX2_X1 U5637 ( .A(n6443), .B(n6594), .S(STATE2_REG_1__SCAN_IN), .Z(n4506)
         );
  NAND2_X1 U5638 ( .A1(n4506), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5639 ( .A1(n4508), .A2(n4507), .ZN(n6458) );
  NOR2_X1 U5640 ( .A1(n4509), .A2(n6458), .ZN(n4589) );
  AOI21_X1 U5641 ( .B1(n4589), .B2(n6594), .A(n6557), .ZN(n4510) );
  NOR2_X1 U5642 ( .A1(n4510), .A2(n4765), .ZN(n6235) );
  XNOR2_X1 U5643 ( .A(n6364), .B(n6237), .ZN(n4512) );
  NAND2_X1 U5644 ( .A1(n6560), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5645 ( .A1(n4512), .A2(n6365), .B1(n4591), .B2(n4317), .ZN(n4514)
         );
  NAND2_X1 U5646 ( .A1(n6235), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4513) );
  OAI21_X1 U5647 ( .B1(n6235), .B2(n4514), .A(n4513), .ZN(U3463) );
  AOI21_X1 U5648 ( .B1(n4516), .B2(n4488), .A(n3909), .ZN(n4530) );
  AND2_X1 U5649 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  OR2_X1 U5650 ( .A1(n4519), .A2(n4553), .ZN(n6192) );
  OAI22_X1 U5651 ( .A1(n6045), .A2(n6192), .B1(n4520), .B2(n6055), .ZN(n4521)
         );
  AOI21_X1 U5652 ( .B1(n4530), .B2(n6052), .A(n4521), .ZN(n4522) );
  INV_X1 U5653 ( .A(n4522), .ZN(U2855) );
  OR2_X1 U5654 ( .A1(n4524), .A2(n4523), .ZN(n4525) );
  NAND2_X1 U5655 ( .A1(n2995), .A2(n4525), .ZN(n6190) );
  NAND2_X1 U5656 ( .A1(n4530), .A2(n6133), .ZN(n4529) );
  OAI22_X1 U5657 ( .A1(n5616), .A2(n5076), .B1(n6191), .B2(n6511), .ZN(n4527)
         );
  AOI21_X1 U5658 ( .B1(n6109), .B2(n5073), .A(n4527), .ZN(n4528) );
  OAI211_X1 U5659 ( .C1(n6190), .C2(n6124), .A(n4529), .B(n4528), .ZN(U2982)
         );
  INV_X1 U5660 ( .A(n4530), .ZN(n5085) );
  OAI222_X1 U5661 ( .A1(n5085), .A2(n5843), .B1(n4668), .B2(n6719), .C1(n5489), 
        .C2(n6092), .ZN(U2887) );
  INV_X1 U5662 ( .A(DATAI_7_), .ZN(n6776) );
  NOR2_X2 U5663 ( .A1(n6776), .A2(n5188), .ZN(n6425) );
  INV_X1 U5664 ( .A(n6425), .ZN(n5194) );
  AND2_X1 U5665 ( .A1(n4315), .A2(n6368), .ZN(n4887) );
  NAND2_X1 U5666 ( .A1(n4317), .A2(n4319), .ZN(n5178) );
  INV_X1 U5667 ( .A(n5178), .ZN(n4531) );
  NAND2_X1 U5668 ( .A1(n6437), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4597) );
  NOR2_X1 U5669 ( .A1(n6446), .A2(n4597), .ZN(n5183) );
  AND2_X1 U5670 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5183), .ZN(n4630)
         );
  AOI21_X1 U5671 ( .B1(n4887), .B2(n4531), .A(n4630), .ZN(n4534) );
  NAND2_X1 U5672 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4532) );
  OAI22_X1 U5673 ( .A1(n4534), .A2(n6371), .B1(n4532), .B2(n4597), .ZN(n4654)
         );
  INV_X1 U5674 ( .A(n4654), .ZN(n4541) );
  NAND2_X1 U5675 ( .A1(n4574), .A2(n3304), .ZN(n5105) );
  NOR2_X1 U5676 ( .A1(n2988), .A2(n4313), .ZN(n4533) );
  NAND2_X1 U5677 ( .A1(n4538), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5754) );
  NAND2_X1 U5678 ( .A1(n4534), .A2(n5754), .ZN(n4537) );
  AOI21_X1 U5679 ( .B1(n5184), .B2(STATE2_REG_3__SCAN_IN), .A(n5188), .ZN(
        n4562) );
  INV_X1 U5680 ( .A(n5183), .ZN(n4535) );
  NAND2_X1 U5681 ( .A1(n6371), .A2(n4535), .ZN(n4536) );
  OAI211_X1 U5682 ( .C1(n6371), .C2(n4537), .A(n4562), .B(n4536), .ZN(n4653)
         );
  AOI22_X1 U5683 ( .A1(n6421), .A2(n4630), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4653), .ZN(n4540) );
  NAND2_X1 U5684 ( .A1(n6133), .A2(DATAI_31_), .ZN(n6430) );
  INV_X1 U5685 ( .A(n6430), .ZN(n6312) );
  NAND2_X1 U5686 ( .A1(n6133), .A2(DATAI_23_), .ZN(n6319) );
  INV_X1 U5687 ( .A(n6319), .ZN(n6423) );
  AOI22_X1 U5688 ( .A1(n6312), .A2(n5228), .B1(n5089), .B2(n6423), .ZN(n4539)
         );
  OAI211_X1 U5689 ( .C1(n5194), .C2(n4541), .A(n4540), .B(n4539), .ZN(U3131)
         );
  OAI21_X1 U5690 ( .B1(n4542), .B2(n4544), .A(n4543), .ZN(n4622) );
  NAND2_X1 U5691 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4545), .ZN(n6220)
         );
  NOR2_X1 U5692 ( .A1(n6211), .A2(n6220), .ZN(n4716) );
  NAND3_X1 U5693 ( .A1(n6189), .A2(n4716), .A3(n4550), .ZN(n4558) );
  NAND2_X1 U5694 ( .A1(n6189), .A2(n6209), .ZN(n4551) );
  NOR2_X1 U5695 ( .A1(n6211), .A2(n6234), .ZN(n4547) );
  INV_X1 U5696 ( .A(n6153), .ZN(n4546) );
  OAI21_X1 U5697 ( .B1(n4548), .B2(n4547), .A(n4546), .ZN(n6217) );
  AOI221_X1 U5698 ( .B1(n4550), .B2(n6221), .C1(n4551), .C2(n6221), .A(n6217), 
        .ZN(n4549) );
  INV_X1 U5699 ( .A(n4549), .ZN(n4719) );
  OAI21_X1 U5700 ( .B1(n5717), .B2(n4551), .A(n4550), .ZN(n4556) );
  OR2_X1 U5701 ( .A1(n4553), .A2(n4552), .ZN(n4554) );
  AND2_X1 U5702 ( .A1(n4663), .A2(n4554), .ZN(n5065) );
  INV_X1 U5703 ( .A(n5065), .ZN(n4635) );
  INV_X1 U5704 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6513) );
  OAI22_X1 U5705 ( .A1(n4635), .A2(n6193), .B1(n6513), .B2(n6191), .ZN(n4555)
         );
  AOI21_X1 U5706 ( .B1(n4719), .B2(n4556), .A(n4555), .ZN(n4557) );
  OAI211_X1 U5707 ( .C1(n4622), .C2(n6201), .A(n4558), .B(n4557), .ZN(U3013)
         );
  INV_X1 U5708 ( .A(n4559), .ZN(n4560) );
  OAI21_X1 U5709 ( .B1(n4560), .B2(n6758), .A(n6365), .ZN(n4565) );
  NOR2_X1 U5710 ( .A1(n4315), .A2(n6321), .ZN(n4768) );
  NAND3_X1 U5711 ( .A1(n6446), .A2(n4844), .A3(n6437), .ZN(n4763) );
  NOR2_X1 U5712 ( .A1(n5184), .A2(n4763), .ZN(n4585) );
  AOI21_X1 U5713 ( .B1(n4768), .B2(n6368), .A(n4585), .ZN(n4566) );
  INV_X1 U5714 ( .A(n4566), .ZN(n4564) );
  AOI21_X1 U5715 ( .B1(n6371), .B2(n4763), .A(n6370), .ZN(n4563) );
  OAI21_X1 U5716 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n4584) );
  OAI22_X1 U5717 ( .A1(n4566), .A2(n4565), .B1(n6374), .B2(n4763), .ZN(n4583)
         );
  AOI22_X1 U5718 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4584), .B1(n6402), 
        .B2(n4583), .ZN(n4568) );
  INV_X1 U5719 ( .A(n6405), .ZN(n6344) );
  AOI22_X1 U5720 ( .A1(n4586), .A2(n6344), .B1(n6400), .B2(n4585), .ZN(n4567)
         );
  OAI211_X1 U5721 ( .C1(n6347), .C2(n4820), .A(n4568), .B(n4567), .ZN(U3032)
         );
  NAND2_X1 U5722 ( .A1(n6133), .A2(DATAI_30_), .ZN(n6353) );
  AOI22_X1 U5723 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4584), .B1(n6415), 
        .B2(n4583), .ZN(n4570) );
  NAND2_X1 U5724 ( .A1(n6133), .A2(DATAI_22_), .ZN(n6419) );
  INV_X1 U5725 ( .A(n6419), .ZN(n6350) );
  NAND2_X1 U5726 ( .A1(n4574), .A2(n2992), .ZN(n5211) );
  AOI22_X1 U5727 ( .A1(n4586), .A2(n6350), .B1(n6412), .B2(n4585), .ZN(n4569)
         );
  OAI211_X1 U5728 ( .C1(n6353), .C2(n4820), .A(n4570), .B(n4569), .ZN(U3034)
         );
  AOI22_X1 U5729 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4584), .B1(n6425), 
        .B2(n4583), .ZN(n4572) );
  AOI22_X1 U5730 ( .A1(n4586), .A2(n6423), .B1(n6421), .B2(n4585), .ZN(n4571)
         );
  OAI211_X1 U5731 ( .C1(n6430), .C2(n4820), .A(n4572), .B(n4571), .ZN(U3035)
         );
  NAND2_X1 U5732 ( .A1(n6133), .A2(DATAI_25_), .ZN(n6339) );
  NOR2_X2 U5733 ( .A1(n4573), .A2(n5188), .ZN(n6384) );
  AOI22_X1 U5734 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4584), .B1(n6384), 
        .B2(n4583), .ZN(n4576) );
  NAND2_X1 U5735 ( .A1(n6133), .A2(DATAI_17_), .ZN(n6387) );
  INV_X1 U5736 ( .A(n6387), .ZN(n6336) );
  NAND2_X1 U5737 ( .A1(n4574), .A2(n3236), .ZN(n5226) );
  AOI22_X1 U5738 ( .A1(n4586), .A2(n6336), .B1(n6382), .B2(n4585), .ZN(n4575)
         );
  OAI211_X1 U5739 ( .C1(n6339), .C2(n4820), .A(n4576), .B(n4575), .ZN(U3029)
         );
  AOI22_X1 U5740 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4584), .B1(n6378), 
        .B2(n4583), .ZN(n4578) );
  INV_X1 U5741 ( .A(n6295), .ZN(n6363) );
  AOI22_X1 U5742 ( .A1(n4586), .A2(n6363), .B1(n6362), .B2(n4585), .ZN(n4577)
         );
  OAI211_X1 U5743 ( .C1(n6381), .C2(n4820), .A(n4578), .B(n4577), .ZN(U3028)
         );
  AOI22_X1 U5744 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4584), .B1(n6390), 
        .B2(n4583), .ZN(n4580) );
  INV_X1 U5745 ( .A(n6301), .ZN(n6389) );
  AOI22_X1 U5746 ( .A1(n4586), .A2(n6389), .B1(n6388), .B2(n4585), .ZN(n4579)
         );
  OAI211_X1 U5747 ( .C1(n6393), .C2(n4820), .A(n4580), .B(n4579), .ZN(U3030)
         );
  AOI22_X1 U5748 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4584), .B1(n6396), 
        .B2(n4583), .ZN(n4582) );
  INV_X1 U5749 ( .A(n6257), .ZN(n6395) );
  AOI22_X1 U5750 ( .A1(n4586), .A2(n6395), .B1(n6394), .B2(n4585), .ZN(n4581)
         );
  OAI211_X1 U5751 ( .C1(n6399), .C2(n4820), .A(n4582), .B(n4581), .ZN(U3031)
         );
  AOI22_X1 U5752 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4584), .B1(n6408), 
        .B2(n4583), .ZN(n4588) );
  INV_X1 U5753 ( .A(n6263), .ZN(n6407) );
  AOI22_X1 U5754 ( .A1(n4586), .A2(n6407), .B1(n6406), .B2(n4585), .ZN(n4587)
         );
  OAI211_X1 U5755 ( .C1(n6411), .C2(n4820), .A(n4588), .B(n4587), .ZN(U3033)
         );
  INV_X1 U5756 ( .A(n6235), .ZN(n4594) );
  INV_X1 U5757 ( .A(n4589), .ZN(n4590) );
  NOR2_X1 U5758 ( .A1(n4590), .A2(n4741), .ZN(n6468) );
  INV_X1 U5759 ( .A(n4591), .ZN(n5756) );
  OAI22_X1 U5760 ( .A1(n4314), .A2(n6371), .B1(n3862), .B2(n5756), .ZN(n4592)
         );
  OAI21_X1 U5761 ( .B1(n6468), .B2(n4592), .A(n4594), .ZN(n4593) );
  OAI21_X1 U5762 ( .B1(n4594), .B2(n5184), .A(n4593), .ZN(U3465) );
  OR3_X1 U5763 ( .A1(n6282), .A2(n2988), .A3(n6758), .ZN(n4595) );
  NAND2_X1 U5764 ( .A1(n4595), .A2(n6365), .ZN(n4601) );
  NOR2_X1 U5765 ( .A1(n5178), .A2(n4596), .ZN(n5015) );
  OR2_X1 U5766 ( .A1(n4597), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5011)
         );
  NOR2_X1 U5767 ( .A1(n5184), .A2(n5011), .ZN(n4625) );
  AOI21_X1 U5768 ( .B1(n5015), .B2(n6368), .A(n4625), .ZN(n4598) );
  OAI22_X1 U5769 ( .A1(n4601), .A2(n4598), .B1(n5011), .B2(n6374), .ZN(n4624)
         );
  INV_X1 U5770 ( .A(n4598), .ZN(n4600) );
  AOI21_X1 U5771 ( .B1(n6371), .B2(n5011), .A(n6370), .ZN(n4599) );
  OAI21_X1 U5772 ( .B1(n4601), .B2(n4600), .A(n4599), .ZN(n4623) );
  AOI22_X1 U5773 ( .A1(n6408), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4604) );
  INV_X1 U5774 ( .A(n6411), .ZN(n6260) );
  AOI22_X1 U5775 ( .A1(n6260), .A2(n4626), .B1(n6406), .B2(n4625), .ZN(n4603)
         );
  OAI211_X1 U5776 ( .C1(n6263), .C2(n4629), .A(n4604), .B(n4603), .ZN(U3065)
         );
  AOI22_X1 U5777 ( .A1(n6402), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4606) );
  INV_X1 U5778 ( .A(n6347), .ZN(n6401) );
  AOI22_X1 U5779 ( .A1(n6401), .A2(n4626), .B1(n6400), .B2(n4625), .ZN(n4605)
         );
  OAI211_X1 U5780 ( .C1(n6405), .C2(n4629), .A(n4606), .B(n4605), .ZN(U3064)
         );
  AOI22_X1 U5781 ( .A1(n6396), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4608) );
  INV_X1 U5782 ( .A(n6399), .ZN(n6254) );
  AOI22_X1 U5783 ( .A1(n6254), .A2(n4626), .B1(n6394), .B2(n4625), .ZN(n4607)
         );
  OAI211_X1 U5784 ( .C1(n6257), .C2(n4629), .A(n4608), .B(n4607), .ZN(U3063)
         );
  AOI22_X1 U5785 ( .A1(n6390), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4610) );
  INV_X1 U5786 ( .A(n6393), .ZN(n6298) );
  AOI22_X1 U5787 ( .A1(n6298), .A2(n4626), .B1(n6388), .B2(n4625), .ZN(n4609)
         );
  OAI211_X1 U5788 ( .C1(n6301), .C2(n4629), .A(n4610), .B(n4609), .ZN(U3062)
         );
  AOI22_X1 U5789 ( .A1(n6384), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4612) );
  INV_X1 U5790 ( .A(n6339), .ZN(n6383) );
  AOI22_X1 U5791 ( .A1(n6383), .A2(n4626), .B1(n6382), .B2(n4625), .ZN(n4611)
         );
  OAI211_X1 U5792 ( .C1(n6387), .C2(n4629), .A(n4612), .B(n4611), .ZN(U3061)
         );
  AOI22_X1 U5793 ( .A1(n6378), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4614) );
  INV_X1 U5794 ( .A(n6381), .ZN(n6284) );
  AOI22_X1 U5795 ( .A1(n6284), .A2(n4626), .B1(n6362), .B2(n4625), .ZN(n4613)
         );
  OAI211_X1 U5796 ( .C1(n6295), .C2(n4629), .A(n4614), .B(n4613), .ZN(U3060)
         );
  AOI22_X1 U5797 ( .A1(n6415), .A2(n4624), .B1(n4623), .B2(
        INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4616) );
  INV_X1 U5798 ( .A(n6353), .ZN(n6413) );
  AOI22_X1 U5799 ( .A1(n6413), .A2(n4626), .B1(n6412), .B2(n4625), .ZN(n4615)
         );
  OAI211_X1 U5800 ( .C1(n6419), .C2(n4629), .A(n4616), .B(n4615), .ZN(U3066)
         );
  OR2_X1 U5801 ( .A1(n4515), .A2(n4617), .ZN(n4660) );
  INV_X1 U5802 ( .A(n4660), .ZN(n4618) );
  AOI21_X1 U5803 ( .B1(n4617), .B2(n4515), .A(n4618), .ZN(n5071) );
  AOI22_X1 U5804 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6199), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4619) );
  OAI21_X1 U5805 ( .B1(n5062), .B2(n6139), .A(n4619), .ZN(n4620) );
  AOI21_X1 U5806 ( .B1(n5071), .B2(n6133), .A(n4620), .ZN(n4621) );
  OAI21_X1 U5807 ( .B1(n6124), .B2(n4622), .A(n4621), .ZN(U2981) );
  AOI22_X1 U5808 ( .A1(n6425), .A2(n4624), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n4623), .ZN(n4628) );
  AOI22_X1 U5809 ( .A1(n6312), .A2(n4626), .B1(n6421), .B2(n4625), .ZN(n4627)
         );
  OAI211_X1 U5810 ( .C1(n6319), .C2(n4629), .A(n4628), .B(n4627), .ZN(U3067)
         );
  INV_X1 U5811 ( .A(n4630), .ZN(n4656) );
  AOI22_X1 U5812 ( .A1(n4654), .A2(n6402), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4653), .ZN(n4631) );
  OAI21_X1 U5813 ( .B1(n5203), .B2(n4656), .A(n4631), .ZN(n4632) );
  AOI21_X1 U5814 ( .B1(n6401), .B2(n5228), .A(n4632), .ZN(n4633) );
  OAI21_X1 U5815 ( .B1(n6405), .B2(n5134), .A(n4633), .ZN(U3128) );
  INV_X1 U5816 ( .A(n5071), .ZN(n4637) );
  OAI222_X1 U5817 ( .A1(n4637), .A2(n5843), .B1(n4668), .B2(n4634), .C1(n5489), 
        .C2(n3898), .ZN(U2886) );
  INV_X1 U5818 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4636) );
  OAI222_X1 U5819 ( .A1(n4637), .A2(n5487), .B1(n4636), .B2(n6055), .C1(n6045), 
        .C2(n4635), .ZN(U2854) );
  AOI22_X1 U5820 ( .A1(n6415), .A2(n4654), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4653), .ZN(n4638) );
  OAI21_X1 U5821 ( .B1(n5211), .B2(n4656), .A(n4638), .ZN(n4639) );
  AOI21_X1 U5822 ( .B1(n6413), .B2(n5228), .A(n4639), .ZN(n4640) );
  OAI21_X1 U5823 ( .B1(n6419), .B2(n5134), .A(n4640), .ZN(U3130) );
  AOI22_X1 U5824 ( .A1(n4654), .A2(n6378), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4653), .ZN(n4641) );
  OAI21_X1 U5825 ( .B1(n5199), .B2(n4656), .A(n4641), .ZN(n4642) );
  AOI21_X1 U5826 ( .B1(n6284), .B2(n5228), .A(n4642), .ZN(n4643) );
  OAI21_X1 U5827 ( .B1(n6295), .B2(n5134), .A(n4643), .ZN(U3124) );
  AOI22_X1 U5828 ( .A1(n4654), .A2(n6384), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4653), .ZN(n4644) );
  OAI21_X1 U5829 ( .B1(n5226), .B2(n4656), .A(n4644), .ZN(n4645) );
  AOI21_X1 U5830 ( .B1(n6383), .B2(n5228), .A(n4645), .ZN(n4646) );
  OAI21_X1 U5831 ( .B1(n6387), .B2(n5134), .A(n4646), .ZN(U3125) );
  AOI22_X1 U5832 ( .A1(n4654), .A2(n6408), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4653), .ZN(n4647) );
  OAI21_X1 U5833 ( .B1(n5207), .B2(n4656), .A(n4647), .ZN(n4648) );
  AOI21_X1 U5834 ( .B1(n6260), .B2(n5228), .A(n4648), .ZN(n4649) );
  OAI21_X1 U5835 ( .B1(n6263), .B2(n5134), .A(n4649), .ZN(U3129) );
  AOI22_X1 U5836 ( .A1(n4654), .A2(n6396), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4653), .ZN(n4650) );
  OAI21_X1 U5837 ( .B1(n5215), .B2(n4656), .A(n4650), .ZN(n4651) );
  AOI21_X1 U5838 ( .B1(n6254), .B2(n5228), .A(n4651), .ZN(n4652) );
  OAI21_X1 U5839 ( .B1(n6257), .B2(n5134), .A(n4652), .ZN(U3127) );
  AOI22_X1 U5840 ( .A1(n4654), .A2(n6390), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4653), .ZN(n4655) );
  OAI21_X1 U5841 ( .B1(n5219), .B2(n4656), .A(n4655), .ZN(n4657) );
  AOI21_X1 U5842 ( .B1(n6298), .B2(n5228), .A(n4657), .ZN(n4658) );
  OAI21_X1 U5843 ( .B1(n6301), .B2(n5134), .A(n4658), .ZN(U3126) );
  AND2_X1 U5844 ( .A1(n3909), .A2(n4659), .ZN(n4706) );
  AOI21_X1 U5845 ( .B1(n4661), .B2(n4660), .A(n4706), .ZN(n6114) );
  INV_X1 U5846 ( .A(n6114), .ZN(n4670) );
  NAND2_X1 U5847 ( .A1(n4663), .A2(n4662), .ZN(n4664) );
  NAND2_X1 U5848 ( .A1(n4709), .A2(n4664), .ZN(n6023) );
  INV_X1 U5849 ( .A(n6023), .ZN(n4665) );
  AOI22_X1 U5850 ( .A1(n4665), .A2(n6051), .B1(EBX_REG_6__SCAN_IN), .B2(n5479), 
        .ZN(n4666) );
  OAI21_X1 U5851 ( .B1(n4670), .B2(n5469), .A(n4666), .ZN(U2853) );
  INV_X1 U5852 ( .A(DATAI_6_), .ZN(n4667) );
  OAI222_X1 U5853 ( .A1(n4670), .A2(n5843), .B1(n5489), .B2(n4669), .C1(n4668), 
        .C2(n4667), .ZN(U2885) );
  NAND2_X1 U5854 ( .A1(n4672), .A2(n4673), .ZN(n4674) );
  AND2_X1 U5855 ( .A1(n4671), .A2(n4674), .ZN(n4988) );
  INV_X1 U5856 ( .A(n4988), .ZN(n4698) );
  AOI22_X1 U5857 ( .A1(n5279), .A2(DATAI_8_), .B1(n6065), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4675) );
  OAI21_X1 U5858 ( .B1(n4698), .B2(n5843), .A(n4675), .ZN(U2883) );
  INV_X1 U5859 ( .A(n6321), .ZN(n4676) );
  NAND3_X1 U5860 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4844), .A3(n6437), .ZN(n6320) );
  NOR2_X1 U5861 ( .A1(n5184), .A2(n6320), .ZN(n4703) );
  AOI21_X1 U5862 ( .B1(n4887), .B2(n4676), .A(n4703), .ZN(n4681) );
  INV_X1 U5863 ( .A(n4681), .ZN(n4679) );
  OAI21_X1 U5864 ( .B1(n4682), .B2(n6758), .A(n6365), .ZN(n4680) );
  AOI21_X1 U5865 ( .B1(n6371), .B2(n6320), .A(n6370), .ZN(n4678) );
  OAI21_X1 U5866 ( .B1(n4679), .B2(n4680), .A(n4678), .ZN(n4702) );
  OAI22_X1 U5867 ( .A1(n4681), .A2(n4680), .B1(n6374), .B2(n6320), .ZN(n4701)
         );
  AOI22_X1 U5868 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4702), .B1(n6415), 
        .B2(n4701), .ZN(n4684) );
  AOI22_X1 U5869 ( .A1(n6356), .A2(n6413), .B1(n6412), .B2(n4703), .ZN(n4683)
         );
  OAI211_X1 U5870 ( .C1(n4849), .C2(n6419), .A(n4684), .B(n4683), .ZN(U3098)
         );
  AOI22_X1 U5871 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4702), .B1(n6425), 
        .B2(n4701), .ZN(n4686) );
  AOI22_X1 U5872 ( .A1(n6356), .A2(n6312), .B1(n6421), .B2(n4703), .ZN(n4685)
         );
  OAI211_X1 U5873 ( .C1(n4849), .C2(n6319), .A(n4686), .B(n4685), .ZN(U3099)
         );
  AOI22_X1 U5874 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4702), .B1(n6408), 
        .B2(n4701), .ZN(n4688) );
  AOI22_X1 U5875 ( .A1(n6356), .A2(n6260), .B1(n6406), .B2(n4703), .ZN(n4687)
         );
  OAI211_X1 U5876 ( .C1(n4849), .C2(n6263), .A(n4688), .B(n4687), .ZN(U3097)
         );
  AOI22_X1 U5877 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4702), .B1(n6396), 
        .B2(n4701), .ZN(n4690) );
  AOI22_X1 U5878 ( .A1(n6356), .A2(n6254), .B1(n6394), .B2(n4703), .ZN(n4689)
         );
  OAI211_X1 U5879 ( .C1(n4849), .C2(n6257), .A(n4690), .B(n4689), .ZN(U3095)
         );
  AOI22_X1 U5880 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4702), .B1(n6402), 
        .B2(n4701), .ZN(n4692) );
  AOI22_X1 U5881 ( .A1(n6356), .A2(n6401), .B1(n6400), .B2(n4703), .ZN(n4691)
         );
  OAI211_X1 U5882 ( .C1(n4849), .C2(n6405), .A(n4692), .B(n4691), .ZN(U3096)
         );
  AOI22_X1 U5883 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4702), .B1(n6378), 
        .B2(n4701), .ZN(n4694) );
  AOI22_X1 U5884 ( .A1(n6356), .A2(n6284), .B1(n6362), .B2(n4703), .ZN(n4693)
         );
  OAI211_X1 U5885 ( .C1(n4849), .C2(n6295), .A(n4694), .B(n4693), .ZN(U3092)
         );
  INV_X1 U5886 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4697) );
  INV_X1 U5887 ( .A(n4810), .ZN(n4695) );
  OAI21_X1 U5888 ( .B1(n3028), .B2(n4696), .A(n4695), .ZN(n6172) );
  OAI222_X1 U5889 ( .A1(n4698), .A2(n5487), .B1(n6055), .B2(n4697), .C1(n6172), 
        .C2(n6045), .ZN(U2851) );
  AOI22_X1 U5890 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4702), .B1(n6390), 
        .B2(n4701), .ZN(n4700) );
  AOI22_X1 U5891 ( .A1(n6356), .A2(n6298), .B1(n6388), .B2(n4703), .ZN(n4699)
         );
  OAI211_X1 U5892 ( .C1(n4849), .C2(n6301), .A(n4700), .B(n4699), .ZN(U3094)
         );
  AOI22_X1 U5893 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4702), .B1(n6384), 
        .B2(n4701), .ZN(n4705) );
  AOI22_X1 U5894 ( .A1(n6356), .A2(n6383), .B1(n6382), .B2(n4703), .ZN(n4704)
         );
  OAI211_X1 U5895 ( .C1(n4849), .C2(n6387), .A(n4705), .B(n4704), .ZN(U3093)
         );
  XOR2_X1 U5896 ( .A(n4707), .B(n4706), .Z(n5008) );
  INV_X1 U5897 ( .A(n5008), .ZN(n4712) );
  AOI22_X1 U5898 ( .A1(n5279), .A2(DATAI_7_), .B1(n6065), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U5899 ( .B1(n4712), .B2(n5843), .A(n4708), .ZN(U2884) );
  AOI21_X1 U5900 ( .B1(n4710), .B2(n4709), .A(n3028), .ZN(n6180) );
  AOI22_X1 U5901 ( .A1(n6180), .A2(n6051), .B1(EBX_REG_7__SCAN_IN), .B2(n5479), 
        .ZN(n4711) );
  OAI21_X1 U5902 ( .B1(n4712), .B2(n5487), .A(n4711), .ZN(U2852) );
  OAI21_X1 U5903 ( .B1(n4715), .B2(n4714), .A(n4713), .ZN(n6113) );
  NOR2_X1 U5904 ( .A1(n6023), .A2(n6193), .ZN(n4722) );
  OR2_X1 U5905 ( .A1(n4716), .A2(n6214), .ZN(n4717) );
  NAND2_X1 U5906 ( .A1(n4717), .A2(n6209), .ZN(n6203) );
  NOR2_X1 U5907 ( .A1(n4718), .A2(n6203), .ZN(n4720) );
  MUX2_X1 U5908 ( .A(n4720), .B(n4719), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4721) );
  AOI211_X1 U5909 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6213), .A(n4722), .B(n4721), 
        .ZN(n4723) );
  OAI21_X1 U5910 ( .B1(n6201), .B2(n6113), .A(n4723), .ZN(U3012) );
  INV_X1 U5911 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5912 ( .A1(n6382), .A2(n6276), .B1(n6384), .B2(n6275), .ZN(n4724)
         );
  OAI21_X1 U5913 ( .B1(n6387), .B2(n6311), .A(n4724), .ZN(n4725) );
  AOI21_X1 U5914 ( .B1(n6383), .B2(n6277), .A(n4725), .ZN(n4726) );
  OAI21_X1 U5915 ( .B1(n4736), .B2(n4727), .A(n4726), .ZN(U3069) );
  INV_X1 U5916 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5917 ( .A1(n6412), .A2(n6276), .B1(n6415), .B2(n6275), .ZN(n4728)
         );
  OAI21_X1 U5918 ( .B1(n6419), .B2(n6311), .A(n4728), .ZN(n4729) );
  AOI21_X1 U5919 ( .B1(n6413), .B2(n6277), .A(n4729), .ZN(n4730) );
  OAI21_X1 U5920 ( .B1(n4736), .B2(n4731), .A(n4730), .ZN(U3074) );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5922 ( .A1(n6425), .A2(n6275), .B1(n6421), .B2(n6276), .ZN(n4732)
         );
  OAI21_X1 U5923 ( .B1(n6319), .B2(n6311), .A(n4732), .ZN(n4733) );
  AOI21_X1 U5924 ( .B1(n6312), .B2(n6277), .A(n4733), .ZN(n4734) );
  OAI21_X1 U5925 ( .B1(n4736), .B2(n4735), .A(n4734), .ZN(U3075) );
  INV_X1 U5926 ( .A(n5769), .ZN(n6433) );
  NAND2_X1 U5927 ( .A1(n6069), .A2(n3006), .ZN(n5160) );
  NOR2_X1 U5928 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4741), .ZN(n6100) );
  AOI22_X1 U5929 ( .A1(n6571), .A2(UWORD_REG_14__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U5930 ( .B1(n4743), .B2(n5160), .A(n4742), .ZN(U2893) );
  AOI22_X1 U5931 ( .A1(n6571), .A2(UWORD_REG_11__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4744) );
  OAI21_X1 U5932 ( .B1(n4745), .B2(n5160), .A(n4744), .ZN(U2896) );
  AOI22_X1 U5933 ( .A1(n6571), .A2(UWORD_REG_10__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4746) );
  OAI21_X1 U5934 ( .B1(n4747), .B2(n5160), .A(n4746), .ZN(U2897) );
  AOI22_X1 U5935 ( .A1(n6571), .A2(UWORD_REG_13__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4748) );
  OAI21_X1 U5936 ( .B1(n4749), .B2(n5160), .A(n4748), .ZN(U2894) );
  AOI22_X1 U5937 ( .A1(n6571), .A2(UWORD_REG_12__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4750) );
  OAI21_X1 U5938 ( .B1(n4751), .B2(n5160), .A(n4750), .ZN(U2895) );
  AOI22_X1 U5939 ( .A1(n6571), .A2(UWORD_REG_9__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5940 ( .B1(n4753), .B2(n5160), .A(n4752), .ZN(U2898) );
  AOI22_X1 U5941 ( .A1(n6571), .A2(UWORD_REG_8__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4754) );
  OAI21_X1 U5942 ( .B1(n4755), .B2(n5160), .A(n4754), .ZN(U2899) );
  AND2_X1 U5943 ( .A1(n4671), .A2(n4756), .ZN(n4758) );
  OR2_X1 U5944 ( .A1(n4758), .A2(n4757), .ZN(n6010) );
  AOI22_X1 U5945 ( .A1(n5279), .A2(DATAI_9_), .B1(n6065), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4759) );
  OAI21_X1 U5946 ( .B1(n6010), .B2(n5843), .A(n4759), .ZN(U2882) );
  NAND2_X1 U5947 ( .A1(n2988), .A2(n4760), .ZN(n6281) );
  NOR2_X1 U5948 ( .A1(n6281), .A2(n4313), .ZN(n4761) );
  NOR2_X1 U5949 ( .A1(n4920), .A2(n6371), .ZN(n4762) );
  INV_X1 U5950 ( .A(n6328), .ZN(n4884) );
  AOI21_X1 U5951 ( .B1(n4820), .B2(n4762), .A(n4884), .ZN(n4767) );
  NOR2_X1 U5952 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4763), .ZN(n4773)
         );
  INV_X1 U5953 ( .A(n4773), .ZN(n4815) );
  INV_X1 U5954 ( .A(n5179), .ZN(n4764) );
  OR2_X1 U5955 ( .A1(n5180), .A2(n4764), .ZN(n5012) );
  INV_X1 U5956 ( .A(n5012), .ZN(n4770) );
  OAI21_X1 U5957 ( .B1(n4770), .B2(n6374), .A(n4765), .ZN(n5016) );
  AOI211_X1 U5958 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4815), .A(n5182), .B(
        n5016), .ZN(n4766) );
  OAI21_X1 U5959 ( .B1(n4768), .B2(n4767), .A(n4766), .ZN(n4813) );
  INV_X1 U5960 ( .A(n4920), .ZN(n4814) );
  INV_X1 U5961 ( .A(n4768), .ZN(n4769) );
  OR2_X1 U5962 ( .A1(n4769), .A2(n6371), .ZN(n4772) );
  NAND2_X1 U5963 ( .A1(n5087), .A2(n4770), .ZN(n4771) );
  NAND2_X1 U5964 ( .A1(n4772), .A2(n4771), .ZN(n4817) );
  AOI22_X1 U5965 ( .A1(n6412), .A2(n4773), .B1(n6415), .B2(n4817), .ZN(n4776)
         );
  INV_X1 U5966 ( .A(n4820), .ZN(n4774) );
  NAND2_X1 U5967 ( .A1(n4774), .A2(n6350), .ZN(n4775) );
  OAI211_X1 U5968 ( .C1(n4814), .C2(n6353), .A(n4776), .B(n4775), .ZN(n4777)
         );
  AOI21_X1 U5969 ( .B1(n4813), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n4777), 
        .ZN(n4778) );
  INV_X1 U5970 ( .A(n4778), .ZN(U3026) );
  NOR2_X1 U5971 ( .A1(n4820), .A2(n6263), .ZN(n4782) );
  NAND2_X1 U5972 ( .A1(n4920), .A2(n6260), .ZN(n4780) );
  NAND2_X1 U5973 ( .A1(n4817), .A2(n6408), .ZN(n4779) );
  OAI211_X1 U5974 ( .C1(n5207), .C2(n4815), .A(n4780), .B(n4779), .ZN(n4781)
         );
  AOI211_X1 U5975 ( .C1(n4813), .C2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n4782), 
        .B(n4781), .ZN(n4783) );
  INV_X1 U5976 ( .A(n4783), .ZN(U3025) );
  NOR2_X1 U5977 ( .A1(n4820), .A2(n6257), .ZN(n4787) );
  NAND2_X1 U5978 ( .A1(n4920), .A2(n6254), .ZN(n4785) );
  NAND2_X1 U5979 ( .A1(n4817), .A2(n6396), .ZN(n4784) );
  OAI211_X1 U5980 ( .C1(n5215), .C2(n4815), .A(n4785), .B(n4784), .ZN(n4786)
         );
  AOI211_X1 U5981 ( .C1(n4813), .C2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n4787), 
        .B(n4786), .ZN(n4788) );
  INV_X1 U5982 ( .A(n4788), .ZN(U3023) );
  NOR2_X1 U5983 ( .A1(n4820), .A2(n6387), .ZN(n4792) );
  NAND2_X1 U5984 ( .A1(n4920), .A2(n6383), .ZN(n4790) );
  NAND2_X1 U5985 ( .A1(n4817), .A2(n6384), .ZN(n4789) );
  OAI211_X1 U5986 ( .C1(n5226), .C2(n4815), .A(n4790), .B(n4789), .ZN(n4791)
         );
  AOI211_X1 U5987 ( .C1(n4813), .C2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n4792), 
        .B(n4791), .ZN(n4793) );
  INV_X1 U5988 ( .A(n4793), .ZN(U3021) );
  NOR2_X1 U5989 ( .A1(n4820), .A2(n6405), .ZN(n4797) );
  NAND2_X1 U5990 ( .A1(n4920), .A2(n6401), .ZN(n4795) );
  NAND2_X1 U5991 ( .A1(n4817), .A2(n6402), .ZN(n4794) );
  OAI211_X1 U5992 ( .C1(n5203), .C2(n4815), .A(n4795), .B(n4794), .ZN(n4796)
         );
  AOI211_X1 U5993 ( .C1(n4813), .C2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n4797), 
        .B(n4796), .ZN(n4798) );
  INV_X1 U5994 ( .A(n4798), .ZN(U3024) );
  NOR2_X1 U5995 ( .A1(n4820), .A2(n6301), .ZN(n4802) );
  NAND2_X1 U5996 ( .A1(n4920), .A2(n6298), .ZN(n4800) );
  NAND2_X1 U5997 ( .A1(n4817), .A2(n6390), .ZN(n4799) );
  OAI211_X1 U5998 ( .C1(n5219), .C2(n4815), .A(n4800), .B(n4799), .ZN(n4801)
         );
  AOI211_X1 U5999 ( .C1(n4813), .C2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n4802), 
        .B(n4801), .ZN(n4803) );
  INV_X1 U6000 ( .A(n4803), .ZN(U3022) );
  NOR2_X1 U6001 ( .A1(n4820), .A2(n6295), .ZN(n4807) );
  NAND2_X1 U6002 ( .A1(n4920), .A2(n6284), .ZN(n4805) );
  NAND2_X1 U6003 ( .A1(n4817), .A2(n6378), .ZN(n4804) );
  OAI211_X1 U6004 ( .C1(n5199), .C2(n4815), .A(n4805), .B(n4804), .ZN(n4806)
         );
  AOI211_X1 U6005 ( .C1(n4813), .C2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n4807), 
        .B(n4806), .ZN(n4808) );
  INV_X1 U6006 ( .A(n4808), .ZN(U3020) );
  INV_X1 U6007 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4812) );
  OR2_X1 U6008 ( .A1(n4810), .A2(n4809), .ZN(n4811) );
  NAND2_X1 U6009 ( .A1(n5976), .A2(n4811), .ZN(n6164) );
  OAI222_X1 U6010 ( .A1(n6010), .A2(n5487), .B1(n4812), .B2(n6055), .C1(n6045), 
        .C2(n6164), .ZN(U2850) );
  NAND2_X1 U6011 ( .A1(n4813), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4819) );
  OAI22_X1 U6012 ( .A1(n5105), .A2(n4815), .B1(n4814), .B2(n6430), .ZN(n4816)
         );
  AOI21_X1 U6013 ( .B1(n6425), .B2(n4817), .A(n4816), .ZN(n4818) );
  OAI211_X1 U6014 ( .C1(n4820), .C2(n6319), .A(n4819), .B(n4818), .ZN(U3027)
         );
  NOR2_X1 U6015 ( .A1(n4827), .A2(n4267), .ZN(n4821) );
  NAND3_X1 U6016 ( .A1(n3006), .A2(n5413), .A3(n4822), .ZN(n4823) );
  AND2_X1 U6017 ( .A1(n4824), .A2(n4823), .ZN(n4825) );
  NAND2_X1 U6018 ( .A1(n3307), .A2(n3236), .ZN(n4826) );
  OR2_X1 U6019 ( .A1(n4827), .A2(n4826), .ZN(n6037) );
  OAI22_X1 U6020 ( .A1(n4828), .A2(n6016), .B1(n6037), .B2(n4319), .ZN(n4829)
         );
  AOI21_X1 U6021 ( .B1(n6041), .B2(n4830), .A(n4829), .ZN(n4837) );
  INV_X1 U6022 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4833) );
  INV_X1 U6023 ( .A(n5269), .ZN(n5075) );
  AOI22_X1 U6024 ( .A1(n6032), .A2(n4833), .B1(n5075), .B2(REIP_REG_1__SCAN_IN), .ZN(n4836) );
  NOR2_X1 U6025 ( .A1(n5267), .A2(REIP_REG_1__SCAN_IN), .ZN(n4929) );
  INV_X1 U6026 ( .A(n4929), .ZN(n4835) );
  NAND2_X1 U6027 ( .A1(n6031), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4834)
         );
  AND4_X1 U6028 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4838)
         );
  OAI21_X1 U6029 ( .B1(n4839), .B2(n6038), .A(n4838), .ZN(U2826) );
  NAND2_X1 U6030 ( .A1(n4849), .A2(n6429), .ZN(n4841) );
  AOI21_X1 U6031 ( .B1(n4841), .B2(STATEBS16_REG_SCAN_IN), .A(n6371), .ZN(
        n4846) );
  INV_X1 U6032 ( .A(n5087), .ZN(n6324) );
  NOR2_X1 U6033 ( .A1(n6324), .A2(n6446), .ZN(n4843) );
  AOI22_X1 U6034 ( .A1(n4846), .A2(n6369), .B1(n5180), .B2(n4843), .ZN(n4877)
         );
  INV_X1 U6035 ( .A(n6369), .ZN(n4845) );
  NAND3_X1 U6036 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4844), .ZN(n6375) );
  OR2_X1 U6037 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6375), .ZN(n4872)
         );
  AOI22_X1 U6038 ( .A1(n4846), .A2(n4845), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4872), .ZN(n4847) );
  NAND2_X1 U6039 ( .A1(n4871), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4852)
         );
  OAI22_X1 U6040 ( .A1(n6429), .A2(n6301), .B1(n5219), .B2(n4872), .ZN(n4850)
         );
  AOI21_X1 U6041 ( .B1(n4874), .B2(n6298), .A(n4850), .ZN(n4851) );
  OAI211_X1 U6042 ( .C1(n4877), .C2(n5128), .A(n4852), .B(n4851), .ZN(U3102)
         );
  NAND2_X1 U6043 ( .A1(n4871), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4855)
         );
  OAI22_X1 U6044 ( .A1(n6429), .A2(n6319), .B1(n5105), .B2(n4872), .ZN(n4853)
         );
  AOI21_X1 U6045 ( .B1(n4874), .B2(n6312), .A(n4853), .ZN(n4854) );
  OAI211_X1 U6046 ( .C1(n4877), .C2(n5194), .A(n4855), .B(n4854), .ZN(U3107)
         );
  NAND2_X1 U6047 ( .A1(n4871), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4858)
         );
  OAI22_X1 U6048 ( .A1(n6429), .A2(n6263), .B1(n5207), .B2(n4872), .ZN(n4856)
         );
  AOI21_X1 U6049 ( .B1(n4874), .B2(n6260), .A(n4856), .ZN(n4857) );
  OAI211_X1 U6050 ( .C1(n4877), .C2(n5100), .A(n4858), .B(n4857), .ZN(U3105)
         );
  INV_X1 U6051 ( .A(n6384), .ZN(n5114) );
  NAND2_X1 U6052 ( .A1(n4871), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4861)
         );
  OAI22_X1 U6053 ( .A1(n6429), .A2(n6387), .B1(n5226), .B2(n4872), .ZN(n4859)
         );
  AOI21_X1 U6054 ( .B1(n4874), .B2(n6383), .A(n4859), .ZN(n4860) );
  OAI211_X1 U6055 ( .C1(n4877), .C2(n5114), .A(n4861), .B(n4860), .ZN(U3101)
         );
  NAND2_X1 U6056 ( .A1(n4871), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4864)
         );
  OAI22_X1 U6057 ( .A1(n6429), .A2(n6257), .B1(n5215), .B2(n4872), .ZN(n4862)
         );
  AOI21_X1 U6058 ( .B1(n4874), .B2(n6254), .A(n4862), .ZN(n4863) );
  OAI211_X1 U6059 ( .C1(n4877), .C2(n5110), .A(n4864), .B(n4863), .ZN(U3103)
         );
  INV_X1 U6060 ( .A(n6415), .ZN(n5118) );
  NAND2_X1 U6061 ( .A1(n4871), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4867)
         );
  OAI22_X1 U6062 ( .A1(n6429), .A2(n6419), .B1(n5211), .B2(n4872), .ZN(n4865)
         );
  AOI21_X1 U6063 ( .B1(n4874), .B2(n6413), .A(n4865), .ZN(n4866) );
  OAI211_X1 U6064 ( .C1(n4877), .C2(n5118), .A(n4867), .B(n4866), .ZN(U3106)
         );
  NAND2_X1 U6065 ( .A1(n4871), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4870)
         );
  OAI22_X1 U6066 ( .A1(n6429), .A2(n6405), .B1(n5203), .B2(n4872), .ZN(n4868)
         );
  AOI21_X1 U6067 ( .B1(n4874), .B2(n6401), .A(n4868), .ZN(n4869) );
  OAI211_X1 U6068 ( .C1(n4877), .C2(n5122), .A(n4870), .B(n4869), .ZN(U3104)
         );
  NAND2_X1 U6069 ( .A1(n4871), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4876)
         );
  OAI22_X1 U6070 ( .A1(n6429), .A2(n6295), .B1(n5199), .B2(n4872), .ZN(n4873)
         );
  AOI21_X1 U6071 ( .B1(n4874), .B2(n6284), .A(n4873), .ZN(n4875) );
  OAI211_X1 U6072 ( .C1(n4877), .C2(n5096), .A(n4876), .B(n4875), .ZN(U3100)
         );
  OAI21_X1 U6073 ( .B1(n4878), .B2(n4880), .A(n4879), .ZN(n6181) );
  NAND2_X1 U6074 ( .A1(n6109), .A2(n4998), .ZN(n4881) );
  NAND2_X1 U6075 ( .A1(n6199), .A2(REIP_REG_7__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U6076 ( .C1(n5616), .C2(n4997), .A(n4881), .B(n6178), .ZN(n4882)
         );
  AOI21_X1 U6077 ( .B1(n5008), .B2(n6133), .A(n4882), .ZN(n4883) );
  OAI21_X1 U6078 ( .B1(n6124), .B2(n6181), .A(n4883), .ZN(U2979) );
  NAND3_X1 U6079 ( .A1(n4312), .A2(n3410), .A3(n2988), .ZN(n4885) );
  AOI21_X1 U6080 ( .B1(n4885), .B2(n6133), .A(n4884), .ZN(n4890) );
  INV_X1 U6081 ( .A(n5093), .ZN(n4886) );
  INV_X1 U6082 ( .A(n4917), .ZN(n4893) );
  AOI21_X1 U6083 ( .B1(n4887), .B2(n4886), .A(n4893), .ZN(n4891) );
  INV_X1 U6084 ( .A(n4891), .ZN(n4889) );
  AOI21_X1 U6085 ( .B1(n5086), .B2(n6371), .A(n6370), .ZN(n4888) );
  INV_X1 U6086 ( .A(n4921), .ZN(n4897) );
  INV_X1 U6087 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4896) );
  OAI22_X1 U6088 ( .A1(n4891), .A2(n6371), .B1(n5086), .B2(n6374), .ZN(n4898)
         );
  AOI22_X1 U6089 ( .A1(n6425), .A2(n4898), .B1(n6312), .B2(n2987), .ZN(n4895)
         );
  AOI22_X1 U6090 ( .A1(n6421), .A2(n4893), .B1(n6423), .B2(n4920), .ZN(n4894)
         );
  OAI211_X1 U6091 ( .C1(n4897), .C2(n4896), .A(n4895), .B(n4894), .ZN(U3147)
         );
  INV_X1 U6092 ( .A(n4898), .ZN(n4918) );
  OAI22_X1 U6093 ( .A1(n5226), .A2(n4917), .B1(n4918), .B2(n5114), .ZN(n4899)
         );
  AOI21_X1 U6094 ( .B1(n6336), .B2(n4920), .A(n4899), .ZN(n4901) );
  NAND2_X1 U6095 ( .A1(n4921), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4900)
         );
  OAI211_X1 U6096 ( .C1(n6785), .C2(n6339), .A(n4901), .B(n4900), .ZN(U3141)
         );
  OAI22_X1 U6097 ( .A1(n5219), .A2(n4917), .B1(n4918), .B2(n5128), .ZN(n4902)
         );
  AOI21_X1 U6098 ( .B1(n6389), .B2(n4920), .A(n4902), .ZN(n4904) );
  NAND2_X1 U6099 ( .A1(n4921), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4903)
         );
  OAI211_X1 U6100 ( .C1(n6785), .C2(n6393), .A(n4904), .B(n4903), .ZN(U3142)
         );
  OAI22_X1 U6101 ( .A1(n5207), .A2(n4917), .B1(n4918), .B2(n5100), .ZN(n4905)
         );
  AOI21_X1 U6102 ( .B1(n6407), .B2(n4920), .A(n4905), .ZN(n4907) );
  NAND2_X1 U6103 ( .A1(n4921), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4906)
         );
  OAI211_X1 U6104 ( .C1(n6785), .C2(n6411), .A(n4907), .B(n4906), .ZN(U3145)
         );
  OAI22_X1 U6105 ( .A1(n5199), .A2(n4917), .B1(n4918), .B2(n5096), .ZN(n4908)
         );
  AOI21_X1 U6106 ( .B1(n6363), .B2(n4920), .A(n4908), .ZN(n4910) );
  NAND2_X1 U6107 ( .A1(n4921), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4909)
         );
  OAI211_X1 U6108 ( .C1(n6785), .C2(n6381), .A(n4910), .B(n4909), .ZN(U3140)
         );
  OAI22_X1 U6109 ( .A1(n5203), .A2(n4917), .B1(n4918), .B2(n5122), .ZN(n4911)
         );
  AOI21_X1 U6110 ( .B1(n6344), .B2(n4920), .A(n4911), .ZN(n4913) );
  NAND2_X1 U6111 ( .A1(n4921), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4912)
         );
  OAI211_X1 U6112 ( .C1(n6785), .C2(n6347), .A(n4913), .B(n4912), .ZN(U3144)
         );
  OAI22_X1 U6113 ( .A1(n5215), .A2(n4917), .B1(n4918), .B2(n5110), .ZN(n4914)
         );
  AOI21_X1 U6114 ( .B1(n6395), .B2(n4920), .A(n4914), .ZN(n4916) );
  NAND2_X1 U6115 ( .A1(n4921), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4915)
         );
  OAI211_X1 U6116 ( .C1(n6785), .C2(n6399), .A(n4916), .B(n4915), .ZN(U3143)
         );
  OAI22_X1 U6117 ( .A1(n5118), .A2(n4918), .B1(n4917), .B2(n5211), .ZN(n4919)
         );
  AOI21_X1 U6118 ( .B1(n6350), .B2(n4920), .A(n4919), .ZN(n4923) );
  NAND2_X1 U6119 ( .A1(n4921), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4922)
         );
  OAI211_X1 U6120 ( .C1(n6785), .C2(n6353), .A(n4923), .B(n4922), .ZN(U3146)
         );
  OAI21_X1 U6121 ( .B1(n4757), .B2(n4926), .A(n4925), .ZN(n5999) );
  AOI22_X1 U6122 ( .A1(n5279), .A2(DATAI_10_), .B1(n6065), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4927) );
  OAI21_X1 U6123 ( .B1(n5999), .B2(n5843), .A(n4927), .ZN(U2881) );
  XNOR2_X1 U6124 ( .A(n5976), .B(n5978), .ZN(n6151) );
  AOI22_X1 U6125 ( .A1(n6151), .A2(n6051), .B1(EBX_REG_10__SCAN_IN), .B2(n5479), .ZN(n4928) );
  OAI21_X1 U6126 ( .B1(n5999), .B2(n5487), .A(n4928), .ZN(U2849) );
  NOR2_X1 U6127 ( .A1(n4929), .A2(n5075), .ZN(n6030) );
  INV_X1 U6128 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U6129 ( .A1(n6134), .A2(n5070), .ZN(n4937) );
  NAND2_X1 U6130 ( .A1(n6034), .A2(EBX_REG_2__SCAN_IN), .ZN(n4934) );
  INV_X1 U6131 ( .A(n6037), .ZN(n4977) );
  NAND2_X1 U6132 ( .A1(n4977), .A2(n4317), .ZN(n4933) );
  INV_X1 U6133 ( .A(n6138), .ZN(n4930) );
  AOI22_X1 U6134 ( .A1(n6031), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6032), 
        .B2(n4930), .ZN(n4932) );
  NAND3_X1 U6135 ( .A1(n5061), .A2(REIP_REG_1__SCAN_IN), .A3(n4938), .ZN(n4931) );
  NAND4_X1 U6136 ( .A1(n4934), .A2(n4933), .A3(n4932), .A4(n4931), .ZN(n4935)
         );
  AOI21_X1 U6137 ( .B1(n6041), .B2(n6212), .A(n4935), .ZN(n4936) );
  OAI211_X1 U6138 ( .C1(n6030), .C2(n4938), .A(n4937), .B(n4936), .ZN(U2825)
         );
  NAND2_X1 U6139 ( .A1(n4958), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4942) );
  INV_X1 U6140 ( .A(n4959), .ZN(n4940) );
  OAI22_X1 U6141 ( .A1(n5105), .A2(n4960), .B1(n6267), .B2(n6319), .ZN(n4939)
         );
  AOI21_X1 U6142 ( .B1(n6425), .B2(n4940), .A(n4939), .ZN(n4941) );
  OAI211_X1 U6143 ( .C1(n4964), .C2(n6430), .A(n4942), .B(n4941), .ZN(U3043)
         );
  NAND2_X1 U6144 ( .A1(n4958), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4945) );
  OAI22_X1 U6145 ( .A1(n5203), .A2(n4960), .B1(n4959), .B2(n5122), .ZN(n4943)
         );
  AOI21_X1 U6146 ( .B1(n6344), .B2(n6268), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6147 ( .C1(n4964), .C2(n6347), .A(n4945), .B(n4944), .ZN(U3040)
         );
  NAND2_X1 U6148 ( .A1(n4958), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4948) );
  OAI22_X1 U6149 ( .A1(n5219), .A2(n4960), .B1(n4959), .B2(n5128), .ZN(n4946)
         );
  AOI21_X1 U6150 ( .B1(n6389), .B2(n6268), .A(n4946), .ZN(n4947) );
  OAI211_X1 U6151 ( .C1(n4964), .C2(n6393), .A(n4948), .B(n4947), .ZN(U3038)
         );
  NAND2_X1 U6152 ( .A1(n4958), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4951) );
  OAI22_X1 U6153 ( .A1(n5207), .A2(n4960), .B1(n4959), .B2(n5100), .ZN(n4949)
         );
  AOI21_X1 U6154 ( .B1(n6407), .B2(n6268), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6155 ( .C1(n4964), .C2(n6411), .A(n4951), .B(n4950), .ZN(U3041)
         );
  NAND2_X1 U6156 ( .A1(n4958), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4954) );
  OAI22_X1 U6157 ( .A1(n5226), .A2(n4960), .B1(n4959), .B2(n5114), .ZN(n4952)
         );
  AOI21_X1 U6158 ( .B1(n6336), .B2(n6268), .A(n4952), .ZN(n4953) );
  OAI211_X1 U6159 ( .C1(n4964), .C2(n6339), .A(n4954), .B(n4953), .ZN(U3037)
         );
  NAND2_X1 U6160 ( .A1(n4958), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4957) );
  OAI22_X1 U6161 ( .A1(n5118), .A2(n4959), .B1(n5211), .B2(n4960), .ZN(n4955)
         );
  AOI21_X1 U6162 ( .B1(n6350), .B2(n6268), .A(n4955), .ZN(n4956) );
  OAI211_X1 U6163 ( .C1(n4964), .C2(n6353), .A(n4957), .B(n4956), .ZN(U3042)
         );
  NAND2_X1 U6164 ( .A1(n4958), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4963) );
  OAI22_X1 U6165 ( .A1(n5215), .A2(n4960), .B1(n4959), .B2(n5110), .ZN(n4961)
         );
  AOI21_X1 U6166 ( .B1(n6395), .B2(n6268), .A(n4961), .ZN(n4962) );
  OAI211_X1 U6167 ( .C1(n4964), .C2(n6399), .A(n4963), .B(n4962), .ZN(U3039)
         );
  OAI21_X1 U6168 ( .B1(n4967), .B2(n4966), .A(n4965), .ZN(n6171) );
  AOI22_X1 U6169 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6199), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4968) );
  OAI21_X1 U6170 ( .B1(n4985), .B2(n6139), .A(n4968), .ZN(n4969) );
  AOI21_X1 U6171 ( .B1(n4988), .B2(n6133), .A(n4969), .ZN(n4970) );
  OAI21_X1 U6172 ( .B1(n6171), .B2(n6124), .A(n4970), .ZN(U2978) );
  OAI21_X1 U6173 ( .B1(n6031), .B2(n6032), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4971) );
  OAI21_X1 U6174 ( .B1(n4972), .B2(n6016), .A(n4971), .ZN(n4976) );
  INV_X1 U6175 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4973) );
  OAI22_X1 U6176 ( .A1(n6024), .A2(n4974), .B1(n5403), .B2(n4973), .ZN(n4975)
         );
  AOI211_X1 U6177 ( .C1(n6368), .C2(n4977), .A(n4976), .B(n4975), .ZN(n4978)
         );
  OAI21_X1 U6178 ( .B1(n6038), .B2(n4979), .A(n4978), .ZN(U2827) );
  AOI22_X1 U6179 ( .A1(EBX_REG_8__SCAN_IN), .A2(n6034), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6031), .ZN(n4981) );
  NAND2_X1 U6180 ( .A1(n5269), .A2(n4980), .ZN(n5994) );
  OAI211_X1 U6181 ( .C1(n6024), .C2(n6172), .A(n4981), .B(n5994), .ZN(n4987)
         );
  NOR2_X1 U6182 ( .A1(n5267), .A2(n4982), .ZN(n5986) );
  NAND2_X1 U6183 ( .A1(n4983), .A2(n5269), .ZN(n5993) );
  OAI211_X1 U6184 ( .C1(REIP_REG_8__SCAN_IN), .C2(n5986), .A(n5993), .B(n5992), 
        .ZN(n4984) );
  OAI21_X1 U6185 ( .B1(n6029), .B2(n4985), .A(n4984), .ZN(n4986) );
  AOI211_X1 U6186 ( .C1(n4988), .C2(n6026), .A(n4987), .B(n4986), .ZN(n4989)
         );
  INV_X1 U6187 ( .A(n4989), .ZN(U2819) );
  INV_X1 U6188 ( .A(n4990), .ZN(n4993) );
  AOI21_X1 U6189 ( .B1(n4993), .B2(n4925), .A(n3984), .ZN(n6110) );
  INV_X1 U6190 ( .A(n6110), .ZN(n4995) );
  AOI22_X1 U6191 ( .A1(n5279), .A2(DATAI_11_), .B1(n6065), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6192 ( .B1(n4995), .B2(n5843), .A(n4994), .ZN(U2880) );
  AOI22_X1 U6193 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6034), .B1(n6041), .B2(n6180), 
        .ZN(n4996) );
  OAI211_X1 U6194 ( .C1(n6005), .C2(n4997), .A(n4996), .B(n5994), .ZN(n5007)
         );
  INV_X1 U6195 ( .A(n4998), .ZN(n5005) );
  NOR3_X1 U6196 ( .A1(n5267), .A2(REIP_REG_6__SCAN_IN), .A3(n4999), .ZN(n6019)
         );
  INV_X1 U6197 ( .A(n4999), .ZN(n5000) );
  OAI21_X1 U6198 ( .B1(n5267), .B2(n5000), .A(n5269), .ZN(n6020) );
  OAI21_X1 U6199 ( .B1(n6019), .B2(n6020), .A(REIP_REG_7__SCAN_IN), .ZN(n5004)
         );
  INV_X1 U6200 ( .A(n5001), .ZN(n5002) );
  OR3_X1 U6201 ( .A1(n5267), .A2(REIP_REG_7__SCAN_IN), .A3(n5002), .ZN(n5003)
         );
  OAI211_X1 U6202 ( .C1(n6029), .C2(n5005), .A(n5004), .B(n5003), .ZN(n5006)
         );
  AOI211_X1 U6203 ( .C1(n5008), .C2(n6026), .A(n5007), .B(n5006), .ZN(n5009)
         );
  INV_X1 U6204 ( .A(n5009), .ZN(U2820) );
  INV_X1 U6205 ( .A(n6281), .ZN(n5176) );
  AND2_X1 U6206 ( .A1(n5176), .A2(n3873), .ZN(n5010) );
  NOR2_X1 U6207 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5011), .ZN(n5022)
         );
  INV_X1 U6208 ( .A(n5022), .ZN(n5044) );
  NAND2_X1 U6209 ( .A1(n6322), .A2(n6365), .ZN(n5013) );
  INV_X1 U6210 ( .A(n5182), .ZN(n6331) );
  OAI22_X1 U6211 ( .A1(n5013), .A2(n5178), .B1(n6331), .B2(n5012), .ZN(n5042)
         );
  AOI21_X1 U6212 ( .B1(n5047), .B2(n6274), .A(n6758), .ZN(n5014) );
  NOR3_X1 U6213 ( .A1(n5015), .A2(n5014), .A3(n6371), .ZN(n5017) );
  NOR3_X1 U6214 ( .A1(n5087), .A2(n5017), .A3(n5016), .ZN(n5018) );
  AOI22_X1 U6215 ( .A1(n5042), .A2(n6402), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5041), .ZN(n5019) );
  OAI21_X1 U6216 ( .B1(n5203), .B2(n5044), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6217 ( .B1(n6401), .B2(n6264), .A(n5020), .ZN(n5021) );
  OAI21_X1 U6218 ( .B1(n6405), .B2(n5047), .A(n5021), .ZN(U3056) );
  AOI22_X1 U6219 ( .A1(n6421), .A2(n5022), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5041), .ZN(n5023) );
  OAI21_X1 U6220 ( .B1(n6430), .B2(n6274), .A(n5023), .ZN(n5024) );
  AOI21_X1 U6221 ( .B1(n6425), .B2(n5042), .A(n5024), .ZN(n5025) );
  OAI21_X1 U6222 ( .B1(n6319), .B2(n5047), .A(n5025), .ZN(U3059) );
  AOI22_X1 U6223 ( .A1(n6415), .A2(n5042), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5041), .ZN(n5026) );
  OAI21_X1 U6224 ( .B1(n5211), .B2(n5044), .A(n5026), .ZN(n5027) );
  AOI21_X1 U6225 ( .B1(n6413), .B2(n6264), .A(n5027), .ZN(n5028) );
  OAI21_X1 U6226 ( .B1(n6419), .B2(n5047), .A(n5028), .ZN(U3058) );
  AOI22_X1 U6227 ( .A1(n5042), .A2(n6378), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5041), .ZN(n5029) );
  OAI21_X1 U6228 ( .B1(n5199), .B2(n5044), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6229 ( .B1(n6284), .B2(n6264), .A(n5030), .ZN(n5031) );
  OAI21_X1 U6230 ( .B1(n6295), .B2(n5047), .A(n5031), .ZN(U3052) );
  AOI22_X1 U6231 ( .A1(n5042), .A2(n6384), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5041), .ZN(n5032) );
  OAI21_X1 U6232 ( .B1(n5226), .B2(n5044), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6233 ( .B1(n6383), .B2(n6264), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6234 ( .B1(n6387), .B2(n5047), .A(n5034), .ZN(U3053) );
  AOI22_X1 U6235 ( .A1(n5042), .A2(n6396), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5041), .ZN(n5035) );
  OAI21_X1 U6236 ( .B1(n5215), .B2(n5044), .A(n5035), .ZN(n5036) );
  AOI21_X1 U6237 ( .B1(n6254), .B2(n6264), .A(n5036), .ZN(n5037) );
  OAI21_X1 U6238 ( .B1(n6257), .B2(n5047), .A(n5037), .ZN(U3055) );
  AOI22_X1 U6239 ( .A1(n5042), .A2(n6408), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5041), .ZN(n5038) );
  OAI21_X1 U6240 ( .B1(n5207), .B2(n5044), .A(n5038), .ZN(n5039) );
  AOI21_X1 U6241 ( .B1(n6260), .B2(n6264), .A(n5039), .ZN(n5040) );
  OAI21_X1 U6242 ( .B1(n6263), .B2(n5047), .A(n5040), .ZN(U3057) );
  AOI22_X1 U6243 ( .A1(n5042), .A2(n6390), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5041), .ZN(n5043) );
  OAI21_X1 U6244 ( .B1(n5219), .B2(n5044), .A(n5043), .ZN(n5045) );
  AOI21_X1 U6245 ( .B1(n6298), .B2(n6264), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6246 ( .B1(n6301), .B2(n5047), .A(n5046), .ZN(U3054) );
  XOR2_X1 U6247 ( .A(n5048), .B(n4992), .Z(n5256) );
  INV_X1 U6248 ( .A(n5254), .ZN(n5057) );
  INV_X1 U6249 ( .A(n5049), .ZN(n5052) );
  NAND2_X1 U6250 ( .A1(n5061), .A2(n5052), .ZN(n5965) );
  AND2_X1 U6251 ( .A1(n5980), .A2(n5050), .ZN(n5051) );
  OR2_X1 U6252 ( .A1(n5051), .A2(n5901), .ZN(n5247) );
  OAI22_X1 U6253 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5965), .B1(n6024), .B2(
        n5247), .ZN(n5056) );
  OAI21_X1 U6254 ( .B1(n5267), .B2(n5052), .A(n5269), .ZN(n5985) );
  AOI22_X1 U6255 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6034), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5985), .ZN(n5053) );
  OAI211_X1 U6256 ( .C1(n6005), .C2(n5054), .A(n5053), .B(n5994), .ZN(n5055)
         );
  AOI211_X1 U6257 ( .C1(n6032), .C2(n5057), .A(n5056), .B(n5055), .ZN(n5058)
         );
  OAI21_X1 U6258 ( .B1(n5135), .B2(n6009), .A(n5058), .ZN(U2815) );
  AOI22_X1 U6259 ( .A1(n5279), .A2(DATAI_12_), .B1(n6065), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5059) );
  OAI21_X1 U6260 ( .B1(n5135), .B2(n5843), .A(n5059), .ZN(U2879) );
  INV_X1 U6261 ( .A(n6020), .ZN(n5064) );
  AOI21_X1 U6262 ( .B1(n5061), .B2(n5060), .A(REIP_REG_5__SCAN_IN), .ZN(n5063)
         );
  OAI22_X1 U6263 ( .A1(n5064), .A2(n5063), .B1(n5062), .B2(n6029), .ZN(n5069)
         );
  INV_X1 U6264 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U6265 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6034), .B1(n6041), .B2(n5065), 
        .ZN(n5066) );
  OAI211_X1 U6266 ( .C1(n6005), .C2(n5067), .A(n5066), .B(n5994), .ZN(n5068)
         );
  AOI211_X1 U6267 ( .C1(n5071), .C2(n5070), .A(n5069), .B(n5068), .ZN(n5072)
         );
  INV_X1 U6268 ( .A(n5072), .ZN(U2822) );
  NOR3_X1 U6269 ( .A1(n5267), .A2(REIP_REG_4__SCAN_IN), .A3(n5074), .ZN(n5083)
         );
  INV_X1 U6270 ( .A(n5073), .ZN(n5081) );
  OAI21_X1 U6271 ( .B1(n5075), .B2(n5074), .A(n5992), .ZN(n6044) );
  OAI22_X1 U6272 ( .A1(n5076), .A2(n6005), .B1(n6511), .B2(n6044), .ZN(n5079)
         );
  OAI22_X1 U6273 ( .A1(n6024), .A2(n6192), .B1(n5077), .B2(n6037), .ZN(n5078)
         );
  NOR3_X1 U6274 ( .A1(n6021), .A2(n5079), .A3(n5078), .ZN(n5080) );
  OAI21_X1 U6275 ( .B1(n5081), .B2(n6029), .A(n5080), .ZN(n5082) );
  AOI211_X1 U6276 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6034), .A(n5083), .B(n5082), 
        .ZN(n5084) );
  OAI21_X1 U6277 ( .B1(n5085), .B2(n6038), .A(n5084), .ZN(U2823) );
  NOR2_X1 U6278 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5086), .ZN(n5095)
         );
  NOR3_X1 U6279 ( .A1(n5088), .A2(n6446), .A3(n5087), .ZN(n5092) );
  OAI21_X1 U6280 ( .B1(n2987), .B2(n5089), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5090) );
  NAND3_X1 U6281 ( .A1(n5093), .A2(n6365), .A3(n5090), .ZN(n5091) );
  NAND2_X1 U6282 ( .A1(n5126), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5099)
         );
  INV_X1 U6283 ( .A(n5180), .ZN(n5094) );
  OAI33_X1 U6284 ( .A1(n6446), .A2(n5094), .A3(n6331), .B1(n5093), .B2(n6371), 
        .B3(n6322), .ZN(n5107) );
  INV_X1 U6285 ( .A(n5107), .ZN(n5129) );
  INV_X1 U6286 ( .A(n5095), .ZN(n5127) );
  OAI22_X1 U6287 ( .A1(n5129), .A2(n5096), .B1(n5199), .B2(n5127), .ZN(n5097)
         );
  AOI21_X1 U6288 ( .B1(n6363), .B2(n2987), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6289 ( .C1(n5134), .C2(n6381), .A(n5099), .B(n5098), .ZN(U3132)
         );
  NAND2_X1 U6290 ( .A1(n5126), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5103)
         );
  OAI22_X1 U6291 ( .A1(n5129), .A2(n5100), .B1(n5207), .B2(n5127), .ZN(n5101)
         );
  AOI21_X1 U6292 ( .B1(n6407), .B2(n2987), .A(n5101), .ZN(n5102) );
  OAI211_X1 U6293 ( .C1(n5134), .C2(n6411), .A(n5103), .B(n5102), .ZN(U3137)
         );
  NAND2_X1 U6294 ( .A1(n5126), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5109)
         );
  OAI22_X1 U6295 ( .A1(n5105), .A2(n5127), .B1(n6319), .B2(n6785), .ZN(n5106)
         );
  AOI21_X1 U6296 ( .B1(n6425), .B2(n5107), .A(n5106), .ZN(n5108) );
  OAI211_X1 U6297 ( .C1(n5134), .C2(n6430), .A(n5109), .B(n5108), .ZN(U3139)
         );
  NAND2_X1 U6298 ( .A1(n5126), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5113)
         );
  OAI22_X1 U6299 ( .A1(n5129), .A2(n5110), .B1(n5215), .B2(n5127), .ZN(n5111)
         );
  AOI21_X1 U6300 ( .B1(n6395), .B2(n2987), .A(n5111), .ZN(n5112) );
  OAI211_X1 U6301 ( .C1(n5134), .C2(n6399), .A(n5113), .B(n5112), .ZN(U3135)
         );
  NAND2_X1 U6302 ( .A1(n5126), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5117)
         );
  OAI22_X1 U6303 ( .A1(n5129), .A2(n5114), .B1(n5226), .B2(n5127), .ZN(n5115)
         );
  AOI21_X1 U6304 ( .B1(n6336), .B2(n2987), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6305 ( .C1(n5134), .C2(n6339), .A(n5117), .B(n5116), .ZN(U3133)
         );
  NAND2_X1 U6306 ( .A1(n5126), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5121)
         );
  OAI22_X1 U6307 ( .A1(n5129), .A2(n5118), .B1(n5211), .B2(n5127), .ZN(n5119)
         );
  AOI21_X1 U6308 ( .B1(n6350), .B2(n2987), .A(n5119), .ZN(n5120) );
  OAI211_X1 U6309 ( .C1(n5134), .C2(n6353), .A(n5121), .B(n5120), .ZN(U3138)
         );
  NAND2_X1 U6310 ( .A1(n5126), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5125)
         );
  OAI22_X1 U6311 ( .A1(n5129), .A2(n5122), .B1(n5203), .B2(n5127), .ZN(n5123)
         );
  AOI21_X1 U6312 ( .B1(n6344), .B2(n2987), .A(n5123), .ZN(n5124) );
  OAI211_X1 U6313 ( .C1(n5134), .C2(n6347), .A(n5125), .B(n5124), .ZN(U3136)
         );
  NAND2_X1 U6314 ( .A1(n5126), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5133)
         );
  OAI22_X1 U6315 ( .A1(n5129), .A2(n5128), .B1(n5219), .B2(n5127), .ZN(n5130)
         );
  AOI21_X1 U6316 ( .B1(n6389), .B2(n2987), .A(n5130), .ZN(n5132) );
  OAI211_X1 U6317 ( .C1(n5134), .C2(n6393), .A(n5133), .B(n5132), .ZN(U3134)
         );
  INV_X1 U6318 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5136) );
  OAI222_X1 U6319 ( .A1(n6045), .A2(n5247), .B1(n6055), .B2(n5136), .C1(n5487), 
        .C2(n5135), .ZN(U2847) );
  NAND2_X1 U6320 ( .A1(n5139), .A2(n5138), .ZN(n5140) );
  XNOR2_X1 U6321 ( .A(n5137), .B(n5140), .ZN(n6167) );
  NAND2_X1 U6322 ( .A1(n6167), .A2(n6135), .ZN(n5144) );
  NAND2_X1 U6323 ( .A1(n6213), .A2(REIP_REG_9__SCAN_IN), .ZN(n6163) );
  OAI21_X1 U6324 ( .B1(n5616), .B2(n6006), .A(n6163), .ZN(n5141) );
  AOI21_X1 U6325 ( .B1(n6109), .B2(n5142), .A(n5141), .ZN(n5143) );
  OAI211_X1 U6326 ( .C1(n6122), .C2(n6010), .A(n5144), .B(n5143), .ZN(U2977)
         );
  AOI22_X1 U6327 ( .A1(n6100), .A2(UWORD_REG_0__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5145) );
  OAI21_X1 U6328 ( .B1(n5146), .B2(n5160), .A(n5145), .ZN(U2907) );
  AOI22_X1 U6329 ( .A1(n6100), .A2(UWORD_REG_1__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5147) );
  OAI21_X1 U6330 ( .B1(n5148), .B2(n5160), .A(n5147), .ZN(U2906) );
  AOI22_X1 U6331 ( .A1(n6571), .A2(UWORD_REG_5__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5149) );
  OAI21_X1 U6332 ( .B1(n5150), .B2(n5160), .A(n5149), .ZN(U2902) );
  AOI22_X1 U6333 ( .A1(n6571), .A2(UWORD_REG_2__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5151) );
  OAI21_X1 U6334 ( .B1(n5152), .B2(n5160), .A(n5151), .ZN(U2905) );
  AOI22_X1 U6335 ( .A1(n6571), .A2(UWORD_REG_3__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5153) );
  OAI21_X1 U6336 ( .B1(n5154), .B2(n5160), .A(n5153), .ZN(U2904) );
  AOI22_X1 U6337 ( .A1(n6571), .A2(UWORD_REG_4__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5155) );
  OAI21_X1 U6338 ( .B1(n5156), .B2(n5160), .A(n5155), .ZN(U2903) );
  AOI22_X1 U6339 ( .A1(n6571), .A2(UWORD_REG_6__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5157) );
  OAI21_X1 U6340 ( .B1(n5158), .B2(n5160), .A(n5157), .ZN(U2901) );
  AOI22_X1 U6341 ( .A1(n6571), .A2(UWORD_REG_7__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5159) );
  OAI21_X1 U6342 ( .B1(n5161), .B2(n5160), .A(n5159), .ZN(U2900) );
  NAND2_X1 U6343 ( .A1(n6104), .A2(n5163), .ZN(n5164) );
  XNOR2_X1 U6344 ( .A(n5162), .B(n5164), .ZN(n6159) );
  NAND2_X1 U6345 ( .A1(n6159), .A2(n6135), .ZN(n5167) );
  NAND2_X1 U6346 ( .A1(n6213), .A2(REIP_REG_10__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U6347 ( .B1(n5616), .B2(n5996), .A(n6149), .ZN(n5165) );
  AOI21_X1 U6348 ( .B1(n6109), .B2(n6001), .A(n5165), .ZN(n5166) );
  OAI211_X1 U6349 ( .C1(n6122), .C2(n5999), .A(n5167), .B(n5166), .ZN(U2976)
         );
  INV_X1 U6350 ( .A(n5168), .ZN(n5171) );
  INV_X1 U6351 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6352 ( .A1(n5171), .A2(n5170), .ZN(n5173) );
  INV_X1 U6353 ( .A(n6048), .ZN(n5175) );
  AOI22_X1 U6354 ( .A1(n5279), .A2(DATAI_13_), .B1(n6065), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5174) );
  OAI21_X1 U6355 ( .B1(n5175), .B2(n5843), .A(n5174), .ZN(U2878) );
  NOR2_X1 U6356 ( .A1(n6322), .A2(n5178), .ZN(n5186) );
  OR2_X1 U6357 ( .A1(n5180), .A2(n5179), .ZN(n6323) );
  INV_X1 U6358 ( .A(n6323), .ZN(n5181) );
  AOI22_X1 U6359 ( .A1(n5186), .A2(n6365), .B1(n5182), .B2(n5181), .ZN(n5197)
         );
  NAND2_X1 U6360 ( .A1(n5184), .A2(n5183), .ZN(n5225) );
  INV_X1 U6361 ( .A(n5225), .ZN(n5192) );
  INV_X1 U6362 ( .A(n5228), .ZN(n5185) );
  AOI21_X1 U6363 ( .B1(n6418), .B2(n5185), .A(n6758), .ZN(n5187) );
  NOR3_X1 U6364 ( .A1(n5187), .A2(n5186), .A3(n6371), .ZN(n5190) );
  AOI21_X1 U6365 ( .B1(n6323), .B2(STATE2_REG_2__SCAN_IN), .A(n5188), .ZN(
        n6330) );
  INV_X1 U6366 ( .A(n6330), .ZN(n5189) );
  AOI211_X1 U6367 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5225), .A(n5190), .B(
        n5189), .ZN(n5191) );
  NAND2_X1 U6368 ( .A1(n5191), .A2(n6324), .ZN(n5222) );
  AOI22_X1 U6369 ( .A1(n6421), .A2(n5192), .B1(INSTQUEUE_REG_12__7__SCAN_IN), 
        .B2(n5222), .ZN(n5193) );
  OAI21_X1 U6370 ( .B1(n5194), .B2(n5197), .A(n5193), .ZN(n5195) );
  AOI21_X1 U6371 ( .B1(n6423), .B2(n5228), .A(n5195), .ZN(n5196) );
  OAI21_X1 U6372 ( .B1(n6430), .B2(n6418), .A(n5196), .ZN(U3123) );
  AOI22_X1 U6373 ( .A1(n5223), .A2(n6378), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5222), .ZN(n5198) );
  OAI21_X1 U6374 ( .B1(n5199), .B2(n5225), .A(n5198), .ZN(n5200) );
  AOI21_X1 U6375 ( .B1(n6363), .B2(n5228), .A(n5200), .ZN(n5201) );
  OAI21_X1 U6376 ( .B1(n6381), .B2(n6418), .A(n5201), .ZN(U3116) );
  AOI22_X1 U6377 ( .A1(n5223), .A2(n6402), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n5222), .ZN(n5202) );
  OAI21_X1 U6378 ( .B1(n5203), .B2(n5225), .A(n5202), .ZN(n5204) );
  AOI21_X1 U6379 ( .B1(n6344), .B2(n5228), .A(n5204), .ZN(n5205) );
  OAI21_X1 U6380 ( .B1(n6347), .B2(n6418), .A(n5205), .ZN(U3120) );
  AOI22_X1 U6381 ( .A1(n5223), .A2(n6408), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n5222), .ZN(n5206) );
  OAI21_X1 U6382 ( .B1(n5207), .B2(n5225), .A(n5206), .ZN(n5208) );
  AOI21_X1 U6383 ( .B1(n6407), .B2(n5228), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6384 ( .B1(n6411), .B2(n6418), .A(n5209), .ZN(U3121) );
  AOI22_X1 U6385 ( .A1(n6415), .A2(n5223), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5222), .ZN(n5210) );
  OAI21_X1 U6386 ( .B1(n5211), .B2(n5225), .A(n5210), .ZN(n5212) );
  AOI21_X1 U6387 ( .B1(n6350), .B2(n5228), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6388 ( .B1(n6353), .B2(n6418), .A(n5213), .ZN(U3122) );
  AOI22_X1 U6389 ( .A1(n5223), .A2(n6396), .B1(INSTQUEUE_REG_12__3__SCAN_IN), 
        .B2(n5222), .ZN(n5214) );
  OAI21_X1 U6390 ( .B1(n5215), .B2(n5225), .A(n5214), .ZN(n5216) );
  AOI21_X1 U6391 ( .B1(n6395), .B2(n5228), .A(n5216), .ZN(n5217) );
  OAI21_X1 U6392 ( .B1(n6399), .B2(n6418), .A(n5217), .ZN(U3119) );
  AOI22_X1 U6393 ( .A1(n5223), .A2(n6390), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n5222), .ZN(n5218) );
  OAI21_X1 U6394 ( .B1(n5219), .B2(n5225), .A(n5218), .ZN(n5220) );
  AOI21_X1 U6395 ( .B1(n6389), .B2(n5228), .A(n5220), .ZN(n5221) );
  OAI21_X1 U6396 ( .B1(n6393), .B2(n6418), .A(n5221), .ZN(U3118) );
  AOI22_X1 U6397 ( .A1(n5223), .A2(n6384), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n5222), .ZN(n5224) );
  OAI21_X1 U6398 ( .B1(n5226), .B2(n5225), .A(n5224), .ZN(n5227) );
  AOI21_X1 U6399 ( .B1(n6336), .B2(n5228), .A(n5227), .ZN(n5229) );
  OAI21_X1 U6400 ( .B1(n6339), .B2(n6418), .A(n5229), .ZN(U3117) );
  OAI21_X1 U6401 ( .B1(n5230), .B2(n5232), .A(n5231), .ZN(n5958) );
  AOI22_X1 U6402 ( .A1(n5279), .A2(DATAI_14_), .B1(n6065), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5233) );
  OAI21_X1 U6403 ( .B1(n5958), .B2(n5843), .A(n5233), .ZN(U2877) );
  INV_X1 U6404 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5235) );
  OAI21_X1 U6405 ( .B1(n5903), .B2(n5234), .A(n5262), .ZN(n5736) );
  OAI222_X1 U6406 ( .A1(n5958), .A2(n5487), .B1(n5235), .B2(n6055), .C1(n6045), 
        .C2(n5736), .ZN(U2845) );
  INV_X1 U6407 ( .A(n5237), .ZN(n5239) );
  NAND2_X1 U6408 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  XNOR2_X1 U6409 ( .A(n5236), .B(n5240), .ZN(n5251) );
  INV_X1 U6410 ( .A(n6141), .ZN(n5893) );
  NOR2_X1 U6411 ( .A1(n5893), .A2(n3515), .ZN(n5246) );
  OAI21_X1 U6412 ( .B1(n5241), .B2(n5717), .A(n5242), .ZN(n6142) );
  NAND3_X1 U6413 ( .A1(n5242), .A2(n5875), .A3(n5717), .ZN(n5243) );
  OAI21_X1 U6414 ( .B1(n6142), .B2(n3515), .A(n5243), .ZN(n5244) );
  INV_X1 U6415 ( .A(n5244), .ZN(n5245) );
  MUX2_X1 U6416 ( .A(n5246), .B(n5245), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5249) );
  NAND2_X1 U6417 ( .A1(n6213), .A2(REIP_REG_12__SCAN_IN), .ZN(n5253) );
  OAI21_X1 U6418 ( .B1(n5247), .B2(n6193), .A(n5253), .ZN(n5248) );
  AOI211_X1 U6419 ( .C1(n5251), .C2(n6229), .A(n5249), .B(n5248), .ZN(n5250)
         );
  INV_X1 U6420 ( .A(n5250), .ZN(U3006) );
  INV_X1 U6421 ( .A(n5251), .ZN(n5258) );
  NAND2_X1 U6422 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5252)
         );
  OAI211_X1 U6423 ( .C1(n6139), .C2(n5254), .A(n5253), .B(n5252), .ZN(n5255)
         );
  AOI21_X1 U6424 ( .B1(n5256), .B2(n6133), .A(n5255), .ZN(n5257) );
  OAI21_X1 U6425 ( .B1(n5258), .B2(n6124), .A(n5257), .ZN(U2974) );
  AND2_X1 U6426 ( .A1(n5231), .A2(n5259), .ZN(n5260) );
  OR2_X1 U6427 ( .A1(n5260), .A2(n3012), .ZN(n5611) );
  AND2_X1 U6428 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  OR2_X1 U6429 ( .A1(n3029), .A2(n5263), .ZN(n5276) );
  INV_X1 U6430 ( .A(n5276), .ZN(n5891) );
  NOR2_X1 U6431 ( .A1(n5267), .A2(n5265), .ZN(n5943) );
  AND2_X1 U6432 ( .A1(n5943), .A2(n6528), .ZN(n5945) );
  INV_X1 U6433 ( .A(n5945), .ZN(n5264) );
  OAI21_X1 U6434 ( .B1(n5607), .B2(n6029), .A(n5264), .ZN(n5273) );
  INV_X1 U6435 ( .A(n5265), .ZN(n5266) );
  NOR2_X1 U6436 ( .A1(n5267), .A2(n5266), .ZN(n5956) );
  INV_X1 U6437 ( .A(n5956), .ZN(n5268) );
  NAND2_X1 U6438 ( .A1(n5269), .A2(n5268), .ZN(n5954) );
  AOI22_X1 U6439 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6034), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5954), .ZN(n5270) );
  OAI211_X1 U6440 ( .C1(n6005), .C2(n5271), .A(n5270), .B(n5994), .ZN(n5272)
         );
  AOI211_X1 U6441 ( .C1(n5891), .C2(n6041), .A(n5273), .B(n5272), .ZN(n5274)
         );
  OAI21_X1 U6442 ( .B1(n5611), .B2(n6009), .A(n5274), .ZN(U2812) );
  OAI22_X1 U6443 ( .A1(n5276), .A2(n6045), .B1(n5275), .B2(n6055), .ZN(n5277)
         );
  INV_X1 U6444 ( .A(n5277), .ZN(n5278) );
  OAI21_X1 U6445 ( .B1(n5611), .B2(n5487), .A(n5278), .ZN(U2844) );
  AOI22_X1 U6446 ( .A1(n5279), .A2(DATAI_15_), .B1(n6065), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U6447 ( .B1(n5611), .B2(n5843), .A(n5280), .ZN(U2876) );
  INV_X1 U6448 ( .A(n5311), .ZN(n5281) );
  NOR2_X1 U6449 ( .A1(n5315), .A2(n5281), .ZN(n5759) );
  XNOR2_X1 U6450 ( .A(n4408), .B(n2996), .ZN(n5282) );
  NOR2_X1 U6451 ( .A1(n5759), .A2(n5282), .ZN(n5286) );
  XNOR2_X1 U6452 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5284) );
  INV_X1 U6453 ( .A(n5282), .ZN(n5283) );
  OAI22_X1 U6454 ( .A1(n6433), .A2(n5284), .B1(n5771), .B2(n5283), .ZN(n5285)
         );
  AOI211_X1 U6455 ( .C1(n4317), .C2(n5758), .A(n5286), .B(n5285), .ZN(n6440)
         );
  INV_X1 U6456 ( .A(n6440), .ZN(n5292) );
  NOR3_X1 U6457 ( .A1(n6465), .A2(n5288), .A3(n5287), .ZN(n5291) );
  INV_X1 U6458 ( .A(n4408), .ZN(n5289) );
  NOR3_X1 U6459 ( .A1(n5778), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5289), 
        .ZN(n5290) );
  AOI211_X1 U6460 ( .C1(n5292), .C2(n5777), .A(n5291), .B(n5290), .ZN(n5295)
         );
  OAI21_X1 U6461 ( .B1(n5299), .B2(n5293), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n5294) );
  OAI21_X1 U6462 ( .B1(n5295), .B2(n5299), .A(n5294), .ZN(U3459) );
  AOI21_X1 U6463 ( .B1(n5777), .B2(n5769), .A(n5299), .ZN(n5301) );
  OAI22_X1 U6464 ( .A1(n3862), .A2(n5297), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5296), .ZN(n6431) );
  OAI22_X1 U6465 ( .A1(n5778), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6465), .ZN(n5298) );
  AOI21_X1 U6466 ( .B1(n5777), .B2(n6431), .A(n5298), .ZN(n5300) );
  OAI22_X1 U6467 ( .A1(n5301), .A2(n3047), .B1(n5300), .B2(n5299), .ZN(U3461)
         );
  INV_X1 U6468 ( .A(n5302), .ZN(n5338) );
  AOI22_X1 U6469 ( .A1(n6062), .A2(DATAI_29_), .B1(n6065), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6470 ( .A1(n6066), .A2(DATAI_13_), .ZN(n5303) );
  OAI211_X1 U6471 ( .C1(n5302), .C2(n5843), .A(n5304), .B(n5303), .ZN(U2862)
         );
  INV_X1 U6472 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5341) );
  INV_X1 U6473 ( .A(n5305), .ZN(n5306) );
  OAI211_X1 U6474 ( .C1(n5461), .C2(n5307), .A(n5351), .B(n5306), .ZN(n5308)
         );
  NAND2_X1 U6475 ( .A1(n5309), .A2(n5308), .ZN(n5630) );
  OAI222_X1 U6476 ( .A1(n5469), .A2(n5302), .B1(n5341), .B2(n6055), .C1(n5630), 
        .C2(n6045), .ZN(U2830) );
  NAND3_X1 U6477 ( .A1(n5311), .A2(n6455), .A3(n5310), .ZN(n5313) );
  AOI22_X1 U6478 ( .A1(n5314), .A2(n5313), .B1(n3597), .B2(n5312), .ZN(n5317)
         );
  INV_X1 U6479 ( .A(n5314), .ZN(n5320) );
  NAND2_X1 U6480 ( .A1(n5320), .A2(n5315), .ZN(n5316) );
  AND2_X1 U6481 ( .A1(n5317), .A2(n5316), .ZN(n6454) );
  INV_X1 U6482 ( .A(n6454), .ZN(n5322) );
  OAI22_X1 U6483 ( .A1(n5320), .A2(n5319), .B1(n4280), .B2(n5318), .ZN(n5915)
         );
  AOI21_X1 U6484 ( .B1(n5321), .B2(n6495), .A(READY_N), .ZN(n6572) );
  NOR2_X1 U6485 ( .A1(n5915), .A2(n6572), .ZN(n6453) );
  NOR2_X1 U6486 ( .A1(n6453), .A2(n6477), .ZN(n5920) );
  MUX2_X1 U6487 ( .A(MORE_REG_SCAN_IN), .B(n5322), .S(n5920), .Z(U3471) );
  INV_X1 U6488 ( .A(n5327), .ZN(n5323) );
  AOI21_X1 U6489 ( .B1(n5325), .B2(n5324), .A(n5323), .ZN(n5330) );
  AOI211_X1 U6490 ( .C1(n5461), .C2(n5351), .A(n5327), .B(n5326), .ZN(n5328)
         );
  AOI21_X1 U6491 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(n5627) );
  NOR3_X1 U6492 ( .A1(n5346), .A2(REIP_REG_30__SCAN_IN), .A3(n6549), .ZN(n5336) );
  OAI22_X1 U6493 ( .A1(n5331), .A2(n6005), .B1(n6029), .B2(n5513), .ZN(n5332)
         );
  AOI21_X1 U6494 ( .B1(EBX_REG_30__SCAN_IN), .B2(n6034), .A(n5332), .ZN(n5333)
         );
  OAI21_X1 U6495 ( .B1(n5334), .B2(n6587), .A(n5333), .ZN(n5335) );
  AOI211_X1 U6496 ( .C1(n5627), .C2(n6041), .A(n5336), .B(n5335), .ZN(n5337)
         );
  OAI21_X1 U6497 ( .B1(n5416), .B2(n6009), .A(n5337), .ZN(U2797) );
  NAND2_X1 U6498 ( .A1(n5338), .A2(n6026), .ZN(n5345) );
  AOI22_X1 U6499 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6031), .B1(n6032), 
        .B2(n5339), .ZN(n5340) );
  OAI21_X1 U6500 ( .B1(n6016), .B2(n5341), .A(n5340), .ZN(n5343) );
  NOR2_X1 U6501 ( .A1(n5630), .A2(n6024), .ZN(n5342) );
  AOI211_X1 U6502 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5354), .A(n5343), .B(n5342), .ZN(n5344) );
  OAI211_X1 U6503 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5346), .A(n5345), .B(n5344), .ZN(U2798) );
  AOI21_X1 U6504 ( .B1(n5348), .B2(n5347), .A(n4221), .ZN(n5525) );
  INV_X1 U6505 ( .A(n5525), .ZN(n5496) );
  INV_X1 U6506 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6692) );
  OR2_X1 U6507 ( .A1(n5364), .A2(n5349), .ZN(n5350) );
  NAND2_X1 U6508 ( .A1(n5351), .A2(n5350), .ZN(n5646) );
  OAI22_X1 U6509 ( .A1(n5352), .A2(n6005), .B1(n6029), .B2(n5523), .ZN(n5353)
         );
  AOI21_X1 U6510 ( .B1(n6034), .B2(EBX_REG_28__SCAN_IN), .A(n5353), .ZN(n5356)
         );
  NAND2_X1 U6511 ( .A1(n5354), .A2(REIP_REG_28__SCAN_IN), .ZN(n5355) );
  OAI211_X1 U6512 ( .C1(n5646), .C2(n6024), .A(n5356), .B(n5355), .ZN(n5357)
         );
  AOI21_X1 U6513 ( .B1(n5358), .B2(n6692), .A(n5357), .ZN(n5359) );
  OAI21_X1 U6514 ( .B1(n5496), .B2(n6009), .A(n5359), .ZN(U2799) );
  OAI21_X2 U6515 ( .B1(n5360), .B2(n5361), .A(n5347), .ZN(n5531) );
  AND2_X1 U6516 ( .A1(n3023), .A2(n5362), .ZN(n5363) );
  OR2_X1 U6517 ( .A1(n5364), .A2(n5363), .ZN(n5652) );
  AOI22_X1 U6518 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6034), .B1(n5534), .B2(n6032), .ZN(n5365) );
  OAI21_X1 U6519 ( .B1(n5530), .B2(n6005), .A(n5365), .ZN(n5366) );
  AOI21_X1 U6520 ( .B1(n5373), .B2(REIP_REG_27__SCAN_IN), .A(n5366), .ZN(n5370) );
  INV_X1 U6521 ( .A(n5788), .ZN(n5368) );
  INV_X1 U6522 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6706) );
  NAND3_X1 U6523 ( .A1(n5368), .A2(n6706), .A3(n5367), .ZN(n5369) );
  OAI211_X1 U6524 ( .C1(n5652), .C2(n6024), .A(n5370), .B(n5369), .ZN(n5371)
         );
  INV_X1 U6525 ( .A(n5371), .ZN(n5372) );
  OAI21_X1 U6526 ( .B1(n5531), .B2(n6009), .A(n5372), .ZN(U2800) );
  INV_X1 U6527 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U6528 ( .A1(n6739), .A2(n5788), .ZN(n5784) );
  AOI21_X1 U6529 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5784), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5384) );
  INV_X1 U6530 ( .A(n5373), .ZN(n5383) );
  AOI21_X1 U6531 ( .B1(n5375), .B2(n5374), .A(n5360), .ZN(n5540) );
  NAND2_X1 U6532 ( .A1(n5540), .A2(n6026), .ZN(n5382) );
  INV_X1 U6533 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5376) );
  OAI22_X1 U6534 ( .A1(n5376), .A2(n6005), .B1(n6029), .B2(n5538), .ZN(n5380)
         );
  OR2_X1 U6535 ( .A1(n5426), .A2(n5377), .ZN(n5378) );
  NAND2_X1 U6536 ( .A1(n3023), .A2(n5378), .ZN(n5662) );
  NOR2_X1 U6537 ( .A1(n5662), .A2(n6024), .ZN(n5379) );
  AOI211_X1 U6538 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6034), .A(n5380), .B(n5379), 
        .ZN(n5381) );
  OAI211_X1 U6539 ( .C1(n5384), .C2(n5383), .A(n5382), .B(n5381), .ZN(U2801)
         );
  NOR2_X1 U6540 ( .A1(n5386), .A2(n5387), .ZN(n5388) );
  OR2_X1 U6541 ( .A1(n5385), .A2(n5388), .ZN(n5568) );
  INV_X1 U6542 ( .A(n5811), .ZN(n5822) );
  NAND2_X1 U6543 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5810) );
  INV_X1 U6544 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6540) );
  OAI21_X1 U6545 ( .B1(n5822), .B2(n5810), .A(n6540), .ZN(n5395) );
  NOR2_X1 U6546 ( .A1(n5403), .A2(n5389), .ZN(n5793) );
  NAND2_X1 U6547 ( .A1(n3018), .A2(n5390), .ZN(n5391) );
  NAND2_X1 U6548 ( .A1(n5431), .A2(n5391), .ZN(n5685) );
  OAI22_X1 U6549 ( .A1(n5435), .A2(n6016), .B1(n5567), .B2(n6005), .ZN(n5392)
         );
  AOI21_X1 U6550 ( .B1(n6032), .B2(n5571), .A(n5392), .ZN(n5393) );
  OAI21_X1 U6551 ( .B1(n5685), .B2(n6024), .A(n5393), .ZN(n5394) );
  AOI21_X1 U6552 ( .B1(n5395), .B2(n5793), .A(n5394), .ZN(n5396) );
  OAI21_X1 U6553 ( .B1(n5568), .B2(n6009), .A(n5396), .ZN(U2804) );
  INV_X1 U6554 ( .A(n5399), .ZN(n5400) );
  AOI21_X1 U6555 ( .B1(n5401), .B2(n5398), .A(n5400), .ZN(n6059) );
  INV_X1 U6556 ( .A(n6059), .ZN(n5481) );
  NOR2_X1 U6557 ( .A1(n5403), .A2(n5402), .ZN(n5938) );
  NAND2_X1 U6558 ( .A1(n6533), .A2(n5404), .ZN(n5408) );
  OAI22_X1 U6559 ( .A1(n5406), .A2(n6016), .B1(n5405), .B2(n6005), .ZN(n5407)
         );
  AOI211_X1 U6560 ( .C1(n5938), .C2(n5408), .A(n6021), .B(n5407), .ZN(n5412)
         );
  INV_X1 U6561 ( .A(n5473), .ZN(n5409) );
  AOI21_X1 U6562 ( .B1(n5410), .B2(n5485), .A(n5409), .ZN(n5882) );
  AOI22_X1 U6563 ( .A1(n5882), .A2(n6041), .B1(n6032), .B2(n5867), .ZN(n5411)
         );
  OAI211_X1 U6564 ( .C1(n5481), .C2(n6009), .A(n5412), .B(n5411), .ZN(U2810)
         );
  OAI22_X1 U6565 ( .A1(n5414), .A2(n6045), .B1(n6055), .B2(n5413), .ZN(U2828)
         );
  AOI22_X1 U6566 ( .A1(n5627), .A2(n6051), .B1(EBX_REG_30__SCAN_IN), .B2(n5479), .ZN(n5415) );
  OAI21_X1 U6567 ( .B1(n5416), .B2(n5487), .A(n5415), .ZN(U2829) );
  INV_X1 U6568 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5417) );
  OAI222_X1 U6569 ( .A1(n5469), .A2(n5496), .B1(n5417), .B2(n6055), .C1(n5646), 
        .C2(n6045), .ZN(U2831) );
  INV_X1 U6570 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5418) );
  OAI222_X1 U6571 ( .A1(n5469), .A2(n5531), .B1(n5418), .B2(n6055), .C1(n5652), 
        .C2(n6045), .ZN(U2832) );
  INV_X1 U6572 ( .A(n5540), .ZN(n5501) );
  INV_X1 U6573 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5419) );
  OAI222_X1 U6574 ( .A1(n5469), .A2(n5501), .B1(n5419), .B2(n6055), .C1(n5662), 
        .C2(n6045), .ZN(U2833) );
  NAND2_X1 U6575 ( .A1(n5421), .A2(n5422), .ZN(n5423) );
  AND2_X1 U6576 ( .A1(n5374), .A2(n5423), .ZN(n5844) );
  INV_X1 U6577 ( .A(n5844), .ZN(n5428) );
  NOR2_X1 U6578 ( .A1(n5432), .A2(n5424), .ZN(n5425) );
  OR2_X1 U6579 ( .A1(n5426), .A2(n5425), .ZN(n5786) );
  OAI222_X1 U6580 ( .A1(n5428), .A2(n5487), .B1(n5427), .B2(n6055), .C1(n6045), 
        .C2(n5786), .ZN(U2834) );
  OAI21_X1 U6581 ( .B1(n5385), .B2(n5429), .A(n5421), .ZN(n5798) );
  INV_X1 U6582 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5434) );
  AND2_X1 U6583 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  OR2_X1 U6584 ( .A1(n5433), .A2(n5432), .ZN(n5802) );
  OAI222_X1 U6585 ( .A1(n5469), .A2(n5798), .B1(n6055), .B2(n5434), .C1(n5802), 
        .C2(n6045), .ZN(U2835) );
  OAI22_X1 U6586 ( .A1(n5685), .A2(n6045), .B1(n5435), .B2(n6055), .ZN(n5436)
         );
  INV_X1 U6587 ( .A(n5436), .ZN(n5437) );
  OAI21_X1 U6588 ( .B1(n5568), .B2(n5469), .A(n5437), .ZN(U2836) );
  AOI21_X1 U6589 ( .B1(n5439), .B2(n5438), .A(n5386), .ZN(n5847) );
  INV_X1 U6590 ( .A(n5847), .ZN(n5443) );
  INV_X1 U6591 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6592 ( .A1(n3022), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6593 ( .A1(n3018), .A2(n5441), .ZN(n5814) );
  OAI222_X1 U6594 ( .A1(n5469), .A2(n5443), .B1(n6055), .B2(n5442), .C1(n5814), 
        .C2(n6045), .ZN(U2837) );
  INV_X1 U6595 ( .A(n5438), .ZN(n5445) );
  AOI21_X1 U6596 ( .B1(n5446), .B2(n5444), .A(n5445), .ZN(n5850) );
  INV_X1 U6597 ( .A(n5850), .ZN(n5451) );
  INV_X1 U6598 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5450) );
  OR2_X1 U6599 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6600 ( .A1(n3022), .A2(n5449), .ZN(n5818) );
  OAI222_X1 U6601 ( .A1(n5451), .A2(n5487), .B1(n5450), .B2(n6055), .C1(n6045), 
        .C2(n5818), .ZN(U2838) );
  OAI21_X1 U6602 ( .B1(n5452), .B2(n5453), .A(n5444), .ZN(n5589) );
  MUX2_X1 U6603 ( .A(n5463), .B(n5454), .S(n3024), .Z(n5456) );
  XNOR2_X1 U6604 ( .A(n5456), .B(n5455), .ZN(n5829) );
  AOI22_X1 U6605 ( .A1(n5829), .A2(n6051), .B1(EBX_REG_20__SCAN_IN), .B2(n5479), .ZN(n5457) );
  OAI21_X1 U6606 ( .B1(n5589), .B2(n5469), .A(n5457), .ZN(U2839) );
  AND2_X1 U6607 ( .A1(n5458), .A2(n5459), .ZN(n5460) );
  OR2_X1 U6608 ( .A1(n5460), .A2(n5452), .ZN(n5837) );
  MUX2_X1 U6609 ( .A(n5463), .B(n5462), .S(n5461), .Z(n5472) );
  OR2_X1 U6610 ( .A1(n3024), .A2(n5472), .ZN(n5466) );
  OR2_X1 U6611 ( .A1(n5473), .A2(n5472), .ZN(n5475) );
  NAND2_X1 U6612 ( .A1(n5475), .A2(n5464), .ZN(n5465) );
  NAND2_X1 U6613 ( .A1(n5466), .A2(n5465), .ZN(n5836) );
  OAI22_X1 U6614 ( .A1(n5836), .A2(n6045), .B1(n5842), .B2(n6055), .ZN(n5467)
         );
  INV_X1 U6615 ( .A(n5467), .ZN(n5468) );
  OAI21_X1 U6616 ( .B1(n5837), .B2(n5469), .A(n5468), .ZN(U2840) );
  NAND2_X1 U6617 ( .A1(n5399), .A2(n5470), .ZN(n5471) );
  INV_X1 U6618 ( .A(n6056), .ZN(n5478) );
  NAND2_X1 U6619 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  INV_X1 U6620 ( .A(n5939), .ZN(n5476) );
  OAI222_X1 U6621 ( .A1(n5478), .A2(n5487), .B1(n5477), .B2(n6055), .C1(n6045), 
        .C2(n5476), .ZN(U2841) );
  AOI22_X1 U6622 ( .A1(n5882), .A2(n6051), .B1(EBX_REG_17__SCAN_IN), .B2(n5479), .ZN(n5480) );
  OAI21_X1 U6623 ( .B1(n5481), .B2(n5487), .A(n5480), .ZN(U2842) );
  OAI21_X1 U6624 ( .B1(n3012), .B2(n5482), .A(n5398), .ZN(n5949) );
  INV_X1 U6625 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5486) );
  OR2_X1 U6626 ( .A1(n3029), .A2(n5483), .ZN(n5484) );
  NAND2_X1 U6627 ( .A1(n5485), .A2(n5484), .ZN(n5953) );
  OAI222_X1 U6628 ( .A1(n5949), .A2(n5487), .B1(n5486), .B2(n6055), .C1(n6045), 
        .C2(n5953), .ZN(U2843) );
  NAND2_X1 U6629 ( .A1(n5491), .A2(n5490), .ZN(n5493) );
  AOI22_X1 U6630 ( .A1(n6062), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6065), .ZN(n5492) );
  NAND2_X1 U6631 ( .A1(n5493), .A2(n5492), .ZN(U2860) );
  AOI22_X1 U6632 ( .A1(n6062), .A2(DATAI_28_), .B1(n6065), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6633 ( .A1(n6066), .A2(DATAI_12_), .ZN(n5494) );
  OAI211_X1 U6634 ( .C1(n5496), .C2(n5843), .A(n5495), .B(n5494), .ZN(U2863)
         );
  AOI22_X1 U6635 ( .A1(n6062), .A2(DATAI_27_), .B1(n6065), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6636 ( .A1(n6066), .A2(DATAI_11_), .ZN(n5497) );
  OAI211_X1 U6637 ( .C1(n5531), .C2(n5843), .A(n5498), .B(n5497), .ZN(U2864)
         );
  AOI22_X1 U6638 ( .A1(n6062), .A2(DATAI_26_), .B1(n6065), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6639 ( .A1(n6066), .A2(DATAI_10_), .ZN(n5499) );
  OAI211_X1 U6640 ( .C1(n5501), .C2(n5843), .A(n5500), .B(n5499), .ZN(U2865)
         );
  AOI22_X1 U6641 ( .A1(n6062), .A2(DATAI_24_), .B1(n6065), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6642 ( .A1(n6066), .A2(DATAI_8_), .ZN(n5502) );
  OAI211_X1 U6643 ( .C1(n5798), .C2(n5843), .A(n5503), .B(n5502), .ZN(U2867)
         );
  AOI22_X1 U6644 ( .A1(n6062), .A2(DATAI_23_), .B1(n6065), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6645 ( .A1(n6066), .A2(DATAI_7_), .ZN(n5504) );
  OAI211_X1 U6646 ( .C1(n5568), .C2(n5843), .A(n5505), .B(n5504), .ZN(U2868)
         );
  AOI22_X1 U6647 ( .A1(n6062), .A2(DATAI_19_), .B1(n6065), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6648 ( .A1(n6066), .A2(DATAI_3_), .ZN(n5506) );
  OAI211_X1 U6649 ( .C1(n5837), .C2(n5843), .A(n5507), .B(n5506), .ZN(U2872)
         );
  NAND2_X1 U6650 ( .A1(n5508), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5509) );
  OAI21_X1 U6651 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5510), .A(n5509), 
        .ZN(n5511) );
  XNOR2_X1 U6652 ( .A(n5511), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5629)
         );
  NAND2_X1 U6653 ( .A1(n6213), .A2(REIP_REG_30__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U6654 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5512)
         );
  OAI211_X1 U6655 ( .C1(n6139), .C2(n5513), .A(n5623), .B(n5512), .ZN(n5514)
         );
  AOI21_X1 U6656 ( .B1(n5515), .B2(n6133), .A(n5514), .ZN(n5516) );
  OAI21_X1 U6657 ( .B1(n5629), .B2(n6124), .A(n5516), .ZN(U2956) );
  NAND3_X1 U6658 ( .A1(n4224), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3512), .ZN(n5520) );
  NOR2_X1 U6659 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U6660 ( .A1(n5857), .A2(n5658), .ZN(n5518) );
  OR2_X1 U6661 ( .A1(n5517), .A2(n5518), .ZN(n5527) );
  AOI22_X1 U6662 ( .A1(n5520), .A2(n5527), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5519), .ZN(n5521) );
  XNOR2_X1 U6663 ( .A(n5521), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5649)
         );
  NAND2_X1 U6664 ( .A1(n6213), .A2(REIP_REG_28__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6665 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5522)
         );
  OAI211_X1 U6666 ( .C1(n6139), .C2(n5523), .A(n5639), .B(n5522), .ZN(n5524)
         );
  AOI21_X1 U6667 ( .B1(n5525), .B2(n6133), .A(n5524), .ZN(n5526) );
  OAI21_X1 U6668 ( .B1(n6124), .B2(n5649), .A(n5526), .ZN(U2958) );
  NAND2_X1 U6669 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U6670 ( .A(n5529), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5657)
         );
  NAND2_X1 U6671 ( .A1(n6213), .A2(REIP_REG_27__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U6672 ( .B1(n5616), .B2(n5530), .A(n5651), .ZN(n5533) );
  NOR2_X1 U6673 ( .A1(n5531), .A2(n6122), .ZN(n5532) );
  AOI211_X2 U6674 ( .C1(n5534), .C2(n6109), .A(n5533), .B(n5532), .ZN(n5535)
         );
  OAI21_X1 U6675 ( .B1(n5657), .B2(n6124), .A(n5535), .ZN(U2959) );
  XNOR2_X1 U6676 ( .A(n3512), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5536)
         );
  XNOR2_X1 U6677 ( .A(n4224), .B(n5536), .ZN(n5666) );
  NAND2_X1 U6678 ( .A1(n6213), .A2(REIP_REG_26__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U6679 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5537)
         );
  OAI211_X1 U6680 ( .C1(n6139), .C2(n5538), .A(n5661), .B(n5537), .ZN(n5539)
         );
  AOI21_X1 U6681 ( .B1(n5540), .B2(n6133), .A(n5539), .ZN(n5541) );
  OAI21_X1 U6682 ( .B1(n6124), .B2(n5666), .A(n5541), .ZN(U2960) );
  AOI21_X1 U6683 ( .B1(n5543), .B2(n5517), .A(n5542), .ZN(n5673) );
  INV_X1 U6684 ( .A(n5785), .ZN(n5545) );
  NAND2_X1 U6685 ( .A1(n6213), .A2(REIP_REG_25__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6686 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5544)
         );
  OAI211_X1 U6687 ( .C1(n6139), .C2(n5545), .A(n5668), .B(n5544), .ZN(n5546)
         );
  AOI21_X1 U6688 ( .B1(n5844), .B2(n6133), .A(n5546), .ZN(n5547) );
  OAI21_X1 U6689 ( .B1(n5673), .B2(n6124), .A(n5547), .ZN(U2961) );
  INV_X1 U6690 ( .A(n5548), .ZN(n5594) );
  NAND2_X1 U6691 ( .A1(n5594), .A2(n5721), .ZN(n5593) );
  OAI21_X1 U6692 ( .B1(n5549), .B2(n5721), .A(n3512), .ZN(n5550) );
  NAND2_X1 U6693 ( .A1(n5593), .A2(n5550), .ZN(n5587) );
  INV_X1 U6694 ( .A(n5587), .ZN(n5553) );
  INV_X1 U6695 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5551) );
  XNOR2_X1 U6696 ( .A(n3512), .B(n5551), .ZN(n5586) );
  NAND2_X1 U6697 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5554) );
  NAND2_X2 U6698 ( .A1(n5563), .A2(n5554), .ZN(n5580) );
  INV_X1 U6699 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U6700 ( .A(n3512), .B(n5555), .ZN(n5581) );
  NOR2_X2 U6701 ( .A1(n5580), .A2(n5581), .ZN(n5579) );
  INV_X1 U6702 ( .A(n5579), .ZN(n5556) );
  OAI21_X1 U6703 ( .B1(n5857), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5556), 
        .ZN(n5575) );
  NAND3_X1 U6704 ( .A1(n3512), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5557) );
  NOR2_X1 U6705 ( .A1(n3512), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5573)
         );
  NAND2_X1 U6706 ( .A1(n5579), .A2(n5573), .ZN(n5564) );
  XNOR2_X1 U6707 ( .A(n5558), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5683)
         );
  INV_X1 U6708 ( .A(n5798), .ZN(n5561) );
  NAND2_X1 U6709 ( .A1(n6213), .A2(REIP_REG_24__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6710 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5559)
         );
  OAI211_X1 U6711 ( .C1(n6139), .C2(n5795), .A(n5679), .B(n5559), .ZN(n5560)
         );
  AOI21_X1 U6712 ( .B1(n5561), .B2(n6133), .A(n5560), .ZN(n5562) );
  OAI21_X1 U6713 ( .B1(n5683), .B2(n6124), .A(n5562), .ZN(U2962) );
  OAI21_X1 U6714 ( .B1(n5563), .B2(n5565), .A(n5564), .ZN(n5566) );
  XNOR2_X1 U6715 ( .A(n5566), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5691)
         );
  NAND2_X1 U6716 ( .A1(n6213), .A2(REIP_REG_23__SCAN_IN), .ZN(n5684) );
  OAI21_X1 U6717 ( .B1(n5616), .B2(n5567), .A(n5684), .ZN(n5570) );
  NOR2_X1 U6718 ( .A1(n5568), .A2(n6122), .ZN(n5569) );
  AOI211_X1 U6719 ( .C1(n6109), .C2(n5571), .A(n5570), .B(n5569), .ZN(n5572)
         );
  OAI21_X1 U6720 ( .B1(n5691), .B2(n6124), .A(n5572), .ZN(U2963) );
  AOI21_X1 U6721 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3512), .A(n5573), 
        .ZN(n5574) );
  XNOR2_X1 U6722 ( .A(n5575), .B(n5574), .ZN(n5699) );
  NAND2_X1 U6723 ( .A1(n6213), .A2(REIP_REG_22__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6724 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5576)
         );
  OAI211_X1 U6725 ( .C1(n6139), .C2(n5804), .A(n5693), .B(n5576), .ZN(n5577)
         );
  AOI21_X1 U6726 ( .B1(n5847), .B2(n6133), .A(n5577), .ZN(n5578) );
  OAI21_X1 U6727 ( .B1(n5699), .B2(n6124), .A(n5578), .ZN(U2964) );
  AOI21_X1 U6728 ( .B1(n5581), .B2(n5580), .A(n5579), .ZN(n5706) );
  INV_X1 U6729 ( .A(n5817), .ZN(n5583) );
  NAND2_X1 U6730 ( .A1(n6129), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5582)
         );
  NAND2_X1 U6731 ( .A1(n6213), .A2(REIP_REG_21__SCAN_IN), .ZN(n5700) );
  OAI211_X1 U6732 ( .C1(n6139), .C2(n5583), .A(n5582), .B(n5700), .ZN(n5584)
         );
  AOI21_X1 U6733 ( .B1(n5850), .B2(n6133), .A(n5584), .ZN(n5585) );
  OAI21_X1 U6734 ( .B1(n5706), .B2(n6124), .A(n5585), .ZN(U2965) );
  NAND2_X1 U6735 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  NAND2_X1 U6736 ( .A1(n5563), .A2(n5588), .ZN(n5720) );
  INV_X1 U6737 ( .A(n5589), .ZN(n5853) );
  AND2_X1 U6738 ( .A1(n6199), .A2(REIP_REG_20__SCAN_IN), .ZN(n5709) );
  AOI21_X1 U6739 ( .B1(n6129), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5709), 
        .ZN(n5590) );
  OAI21_X1 U6740 ( .B1(n5825), .B2(n6139), .A(n5590), .ZN(n5591) );
  AOI21_X1 U6741 ( .B1(n5853), .B2(n6133), .A(n5591), .ZN(n5592) );
  OAI21_X1 U6742 ( .B1(n5720), .B2(n6124), .A(n5592), .ZN(U2966) );
  OAI21_X1 U6743 ( .B1(n5594), .B2(n5721), .A(n5593), .ZN(n5595) );
  XNOR2_X1 U6744 ( .A(n5595), .B(n3512), .ZN(n5728) );
  NAND2_X1 U6745 ( .A1(n6213), .A2(REIP_REG_19__SCAN_IN), .ZN(n5723) );
  OAI21_X1 U6746 ( .B1(n5616), .B2(n5834), .A(n5723), .ZN(n5597) );
  NOR2_X1 U6747 ( .A1(n5837), .A2(n6122), .ZN(n5596) );
  AOI211_X1 U6748 ( .C1(n6109), .C2(n5839), .A(n5597), .B(n5596), .ZN(n5598)
         );
  OAI21_X1 U6749 ( .B1(n6124), .B2(n5728), .A(n5598), .ZN(U2967) );
  XNOR2_X1 U6750 ( .A(n3512), .B(n5856), .ZN(n5600) );
  XNOR2_X1 U6751 ( .A(n5599), .B(n5600), .ZN(n5735) );
  INV_X1 U6752 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U6753 ( .A1(n6213), .A2(REIP_REG_16__SCAN_IN), .ZN(n5729) );
  OAI21_X1 U6754 ( .B1(n5616), .B2(n5601), .A(n5729), .ZN(n5603) );
  NOR2_X1 U6755 ( .A1(n5949), .A2(n6122), .ZN(n5602) );
  AOI211_X1 U6756 ( .C1(n6109), .C2(n5950), .A(n5603), .B(n5602), .ZN(n5604)
         );
  OAI21_X1 U6757 ( .B1(n6124), .B2(n5735), .A(n5604), .ZN(U2970) );
  XNOR2_X1 U6758 ( .A(n3512), .B(n5898), .ZN(n5606) );
  XNOR2_X1 U6759 ( .A(n5605), .B(n5606), .ZN(n5895) );
  NAND2_X1 U6760 ( .A1(n5895), .A2(n6135), .ZN(n5610) );
  AND2_X1 U6761 ( .A1(n6199), .A2(REIP_REG_15__SCAN_IN), .ZN(n5890) );
  NOR2_X1 U6762 ( .A1(n6139), .A2(n5607), .ZN(n5608) );
  AOI211_X1 U6763 ( .C1(n6129), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5890), 
        .B(n5608), .ZN(n5609) );
  OAI211_X1 U6764 ( .C1(n6122), .C2(n5611), .A(n5610), .B(n5609), .ZN(U2971)
         );
  XNOR2_X1 U6765 ( .A(n3512), .B(n5613), .ZN(n5614) );
  XNOR2_X1 U6766 ( .A(n5612), .B(n5614), .ZN(n5750) );
  INV_X1 U6767 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U6768 ( .A1(n6213), .A2(REIP_REG_14__SCAN_IN), .ZN(n5737) );
  OAI21_X1 U6769 ( .B1(n5616), .B2(n5615), .A(n5737), .ZN(n5618) );
  NOR2_X1 U6770 ( .A1(n5958), .A2(n6122), .ZN(n5617) );
  AOI211_X1 U6771 ( .C1(n6109), .C2(n5959), .A(n5618), .B(n5617), .ZN(n5619)
         );
  OAI21_X1 U6772 ( .B1(n6124), .B2(n5750), .A(n5619), .ZN(U2972) );
  INV_X1 U6773 ( .A(n5620), .ZN(n5625) );
  NAND2_X1 U6774 ( .A1(n5621), .A2(n5624), .ZN(n5622) );
  OAI211_X1 U6775 ( .C1(n5625), .C2(n5624), .A(n5623), .B(n5622), .ZN(n5626)
         );
  AOI21_X1 U6776 ( .B1(n5627), .B2(n6223), .A(n5626), .ZN(n5628) );
  OAI21_X1 U6777 ( .B1(n5629), .B2(n6201), .A(n5628), .ZN(U2988) );
  INV_X1 U6778 ( .A(n5630), .ZN(n5636) );
  NOR3_X1 U6779 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5641), 
        .ZN(n5635) );
  OAI21_X1 U6780 ( .B1(n5633), .B2(n5632), .A(n5631), .ZN(n5634) );
  AOI211_X1 U6781 ( .C1(n5636), .C2(n6223), .A(n5635), .B(n5634), .ZN(n5637)
         );
  OAI21_X1 U6782 ( .B1(n5638), .B2(n6201), .A(n5637), .ZN(U2989) );
  INV_X1 U6783 ( .A(n5639), .ZN(n5640) );
  AOI21_X1 U6784 ( .B1(n5655), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5640), 
        .ZN(n5645) );
  INV_X1 U6785 ( .A(n5641), .ZN(n5642) );
  OR3_X1 U6786 ( .A1(n5650), .A2(n5643), .A3(n5642), .ZN(n5644) );
  OAI211_X1 U6787 ( .C1(n5646), .C2(n6193), .A(n5645), .B(n5644), .ZN(n5647)
         );
  INV_X1 U6788 ( .A(n5647), .ZN(n5648) );
  OAI21_X1 U6789 ( .B1(n5649), .B2(n6201), .A(n5648), .ZN(U2990) );
  NOR2_X1 U6790 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5654)
         );
  OAI21_X1 U6791 ( .B1(n5652), .B2(n6193), .A(n5651), .ZN(n5653) );
  AOI211_X1 U6792 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5655), .A(n5654), .B(n5653), .ZN(n5656) );
  OAI21_X1 U6793 ( .B1(n5657), .B2(n6201), .A(n5656), .ZN(U2991) );
  INV_X1 U6794 ( .A(n5671), .ZN(n5660) );
  NOR3_X1 U6795 ( .A1(n5660), .A2(n5659), .A3(n5658), .ZN(n5664) );
  OAI21_X1 U6796 ( .B1(n5662), .B2(n6193), .A(n5661), .ZN(n5663) );
  AOI211_X1 U6797 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5676), .A(n5664), .B(n5663), .ZN(n5665) );
  OAI21_X1 U6798 ( .B1(n5666), .B2(n6201), .A(n5665), .ZN(U2992) );
  NAND2_X1 U6799 ( .A1(n5676), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U6800 ( .C1(n5786), .C2(n6193), .A(n5668), .B(n5667), .ZN(n5669)
         );
  AOI21_X1 U6801 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5672) );
  OAI21_X1 U6802 ( .B1(n5673), .B2(n6201), .A(n5672), .ZN(U2993) );
  INV_X1 U6803 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6804 ( .A1(n5686), .A2(n5674), .ZN(n5678) );
  INV_X1 U6805 ( .A(n5675), .ZN(n5677) );
  NAND3_X1 U6806 ( .A1(n5678), .A2(n5677), .A3(n5676), .ZN(n5680) );
  OAI211_X1 U6807 ( .C1(n5802), .C2(n6193), .A(n5680), .B(n5679), .ZN(n5681)
         );
  INV_X1 U6808 ( .A(n5681), .ZN(n5682) );
  OAI21_X1 U6809 ( .B1(n5683), .B2(n6201), .A(n5682), .ZN(U2994) );
  OAI21_X1 U6810 ( .B1(n5685), .B2(n6193), .A(n5684), .ZN(n5688) );
  NOR2_X1 U6811 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5687)
         );
  AOI211_X1 U6812 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5689), .A(n5688), .B(n5687), .ZN(n5690) );
  OAI21_X1 U6813 ( .B1(n5691), .B2(n6201), .A(n5690), .ZN(U2995) );
  INV_X1 U6814 ( .A(n5692), .ZN(n5704) );
  OAI21_X1 U6815 ( .B1(n5814), .B2(n6193), .A(n5693), .ZN(n5697) );
  NOR3_X1 U6816 ( .A1(n5701), .A2(n5695), .A3(n5694), .ZN(n5696) );
  AOI211_X1 U6817 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5704), .A(n5697), .B(n5696), .ZN(n5698) );
  OAI21_X1 U6818 ( .B1(n5699), .B2(n6201), .A(n5698), .ZN(U2996) );
  OAI21_X1 U6819 ( .B1(n5818), .B2(n6193), .A(n5700), .ZN(n5703) );
  NOR2_X1 U6820 ( .A1(n5701), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5702)
         );
  AOI211_X1 U6821 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5704), .A(n5703), .B(n5702), .ZN(n5705) );
  OAI21_X1 U6822 ( .B1(n5706), .B2(n6201), .A(n5705), .ZN(U2997) );
  NOR2_X1 U6823 ( .A1(n5708), .A2(n5707), .ZN(n5710) );
  AOI21_X1 U6824 ( .B1(n5722), .B2(n5710), .A(n5709), .ZN(n5719) );
  NOR2_X1 U6825 ( .A1(n5711), .A2(n5874), .ZN(n5712) );
  NOR2_X1 U6826 ( .A1(n5717), .A2(n5712), .ZN(n5713) );
  NOR2_X1 U6827 ( .A1(n5714), .A2(n5713), .ZN(n5881) );
  NAND2_X1 U6828 ( .A1(n6156), .A2(n5715), .ZN(n5716) );
  OAI211_X1 U6829 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5717), .A(n5881), .B(n5716), .ZN(n5726) );
  AOI22_X1 U6830 ( .A1(n5726), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n5829), .B2(n6223), .ZN(n5718) );
  OAI211_X1 U6831 ( .C1(n5720), .C2(n6201), .A(n5719), .B(n5718), .ZN(U2998)
         );
  NAND2_X1 U6832 ( .A1(n5722), .A2(n5721), .ZN(n5724) );
  OAI211_X1 U6833 ( .C1(n6193), .C2(n5836), .A(n5724), .B(n5723), .ZN(n5725)
         );
  AOI21_X1 U6834 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5726), .A(n5725), 
        .ZN(n5727) );
  OAI21_X1 U6835 ( .B1(n5728), .B2(n6201), .A(n5727), .ZN(U2999) );
  AOI211_X1 U6836 ( .C1(n5898), .C2(n5856), .A(n5893), .B(n5892), .ZN(n5732)
         );
  OAI21_X1 U6837 ( .B1(n5953), .B2(n6193), .A(n5729), .ZN(n5731) );
  AOI21_X1 U6838 ( .B1(n5892), .B2(n6221), .A(n6142), .ZN(n5899) );
  NOR2_X1 U6839 ( .A1(n5899), .A2(n5856), .ZN(n5730) );
  AOI211_X1 U6840 ( .C1(n5733), .C2(n5732), .A(n5731), .B(n5730), .ZN(n5734)
         );
  OAI21_X1 U6841 ( .B1(n5735), .B2(n6201), .A(n5734), .ZN(U3002) );
  INV_X1 U6842 ( .A(n5736), .ZN(n5955) );
  NAND2_X1 U6843 ( .A1(n5742), .A2(n6141), .ZN(n5738) );
  OAI21_X1 U6844 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5738), .A(n5737), 
        .ZN(n5739) );
  AOI21_X1 U6845 ( .B1(n5955), .B2(n6223), .A(n5739), .ZN(n5749) );
  AOI21_X1 U6846 ( .B1(n5904), .B2(n5740), .A(n6142), .ZN(n5741) );
  OAI21_X1 U6847 ( .B1(n5742), .B2(n5906), .A(n5741), .ZN(n5908) );
  INV_X1 U6848 ( .A(n5743), .ZN(n5745) );
  NAND3_X1 U6849 ( .A1(n5745), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5744), 
        .ZN(n5746) );
  AOI211_X1 U6850 ( .C1(n5747), .C2(n5746), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5904), .ZN(n5910) );
  OAI21_X1 U6851 ( .B1(n5908), .B2(n5910), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5748) );
  OAI211_X1 U6852 ( .C1(n5750), .C2(n6201), .A(n5749), .B(n5748), .ZN(U3004)
         );
  OAI21_X1 U6853 ( .B1(n2988), .B2(STATEBS16_REG_SCAN_IN), .A(n6365), .ZN(
        n5751) );
  OAI22_X1 U6854 ( .A1(n6364), .A2(n5751), .B1(n4319), .B2(n5756), .ZN(n5752)
         );
  MUX2_X1 U6855 ( .A(n5752), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n6235), 
        .Z(U3464) );
  INV_X1 U6856 ( .A(n6282), .ZN(n5753) );
  NAND2_X1 U6857 ( .A1(n5753), .A2(n6364), .ZN(n6287) );
  NAND3_X1 U6858 ( .A1(n6287), .A2(n6366), .A3(n5754), .ZN(n6239) );
  INV_X1 U6859 ( .A(n6239), .ZN(n5755) );
  MUX2_X1 U6860 ( .A(n5757), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(n6235), 
        .Z(U3462) );
  NAND2_X1 U6861 ( .A1(n4315), .A2(n5758), .ZN(n5776) );
  INV_X1 U6862 ( .A(n5759), .ZN(n5774) );
  MUX2_X1 U6863 ( .A(n5760), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4408), 
        .Z(n5761) );
  NOR2_X1 U6864 ( .A1(n5761), .A2(n4503), .ZN(n5773) );
  INV_X1 U6865 ( .A(n5762), .ZN(n5763) );
  OAI21_X1 U6866 ( .B1(n4408), .B2(n3111), .A(n5763), .ZN(n5765) );
  NOR2_X1 U6867 ( .A1(n5765), .A2(n5764), .ZN(n5779) );
  NAND2_X1 U6868 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5766) );
  INV_X1 U6869 ( .A(n5766), .ZN(n5767) );
  MUX2_X1 U6870 ( .A(n5767), .B(n5766), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5768) );
  NAND2_X1 U6871 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  OAI21_X1 U6872 ( .B1(n5779), .B2(n5771), .A(n5770), .ZN(n5772) );
  AOI21_X1 U6873 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5775) );
  NAND2_X1 U6874 ( .A1(n5776), .A2(n5775), .ZN(n6445) );
  INV_X1 U6875 ( .A(n6445), .ZN(n5781) );
  INV_X1 U6876 ( .A(n5777), .ZN(n5780) );
  OAI22_X1 U6877 ( .A1(n5781), .A2(n5780), .B1(n5779), .B2(n5778), .ZN(n5783)
         );
  MUX2_X1 U6878 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5783), .S(n5782), 
        .Z(U3456) );
  AND2_X1 U6879 ( .A1(n6090), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6880 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6034), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6031), .ZN(n5792) );
  INV_X1 U6881 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U6882 ( .A1(n5785), .A2(n6032), .B1(n5784), .B2(n6745), .ZN(n5791)
         );
  NOR2_X1 U6883 ( .A1(n5786), .A2(n6024), .ZN(n5787) );
  AOI21_X1 U6884 ( .B1(n5844), .B2(n6026), .A(n5787), .ZN(n5790) );
  NOR2_X1 U6885 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5788), .ZN(n5799) );
  OAI21_X1 U6886 ( .B1(n5793), .B2(n5799), .A(REIP_REG_25__SCAN_IN), .ZN(n5789) );
  NAND4_X1 U6887 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(U2802)
         );
  AOI22_X1 U6888 ( .A1(n6031), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(n5793), .ZN(n5794) );
  OAI21_X1 U6889 ( .B1(n6029), .B2(n5795), .A(n5794), .ZN(n5796) );
  AOI21_X1 U6890 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6034), .A(n5796), .ZN(n5797)
         );
  OAI21_X1 U6891 ( .B1(n5798), .B2(n6009), .A(n5797), .ZN(n5800) );
  NOR2_X1 U6892 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  OAI21_X1 U6893 ( .B1(n5802), .B2(n6024), .A(n5801), .ZN(U2803) );
  NAND2_X1 U6894 ( .A1(n5992), .A2(n5803), .ZN(n5823) );
  INV_X1 U6895 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5808) );
  INV_X1 U6896 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5805) );
  OAI22_X1 U6897 ( .A1(n5805), .A2(n6005), .B1(n6029), .B2(n5804), .ZN(n5806)
         );
  AOI21_X1 U6898 ( .B1(n6034), .B2(EBX_REG_22__SCAN_IN), .A(n5806), .ZN(n5807)
         );
  OAI21_X1 U6899 ( .B1(n5823), .B2(n5808), .A(n5807), .ZN(n5809) );
  AOI21_X1 U6900 ( .B1(n5847), .B2(n6026), .A(n5809), .ZN(n5813) );
  OAI211_X1 U6901 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5811), .B(n5810), .ZN(n5812) );
  OAI211_X1 U6902 ( .C1(n6024), .C2(n5814), .A(n5813), .B(n5812), .ZN(U2805)
         );
  INV_X1 U6903 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6697) );
  AOI22_X1 U6904 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6034), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6031), .ZN(n5815) );
  OAI21_X1 U6905 ( .B1(n6697), .B2(n5823), .A(n5815), .ZN(n5816) );
  AOI21_X1 U6906 ( .B1(n5817), .B2(n6032), .A(n5816), .ZN(n5821) );
  INV_X1 U6907 ( .A(n5818), .ZN(n5819) );
  AOI22_X1 U6908 ( .A1(n5850), .A2(n6026), .B1(n6041), .B2(n5819), .ZN(n5820)
         );
  OAI211_X1 U6909 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5822), .A(n5821), .B(n5820), .ZN(U2806) );
  AOI21_X1 U6910 ( .B1(n6703), .B2(n5824), .A(n5823), .ZN(n5828) );
  INV_X1 U6911 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5826) );
  OAI22_X1 U6912 ( .A1(n5826), .A2(n6005), .B1(n5825), .B2(n6029), .ZN(n5827)
         );
  AOI211_X1 U6913 ( .C1(n6034), .C2(EBX_REG_20__SCAN_IN), .A(n5828), .B(n5827), 
        .ZN(n5831) );
  AOI22_X1 U6914 ( .A1(n5853), .A2(n6026), .B1(n6041), .B2(n5829), .ZN(n5830)
         );
  NAND2_X1 U6915 ( .A1(n5831), .A2(n5830), .ZN(U2807) );
  NAND2_X1 U6916 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5832) );
  OAI211_X1 U6917 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5935), .B(n5832), .ZN(n5833) );
  OAI211_X1 U6918 ( .C1(n6005), .C2(n5834), .A(n5833), .B(n5994), .ZN(n5835)
         );
  AOI21_X1 U6919 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5938), .A(n5835), .ZN(n5841) );
  OAI22_X1 U6920 ( .A1(n5837), .A2(n6009), .B1(n6024), .B2(n5836), .ZN(n5838)
         );
  AOI21_X1 U6921 ( .B1(n5839), .B2(n6032), .A(n5838), .ZN(n5840) );
  OAI211_X1 U6922 ( .C1(n5842), .C2(n6016), .A(n5841), .B(n5840), .ZN(U2808)
         );
  AOI22_X1 U6923 ( .A1(n5844), .A2(n6063), .B1(n6062), .B2(DATAI_25_), .ZN(
        n5846) );
  AOI22_X1 U6924 ( .A1(n6066), .A2(DATAI_9_), .B1(n6065), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6925 ( .A1(n5846), .A2(n5845), .ZN(U2866) );
  AOI22_X1 U6926 ( .A1(n5847), .A2(n6063), .B1(n6062), .B2(DATAI_22_), .ZN(
        n5849) );
  AOI22_X1 U6927 ( .A1(n6066), .A2(DATAI_6_), .B1(n6065), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U6928 ( .A1(n5849), .A2(n5848), .ZN(U2869) );
  AOI22_X1 U6929 ( .A1(n5850), .A2(n6063), .B1(n6062), .B2(DATAI_21_), .ZN(
        n5852) );
  AOI22_X1 U6930 ( .A1(n6066), .A2(DATAI_5_), .B1(n6065), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6931 ( .A1(n5852), .A2(n5851), .ZN(U2870) );
  AOI22_X1 U6932 ( .A1(n5853), .A2(n6063), .B1(n6062), .B2(DATAI_20_), .ZN(
        n5855) );
  AOI22_X1 U6933 ( .A1(n6066), .A2(DATAI_4_), .B1(n6065), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6934 ( .A1(n5855), .A2(n5854), .ZN(U2871) );
  AOI22_X1 U6935 ( .A1(n6199), .A2(REIP_REG_18__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5862) );
  NAND3_X1 U6936 ( .A1(n5599), .A2(n5857), .A3(n5856), .ZN(n5863) );
  NOR3_X1 U6937 ( .A1(n5599), .A2(n5857), .A3(n5856), .ZN(n5865) );
  NAND2_X1 U6938 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5858) );
  OAI21_X1 U6939 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5863), .A(n5858), 
        .ZN(n5860) );
  XNOR2_X1 U6940 ( .A(n5860), .B(n5859), .ZN(n5877) );
  AOI22_X1 U6941 ( .A1(n5877), .A2(n6135), .B1(n6133), .B2(n6056), .ZN(n5861)
         );
  OAI211_X1 U6942 ( .C1(n6139), .C2(n5942), .A(n5862), .B(n5861), .ZN(U2968)
         );
  INV_X1 U6943 ( .A(n5863), .ZN(n5864) );
  NOR2_X1 U6944 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  XNOR2_X1 U6945 ( .A(n5866), .B(n5874), .ZN(n5889) );
  AOI22_X1 U6946 ( .A1(n6199), .A2(REIP_REG_17__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5869) );
  AOI22_X1 U6947 ( .A1(n6059), .A2(n6133), .B1(n6109), .B2(n5867), .ZN(n5868)
         );
  OAI211_X1 U6948 ( .C1(n5889), .C2(n6124), .A(n5869), .B(n5868), .ZN(U2969)
         );
  AOI22_X1 U6949 ( .A1(n6199), .A2(REIP_REG_13__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U6950 ( .A(n5871), .B(n5870), .ZN(n5909) );
  AOI22_X1 U6951 ( .A1(n5909), .A2(n6135), .B1(n6133), .B2(n6048), .ZN(n5872)
         );
  OAI211_X1 U6952 ( .C1(n6139), .C2(n5975), .A(n5873), .B(n5872), .ZN(U2973)
         );
  OR2_X1 U6953 ( .A1(n5874), .A2(n5885), .ZN(n5880) );
  OAI21_X1 U6954 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5875), .A(n5881), 
        .ZN(n5876) );
  AOI22_X1 U6955 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5876), .B1(n6199), .B2(REIP_REG_18__SCAN_IN), .ZN(n5879) );
  AOI22_X1 U6956 ( .A1(n5877), .A2(n6229), .B1(n6223), .B2(n5939), .ZN(n5878)
         );
  OAI211_X1 U6957 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5880), .A(n5879), .B(n5878), .ZN(U3000) );
  INV_X1 U6958 ( .A(n5881), .ZN(n5887) );
  NAND2_X1 U6959 ( .A1(n5882), .A2(n6223), .ZN(n5884) );
  NAND2_X1 U6960 ( .A1(n6199), .A2(REIP_REG_17__SCAN_IN), .ZN(n5883) );
  OAI211_X1 U6961 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5885), .A(n5884), .B(n5883), .ZN(n5886) );
  AOI21_X1 U6962 ( .B1(n5887), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5886), 
        .ZN(n5888) );
  OAI21_X1 U6963 ( .B1(n5889), .B2(n6201), .A(n5888), .ZN(U3001) );
  AOI21_X1 U6964 ( .B1(n5891), .B2(n6223), .A(n5890), .ZN(n5897) );
  NOR2_X1 U6965 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  AOI22_X1 U6966 ( .A1(n5895), .A2(n6229), .B1(n5894), .B2(n5898), .ZN(n5896)
         );
  OAI211_X1 U6967 ( .C1(n5899), .C2(n5898), .A(n5897), .B(n5896), .ZN(U3003)
         );
  NOR2_X1 U6968 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  OR2_X1 U6969 ( .A1(n5903), .A2(n5902), .ZN(n6046) );
  INV_X1 U6970 ( .A(n6046), .ZN(n5970) );
  NOR4_X1 U6971 ( .A1(n5906), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5905), 
        .A4(n5904), .ZN(n5907) );
  AOI21_X1 U6972 ( .B1(n5970), .B2(n6223), .A(n5907), .ZN(n5914) );
  AOI22_X1 U6973 ( .A1(n5909), .A2(n6229), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5908), .ZN(n5913) );
  INV_X1 U6974 ( .A(n5910), .ZN(n5912) );
  NAND2_X1 U6975 ( .A1(n6199), .A2(REIP_REG_13__SCAN_IN), .ZN(n5911) );
  NAND4_X1 U6976 ( .A1(n5914), .A2(n5913), .A3(n5912), .A4(n5911), .ZN(U3005)
         );
  INV_X1 U6977 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6498) );
  INV_X1 U6978 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6609) );
  INV_X1 U6979 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6488) );
  AOI221_X1 U6980 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6488), .C2(STATE_REG_0__SCAN_IN), .A(n6581), .ZN(n6556) );
  OAI21_X1 U6981 ( .B1(n6581), .B2(n6609), .A(n6487), .ZN(U2789) );
  OAI21_X1 U6982 ( .B1(n5915), .B2(n6477), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5916) );
  OAI21_X1 U6983 ( .B1(n5917), .B2(n6466), .A(n5916), .ZN(U2790) );
  INV_X1 U6984 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6754) );
  NOR2_X1 U6985 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5919) );
  NOR2_X1 U6986 ( .A1(n6581), .A2(n5919), .ZN(n5918) );
  AOI22_X1 U6987 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6581), .B1(n6754), .B2(
        n5918), .ZN(U2791) );
  OAI21_X1 U6988 ( .B1(BS16_N), .B2(n5919), .A(n6556), .ZN(n6554) );
  OAI21_X1 U6989 ( .B1(n6556), .B2(n6758), .A(n6554), .ZN(U2792) );
  OAI21_X1 U6990 ( .B1(n5920), .B2(n6594), .A(n6124), .ZN(U2793) );
  NOR4_X1 U6991 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5924) );
  NOR4_X1 U6992 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5923) );
  NOR4_X1 U6993 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5922) );
  NOR4_X1 U6994 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5921) );
  NAND4_X1 U6995 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n5930)
         );
  NOR4_X1 U6996 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5928) );
  AOI211_X1 U6997 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5927) );
  NOR4_X1 U6998 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5926) );
  NOR4_X1 U6999 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5925) );
  NAND4_X1 U7000 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n5929)
         );
  NOR2_X1 U7001 ( .A1(n5930), .A2(n5929), .ZN(n6566) );
  INV_X1 U7002 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6685) );
  NOR3_X1 U7003 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5932) );
  OAI21_X1 U7004 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5932), .A(n6566), .ZN(n5931)
         );
  OAI21_X1 U7005 ( .B1(n6566), .B2(n6685), .A(n5931), .ZN(U2794) );
  INV_X1 U7006 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6561) );
  INV_X1 U7007 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6555) );
  AOI21_X1 U7008 ( .B1(n6561), .B2(n6555), .A(n5932), .ZN(n5933) );
  INV_X1 U7009 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6718) );
  INV_X1 U7010 ( .A(n6566), .ZN(n6563) );
  AOI22_X1 U7011 ( .A1(n6566), .A2(n5933), .B1(n6718), .B2(n6563), .ZN(U2795)
         );
  INV_X1 U7012 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5934) );
  AOI22_X1 U7013 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6034), .B1(n5935), .B2(n5934), .ZN(n5936) );
  OAI211_X1 U7014 ( .C1(n6005), .C2(n4086), .A(n5936), .B(n5994), .ZN(n5937)
         );
  AOI21_X1 U7015 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5938), .A(n5937), .ZN(n5941) );
  AOI22_X1 U7016 ( .A1(n6056), .A2(n6026), .B1(n6041), .B2(n5939), .ZN(n5940)
         );
  OAI211_X1 U7017 ( .C1(n5942), .C2(n6029), .A(n5941), .B(n5940), .ZN(U2809)
         );
  INV_X1 U7018 ( .A(n5943), .ZN(n5944) );
  NOR3_X1 U7019 ( .A1(n5944), .A2(REIP_REG_16__SCAN_IN), .A3(n6528), .ZN(n5948) );
  OAI21_X1 U7020 ( .B1(n5945), .B2(n5954), .A(REIP_REG_16__SCAN_IN), .ZN(n5946) );
  OAI211_X1 U7021 ( .C1(n6005), .C2(n5601), .A(n5994), .B(n5946), .ZN(n5947)
         );
  AOI211_X1 U7022 ( .C1(n6034), .C2(EBX_REG_16__SCAN_IN), .A(n5948), .B(n5947), 
        .ZN(n5952) );
  INV_X1 U7023 ( .A(n5949), .ZN(n6064) );
  AOI22_X1 U7024 ( .A1(n6064), .A2(n6026), .B1(n6032), .B2(n5950), .ZN(n5951)
         );
  OAI211_X1 U7025 ( .C1(n6024), .C2(n5953), .A(n5952), .B(n5951), .ZN(U2811)
         );
  AOI22_X1 U7026 ( .A1(n6041), .A2(n5955), .B1(REIP_REG_14__SCAN_IN), .B2(
        n5954), .ZN(n5964) );
  AOI22_X1 U7027 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6031), .B1(n5957), 
        .B2(n5956), .ZN(n5963) );
  AOI21_X1 U7028 ( .B1(n6034), .B2(EBX_REG_14__SCAN_IN), .A(n6021), .ZN(n5962)
         );
  INV_X1 U7029 ( .A(n5958), .ZN(n5960) );
  AOI22_X1 U7030 ( .A1(n5960), .A2(n6026), .B1(n6032), .B2(n5959), .ZN(n5961)
         );
  NAND4_X1 U7031 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(U2813)
         );
  INV_X1 U7032 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5967) );
  INV_X1 U7033 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5966) );
  AOI21_X1 U7034 ( .B1(n5967), .B2(n5966), .A(n5965), .ZN(n5969) );
  AOI22_X1 U7035 ( .A1(n6041), .A2(n5970), .B1(n5969), .B2(n5968), .ZN(n5974)
         );
  AOI22_X1 U7036 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6031), .B1(
        REIP_REG_13__SCAN_IN), .B2(n5985), .ZN(n5971) );
  OAI211_X1 U7037 ( .C1(n6016), .C2(n6050), .A(n5971), .B(n5994), .ZN(n5972)
         );
  AOI21_X1 U7038 ( .B1(n6048), .B2(n6026), .A(n5972), .ZN(n5973) );
  OAI211_X1 U7039 ( .C1(n5975), .C2(n6029), .A(n5974), .B(n5973), .ZN(U2814)
         );
  INV_X1 U7040 ( .A(n5976), .ZN(n5979) );
  AOI21_X1 U7041 ( .B1(n5979), .B2(n5978), .A(n5977), .ZN(n5982) );
  INV_X1 U7042 ( .A(n5980), .ZN(n5981) );
  NOR2_X1 U7043 ( .A1(n5982), .A2(n5981), .ZN(n6140) );
  OAI22_X1 U7044 ( .A1(n6054), .A2(n6016), .B1(n5983), .B2(n6005), .ZN(n5984)
         );
  AOI211_X1 U7045 ( .C1(n6041), .C2(n6140), .A(n6021), .B(n5984), .ZN(n5991)
         );
  AOI22_X1 U7046 ( .A1(n6110), .A2(n6026), .B1(n6032), .B2(n6108), .ZN(n5990)
         );
  NAND2_X1 U7047 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5985), .ZN(n5989) );
  INV_X1 U7048 ( .A(n5986), .ZN(n5987) );
  NOR2_X1 U7049 ( .A1(n5987), .A2(n6517), .ZN(n6004) );
  INV_X1 U7050 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6524) );
  NAND4_X1 U7051 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n6004), .A4(n6524), .ZN(n5988) );
  NAND4_X1 U7052 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(U2816)
         );
  NAND2_X1 U7053 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6004), .ZN(n6003) );
  INV_X1 U7054 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6522) );
  INV_X1 U7055 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6519) );
  OAI21_X1 U7056 ( .B1(n6519), .B2(n5993), .A(n5992), .ZN(n6014) );
  NAND2_X1 U7057 ( .A1(n6034), .A2(EBX_REG_10__SCAN_IN), .ZN(n5995) );
  OAI211_X1 U7058 ( .C1(n6005), .C2(n5996), .A(n5995), .B(n5994), .ZN(n5997)
         );
  AOI21_X1 U7059 ( .B1(n6041), .B2(n6151), .A(n5997), .ZN(n5998) );
  OAI21_X1 U7060 ( .B1(n5999), .B2(n6009), .A(n5998), .ZN(n6000) );
  AOI21_X1 U7061 ( .B1(n6001), .B2(n6032), .A(n6000), .ZN(n6002) );
  OAI221_X1 U7062 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6003), .C1(n6522), .C2(
        n6014), .A(n6002), .ZN(U2817) );
  NOR2_X1 U7063 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6004), .ZN(n6015) );
  OAI22_X1 U7064 ( .A1(n6006), .A2(n6005), .B1(n6024), .B2(n6164), .ZN(n6007)
         );
  AOI211_X1 U7065 ( .C1(n6034), .C2(EBX_REG_9__SCAN_IN), .A(n6021), .B(n6007), 
        .ZN(n6013) );
  OAI22_X1 U7066 ( .A1(n6010), .A2(n6009), .B1(n6029), .B2(n6008), .ZN(n6011)
         );
  INV_X1 U7067 ( .A(n6011), .ZN(n6012) );
  OAI211_X1 U7068 ( .C1(n6015), .C2(n6014), .A(n6013), .B(n6012), .ZN(U2818)
         );
  NOR2_X1 U7069 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  AOI211_X1 U7070 ( .C1(n6020), .C2(REIP_REG_6__SCAN_IN), .A(n6019), .B(n6018), 
        .ZN(n6028) );
  AOI21_X1 U7071 ( .B1(n6031), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6021), 
        .ZN(n6022) );
  OAI21_X1 U7072 ( .B1(n6024), .B2(n6023), .A(n6022), .ZN(n6025) );
  AOI21_X1 U7073 ( .B1(n6114), .B2(n6026), .A(n6025), .ZN(n6027) );
  OAI211_X1 U7074 ( .C1(n6118), .C2(n6029), .A(n6028), .B(n6027), .ZN(U2821)
         );
  INV_X1 U7075 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7076 ( .A1(n6030), .A2(REIP_REG_2__SCAN_IN), .ZN(n6043) );
  INV_X1 U7077 ( .A(n6128), .ZN(n6033) );
  AOI22_X1 U7078 ( .A1(n6033), .A2(n6032), .B1(n6031), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7079 ( .A1(n6034), .A2(EBX_REG_3__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7080 ( .C1(n6322), .C2(n6037), .A(n6036), .B(n6035), .ZN(n6040)
         );
  NOR2_X1 U7081 ( .A1(n6123), .A2(n6038), .ZN(n6039) );
  AOI211_X1 U7082 ( .C1(n6041), .C2(n6200), .A(n6040), .B(n6039), .ZN(n6042)
         );
  OAI221_X1 U7083 ( .B1(n6044), .B2(n6509), .C1(n6044), .C2(n6043), .A(n6042), 
        .ZN(U2824) );
  NOR2_X1 U7084 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  AOI21_X1 U7085 ( .B1(n6048), .B2(n6052), .A(n6047), .ZN(n6049) );
  OAI21_X1 U7086 ( .B1(n6055), .B2(n6050), .A(n6049), .ZN(U2846) );
  AOI22_X1 U7087 ( .A1(n6110), .A2(n6052), .B1(n6051), .B2(n6140), .ZN(n6053)
         );
  OAI21_X1 U7088 ( .B1(n6055), .B2(n6054), .A(n6053), .ZN(U2848) );
  AOI22_X1 U7089 ( .A1(n6056), .A2(n6063), .B1(n6062), .B2(DATAI_18_), .ZN(
        n6058) );
  AOI22_X1 U7090 ( .A1(n6066), .A2(DATAI_2_), .B1(n6065), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7091 ( .A1(n6058), .A2(n6057), .ZN(U2873) );
  AOI22_X1 U7092 ( .A1(n6059), .A2(n6063), .B1(n6062), .B2(DATAI_17_), .ZN(
        n6061) );
  AOI22_X1 U7093 ( .A1(n6066), .A2(DATAI_1_), .B1(n6065), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7094 ( .A1(n6061), .A2(n6060), .ZN(U2874) );
  AOI22_X1 U7095 ( .A1(n6064), .A2(n6063), .B1(n6062), .B2(DATAI_16_), .ZN(
        n6068) );
  AOI22_X1 U7096 ( .A1(n6066), .A2(DATAI_0_), .B1(n6065), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7097 ( .A1(n6068), .A2(n6067), .ZN(U2875) );
  AOI22_X1 U7098 ( .A1(n6571), .A2(LWORD_REG_15__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U7099 ( .B1(n6071), .B2(n6102), .A(n6070), .ZN(U2908) );
  AOI22_X1 U7100 ( .A1(n6571), .A2(LWORD_REG_14__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U7101 ( .B1(n6073), .B2(n6102), .A(n6072), .ZN(U2909) );
  AOI22_X1 U7102 ( .A1(n6571), .A2(LWORD_REG_13__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U7103 ( .B1(n6075), .B2(n6102), .A(n6074), .ZN(U2910) );
  AOI22_X1 U7104 ( .A1(n6571), .A2(LWORD_REG_12__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U7105 ( .B1(n6077), .B2(n6102), .A(n6076), .ZN(U2911) );
  AOI22_X1 U7106 ( .A1(n6571), .A2(LWORD_REG_11__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7107 ( .B1(n6079), .B2(n6102), .A(n6078), .ZN(U2912) );
  AOI22_X1 U7108 ( .A1(n6571), .A2(LWORD_REG_10__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7109 ( .B1(n6081), .B2(n6102), .A(n6080), .ZN(U2913) );
  AOI22_X1 U7110 ( .A1(n6571), .A2(LWORD_REG_9__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7111 ( .B1(n6083), .B2(n6102), .A(n6082), .ZN(U2914) );
  AOI22_X1 U7112 ( .A1(n6571), .A2(LWORD_REG_8__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7113 ( .B1(n6085), .B2(n6102), .A(n6084), .ZN(U2915) );
  AOI22_X1 U7114 ( .A1(n6100), .A2(LWORD_REG_7__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7115 ( .B1(n6087), .B2(n6102), .A(n6086), .ZN(U2916) );
  AOI22_X1 U7116 ( .A1(n6100), .A2(LWORD_REG_6__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7117 ( .B1(n4669), .B2(n6102), .A(n6088), .ZN(U2917) );
  AOI22_X1 U7118 ( .A1(n6100), .A2(LWORD_REG_5__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7119 ( .B1(n3898), .B2(n6102), .A(n6089), .ZN(U2918) );
  AOI22_X1 U7120 ( .A1(n6100), .A2(LWORD_REG_4__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7121 ( .B1(n6092), .B2(n6102), .A(n6091), .ZN(U2919) );
  AOI22_X1 U7122 ( .A1(n6100), .A2(LWORD_REG_3__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7123 ( .B1(n6094), .B2(n6102), .A(n6093), .ZN(U2920) );
  AOI22_X1 U7124 ( .A1(n6100), .A2(LWORD_REG_2__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7125 ( .B1(n6096), .B2(n6102), .A(n6095), .ZN(U2921) );
  AOI22_X1 U7126 ( .A1(n6100), .A2(LWORD_REG_1__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7127 ( .B1(n6098), .B2(n6102), .A(n6097), .ZN(U2922) );
  AOI22_X1 U7128 ( .A1(n6100), .A2(LWORD_REG_0__SCAN_IN), .B1(n6099), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7129 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(U2923) );
  NAND2_X1 U7130 ( .A1(n6105), .A2(n6104), .ZN(n6107) );
  XNOR2_X1 U7131 ( .A(n3512), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6106)
         );
  XNOR2_X1 U7132 ( .A(n6107), .B(n6106), .ZN(n6145) );
  AOI22_X1 U7133 ( .A1(n6199), .A2(REIP_REG_11__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6112) );
  AOI22_X1 U7134 ( .A1(n6110), .A2(n6133), .B1(n6109), .B2(n6108), .ZN(n6111)
         );
  OAI211_X1 U7135 ( .C1(n6145), .C2(n6124), .A(n6112), .B(n6111), .ZN(U2975)
         );
  AOI22_X1 U7136 ( .A1(n6199), .A2(REIP_REG_6__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6117) );
  INV_X1 U7137 ( .A(n6113), .ZN(n6115) );
  AOI22_X1 U7138 ( .A1(n6115), .A2(n6135), .B1(n6114), .B2(n6133), .ZN(n6116)
         );
  OAI211_X1 U7139 ( .C1(n6139), .C2(n6118), .A(n6117), .B(n6116), .ZN(U2980)
         );
  AOI22_X1 U7140 ( .A1(n6199), .A2(REIP_REG_3__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7141 ( .B1(n6119), .B2(n6121), .A(n6120), .ZN(n6202) );
  OAI22_X1 U7142 ( .A1(n6202), .A2(n6124), .B1(n6123), .B2(n6122), .ZN(n6125)
         );
  INV_X1 U7143 ( .A(n6125), .ZN(n6126) );
  OAI211_X1 U7144 ( .C1(n6139), .C2(n6128), .A(n6127), .B(n6126), .ZN(U2983)
         );
  AOI22_X1 U7145 ( .A1(n6199), .A2(REIP_REG_2__SCAN_IN), .B1(n6129), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6137) );
  XOR2_X1 U7146 ( .A(n6130), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6132) );
  XNOR2_X1 U7147 ( .A(n6132), .B(n6131), .ZN(n6216) );
  AOI22_X1 U7148 ( .A1(n6135), .A2(n6216), .B1(n6134), .B2(n6133), .ZN(n6136)
         );
  OAI211_X1 U7149 ( .C1(n6139), .C2(n6138), .A(n6137), .B(n6136), .ZN(U2984)
         );
  AOI22_X1 U7150 ( .A1(n6140), .A2(n6223), .B1(n6199), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6144) );
  AOI22_X1 U7151 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6142), .B1(n6141), .B2(n3515), .ZN(n6143) );
  OAI211_X1 U7152 ( .C1(n6145), .C2(n6201), .A(n6144), .B(n6143), .ZN(U3007)
         );
  INV_X1 U7153 ( .A(n6203), .ZN(n6146) );
  NAND2_X1 U7154 ( .A1(n6158), .A2(n6182), .ZN(n6170) );
  AOI22_X1 U7155 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3514), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6148), .ZN(n6162) );
  INV_X1 U7156 ( .A(n6149), .ZN(n6150) );
  AOI21_X1 U7157 ( .B1(n6151), .B2(n6223), .A(n6150), .ZN(n6161) );
  AND2_X1 U7158 ( .A1(n6214), .A2(n6152), .ZN(n6154) );
  AOI211_X1 U7159 ( .C1(n6156), .C2(n6155), .A(n6154), .B(n6153), .ZN(n6187)
         );
  OAI21_X1 U7160 ( .B1(n6158), .B2(n6157), .A(n6187), .ZN(n6166) );
  AOI22_X1 U7161 ( .A1(n6159), .A2(n6229), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6166), .ZN(n6160) );
  OAI211_X1 U7162 ( .C1(n6170), .C2(n6162), .A(n6161), .B(n6160), .ZN(U3008)
         );
  OAI21_X1 U7163 ( .B1(n6164), .B2(n6193), .A(n6163), .ZN(n6165) );
  INV_X1 U7164 ( .A(n6165), .ZN(n6169) );
  AOI22_X1 U7165 ( .A1(n6167), .A2(n6229), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6166), .ZN(n6168) );
  OAI211_X1 U7166 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6170), .A(n6169), 
        .B(n6168), .ZN(U3009) );
  OAI222_X1 U7167 ( .A1(n6172), .A2(n6193), .B1(n6191), .B2(n6517), .C1(n6201), 
        .C2(n6171), .ZN(n6173) );
  INV_X1 U7168 ( .A(n6173), .ZN(n6176) );
  OAI211_X1 U7169 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6182), .B(n6174), .ZN(n6175) );
  OAI211_X1 U7170 ( .C1(n6187), .C2(n6177), .A(n6176), .B(n6175), .ZN(U3010)
         );
  INV_X1 U7171 ( .A(n6178), .ZN(n6179) );
  AOI21_X1 U7172 ( .B1(n6180), .B2(n6223), .A(n6179), .ZN(n6185) );
  INV_X1 U7173 ( .A(n6181), .ZN(n6183) );
  AOI22_X1 U7174 ( .A1(n6183), .A2(n6229), .B1(n6182), .B2(n6186), .ZN(n6184)
         );
  OAI211_X1 U7175 ( .C1(n6187), .C2(n6186), .A(n6185), .B(n6184), .ZN(U3011)
         );
  INV_X1 U7176 ( .A(n6209), .ZN(n6188) );
  AOI21_X1 U7177 ( .B1(n6214), .B2(n6188), .A(n6217), .ZN(n6208) );
  AOI211_X1 U7178 ( .C1(n6207), .C2(n6198), .A(n6189), .B(n6203), .ZN(n6196)
         );
  NOR2_X1 U7179 ( .A1(n6190), .A2(n6201), .ZN(n6195) );
  OAI22_X1 U7180 ( .A1(n6193), .A2(n6192), .B1(n6511), .B2(n6191), .ZN(n6194)
         );
  NOR3_X1 U7181 ( .A1(n6196), .A2(n6195), .A3(n6194), .ZN(n6197) );
  OAI21_X1 U7182 ( .B1(n6208), .B2(n6198), .A(n6197), .ZN(U3014) );
  AOI22_X1 U7183 ( .A1(n6223), .A2(n6200), .B1(n6199), .B2(REIP_REG_3__SCAN_IN), .ZN(n6206) );
  OAI22_X1 U7184 ( .A1(n6203), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6202), 
        .B2(n6201), .ZN(n6204) );
  INV_X1 U7185 ( .A(n6204), .ZN(n6205) );
  OAI211_X1 U7186 ( .C1(n6208), .C2(n6207), .A(n6206), .B(n6205), .ZN(U3015)
         );
  OAI21_X1 U7187 ( .B1(n6211), .B2(n6210), .A(n6209), .ZN(n6215) );
  AOI222_X1 U7188 ( .A1(n6215), .A2(n6214), .B1(REIP_REG_2__SCAN_IN), .B2(
        n6213), .C1(n6212), .C2(n6223), .ZN(n6219) );
  AOI22_X1 U7189 ( .A1(n6217), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6216), 
        .B2(n6229), .ZN(n6218) );
  OAI211_X1 U7190 ( .C1(INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n6220), .A(n6219), 
        .B(n6218), .ZN(U3016) );
  NAND2_X1 U7191 ( .A1(n6234), .A2(n6221), .ZN(n6226) );
  NAND2_X1 U7192 ( .A1(n6223), .A2(n6222), .ZN(n6225) );
  OAI211_X1 U7193 ( .C1(n6227), .C2(n6226), .A(n6225), .B(n6224), .ZN(n6228)
         );
  AOI21_X1 U7194 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(n6231) );
  OAI221_X1 U7195 ( .B1(n6234), .B2(n6233), .C1(n6234), .C2(n6232), .A(n6231), 
        .ZN(U3017) );
  AND2_X1 U7196 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6235), .ZN(U3019)
         );
  INV_X1 U7197 ( .A(n6361), .ZN(n6236) );
  NAND2_X1 U7198 ( .A1(n6236), .A2(n6446), .ZN(n6241) );
  INV_X1 U7199 ( .A(n6241), .ZN(n6269) );
  AOI22_X1 U7200 ( .A1(n6362), .A2(n6269), .B1(n6264), .B2(n6363), .ZN(n6249)
         );
  NAND2_X1 U7201 ( .A1(n6364), .A2(n6237), .ZN(n6238) );
  OAI21_X1 U7202 ( .B1(n6239), .B2(n6238), .A(n6365), .ZN(n6247) );
  OR2_X1 U7203 ( .A1(n6240), .A2(n3862), .ZN(n6242) );
  INV_X1 U7204 ( .A(n6246), .ZN(n6244) );
  AOI21_X1 U7205 ( .B1(n6371), .B2(n6245), .A(n6370), .ZN(n6243) );
  OAI21_X1 U7206 ( .B1(n6247), .B2(n6244), .A(n6243), .ZN(n6271) );
  OAI22_X1 U7207 ( .A1(n6247), .A2(n6246), .B1(n6245), .B2(n6374), .ZN(n6270)
         );
  AOI22_X1 U7208 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6271), .B1(n6378), 
        .B2(n6270), .ZN(n6248) );
  OAI211_X1 U7209 ( .C1(n6381), .C2(n6267), .A(n6249), .B(n6248), .ZN(U3044)
         );
  AOI22_X1 U7210 ( .A1(n6382), .A2(n6269), .B1(n6268), .B2(n6383), .ZN(n6251)
         );
  AOI22_X1 U7211 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6271), .B1(n6384), 
        .B2(n6270), .ZN(n6250) );
  OAI211_X1 U7212 ( .C1(n6387), .C2(n6274), .A(n6251), .B(n6250), .ZN(U3045)
         );
  AOI22_X1 U7213 ( .A1(n6388), .A2(n6269), .B1(n6268), .B2(n6298), .ZN(n6253)
         );
  AOI22_X1 U7214 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6271), .B1(n6390), 
        .B2(n6270), .ZN(n6252) );
  OAI211_X1 U7215 ( .C1(n6301), .C2(n6274), .A(n6253), .B(n6252), .ZN(U3046)
         );
  AOI22_X1 U7216 ( .A1(n6394), .A2(n6269), .B1(n6268), .B2(n6254), .ZN(n6256)
         );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6271), .B1(n6396), 
        .B2(n6270), .ZN(n6255) );
  OAI211_X1 U7218 ( .C1(n6257), .C2(n6274), .A(n6256), .B(n6255), .ZN(U3047)
         );
  AOI22_X1 U7219 ( .A1(n6400), .A2(n6269), .B1(n6268), .B2(n6401), .ZN(n6259)
         );
  AOI22_X1 U7220 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6271), .B1(n6402), 
        .B2(n6270), .ZN(n6258) );
  OAI211_X1 U7221 ( .C1(n6405), .C2(n6274), .A(n6259), .B(n6258), .ZN(U3048)
         );
  AOI22_X1 U7222 ( .A1(n6406), .A2(n6269), .B1(n6268), .B2(n6260), .ZN(n6262)
         );
  AOI22_X1 U7223 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6271), .B1(n6408), 
        .B2(n6270), .ZN(n6261) );
  OAI211_X1 U7224 ( .C1(n6263), .C2(n6274), .A(n6262), .B(n6261), .ZN(U3049)
         );
  AOI22_X1 U7225 ( .A1(n6412), .A2(n6269), .B1(n6264), .B2(n6350), .ZN(n6266)
         );
  AOI22_X1 U7226 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6271), .B1(n6415), 
        .B2(n6270), .ZN(n6265) );
  OAI211_X1 U7227 ( .C1(n6267), .C2(n6353), .A(n6266), .B(n6265), .ZN(U3050)
         );
  AOI22_X1 U7228 ( .A1(n6421), .A2(n6269), .B1(n6268), .B2(n6312), .ZN(n6273)
         );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6271), .B1(n6425), 
        .B2(n6270), .ZN(n6272) );
  OAI211_X1 U7230 ( .C1(n6319), .C2(n6274), .A(n6273), .B(n6272), .ZN(U3051)
         );
  AOI22_X1 U7231 ( .A1(n6362), .A2(n6276), .B1(n6378), .B2(n6275), .ZN(n6280)
         );
  AOI22_X1 U7232 ( .A1(n6278), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6284), 
        .B2(n6277), .ZN(n6279) );
  OAI211_X1 U7233 ( .C1(n6295), .C2(n6311), .A(n6280), .B(n6279), .ZN(U3068)
         );
  INV_X1 U7234 ( .A(n6283), .ZN(n6314) );
  AOI22_X1 U7235 ( .A1(n6362), .A2(n6314), .B1(n6313), .B2(n6284), .ZN(n6294)
         );
  INV_X1 U7236 ( .A(n6285), .ZN(n6286) );
  AOI21_X1 U7237 ( .B1(n6286), .B2(n6368), .A(n6314), .ZN(n6292) );
  INV_X1 U7238 ( .A(n6292), .ZN(n6289) );
  NAND2_X1 U7239 ( .A1(n6365), .A2(n6287), .ZN(n6291) );
  AOI21_X1 U7240 ( .B1(n6290), .B2(n6371), .A(n6370), .ZN(n6288) );
  OAI21_X1 U7241 ( .B1(n6289), .B2(n6291), .A(n6288), .ZN(n6316) );
  OAI22_X1 U7242 ( .A1(n6292), .A2(n6291), .B1(n6374), .B2(n6290), .ZN(n6315)
         );
  AOI22_X1 U7243 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6316), .B1(n6378), 
        .B2(n6315), .ZN(n6293) );
  OAI211_X1 U7244 ( .C1(n6295), .C2(n6360), .A(n6294), .B(n6293), .ZN(U3076)
         );
  INV_X1 U7245 ( .A(n6360), .ZN(n6308) );
  AOI22_X1 U7246 ( .A1(n6382), .A2(n6314), .B1(n6308), .B2(n6336), .ZN(n6297)
         );
  AOI22_X1 U7247 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6316), .B1(n6384), 
        .B2(n6315), .ZN(n6296) );
  OAI211_X1 U7248 ( .C1(n6339), .C2(n6311), .A(n6297), .B(n6296), .ZN(U3077)
         );
  AOI22_X1 U7249 ( .A1(n6388), .A2(n6314), .B1(n6313), .B2(n6298), .ZN(n6300)
         );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6316), .B1(n6390), 
        .B2(n6315), .ZN(n6299) );
  OAI211_X1 U7251 ( .C1(n6301), .C2(n6360), .A(n6300), .B(n6299), .ZN(U3078)
         );
  AOI22_X1 U7252 ( .A1(n6394), .A2(n6314), .B1(n6308), .B2(n6395), .ZN(n6303)
         );
  AOI22_X1 U7253 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6316), .B1(n6396), 
        .B2(n6315), .ZN(n6302) );
  OAI211_X1 U7254 ( .C1(n6399), .C2(n6311), .A(n6303), .B(n6302), .ZN(U3079)
         );
  AOI22_X1 U7255 ( .A1(n6400), .A2(n6314), .B1(n6308), .B2(n6344), .ZN(n6305)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6316), .B1(n6402), 
        .B2(n6315), .ZN(n6304) );
  OAI211_X1 U7257 ( .C1(n6347), .C2(n6311), .A(n6305), .B(n6304), .ZN(U3080)
         );
  AOI22_X1 U7258 ( .A1(n6406), .A2(n6314), .B1(n6308), .B2(n6407), .ZN(n6307)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6316), .B1(n6408), 
        .B2(n6315), .ZN(n6306) );
  OAI211_X1 U7260 ( .C1(n6411), .C2(n6311), .A(n6307), .B(n6306), .ZN(U3081)
         );
  AOI22_X1 U7261 ( .A1(n6412), .A2(n6314), .B1(n6308), .B2(n6350), .ZN(n6310)
         );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6316), .B1(n6415), 
        .B2(n6315), .ZN(n6309) );
  OAI211_X1 U7263 ( .C1(n6353), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3082)
         );
  AOI22_X1 U7264 ( .A1(n6421), .A2(n6314), .B1(n6313), .B2(n6312), .ZN(n6318)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6316), .B1(n6425), 
        .B2(n6315), .ZN(n6317) );
  OAI211_X1 U7266 ( .C1(n6319), .C2(n6360), .A(n6318), .B(n6317), .ZN(U3083)
         );
  NOR2_X1 U7267 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6320), .ZN(n6354)
         );
  NOR2_X1 U7268 ( .A1(n6322), .A2(n6321), .ZN(n6327) );
  INV_X1 U7269 ( .A(n6327), .ZN(n6325) );
  OAI22_X1 U7270 ( .A1(n6325), .A2(n6371), .B1(n6324), .B2(n6323), .ZN(n6355)
         );
  AOI22_X1 U7271 ( .A1(n6362), .A2(n6354), .B1(n6378), .B2(n6355), .ZN(n6335)
         );
  INV_X1 U7272 ( .A(n6356), .ZN(n6326) );
  NAND3_X1 U7273 ( .A1(n6326), .A2(n6365), .A3(n6360), .ZN(n6329) );
  AOI21_X1 U7274 ( .B1(n6329), .B2(n6328), .A(n6327), .ZN(n6333) );
  OAI211_X1 U7275 ( .C1(n6560), .C2(n6354), .A(n6331), .B(n6330), .ZN(n6332)
         );
  AOI22_X1 U7276 ( .A1(n6357), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6363), 
        .B2(n6356), .ZN(n6334) );
  OAI211_X1 U7277 ( .C1(n6381), .C2(n6360), .A(n6335), .B(n6334), .ZN(U3084)
         );
  AOI22_X1 U7278 ( .A1(n6382), .A2(n6354), .B1(n6384), .B2(n6355), .ZN(n6338)
         );
  AOI22_X1 U7279 ( .A1(n6357), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6336), 
        .B2(n6356), .ZN(n6337) );
  OAI211_X1 U7280 ( .C1(n6339), .C2(n6360), .A(n6338), .B(n6337), .ZN(U3085)
         );
  AOI22_X1 U7281 ( .A1(n6388), .A2(n6354), .B1(n6390), .B2(n6355), .ZN(n6341)
         );
  AOI22_X1 U7282 ( .A1(n6357), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6389), 
        .B2(n6356), .ZN(n6340) );
  OAI211_X1 U7283 ( .C1(n6393), .C2(n6360), .A(n6341), .B(n6340), .ZN(U3086)
         );
  AOI22_X1 U7284 ( .A1(n6394), .A2(n6354), .B1(n6396), .B2(n6355), .ZN(n6343)
         );
  AOI22_X1 U7285 ( .A1(n6357), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6395), 
        .B2(n6356), .ZN(n6342) );
  OAI211_X1 U7286 ( .C1(n6399), .C2(n6360), .A(n6343), .B(n6342), .ZN(U3087)
         );
  AOI22_X1 U7287 ( .A1(n6400), .A2(n6354), .B1(n6402), .B2(n6355), .ZN(n6346)
         );
  AOI22_X1 U7288 ( .A1(n6357), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6344), 
        .B2(n6356), .ZN(n6345) );
  OAI211_X1 U7289 ( .C1(n6347), .C2(n6360), .A(n6346), .B(n6345), .ZN(U3088)
         );
  AOI22_X1 U7290 ( .A1(n6406), .A2(n6354), .B1(n6408), .B2(n6355), .ZN(n6349)
         );
  AOI22_X1 U7291 ( .A1(n6357), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6407), 
        .B2(n6356), .ZN(n6348) );
  OAI211_X1 U7292 ( .C1(n6411), .C2(n6360), .A(n6349), .B(n6348), .ZN(U3089)
         );
  AOI22_X1 U7293 ( .A1(n6412), .A2(n6354), .B1(n6415), .B2(n6355), .ZN(n6352)
         );
  AOI22_X1 U7294 ( .A1(n6357), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6350), 
        .B2(n6356), .ZN(n6351) );
  OAI211_X1 U7295 ( .C1(n6353), .C2(n6360), .A(n6352), .B(n6351), .ZN(U3090)
         );
  AOI22_X1 U7296 ( .A1(n6425), .A2(n6355), .B1(n6421), .B2(n6354), .ZN(n6359)
         );
  AOI22_X1 U7297 ( .A1(n6357), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6423), 
        .B2(n6356), .ZN(n6358) );
  OAI211_X1 U7298 ( .C1(n6430), .C2(n6360), .A(n6359), .B(n6358), .ZN(U3091)
         );
  INV_X1 U7299 ( .A(n6418), .ZN(n6422) );
  NOR2_X1 U7300 ( .A1(n6361), .A2(n6446), .ZN(n6420) );
  AOI22_X1 U7301 ( .A1(n6363), .A2(n6422), .B1(n6362), .B2(n6420), .ZN(n6380)
         );
  INV_X1 U7302 ( .A(n6364), .ZN(n6367) );
  OAI21_X1 U7303 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6377) );
  AOI21_X1 U7304 ( .B1(n6369), .B2(n6368), .A(n6420), .ZN(n6376) );
  INV_X1 U7305 ( .A(n6376), .ZN(n6373) );
  AOI21_X1 U7306 ( .B1(n6371), .B2(n6375), .A(n6370), .ZN(n6372) );
  OAI21_X1 U7307 ( .B1(n6377), .B2(n6373), .A(n6372), .ZN(n6426) );
  OAI22_X1 U7308 ( .A1(n6377), .A2(n6376), .B1(n6375), .B2(n6374), .ZN(n6424)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6426), .B1(n6378), 
        .B2(n6424), .ZN(n6379) );
  OAI211_X1 U7310 ( .C1(n6381), .C2(n6429), .A(n6380), .B(n6379), .ZN(U3108)
         );
  INV_X1 U7311 ( .A(n6429), .ZN(n6414) );
  AOI22_X1 U7312 ( .A1(n6414), .A2(n6383), .B1(n6382), .B2(n6420), .ZN(n6386)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6426), .B1(n6384), 
        .B2(n6424), .ZN(n6385) );
  OAI211_X1 U7314 ( .C1(n6387), .C2(n6418), .A(n6386), .B(n6385), .ZN(U3109)
         );
  AOI22_X1 U7315 ( .A1(n6389), .A2(n6422), .B1(n6388), .B2(n6420), .ZN(n6392)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6426), .B1(n6390), 
        .B2(n6424), .ZN(n6391) );
  OAI211_X1 U7317 ( .C1(n6393), .C2(n6429), .A(n6392), .B(n6391), .ZN(U3110)
         );
  AOI22_X1 U7318 ( .A1(n6395), .A2(n6422), .B1(n6394), .B2(n6420), .ZN(n6398)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6426), .B1(n6396), 
        .B2(n6424), .ZN(n6397) );
  OAI211_X1 U7320 ( .C1(n6399), .C2(n6429), .A(n6398), .B(n6397), .ZN(U3111)
         );
  AOI22_X1 U7321 ( .A1(n6414), .A2(n6401), .B1(n6400), .B2(n6420), .ZN(n6404)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6426), .B1(n6402), 
        .B2(n6424), .ZN(n6403) );
  OAI211_X1 U7323 ( .C1(n6405), .C2(n6418), .A(n6404), .B(n6403), .ZN(U3112)
         );
  AOI22_X1 U7324 ( .A1(n6407), .A2(n6422), .B1(n6406), .B2(n6420), .ZN(n6410)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6426), .B1(n6408), 
        .B2(n6424), .ZN(n6409) );
  OAI211_X1 U7326 ( .C1(n6411), .C2(n6429), .A(n6410), .B(n6409), .ZN(U3113)
         );
  AOI22_X1 U7327 ( .A1(n6414), .A2(n6413), .B1(n6412), .B2(n6420), .ZN(n6417)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6426), .B1(n6415), 
        .B2(n6424), .ZN(n6416) );
  OAI211_X1 U7329 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n6416), .ZN(U3114)
         );
  AOI22_X1 U7330 ( .A1(n6423), .A2(n6422), .B1(n6421), .B2(n6420), .ZN(n6428)
         );
  AOI22_X1 U7331 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6426), .B1(n6425), 
        .B2(n6424), .ZN(n6427) );
  OAI211_X1 U7332 ( .C1(n6430), .C2(n6429), .A(n6428), .B(n6427), .ZN(U3115)
         );
  INV_X1 U7333 ( .A(n6431), .ZN(n6432) );
  OAI211_X1 U7334 ( .C1(n3047), .C2(n6433), .A(n6432), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6438) );
  AOI22_X1 U7335 ( .A1(n6438), .A2(n6437), .B1(n6434), .B2(n6439), .ZN(n6435)
         );
  INV_X1 U7336 ( .A(n6435), .ZN(n6436) );
  OAI21_X1 U7337 ( .B1(n6438), .B2(n6437), .A(n6436), .ZN(n6442) );
  MUX2_X1 U7338 ( .A(n2996), .B(n6440), .S(n6439), .Z(n6452) );
  AOI222_X1 U7339 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6442), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6452), .C1(n6442), .C2(n6452), 
        .ZN(n6447) );
  MUX2_X1 U7340 ( .A(n6445), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6443), 
        .Z(n6450) );
  OAI21_X1 U7341 ( .B1(n6447), .B2(n6446), .A(n6450), .ZN(n6449) );
  NAND2_X1 U7342 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  AOI21_X1 U7343 ( .B1(n6449), .B2(n6448), .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .ZN(n6460) );
  INV_X1 U7344 ( .A(n6450), .ZN(n6451) );
  NOR2_X1 U7345 ( .A1(n6452), .A2(n6451), .ZN(n6459) );
  OAI21_X1 U7346 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6453), 
        .ZN(n6456) );
  NAND3_X1 U7347 ( .A1(n6456), .A2(n6455), .A3(n6454), .ZN(n6457) );
  NOR4_X1 U7348 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6474)
         );
  OR3_X1 U7349 ( .A1(n6462), .A2(n6573), .A3(n6461), .ZN(n6463) );
  NAND2_X1 U7350 ( .A1(n6463), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6464) );
  AOI221_X1 U7351 ( .B1(n6465), .B2(n6466), .C1(n4287), .C2(n6466), .A(n6464), 
        .ZN(n6469) );
  OAI221_X1 U7352 ( .B1(n6466), .B2(n6474), .C1(n6466), .C2(n6465), .A(n6469), 
        .ZN(n6559) );
  OAI21_X1 U7353 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4287), .A(n6559), .ZN(
        n6475) );
  AOI221_X1 U7354 ( .B1(n6468), .B2(STATE2_REG_0__SCAN_IN), .C1(n6475), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6467), .ZN(n6473) );
  AOI211_X1 U7355 ( .C1(n6574), .C2(n6470), .A(STATE2_REG_0__SCAN_IN), .B(
        n6469), .ZN(n6471) );
  INV_X1 U7356 ( .A(n6471), .ZN(n6472) );
  OAI211_X1 U7357 ( .C1(n6474), .C2(n6477), .A(n6473), .B(n6472), .ZN(U3148)
         );
  NAND3_X1 U7358 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6476), .A3(n6475), .ZN(
        n6482) );
  OAI21_X1 U7359 ( .B1(READY_N), .B2(n6478), .A(n6477), .ZN(n6480) );
  AOI21_X1 U7360 ( .B1(n6480), .B2(n6559), .A(n6479), .ZN(n6481) );
  NAND2_X1 U7361 ( .A1(n6482), .A2(n6481), .ZN(U3149) );
  OAI211_X1 U7362 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4287), .A(n6557), .B(
        n6483), .ZN(n6485) );
  OAI21_X1 U7363 ( .B1(n6486), .B2(n6485), .A(n6484), .ZN(U3150) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6487), .ZN(U3151) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6487), .ZN(U3152) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6487), .ZN(U3153) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6487), .ZN(U3154) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6487), .ZN(U3155) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6487), .ZN(U3156) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6487), .ZN(U3157) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6487), .ZN(U3158) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6487), .ZN(U3159) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6487), .ZN(U3160) );
  AND2_X1 U7374 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6487), .ZN(U3161) );
  AND2_X1 U7375 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6487), .ZN(U3162) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6487), .ZN(U3163) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6487), .ZN(U3164) );
  AND2_X1 U7378 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6487), .ZN(U3165) );
  AND2_X1 U7379 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6487), .ZN(U3166) );
  AND2_X1 U7380 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6487), .ZN(U3167) );
  AND2_X1 U7381 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6487), .ZN(U3168) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6487), .ZN(U3169) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6487), .ZN(U3170) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6487), .ZN(U3171) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6487), .ZN(U3172) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6487), .ZN(U3173) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6487), .ZN(U3174) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6487), .ZN(U3175) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6487), .ZN(U3176) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6487), .ZN(U3177) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6487), .ZN(U3178) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6487), .ZN(U3179) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6487), .ZN(U3180) );
  INV_X1 U7394 ( .A(HOLD), .ZN(n6702) );
  NOR2_X1 U7395 ( .A1(n6488), .A2(n6702), .ZN(n6494) );
  INV_X1 U7396 ( .A(n6494), .ZN(n6492) );
  NAND2_X1 U7397 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6493) );
  NAND2_X1 U7398 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U7399 ( .A1(n6493), .A2(n6500), .ZN(n6489) );
  INV_X1 U7400 ( .A(NA_N), .ZN(n6610) );
  AOI221_X1 U7401 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6610), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6505) );
  AOI21_X1 U7402 ( .B1(n6490), .B2(n6489), .A(n6505), .ZN(n6491) );
  OAI221_X1 U7403 ( .B1(n6581), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6581), 
        .C2(n6492), .A(n6491), .ZN(U3181) );
  INV_X1 U7404 ( .A(n6493), .ZN(n6497) );
  AOI21_X1 U7405 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6494), .ZN(n6496) );
  OAI211_X1 U7406 ( .C1(n6497), .C2(n6496), .A(n6495), .B(n6500), .ZN(U3182)
         );
  AOI221_X1 U7407 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4287), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6499) );
  AOI221_X1 U7408 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6499), .C2(HOLD), .A(n6498), .ZN(n6504) );
  INV_X1 U7409 ( .A(n6500), .ZN(n6501) );
  NAND4_X1 U7410 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6501), .A4(n6610), .ZN(n6503) );
  NAND3_X1 U7411 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6502) );
  OAI211_X1 U7412 ( .C1(n6505), .C2(n6504), .A(n6503), .B(n6502), .ZN(U3183)
         );
  NAND2_X1 U7413 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6581), .ZN(n6552) );
  INV_X2 U7414 ( .A(n6581), .ZN(n6580) );
  NOR2_X2 U7415 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6580), .ZN(n6550) );
  AOI22_X1 U7416 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6580), .ZN(n6506) );
  OAI21_X1 U7417 ( .B1(n6561), .B2(n6552), .A(n6506), .ZN(U3184) );
  AOI22_X1 U7418 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6580), .ZN(n6507) );
  OAI21_X1 U7419 ( .B1(n4938), .B2(n6552), .A(n6507), .ZN(U3185) );
  AOI22_X1 U7420 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6580), .ZN(n6508) );
  OAI21_X1 U7421 ( .B1(n6509), .B2(n6552), .A(n6508), .ZN(U3186) );
  AOI22_X1 U7422 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6580), .ZN(n6510) );
  OAI21_X1 U7423 ( .B1(n6511), .B2(n6552), .A(n6510), .ZN(U3187) );
  AOI22_X1 U7424 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6580), .ZN(n6512) );
  OAI21_X1 U7425 ( .B1(n6513), .B2(n6552), .A(n6512), .ZN(U3188) );
  AOI22_X1 U7426 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6580), .ZN(n6514) );
  OAI21_X1 U7427 ( .B1(n6515), .B2(n6552), .A(n6514), .ZN(U3189) );
  INV_X1 U7428 ( .A(n6552), .ZN(n6545) );
  AOI22_X1 U7429 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6580), .ZN(n6516) );
  OAI21_X1 U7430 ( .B1(n6517), .B2(n6547), .A(n6516), .ZN(U3190) );
  AOI22_X1 U7431 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6580), .ZN(n6518) );
  OAI21_X1 U7432 ( .B1(n6519), .B2(n6547), .A(n6518), .ZN(U3191) );
  AOI22_X1 U7433 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6580), .ZN(n6520) );
  OAI21_X1 U7434 ( .B1(n6522), .B2(n6547), .A(n6520), .ZN(U3192) );
  AOI22_X1 U7435 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6580), .ZN(n6521) );
  OAI21_X1 U7436 ( .B1(n6522), .B2(n6552), .A(n6521), .ZN(U3193) );
  AOI22_X1 U7437 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6580), .ZN(n6523) );
  OAI21_X1 U7438 ( .B1(n6524), .B2(n6552), .A(n6523), .ZN(U3194) );
  AOI22_X1 U7439 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6580), .ZN(n6525) );
  OAI21_X1 U7440 ( .B1(n5966), .B2(n6547), .A(n6525), .ZN(U3195) );
  AOI22_X1 U7441 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6580), .ZN(n6526) );
  OAI21_X1 U7442 ( .B1(n5966), .B2(n6552), .A(n6526), .ZN(U3196) );
  AOI22_X1 U7443 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6580), .ZN(n6527) );
  OAI21_X1 U7444 ( .B1(n6528), .B2(n6547), .A(n6527), .ZN(U3197) );
  AOI22_X1 U7445 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6580), .ZN(n6529) );
  OAI21_X1 U7446 ( .B1(n6531), .B2(n6547), .A(n6529), .ZN(U3198) );
  AOI22_X1 U7447 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6580), .ZN(n6530) );
  OAI21_X1 U7448 ( .B1(n6531), .B2(n6552), .A(n6530), .ZN(U3199) );
  AOI22_X1 U7449 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6580), .ZN(n6532) );
  OAI21_X1 U7450 ( .B1(n6533), .B2(n6552), .A(n6532), .ZN(U3200) );
  INV_X1 U7451 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7452 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6580), .ZN(n6534) );
  OAI21_X1 U7453 ( .B1(n6736), .B2(n6547), .A(n6534), .ZN(U3201) );
  AOI22_X1 U7454 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6580), .ZN(n6535) );
  OAI21_X1 U7455 ( .B1(n6736), .B2(n6552), .A(n6535), .ZN(U3202) );
  AOI22_X1 U7456 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6580), .ZN(n6536) );
  OAI21_X1 U7457 ( .B1(n6703), .B2(n6552), .A(n6536), .ZN(U3203) );
  AOI22_X1 U7458 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6580), .ZN(n6537) );
  OAI21_X1 U7459 ( .B1(n6697), .B2(n6552), .A(n6537), .ZN(U3204) );
  AOI22_X1 U7460 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6580), .ZN(n6538) );
  OAI21_X1 U7461 ( .B1(n6540), .B2(n6547), .A(n6538), .ZN(U3205) );
  AOI22_X1 U7462 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6580), .ZN(n6539) );
  OAI21_X1 U7463 ( .B1(n6540), .B2(n6552), .A(n6539), .ZN(U3206) );
  AOI22_X1 U7464 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6580), .ZN(n6541) );
  OAI21_X1 U7465 ( .B1(n6745), .B2(n6547), .A(n6541), .ZN(U3207) );
  AOI22_X1 U7466 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6580), .ZN(n6542) );
  OAI21_X1 U7467 ( .B1(n6745), .B2(n6552), .A(n6542), .ZN(U3208) );
  AOI22_X1 U7468 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6580), .ZN(n6543) );
  OAI21_X1 U7469 ( .B1(n6706), .B2(n6547), .A(n6543), .ZN(U3209) );
  AOI22_X1 U7470 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6580), .ZN(n6544) );
  OAI21_X1 U7471 ( .B1(n6692), .B2(n6547), .A(n6544), .ZN(U3210) );
  AOI22_X1 U7472 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6545), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6580), .ZN(n6546) );
  OAI21_X1 U7473 ( .B1(n6549), .B2(n6547), .A(n6546), .ZN(U3211) );
  AOI22_X1 U7474 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6580), .ZN(n6548) );
  OAI21_X1 U7475 ( .B1(n6549), .B2(n6552), .A(n6548), .ZN(U3212) );
  AOI22_X1 U7476 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6580), .ZN(n6551) );
  OAI21_X1 U7477 ( .B1(n6587), .B2(n6552), .A(n6551), .ZN(U3213) );
  MUX2_X1 U7478 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6580), .Z(U3446) );
  MUX2_X1 U7479 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6580), .Z(U3447) );
  MUX2_X1 U7480 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6580), .Z(U3448) );
  OAI21_X1 U7481 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6556), .A(n6554), .ZN(
        n6553) );
  INV_X1 U7482 ( .A(n6553), .ZN(U3451) );
  OAI21_X1 U7483 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(U3452) );
  OAI211_X1 U7484 ( .C1(n6560), .C2(n6559), .A(n6558), .B(n6557), .ZN(U3453)
         );
  AOI21_X1 U7485 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U7486 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6562), .B2(n6561), .ZN(n6564) );
  INV_X1 U7487 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6691) );
  AOI22_X1 U7488 ( .A1(n6566), .A2(n6564), .B1(n6691), .B2(n6563), .ZN(U3468)
         );
  INV_X1 U7489 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6751) );
  OAI21_X1 U7490 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6566), .ZN(n6565) );
  OAI21_X1 U7491 ( .B1(n6566), .B2(n6751), .A(n6565), .ZN(U3469) );
  INV_X1 U7492 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6567) );
  OAI22_X1 U7493 ( .A1(n6580), .A2(n6567), .B1(W_R_N_REG_SCAN_IN), .B2(n6581), 
        .ZN(n6568) );
  INV_X1 U7494 ( .A(n6568), .ZN(U3470) );
  AOI211_X1 U7495 ( .C1(n6571), .C2(n4287), .A(n6570), .B(n6569), .ZN(n6578)
         );
  OAI211_X1 U7496 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6573), .A(n6572), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6575) );
  AOI21_X1 U7497 ( .B1(n6575), .B2(STATE2_REG_0__SCAN_IN), .A(n6574), .ZN(
        n6577) );
  NAND2_X1 U7498 ( .A1(n6578), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6576) );
  OAI21_X1 U7499 ( .B1(n6578), .B2(n6577), .A(n6576), .ZN(U3472) );
  INV_X1 U7500 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7501 ( .A1(n6581), .A2(n6579), .B1(n6601), .B2(n6580), .ZN(U3473)
         );
  AOI22_X1 U7502 ( .A1(n6581), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6580), .ZN(n6784) );
  AOI22_X1 U7503 ( .A1(n6719), .A2(keyinput_g27), .B1(n6692), .B2(keyinput_g54), .ZN(n6582) );
  OAI221_X1 U7504 ( .B1(n6719), .B2(keyinput_g27), .C1(n6692), .C2(
        keyinput_g54), .A(n6582), .ZN(n6591) );
  INV_X1 U7505 ( .A(DATAI_27_), .ZN(n6699) );
  AOI22_X1 U7506 ( .A1(n6699), .A2(keyinput_g4), .B1(n6758), .B2(keyinput_g43), 
        .ZN(n6583) );
  OAI221_X1 U7507 ( .B1(n6699), .B2(keyinput_g4), .C1(n6758), .C2(keyinput_g43), .A(n6583), .ZN(n6590) );
  INV_X1 U7508 ( .A(DATAI_30_), .ZN(n6585) );
  AOI22_X1 U7509 ( .A1(n6760), .A2(keyinput_g31), .B1(n6585), .B2(keyinput_g1), 
        .ZN(n6584) );
  OAI221_X1 U7510 ( .B1(n6760), .B2(keyinput_g31), .C1(n6585), .C2(keyinput_g1), .A(n6584), .ZN(n6589) );
  AOI22_X1 U7511 ( .A1(n6706), .A2(keyinput_g55), .B1(n6587), .B2(keyinput_g52), .ZN(n6586) );
  OAI221_X1 U7512 ( .B1(n6706), .B2(keyinput_g55), .C1(n6587), .C2(
        keyinput_g52), .A(n6586), .ZN(n6588) );
  NOR4_X1 U7513 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6631)
         );
  INV_X1 U7514 ( .A(BS16_N), .ZN(n6593) );
  AOI22_X1 U7515 ( .A1(n6594), .A2(keyinput_g45), .B1(keyinput_g34), .B2(n6593), .ZN(n6592) );
  OAI221_X1 U7516 ( .B1(n6594), .B2(keyinput_g45), .C1(n6593), .C2(
        keyinput_g34), .A(n6592), .ZN(n6605) );
  INV_X1 U7517 ( .A(DATAI_19_), .ZN(n6596) );
  AOI22_X1 U7518 ( .A1(n6596), .A2(keyinput_g12), .B1(keyinput_g47), .B2(n6751), .ZN(n6595) );
  OAI221_X1 U7519 ( .B1(n6596), .B2(keyinput_g12), .C1(n6751), .C2(
        keyinput_g47), .A(n6595), .ZN(n6604) );
  INV_X1 U7520 ( .A(DATAI_24_), .ZN(n6599) );
  INV_X1 U7521 ( .A(DATAI_26_), .ZN(n6598) );
  AOI22_X1 U7522 ( .A1(n6599), .A2(keyinput_g7), .B1(n6598), .B2(keyinput_g5), 
        .ZN(n6597) );
  OAI221_X1 U7523 ( .B1(n6599), .B2(keyinput_g7), .C1(n6598), .C2(keyinput_g5), 
        .A(n6597), .ZN(n6603) );
  INV_X1 U7524 ( .A(MORE_REG_SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7525 ( .A1(n6601), .A2(keyinput_g40), .B1(n6757), .B2(keyinput_g44), .ZN(n6600) );
  OAI221_X1 U7526 ( .B1(n6601), .B2(keyinput_g40), .C1(n6757), .C2(
        keyinput_g44), .A(n6600), .ZN(n6602) );
  NOR4_X1 U7527 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n6630)
         );
  INV_X1 U7528 ( .A(DATAI_11_), .ZN(n6607) );
  AOI22_X1 U7529 ( .A1(n6607), .A2(keyinput_g20), .B1(n6739), .B2(keyinput_g58), .ZN(n6606) );
  OAI221_X1 U7530 ( .B1(n6607), .B2(keyinput_g20), .C1(n6739), .C2(
        keyinput_g58), .A(n6606), .ZN(n6616) );
  AOI22_X1 U7531 ( .A1(n6610), .A2(keyinput_g33), .B1(n6609), .B2(keyinput_g38), .ZN(n6608) );
  OAI221_X1 U7532 ( .B1(n6610), .B2(keyinput_g33), .C1(n6609), .C2(
        keyinput_g38), .A(n6608), .ZN(n6615) );
  AOI22_X1 U7533 ( .A1(n6697), .A2(keyinput_g61), .B1(keyinput_g28), .B2(n6738), .ZN(n6611) );
  OAI221_X1 U7534 ( .B1(n6697), .B2(keyinput_g61), .C1(n6738), .C2(
        keyinput_g28), .A(n6611), .ZN(n6614) );
  AOI22_X1 U7535 ( .A1(n6745), .A2(keyinput_g57), .B1(keyinput_g50), .B2(n6718), .ZN(n6612) );
  OAI221_X1 U7536 ( .B1(n6745), .B2(keyinput_g57), .C1(n6718), .C2(
        keyinput_g50), .A(n6612), .ZN(n6613) );
  NOR4_X1 U7537 ( .A1(n6616), .A2(n6615), .A3(n6614), .A4(n6613), .ZN(n6629)
         );
  INV_X1 U7538 ( .A(DATAI_20_), .ZN(n6618) );
  AOI22_X1 U7539 ( .A1(n4287), .A2(keyinput_g35), .B1(keyinput_g11), .B2(n6618), .ZN(n6617) );
  OAI221_X1 U7540 ( .B1(n4287), .B2(keyinput_g35), .C1(n6618), .C2(
        keyinput_g11), .A(n6617), .ZN(n6627) );
  INV_X1 U7541 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7542 ( .A1(n6691), .A2(keyinput_g49), .B1(n6742), .B2(keyinput_g56), .ZN(n6619) );
  OAI221_X1 U7543 ( .B1(n6691), .B2(keyinput_g49), .C1(n6742), .C2(
        keyinput_g56), .A(n6619), .ZN(n6626) );
  INV_X1 U7544 ( .A(DATAI_17_), .ZN(n6721) );
  INV_X1 U7545 ( .A(DATAI_10_), .ZN(n6621) );
  AOI22_X1 U7546 ( .A1(n6721), .A2(keyinput_g14), .B1(n6621), .B2(keyinput_g21), .ZN(n6620) );
  OAI221_X1 U7547 ( .B1(n6721), .B2(keyinput_g14), .C1(n6621), .C2(
        keyinput_g21), .A(n6620), .ZN(n6625) );
  INV_X1 U7548 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6689) );
  INV_X1 U7549 ( .A(DATAI_8_), .ZN(n6623) );
  AOI22_X1 U7550 ( .A1(n6689), .A2(keyinput_g51), .B1(keyinput_g23), .B2(n6623), .ZN(n6622) );
  OAI221_X1 U7551 ( .B1(n6689), .B2(keyinput_g51), .C1(n6623), .C2(
        keyinput_g23), .A(n6622), .ZN(n6624) );
  NOR4_X1 U7552 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6628)
         );
  NAND4_X1 U7553 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6782)
         );
  AOI22_X1 U7554 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(REIP_REG_23__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n6632) );
  OAI221_X1 U7555 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6632), .ZN(n6639) );
  AOI22_X1 U7556 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        DATAI_21_), .B2(keyinput_g10), .ZN(n6633) );
  OAI221_X1 U7557 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        DATAI_21_), .C2(keyinput_g10), .A(n6633), .ZN(n6638) );
  AOI22_X1 U7558 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        DATAI_22_), .B2(keyinput_g9), .ZN(n6634) );
  OAI221_X1 U7559 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        DATAI_22_), .C2(keyinput_g9), .A(n6634), .ZN(n6637) );
  AOI22_X1 U7560 ( .A1(HOLD), .A2(keyinput_g36), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n6635) );
  OAI221_X1 U7561 ( .B1(HOLD), .B2(keyinput_g36), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n6635), .ZN(n6636) );
  NOR4_X1 U7562 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6666)
         );
  INV_X1 U7563 ( .A(DATAI_12_), .ZN(n6684) );
  XNOR2_X1 U7564 ( .A(n6684), .B(keyinput_g19), .ZN(n6646) );
  AOI22_X1 U7565 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_g63), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6640) );
  OAI221_X1 U7566 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6640), .ZN(n6645) );
  AOI22_X1 U7567 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n6641) );
  OAI221_X1 U7568 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n6641), .ZN(n6644) );
  AOI22_X1 U7569 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAI_25_), .B2(keyinput_g6), .ZN(n6642) );
  OAI221_X1 U7570 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        DATAI_25_), .C2(keyinput_g6), .A(n6642), .ZN(n6643) );
  NOR4_X1 U7571 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6665)
         );
  AOI22_X1 U7572 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6647) );
  OAI221_X1 U7573 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6647), .ZN(n6654) );
  AOI22_X1 U7574 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        DATAI_13_), .B2(keyinput_g18), .ZN(n6648) );
  OAI221_X1 U7575 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        DATAI_13_), .C2(keyinput_g18), .A(n6648), .ZN(n6653) );
  INV_X1 U7576 ( .A(DATAI_9_), .ZN(n6761) );
  AOI22_X1 U7577 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(n6761), .B2(
        keyinput_g22), .ZN(n6649) );
  OAI221_X1 U7578 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(n6761), .C2(
        keyinput_g22), .A(n6649), .ZN(n6652) );
  AOI22_X1 U7579 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(DATAI_6_), 
        .B2(keyinput_g25), .ZN(n6650) );
  OAI221_X1 U7580 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(DATAI_6_), 
        .C2(keyinput_g25), .A(n6650), .ZN(n6651) );
  NOR4_X1 U7581 ( .A1(n6654), .A2(n6653), .A3(n6652), .A4(n6651), .ZN(n6664)
         );
  AOI22_X1 U7582 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(DATAI_1_), .B2(keyinput_g30), .ZN(n6655) );
  OAI221_X1 U7583 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_1_), .C2(keyinput_g30), .A(n6655), .ZN(n6662) );
  AOI22_X1 U7584 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        REIP_REG_29__SCAN_IN), .B2(keyinput_g53), .ZN(n6656) );
  OAI221_X1 U7585 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_g53), .A(n6656), .ZN(n6661) );
  AOI22_X1 U7586 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_31_), .B2(
        keyinput_g0), .ZN(n6657) );
  OAI221_X1 U7587 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n6657), .ZN(n6660) );
  AOI22_X1 U7588 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n6658) );
  OAI221_X1 U7589 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(DATAI_23_), .C2(
        keyinput_g8), .A(n6658), .ZN(n6659) );
  NOR4_X1 U7590 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6663)
         );
  NAND4_X1 U7591 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6781)
         );
  INV_X1 U7592 ( .A(keyinput_f24), .ZN(n6774) );
  OAI22_X1 U7593 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f40), .B2(M_IO_N_REG_SCAN_IN), .ZN(n6667) );
  AOI221_X1 U7594 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_f40), .A(n6667), .ZN(n6674) );
  OAI22_X1 U7595 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(keyinput_f38), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6668) );
  AOI221_X1 U7596 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_f38), .A(n6668), .ZN(n6673) );
  OAI22_X1 U7597 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(keyinput_f7), .B2(
        DATAI_24_), .ZN(n6669) );
  AOI221_X1 U7598 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(DATAI_24_), .C2(
        keyinput_f7), .A(n6669), .ZN(n6672) );
  OAI22_X1 U7599 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(
        READREQUEST_REG_SCAN_IN), .B2(keyinput_f37), .ZN(n6670) );
  AOI221_X1 U7600 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(keyinput_f37), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6670), .ZN(n6671) );
  NAND4_X1 U7601 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6773)
         );
  OAI22_X1 U7602 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(keyinput_f42), .B2(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6675) );
  AOI221_X1 U7603 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f42), .A(n6675), .ZN(n6681)
         );
  OAI22_X1 U7604 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .ZN(n6676) );
  AOI221_X1 U7605 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(keyinput_f32), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6676), .ZN(n6680) );
  OAI22_X1 U7606 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(keyinput_f25), .B2(
        DATAI_6_), .ZN(n6677) );
  AOI221_X1 U7607 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(DATAI_6_), .C2(
        keyinput_f25), .A(n6677), .ZN(n6679) );
  XNOR2_X1 U7608 ( .A(DATAI_31_), .B(keyinput_f0), .ZN(n6678) );
  NAND4_X1 U7609 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6772)
         );
  OAI22_X1 U7610 ( .A1(n6684), .A2(keyinput_f19), .B1(n6683), .B2(keyinput_f29), .ZN(n6682) );
  AOI221_X1 U7611 ( .B1(n6684), .B2(keyinput_f19), .C1(keyinput_f29), .C2(
        n6683), .A(n6682), .ZN(n6687) );
  XOR2_X1 U7612 ( .A(keyinput_f48), .B(n6685), .Z(n6686) );
  OAI211_X1 U7613 ( .C1(n6689), .C2(keyinput_f51), .A(n6687), .B(n6686), .ZN(
        n6688) );
  AOI21_X1 U7614 ( .B1(n6689), .B2(keyinput_f51), .A(n6688), .ZN(n6714) );
  OAI22_X1 U7615 ( .A1(n6692), .A2(keyinput_f54), .B1(n6691), .B2(keyinput_f49), .ZN(n6690) );
  AOI221_X1 U7616 ( .B1(n6692), .B2(keyinput_f54), .C1(keyinput_f49), .C2(
        n6691), .A(n6690), .ZN(n6713) );
  INV_X1 U7617 ( .A(DATAI_14_), .ZN(n6694) );
  OAI22_X1 U7618 ( .A1(n4287), .A2(keyinput_f35), .B1(n6694), .B2(keyinput_f17), .ZN(n6693) );
  AOI221_X1 U7619 ( .B1(n4287), .B2(keyinput_f35), .C1(keyinput_f17), .C2(
        n6694), .A(n6693), .ZN(n6712) );
  INV_X1 U7620 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6696) );
  AOI22_X1 U7621 ( .A1(n6697), .A2(keyinput_f61), .B1(keyinput_f39), .B2(n6696), .ZN(n6695) );
  OAI221_X1 U7622 ( .B1(n6697), .B2(keyinput_f61), .C1(n6696), .C2(
        keyinput_f39), .A(n6695), .ZN(n6710) );
  INV_X1 U7623 ( .A(DATAI_25_), .ZN(n6700) );
  AOI22_X1 U7624 ( .A1(n6700), .A2(keyinput_f6), .B1(n6699), .B2(keyinput_f4), 
        .ZN(n6698) );
  OAI221_X1 U7625 ( .B1(n6700), .B2(keyinput_f6), .C1(n6699), .C2(keyinput_f4), 
        .A(n6698), .ZN(n6709) );
  AOI22_X1 U7626 ( .A1(n6703), .A2(keyinput_f62), .B1(keyinput_f36), .B2(n6702), .ZN(n6701) );
  OAI221_X1 U7627 ( .B1(n6703), .B2(keyinput_f62), .C1(n6702), .C2(
        keyinput_f36), .A(n6701), .ZN(n6708) );
  INV_X1 U7628 ( .A(DATAI_28_), .ZN(n6705) );
  AOI22_X1 U7629 ( .A1(n6706), .A2(keyinput_f55), .B1(keyinput_f3), .B2(n6705), 
        .ZN(n6704) );
  OAI221_X1 U7630 ( .B1(n6706), .B2(keyinput_f55), .C1(n6705), .C2(keyinput_f3), .A(n6704), .ZN(n6707) );
  NOR4_X1 U7631 ( .A1(n6710), .A2(n6709), .A3(n6708), .A4(n6707), .ZN(n6711)
         );
  NAND4_X1 U7632 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6771)
         );
  AOI22_X1 U7633 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_30_), .B2(
        keyinput_f1), .ZN(n6715) );
  OAI221_X1 U7634 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(DATAI_30_), .C2(
        keyinput_f1), .A(n6715), .ZN(n6725) );
  AOI22_X1 U7635 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(DATAI_15_), 
        .B2(keyinput_f16), .ZN(n6716) );
  OAI221_X1 U7636 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(DATAI_15_), 
        .C2(keyinput_f16), .A(n6716), .ZN(n6724) );
  AOI22_X1 U7637 ( .A1(n6719), .A2(keyinput_f27), .B1(keyinput_f50), .B2(n6718), .ZN(n6717) );
  OAI221_X1 U7638 ( .B1(n6719), .B2(keyinput_f27), .C1(n6718), .C2(
        keyinput_f50), .A(n6717), .ZN(n6723) );
  AOI22_X1 U7639 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(n6721), .B2(
        keyinput_f14), .ZN(n6720) );
  OAI221_X1 U7640 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(n6721), .C2(
        keyinput_f14), .A(n6720), .ZN(n6722) );
  NOR4_X1 U7641 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6769)
         );
  AOI22_X1 U7642 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .ZN(n6726) );
  OAI221_X1 U7643 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_f53), .A(n6726), .ZN(n6733) );
  AOI22_X1 U7644 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_f45), .B1(DATAI_1_), 
        .B2(keyinput_f30), .ZN(n6727) );
  OAI221_X1 U7645 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_f45), .C1(DATAI_1_), 
        .C2(keyinput_f30), .A(n6727), .ZN(n6732) );
  AOI22_X1 U7646 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_f59), .ZN(n6728) );
  OAI221_X1 U7647 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_f59), .A(n6728), .ZN(n6731) );
  AOI22_X1 U7648 ( .A1(keyinput_f34), .A2(BS16_N), .B1(DATAI_26_), .B2(
        keyinput_f5), .ZN(n6729) );
  OAI221_X1 U7649 ( .B1(keyinput_f34), .B2(BS16_N), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n6729), .ZN(n6730) );
  NOR4_X1 U7650 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6768)
         );
  INV_X1 U7651 ( .A(keyinput_f33), .ZN(n6735) );
  AOI22_X1 U7652 ( .A1(n6736), .A2(keyinput_f63), .B1(NA_N), .B2(n6735), .ZN(
        n6734) );
  OAI221_X1 U7653 ( .B1(n6736), .B2(keyinput_f63), .C1(n6735), .C2(NA_N), .A(
        n6734), .ZN(n6749) );
  AOI22_X1 U7654 ( .A1(n6739), .A2(keyinput_f58), .B1(keyinput_f28), .B2(n6738), .ZN(n6737) );
  OAI221_X1 U7655 ( .B1(n6739), .B2(keyinput_f58), .C1(n6738), .C2(
        keyinput_f28), .A(n6737), .ZN(n6748) );
  INV_X1 U7656 ( .A(DATAI_16_), .ZN(n6741) );
  AOI22_X1 U7657 ( .A1(n6742), .A2(keyinput_f56), .B1(keyinput_f15), .B2(n6741), .ZN(n6740) );
  OAI221_X1 U7658 ( .B1(n6742), .B2(keyinput_f56), .C1(n6741), .C2(
        keyinput_f15), .A(n6740), .ZN(n6747) );
  INV_X1 U7659 ( .A(DATAI_18_), .ZN(n6744) );
  AOI22_X1 U7660 ( .A1(n6745), .A2(keyinput_f57), .B1(keyinput_f13), .B2(n6744), .ZN(n6743) );
  OAI221_X1 U7661 ( .B1(n6745), .B2(keyinput_f57), .C1(n6744), .C2(
        keyinput_f13), .A(n6743), .ZN(n6746) );
  NOR4_X1 U7662 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n6767)
         );
  INV_X1 U7663 ( .A(DATAI_22_), .ZN(n6752) );
  AOI22_X1 U7664 ( .A1(n6752), .A2(keyinput_f9), .B1(keyinput_f47), .B2(n6751), 
        .ZN(n6750) );
  OAI221_X1 U7665 ( .B1(n6752), .B2(keyinput_f9), .C1(n6751), .C2(keyinput_f47), .A(n6750), .ZN(n6765) );
  INV_X1 U7666 ( .A(DATAI_21_), .ZN(n6755) );
  AOI22_X1 U7667 ( .A1(n6755), .A2(keyinput_f10), .B1(keyinput_f41), .B2(n6754), .ZN(n6753) );
  OAI221_X1 U7668 ( .B1(n6755), .B2(keyinput_f10), .C1(n6754), .C2(
        keyinput_f41), .A(n6753), .ZN(n6764) );
  AOI22_X1 U7669 ( .A1(n6758), .A2(keyinput_f43), .B1(keyinput_f44), .B2(n6757), .ZN(n6756) );
  OAI221_X1 U7670 ( .B1(n6758), .B2(keyinput_f43), .C1(n6757), .C2(
        keyinput_f44), .A(n6756), .ZN(n6763) );
  AOI22_X1 U7671 ( .A1(n6761), .A2(keyinput_f22), .B1(keyinput_f31), .B2(n6760), .ZN(n6759) );
  OAI221_X1 U7672 ( .B1(n6761), .B2(keyinput_f22), .C1(n6760), .C2(
        keyinput_f31), .A(n6759), .ZN(n6762) );
  NOR4_X1 U7673 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  NAND4_X1 U7674 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6770)
         );
  NOR4_X1 U7675 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6777)
         );
  OAI211_X1 U7676 ( .C1(n6774), .C2(n6777), .A(DATAI_7_), .B(keyinput_g24), 
        .ZN(n6779) );
  INV_X1 U7677 ( .A(keyinput_g24), .ZN(n6775) );
  OAI211_X1 U7678 ( .C1(n6777), .C2(keyinput_f24), .A(n6776), .B(n6775), .ZN(
        n6778) );
  NAND2_X1 U7679 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  OAI21_X1 U7680 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n6783) );
  XOR2_X1 U7681 ( .A(n6784), .B(n6783), .Z(U3445) );
  CLKBUF_X1 U34480 ( .A(n3180), .Z(n4114) );
  CLKBUF_X1 U3450 ( .A(n3626), .Z(n5454) );
  CLKBUF_X1 U34550 ( .A(n6100), .Z(n6571) );
  CLKBUF_X1 U3457 ( .A(n6099), .Z(n6090) );
  INV_X1 U3552 ( .A(n6069), .ZN(n6102) );
  OR3_X1 U3744 ( .A1(n6237), .A2(n4892), .A3(n4313), .ZN(n6785) );
endmodule

