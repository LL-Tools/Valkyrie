

module b21_C_SARLock_k_64_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4253, n4254, n4255, n4256, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063;

  INV_X4 U4759 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  BUF_X2 U4760 ( .A(n5784), .Z(n7527) );
  NAND2_X1 U4761 ( .A1(n5611), .A2(n5613), .ZN(n6844) );
  INV_X1 U4762 ( .A(n7848), .ZN(n7813) );
  CLKBUF_X2 U4763 ( .A(n5054), .Z(n4279) );
  INV_X2 U4764 ( .A(n5104), .ZN(n5446) );
  INV_X1 U4765 ( .A(n6488), .ZN(n7808) );
  NOR2_X1 U4766 ( .A1(n7012), .A2(n7286), .ZN(n7197) );
  AND2_X1 U4767 ( .A1(n5758), .A2(n6590), .ZN(n5843) );
  INV_X1 U4768 ( .A(n5463), .ZN(n5054) );
  XOR2_X1 U4769 ( .A(n8369), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8372) );
  CLKBUF_X2 U4770 ( .A(n5076), .Z(n5576) );
  CLKBUF_X3 U4771 ( .A(n7655), .Z(n4272) );
  INV_X1 U4772 ( .A(n9666), .ZN(n6777) );
  XNOR2_X1 U4773 ( .A(n9629), .B(n9651), .ZN(n7978) );
  INV_X1 U4774 ( .A(n6501), .ZN(n9675) );
  INV_X2 U4775 ( .A(n5067), .ZN(n5581) );
  INV_X1 U4776 ( .A(n5027), .ZN(n5510) );
  BUF_X1 U4777 ( .A(n6230), .Z(n7636) );
  NOR2_X1 U4778 ( .A1(n9368), .A2(n4468), .ZN(n9244) );
  BUF_X1 U4779 ( .A(n6184), .Z(n9651) );
  OAI21_X1 U4780 ( .B1(n4274), .B2(n6133), .A(n6085), .ZN(n6290) );
  OR2_X1 U4781 ( .A1(n6179), .A2(n6178), .ZN(n9629) );
  INV_X1 U4782 ( .A(n6096), .ZN(n6098) );
  AND3_X1 U4783 ( .A1(n4319), .A2(n4423), .A3(n4371), .ZN(n4253) );
  AND2_X1 U4784 ( .A1(n7710), .A2(n7709), .ZN(n4254) );
  OR2_X1 U4785 ( .A1(n5508), .A2(n5604), .ZN(n5721) );
  OAI21_X2 U4786 ( .B1(n7421), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7420), .ZN(
        n7463) );
  INV_X1 U4787 ( .A(n7957), .ZN(n7649) );
  XNOR2_X2 U4788 ( .A(n5473), .B(n5472), .ZN(n8433) );
  XNOR2_X2 U4789 ( .A(n5478), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5480) );
  OAI211_X2 U4790 ( .C1(n7569), .C2(n9496), .A(n6162), .B(n6161), .ZN(n6163)
         );
  INV_X2 U4791 ( .A(n5099), .ZN(n5027) );
  NOR2_X2 U4792 ( .A1(n6424), .A2(n6423), .ZN(n6436) );
  AOI21_X2 U4793 ( .B1(n8311), .B2(P2_REG1_REG_5__SCAN_IN), .A(n8312), .ZN(
        n6424) );
  AND2_X2 U4794 ( .A1(n6689), .A2(n6688), .ZN(n8327) );
  AND2_X4 U4795 ( .A1(n5007), .A2(n8781), .ZN(n5067) );
  AOI21_X2 U4796 ( .B1(n6437), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6436), .ZN(
        n6466) );
  NAND2_X1 U4797 ( .A1(n4254), .A2(n4255), .ZN(n8879) );
  CLKBUF_X1 U4798 ( .A(n8817), .Z(n4262) );
  CLKBUF_X1 U4799 ( .A(n8846), .Z(n4263) );
  NAND2_X1 U4800 ( .A1(n8503), .A2(n5506), .ZN(n8490) );
  NAND2_X1 U4801 ( .A1(n8520), .A2(n5503), .ZN(n8521) );
  MUX2_X1 U4802 ( .A(n7924), .B(n7923), .S(n7964), .Z(n7930) );
  NAND2_X1 U4803 ( .A1(n4857), .A2(n4854), .ZN(n9447) );
  NAND2_X1 U4804 ( .A1(n7755), .A2(n7754), .ZN(n9319) );
  INV_X1 U4805 ( .A(n9164), .ZN(n9127) );
  NOR3_X2 U4806 ( .A1(n7223), .A2(n7448), .A3(n4600), .ZN(n4597) );
  NAND2_X1 U4807 ( .A1(n6586), .A2(n4741), .ZN(n6925) );
  NAND2_X1 U4808 ( .A1(n7629), .A2(n7628), .ZN(n9354) );
  NAND2_X1 U4809 ( .A1(n6148), .A2(n9635), .ZN(n8894) );
  INV_X1 U4810 ( .A(n6629), .ZN(n9660) );
  INV_X2 U4811 ( .A(n7798), .ZN(n7824) );
  CLKBUF_X2 U4812 ( .A(n6227), .Z(n7848) );
  CLKBUF_X2 U4813 ( .A(n7858), .Z(n4276) );
  AND2_X2 U4814 ( .A1(n6238), .A2(n6164), .ZN(n7801) );
  INV_X1 U4815 ( .A(n6167), .ZN(n7798) );
  NAND2_X1 U4816 ( .A1(n6098), .A2(n6097), .ZN(n7858) );
  NAND2_X1 U4817 ( .A1(n6097), .A2(n6096), .ZN(n7655) );
  INV_X4 U4818 ( .A(n6156), .ZN(n6158) );
  NOR2_X1 U4819 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4419) );
  NAND2_X1 U4820 ( .A1(n7746), .A2(n7747), .ZN(n8805) );
  OAI21_X1 U4821 ( .B1(n7523), .B2(n8138), .A(n5866), .ZN(n8141) );
  OR2_X1 U4822 ( .A1(n5725), .A2(n4377), .ZN(n4376) );
  AOI21_X1 U4823 ( .B1(n5894), .B2(n9745), .A(n5893), .ZN(n8403) );
  NAND2_X1 U4824 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  AND2_X1 U4825 ( .A1(n8638), .A2(n8641), .ZN(n8720) );
  AND2_X1 U4826 ( .A1(n7953), .A2(n7952), .ZN(n7961) );
  NAND2_X1 U4827 ( .A1(n8490), .A2(n4308), .ZN(n8464) );
  NAND2_X1 U4828 ( .A1(n9145), .A2(n9144), .ZN(n9143) );
  NAND2_X1 U4829 ( .A1(n7860), .A2(n7859), .ZN(n7963) );
  NAND2_X1 U4830 ( .A1(n4776), .A2(n4785), .ZN(n8795) );
  OAI21_X1 U4831 ( .B1(n4444), .B2(n4443), .A(n7936), .ZN(n7944) );
  NAND2_X1 U4832 ( .A1(n8536), .A2(n5501), .ZN(n8520) );
  AOI21_X1 U4833 ( .B1(n4842), .B2(n4845), .A(n4841), .ZN(n4840) );
  NAND2_X1 U4834 ( .A1(n5456), .A2(n5455), .ZN(n7532) );
  NOR2_X1 U4835 ( .A1(n9265), .A2(n9264), .ZN(n9368) );
  AOI21_X1 U4836 ( .B1(n7362), .B2(n7361), .A(n7360), .ZN(n7363) );
  OAI21_X1 U4837 ( .B1(n5562), .B2(n4677), .A(n4675), .ZN(n5590) );
  XNOR2_X1 U4838 ( .A(n5562), .B(n5561), .ZN(n7805) );
  AND2_X1 U4839 ( .A1(n7440), .A2(n5285), .ZN(n8616) );
  NAND2_X1 U4840 ( .A1(n4761), .A2(n4762), .ZN(n7362) );
  AOI21_X1 U4841 ( .B1(n9447), .B2(n9448), .A(n9012), .ZN(n9277) );
  NAND2_X1 U4842 ( .A1(n5454), .A2(n5453), .ZN(n5562) );
  NAND2_X1 U4843 ( .A1(n5432), .A2(n5431), .ZN(n5452) );
  AND2_X1 U4844 ( .A1(n4549), .A2(n4548), .ZN(n9457) );
  NAND2_X1 U4845 ( .A1(n7545), .A2(n7544), .ZN(n9323) );
  INV_X1 U4846 ( .A(n7728), .ZN(n4255) );
  NAND2_X1 U4847 ( .A1(n7733), .A2(n7732), .ZN(n9328) );
  AND2_X1 U4848 ( .A1(n4459), .A2(n4458), .ZN(n6861) );
  NAND2_X1 U4849 ( .A1(n5802), .A2(n4735), .ZN(n6990) );
  NOR2_X1 U4850 ( .A1(n6729), .A2(n6728), .ZN(n6860) );
  NAND2_X1 U4851 ( .A1(n6925), .A2(n5795), .ZN(n6928) );
  OAI21_X1 U4852 ( .B1(n4833), .B2(n6636), .A(n4454), .ZN(n6729) );
  OR2_X2 U4853 ( .A1(n7222), .A2(n7226), .ZN(n7223) );
  NAND2_X1 U4854 ( .A1(n7610), .A2(n7609), .ZN(n9359) );
  AND2_X1 U4855 ( .A1(n9371), .A2(n9262), .ZN(n9046) );
  NAND2_X1 U4856 ( .A1(n7572), .A2(n7571), .ZN(n9371) );
  NAND2_X1 U4857 ( .A1(n4955), .A2(n4954), .ZN(n5303) );
  NAND2_X1 U4858 ( .A1(n5187), .A2(n5186), .ZN(n7157) );
  NAND2_X1 U4859 ( .A1(n6732), .A2(n6731), .ZN(n7063) );
  OR2_X1 U4860 ( .A1(n5485), .A2(n6911), .ZN(n5486) );
  AND2_X1 U4861 ( .A1(n5620), .A2(n6910), .ZN(n5484) );
  NAND2_X1 U4862 ( .A1(n6865), .A2(n6864), .ZN(n7123) );
  NAND2_X1 U4863 ( .A1(n5246), .A2(n4869), .ZN(n4940) );
  XNOR2_X1 U4864 ( .A(n5195), .B(n5194), .ZN(n6862) );
  NAND2_X1 U4865 ( .A1(n6647), .A2(n6646), .ZN(n7131) );
  NAND2_X1 U4866 ( .A1(n4471), .A2(n4474), .ZN(n4470) );
  NAND2_X1 U4867 ( .A1(n4805), .A2(n6543), .ZN(n9678) );
  OR2_X1 U4868 ( .A1(n5191), .A2(n5176), .ZN(n5178) );
  OAI211_X2 U4869 ( .C1(n5999), .C2(n5134), .A(n5133), .B(n5132), .ZN(n6839)
         );
  AND2_X1 U4870 ( .A1(n8314), .A2(n8315), .ZN(n8312) );
  NAND2_X1 U4871 ( .A1(n4904), .A2(n4903), .ZN(n5191) );
  INV_X1 U4872 ( .A(n4904), .ZN(n4471) );
  NAND2_X1 U4873 ( .A1(n5147), .A2(n4901), .ZN(n4904) );
  AND3_X1 U4874 ( .A1(n5065), .A2(n5064), .A3(n5063), .ZN(n9789) );
  NAND2_X1 U4875 ( .A1(n6109), .A2(n6108), .ZN(n6241) );
  INV_X1 U4876 ( .A(n6163), .ZN(n6789) );
  OAI211_X1 U4877 ( .C1(n4274), .C2(n6304), .A(n6303), .B(n6302), .ZN(n9666)
         );
  OR2_X1 U4878 ( .A1(n5103), .A2(n4588), .ZN(n9741) );
  OR2_X1 U4879 ( .A1(n6232), .A2(n6231), .ZN(n9627) );
  OR2_X1 U4880 ( .A1(n6194), .A2(n6193), .ZN(n8935) );
  AND4_X2 U4881 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n6847)
         );
  AND4_X1 U4882 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n7146)
         );
  CLKBUF_X1 U4883 ( .A(n5077), .Z(n5320) );
  CLKBUF_X1 U4884 ( .A(n4276), .Z(n7852) );
  INV_X1 U4885 ( .A(n6594), .ZN(n7525) );
  INV_X2 U4886 ( .A(n5077), .ZN(n5596) );
  INV_X1 U4887 ( .A(n5843), .ZN(n5784) );
  AND4_X1 U4888 ( .A1(n5143), .A2(n5142), .A3(n5141), .A4(n5140), .ZN(n7074)
         );
  INV_X1 U4889 ( .A(n5076), .ZN(n5134) );
  AND4_X1 U4890 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n6916)
         );
  INV_X1 U4891 ( .A(n5051), .ZN(n5291) );
  INV_X2 U4892 ( .A(n7798), .ZN(n4256) );
  NAND2_X1 U4893 ( .A1(n5110), .A2(n5109), .ZN(n5124) );
  OR2_X2 U4894 ( .A1(n9777), .A2(n5878), .ZN(n6594) );
  XNOR2_X1 U4895 ( .A(n5110), .B(n5109), .ZN(n6475) );
  AND2_X1 U4896 ( .A1(n6152), .A2(n6199), .ZN(n6164) );
  AND2_X1 U4897 ( .A1(n6658), .A2(n6199), .ZN(n6167) );
  NAND2_X1 U4898 ( .A1(n6132), .A2(n8110), .ZN(n6238) );
  OR3_X2 U4899 ( .A1(n7386), .A2(n7377), .A3(n7167), .ZN(n6199) );
  NAND2_X1 U4900 ( .A1(n6986), .A2(n6936), .ZN(n9777) );
  INV_X1 U4901 ( .A(n5480), .ZN(n6936) );
  NAND2_X1 U4902 ( .A1(n5967), .A2(n5966), .ZN(n4274) );
  XNOR2_X1 U4903 ( .A(n6095), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U4904 ( .A1(n5967), .A2(n5966), .ZN(n7569) );
  AND2_X1 U4905 ( .A1(n6094), .A2(n6093), .ZN(n6097) );
  AND2_X1 U4906 ( .A1(n4921), .A2(n4914), .ZN(n5194) );
  NAND2_X1 U4907 ( .A1(n4989), .A2(n4990), .ZN(n6368) );
  NAND2_X1 U4908 ( .A1(n6094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U4909 ( .A(n8781), .ZN(n5006) );
  OAI21_X1 U4910 ( .B1(n6092), .B2(n6091), .A(n6090), .ZN(n6093) );
  NAND2_X1 U4911 ( .A1(n5921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5922) );
  MUX2_X1 U4912 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4988), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4990) );
  AND2_X1 U4913 ( .A1(n6103), .A2(n6102), .ZN(n6658) );
  NAND2_X1 U4914 ( .A1(n4382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U4915 ( .A1(n5471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  NOR2_X1 U4916 ( .A1(n5527), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4983) );
  XNOR2_X1 U4917 ( .A(n4632), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8781) );
  OR2_X1 U4918 ( .A1(n8773), .A2(n5529), .ZN(n5005) );
  NAND2_X1 U4919 ( .A1(n5958), .A2(n5957), .ZN(n6092) );
  NAND2_X1 U4920 ( .A1(n5004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U4921 ( .A1(n6086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U4922 ( .A1(n4374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  INV_X2 U4923 ( .A(n9398), .ZN(n9402) );
  NAND2_X1 U4924 ( .A1(n4906), .A2(n4905), .ZN(n5177) );
  NAND2_X2 U4925 ( .A1(n6156), .A2(P2_U3152), .ZN(n8783) );
  NOR2_X1 U4926 ( .A1(n5920), .A2(n5996), .ZN(n5927) );
  NOR2_X1 U4927 ( .A1(n6012), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U4928 ( .A1(n4788), .A2(n5907), .ZN(n5996) );
  NOR2_X1 U4929 ( .A1(n4862), .A2(n4321), .ZN(n4861) );
  INV_X1 U4930 ( .A(n4863), .ZN(n4862) );
  XNOR2_X1 U4931 ( .A(n5062), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9423) );
  INV_X1 U4932 ( .A(n5993), .ZN(n4788) );
  NOR2_X1 U4933 ( .A1(n4739), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n4738) );
  AND2_X1 U4934 ( .A1(n5929), .A2(n5925), .ZN(n4863) );
  AND4_X1 U4935 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n5161), .ZN(n4636)
         );
  NAND4_X1 U4936 ( .A1(n4419), .A2(n4819), .A3(n5906), .A4(n4418), .ZN(n5993)
         );
  NOR2_X1 U4937 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5908) );
  INV_X1 U4938 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5929) );
  INV_X1 U4939 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5955) );
  NOR3_X1 U4940 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n4980) );
  INV_X1 U4941 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6121) );
  INV_X1 U4942 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5161) );
  INV_X1 U4943 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6021) );
  INV_X2 U4944 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4945 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6336) );
  NOR2_X1 U4946 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4638) );
  NOR2_X1 U4947 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4639) );
  INV_X1 U4948 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5954) );
  NOR2_X1 U4949 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4637) );
  INV_X1 U4950 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5906) );
  NOR2_X2 U4951 ( .A1(n9460), .A2(n9371), .ZN(n9278) );
  OR2_X1 U4952 ( .A1(n9459), .A2(n10034), .ZN(n9460) );
  NAND2_X1 U4953 ( .A1(n4811), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U4954 ( .A1(n8832), .A2(n4260), .ZN(n4258) );
  AND2_X1 U4955 ( .A1(n4258), .A2(n4259), .ZN(n8878) );
  OR2_X1 U4956 ( .A1(n4255), .A2(n7709), .ZN(n4259) );
  AND2_X1 U4957 ( .A1(n8833), .A2(n7728), .ZN(n4260) );
  CLKBUF_X1 U4958 ( .A(n6207), .Z(n4261) );
  OAI21_X1 U4959 ( .B1(n4268), .B2(n4304), .A(n4771), .ZN(n4264) );
  AOI21_X1 U4960 ( .B1(n7362), .B2(n7361), .A(n7360), .ZN(n4265) );
  AOI21_X1 U4961 ( .B1(n8805), .B2(n8808), .A(n8807), .ZN(n4266) );
  AOI21_X1 U4962 ( .B1(n8805), .B2(n8808), .A(n8807), .ZN(n4267) );
  INV_X1 U4963 ( .A(n4770), .ZN(n4268) );
  INV_X1 U4964 ( .A(n6003), .ZN(n4269) );
  OAI21_X1 U4965 ( .B1(n6493), .B2(n4304), .A(n4771), .ZN(n6799) );
  AOI21_X1 U4966 ( .B1(n8805), .B2(n8808), .A(n8807), .ZN(n8863) );
  OAI21_X1 U4967 ( .B1(n6487), .B2(n6486), .A(n6485), .ZN(n6493) );
  XNOR2_X1 U4968 ( .A(n5922), .B(n5954), .ZN(n7386) );
  AND2_X1 U4969 ( .A1(n6238), .A2(n6164), .ZN(n4270) );
  AND2_X1 U4970 ( .A1(n6658), .A2(n6199), .ZN(n4271) );
  NAND2_X1 U4971 ( .A1(n6212), .A2(n6211), .ZN(n6294) );
  NOR2_X2 U4972 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5038) );
  NAND2_X1 U4973 ( .A1(n5967), .A2(n5966), .ZN(n4273) );
  NAND2_X2 U4974 ( .A1(n5858), .A2(n5857), .ZN(n5861) );
  NAND2_X1 U4975 ( .A1(n5051), .A2(n5367), .ZN(n4275) );
  NAND2_X1 U4976 ( .A1(n5095), .A2(n9803), .ZN(n6912) );
  INV_X1 U4977 ( .A(n5095), .ZN(n6917) );
  AND3_X4 U4978 ( .A1(n4608), .A2(n4607), .A3(n4372), .ZN(n9784) );
  OAI222_X1 U4979 ( .A1(n9402), .A2(n7387), .B1(P1_U3084), .B2(n4269), .C1(
        n7772), .C2(n9404), .ZN(P1_U3327) );
  NAND2_X1 U4980 ( .A1(n6098), .A2(n6097), .ZN(n4277) );
  OAI21_X2 U4981 ( .B1(n6845), .B2(n6844), .A(n5611), .ZN(n6602) );
  NAND2_X1 U4982 ( .A1(n6098), .A2(n7514), .ZN(n6227) );
  OAI21_X2 U4983 ( .B1(n7218), .B2(n5495), .A(n5647), .ZN(n7205) );
  NAND2_X2 U4984 ( .A1(n7688), .A2(n7687), .ZN(n8832) );
  NOR3_X4 U4985 ( .A1(n8481), .A2(n4604), .A3(n8424), .ZN(n4606) );
  XNOR2_X2 U4986 ( .A(n5005), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8778) );
  NOR2_X2 U4987 ( .A1(n5914), .A2(n5913), .ZN(n5947) );
  CLKBUF_X1 U4988 ( .A(n5966), .Z(n4278) );
  XNOR2_X1 U4989 ( .A(n5958), .B(n5956), .ZN(n5966) );
  NAND2_X1 U4990 ( .A1(n6155), .A2(n6154), .ZN(n6172) );
  XNOR2_X1 U4991 ( .A(n6166), .B(n7799), .ZN(n6170) );
  NAND2_X1 U4992 ( .A1(n6096), .A2(n7514), .ZN(n6230) );
  NAND2_X1 U4993 ( .A1(n6299), .A2(n6298), .ZN(n6487) );
  AOI21_X1 U4994 ( .B1(n4573), .B2(n5702), .A(n4572), .ZN(n5703) );
  AND2_X1 U4995 ( .A1(n5701), .A2(n5721), .ZN(n4572) );
  AND2_X1 U4996 ( .A1(n8064), .A2(n8060), .ZN(n4435) );
  INV_X1 U4997 ( .A(n5209), .ZN(n4927) );
  INV_X1 U4998 ( .A(n4923), .ZN(n4475) );
  INV_X1 U4999 ( .A(n5179), .ZN(n4919) );
  AND2_X1 U5000 ( .A1(n4413), .A2(n4412), .ZN(n5714) );
  AOI21_X1 U5001 ( .B1(n8542), .B2(n4657), .A(n5348), .ZN(n4656) );
  INV_X1 U5002 ( .A(n4658), .ZN(n4657) );
  NAND2_X1 U5003 ( .A1(n4932), .A2(n4931), .ZN(n5232) );
  AND2_X1 U5004 ( .A1(n9472), .A2(n9435), .ZN(n9009) );
  NAND2_X1 U5005 ( .A1(n9702), .A2(n7121), .ZN(n4458) );
  INV_X1 U5006 ( .A(n6860), .ZN(n4459) );
  NAND2_X1 U5007 ( .A1(n7890), .A2(n4363), .ZN(n4362) );
  NOR2_X1 U5008 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  INV_X1 U5009 ( .A(n7888), .ZN(n4364) );
  INV_X1 U5010 ( .A(n7889), .ZN(n4365) );
  NAND2_X1 U5011 ( .A1(n4406), .A2(n4408), .ZN(n4404) );
  NAND2_X1 U5012 ( .A1(n5703), .A2(n4406), .ZN(n4405) );
  AND2_X1 U5013 ( .A1(n4407), .A2(n5726), .ZN(n4406) );
  AOI21_X1 U5014 ( .B1(n4285), .B2(n8064), .A(n7964), .ZN(n4425) );
  INV_X1 U5015 ( .A(n9085), .ZN(n4433) );
  NAND2_X1 U5016 ( .A1(n9034), .A2(n8926), .ZN(n9065) );
  NAND2_X1 U5017 ( .A1(n4960), .A2(n4959), .ZN(n4689) );
  INV_X1 U5018 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4984) );
  OR2_X1 U5019 ( .A1(n8400), .A2(n6378), .ZN(n5727) );
  OR2_X1 U5020 ( .A1(n8456), .A2(n8436), .ZN(n5699) );
  INV_X1 U5021 ( .A(n8681), .ZN(n4592) );
  NOR2_X1 U5022 ( .A1(n7318), .A2(n4646), .ZN(n4645) );
  INV_X1 U5023 ( .A(n4648), .ZN(n4646) );
  NAND2_X1 U5024 ( .A1(n8287), .A2(n9820), .ZN(n5631) );
  NAND3_X1 U5025 ( .A1(n5078), .A2(n4636), .A3(n4973), .ZN(n5247) );
  NOR2_X1 U5026 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4973) );
  OR2_X1 U5027 ( .A1(n9442), .A2(n9454), .ZN(n9011) );
  OR2_X1 U5028 ( .A1(n9433), .A2(n9434), .ZN(n4549) );
  NAND2_X1 U5029 ( .A1(n4456), .A2(n7185), .ZN(n7186) );
  OR2_X1 U5030 ( .A1(n7286), .A2(n8928), .ZN(n7185) );
  NAND2_X1 U5031 ( .A1(n4457), .A2(n4823), .ZN(n4456) );
  AOI21_X1 U5032 ( .B1(n4824), .B2(n7009), .A(n4320), .ZN(n4823) );
  NAND2_X1 U5033 ( .A1(n5452), .A2(n5451), .ZN(n5454) );
  OAI21_X1 U5034 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n4692) );
  INV_X1 U5035 ( .A(n5350), .ZN(n4704) );
  AOI21_X1 U5036 ( .B1(n4696), .B2(n4699), .A(n4695), .ZN(n4694) );
  AOI21_X1 U5037 ( .B1(n4698), .B2(n4700), .A(n4697), .ZN(n4696) );
  INV_X1 U5038 ( .A(n4949), .ZN(n4697) );
  INV_X1 U5039 ( .A(n4702), .ZN(n4698) );
  NAND2_X1 U5040 ( .A1(n4933), .A2(n4932), .ZN(n5246) );
  NAND2_X1 U5041 ( .A1(n4470), .A2(n4306), .ZN(n4933) );
  INV_X1 U5042 ( .A(n5232), .ZN(n4479) );
  NOR2_X1 U5043 ( .A1(n4874), .A2(n4922), .ZN(n4923) );
  XNOR2_X1 U5044 ( .A(n4925), .B(SI_11_), .ZN(n5209) );
  NAND2_X1 U5045 ( .A1(n5177), .A2(n4908), .ZN(n5176) );
  AOI21_X2 U5046 ( .B1(n5124), .B2(n4900), .A(n4872), .ZN(n5147) );
  OAI211_X1 U5047 ( .C1(n4809), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4706), .B(
        n4705), .ZN(n4882) );
  OR2_X1 U5048 ( .A1(n4810), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U5049 ( .A1(n5049), .A2(n6083), .ZN(n4880) );
  AND2_X1 U5050 ( .A1(n8138), .A2(n4727), .ZN(n4726) );
  NAND2_X1 U5051 ( .A1(n7516), .A2(n5860), .ZN(n4727) );
  NAND2_X1 U5052 ( .A1(n5586), .A2(n4311), .ZN(n4617) );
  AOI21_X1 U5053 ( .B1(n4571), .B2(n4570), .A(n5747), .ZN(n5725) );
  INV_X1 U5054 ( .A(n5722), .ZN(n4570) );
  NAND2_X1 U5055 ( .A1(n5724), .A2(n5723), .ZN(n4571) );
  AND4_X1 U5056 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), .ZN(n7431)
         );
  NAND2_X2 U5057 ( .A1(n8778), .A2(n5006), .ZN(n5463) );
  NAND2_X1 U5058 ( .A1(n5727), .A2(n5726), .ZN(n5888) );
  AND2_X1 U5059 ( .A1(n8501), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U5060 ( .A1(n4652), .A2(n4651), .ZN(n4650) );
  OR2_X1 U5061 ( .A1(n8511), .A2(n8493), .ZN(n4651) );
  OR2_X1 U5062 ( .A1(n8681), .A2(n8567), .ZN(n8519) );
  AND2_X1 U5063 ( .A1(n8681), .A2(n8276), .ZN(n4658) );
  AOI21_X1 U5064 ( .B1(n4612), .B2(n4614), .A(n4610), .ZN(n4609) );
  NAND2_X1 U5065 ( .A1(n5496), .A2(n4612), .ZN(n4611) );
  INV_X1 U5066 ( .A(n5670), .ZN(n4610) );
  AND2_X1 U5067 ( .A1(n7318), .A2(n5652), .ZN(n4631) );
  AND2_X1 U5068 ( .A1(n5188), .A2(n5168), .ZN(n4668) );
  NAND2_X1 U5069 ( .A1(n5051), .A2(n5367), .ZN(n5077) );
  AND2_X1 U5070 ( .A1(n5051), .A2(n6156), .ZN(n5076) );
  NAND2_X2 U5071 ( .A1(n6359), .A2(n6368), .ZN(n5051) );
  INV_X1 U5073 ( .A(n7747), .ZN(n7748) );
  INV_X1 U5074 ( .A(n7799), .ZN(n7822) );
  INV_X2 U5075 ( .A(n7636), .ZN(n7853) );
  XNOR2_X1 U5076 ( .A(n9314), .B(n8927), .ZN(n9109) );
  AOI21_X1 U5077 ( .B1(n4844), .B2(n4843), .A(n4313), .ZN(n4842) );
  INV_X1 U5078 ( .A(n4848), .ZN(n4843) );
  NOR2_X1 U5079 ( .A1(n9159), .A2(n9060), .ZN(n9145) );
  INV_X1 U5080 ( .A(n9186), .ZN(n4493) );
  AOI21_X1 U5081 ( .B1(n4808), .B2(n9056), .A(n7970), .ZN(n4807) );
  AOI21_X1 U5082 ( .B1(n4283), .B2(n9021), .A(n4345), .ZN(n4851) );
  AOI21_X1 U5083 ( .B1(n9228), .B2(n9238), .A(n4467), .ZN(n9215) );
  AND2_X1 U5084 ( .A1(n9354), .A2(n9017), .ZN(n4467) );
  OAI22_X1 U5085 ( .A1(n9277), .A2(n9013), .B1(n9371), .B2(n9453), .ZN(n9265)
         );
  NAND2_X1 U5086 ( .A1(n6733), .A2(n4834), .ZN(n4833) );
  NAND2_X1 U5087 ( .A1(n4836), .A2(n4455), .ZN(n4454) );
  INV_X1 U5088 ( .A(n4835), .ZN(n4834) );
  OR2_X1 U5089 ( .A1(n8068), .A2(n9512), .ZN(n9289) );
  INV_X1 U5090 ( .A(n9299), .ZN(n4813) );
  NAND2_X1 U5091 ( .A1(n7183), .A2(n7182), .ZN(n9472) );
  NAND2_X1 U5092 ( .A1(n6089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5093 ( .A1(n4870), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U5094 ( .A1(n8222), .A2(n8221), .B1(n5842), .B2(n5841), .ZN(n8174)
         );
  NAND2_X1 U5095 ( .A1(n4309), .A2(n8603), .ZN(n8638) );
  INV_X1 U5096 ( .A(n9147), .ZN(n9112) );
  OAI21_X1 U5097 ( .B1(n7872), .B2(n7871), .A(n8020), .ZN(n4446) );
  NAND2_X1 U5098 ( .A1(n4559), .A2(n4557), .ZN(n5640) );
  AOI21_X1 U5099 ( .B1(n4567), .B2(n5633), .A(n4558), .ZN(n4557) );
  INV_X1 U5100 ( .A(n5643), .ZN(n4558) );
  NAND2_X1 U5101 ( .A1(n4362), .A2(n4361), .ZN(n7894) );
  AND2_X1 U5102 ( .A1(n8038), .A2(n8085), .ZN(n4361) );
  NAND2_X1 U5103 ( .A1(n9252), .A2(n7917), .ZN(n4438) );
  INV_X1 U5104 ( .A(n7870), .ZN(n7918) );
  NOR2_X1 U5105 ( .A1(n4441), .A2(n4440), .ZN(n4439) );
  INV_X1 U5106 ( .A(n9264), .ZN(n4440) );
  INV_X1 U5107 ( .A(n7915), .ZN(n4441) );
  NOR2_X1 U5108 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  NOR2_X1 U5109 ( .A1(n8577), .A2(n5719), .ZN(n4580) );
  INV_X1 U5110 ( .A(n5728), .ZN(n4581) );
  NAND2_X1 U5111 ( .A1(n4394), .A2(n5684), .ZN(n4393) );
  INV_X1 U5112 ( .A(n4395), .ZN(n4394) );
  AOI21_X1 U5113 ( .B1(n4291), .B2(n4398), .A(n4396), .ZN(n4395) );
  INV_X1 U5114 ( .A(n4327), .ZN(n4396) );
  NAND2_X1 U5115 ( .A1(n4583), .A2(n5719), .ZN(n4582) );
  NAND2_X1 U5116 ( .A1(n4585), .A2(n4584), .ZN(n4583) );
  AND2_X1 U5117 ( .A1(n8559), .A2(n5673), .ZN(n4584) );
  AND2_X1 U5118 ( .A1(n4391), .A2(n4579), .ZN(n4387) );
  NOR2_X1 U5119 ( .A1(n8488), .A2(n4392), .ZN(n4391) );
  NAND2_X1 U5120 ( .A1(n4398), .A2(n5684), .ZN(n4392) );
  NAND2_X1 U5121 ( .A1(n7921), .A2(n4442), .ZN(n7920) );
  AND2_X1 U5122 ( .A1(n7974), .A2(n7996), .ZN(n4442) );
  INV_X1 U5123 ( .A(n5707), .ZN(n4414) );
  NAND2_X1 U5124 ( .A1(n4411), .A2(n5708), .ZN(n4410) );
  NAND2_X1 U5125 ( .A1(n4414), .A2(n4415), .ZN(n4411) );
  OR2_X1 U5126 ( .A1(n4410), .A2(n4414), .ZN(n4403) );
  NAND2_X1 U5127 ( .A1(n7944), .A2(n9062), .ZN(n7945) );
  NAND2_X1 U5128 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  INV_X1 U5129 ( .A(n8060), .ZN(n4431) );
  OR2_X1 U5130 ( .A1(n9301), .A2(n9085), .ZN(n8059) );
  OR2_X1 U5131 ( .A1(n9034), .A2(n8926), .ZN(n8053) );
  OR2_X1 U5132 ( .A1(n9339), .A2(n9204), .ZN(n7972) );
  NOR2_X1 U5133 ( .A1(n9310), .A2(n9314), .ZN(n4498) );
  INV_X1 U5134 ( .A(n5566), .ZN(n4679) );
  INV_X1 U5135 ( .A(n5561), .ZN(n4676) );
  AOI21_X1 U5136 ( .B1(n4687), .B2(n4686), .A(n4324), .ZN(n4685) );
  INV_X1 U5137 ( .A(n4959), .ZN(n4686) );
  INV_X1 U5138 ( .A(n4963), .ZN(n4690) );
  OAI21_X1 U5139 ( .B1(n5367), .B2(P1_DATAO_REG_10__SCAN_IN), .A(n4366), .ZN(
        n4912) );
  NAND2_X1 U5140 ( .A1(n5367), .A2(n6024), .ZN(n4366) );
  NAND2_X1 U5141 ( .A1(n8385), .A2(n5480), .ZN(n4619) );
  NAND2_X1 U5142 ( .A1(n5027), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5028) );
  INV_X1 U5143 ( .A(n8778), .ZN(n5007) );
  NAND2_X1 U5144 ( .A1(n4605), .A2(n8734), .ZN(n4604) );
  OR2_X1 U5145 ( .A1(n8443), .A2(n8184), .ZN(n5698) );
  NOR2_X1 U5146 ( .A1(n8456), .A2(n8473), .ZN(n4605) );
  OR2_X1 U5147 ( .A1(n8473), .A2(n8213), .ZN(n5694) );
  NOR2_X1 U5148 ( .A1(n8688), .A2(n8590), .ZN(n4593) );
  OR2_X1 U5149 ( .A1(n8629), .A2(n8595), .ZN(n5670) );
  NOR2_X1 U5150 ( .A1(n7503), .A2(n7210), .ZN(n4601) );
  OR2_X1 U5151 ( .A1(n7210), .A2(n7304), .ZN(n5652) );
  NAND2_X1 U5152 ( .A1(n4587), .A2(n4586), .ZN(n5732) );
  INV_X1 U5153 ( .A(n5103), .ZN(n4587) );
  AND2_X1 U5154 ( .A1(n5106), .A2(n9811), .ZN(n4586) );
  OR2_X1 U5155 ( .A1(n8289), .A2(n9789), .ZN(n5611) );
  OR2_X1 U5156 ( .A1(n7210), .A2(n8282), .ZN(n4648) );
  OR2_X1 U5157 ( .A1(n7208), .A2(n7209), .ZN(n4647) );
  INV_X1 U5158 ( .A(n9784), .ZN(n5041) );
  AND2_X1 U5159 ( .A1(n4786), .A2(n7566), .ZN(n4785) );
  NAND2_X1 U5160 ( .A1(n7555), .A2(n7554), .ZN(n4786) );
  NAND2_X1 U5161 ( .A1(n7861), .A2(n7963), .ZN(n8064) );
  OR2_X1 U5162 ( .A1(n9306), .A2(n9100), .ZN(n9066) );
  NAND2_X1 U5163 ( .A1(n4525), .A2(n4523), .ZN(n9083) );
  AND2_X1 U5164 ( .A1(n4533), .A2(n4524), .ZN(n4523) );
  INV_X1 U5165 ( .A(n4534), .ZN(n4533) );
  AND2_X1 U5166 ( .A1(n9066), .A2(n8055), .ZN(n9082) );
  NAND2_X1 U5167 ( .A1(n4529), .A2(n9062), .ZN(n4528) );
  INV_X1 U5168 ( .A(n4530), .ZN(n4529) );
  NAND2_X1 U5169 ( .A1(n9319), .A2(n9112), .ZN(n7968) );
  OR2_X1 U5170 ( .A1(n9049), .A2(n4803), .ZN(n4800) );
  NOR2_X1 U5171 ( .A1(n4803), .A2(n9046), .ZN(n4802) );
  NAND2_X1 U5172 ( .A1(n7989), .A2(n4825), .ZN(n4824) );
  INV_X1 U5173 ( .A(n4826), .ZN(n4825) );
  OR2_X1 U5174 ( .A1(n7131), .A2(n6655), .ZN(n8038) );
  INV_X1 U5175 ( .A(n6651), .ZN(n6381) );
  NAND2_X1 U5176 ( .A1(n6379), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6555) );
  INV_X1 U5177 ( .A(n6497), .ZN(n6379) );
  NAND2_X1 U5178 ( .A1(n9678), .A2(n6716), .ZN(n7888) );
  NAND2_X1 U5179 ( .A1(n9129), .A2(n4496), .ZN(n9086) );
  XNOR2_X1 U5180 ( .A(n5590), .B(n5589), .ZN(n5587) );
  NAND2_X1 U5181 ( .A1(n4692), .A2(n5430), .ZN(n5432) );
  OAI21_X1 U5182 ( .B1(n5398), .B2(n5397), .A(n5396), .ZN(n5416) );
  NAND2_X1 U5183 ( .A1(n5383), .A2(n5382), .ZN(n5398) );
  NAND2_X1 U5184 ( .A1(n5381), .A2(n5380), .ZN(n5383) );
  NAND2_X1 U5185 ( .A1(n6057), .A2(n6059), .ZN(n4795) );
  NAND2_X1 U5186 ( .A1(n5337), .A2(n5336), .ZN(n5349) );
  NAND2_X1 U5187 ( .A1(n4949), .A2(n4948), .ZN(n5275) );
  XNOR2_X1 U5188 ( .A(n4941), .B(SI_14_), .ZN(n5260) );
  NAND2_X1 U5189 ( .A1(n4910), .A2(SI_9_), .ZN(n5179) );
  NOR2_X1 U5190 ( .A1(n4790), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4789) );
  XNOR2_X1 U5191 ( .A(n4902), .B(SI_7_), .ZN(n5146) );
  XNOR2_X1 U5192 ( .A(n4897), .B(SI_6_), .ZN(n5125) );
  INV_X1 U5193 ( .A(n5059), .ZN(n4450) );
  INV_X1 U5194 ( .A(n4881), .ZN(n4453) );
  NAND2_X1 U5195 ( .A1(n4876), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4811) );
  INV_X1 U5196 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4876) );
  OAI21_X2 U5197 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4812), .ZN(n4809) );
  AND2_X1 U5198 ( .A1(n7524), .A2(n7521), .ZN(n8138) );
  AOI21_X1 U5199 ( .B1(n7301), .B2(n4733), .A(n4732), .ZN(n4731) );
  INV_X1 U5200 ( .A(n5819), .ZN(n4732) );
  NOR2_X1 U5201 ( .A1(n7301), .A2(n4733), .ZN(n4730) );
  XNOR2_X1 U5202 ( .A(n8473), .B(n7527), .ZN(n5853) );
  XNOR2_X1 U5203 ( .A(n6533), .B(n5784), .ZN(n8125) );
  INV_X1 U5204 ( .A(n5934), .ZN(n5774) );
  AND2_X1 U5205 ( .A1(n4718), .A2(n4338), .ZN(n4716) );
  NAND2_X1 U5206 ( .A1(n4719), .A2(n5833), .ZN(n4718) );
  NAND2_X1 U5207 ( .A1(n8206), .A2(n4284), .ZN(n4717) );
  AND2_X1 U5208 ( .A1(n4381), .A2(n4380), .ZN(n4379) );
  INV_X1 U5209 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4380) );
  INV_X1 U5210 ( .A(n5749), .ZN(n4377) );
  NAND2_X1 U5211 ( .A1(n4621), .A2(n4627), .ZN(n4620) );
  INV_X1 U5212 ( .A(n5706), .ZN(n4627) );
  NAND2_X1 U5213 ( .A1(n4624), .A2(n5702), .ZN(n8415) );
  XNOR2_X1 U5214 ( .A(n8424), .B(n8437), .ZN(n8421) );
  AND2_X1 U5215 ( .A1(n5412), .A2(n5411), .ZN(n8436) );
  OR2_X1 U5216 ( .A1(n5424), .A2(n5423), .ZN(n5442) );
  NOR2_X1 U5217 ( .A1(n8481), .A2(n4603), .ZN(n8454) );
  INV_X1 U5218 ( .A(n4605), .ZN(n4603) );
  AND2_X1 U5219 ( .A1(n5694), .A2(n5695), .ZN(n8470) );
  NOR2_X1 U5220 ( .A1(n8481), .A2(n8473), .ZN(n8472) );
  INV_X1 U5221 ( .A(n4656), .ZN(n4655) );
  AOI21_X1 U5222 ( .B1(n4656), .B2(n4658), .A(n4328), .ZN(n4654) );
  AOI21_X1 U5223 ( .B1(n4662), .B2(n4664), .A(n4329), .ZN(n4661) );
  AND2_X1 U5224 ( .A1(n8519), .A2(n5677), .ZN(n8542) );
  INV_X1 U5225 ( .A(n4663), .ZN(n4662) );
  OAI22_X1 U5226 ( .A1(n5331), .A2(n4282), .B1(n8590), .B2(n8277), .ZN(n4663)
         );
  OR2_X1 U5227 ( .A1(n5331), .A2(n8599), .ZN(n4664) );
  NAND2_X1 U5228 ( .A1(n5001), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5324) );
  INV_X1 U5229 ( .A(n5309), .ZN(n5001) );
  AND2_X1 U5230 ( .A1(n8577), .A2(n5673), .ZN(n8599) );
  OR2_X1 U5231 ( .A1(n8600), .A2(n8599), .ZN(n4665) );
  AND4_X1 U5232 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n8622)
         );
  OAI21_X1 U5233 ( .B1(n7208), .B2(n4643), .A(n4641), .ZN(n7441) );
  AOI21_X1 U5234 ( .B1(n5274), .B2(n4289), .A(n4318), .ZN(n4641) );
  OR2_X1 U5235 ( .A1(n7493), .A2(n7446), .ZN(n7442) );
  NAND2_X1 U5236 ( .A1(n4647), .A2(n4645), .ZN(n7484) );
  NOR2_X1 U5237 ( .A1(n5273), .A2(n4630), .ZN(n4629) );
  INV_X1 U5238 ( .A(n5658), .ZN(n4630) );
  AND2_X1 U5239 ( .A1(n5652), .A2(n5651), .ZN(n7209) );
  AOI21_X1 U5240 ( .B1(n5151), .B2(n5150), .A(n4873), .ZN(n7077) );
  INV_X1 U5241 ( .A(n6754), .ZN(n5150) );
  NAND2_X1 U5242 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  OR2_X1 U5243 ( .A1(n9826), .A2(n8433), .ZN(n5870) );
  NOR2_X1 U5244 ( .A1(n8543), .A2(n8542), .ZN(n8685) );
  NAND2_X1 U5245 ( .A1(n5167), .A2(n5166), .ZN(n7233) );
  NAND2_X1 U5246 ( .A1(n4745), .A2(n4744), .ZN(n4743) );
  NOR2_X1 U5247 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4744) );
  NOR2_X1 U5248 ( .A1(n5262), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5276) );
  CLKBUF_X1 U5249 ( .A(n5247), .Z(n5248) );
  NAND2_X1 U5250 ( .A1(n7750), .A2(n7751), .ZN(n4759) );
  NAND3_X1 U5251 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6497) );
  INV_X1 U5252 ( .A(n7111), .ZN(n4765) );
  INV_X1 U5253 ( .A(n7106), .ZN(n4763) );
  NAND2_X1 U5254 ( .A1(n4299), .A2(n6165), .ZN(n6166) );
  INV_X1 U5255 ( .A(n6492), .ZN(n4772) );
  AND2_X1 U5256 ( .A1(n4760), .A2(n4759), .ZN(n4758) );
  OR2_X1 U5257 ( .A1(n8840), .A2(n4757), .ZN(n4756) );
  INV_X1 U5258 ( .A(n4760), .ZN(n4757) );
  INV_X1 U5259 ( .A(n4758), .ZN(n4754) );
  NOR2_X1 U5260 ( .A1(n4755), .A2(n4751), .ZN(n4750) );
  INV_X1 U5261 ( .A(n8865), .ZN(n4751) );
  INV_X1 U5262 ( .A(n4756), .ZN(n4755) );
  NAND2_X1 U5263 ( .A1(n7961), .A2(n4424), .ZN(n4423) );
  AND2_X1 U5264 ( .A1(n9294), .A2(n9002), .ZN(n8104) );
  NOR2_X1 U5265 ( .A1(n9491), .A2(n4305), .ZN(n9506) );
  NOR2_X1 U5266 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4821) );
  NOR2_X1 U5267 ( .A1(n9579), .A2(n4346), .ZN(n9598) );
  OAI21_X1 U5268 ( .B1(n7558), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7294), .ZN(
        n8957) );
  NOR2_X1 U5269 ( .A1(n8982), .A2(n4509), .ZN(n9607) );
  AND2_X1 U5270 ( .A1(n8987), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4509) );
  AND2_X1 U5271 ( .A1(n9129), .A2(n4332), .ZN(n9073) );
  NAND2_X1 U5272 ( .A1(n9062), .A2(n7968), .ZN(n9124) );
  INV_X1 U5273 ( .A(n9026), .ZN(n4846) );
  NOR2_X1 U5274 ( .A1(n4849), .A2(n9027), .ZN(n4848) );
  INV_X1 U5275 ( .A(n9024), .ZN(n4849) );
  AND2_X1 U5276 ( .A1(n4537), .A2(n4331), .ZN(n9159) );
  OAI21_X1 U5278 ( .B1(n4494), .B2(n9054), .A(n9053), .ZN(n9186) );
  NOR2_X1 U5279 ( .A1(n9186), .A2(n9187), .ZN(n9185) );
  NAND2_X1 U5280 ( .A1(n9212), .A2(n9219), .ZN(n4852) );
  OAI22_X1 U5281 ( .A1(n9215), .A2(n9019), .B1(n9225), .B2(n9241), .ZN(n9198)
         );
  NOR2_X1 U5282 ( .A1(n4505), .A2(n9048), .ZN(n4804) );
  NOR2_X1 U5283 ( .A1(n9044), .A2(n9046), .ZN(n4505) );
  INV_X1 U5284 ( .A(n9047), .ZN(n4803) );
  NOR2_X1 U5285 ( .A1(n9448), .A2(n9449), .ZN(n4548) );
  INV_X1 U5286 ( .A(n4804), .ZN(n4797) );
  AND2_X1 U5287 ( .A1(n8023), .A2(n9050), .ZN(n9252) );
  AND2_X1 U5288 ( .A1(n9365), .A2(n9014), .ZN(n4468) );
  NOR2_X1 U5289 ( .A1(n9283), .A2(n9046), .ZN(n9259) );
  OR2_X1 U5290 ( .A1(n7576), .A2(n7575), .ZN(n7594) );
  INV_X1 U5291 ( .A(n9436), .ZN(n9286) );
  INV_X1 U5292 ( .A(n4855), .ZN(n4854) );
  OAI21_X1 U5293 ( .B1(n4859), .B2(n4856), .A(n9011), .ZN(n4855) );
  OR2_X1 U5294 ( .A1(n7190), .A2(n7189), .ZN(n7404) );
  NAND2_X1 U5295 ( .A1(n9434), .A2(n4860), .ZN(n4859) );
  INV_X1 U5296 ( .A(n9009), .ZN(n4860) );
  NOR2_X1 U5297 ( .A1(n7186), .A2(n7992), .ZN(n9010) );
  AND2_X1 U5298 ( .A1(n7903), .A2(n7902), .ZN(n7992) );
  OR2_X1 U5299 ( .A1(n7123), .A2(n8929), .ZN(n7009) );
  OR2_X1 U5300 ( .A1(n6861), .A2(n4824), .ZN(n7010) );
  OAI21_X1 U5301 ( .B1(n6734), .B2(n6733), .A(n8038), .ZN(n6995) );
  AND2_X1 U5302 ( .A1(n7131), .A2(n8931), .ZN(n6728) );
  NAND2_X1 U5303 ( .A1(n8038), .A2(n7891), .ZN(n6733) );
  OAI21_X1 U5304 ( .B1(n6635), .B2(n4837), .A(n6707), .ZN(n4836) );
  NAND2_X1 U5305 ( .A1(n6638), .A2(n4281), .ZN(n4835) );
  NAND2_X1 U5306 ( .A1(n6700), .A2(n7889), .ZN(n6734) );
  NAND2_X1 U5307 ( .A1(n6770), .A2(n6772), .ZN(n4822) );
  NAND2_X1 U5308 ( .A1(n8073), .A2(n6163), .ZN(n4420) );
  NAND2_X1 U5309 ( .A1(n6628), .A2(n6627), .ZN(n7023) );
  NAND2_X1 U5310 ( .A1(n4274), .A2(n6156), .ZN(n6215) );
  INV_X1 U5311 ( .A(n7979), .ZN(n6242) );
  AND2_X1 U5312 ( .A1(n9301), .A2(n9679), .ZN(n4818) );
  XNOR2_X1 U5313 ( .A(n5587), .B(SI_30_), .ZN(n7845) );
  XNOR2_X1 U5314 ( .A(n5416), .B(n5415), .ZN(n7752) );
  INV_X1 U5315 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U5316 ( .A1(n4691), .A2(n4963), .ZN(n5013) );
  NAND2_X1 U5317 ( .A1(n4684), .A2(n4687), .ZN(n4691) );
  NAND2_X1 U5318 ( .A1(n5303), .A2(n4959), .ZN(n4684) );
  OAI21_X1 U5319 ( .B1(n4940), .B2(n4699), .A(n4696), .ZN(n5287) );
  NAND2_X1 U5320 ( .A1(n4470), .A2(n4472), .ZN(n5233) );
  NAND2_X1 U5321 ( .A1(n4476), .A2(n4923), .ZN(n5210) );
  NAND2_X1 U5322 ( .A1(n4904), .A2(n4477), .ZN(n4476) );
  XNOR2_X1 U5323 ( .A(n5191), .B(n5176), .ZN(n6644) );
  AOI21_X2 U5324 ( .B1(n5073), .B2(n4889), .A(n4300), .ZN(n5110) );
  INV_X1 U5325 ( .A(n8574), .ZN(n8688) );
  AOI21_X1 U5326 ( .B1(n4723), .B2(n4725), .A(n4348), .ZN(n4720) );
  NAND2_X1 U5327 ( .A1(n4992), .A2(n4991), .ZN(n8681) );
  INV_X1 U5328 ( .A(n7146), .ZN(n8286) );
  NOR2_X1 U5329 ( .A1(n4865), .A2(n5069), .ZN(n5071) );
  NAND2_X1 U5330 ( .A1(n5570), .A2(n5569), .ZN(n8400) );
  NAND2_X1 U5331 ( .A1(n5092), .A2(n4310), .ZN(n5093) );
  OR2_X1 U5332 ( .A1(n9767), .A2(n5870), .ZN(n9755) );
  NAND2_X1 U5333 ( .A1(n5598), .A2(n5597), .ZN(n8386) );
  NAND2_X1 U5334 ( .A1(n8403), .A2(n8397), .ZN(n5896) );
  INV_X1 U5335 ( .A(n8928), .ZN(n7369) );
  INV_X1 U5336 ( .A(n9627), .ZN(n6717) );
  NAND2_X1 U5337 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  AOI21_X1 U5338 ( .B1(n6058), .B2(P1_IR_REG_31__SCAN_IN), .A(n4793), .ZN(
        n4792) );
  AOI21_X1 U5339 ( .B1(n8069), .B2(n8994), .A(n8111), .ZN(n4670) );
  INV_X1 U5340 ( .A(n8120), .ZN(n4360) );
  NAND2_X1 U5341 ( .A1(n7552), .A2(n7551), .ZN(n9164) );
  OR2_X1 U5342 ( .A1(n7007), .A2(n7006), .ZN(n9435) );
  OR2_X1 U5343 ( .A1(n7293), .A2(n9975), .ZN(n4515) );
  INV_X1 U5344 ( .A(n4831), .ZN(n4830) );
  AOI21_X1 U5345 ( .B1(n4831), .B2(n4829), .A(n4322), .ZN(n4828) );
  NAND2_X1 U5346 ( .A1(n9036), .A2(n4314), .ZN(n4827) );
  NAND2_X1 U5347 ( .A1(n4814), .A2(n9072), .ZN(n9299) );
  NAND2_X1 U5348 ( .A1(n4815), .A2(n9451), .ZN(n4814) );
  NAND2_X1 U5349 ( .A1(n4527), .A2(n9062), .ZN(n9110) );
  INV_X1 U5350 ( .A(n6103), .ZN(n8062) );
  INV_X1 U5351 ( .A(n6751), .ZN(n4564) );
  NAND2_X1 U5352 ( .A1(n6751), .A2(n5721), .ZN(n4566) );
  NAND2_X1 U5353 ( .A1(n4561), .A2(n4560), .ZN(n4568) );
  AOI21_X1 U5354 ( .B1(n4302), .B2(n5628), .A(n5721), .ZN(n4560) );
  AND2_X1 U5355 ( .A1(n7072), .A2(n5632), .ZN(n4567) );
  AND2_X1 U5356 ( .A1(n7918), .A2(n4439), .ZN(n4436) );
  AND2_X1 U5357 ( .A1(n7918), .A2(n4438), .ZN(n4437) );
  NAND2_X1 U5358 ( .A1(n4386), .A2(n4389), .ZN(n5678) );
  NAND2_X1 U5359 ( .A1(n4390), .A2(n5685), .ZN(n4389) );
  NAND2_X1 U5360 ( .A1(n4393), .A2(n5679), .ZN(n4390) );
  NAND2_X1 U5361 ( .A1(n4417), .A2(n4416), .ZN(n4415) );
  NAND2_X1 U5362 ( .A1(n5704), .A2(n5721), .ZN(n4416) );
  INV_X1 U5363 ( .A(n8421), .ZN(n4417) );
  NAND2_X1 U5364 ( .A1(n5696), .A2(n5741), .ZN(n4577) );
  AND2_X1 U5365 ( .A1(n5698), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5366 ( .A1(n4576), .A2(n5719), .ZN(n4575) );
  INV_X1 U5367 ( .A(n5699), .ZN(n4576) );
  OR2_X1 U5368 ( .A1(n4408), .A2(n4414), .ZN(n4407) );
  NAND2_X1 U5369 ( .A1(n4409), .A2(n7526), .ZN(n4408) );
  NAND2_X1 U5370 ( .A1(n4414), .A2(n4415), .ZN(n4409) );
  INV_X1 U5371 ( .A(n5703), .ZN(n4401) );
  AOI21_X1 U5372 ( .B1(n4403), .B2(n4400), .A(n4316), .ZN(n4399) );
  AND2_X1 U5373 ( .A1(n4410), .A2(n4303), .ZN(n4400) );
  NAND2_X1 U5374 ( .A1(n4403), .A2(n4303), .ZN(n4402) );
  OR2_X1 U5375 ( .A1(n5224), .A2(n7230), .ZN(n5226) );
  NAND2_X1 U5376 ( .A1(n8849), .A2(n7607), .ZN(n4747) );
  AOI21_X1 U5377 ( .B1(n4428), .B2(n4430), .A(n4448), .ZN(n4427) );
  OAI21_X1 U5378 ( .B1(n9097), .B2(n4535), .A(n9065), .ZN(n4534) );
  AND2_X1 U5379 ( .A1(n9096), .A2(n4280), .ZN(n4526) );
  AND2_X1 U5380 ( .A1(n7875), .A2(n7888), .ZN(n8018) );
  NOR2_X1 U5381 ( .A1(n7063), .A2(n4500), .ZN(n4499) );
  OR2_X1 U5382 ( .A1(n4503), .A2(n7123), .ZN(n4500) );
  INV_X1 U5383 ( .A(n5286), .ZN(n4695) );
  NOR2_X1 U5384 ( .A1(n5275), .A2(n4701), .ZN(n4700) );
  INV_X1 U5385 ( .A(n4943), .ZN(n4701) );
  NAND2_X1 U5386 ( .A1(n4946), .A2(n4945), .ZN(n4949) );
  NAND2_X1 U5387 ( .A1(n4912), .A2(n4911), .ZN(n4921) );
  INV_X1 U5388 ( .A(n5125), .ZN(n4898) );
  INV_X1 U5389 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9983) );
  INV_X1 U5390 ( .A(n8245), .ZN(n4719) );
  AND2_X1 U5391 ( .A1(n7430), .A2(n4335), .ZN(n4729) );
  INV_X1 U5392 ( .A(n4622), .ZN(n4621) );
  OR2_X1 U5393 ( .A1(n7532), .A2(n7526), .ZN(n5709) );
  OR2_X1 U5394 ( .A1(n5375), .A2(n8155), .ZN(n5388) );
  OR2_X1 U5395 ( .A1(n5359), .A2(n8230), .ZN(n5375) );
  NAND2_X1 U5396 ( .A1(n5002), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5021) );
  INV_X1 U5397 ( .A(n4613), .ZN(n4612) );
  OAI21_X1 U5398 ( .B1(n5663), .B2(n4614), .A(n5605), .ZN(n4613) );
  INV_X1 U5399 ( .A(n5497), .ZN(n4614) );
  INV_X1 U5400 ( .A(n4645), .ZN(n4642) );
  NAND2_X1 U5401 ( .A1(n4645), .A2(n7209), .ZN(n4644) );
  NAND2_X1 U5402 ( .A1(n8771), .A2(n4601), .ZN(n4600) );
  AND2_X1 U5403 ( .A1(n4635), .A2(n4634), .ZN(n5108) );
  OR2_X1 U5404 ( .A1(n5581), .A2(n5082), .ZN(n5083) );
  AND2_X1 U5405 ( .A1(n8605), .A2(n4288), .ZN(n8527) );
  NAND2_X1 U5406 ( .A1(n8605), .A2(n8754), .ZN(n8587) );
  AND2_X1 U5407 ( .A1(n4982), .A2(n4984), .ZN(n4745) );
  NOR2_X1 U5408 ( .A1(n4290), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4381) );
  INV_X1 U5409 ( .A(n6164), .ZN(n6488) );
  INV_X1 U5410 ( .A(n4780), .ZN(n4779) );
  OAI22_X1 U5411 ( .A1(n4296), .A2(n4782), .B1(n4781), .B2(n7554), .ZN(n4780)
         );
  NAND2_X1 U5412 ( .A1(n4427), .A2(n4429), .ZN(n4422) );
  INV_X1 U5413 ( .A(n4430), .ZN(n4429) );
  INV_X1 U5414 ( .A(n8064), .ZN(n4426) );
  INV_X1 U5415 ( .A(n8104), .ZN(n4434) );
  OR2_X1 U5416 ( .A1(n7967), .A2(n9070), .ZN(n8107) );
  NOR2_X1 U5417 ( .A1(n7027), .A2(n4522), .ZN(n7290) );
  AND2_X1 U5418 ( .A1(n7391), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U5419 ( .A1(n9306), .A2(n4497), .ZN(n4496) );
  INV_X1 U5420 ( .A(n4498), .ZN(n4497) );
  INV_X1 U5421 ( .A(n9124), .ZN(n4841) );
  OR2_X1 U5422 ( .A1(n9354), .A2(n9254), .ZN(n7996) );
  INV_X1 U5423 ( .A(n7992), .ZN(n4856) );
  INV_X1 U5424 ( .A(n4859), .ZN(n4858) );
  OR2_X1 U5425 ( .A1(n9472), .A2(n7281), .ZN(n7903) );
  NOR2_X1 U5426 ( .A1(n6995), .A2(n8037), .ZN(n9042) );
  INV_X1 U5427 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6663) );
  OR2_X1 U5428 ( .A1(n6664), .A2(n6663), .ZN(n6736) );
  AND2_X1 U5429 ( .A1(n6733), .A2(n4281), .ZN(n4455) );
  NAND2_X1 U5430 ( .A1(n6380), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6651) );
  NOR2_X1 U5431 ( .A1(n4469), .A2(n6629), .ZN(n6775) );
  INV_X1 U5432 ( .A(n6213), .ZN(n6160) );
  INV_X1 U5433 ( .A(n6658), .ZN(n6152) );
  AND2_X1 U5434 ( .A1(n7197), .A2(n7374), .ZN(n9443) );
  INV_X1 U5435 ( .A(n4678), .ZN(n4677) );
  AOI21_X1 U5436 ( .B1(n4676), .B2(n4678), .A(n4353), .ZN(n4675) );
  NOR2_X1 U5437 ( .A1(n5574), .A2(n4679), .ZN(n4678) );
  INV_X1 U5438 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6089) );
  AOI21_X1 U5439 ( .B1(n4685), .B2(n4688), .A(n4682), .ZN(n4681) );
  INV_X1 U5440 ( .A(n4968), .ZN(n4682) );
  AND2_X1 U5441 ( .A1(n5336), .A2(n4972), .ZN(n5334) );
  INV_X1 U5442 ( .A(n4700), .ZN(n4699) );
  NOR2_X1 U5443 ( .A1(n4944), .A2(n4703), .ZN(n4702) );
  INV_X1 U5444 ( .A(n4939), .ZN(n4703) );
  AOI21_X1 U5445 ( .B1(n4473), .B2(n4474), .A(n4326), .ZN(n4472) );
  NOR2_X1 U5446 ( .A1(n4915), .A2(n4478), .ZN(n4477) );
  INV_X1 U5447 ( .A(n4903), .ZN(n4478) );
  OR2_X1 U5448 ( .A1(n5190), .A2(n4920), .ZN(n4915) );
  OR2_X1 U5449 ( .A1(n4919), .A2(n4918), .ZN(n5192) );
  OR2_X1 U5450 ( .A1(n5176), .A2(n4919), .ZN(n5190) );
  NAND2_X1 U5451 ( .A1(n5907), .A2(n4791), .ZN(n4790) );
  INV_X1 U5452 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4791) );
  INV_X1 U5453 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4819) );
  INV_X1 U5454 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4418) );
  AOI21_X1 U5455 ( .B1(n4726), .B2(n7522), .A(n4724), .ZN(n4723) );
  INV_X1 U5456 ( .A(n7524), .ZN(n4724) );
  INV_X1 U5457 ( .A(n4726), .ZN(n4725) );
  OR2_X1 U5458 ( .A1(n5021), .A2(n8223), .ZN(n5341) );
  NAND2_X1 U5459 ( .A1(n5340), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5359) );
  INV_X1 U5460 ( .A(n5341), .ZN(n5340) );
  NAND2_X1 U5461 ( .A1(n4709), .A2(n4707), .ZN(n5855) );
  NAND2_X1 U5462 ( .A1(n4994), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5137) );
  INV_X1 U5463 ( .A(n9741), .ZN(n6837) );
  AND2_X1 U5464 ( .A1(n8126), .A2(n4868), .ZN(n5779) );
  AND2_X1 U5465 ( .A1(n9777), .A2(n5757), .ZN(n4569) );
  NAND2_X1 U5466 ( .A1(n6857), .A2(n8433), .ZN(n5878) );
  AND4_X1 U5467 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n8249)
         );
  AND4_X1 U5468 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n7446)
         );
  AND4_X1 U5469 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n7304)
         );
  NAND2_X1 U5470 ( .A1(n5054), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U5471 ( .A1(n6945), .A2(n6946), .ZN(n7093) );
  NAND2_X1 U5472 ( .A1(n7093), .A2(n4373), .ZN(n7099) );
  OR2_X1 U5473 ( .A1(n7094), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5474 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  AOI21_X1 U5475 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8352), .A(n8351), .ZN(
        n8354) );
  NOR2_X1 U5476 ( .A1(n8423), .A2(n7532), .ZN(n5895) );
  INV_X1 U5477 ( .A(n8434), .ZN(n4626) );
  NOR2_X1 U5478 ( .A1(n8421), .A2(n4623), .ZN(n4622) );
  INV_X1 U5479 ( .A(n5702), .ZN(n4623) );
  OR2_X1 U5480 ( .A1(n8425), .A2(n5510), .ZN(n5449) );
  INV_X1 U5481 ( .A(n5406), .ZN(n5405) );
  OR2_X1 U5482 ( .A1(n8456), .A2(n8275), .ZN(n5413) );
  NAND2_X1 U5483 ( .A1(n5699), .A2(n5700), .ZN(n8452) );
  NAND2_X1 U5484 ( .A1(n8665), .A2(n8505), .ZN(n5379) );
  NAND2_X1 U5485 ( .A1(n8527), .A2(n8747), .ZN(n8508) );
  NAND2_X1 U5486 ( .A1(n5690), .A2(n5691), .ZN(n8487) );
  NAND2_X1 U5487 ( .A1(n8605), .A2(n4593), .ZN(n8568) );
  AND4_X1 U5488 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n8567)
         );
  OR2_X1 U5489 ( .A1(n8610), .A2(n8620), .ZN(n8577) );
  OR2_X1 U5490 ( .A1(n5324), .A2(n8250), .ZN(n5326) );
  AND4_X1 U5491 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n8595)
         );
  AND2_X1 U5492 ( .A1(n8627), .A2(n8758), .ZN(n8605) );
  NAND2_X1 U5493 ( .A1(n5000), .A2(n4999), .ZN(n5309) );
  INV_X1 U5494 ( .A(n5295), .ZN(n5000) );
  NAND2_X1 U5495 ( .A1(n7445), .A2(n5497), .ZN(n8618) );
  NAND2_X1 U5496 ( .A1(n5496), .A2(n5663), .ZN(n7445) );
  INV_X1 U5497 ( .A(n4601), .ZN(n4599) );
  NAND2_X1 U5498 ( .A1(n7204), .A2(n5652), .ZN(n7313) );
  NAND2_X1 U5499 ( .A1(n4998), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5254) );
  INV_X1 U5500 ( .A(n5240), .ZN(n4998) );
  OR2_X1 U5501 ( .A1(n5254), .A2(n6947), .ZN(n5267) );
  AND2_X1 U5502 ( .A1(n7152), .A2(n9825), .ZN(n7338) );
  AND4_X1 U5503 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n7331)
         );
  OR2_X1 U5504 ( .A1(n5153), .A2(n5152), .ZN(n5170) );
  NAND2_X1 U5505 ( .A1(n4996), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5217) );
  INV_X1 U5506 ( .A(n5170), .ZN(n4996) );
  AND4_X1 U5507 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n7162)
         );
  NOR2_X1 U5508 ( .A1(n7081), .A2(n7233), .ZN(n7152) );
  OR2_X1 U5509 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  OAI211_X1 U5510 ( .C1(n6354), .C2(n6474), .A(n5149), .B(n5148), .ZN(n6765)
         );
  OR2_X1 U5511 ( .A1(n6831), .A2(n6765), .ZN(n7081) );
  AND2_X1 U5512 ( .A1(n5630), .A2(n5631), .ZN(n6754) );
  INV_X1 U5513 ( .A(n9742), .ZN(n8621) );
  AND2_X1 U5514 ( .A1(n6919), .A2(n8131), .ZN(n6920) );
  NAND2_X1 U5515 ( .A1(n4993), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5116) );
  INV_X1 U5516 ( .A(n5097), .ZN(n4993) );
  OR2_X1 U5517 ( .A1(n5077), .A2(n5989), .ZN(n5081) );
  OR2_X1 U5518 ( .A1(n6851), .A2(n5093), .ZN(n9752) );
  INV_X1 U5519 ( .A(n6214), .ZN(n4667) );
  NAND2_X1 U5520 ( .A1(n5481), .A2(n6595), .ZN(n6971) );
  NAND2_X1 U5521 ( .A1(n5439), .A2(n5438), .ZN(n8424) );
  NAND2_X1 U5522 ( .A1(n7789), .A2(n5576), .ZN(n5439) );
  AND3_X1 U5523 ( .A1(n4287), .A2(n8432), .A3(n8603), .ZN(n8650) );
  NAND2_X1 U5524 ( .A1(n5280), .A2(n5279), .ZN(n7448) );
  NAND2_X1 U5525 ( .A1(n4647), .A2(n4648), .ZN(n7319) );
  OR2_X1 U5526 ( .A1(n5077), .A2(n5988), .ZN(n5065) );
  NOR2_X1 U5527 ( .A1(n5041), .A2(n6595), .ZN(n9781) );
  AND2_X1 U5528 ( .A1(n7310), .A2(n5542), .ZN(n9768) );
  NAND2_X1 U5529 ( .A1(n6351), .A2(n9774), .ZN(n9767) );
  NAND3_X1 U5530 ( .A1(n4736), .A2(n4975), .A3(n4589), .ZN(n5004) );
  NOR2_X1 U5531 ( .A1(n4742), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U5532 ( .A1(n5531), .A2(n4591), .ZN(n4590) );
  INV_X1 U5533 ( .A(n4745), .ZN(n4742) );
  AND2_X1 U5534 ( .A1(n4736), .A2(n4975), .ZN(n5530) );
  INV_X1 U5535 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5531) );
  AND2_X1 U5536 ( .A1(n4738), .A2(n4383), .ZN(n4384) );
  NOR2_X1 U5537 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4383) );
  INV_X1 U5538 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4974) );
  INV_X1 U5539 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U5540 ( .A1(n6156), .A2(n4878), .ZN(n5049) );
  NAND2_X1 U5541 ( .A1(n8818), .A2(n7668), .ZN(n4768) );
  NAND2_X1 U5542 ( .A1(n4268), .A2(n6492), .ZN(n4774) );
  NAND2_X1 U5543 ( .A1(n4770), .A2(n4772), .ZN(n4775) );
  INV_X1 U5544 ( .A(n6493), .ZN(n4770) );
  NAND2_X1 U5545 ( .A1(n4748), .A2(n7604), .ZN(n8847) );
  INV_X1 U5546 ( .A(n4263), .ZN(n4748) );
  NAND2_X1 U5547 ( .A1(n6131), .A2(n6130), .ZN(n6151) );
  NAND2_X1 U5548 ( .A1(n6387), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7673) );
  INV_X1 U5549 ( .A(n7653), .ZN(n6387) );
  OR2_X1 U5550 ( .A1(n7673), .A2(n10001), .ZN(n7694) );
  OR2_X1 U5551 ( .A1(n7694), .A2(n7693), .ZN(n7716) );
  NAND2_X1 U5552 ( .A1(n6388), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7735) );
  INV_X1 U5553 ( .A(n7716), .ZN(n6388) );
  NAND2_X1 U5554 ( .A1(n4778), .A2(n4777), .ZN(n7585) );
  AOI21_X1 U5555 ( .B1(n4296), .B2(n7555), .A(n4782), .ZN(n4777) );
  NAND2_X1 U5556 ( .A1(n4794), .A2(n5948), .ZN(n4793) );
  NAND2_X1 U5557 ( .A1(n4795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4794) );
  INV_X1 U5558 ( .A(n4276), .ZN(n7633) );
  INV_X1 U5559 ( .A(n4272), .ZN(n7797) );
  OR2_X1 U5560 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5962) );
  OR2_X1 U5561 ( .A1(n9506), .A2(n9505), .ZN(n4521) );
  AOI21_X1 U5562 ( .B1(n6276), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9537), .ZN(
        n9551) );
  NOR2_X1 U5563 ( .A1(n9552), .A2(n4340), .ZN(n8946) );
  NAND2_X1 U5564 ( .A1(n8946), .A2(n8947), .ZN(n8945) );
  AOI21_X1 U5565 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6645), .A(n6401), .ZN(
        n9565) );
  NOR2_X1 U5566 ( .A1(n9566), .A2(n4517), .ZN(n9581) );
  NOR2_X1 U5567 ( .A1(n4519), .A2(n4518), .ZN(n4517) );
  INV_X1 U5568 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4518) );
  INV_X1 U5569 ( .A(n9572), .ZN(n4519) );
  NOR2_X1 U5570 ( .A1(n9581), .A2(n9580), .ZN(n9579) );
  NAND2_X1 U5571 ( .A1(n9598), .A2(n9599), .ZN(n9597) );
  NAND2_X1 U5572 ( .A1(n9595), .A2(n9596), .ZN(n9594) );
  NOR2_X1 U5573 ( .A1(n6611), .A2(n4351), .ZN(n6615) );
  NOR2_X1 U5574 ( .A1(n6615), .A2(n6614), .ZN(n7027) );
  NAND2_X1 U5575 ( .A1(n6618), .A2(n6619), .ZN(n7032) );
  XNOR2_X1 U5576 ( .A(n7290), .B(n7289), .ZN(n7029) );
  NAND2_X1 U5577 ( .A1(n7032), .A2(n4368), .ZN(n7033) );
  OR2_X1 U5578 ( .A1(n7391), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4368) );
  AOI21_X1 U5579 ( .B1(n8975), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8974), .ZN(
        n8977) );
  NOR2_X1 U5580 ( .A1(n9607), .A2(n9608), .ZN(n9606) );
  INV_X1 U5581 ( .A(n4297), .ZN(n4829) );
  NOR2_X1 U5582 ( .A1(n9039), .A2(n4298), .ZN(n4831) );
  XNOR2_X1 U5583 ( .A(n4816), .B(n9039), .ZN(n4815) );
  AOI21_X1 U5584 ( .B1(n9083), .B2(n9082), .A(n9067), .ZN(n4816) );
  AND2_X1 U5585 ( .A1(n7792), .A2(n7791), .ZN(n9034) );
  NOR2_X1 U5586 ( .A1(n4532), .A2(n9064), .ZN(n9098) );
  INV_X1 U5587 ( .A(n4536), .ZN(n4532) );
  OAI21_X1 U5588 ( .B1(n9143), .B2(n8005), .A(n4280), .ZN(n4536) );
  OR2_X1 U5589 ( .A1(n7775), .A2(n8903), .ZN(n7811) );
  NOR2_X1 U5590 ( .A1(n9063), .A2(n4531), .ZN(n4530) );
  INV_X1 U5591 ( .A(n9061), .ZN(n4531) );
  NAND2_X1 U5592 ( .A1(n9153), .A2(n9142), .ZN(n9137) );
  NAND2_X1 U5593 ( .A1(n9190), .A2(n9181), .ZN(n9174) );
  NOR2_X1 U5594 ( .A1(n9174), .A2(n9328), .ZN(n9153) );
  INV_X1 U5595 ( .A(n4799), .ZN(n4798) );
  OAI22_X1 U5596 ( .A1(n4804), .A2(n4800), .B1(n9049), .B2(n9050), .ZN(n4799)
         );
  NAND2_X1 U5597 ( .A1(n9245), .A2(n9232), .ZN(n9229) );
  NAND2_X1 U5598 ( .A1(n7996), .A2(n9051), .ZN(n9238) );
  OAI21_X1 U5599 ( .B1(n9244), .B2(n9016), .A(n4347), .ZN(n9228) );
  INV_X1 U5600 ( .A(n7594), .ZN(n6385) );
  OR2_X1 U5601 ( .A1(n7611), .A2(n8857), .ZN(n7631) );
  NOR2_X1 U5602 ( .A1(n9267), .A2(n9359), .ZN(n9245) );
  NAND2_X1 U5603 ( .A1(n9278), .A2(n9272), .ZN(n9267) );
  NOR2_X1 U5604 ( .A1(n9457), .A2(n9045), .ZN(n9283) );
  NAND2_X1 U5605 ( .A1(n7560), .A2(n7559), .ZN(n10034) );
  NAND2_X1 U5606 ( .A1(n6383), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7190) );
  INV_X1 U5607 ( .A(n7001), .ZN(n6383) );
  NAND2_X1 U5608 ( .A1(n4550), .A2(n9040), .ZN(n9433) );
  NAND2_X1 U5609 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5610 ( .A(n9041), .ZN(n4551) );
  INV_X1 U5611 ( .A(n9042), .ZN(n4552) );
  INV_X1 U5612 ( .A(n4549), .ZN(n9450) );
  OR2_X1 U5613 ( .A1(n6736), .A2(n7117), .ZN(n6870) );
  NAND2_X1 U5614 ( .A1(n4502), .A2(n4501), .ZN(n6877) );
  NOR2_X1 U5615 ( .A1(n7063), .A2(n4503), .ZN(n4501) );
  NOR2_X1 U5616 ( .A1(n6887), .A2(n4503), .ZN(n6744) );
  NAND2_X1 U5617 ( .A1(n4545), .A2(n4543), .ZN(n6700) );
  INV_X1 U5618 ( .A(n8084), .ZN(n4544) );
  NOR2_X1 U5619 ( .A1(n6887), .A2(n6803), .ZN(n6702) );
  AND2_X1 U5620 ( .A1(n7888), .A2(n7877), .ZN(n7874) );
  AND2_X1 U5621 ( .A1(n6777), .A2(n6775), .ZN(n6776) );
  NAND2_X1 U5622 ( .A1(n8081), .A2(n8031), .ZN(n9626) );
  NAND2_X1 U5623 ( .A1(n6789), .A2(n8071), .ZN(n7019) );
  AND2_X1 U5624 ( .A1(n8937), .A2(n6290), .ZN(n6243) );
  INV_X1 U5625 ( .A(n9307), .ZN(n4466) );
  NOR2_X1 U5626 ( .A1(n9309), .A2(n4488), .ZN(n4487) );
  AND2_X1 U5627 ( .A1(n9310), .A2(n9679), .ZN(n4488) );
  NAND2_X1 U5628 ( .A1(n7771), .A2(n6643), .ZN(n7774) );
  NAND2_X1 U5629 ( .A1(n6541), .A2(n6643), .ZN(n4805) );
  OR2_X1 U5630 ( .A1(n6286), .A2(n8110), .ZN(n9701) );
  INV_X1 U5631 ( .A(n9701), .ZN(n9679) );
  XNOR2_X1 U5632 ( .A(n5575), .B(n5568), .ZN(n7955) );
  NAND2_X1 U5633 ( .A1(n4680), .A2(n5566), .ZN(n5575) );
  NAND2_X1 U5634 ( .A1(n5562), .A2(n5561), .ZN(n4680) );
  XNOR2_X1 U5635 ( .A(n5452), .B(n5451), .ZN(n7789) );
  OAI21_X1 U5636 ( .B1(n5366), .B2(n5365), .A(n5364), .ZN(n5381) );
  AND2_X1 U5637 ( .A1(n5382), .A2(n5372), .ZN(n5380) );
  OAI21_X1 U5638 ( .B1(n5303), .B2(n4960), .A(n4959), .ZN(n5317) );
  XNOR2_X1 U5639 ( .A(n4480), .B(n5275), .ZN(n7567) );
  NAND2_X1 U5640 ( .A1(n4481), .A2(n4943), .ZN(n4480) );
  NAND2_X1 U5641 ( .A1(n4940), .A2(n4702), .ZN(n4481) );
  OR2_X1 U5642 ( .A1(n6052), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6118) );
  AND2_X1 U5643 ( .A1(n6023), .A2(n6029), .ZN(n6863) );
  XNOR2_X1 U5644 ( .A(n5182), .B(n5181), .ZN(n6730) );
  XNOR2_X1 U5645 ( .A(n5147), .B(n5146), .ZN(n6639) );
  XNOR2_X1 U5646 ( .A(n4891), .B(SI_4_), .ZN(n5074) );
  NAND2_X1 U5647 ( .A1(n4885), .A2(n4884), .ZN(n5088) );
  XNOR2_X1 U5648 ( .A(n4886), .B(SI_3_), .ZN(n5087) );
  XNOR2_X1 U5649 ( .A(n5960), .B(P1_IR_REG_1__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U5650 ( .A1(n6586), .A2(n5789), .ZN(n5942) );
  NAND2_X1 U5651 ( .A1(n4722), .A2(n4726), .ZN(n8142) );
  NAND2_X1 U5652 ( .A1(n5861), .A2(n7516), .ZN(n4722) );
  AOI21_X1 U5653 ( .B1(n5820), .B2(n4731), .A(n4730), .ZN(n4728) );
  NAND2_X1 U5654 ( .A1(n5266), .A2(n5265), .ZN(n7493) );
  AND2_X1 U5655 ( .A1(n4717), .A2(n4716), .ZN(n8165) );
  AND4_X1 U5656 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n7332)
         );
  NAND2_X1 U5657 ( .A1(n5239), .A2(n5238), .ZN(n7210) );
  NAND2_X1 U5658 ( .A1(n5293), .A2(n5292), .ZN(n8629) );
  NAND2_X1 U5659 ( .A1(n8206), .A2(n8205), .ZN(n8246) );
  NAND2_X1 U5660 ( .A1(n5385), .A2(n5384), .ZN(n8473) );
  CLKBUF_X1 U5661 ( .A(n5932), .Z(n6529) );
  INV_X1 U5662 ( .A(n5481), .ZN(n6570) );
  NAND2_X1 U5663 ( .A1(n4713), .A2(n4715), .ZN(n4712) );
  NAND2_X1 U5664 ( .A1(n4716), .A2(n8164), .ZN(n4713) );
  NAND2_X1 U5665 ( .A1(n5820), .A2(n5819), .ZN(n7303) );
  NAND2_X1 U5666 ( .A1(n5358), .A2(n5357), .ZN(n8511) );
  NAND2_X1 U5667 ( .A1(n5869), .A2(n9755), .ZN(n8238) );
  INV_X1 U5668 ( .A(n8199), .ZN(n8233) );
  CLKBUF_X1 U5669 ( .A(n6579), .Z(n8137) );
  INV_X1 U5670 ( .A(n8238), .ZN(n8270) );
  AND2_X1 U5671 ( .A1(n5877), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8266) );
  NAND2_X1 U5672 ( .A1(n5725), .A2(n4569), .ZN(n5750) );
  AND2_X1 U5673 ( .A1(n5515), .A2(n5514), .ZN(n6378) );
  NOR2_X1 U5674 ( .A1(n7466), .A2(n7465), .ZN(n7468) );
  INV_X1 U5675 ( .A(n9418), .ZN(n9724) );
  NAND2_X1 U5676 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  NAND2_X1 U5677 ( .A1(n5422), .A2(n5421), .ZN(n8443) );
  NAND2_X1 U5678 ( .A1(n8490), .A2(n5691), .ZN(n8466) );
  OAI21_X1 U5679 ( .B1(n8543), .B2(n4655), .A(n4654), .ZN(n8499) );
  NOR2_X1 U5680 ( .A1(n8685), .A2(n4658), .ZN(n8518) );
  AND2_X1 U5681 ( .A1(n5018), .A2(n5017), .ZN(n8574) );
  NAND2_X1 U5682 ( .A1(n4660), .A2(n4662), .ZN(n8556) );
  OR2_X1 U5683 ( .A1(n8600), .A2(n4664), .ZN(n4660) );
  AND2_X1 U5684 ( .A1(n4665), .A2(n4282), .ZN(n8582) );
  NAND2_X1 U5685 ( .A1(n7315), .A2(n5658), .ZN(n7489) );
  NAND2_X1 U5686 ( .A1(n5252), .A2(n5251), .ZN(n7503) );
  NAND2_X1 U5687 ( .A1(n5214), .A2(n5213), .ZN(n7226) );
  NAND2_X1 U5688 ( .A1(n7075), .A2(n5168), .ZN(n7143) );
  NAND2_X1 U5689 ( .A1(n5291), .A2(n9410), .ZN(n4607) );
  NAND2_X1 U5690 ( .A1(n5076), .A2(n5036), .ZN(n4608) );
  INV_X1 U5691 ( .A(n8609), .ZN(n9762) );
  AND2_X1 U5692 ( .A1(n9757), .A2(n6591), .ZN(n9764) );
  AND2_X1 U5693 ( .A1(n9757), .A2(n6593), .ZN(n8609) );
  AND2_X1 U5694 ( .A1(n5578), .A2(n5577), .ZN(n8726) );
  AND2_X1 U5695 ( .A1(n8642), .A2(n8641), .ZN(n8723) );
  AOI211_X1 U5696 ( .C1(n8405), .C2(n9838), .A(n8411), .B(n8404), .ZN(n5555)
         );
  INV_X1 U5697 ( .A(n8424), .ZN(n8730) );
  INV_X1 U5698 ( .A(n9769), .ZN(n9772) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9928) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9959) );
  OR3_X1 U5701 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5702 ( .A1(n7107), .A2(n7106), .ZN(n4766) );
  XNOR2_X1 U5703 ( .A(n6297), .B(n6295), .ZN(n6293) );
  NAND2_X1 U5704 ( .A1(n7651), .A2(n7650), .ZN(n9349) );
  NAND2_X1 U5705 ( .A1(n7592), .A2(n7591), .ZN(n9365) );
  NAND2_X1 U5706 ( .A1(n8847), .A2(n7607), .ZN(n8856) );
  AND2_X1 U5707 ( .A1(n7757), .A2(n7546), .ZN(n9140) );
  NAND2_X1 U5708 ( .A1(n8815), .A2(n7668), .ZN(n8872) );
  NAND2_X1 U5709 ( .A1(n7714), .A2(n7713), .ZN(n9334) );
  AOI21_X1 U5710 ( .B1(n4764), .B2(n4763), .A(n4323), .ZN(n4762) );
  INV_X1 U5711 ( .A(n8904), .ZN(n8918) );
  AND2_X1 U5712 ( .A1(n6195), .A2(n9512), .ZN(n8901) );
  NAND2_X1 U5713 ( .A1(n4772), .A2(n6494), .ZN(n4771) );
  INV_X1 U5714 ( .A(n6494), .ZN(n4773) );
  NAND2_X1 U5715 ( .A1(n8864), .A2(n4758), .ZN(n4752) );
  NAND2_X1 U5716 ( .A1(n4756), .A2(n4754), .ZN(n4753) );
  NAND2_X1 U5717 ( .A1(n7764), .A2(n7763), .ZN(n9147) );
  OR2_X1 U5718 ( .A1(n7579), .A2(n7578), .ZN(n9453) );
  OR2_X1 U5719 ( .A1(n7193), .A2(n7192), .ZN(n9454) );
  OR2_X1 U5720 ( .A1(n6873), .A2(n6872), .ZN(n8928) );
  OR2_X1 U5721 ( .A1(n6654), .A2(n6653), .ZN(n8931) );
  OR2_X1 U5722 ( .A1(n6500), .A2(n6499), .ZN(n8933) );
  OR2_X1 U5723 ( .A1(n6319), .A2(n6318), .ZN(n8934) );
  OAI22_X1 U5724 ( .A1(n6230), .A2(n6106), .B1(n4277), .B2(n6260), .ZN(n6107)
         );
  AND2_X1 U5725 ( .A1(n4521), .A2(n4520), .ZN(n5969) );
  NAND2_X1 U5726 ( .A1(n9515), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4520) );
  AOI21_X1 U5727 ( .B1(n9515), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9500), .ZN(
        n5977) );
  AND2_X1 U5728 ( .A1(n4820), .A2(n4821), .ZN(n5991) );
  NOR2_X1 U5729 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4820) );
  NAND2_X1 U5730 ( .A1(n6269), .A2(n6268), .ZN(n6409) );
  NAND2_X1 U5731 ( .A1(n8945), .A2(n4510), .ZN(n6269) );
  NAND2_X1 U5732 ( .A1(n8938), .A2(n4511), .ZN(n4510) );
  INV_X1 U5733 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U5734 ( .A1(n9594), .A2(n4367), .ZN(n6404) );
  NAND2_X1 U5735 ( .A1(n6400), .A2(n9482), .ZN(n4367) );
  NOR2_X1 U5736 ( .A1(n8960), .A2(n8959), .ZN(n8962) );
  OAI21_X1 U5737 ( .B1(n7293), .B2(n4513), .A(n4512), .ZN(n8969) );
  NAND2_X1 U5738 ( .A1(n4516), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5739 ( .A1(n8954), .A2(n4516), .ZN(n4512) );
  INV_X1 U5740 ( .A(n8956), .ZN(n4516) );
  INV_X1 U5741 ( .A(n8954), .ZN(n4514) );
  XNOR2_X1 U5742 ( .A(n4369), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U5743 ( .A1(n9616), .A2(n4370), .ZN(n4369) );
  OR2_X1 U5744 ( .A1(n8988), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4370) );
  XNOR2_X1 U5745 ( .A(n4507), .B(n4506), .ZN(n8993) );
  INV_X1 U5746 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4506) );
  OR2_X1 U5747 ( .A1(n9606), .A2(n4508), .ZN(n4507) );
  AND2_X1 U5748 ( .A1(n8988), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4508) );
  INV_X1 U5749 ( .A(n7963), .ZN(n9294) );
  INV_X1 U5750 ( .A(n7967), .ZN(n9297) );
  AOI21_X1 U5751 ( .B1(n9630), .B2(n8926), .A(n4541), .ZN(n4540) );
  OR2_X1 U5752 ( .A1(n9084), .A2(n9632), .ZN(n4542) );
  NOR2_X1 U5753 ( .A1(n9085), .A2(n9289), .ZN(n4541) );
  NAND2_X1 U5754 ( .A1(n4492), .A2(n4490), .ZN(n9308) );
  INV_X1 U5755 ( .A(n4491), .ZN(n4490) );
  OR2_X1 U5756 ( .A1(n9099), .A2(n9632), .ZN(n4492) );
  OAI22_X1 U5757 ( .A1(n9128), .A2(n9287), .B1(n9100), .B2(n9289), .ZN(n4491)
         );
  NAND2_X1 U5758 ( .A1(n7752), .A2(n6643), .ZN(n7755) );
  NAND2_X1 U5759 ( .A1(n9143), .A2(n9061), .ZN(n9125) );
  NAND2_X1 U5760 ( .A1(n4839), .A2(n4842), .ZN(n9123) );
  OR2_X1 U5761 ( .A1(n9025), .A2(n4845), .ZN(n4839) );
  NAND2_X1 U5762 ( .A1(n4847), .A2(n9026), .ZN(n9136) );
  NAND2_X1 U5763 ( .A1(n4537), .A2(n4807), .ZN(n9160) );
  NAND2_X1 U5764 ( .A1(n9025), .A2(n9024), .ZN(n9152) );
  INV_X1 U5765 ( .A(n9334), .ZN(n9181) );
  NOR2_X1 U5766 ( .A1(n9185), .A2(n9056), .ZN(n9171) );
  NAND2_X1 U5767 ( .A1(n7692), .A2(n7691), .ZN(n9339) );
  NAND2_X1 U5768 ( .A1(n4853), .A2(n4283), .ZN(n9184) );
  OR2_X1 U5769 ( .A1(n9198), .A2(n9021), .ZN(n4853) );
  OAI21_X1 U5770 ( .B1(n9457), .B2(n4797), .A(n4796), .ZN(n9251) );
  AOI21_X1 U5771 ( .B1(n4804), .B2(n9046), .A(n4803), .ZN(n4796) );
  OR2_X1 U5772 ( .A1(n9010), .A2(n4859), .ZN(n9431) );
  NOR2_X1 U5773 ( .A1(n9010), .A2(n9009), .ZN(n9432) );
  NAND2_X1 U5774 ( .A1(n7393), .A2(n7392), .ZN(n9442) );
  NAND2_X1 U5775 ( .A1(n6998), .A2(n6997), .ZN(n7286) );
  NAND2_X1 U5776 ( .A1(n7010), .A2(n7009), .ZN(n7184) );
  OR2_X1 U5777 ( .A1(n9648), .A2(n6673), .ZN(n9638) );
  OAI21_X1 U5778 ( .B1(n6636), .B2(n4835), .A(n4832), .ZN(n6656) );
  NAND2_X1 U5779 ( .A1(n4836), .A2(n4281), .ZN(n4832) );
  NAND2_X1 U5780 ( .A1(n6644), .A2(n6643), .ZN(n6647) );
  NAND2_X1 U5781 ( .A1(n6883), .A2(n6638), .ZN(n6708) );
  INV_X1 U5782 ( .A(n6713), .ZN(n6633) );
  INV_X1 U5783 ( .A(n9638), .ZN(n10033) );
  OR2_X1 U5784 ( .A1(n9458), .A2(n6147), .ZN(n9635) );
  AND2_X1 U5785 ( .A1(n4817), .A2(n4813), .ZN(n9302) );
  NOR2_X1 U5786 ( .A1(n9300), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5787 ( .A1(n4465), .A2(n4463), .ZN(n9379) );
  NOR2_X1 U5788 ( .A1(n4464), .A2(n9304), .ZN(n4463) );
  NAND2_X1 U5789 ( .A1(n4466), .A2(n9705), .ZN(n4465) );
  OR2_X1 U5790 ( .A1(n9305), .A2(n4350), .ZN(n4464) );
  NAND2_X1 U5791 ( .A1(n4489), .A2(n4485), .ZN(n9380) );
  INV_X1 U5792 ( .A(n9308), .ZN(n4489) );
  INV_X1 U5793 ( .A(n4486), .ZN(n4485) );
  OAI21_X1 U5794 ( .B1(n9311), .B2(n9373), .A(n4487), .ZN(n4486) );
  INV_X1 U5795 ( .A(n6097), .ZN(n7514) );
  CLKBUF_X1 U5796 ( .A(n5967), .Z(n8123) );
  NAND2_X1 U5797 ( .A1(n5927), .A2(n5929), .ZN(n5924) );
  XNOR2_X1 U5798 ( .A(n5381), .B(n5380), .ZN(n7730) );
  CLKBUF_X1 U5799 ( .A(n6102), .Z(n8111) );
  AND2_X1 U5800 ( .A1(n6523), .A2(n6338), .ZN(n8987) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6024) );
  INV_X1 U5802 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6301) );
  INV_X1 U5803 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5804 ( .A1(n4452), .A2(n4881), .ZN(n5060) );
  NAND2_X1 U5805 ( .A1(n5035), .A2(n5034), .ZN(n4452) );
  INV_X1 U5806 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6181) );
  NOR2_X1 U5807 ( .A1(n7264), .A2(n10053), .ZN(n9884) );
  INV_X1 U5808 ( .A(n5903), .ZN(n5904) );
  OAI21_X1 U5809 ( .B1(n8720), .B2(n5900), .A(n4595), .ZN(P2_U3519) );
  AOI21_X1 U5810 ( .B1(n8386), .B2(n6840), .A(n4596), .ZN(n4595) );
  NOR2_X1 U5811 ( .A1(n9840), .A2(n8721), .ZN(n4596) );
  NOR2_X1 U5812 ( .A1(n4342), .A2(n5898), .ZN(n5899) );
  OR2_X1 U5813 ( .A1(n8119), .A2(n8118), .ZN(n4358) );
  INV_X1 U5814 ( .A(n4515), .ZN(n8953) );
  NAND2_X1 U5815 ( .A1(n4539), .A2(n4538), .ZN(P1_U3551) );
  OR2_X1 U5816 ( .A1(n9721), .A2(n7816), .ZN(n4538) );
  NAND2_X1 U5817 ( .A1(n9379), .A2(n9721), .ZN(n4539) );
  NAND2_X1 U5818 ( .A1(n4462), .A2(n4460), .ZN(P1_U3519) );
  OR2_X1 U5819 ( .A1(n9709), .A2(n4461), .ZN(n4460) );
  NAND2_X1 U5820 ( .A1(n9379), .A2(n9709), .ZN(n4462) );
  INV_X1 U5821 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U5822 ( .A1(n4484), .A2(n4482), .ZN(P1_U3518) );
  OR2_X1 U5823 ( .A1(n9709), .A2(n4483), .ZN(n4482) );
  NAND2_X1 U5824 ( .A1(n9380), .A2(n9709), .ZN(n4484) );
  INV_X1 U5825 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n4483) );
  AND2_X1 U5826 ( .A1(n9109), .A2(n4528), .ZN(n4280) );
  OR2_X1 U5827 ( .A1(n6803), .A2(n8932), .ZN(n4281) );
  OR2_X1 U5828 ( .A1(n8610), .A2(n5315), .ZN(n4282) );
  AND2_X1 U5829 ( .A1(n9187), .A2(n4852), .ZN(n4283) );
  XNOR2_X1 U5830 ( .A(n5950), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6075) );
  AND2_X1 U5831 ( .A1(n4719), .A2(n8205), .ZN(n4284) );
  NAND2_X1 U5832 ( .A1(n4435), .A2(n4433), .ZN(n4285) );
  NAND2_X1 U5833 ( .A1(n4493), .A2(n4808), .ZN(n4537) );
  AND2_X1 U5834 ( .A1(n4593), .A2(n4592), .ZN(n4286) );
  OR2_X1 U5835 ( .A1(n8481), .A2(n4604), .ZN(n4287) );
  AND2_X1 U5836 ( .A1(n4286), .A2(n8532), .ZN(n4288) );
  AND2_X1 U5837 ( .A1(n4644), .A2(n4642), .ZN(n4289) );
  NAND2_X1 U5838 ( .A1(n5472), .A2(n5475), .ZN(n4290) );
  INV_X1 U5839 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4385) );
  OR2_X1 U5840 ( .A1(n5680), .A2(n5675), .ZN(n4291) );
  AND2_X1 U5841 ( .A1(n4710), .A2(n5852), .ZN(n4292) );
  AND2_X1 U5842 ( .A1(n4284), .A2(n4715), .ZN(n4293) );
  INV_X1 U5843 ( .A(n9113), .ZN(n8926) );
  OR2_X1 U5844 ( .A1(n7223), .A2(n4599), .ZN(n4294) );
  INV_X1 U5845 ( .A(n9301), .ZN(n4495) );
  NAND2_X1 U5846 ( .A1(n4975), .A2(n4341), .ZN(n4295) );
  NAND2_X1 U5847 ( .A1(n9695), .A2(n4504), .ZN(n4503) );
  AND2_X1 U5848 ( .A1(n7875), .A2(n8020), .ZN(n6713) );
  NAND2_X1 U5849 ( .A1(n4354), .A2(n4775), .ZN(n6540) );
  XNOR2_X1 U5850 ( .A(n5595), .B(n5594), .ZN(n8772) );
  AND2_X1 U5851 ( .A1(n4787), .A2(n7554), .ZN(n4296) );
  NAND2_X1 U5852 ( .A1(n8778), .A2(n8781), .ZN(n5099) );
  AND2_X1 U5853 ( .A1(n5038), .A2(n4640), .ZN(n5078) );
  NAND4_X1 U5854 ( .A1(n4866), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5481)
         );
  AND2_X1 U5855 ( .A1(n9037), .A2(n9035), .ZN(n4297) );
  AOI21_X1 U5856 ( .B1(n8543), .B2(n4653), .A(n4650), .ZN(n4649) );
  AND2_X1 U5857 ( .A1(n9306), .A2(n9038), .ZN(n4298) );
  INV_X1 U5858 ( .A(n8456), .ZN(n8738) );
  NAND2_X1 U5859 ( .A1(n5404), .A2(n5403), .ZN(n8456) );
  NAND2_X1 U5860 ( .A1(n5698), .A2(n5702), .ZN(n8441) );
  INV_X1 U5861 ( .A(n8441), .ZN(n4625) );
  OR2_X1 U5862 ( .A1(n6789), .A2(n6488), .ZN(n4299) );
  NOR2_X1 U5863 ( .A1(n4892), .A2(n5074), .ZN(n4300) );
  AND2_X1 U5864 ( .A1(n5601), .A2(n5712), .ZN(n4301) );
  AND2_X1 U5865 ( .A1(n6751), .A2(n5731), .ZN(n4302) );
  AND2_X1 U5866 ( .A1(n5727), .A2(n5709), .ZN(n4303) );
  INV_X1 U5867 ( .A(n4845), .ZN(n4844) );
  OR2_X1 U5868 ( .A1(n9028), .A2(n4846), .ZN(n4845) );
  AND2_X1 U5869 ( .A1(n8059), .A2(n8101), .ZN(n9039) );
  AND2_X1 U5870 ( .A1(n6492), .A2(n4773), .ZN(n4304) );
  AND2_X1 U5871 ( .A1(n5986), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4305) );
  AND2_X1 U5872 ( .A1(n5323), .A2(n5322), .ZN(n8754) );
  INV_X1 U5873 ( .A(n8754), .ZN(n8590) );
  NAND2_X1 U5874 ( .A1(n8053), .A2(n9065), .ZN(n9097) );
  INV_X1 U5875 ( .A(n9097), .ZN(n9096) );
  NAND2_X1 U5876 ( .A1(n4769), .A2(n7665), .ZN(n8815) );
  NOR2_X1 U5877 ( .A1(n9217), .A2(n9216), .ZN(n4494) );
  INV_X1 U5878 ( .A(n9161), .ZN(n4806) );
  AND2_X1 U5879 ( .A1(n4472), .A2(n4479), .ZN(n4306) );
  AND2_X1 U5880 ( .A1(n5685), .A2(n5679), .ZN(n8498) );
  NAND2_X1 U5881 ( .A1(n7807), .A2(n7806), .ZN(n9306) );
  AND2_X1 U5882 ( .A1(n5687), .A2(n5688), .ZN(n4307) );
  AND2_X1 U5883 ( .A1(n8470), .A2(n5691), .ZN(n4308) );
  AOI21_X1 U5884 ( .B1(n9187), .B2(n7971), .A(n9058), .ZN(n4808) );
  INV_X1 U5885 ( .A(n8610), .ZN(n8758) );
  NAND2_X1 U5886 ( .A1(n5308), .A2(n5307), .ZN(n8610) );
  OR2_X1 U5887 ( .A1(n8511), .A2(n8526), .ZN(n5685) );
  XOR2_X1 U5888 ( .A(n8389), .B(n8386), .Z(n4309) );
  NOR2_X1 U5889 ( .A1(n4475), .A2(n4927), .ZN(n4474) );
  INV_X1 U5890 ( .A(n4688), .ZN(n4687) );
  NAND2_X1 U5891 ( .A1(n4689), .A2(n4961), .ZN(n4688) );
  AND2_X1 U5892 ( .A1(n5091), .A2(n4666), .ZN(n4310) );
  AND2_X1 U5893 ( .A1(n4301), .A2(n8726), .ZN(n4311) );
  AND2_X1 U5894 ( .A1(n4853), .A2(n4852), .ZN(n4312) );
  NAND2_X1 U5895 ( .A1(n5339), .A2(n5338), .ZN(n8676) );
  INV_X1 U5896 ( .A(n7526), .ZN(n8272) );
  AND2_X1 U5897 ( .A1(n5466), .A2(n5465), .ZN(n7526) );
  AND2_X1 U5898 ( .A1(n9142), .A2(n9127), .ZN(n4313) );
  AND2_X1 U5899 ( .A1(n4297), .A2(n9039), .ZN(n4314) );
  AND2_X1 U5900 ( .A1(n4301), .A2(n4619), .ZN(n4315) );
  AND2_X1 U5901 ( .A1(n5711), .A2(n8406), .ZN(n4316) );
  OR2_X1 U5902 ( .A1(n10034), .A2(n9286), .ZN(n9044) );
  AND2_X1 U5903 ( .A1(n5606), .A2(n5643), .ZN(n7144) );
  INV_X1 U5904 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4591) );
  AND2_X1 U5905 ( .A1(n5626), .A2(n6910), .ZN(n4317) );
  NOR2_X1 U5906 ( .A1(n7493), .A2(n8280), .ZN(n4318) );
  XNOR2_X1 U5907 ( .A(n5843), .B(n9784), .ZN(n5761) );
  AND3_X1 U5908 ( .A1(n4422), .A2(n4421), .A3(n4434), .ZN(n4319) );
  NOR2_X1 U5909 ( .A1(n9479), .A2(n7369), .ZN(n4320) );
  NAND2_X1 U5910 ( .A1(n5955), .A2(n5954), .ZN(n4321) );
  NAND2_X1 U5911 ( .A1(n4542), .A2(n4540), .ZN(n9304) );
  AND2_X1 U5912 ( .A1(n9039), .A2(n4298), .ZN(n4322) );
  INV_X1 U5913 ( .A(n8108), .ZN(n4432) );
  AND2_X1 U5914 ( .A1(n7274), .A2(n7273), .ZN(n4323) );
  INV_X1 U5915 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9970) );
  INV_X1 U5916 ( .A(n5851), .ZN(n4710) );
  OR2_X1 U5917 ( .A1(n5012), .A2(n4690), .ZN(n4324) );
  INV_X1 U5918 ( .A(n6638), .ZN(n4837) );
  NAND2_X1 U5919 ( .A1(n4625), .A2(n4627), .ZN(n4325) );
  AND2_X1 U5920 ( .A1(n4926), .A2(SI_11_), .ZN(n4326) );
  AND2_X1 U5921 ( .A1(n8500), .A2(n5677), .ZN(n4327) );
  NOR2_X1 U5922 ( .A1(n8532), .A2(n8232), .ZN(n4328) );
  NOR2_X1 U5923 ( .A1(n8574), .A2(n8249), .ZN(n4329) );
  AND2_X1 U5924 ( .A1(n7972), .A2(n7971), .ZN(n9055) );
  AND2_X1 U5925 ( .A1(n8855), .A2(n4747), .ZN(n4330) );
  AND2_X1 U5926 ( .A1(n4807), .A2(n4806), .ZN(n4331) );
  AND2_X1 U5927 ( .A1(n4496), .A2(n4495), .ZN(n4332) );
  AND2_X1 U5928 ( .A1(n7442), .A2(n5661), .ZN(n7485) );
  AND2_X1 U5929 ( .A1(n4768), .A2(n8871), .ZN(n4333) );
  AND2_X1 U5930 ( .A1(n4624), .A2(n4622), .ZN(n4334) );
  OR2_X1 U5931 ( .A1(n4731), .A2(n4730), .ZN(n4335) );
  AND2_X1 U5932 ( .A1(n4753), .A2(n8900), .ZN(n4336) );
  NAND2_X1 U5933 ( .A1(n7959), .A2(n7958), .ZN(n9301) );
  NAND2_X1 U5934 ( .A1(n4273), .A2(n6158), .ZN(n6213) );
  AND2_X1 U5935 ( .A1(n5659), .A2(n5658), .ZN(n7318) );
  AND2_X1 U5936 ( .A1(n5531), .A2(n4591), .ZN(n4337) );
  NOR2_X1 U5937 ( .A1(n7275), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5938 ( .A1(n5836), .A2(n5837), .ZN(n4338) );
  INV_X1 U5939 ( .A(n5106), .ZN(n4588) );
  OR2_X1 U5940 ( .A1(n8381), .A2(n8380), .ZN(P2_U3264) );
  AND2_X1 U5941 ( .A1(n7141), .A2(n5189), .ZN(n7227) );
  INV_X1 U5942 ( .A(n7532), .ZN(n8406) );
  XNOR2_X1 U5943 ( .A(n5951), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6103) );
  INV_X1 U5944 ( .A(n4728), .ZN(n7429) );
  AND2_X1 U5945 ( .A1(n6542), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4340) );
  INV_X1 U5946 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U5947 ( .A1(n7672), .A2(n7671), .ZN(n9344) );
  NAND2_X1 U5948 ( .A1(n4975), .A2(n4738), .ZN(n5288) );
  AND2_X1 U5949 ( .A1(n4738), .A2(n4385), .ZN(n4341) );
  NAND2_X1 U5950 ( .A1(n4975), .A2(n4974), .ZN(n5262) );
  NOR2_X1 U5951 ( .A1(n5902), .A2(n8770), .ZN(n4342) );
  NOR2_X1 U5952 ( .A1(n8239), .A2(n5846), .ZN(n8229) );
  NAND2_X1 U5953 ( .A1(n8605), .A2(n4286), .ZN(n4594) );
  AND2_X1 U5954 ( .A1(n4717), .A2(n4718), .ZN(n4343) );
  AND2_X1 U5955 ( .A1(n4515), .A2(n4514), .ZN(n4344) );
  AND2_X1 U5956 ( .A1(n9339), .A2(n9022), .ZN(n4345) );
  INV_X1 U5957 ( .A(n4602), .ZN(n7324) );
  NOR2_X1 U5958 ( .A1(n7223), .A2(n7210), .ZN(n4602) );
  INV_X1 U5959 ( .A(n4598), .ZN(n7492) );
  NOR2_X1 U5960 ( .A1(n7223), .A2(n4600), .ZN(n4598) );
  AND2_X1 U5961 ( .A1(n6863), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4346) );
  INV_X1 U5962 ( .A(n9314), .ZN(n9120) );
  NAND2_X1 U5963 ( .A1(n7774), .A2(n7773), .ZN(n9314) );
  OR2_X1 U5964 ( .A1(n9246), .A2(n9263), .ZN(n4347) );
  NOR2_X1 U5965 ( .A1(n7534), .A2(n7533), .ZN(n4348) );
  NAND2_X1 U5966 ( .A1(n5374), .A2(n5373), .ZN(n8665) );
  OR2_X1 U5967 ( .A1(n7788), .A2(n7787), .ZN(n4349) );
  AND2_X1 U5968 ( .A1(n9306), .A2(n9679), .ZN(n4350) );
  INV_X1 U5969 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U5970 ( .A1(n7058), .A2(n7127), .ZN(n7107) );
  NAND2_X1 U5971 ( .A1(n7111), .A2(n4766), .ZN(n7276) );
  INV_X1 U5972 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n4740) );
  INV_X1 U5973 ( .A(n7555), .ZN(n4784) );
  NAND2_X1 U5974 ( .A1(n6636), .A2(n6635), .ZN(n6883) );
  AND2_X1 U5975 ( .A1(n7181), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5976 ( .A1(n4822), .A2(n6632), .ZN(n6724) );
  AND2_X1 U5977 ( .A1(n4545), .A2(n8084), .ZN(n4352) );
  OR2_X1 U5978 ( .A1(n6886), .A2(n9678), .ZN(n6887) );
  INV_X1 U5979 ( .A(n6887), .ZN(n4502) );
  INV_X1 U5980 ( .A(n8163), .ZN(n4715) );
  AND2_X1 U5981 ( .A1(n5573), .A2(SI_29_), .ZN(n4353) );
  AND2_X1 U5982 ( .A1(n4774), .A2(n6494), .ZN(n4354) );
  NOR2_X1 U5983 ( .A1(n6861), .A2(n4826), .ZN(n4355) );
  AND2_X1 U5984 ( .A1(n4775), .A2(n4774), .ZN(n4356) );
  INV_X1 U5985 ( .A(n6803), .ZN(n4504) );
  OR2_X1 U5986 ( .A1(n9777), .A2(n5747), .ZN(n9826) );
  AND2_X1 U5987 ( .A1(n6246), .A2(n6245), .ZN(n9632) );
  OR2_X1 U5988 ( .A1(n8068), .A2(n8123), .ZN(n9287) );
  INV_X1 U5989 ( .A(n7964), .ZN(n4448) );
  AND2_X1 U5990 ( .A1(n6550), .A2(n6549), .ZN(n4357) );
  INV_X1 U5991 ( .A(n4469), .ZN(n9642) );
  OR2_X1 U5992 ( .A1(n7019), .A2(n9651), .ZN(n4469) );
  NOR2_X1 U5993 ( .A1(n5525), .A2(n4743), .ZN(n8773) );
  INV_X1 U5994 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U5995 ( .A1(n4359), .A2(n4358), .ZN(P1_U3240) );
  OAI21_X1 U5996 ( .B1(n8070), .B2(n4669), .A(n4360), .ZN(n4359) );
  NAND2_X1 U5997 ( .A1(n6662), .A2(n8081), .ZN(n6771) );
  MUX2_X1 U5998 ( .A(n7897), .B(n7896), .S(n4448), .Z(n7908) );
  NAND2_X1 U5999 ( .A1(n6160), .A2(n5036), .ZN(n6161) );
  NAND2_X1 U6000 ( .A1(n6247), .A2(n7979), .ZN(n6660) );
  NAND2_X1 U6001 ( .A1(n7978), .A2(n8078), .ZN(n6661) );
  NAND2_X1 U6002 ( .A1(n7965), .A2(n7966), .ZN(n4371) );
  NAND2_X1 U6003 ( .A1(n7873), .A2(n4448), .ZN(n4447) );
  NAND2_X2 U6004 ( .A1(n7205), .A2(n7209), .ZN(n7204) );
  NAND2_X1 U6005 ( .A1(n4611), .A2(n4609), .ZN(n8594) );
  AOI21_X1 U6006 ( .B1(n4881), .B2(n4451), .A(n4450), .ZN(n4449) );
  INV_X1 U6007 ( .A(n5752), .ZN(n4378) );
  NAND2_X1 U6008 ( .A1(n7330), .A2(n5607), .ZN(n4628) );
  NAND2_X1 U6009 ( .A1(n4375), .A2(n5751), .ZN(n5756) );
  OAI21_X2 U6010 ( .B1(n8180), .B2(n8182), .A(n8181), .ZN(n5858) );
  OAI21_X1 U6011 ( .B1(n5820), .B2(n4730), .A(n4729), .ZN(n5825) );
  NAND2_X1 U6012 ( .A1(n4714), .A2(n4712), .ZN(n8222) );
  NOR2_X2 U6013 ( .A1(n5861), .A2(n5860), .ZN(n7523) );
  INV_X1 U6014 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6015 ( .A1(n4734), .A2(n5810), .ZN(n7160) );
  NAND2_X1 U6016 ( .A1(n5765), .A2(n6506), .ZN(n6513) );
  NAND2_X1 U6017 ( .A1(n4976), .A2(n4740), .ZN(n4739) );
  AOI21_X1 U6018 ( .B1(n5932), .B2(n5780), .A(n5779), .ZN(n6579) );
  OR2_X1 U6019 ( .A1(n4275), .A2(n5033), .ZN(n4372) );
  NAND2_X4 U6020 ( .A1(n4810), .A2(n4809), .ZN(n6156) );
  INV_X1 U6021 ( .A(n4477), .ZN(n4473) );
  INV_X1 U6022 ( .A(n5194), .ZN(n4920) );
  NAND2_X1 U6023 ( .A1(n5335), .A2(n5334), .ZN(n5337) );
  NAND2_X1 U6024 ( .A1(n4425), .A2(n4426), .ZN(n4421) );
  OAI21_X1 U6025 ( .B1(n5349), .B2(n4704), .A(n5353), .ZN(n5366) );
  INV_X1 U6026 ( .A(n5920), .ZN(n4547) );
  NAND2_X1 U6027 ( .A1(n4752), .A2(n4756), .ZN(n8897) );
  NAND3_X1 U6028 ( .A1(n7585), .A2(n8795), .A3(n7586), .ZN(n8912) );
  NAND2_X1 U6029 ( .A1(n4683), .A2(n4681), .ZN(n5335) );
  NAND2_X1 U6030 ( .A1(n4435), .A2(n9301), .ZN(n4428) );
  INV_X1 U6031 ( .A(n7057), .ZN(n7054) );
  NAND2_X1 U6032 ( .A1(n7048), .A2(n7047), .ZN(n7057) );
  NAND2_X1 U6033 ( .A1(n8864), .A2(n4759), .ZN(n8839) );
  NAND2_X1 U6034 ( .A1(n5088), .A2(n5087), .ZN(n5073) );
  NAND2_X1 U6035 ( .A1(n6990), .A2(n6989), .ZN(n4734) );
  NAND2_X1 U6036 ( .A1(n5825), .A2(n5824), .ZN(n8192) );
  NAND2_X1 U6037 ( .A1(n5530), .A2(n4337), .ZN(n5527) );
  AOI21_X2 U6038 ( .B1(n6443), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6464), .ZN(
        n6441) );
  AOI21_X2 U6039 ( .B1(n6452), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6451), .ZN(
        n6454) );
  AOI21_X2 U6040 ( .B1(n8325), .B2(P2_REG1_REG_10__SCAN_IN), .A(n8326), .ZN(
        n6694) );
  NAND2_X2 U6041 ( .A1(n7389), .A2(n7388), .ZN(n7556) );
  NAND2_X1 U6042 ( .A1(n5927), .A2(n4863), .ZN(n4374) );
  NAND3_X1 U6043 ( .A1(n5750), .A2(n4378), .A3(n4376), .ZN(n4375) );
  NAND2_X1 U6044 ( .A1(n5015), .A2(n5014), .ZN(n5471) );
  NAND2_X1 U6045 ( .A1(n5015), .A2(n4381), .ZN(n5477) );
  NAND2_X1 U6046 ( .A1(n5015), .A2(n4379), .ZN(n4382) );
  NAND2_X1 U6047 ( .A1(n4384), .A2(n4975), .ZN(n5318) );
  NAND3_X1 U6048 ( .A1(n4582), .A2(n4387), .A3(n4388), .ZN(n4386) );
  AND2_X1 U6049 ( .A1(n4388), .A2(n4579), .ZN(n4397) );
  OR2_X1 U6050 ( .A1(n4585), .A2(n5674), .ZN(n4388) );
  NAND2_X1 U6051 ( .A1(n4582), .A2(n4397), .ZN(n5681) );
  INV_X1 U6052 ( .A(n5682), .ZN(n4398) );
  OAI21_X1 U6053 ( .B1(n4402), .B2(n4401), .A(n4399), .ZN(n4412) );
  NAND3_X1 U6054 ( .A1(n4405), .A2(n4404), .A3(n5721), .ZN(n4413) );
  NAND2_X1 U6055 ( .A1(n6660), .A2(n4420), .ZN(n8078) );
  XNOR2_X1 U6056 ( .A(n6241), .B(n6163), .ZN(n7979) );
  OR2_X1 U6057 ( .A1(n4425), .A2(n4427), .ZN(n4424) );
  XNOR2_X2 U6058 ( .A(n6092), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5967) );
  AOI21_X1 U6059 ( .B1(n7916), .B2(n4436), .A(n4437), .ZN(n7921) );
  OAI21_X1 U6060 ( .B1(n7932), .B2(n4448), .A(n7935), .ZN(n4443) );
  NOR2_X1 U6061 ( .A1(n7933), .A2(n7964), .ZN(n4444) );
  NAND2_X1 U6062 ( .A1(n4447), .A2(n4445), .ZN(n7890) );
  AOI21_X1 U6063 ( .B1(n4446), .B2(n7964), .A(n7876), .ZN(n4445) );
  NAND2_X1 U6064 ( .A1(n6714), .A2(n8017), .ZN(n7872) );
  OAI21_X1 U6065 ( .B1(n4453), .B2(n5035), .A(n4449), .ZN(n4885) );
  INV_X1 U6066 ( .A(n5034), .ZN(n4451) );
  XNOR2_X1 U6067 ( .A(n4880), .B(n4879), .ZN(n5035) );
  NAND2_X1 U6068 ( .A1(n6861), .A2(n7009), .ZN(n4457) );
  NOR2_X2 U6069 ( .A1(n9205), .A2(n9339), .ZN(n9190) );
  NOR2_X2 U6070 ( .A1(n9229), .A2(n9349), .ZN(n9220) );
  AND2_X1 U6071 ( .A1(n9129), .A2(n4498), .ZN(n9101) );
  NAND2_X1 U6072 ( .A1(n9129), .A2(n9120), .ZN(n9114) );
  NAND2_X1 U6073 ( .A1(n4502), .A2(n4499), .ZN(n7012) );
  MUX2_X1 U6074 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n6156), .Z(n5034) );
  MUX2_X1 U6075 ( .A(n6301), .B(n5989), .S(n6156), .Z(n4891) );
  MUX2_X1 U6076 ( .A(n6014), .B(n9959), .S(n6156), .Z(n4906) );
  MUX2_X1 U6077 ( .A(n4909), .B(n6026), .S(n6156), .Z(n4917) );
  MUX2_X1 U6078 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6156), .Z(n4902) );
  MUX2_X1 U6079 ( .A(n6031), .B(n4924), .S(n6156), .Z(n4925) );
  MUX2_X1 U6080 ( .A(n6124), .B(n6126), .S(n6156), .Z(n4941) );
  MUX2_X1 U6081 ( .A(n4956), .B(n6342), .S(n6156), .Z(n4957) );
  MUX2_X1 U6082 ( .A(n7670), .B(n6859), .S(n6156), .Z(n4970) );
  MUX2_X1 U6083 ( .A(n7712), .B(n6988), .S(n6156), .Z(n5354) );
  MUX2_X1 U6084 ( .A(n10002), .B(n7177), .S(n6156), .Z(n5394) );
  XNOR2_X1 U6085 ( .A(n8952), .B(n8958), .ZN(n7293) );
  INV_X1 U6086 ( .A(n4521), .ZN(n9504) );
  NOR2_X1 U6087 ( .A1(n5969), .A2(n5968), .ZN(n6263) );
  NAND2_X1 U6088 ( .A1(n9143), .A2(n4526), .ZN(n4525) );
  NAND2_X1 U6089 ( .A1(n9143), .A2(n4530), .ZN(n4527) );
  NAND3_X1 U6090 ( .A1(n9096), .A2(n4280), .A3(n8005), .ZN(n4524) );
  INV_X1 U6091 ( .A(n9064), .ZN(n4535) );
  NOR2_X1 U6092 ( .A1(n6707), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U6093 ( .A1(n6714), .A2(n8083), .ZN(n4545) );
  INV_X1 U6094 ( .A(n5996), .ZN(n4546) );
  NAND3_X1 U6095 ( .A1(n4547), .A2(n4546), .A3(n4861), .ZN(n6086) );
  NAND3_X1 U6096 ( .A1(n9457), .A2(n4802), .A3(n8023), .ZN(n4801) );
  NAND2_X1 U6097 ( .A1(n4554), .A2(n4553), .ZN(n5664) );
  AND2_X1 U6098 ( .A1(n5660), .A2(n7485), .ZN(n4553) );
  NAND2_X1 U6099 ( .A1(n4555), .A2(n7318), .ZN(n4554) );
  OAI21_X1 U6100 ( .B1(n5657), .B2(n4556), .A(n5656), .ZN(n4555) );
  NAND2_X1 U6101 ( .A1(n5646), .A2(n7209), .ZN(n4556) );
  NAND2_X1 U6102 ( .A1(n5629), .A2(n4302), .ZN(n4561) );
  NAND4_X1 U6103 ( .A1(n4565), .A2(n4568), .A3(n4562), .A4(n4567), .ZN(n4559)
         );
  NAND2_X1 U6104 ( .A1(n4317), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U6105 ( .A1(n5625), .A2(n4564), .ZN(n4563) );
  OR2_X1 U6106 ( .A1(n5624), .A2(n4566), .ZN(n4565) );
  OAI21_X1 U6107 ( .B1(n4578), .B2(n4577), .A(n4574), .ZN(n4573) );
  AOI21_X1 U6108 ( .B1(n5689), .B2(n4307), .A(n5697), .ZN(n4578) );
  OR2_X1 U6109 ( .A1(n5672), .A2(n5671), .ZN(n4585) );
  NAND3_X1 U6110 ( .A1(n4736), .A2(n4975), .A3(n5531), .ZN(n5525) );
  INV_X1 U6111 ( .A(n4594), .ZN(n8547) );
  INV_X1 U6112 ( .A(n4597), .ZN(n8628) );
  INV_X1 U6113 ( .A(n4606), .ZN(n8423) );
  NAND2_X1 U6114 ( .A1(n4615), .A2(n4315), .ZN(n4618) );
  NAND2_X1 U6115 ( .A1(n5585), .A2(n5716), .ZN(n4615) );
  XNOR2_X1 U6116 ( .A(n4616), .B(n8433), .ZN(n5602) );
  NAND3_X1 U6117 ( .A1(n4618), .A2(n4617), .A3(n5715), .ZN(n4616) );
  OAI21_X2 U6118 ( .B1(n8434), .B2(n4325), .A(n4620), .ZN(n5509) );
  NAND2_X2 U6119 ( .A1(n4628), .A2(n5644), .ZN(n7218) );
  NAND2_X2 U6120 ( .A1(n7315), .A2(n4629), .ZN(n7487) );
  NAND2_X2 U6121 ( .A1(n7204), .A2(n4631), .ZN(n7315) );
  OAI21_X2 U6122 ( .B1(n5571), .B2(n5710), .A(n5726), .ZN(n5585) );
  NOR2_X2 U6123 ( .A1(n5560), .A2(n5559), .ZN(n5887) );
  NAND2_X1 U6124 ( .A1(n5730), .A2(n6972), .ZN(n6975) );
  NAND2_X1 U6125 ( .A1(n5042), .A2(n5041), .ZN(n5483) );
  NOR2_X1 U6126 ( .A1(n5509), .A2(n5743), .ZN(n5560) );
  NAND2_X1 U6127 ( .A1(n5492), .A2(n5491), .ZN(n7073) );
  NAND3_X1 U6128 ( .A1(n5487), .A2(n5732), .A3(n5486), .ZN(n6835) );
  NAND2_X1 U6129 ( .A1(n6975), .A2(n5615), .ZN(n6845) );
  NAND2_X1 U6130 ( .A1(n5483), .A2(n5482), .ZN(n6970) );
  NAND2_X1 U6131 ( .A1(n5494), .A2(n5643), .ZN(n7330) );
  NAND2_X1 U6132 ( .A1(n4633), .A2(n9811), .ZN(n5114) );
  NAND3_X1 U6133 ( .A1(n5107), .A2(n5108), .A3(n6837), .ZN(n4633) );
  NAND3_X1 U6134 ( .A1(n6598), .A2(n4875), .A3(n6599), .ZN(n4634) );
  NAND2_X1 U6135 ( .A1(n6910), .A2(n4875), .ZN(n4635) );
  INV_X2 U6136 ( .A(n5247), .ZN(n4975) );
  NOR2_X1 U6137 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4640) );
  NAND2_X1 U6138 ( .A1(n5274), .A2(n4644), .ZN(n4643) );
  NAND3_X1 U6139 ( .A1(n8501), .A2(n4654), .A3(n4655), .ZN(n4652) );
  NAND2_X1 U6140 ( .A1(n4659), .A2(n4661), .ZN(n5333) );
  NAND2_X1 U6141 ( .A1(n8600), .A2(n4662), .ZN(n4659) );
  INV_X1 U6142 ( .A(n4665), .ZN(n8602) );
  NAND2_X1 U6143 ( .A1(n5076), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U6144 ( .A1(n7075), .A2(n4668), .ZN(n7141) );
  NAND2_X1 U6145 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  NAND2_X1 U6146 ( .A1(n4672), .A2(n9193), .ZN(n4671) );
  NAND2_X1 U6147 ( .A1(n4673), .A2(n8067), .ZN(n4672) );
  NAND2_X1 U6148 ( .A1(n4253), .A2(n4674), .ZN(n4673) );
  INV_X1 U6149 ( .A(n8068), .ZN(n4674) );
  NAND2_X1 U6150 ( .A1(n5303), .A2(n4685), .ZN(n4683) );
  XNOR2_X1 U6151 ( .A(n4692), .B(n5430), .ZN(n7771) );
  NAND2_X1 U6152 ( .A1(n4940), .A2(n4696), .ZN(n4693) );
  NAND2_X1 U6153 ( .A1(n4693), .A2(n4694), .ZN(n4955) );
  NAND2_X1 U6154 ( .A1(n4940), .A2(n4939), .ZN(n5261) );
  INV_X2 U6155 ( .A(n6156), .ZN(n5367) );
  NAND3_X1 U6156 ( .A1(n4809), .A2(n4810), .A3(n6181), .ZN(n4705) );
  OAI21_X1 U6157 ( .B1(n8229), .B2(n5851), .A(n4708), .ZN(n4707) );
  INV_X1 U6158 ( .A(n4707), .ZN(n8151) );
  INV_X1 U6159 ( .A(n8229), .ZN(n4711) );
  NAND2_X1 U6160 ( .A1(n4711), .A2(n4292), .ZN(n8149) );
  INV_X1 U6161 ( .A(n5852), .ZN(n4708) );
  NAND2_X1 U6162 ( .A1(n8149), .A2(n8152), .ZN(n4709) );
  NAND2_X1 U6163 ( .A1(n8206), .A2(n4293), .ZN(n4714) );
  OAI21_X1 U6164 ( .B1(n5861), .B2(n4725), .A(n4723), .ZN(n7538) );
  NAND2_X1 U6165 ( .A1(n4721), .A2(n4720), .ZN(n7536) );
  NAND2_X1 U6166 ( .A1(n5861), .A2(n4723), .ZN(n4721) );
  INV_X1 U6167 ( .A(n7300), .ZN(n4733) );
  AND2_X1 U6168 ( .A1(n5801), .A2(n6953), .ZN(n4735) );
  NOR2_X2 U6169 ( .A1(n4737), .A2(n4981), .ZN(n4736) );
  AND2_X1 U6170 ( .A1(n5794), .A2(n5789), .ZN(n4741) );
  NAND2_X2 U6171 ( .A1(n5785), .A2(n6580), .ZN(n6586) );
  NAND2_X1 U6172 ( .A1(n8846), .A2(n7607), .ZN(n4746) );
  NAND2_X1 U6173 ( .A1(n4746), .A2(n4330), .ZN(n7626) );
  NAND2_X1 U6174 ( .A1(n8863), .A2(n8865), .ZN(n8864) );
  NAND2_X1 U6175 ( .A1(n4749), .A2(n4336), .ZN(n8899) );
  NAND2_X1 U6176 ( .A1(n4266), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U6177 ( .A1(n7770), .A2(n7769), .ZN(n4760) );
  NAND3_X1 U6178 ( .A1(n7058), .A2(n4764), .A3(n7127), .ZN(n4761) );
  INV_X1 U6179 ( .A(n4262), .ZN(n4769) );
  NAND2_X1 U6180 ( .A1(n4767), .A2(n4333), .ZN(n7688) );
  NAND2_X1 U6181 ( .A1(n8817), .A2(n7668), .ZN(n4767) );
  NAND2_X1 U6182 ( .A1(n7556), .A2(n7554), .ZN(n4776) );
  OAI21_X1 U6183 ( .B1(n7556), .B2(n7555), .A(n4296), .ZN(n8796) );
  NAND2_X1 U6184 ( .A1(n7556), .A2(n4296), .ZN(n4778) );
  OAI21_X1 U6185 ( .B1(n7556), .B2(n4783), .A(n4779), .ZN(n7588) );
  INV_X1 U6186 ( .A(n4785), .ZN(n4781) );
  INV_X1 U6187 ( .A(n8798), .ZN(n4782) );
  AOI21_X1 U6188 ( .B1(n8798), .B2(n4784), .A(n4785), .ZN(n4783) );
  INV_X1 U6189 ( .A(n7566), .ZN(n4787) );
  NAND2_X1 U6190 ( .A1(n4789), .A2(n4788), .ZN(n6012) );
  NOR2_X1 U6191 ( .A1(n5993), .A2(n4790), .ZN(n6007) );
  OAI21_X1 U6192 ( .B1(n6058), .B2(n4795), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5951) );
  INV_X1 U6193 ( .A(n4792), .ZN(n5949) );
  OAI21_X1 U6194 ( .B1(n6058), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U6195 ( .A1(n4801), .A2(n4798), .ZN(n9239) );
  NAND3_X1 U6196 ( .A1(n4809), .A2(n4810), .A3(n4877), .ZN(n6083) );
  NAND3_X1 U6197 ( .A1(n4822), .A2(n6632), .A3(n6633), .ZN(n6723) );
  AND2_X1 U6198 ( .A1(n7063), .A2(n8930), .ZN(n4826) );
  NAND2_X1 U6199 ( .A1(n9036), .A2(n4297), .ZN(n9081) );
  OAI211_X1 U6200 ( .C1(n9036), .C2(n4830), .A(n4828), .B(n4827), .ZN(n9298)
         );
  AND2_X1 U6201 ( .A1(n9036), .A2(n9035), .ZN(n4864) );
  NAND2_X1 U6202 ( .A1(n4838), .A2(n4840), .ZN(n9030) );
  NAND2_X1 U6203 ( .A1(n9025), .A2(n4842), .ZN(n4838) );
  NAND2_X1 U6204 ( .A1(n9025), .A2(n4848), .ZN(n4847) );
  NAND2_X1 U6205 ( .A1(n9198), .A2(n4283), .ZN(n4850) );
  NAND2_X1 U6206 ( .A1(n4850), .A2(n4851), .ZN(n9168) );
  INV_X1 U6207 ( .A(n9168), .ZN(n9023) );
  NAND2_X1 U6208 ( .A1(n7186), .A2(n4858), .ZN(n4857) );
  OR2_X1 U6209 ( .A1(n9777), .A2(n5550), .ZN(n9835) );
  NAND2_X1 U6210 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  CLKBUF_X1 U6211 ( .A(n6505), .Z(n8290) );
  NAND2_X2 U6212 ( .A1(n8521), .A2(n5505), .ZN(n8503) );
  NAND2_X1 U6213 ( .A1(n6513), .A2(n5769), .ZN(n5935) );
  NOR2_X1 U6214 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  AOI21_X2 U6215 ( .B1(n8192), .B2(n5831), .A(n5830), .ZN(n8206) );
  NAND2_X1 U6216 ( .A1(n9023), .A2(n4871), .ZN(n9025) );
  INV_X1 U6217 ( .A(n6016), .ZN(n6019) );
  OAI22_X2 U6218 ( .A1(n8174), .A2(n8173), .B1(n5845), .B2(n5844), .ZN(n5847)
         );
  NOR2_X1 U6219 ( .A1(n5463), .A2(n5066), .ZN(n4865) );
  OR2_X1 U6220 ( .A1(n5463), .A2(n5043), .ZN(n4866) );
  OR2_X1 U6221 ( .A1(n6215), .A2(n6181), .ZN(n4867) );
  INV_X1 U6222 ( .A(n8923), .ZN(n8898) );
  INV_X1 U6223 ( .A(n10037), .ZN(n9644) );
  INV_X1 U6224 ( .A(n6075), .ZN(n6132) );
  INV_X1 U6225 ( .A(n8927), .ZN(n9128) );
  AND2_X1 U6226 ( .A1(n5778), .A2(n5777), .ZN(n4868) );
  INV_X1 U6227 ( .A(n8526), .ZN(n8493) );
  AND3_X1 U6228 ( .A1(n5363), .A2(n5362), .A3(n5361), .ZN(n8526) );
  AND2_X1 U6229 ( .A1(n4939), .A2(n4938), .ZN(n4869) );
  NAND2_X1 U6230 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4870) );
  OR2_X1 U6231 ( .A1(n9181), .A2(n9189), .ZN(n4871) );
  NOR2_X1 U6232 ( .A1(n4899), .A2(n4898), .ZN(n4872) );
  AND2_X1 U6233 ( .A1(n7074), .A2(n9820), .ZN(n4873) );
  NOR2_X1 U6234 ( .A1(n4920), .A2(n5192), .ZN(n4874) );
  INV_X1 U6235 ( .A(n9292), .ZN(n10041) );
  INV_X1 U6236 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5989) );
  AND2_X1 U6237 ( .A1(n7819), .A2(n7818), .ZN(n9100) );
  AOI21_X1 U6238 ( .B1(n8439), .B2(n5027), .A(n5428), .ZN(n8184) );
  NAND2_X1 U6239 ( .A1(n9840), .A2(n9812), .ZN(n8770) );
  AND2_X2 U6240 ( .A1(n5554), .A2(n6589), .ZN(n9840) );
  INV_X1 U6241 ( .A(n9840), .ZN(n5900) );
  AND4_X1 U6242 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8620)
         );
  AND2_X1 U6243 ( .A1(n5094), .A2(n9748), .ZN(n4875) );
  INV_X1 U6244 ( .A(n8244), .ZN(n5866) );
  OR2_X1 U6245 ( .A1(n5879), .A2(n5865), .ZN(n8244) );
  INV_X1 U6246 ( .A(n8719), .ZN(n5551) );
  AND2_X1 U6247 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  AND2_X1 U6248 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  INV_X1 U6249 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6250 ( .A1(n9314), .A2(n8927), .ZN(n9031) );
  INV_X1 U6251 ( .A(n9100), .ZN(n9038) );
  AND2_X1 U6252 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  INV_X1 U6253 ( .A(n5326), .ZN(n5002) );
  INV_X1 U6254 ( .A(n5388), .ZN(n5386) );
  OR2_X1 U6255 ( .A1(n8424), .A2(n8273), .ZN(n5450) );
  INV_X1 U6256 ( .A(n8620), .ZN(n5315) );
  INV_X1 U6257 ( .A(n5116), .ZN(n4994) );
  INV_X1 U6258 ( .A(n6488), .ZN(n7793) );
  INV_X1 U6259 ( .A(n7735), .ZN(n6389) );
  INV_X1 U6260 ( .A(n6555), .ZN(n6380) );
  OR2_X1 U6261 ( .A1(n9319), .A2(n9147), .ZN(n9029) );
  INV_X1 U6262 ( .A(n7631), .ZN(n6386) );
  INV_X1 U6263 ( .A(n6870), .ZN(n6382) );
  INV_X1 U6264 ( .A(n7874), .ZN(n6635) );
  OR2_X1 U6265 ( .A1(n6075), .A2(n8994), .ZN(n7964) );
  INV_X1 U6266 ( .A(n4921), .ZN(n4922) );
  INV_X1 U6267 ( .A(n5146), .ZN(n4901) );
  INV_X1 U6268 ( .A(n5137), .ZN(n4995) );
  NAND2_X1 U6269 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5097) );
  NAND2_X1 U6270 ( .A1(n5386), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6271 ( .A1(n4279), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6272 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4984), .ZN(n4985) );
  NAND2_X1 U6273 ( .A1(n5709), .A2(n5708), .ZN(n5743) );
  NAND2_X1 U6274 ( .A1(n5405), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5424) );
  OR2_X1 U6275 ( .A1(n5267), .A2(n7100), .ZN(n5295) );
  OR2_X1 U6276 ( .A1(n5217), .A2(n4997), .ZN(n5240) );
  OR2_X1 U6277 ( .A1(n8688), .A2(n8539), .ZN(n5332) );
  OAI21_X1 U6278 ( .B1(n6909), .B2(n6837), .A(n5114), .ZN(n6829) );
  INV_X1 U6279 ( .A(n7404), .ZN(n6384) );
  INV_X1 U6280 ( .A(n8849), .ZN(n7604) );
  INV_X1 U6281 ( .A(n8818), .ZN(n7665) );
  NAND2_X1 U6282 ( .A1(n6389), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U6283 ( .A1(n6385), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U6284 ( .A1(n6390), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U6285 ( .A1(n6386), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U6286 ( .A1(n6382), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U6287 ( .A1(n6381), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6664) );
  INV_X1 U6288 ( .A(n5260), .ZN(n4944) );
  NAND2_X1 U6289 ( .A1(n4929), .A2(n4928), .ZN(n4932) );
  INV_X1 U6290 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6291 ( .A1(n4995), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5153) );
  AND2_X1 U6292 ( .A1(n5776), .A2(n6527), .ZN(n6528) );
  AND2_X1 U6293 ( .A1(n5840), .A2(n5839), .ZN(n8163) );
  NOR2_X1 U6294 ( .A1(n8526), .A2(n7525), .ZN(n5846) );
  OR2_X1 U6295 ( .A1(n8408), .A2(n5510), .ZN(n5466) );
  NOR2_X1 U6296 ( .A1(n8327), .A2(n8328), .ZN(n8326) );
  NAND2_X1 U6297 ( .A1(n8383), .A2(n8271), .ZN(n5891) );
  AND2_X1 U6298 ( .A1(n5728), .A2(n8559), .ZN(n8583) );
  AND2_X1 U6299 ( .A1(n5508), .A2(n5480), .ZN(n6353) );
  INV_X1 U6300 ( .A(n8400), .ZN(n5902) );
  AND2_X1 U6301 ( .A1(n9768), .A2(n9771), .ZN(n5548) );
  NAND2_X1 U6302 ( .A1(n6384), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7576) );
  OR2_X1 U6303 ( .A1(n7737), .A2(n9958), .ZN(n7757) );
  INV_X1 U6304 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7117) );
  INV_X1 U6305 ( .A(n9306), .ZN(n9092) );
  INV_X1 U6306 ( .A(n9158), .ZN(n9189) );
  INV_X1 U6307 ( .A(n9453), .ZN(n9262) );
  NOR2_X1 U6308 ( .A1(n10034), .A2(n9436), .ZN(n9012) );
  INV_X1 U6309 ( .A(n8930), .ZN(n7121) );
  OR2_X1 U6310 ( .A1(n6286), .A2(n6244), .ZN(n9458) );
  NAND2_X1 U6311 ( .A1(n7569), .A2(n9405), .ZN(n6085) );
  AND2_X1 U6312 ( .A1(n8045), .A2(n9047), .ZN(n9264) );
  NAND2_X1 U6313 ( .A1(n9044), .A2(n8024), .ZN(n9448) );
  INV_X1 U6314 ( .A(n7063), .ZN(n9702) );
  INV_X1 U6315 ( .A(n8935), .ZN(n6774) );
  AND2_X1 U6316 ( .A1(n4954), .A2(n4953), .ZN(n5286) );
  OR3_X1 U6317 ( .A1(n7179), .A2(n5547), .A3(n7375), .ZN(n6351) );
  NAND2_X1 U6318 ( .A1(n8141), .A2(n8140), .ZN(n8143) );
  INV_X1 U6319 ( .A(n8266), .ZN(n8251) );
  OR2_X1 U6320 ( .A1(n5871), .A2(n9767), .ZN(n5879) );
  AND2_X1 U6321 ( .A1(n5449), .A2(n5448), .ZN(n8437) );
  AND4_X1 U6322 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n8596)
         );
  INV_X1 U6323 ( .A(n6344), .ZN(n9410) );
  INV_X1 U6324 ( .A(n8370), .ZN(n9722) );
  AND2_X1 U6325 ( .A1(n5442), .A2(n5425), .ZN(n8439) );
  INV_X1 U6326 ( .A(n8612), .ZN(n8634) );
  AND2_X1 U6327 ( .A1(n6353), .A2(n6350), .ZN(n9742) );
  OAI21_X1 U6328 ( .B1(n5902), .B2(n8719), .A(n5901), .ZN(n5903) );
  NOR2_X1 U6329 ( .A1(n9770), .A2(n5548), .ZN(n5864) );
  INV_X1 U6330 ( .A(n9835), .ZN(n9812) );
  NOR2_X1 U6331 ( .A1(n5546), .A2(n5863), .ZN(n5554) );
  INV_X1 U6332 ( .A(n7569), .ZN(n7648) );
  AND2_X1 U6333 ( .A1(n7811), .A2(n7776), .ZN(n9117) );
  OR2_X1 U6334 ( .A1(n9130), .A2(n4272), .ZN(n7764) );
  INV_X1 U6335 ( .A(n9034), .ZN(n9310) );
  AND2_X1 U6336 ( .A1(n8025), .A2(n9257), .ZN(n9284) );
  NAND2_X1 U6337 ( .A1(n6132), .A2(n8062), .ZN(n6286) );
  INV_X1 U6338 ( .A(n9705), .ZN(n9373) );
  NAND2_X1 U6339 ( .A1(n9656), .A2(n9682), .ZN(n9705) );
  AND2_X1 U6340 ( .A1(n6080), .A2(n6079), .ZN(n6257) );
  XNOR2_X1 U6341 ( .A(n6056), .B(n6057), .ZN(n6102) );
  AND2_X1 U6342 ( .A1(n6053), .A2(n6118), .ZN(n7181) );
  XNOR2_X1 U6343 ( .A(n4894), .B(SI_5_), .ZN(n5109) );
  INV_X1 U6344 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8379) );
  INV_X1 U6345 ( .A(n9731), .ZN(n9417) );
  OR2_X1 U6346 ( .A1(n5879), .A2(n5878), .ZN(n8264) );
  OR2_X1 U6347 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  INV_X1 U6348 ( .A(n8436), .ZN(n8275) );
  INV_X1 U6349 ( .A(n9424), .ZN(n9726) );
  INV_X1 U6350 ( .A(n9764), .ZN(n8584) );
  NAND2_X1 U6351 ( .A1(n9855), .A2(n9812), .ZN(n8719) );
  INV_X1 U6352 ( .A(n9855), .ZN(n9853) );
  INV_X1 U6353 ( .A(n8443), .ZN(n8734) );
  NOR2_X1 U6354 ( .A1(n5872), .A2(P2_U3152), .ZN(n9774) );
  XNOR2_X1 U6355 ( .A(n5540), .B(n5539), .ZN(n7179) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6117) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6026) );
  INV_X1 U6358 ( .A(n9323), .ZN(n9142) );
  AND2_X1 U6359 ( .A1(n6398), .A2(n6397), .ZN(n9085) );
  NAND2_X1 U6360 ( .A1(n7782), .A2(n7781), .ZN(n8927) );
  OR2_X1 U6361 ( .A1(n7617), .A2(n7616), .ZN(n9015) );
  INV_X1 U6362 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9518) );
  OAI21_X1 U6363 ( .B1(n4864), .B2(n9037), .A(n9081), .ZN(n9307) );
  OR2_X1 U6364 ( .A1(n9648), .A2(n6710), .ZN(n9292) );
  INV_X1 U6365 ( .A(n9721), .ZN(n9718) );
  INV_X1 U6366 ( .A(n9709), .ZN(n9707) );
  INV_X1 U6367 ( .A(n9393), .ZN(n6146) );
  INV_X1 U6368 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U6369 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  AND2_X1 U6370 ( .A1(n5931), .A2(n9774), .ZN(P2_U3966) );
  OAI21_X1 U6371 ( .B1(n7523), .B2(n5884), .A(n5883), .ZN(P2_U3242) );
  INV_X1 U6372 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5549) );
  AND2_X1 U6373 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4877) );
  AND2_X1 U6374 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4878) );
  INV_X1 U6375 ( .A(SI_1_), .ZN(n4879) );
  NAND2_X1 U6376 ( .A1(n4880), .A2(SI_1_), .ZN(n4881) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U6378 ( .A(n4882), .B(SI_2_), .ZN(n5059) );
  INV_X1 U6379 ( .A(n4882), .ZN(n4883) );
  NAND2_X1 U6380 ( .A1(n4883), .A2(SI_2_), .ZN(n4884) );
  MUX2_X1 U6381 ( .A(n9983), .B(n6216), .S(n6158), .Z(n4886) );
  INV_X1 U6382 ( .A(n4886), .ZN(n4887) );
  NAND2_X1 U6383 ( .A1(n4887), .A2(SI_3_), .ZN(n5072) );
  INV_X1 U6384 ( .A(n4891), .ZN(n4888) );
  NAND2_X1 U6385 ( .A1(n4888), .A2(SI_4_), .ZN(n4890) );
  AND2_X1 U6386 ( .A1(n5072), .A2(n4890), .ZN(n4889) );
  INV_X1 U6387 ( .A(n4890), .ZN(n4892) );
  INV_X1 U6388 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4893) );
  INV_X1 U6389 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6476) );
  MUX2_X1 U6390 ( .A(n4893), .B(n6476), .S(n6158), .Z(n4894) );
  INV_X1 U6391 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6392 ( .A1(n4895), .A2(SI_5_), .ZN(n5123) );
  MUX2_X1 U6393 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5367), .Z(n4897) );
  NAND2_X1 U6394 ( .A1(n4897), .A2(SI_6_), .ZN(n4896) );
  AND2_X1 U6395 ( .A1(n5123), .A2(n4896), .ZN(n4900) );
  INV_X1 U6396 ( .A(n4896), .ZN(n4899) );
  NAND2_X1 U6397 ( .A1(n4902), .A2(SI_7_), .ZN(n4903) );
  INV_X1 U6398 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6014) );
  INV_X1 U6399 ( .A(SI_8_), .ZN(n4905) );
  INV_X1 U6400 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6401 ( .A1(n4907), .A2(SI_8_), .ZN(n4908) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4909) );
  INV_X1 U6403 ( .A(n4917), .ZN(n4910) );
  INV_X1 U6404 ( .A(SI_10_), .ZN(n4911) );
  INV_X1 U6405 ( .A(n4912), .ZN(n4913) );
  NAND2_X1 U6406 ( .A1(n4913), .A2(SI_10_), .ZN(n4914) );
  INV_X1 U6407 ( .A(SI_9_), .ZN(n4916) );
  NAND2_X1 U6408 ( .A1(n4917), .A2(n4916), .ZN(n5180) );
  AND2_X1 U6409 ( .A1(n5177), .A2(n5180), .ZN(n4918) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4924) );
  INV_X1 U6411 ( .A(n4925), .ZN(n4926) );
  INV_X1 U6412 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6055) );
  MUX2_X1 U6413 ( .A(n9928), .B(n6055), .S(n6158), .Z(n4929) );
  INV_X1 U6414 ( .A(SI_12_), .ZN(n4928) );
  INV_X1 U6415 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6416 ( .A1(n4930), .A2(SI_12_), .ZN(n4931) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U6418 ( .A(n6117), .B(n4934), .S(n5367), .Z(n4936) );
  INV_X1 U6419 ( .A(SI_13_), .ZN(n4935) );
  NAND2_X1 U6420 ( .A1(n4936), .A2(n4935), .ZN(n4939) );
  INV_X1 U6421 ( .A(n4936), .ZN(n4937) );
  NAND2_X1 U6422 ( .A1(n4937), .A2(SI_13_), .ZN(n4938) );
  INV_X1 U6423 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6126) );
  INV_X1 U6424 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6124) );
  INV_X1 U6425 ( .A(n4941), .ZN(n4942) );
  NAND2_X1 U6426 ( .A1(n4942), .A2(SI_14_), .ZN(n4943) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6327) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7568) );
  MUX2_X1 U6429 ( .A(n6327), .B(n7568), .S(n6158), .Z(n4946) );
  INV_X1 U6430 ( .A(SI_15_), .ZN(n4945) );
  INV_X1 U6431 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6432 ( .A1(n4947), .A2(SI_15_), .ZN(n4948) );
  INV_X1 U6433 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6328) );
  INV_X1 U6434 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U6435 ( .A(n6328), .B(n6333), .S(n5367), .Z(n4951) );
  INV_X1 U6436 ( .A(SI_16_), .ZN(n4950) );
  NAND2_X1 U6437 ( .A1(n4951), .A2(n4950), .ZN(n4954) );
  INV_X1 U6438 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6439 ( .A1(n4952), .A2(SI_16_), .ZN(n4953) );
  INV_X1 U6440 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6342) );
  INV_X1 U6441 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4956) );
  XNOR2_X1 U6442 ( .A(n4957), .B(SI_17_), .ZN(n5302) );
  INV_X1 U6443 ( .A(n5302), .ZN(n4960) );
  INV_X1 U6444 ( .A(n4957), .ZN(n4958) );
  NAND2_X1 U6445 ( .A1(n4958), .A2(SI_17_), .ZN(n4959) );
  MUX2_X1 U6446 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6158), .Z(n4962) );
  XNOR2_X1 U6447 ( .A(n4962), .B(SI_18_), .ZN(n5316) );
  INV_X1 U6448 ( .A(n5316), .ZN(n4961) );
  NAND2_X1 U6449 ( .A1(n4962), .A2(SI_18_), .ZN(n4963) );
  INV_X1 U6450 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6624) );
  INV_X1 U6451 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6626) );
  MUX2_X1 U6452 ( .A(n6624), .B(n6626), .S(n5367), .Z(n4965) );
  INV_X1 U6453 ( .A(SI_19_), .ZN(n4964) );
  NAND2_X1 U6454 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  INV_X1 U6455 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6456 ( .A1(n4966), .A2(SI_19_), .ZN(n4967) );
  NAND2_X1 U6457 ( .A1(n4968), .A2(n4967), .ZN(n5012) );
  INV_X1 U6458 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6859) );
  INV_X1 U6459 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7670) );
  INV_X1 U6460 ( .A(SI_20_), .ZN(n4969) );
  NAND2_X1 U6461 ( .A1(n4970), .A2(n4969), .ZN(n5336) );
  INV_X1 U6462 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6463 ( .A1(n4971), .A2(SI_20_), .ZN(n4972) );
  XNOR2_X1 U6464 ( .A(n5335), .B(n5334), .ZN(n7669) );
  NOR2_X1 U6465 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4979) );
  NOR2_X1 U6466 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4978) );
  NOR2_X1 U6467 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4977) );
  NAND4_X1 U6468 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n4981)
         );
  INV_X1 U6469 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4982) );
  INV_X1 U6470 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5529) );
  OAI21_X1 U6471 ( .B1(n4983), .B2(n5529), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n4986) );
  NAND2_X2 U6472 ( .A1(n4987), .A2(n5004), .ZN(n6359) );
  NAND2_X1 U6473 ( .A1(n5527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4988) );
  INV_X1 U6474 ( .A(n4983), .ZN(n4989) );
  NAND2_X1 U6475 ( .A1(n7669), .A2(n5576), .ZN(n4992) );
  NAND2_X1 U6476 ( .A1(n5596), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n4991) );
  INV_X1 U6477 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6478 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n4997) );
  INV_X1 U6479 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6947) );
  INV_X1 U6480 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7100) );
  AND2_X1 U6481 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n4999) );
  INV_X1 U6482 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8250) );
  INV_X1 U6483 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U6484 ( .A1(n5021), .A2(n8223), .ZN(n5003) );
  AND2_X1 U6485 ( .A1(n5341), .A2(n5003), .ZN(n8548) );
  NAND2_X1 U6486 ( .A1(n8548), .A2(n5027), .ZN(n5011) );
  NAND2_X1 U6487 ( .A1(n5067), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6488 ( .A1(n4279), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5009) );
  AND2_X4 U6489 ( .A1(n5007), .A2(n5006), .ZN(n5104) );
  NAND2_X1 U6490 ( .A1(n5104), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5008) );
  INV_X1 U6491 ( .A(n8567), .ZN(n8276) );
  XNOR2_X1 U6492 ( .A(n5013), .B(n5012), .ZN(n7647) );
  NAND2_X1 U6493 ( .A1(n7647), .A2(n5576), .ZN(n5018) );
  INV_X1 U6494 ( .A(n5318), .ZN(n5015) );
  INV_X1 U6495 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5014) );
  INV_X1 U6496 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5472) );
  OAI22_X1 U6497 ( .A1(n5320), .A2(n6624), .B1(n6354), .B2(n8433), .ZN(n5016)
         );
  INV_X1 U6498 ( .A(n5016), .ZN(n5017) );
  NAND2_X1 U6499 ( .A1(n5104), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5026) );
  INV_X1 U6500 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8365) );
  OR2_X1 U6501 ( .A1(n5463), .A2(n8365), .ZN(n5025) );
  INV_X1 U6502 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6503 ( .A1(n5326), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U6504 ( .A1(n5021), .A2(n5020), .ZN(n8168) );
  OR2_X1 U6505 ( .A1(n5510), .A2(n8168), .ZN(n5024) );
  INV_X1 U6506 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5022) );
  OR2_X1 U6507 ( .A1(n5581), .A2(n5022), .ZN(n5023) );
  NAND2_X1 U6508 ( .A1(n5104), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6509 ( .A1(n5067), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5029) );
  AND3_X1 U6510 ( .A1(n5030), .A2(n5029), .A3(n5028), .ZN(n5032) );
  NAND2_X1 U6511 ( .A1(n5032), .A2(n5031), .ZN(n6505) );
  INV_X1 U6512 ( .A(n6505), .ZN(n5042) );
  INV_X1 U6513 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5033) );
  XNOR2_X1 U6514 ( .A(n5035), .B(n5034), .ZN(n6159) );
  INV_X1 U6515 ( .A(n6159), .ZN(n5036) );
  NAND2_X1 U6516 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5037) );
  MUX2_X1 U6517 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5037), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5040) );
  INV_X1 U6518 ( .A(n5038), .ZN(n5039) );
  NAND2_X1 U6519 ( .A1(n5040), .A2(n5039), .ZN(n6344) );
  NAND2_X1 U6520 ( .A1(n6505), .A2(n9784), .ZN(n5482) );
  INV_X1 U6521 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6522 ( .A1(n5027), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6523 ( .A1(n5104), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6524 ( .A1(n5067), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6525 ( .A1(n6156), .A2(SI_0_), .ZN(n5048) );
  INV_X1 U6526 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6527 ( .A1(n5048), .A2(n5047), .ZN(n5050) );
  AND2_X1 U6528 ( .A1(n5050), .A2(n5049), .ZN(n8785) );
  MUX2_X1 U6529 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8785), .S(n5051), .Z(n6595) );
  NAND2_X1 U6530 ( .A1(n6970), .A2(n6971), .ZN(n5053) );
  OR2_X1 U6531 ( .A1(n6505), .A2(n5041), .ZN(n5052) );
  NAND2_X1 U6532 ( .A1(n5053), .A2(n5052), .ZN(n6843) );
  NAND2_X1 U6533 ( .A1(n4279), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6534 ( .A1(n5027), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6535 ( .A1(n5104), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6536 ( .A1(n5067), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5055) );
  NAND4_X2 U6537 ( .A1(n5058), .A2(n5057), .A3(n5056), .A4(n5055), .ZN(n8289)
         );
  XNOR2_X1 U6538 ( .A(n5059), .B(n5060), .ZN(n6180) );
  INV_X1 U6539 ( .A(n6180), .ZN(n5061) );
  NAND2_X1 U6540 ( .A1(n5076), .A2(n5061), .ZN(n5064) );
  OR2_X1 U6541 ( .A1(n5038), .A2(n5529), .ZN(n5062) );
  NAND2_X1 U6542 ( .A1(n5291), .A2(n9423), .ZN(n5063) );
  NAND2_X1 U6543 ( .A1(n8289), .A2(n9789), .ZN(n5613) );
  NAND2_X1 U6544 ( .A1(n6843), .A2(n6844), .ZN(n6598) );
  INV_X1 U6545 ( .A(n9789), .ZN(n6854) );
  OR2_X1 U6546 ( .A1(n8289), .A2(n6854), .ZN(n6599) );
  INV_X1 U6547 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5066) );
  INV_X1 U6548 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U6549 ( .A1(n5104), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5068) );
  OAI21_X1 U6550 ( .B1(n5581), .B2(n6361), .A(n5068), .ZN(n5069) );
  OAI21_X1 U6551 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5097), .ZN(n9756) );
  OR2_X1 U6552 ( .A1(n5099), .A2(n9756), .ZN(n5070) );
  NAND2_X1 U6553 ( .A1(n5071), .A2(n5070), .ZN(n5095) );
  NAND2_X1 U6554 ( .A1(n5073), .A2(n5072), .ZN(n5075) );
  XNOR2_X1 U6555 ( .A(n5075), .B(n5074), .ZN(n6300) );
  OR2_X1 U6556 ( .A1(n5078), .A2(n5529), .ZN(n5079) );
  XNOR2_X1 U6557 ( .A(n5079), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U6558 ( .A1(n5291), .A2(n6428), .ZN(n5080) );
  OAI211_X2 U6559 ( .C1(n6300), .C2(n5134), .A(n5081), .B(n5080), .ZN(n6533)
         );
  INV_X1 U6560 ( .A(n6533), .ZN(n9803) );
  NAND2_X1 U6561 ( .A1(n6917), .A2(n9803), .ZN(n5094) );
  NAND2_X1 U6562 ( .A1(n5104), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5086) );
  INV_X1 U6563 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6343) );
  OR2_X1 U6564 ( .A1(n5463), .A2(n6343), .ZN(n5085) );
  OR2_X1 U6565 ( .A1(n5099), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5084) );
  INV_X1 U6566 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6567 ( .A1(n5596), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U6568 ( .A(n5088), .B(n5087), .ZN(n6214) );
  NAND2_X1 U6569 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5089), .ZN(n5090) );
  XNOR2_X1 U6570 ( .A(n5090), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U6571 ( .A1(n5291), .A2(n8297), .ZN(n5091) );
  INV_X1 U6572 ( .A(n5093), .ZN(n9797) );
  NAND2_X1 U6573 ( .A1(n6847), .A2(n9797), .ZN(n9748) );
  NAND2_X1 U6574 ( .A1(n6847), .A2(n5093), .ZN(n9737) );
  INV_X1 U6575 ( .A(n6847), .ZN(n9743) );
  NAND2_X1 U6576 ( .A1(n9743), .A2(n9797), .ZN(n5627) );
  NAND2_X1 U6577 ( .A1(n9737), .A2(n5627), .ZN(n9746) );
  INV_X1 U6578 ( .A(n5094), .ZN(n5096) );
  NAND2_X1 U6579 ( .A1(n6917), .A2(n6533), .ZN(n5619) );
  NAND2_X1 U6580 ( .A1(n5619), .A2(n6912), .ZN(n9751) );
  OR2_X1 U6581 ( .A1(n5096), .A2(n9751), .ZN(n5107) );
  AND2_X1 U6582 ( .A1(n5108), .A2(n5107), .ZN(n6909) );
  INV_X1 U6583 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U6584 ( .A1(n5097), .A2(n8309), .ZN(n5098) );
  NAND2_X1 U6585 ( .A1(n5116), .A2(n5098), .ZN(n8130) );
  OR2_X1 U6586 ( .A1(n5099), .A2(n8130), .ZN(n5102) );
  NAND2_X1 U6587 ( .A1(n5067), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5100) );
  NAND3_X1 U6588 ( .A1(n5102), .A2(n5101), .A3(n5100), .ZN(n5103) );
  INV_X1 U6589 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5105) );
  OR2_X1 U6590 ( .A1(n5446), .A2(n5105), .ZN(n5106) );
  NAND2_X1 U6591 ( .A1(n5596), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5113) );
  INV_X1 U6592 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6593 ( .A1(n5078), .A2(n5162), .ZN(n5111) );
  NAND2_X1 U6594 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6595 ( .A(n5127), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U6596 ( .A1(n5291), .A2(n8311), .ZN(n5112) );
  OAI211_X2 U6597 ( .C1(n6475), .C2(n5134), .A(n5113), .B(n5112), .ZN(n9811)
         );
  NAND2_X1 U6598 ( .A1(n5067), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5122) );
  INV_X1 U6599 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6901) );
  OR2_X1 U6600 ( .A1(n5463), .A2(n6901), .ZN(n5121) );
  INV_X1 U6601 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6602 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6603 ( .A1(n5137), .A2(n5117), .ZN(n6902) );
  OR2_X1 U6604 ( .A1(n5510), .A2(n6902), .ZN(n5120) );
  INV_X1 U6605 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5118) );
  OR2_X1 U6606 ( .A1(n5446), .A2(n5118), .ZN(n5119) );
  NAND2_X1 U6607 ( .A1(n5124), .A2(n5123), .ZN(n5126) );
  XNOR2_X1 U6608 ( .A(n5126), .B(n5125), .ZN(n6541) );
  INV_X1 U6609 ( .A(n6541), .ZN(n5999) );
  NAND2_X1 U6610 ( .A1(n5596), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5133) );
  INV_X1 U6611 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U6612 ( .A1(n5127), .A2(n9937), .ZN(n5128) );
  NAND2_X1 U6613 ( .A1(n5128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6614 ( .A1(n5130), .A2(n5129), .ZN(n5144) );
  OR2_X1 U6615 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  AND2_X1 U6616 ( .A1(n5144), .A2(n5131), .ZN(n6437) );
  NAND2_X1 U6617 ( .A1(n5291), .A2(n6437), .ZN(n5132) );
  NAND2_X1 U6618 ( .A1(n6916), .A2(n6839), .ZN(n6752) );
  INV_X1 U6619 ( .A(n6916), .ZN(n8288) );
  INV_X1 U6620 ( .A(n6839), .ZN(n6903) );
  NAND2_X1 U6621 ( .A1(n8288), .A2(n6903), .ZN(n6751) );
  NAND2_X1 U6622 ( .A1(n6752), .A2(n6751), .ZN(n6834) );
  NAND2_X1 U6623 ( .A1(n6829), .A2(n6834), .ZN(n5136) );
  NAND2_X1 U6624 ( .A1(n8288), .A2(n6839), .ZN(n5135) );
  NAND2_X1 U6625 ( .A1(n5136), .A2(n5135), .ZN(n6750) );
  INV_X1 U6626 ( .A(n6750), .ZN(n5151) );
  NAND2_X1 U6627 ( .A1(n5067), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5143) );
  INV_X1 U6628 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6763) );
  OR2_X1 U6629 ( .A1(n5463), .A2(n6763), .ZN(n5142) );
  INV_X1 U6630 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U6631 ( .A1(n5137), .A2(n6463), .ZN(n5138) );
  NAND2_X1 U6632 ( .A1(n5153), .A2(n5138), .ZN(n6762) );
  OR2_X1 U6633 ( .A1(n5510), .A2(n6762), .ZN(n5141) );
  INV_X1 U6634 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5139) );
  OR2_X1 U6635 ( .A1(n5446), .A2(n5139), .ZN(n5140) );
  NAND2_X1 U6636 ( .A1(n5144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5145) );
  XNOR2_X1 U6637 ( .A(n5145), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6443) );
  INV_X1 U6638 ( .A(n6443), .ZN(n6474) );
  NAND2_X1 U6639 ( .A1(n6639), .A2(n5576), .ZN(n5149) );
  NAND2_X1 U6640 ( .A1(n5596), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6641 ( .A1(n7074), .A2(n6765), .ZN(n5630) );
  INV_X1 U6642 ( .A(n7074), .ZN(n8287) );
  INV_X1 U6643 ( .A(n6765), .ZN(n9820) );
  NAND2_X1 U6644 ( .A1(n5067), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5159) );
  INV_X1 U6645 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6446) );
  OR2_X1 U6646 ( .A1(n5463), .A2(n6446), .ZN(n5158) );
  NAND2_X1 U6647 ( .A1(n5153), .A2(n5152), .ZN(n5154) );
  NAND2_X1 U6648 ( .A1(n5170), .A2(n5154), .ZN(n6931) );
  OR2_X1 U6649 ( .A1(n5510), .A2(n6931), .ZN(n5157) );
  INV_X1 U6650 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5155) );
  OR2_X1 U6651 ( .A1(n5446), .A2(n5155), .ZN(n5156) );
  NAND2_X1 U6652 ( .A1(n6644), .A2(n5576), .ZN(n5167) );
  AND4_X1 U6653 ( .A1(n9937), .A2(n5162), .A3(n5129), .A4(n5161), .ZN(n5163)
         );
  NAND2_X1 U6654 ( .A1(n5078), .A2(n5163), .ZN(n5183) );
  NAND2_X1 U6655 ( .A1(n5183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6656 ( .A(n5160), .B(n5164), .ZN(n6458) );
  OAI22_X1 U6657 ( .A1(n5320), .A2(n9959), .B1(n6354), .B2(n6458), .ZN(n5165)
         );
  INV_X1 U6658 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6659 ( .A1(n7146), .A2(n7233), .ZN(n5634) );
  INV_X1 U6660 ( .A(n7233), .ZN(n7084) );
  NAND2_X1 U6661 ( .A1(n7084), .A2(n8286), .ZN(n5642) );
  NAND2_X1 U6662 ( .A1(n5634), .A2(n5642), .ZN(n7076) );
  NAND2_X1 U6663 ( .A1(n8286), .A2(n7233), .ZN(n5168) );
  NAND2_X1 U6664 ( .A1(n5104), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5175) );
  INV_X1 U6665 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7151) );
  OR2_X1 U6666 ( .A1(n5463), .A2(n7151), .ZN(n5174) );
  INV_X1 U6667 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6668 ( .A1(n5170), .A2(n5169), .ZN(n5171) );
  NAND2_X1 U6669 ( .A1(n5217), .A2(n5171), .ZN(n7150) );
  OR2_X1 U6670 ( .A1(n5510), .A2(n7150), .ZN(n5173) );
  INV_X1 U6671 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6685) );
  OR2_X1 U6672 ( .A1(n5581), .A2(n6685), .ZN(n5172) );
  NAND2_X1 U6673 ( .A1(n5178), .A2(n5177), .ZN(n5182) );
  AND2_X1 U6674 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  NAND2_X1 U6675 ( .A1(n6730), .A2(n5576), .ZN(n5187) );
  NOR2_X1 U6676 ( .A1(n5183), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6677 ( .A1(n5197), .A2(n5529), .ZN(n5184) );
  XNOR2_X1 U6678 ( .A(n5184), .B(n5196), .ZN(n6686) );
  OAI22_X1 U6679 ( .A1(n5320), .A2(n6026), .B1(n6354), .B2(n6686), .ZN(n5185)
         );
  INV_X1 U6680 ( .A(n5185), .ZN(n5186) );
  OR2_X1 U6681 ( .A1(n7332), .A2(n7157), .ZN(n5606) );
  NAND2_X1 U6682 ( .A1(n7157), .A2(n7332), .ZN(n5643) );
  INV_X1 U6683 ( .A(n7144), .ZN(n5188) );
  INV_X1 U6684 ( .A(n7332), .ZN(n8285) );
  OR2_X1 U6685 ( .A1(n8285), .A2(n7157), .ZN(n5189) );
  OR2_X1 U6686 ( .A1(n5191), .A2(n5190), .ZN(n5193) );
  NAND2_X1 U6687 ( .A1(n5193), .A2(n5192), .ZN(n5195) );
  NAND2_X1 U6688 ( .A1(n6862), .A2(n5576), .ZN(n5203) );
  NAND2_X1 U6689 ( .A1(n5197), .A2(n5196), .ZN(n5234) );
  NAND2_X1 U6690 ( .A1(n5234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5199) );
  INV_X1 U6691 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6692 ( .A1(n5199), .A2(n5198), .ZN(n5211) );
  OR2_X1 U6693 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6694 ( .A1(n5211), .A2(n5200), .ZN(n6690) );
  OAI22_X1 U6695 ( .A1(n5320), .A2(n9970), .B1(n6354), .B2(n6690), .ZN(n5201)
         );
  INV_X1 U6696 ( .A(n5201), .ZN(n5202) );
  NAND2_X1 U6697 ( .A1(n5203), .A2(n5202), .ZN(n7455) );
  NAND2_X1 U6698 ( .A1(n5067), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5208) );
  INV_X1 U6699 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6681) );
  OR2_X1 U6700 ( .A1(n5463), .A2(n6681), .ZN(n5207) );
  INV_X1 U6701 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6702 ( .A(n5217), .B(n5216), .ZN(n7341) );
  OR2_X1 U6703 ( .A1(n5510), .A2(n7341), .ZN(n5206) );
  INV_X1 U6704 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5204) );
  OR2_X1 U6705 ( .A1(n5446), .A2(n5204), .ZN(n5205) );
  OR2_X1 U6706 ( .A1(n7455), .A2(n7162), .ZN(n5607) );
  NAND2_X1 U6707 ( .A1(n7455), .A2(n7162), .ZN(n5644) );
  NAND2_X1 U6708 ( .A1(n5607), .A2(n5644), .ZN(n7334) );
  XNOR2_X1 U6709 ( .A(n5210), .B(n5209), .ZN(n6996) );
  NAND2_X1 U6710 ( .A1(n6996), .A2(n5576), .ZN(n5214) );
  NAND2_X1 U6711 ( .A1(n5211), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5212) );
  XNOR2_X1 U6712 ( .A(n5212), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6818) );
  AOI22_X1 U6713 ( .A1(n5596), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5291), .B2(
        n6818), .ZN(n5213) );
  NAND2_X1 U6714 ( .A1(n5067), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5223) );
  INV_X1 U6715 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7221) );
  OR2_X1 U6716 ( .A1(n5463), .A2(n7221), .ZN(n5222) );
  INV_X1 U6717 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5215) );
  OAI21_X1 U6718 ( .B1(n5217), .B2(n5216), .A(n5215), .ZN(n5218) );
  NAND2_X1 U6719 ( .A1(n5218), .A2(n5240), .ZN(n7220) );
  OR2_X1 U6720 ( .A1(n5510), .A2(n7220), .ZN(n5221) );
  INV_X1 U6721 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5219) );
  OR2_X1 U6722 ( .A1(n5446), .A2(n5219), .ZN(n5220) );
  INV_X1 U6723 ( .A(n7331), .ZN(n8283) );
  NAND2_X1 U6724 ( .A1(n7226), .A2(n8283), .ZN(n5227) );
  INV_X1 U6725 ( .A(n5227), .ZN(n5224) );
  OR2_X1 U6726 ( .A1(n7226), .A2(n7331), .ZN(n5647) );
  NAND2_X1 U6727 ( .A1(n7226), .A2(n7331), .ZN(n5650) );
  NAND2_X1 U6728 ( .A1(n5647), .A2(n5650), .ZN(n7230) );
  AND2_X1 U6729 ( .A1(n7334), .A2(n5226), .ZN(n5225) );
  NAND2_X1 U6730 ( .A1(n7227), .A2(n5225), .ZN(n5231) );
  INV_X1 U6731 ( .A(n5226), .ZN(n5229) );
  INV_X1 U6732 ( .A(n7162), .ZN(n8284) );
  NAND2_X1 U6733 ( .A1(n7455), .A2(n8284), .ZN(n7228) );
  AND2_X1 U6734 ( .A1(n7228), .A2(n5227), .ZN(n5228) );
  OR2_X1 U6735 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U6736 ( .A1(n5231), .A2(n5230), .ZN(n7208) );
  XNOR2_X1 U6737 ( .A(n5233), .B(n5232), .ZN(n7180) );
  NAND2_X1 U6738 ( .A1(n7180), .A2(n5576), .ZN(n5239) );
  OR3_X1 U6739 ( .A1(n5234), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6740 ( .A1(n5235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5236) );
  XNOR2_X1 U6741 ( .A(n5236), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6944) );
  INV_X1 U6742 ( .A(n6944), .ZN(n6828) );
  OAI22_X1 U6743 ( .A1(n5320), .A2(n9928), .B1(n6354), .B2(n6828), .ZN(n5237)
         );
  INV_X1 U6744 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6745 ( .A1(n5104), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5245) );
  INV_X1 U6746 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7212) );
  OR2_X1 U6747 ( .A1(n5463), .A2(n7212), .ZN(n5244) );
  INV_X1 U6748 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6819) );
  OR2_X1 U6749 ( .A1(n5581), .A2(n6819), .ZN(n5243) );
  INV_X1 U6750 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U6751 ( .A1(n5240), .A2(n7172), .ZN(n5241) );
  NAND2_X1 U6752 ( .A1(n5254), .A2(n5241), .ZN(n7211) );
  OR2_X1 U6753 ( .A1(n5510), .A2(n7211), .ZN(n5242) );
  NAND2_X1 U6754 ( .A1(n7210), .A2(n7304), .ZN(n5651) );
  INV_X1 U6755 ( .A(n7304), .ZN(n8282) );
  XNOR2_X1 U6756 ( .A(n5246), .B(n4869), .ZN(n7390) );
  NAND2_X1 U6757 ( .A1(n7390), .A2(n5576), .ZN(n5252) );
  NAND2_X1 U6758 ( .A1(n5248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6759 ( .A(n5249), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7094) );
  INV_X1 U6760 ( .A(n7094), .ZN(n7089) );
  OAI22_X1 U6761 ( .A1(n5320), .A2(n6117), .B1(n6354), .B2(n7089), .ZN(n5250)
         );
  INV_X1 U6762 ( .A(n5250), .ZN(n5251) );
  NAND2_X1 U6763 ( .A1(n5104), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5259) );
  INV_X1 U6764 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6765 ( .A1(n5581), .A2(n5253), .ZN(n5258) );
  INV_X1 U6766 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7323) );
  OR2_X1 U6767 ( .A1(n5463), .A2(n7323), .ZN(n5257) );
  NAND2_X1 U6768 ( .A1(n5254), .A2(n6947), .ZN(n5255) );
  NAND2_X1 U6769 ( .A1(n5267), .A2(n5255), .ZN(n7322) );
  OR2_X1 U6770 ( .A1(n5510), .A2(n7322), .ZN(n5256) );
  OR2_X1 U6771 ( .A1(n7503), .A2(n7431), .ZN(n5659) );
  NAND2_X1 U6772 ( .A1(n7503), .A2(n7431), .ZN(n5658) );
  XNOR2_X1 U6773 ( .A(n5261), .B(n5260), .ZN(n7557) );
  NAND2_X1 U6774 ( .A1(n7557), .A2(n5576), .ZN(n5266) );
  NAND2_X1 U6775 ( .A1(n5262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6776 ( .A(n5263), .B(n4740), .ZN(n7419) );
  OAI22_X1 U6777 ( .A1(n5320), .A2(n6126), .B1(n6354), .B2(n7419), .ZN(n5264)
         );
  INV_X1 U6778 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6779 ( .A1(n5104), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5272) );
  INV_X1 U6780 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7096) );
  OR2_X1 U6781 ( .A1(n5581), .A2(n7096), .ZN(n5271) );
  INV_X1 U6782 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7495) );
  OR2_X1 U6783 ( .A1(n5463), .A2(n7495), .ZN(n5270) );
  NAND2_X1 U6784 ( .A1(n5267), .A2(n7100), .ZN(n5268) );
  NAND2_X1 U6785 ( .A1(n5295), .A2(n5268), .ZN(n7494) );
  OR2_X1 U6786 ( .A1(n5510), .A2(n7494), .ZN(n5269) );
  NAND2_X1 U6787 ( .A1(n7493), .A2(n7446), .ZN(n5661) );
  INV_X1 U6788 ( .A(n7485), .ZN(n5273) );
  INV_X1 U6789 ( .A(n7431), .ZN(n8281) );
  NAND2_X1 U6790 ( .A1(n7503), .A2(n8281), .ZN(n7483) );
  AND2_X1 U6791 ( .A1(n5273), .A2(n7483), .ZN(n5274) );
  INV_X1 U6792 ( .A(n7446), .ZN(n8280) );
  NAND2_X1 U6793 ( .A1(n7567), .A2(n5576), .ZN(n5280) );
  OR2_X1 U6794 ( .A1(n5276), .A2(n5529), .ZN(n5277) );
  XNOR2_X1 U6795 ( .A(n5277), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7470) );
  INV_X1 U6796 ( .A(n7470), .ZN(n7464) );
  OAI22_X1 U6797 ( .A1(n5320), .A2(n6327), .B1(n6354), .B2(n7464), .ZN(n5278)
         );
  INV_X1 U6798 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6799 ( .A1(n4279), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5284) );
  INV_X1 U6800 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8713) );
  OR2_X1 U6801 ( .A1(n5581), .A2(n8713), .ZN(n5283) );
  INV_X1 U6802 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8262) );
  XNOR2_X1 U6803 ( .A(n5295), .B(n8262), .ZN(n7449) );
  OR2_X1 U6804 ( .A1(n5510), .A2(n7449), .ZN(n5282) );
  INV_X1 U6805 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8764) );
  OR2_X1 U6806 ( .A1(n5446), .A2(n8764), .ZN(n5281) );
  XNOR2_X1 U6807 ( .A(n7448), .B(n8622), .ZN(n7443) );
  NAND2_X1 U6808 ( .A1(n7441), .A2(n7443), .ZN(n7440) );
  INV_X1 U6809 ( .A(n8622), .ZN(n8279) );
  OR2_X1 U6810 ( .A1(n7448), .A2(n8279), .ZN(n5285) );
  XNOR2_X1 U6811 ( .A(n5287), .B(n5286), .ZN(n7590) );
  NAND2_X1 U6812 ( .A1(n7590), .A2(n5576), .ZN(n5293) );
  NAND2_X1 U6813 ( .A1(n5288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5289) );
  MUX2_X1 U6814 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5289), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5290) );
  AND2_X1 U6815 ( .A1(n5290), .A2(n4295), .ZN(n8340) );
  AOI22_X1 U6816 ( .A1(n5596), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5291), .B2(
        n8340), .ZN(n5292) );
  NAND2_X1 U6817 ( .A1(n5104), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5300) );
  INV_X1 U6818 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8708) );
  OR2_X1 U6819 ( .A1(n5581), .A2(n8708), .ZN(n5299) );
  INV_X1 U6820 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8631) );
  OR2_X1 U6821 ( .A1(n5463), .A2(n8631), .ZN(n5298) );
  INV_X1 U6822 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5294) );
  OAI21_X1 U6823 ( .B1(n5295), .B2(n8262), .A(n5294), .ZN(n5296) );
  NAND2_X1 U6824 ( .A1(n5309), .A2(n5296), .ZN(n8630) );
  OR2_X1 U6825 ( .A1(n5510), .A2(n8630), .ZN(n5297) );
  NAND2_X1 U6826 ( .A1(n8629), .A2(n8595), .ZN(n5605) );
  NAND2_X1 U6827 ( .A1(n5670), .A2(n5605), .ZN(n8617) );
  NAND2_X1 U6828 ( .A1(n8616), .A2(n8617), .ZN(n8615) );
  INV_X1 U6829 ( .A(n8595), .ZN(n8278) );
  NAND2_X1 U6830 ( .A1(n8629), .A2(n8278), .ZN(n5301) );
  NAND2_X1 U6831 ( .A1(n8615), .A2(n5301), .ZN(n8600) );
  XNOR2_X1 U6832 ( .A(n5303), .B(n5302), .ZN(n7608) );
  NAND2_X1 U6833 ( .A1(n7608), .A2(n5576), .ZN(n5308) );
  NAND2_X1 U6834 ( .A1(n4295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5304) );
  MUX2_X1 U6835 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5304), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5305) );
  NAND2_X1 U6836 ( .A1(n5305), .A2(n5318), .ZN(n8350) );
  OAI22_X1 U6837 ( .A1(n5320), .A2(n6342), .B1(n6354), .B2(n8350), .ZN(n5306)
         );
  INV_X1 U6838 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6839 ( .A1(n5104), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5314) );
  INV_X1 U6840 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8341) );
  OR2_X1 U6841 ( .A1(n5581), .A2(n8341), .ZN(n5313) );
  INV_X1 U6842 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8607) );
  OR2_X1 U6843 ( .A1(n5463), .A2(n8607), .ZN(n5312) );
  INV_X1 U6844 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U6845 ( .A1(n5309), .A2(n8338), .ZN(n5310) );
  NAND2_X1 U6846 ( .A1(n5324), .A2(n5310), .ZN(n8606) );
  OR2_X1 U6847 ( .A1(n5510), .A2(n8606), .ZN(n5311) );
  NAND2_X1 U6848 ( .A1(n8610), .A2(n8620), .ZN(n5673) );
  XNOR2_X1 U6849 ( .A(n5317), .B(n5316), .ZN(n7627) );
  NAND2_X1 U6850 ( .A1(n7627), .A2(n5576), .ZN(n5323) );
  INV_X1 U6851 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U6852 ( .A1(n5318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U6853 ( .A(n5319), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8368) );
  INV_X1 U6854 ( .A(n8368), .ZN(n8357) );
  OAI22_X1 U6855 ( .A1(n5320), .A2(n6522), .B1(n6354), .B2(n8357), .ZN(n5321)
         );
  INV_X1 U6856 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6857 ( .A1(n5104), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5330) );
  INV_X1 U6858 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8695) );
  OR2_X1 U6859 ( .A1(n5581), .A2(n8695), .ZN(n5329) );
  INV_X1 U6860 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8586) );
  OR2_X1 U6861 ( .A1(n5463), .A2(n8586), .ZN(n5328) );
  NAND2_X1 U6862 ( .A1(n5324), .A2(n8250), .ZN(n5325) );
  NAND2_X1 U6863 ( .A1(n5326), .A2(n5325), .ZN(n8585) );
  OR2_X1 U6864 ( .A1(n5510), .A2(n8585), .ZN(n5327) );
  NOR2_X1 U6865 ( .A1(n8754), .A2(n8596), .ZN(n5331) );
  INV_X1 U6866 ( .A(n8596), .ZN(n8277) );
  INV_X1 U6867 ( .A(n8249), .ZN(n8539) );
  NAND2_X1 U6868 ( .A1(n5333), .A2(n5332), .ZN(n8543) );
  NAND2_X1 U6869 ( .A1(n8681), .A2(n8567), .ZN(n5677) );
  INV_X1 U6870 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6938) );
  INV_X1 U6871 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7690) );
  MUX2_X1 U6872 ( .A(n6938), .B(n7690), .S(n6158), .Z(n5351) );
  XNOR2_X1 U6873 ( .A(n5351), .B(SI_21_), .ZN(n5350) );
  XNOR2_X1 U6874 ( .A(n5349), .B(n5350), .ZN(n7689) );
  NAND2_X1 U6875 ( .A1(n7689), .A2(n5576), .ZN(n5339) );
  NAND2_X1 U6876 ( .A1(n5596), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5338) );
  INV_X1 U6877 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5347) );
  INV_X1 U6878 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U6879 ( .A1(n5341), .A2(n8175), .ZN(n5342) );
  NAND2_X1 U6880 ( .A1(n5359), .A2(n5342), .ZN(n8528) );
  OR2_X1 U6881 ( .A1(n8528), .A2(n5510), .ZN(n5346) );
  NAND2_X1 U6882 ( .A1(n5067), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6883 ( .A1(n4279), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5343) );
  AND2_X1 U6884 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  OAI211_X1 U6885 ( .C1(n5446), .C2(n5347), .A(n5346), .B(n5345), .ZN(n8540)
         );
  NOR2_X1 U6886 ( .A1(n8676), .A2(n8540), .ZN(n5348) );
  INV_X1 U6887 ( .A(n8676), .ZN(n8532) );
  INV_X1 U6888 ( .A(n8540), .ZN(n8232) );
  INV_X1 U6889 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6890 ( .A1(n5352), .A2(SI_21_), .ZN(n5353) );
  INV_X1 U6891 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6988) );
  INV_X1 U6892 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7712) );
  INV_X1 U6893 ( .A(SI_22_), .ZN(n10008) );
  NAND2_X1 U6894 ( .A1(n5354), .A2(n10008), .ZN(n5364) );
  INV_X1 U6895 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6896 ( .A1(n5355), .A2(SI_22_), .ZN(n5356) );
  NAND2_X1 U6897 ( .A1(n5364), .A2(n5356), .ZN(n5365) );
  XNOR2_X1 U6898 ( .A(n5366), .B(n5365), .ZN(n7711) );
  NAND2_X1 U6899 ( .A1(n7711), .A2(n5576), .ZN(n5358) );
  NAND2_X1 U6900 ( .A1(n5596), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5357) );
  INV_X1 U6901 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U6902 ( .A1(n5359), .A2(n8230), .ZN(n5360) );
  AND2_X1 U6903 ( .A1(n5375), .A2(n5360), .ZN(n8512) );
  NAND2_X1 U6904 ( .A1(n8512), .A2(n5027), .ZN(n5363) );
  AOI22_X1 U6905 ( .A1(n5067), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n4279), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6906 ( .A1(n5104), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6907 ( .A1(n8511), .A2(n8526), .ZN(n5679) );
  INV_X1 U6908 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5368) );
  INV_X1 U6909 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7731) );
  MUX2_X1 U6910 ( .A(n5368), .B(n7731), .S(n5367), .Z(n5370) );
  INV_X1 U6911 ( .A(SI_23_), .ZN(n5369) );
  NAND2_X1 U6912 ( .A1(n5370), .A2(n5369), .ZN(n5382) );
  INV_X1 U6913 ( .A(n5370), .ZN(n5371) );
  NAND2_X1 U6914 ( .A1(n5371), .A2(SI_23_), .ZN(n5372) );
  NAND2_X1 U6915 ( .A1(n7730), .A2(n5576), .ZN(n5374) );
  NAND2_X1 U6916 ( .A1(n5596), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5373) );
  INV_X1 U6917 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U6918 ( .A1(n5375), .A2(n8155), .ZN(n5376) );
  NAND2_X1 U6919 ( .A1(n5388), .A2(n5376), .ZN(n8483) );
  AOI22_X1 U6920 ( .A1(n5067), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n4279), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6921 ( .A1(n5104), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5377) );
  OAI211_X1 U6922 ( .C1(n8483), .C2(n5510), .A(n5378), .B(n5377), .ZN(n8505)
         );
  INV_X1 U6923 ( .A(n8505), .ZN(n8235) );
  OR2_X1 U6924 ( .A1(n8665), .A2(n8235), .ZN(n5690) );
  NAND2_X1 U6925 ( .A1(n8665), .A2(n8235), .ZN(n5691) );
  NAND2_X1 U6926 ( .A1(n4649), .A2(n8487), .ZN(n8480) );
  INV_X1 U6927 ( .A(n8665), .ZN(n8486) );
  NAND2_X1 U6928 ( .A1(n8480), .A2(n5379), .ZN(n8471) );
  INV_X1 U6929 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7177) );
  INV_X1 U6930 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10002) );
  XNOR2_X1 U6931 ( .A(n5394), .B(SI_24_), .ZN(n5393) );
  XNOR2_X1 U6932 ( .A(n5398), .B(n5393), .ZN(n7543) );
  NAND2_X1 U6933 ( .A1(n7543), .A2(n5576), .ZN(n5385) );
  NAND2_X1 U6934 ( .A1(n5596), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5384) );
  INV_X1 U6935 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6936 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  AND2_X1 U6937 ( .A1(n5406), .A2(n5389), .ZN(n8474) );
  INV_X1 U6938 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U6939 ( .A1(n4279), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6940 ( .A1(n5067), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5390) );
  OAI211_X1 U6941 ( .C1(n5446), .C2(n8740), .A(n5391), .B(n5390), .ZN(n5392)
         );
  AOI21_X1 U6942 ( .B1(n8474), .B2(n5027), .A(n5392), .ZN(n8213) );
  NAND2_X1 U6943 ( .A1(n8473), .A2(n8213), .ZN(n5695) );
  INV_X1 U6944 ( .A(n8213), .ZN(n8492) );
  OAI22_X1 U6945 ( .A1(n8471), .A2(n8470), .B1(n8473), .B2(n8492), .ZN(n8453)
         );
  INV_X1 U6946 ( .A(n5393), .ZN(n5397) );
  INV_X1 U6947 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6948 ( .A1(n5395), .A2(SI_24_), .ZN(n5396) );
  INV_X1 U6949 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10016) );
  INV_X1 U6950 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7753) );
  MUX2_X1 U6951 ( .A(n10016), .B(n7753), .S(n6158), .Z(n5400) );
  INV_X1 U6952 ( .A(SI_25_), .ZN(n5399) );
  NAND2_X1 U6953 ( .A1(n5400), .A2(n5399), .ZN(n5414) );
  INV_X1 U6954 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6955 ( .A1(n5401), .A2(SI_25_), .ZN(n5402) );
  NAND2_X1 U6956 ( .A1(n5414), .A2(n5402), .ZN(n5415) );
  NAND2_X1 U6957 ( .A1(n7752), .A2(n5576), .ZN(n5404) );
  NAND2_X1 U6958 ( .A1(n5596), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5403) );
  INV_X1 U6959 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U6960 ( .A1(n5406), .A2(n9997), .ZN(n5407) );
  NAND2_X1 U6961 ( .A1(n5424), .A2(n5407), .ZN(n8457) );
  OR2_X1 U6962 ( .A1(n8457), .A2(n5510), .ZN(n5412) );
  INV_X1 U6963 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U6964 ( .A1(n5067), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6965 ( .A1(n4279), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5408) );
  OAI211_X1 U6966 ( .C1(n8736), .C2(n5446), .A(n5409), .B(n5408), .ZN(n5410)
         );
  INV_X1 U6967 ( .A(n5410), .ZN(n5411) );
  NAND2_X1 U6968 ( .A1(n8456), .A2(n8436), .ZN(n5700) );
  NAND2_X1 U6969 ( .A1(n8453), .A2(n8452), .ZN(n8451) );
  NAND2_X1 U6970 ( .A1(n8451), .A2(n5413), .ZN(n8442) );
  INV_X1 U6971 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5417) );
  INV_X1 U6972 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7772) );
  MUX2_X1 U6973 ( .A(n5417), .B(n7772), .S(n6158), .Z(n5418) );
  NAND2_X1 U6974 ( .A1(n5418), .A2(n9925), .ZN(n5431) );
  INV_X1 U6975 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6976 ( .A1(n5419), .A2(SI_26_), .ZN(n5420) );
  AND2_X1 U6977 ( .A1(n5431), .A2(n5420), .ZN(n5430) );
  NAND2_X1 U6978 ( .A1(n7771), .A2(n5576), .ZN(n5422) );
  NAND2_X1 U6979 ( .A1(n5596), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5421) );
  INV_X1 U6980 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6981 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  INV_X1 U6982 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U6983 ( .A1(n5067), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6984 ( .A1(n4279), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5426) );
  OAI211_X1 U6985 ( .C1(n8732), .C2(n5446), .A(n5427), .B(n5426), .ZN(n5428)
         );
  NAND2_X1 U6986 ( .A1(n8443), .A2(n8184), .ZN(n5702) );
  NAND2_X1 U6987 ( .A1(n8442), .A2(n8441), .ZN(n8440) );
  INV_X1 U6988 ( .A(n8184), .ZN(n8274) );
  NAND2_X1 U6989 ( .A1(n8734), .A2(n8184), .ZN(n5429) );
  NAND2_X1 U6990 ( .A1(n8440), .A2(n5429), .ZN(n8422) );
  INV_X1 U6991 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5433) );
  INV_X1 U6992 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7790) );
  MUX2_X1 U6993 ( .A(n5433), .B(n7790), .S(n6158), .Z(n5435) );
  INV_X1 U6994 ( .A(SI_27_), .ZN(n5434) );
  NAND2_X1 U6995 ( .A1(n5435), .A2(n5434), .ZN(n5453) );
  INV_X1 U6996 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6997 ( .A1(n5436), .A2(SI_27_), .ZN(n5437) );
  AND2_X1 U6998 ( .A1(n5453), .A2(n5437), .ZN(n5451) );
  NAND2_X1 U6999 ( .A1(n5596), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5438) );
  INV_X1 U7000 ( .A(n5442), .ZN(n5440) );
  NAND2_X1 U7001 ( .A1(n5440), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5459) );
  INV_X1 U7002 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7003 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  NAND2_X1 U7004 ( .A1(n5459), .A2(n5443), .ZN(n8425) );
  INV_X1 U7005 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U7006 ( .A1(n5067), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7007 ( .A1(n4279), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5444) );
  OAI211_X1 U7008 ( .C1(n8728), .C2(n5446), .A(n5445), .B(n5444), .ZN(n5447)
         );
  INV_X1 U7009 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U7010 ( .A1(n8422), .A2(n8421), .ZN(n8420) );
  INV_X1 U7011 ( .A(n8437), .ZN(n8273) );
  NAND2_X1 U7012 ( .A1(n8420), .A2(n5450), .ZN(n5467) );
  MUX2_X1 U7013 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6156), .Z(n5563) );
  INV_X1 U7014 ( .A(SI_28_), .ZN(n5564) );
  XNOR2_X1 U7015 ( .A(n5563), .B(n5564), .ZN(n5561) );
  NAND2_X1 U7016 ( .A1(n7805), .A2(n5576), .ZN(n5456) );
  NAND2_X1 U7017 ( .A1(n5596), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5455) );
  INV_X1 U7018 ( .A(n5459), .ZN(n5457) );
  NAND2_X1 U7019 ( .A1(n5457), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8396) );
  INV_X1 U7020 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7021 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  NAND2_X1 U7022 ( .A1(n8396), .A2(n5460), .ZN(n8408) );
  INV_X1 U7023 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U7024 ( .A1(n5067), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7025 ( .A1(n5104), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5461) );
  OAI211_X1 U7026 ( .C1(n5463), .C2(n8407), .A(n5462), .B(n5461), .ZN(n5464)
         );
  INV_X1 U7027 ( .A(n5464), .ZN(n5465) );
  NAND2_X1 U7028 ( .A1(n7532), .A2(n7526), .ZN(n5708) );
  NAND2_X1 U7029 ( .A1(n5467), .A2(n5743), .ZN(n5885) );
  INV_X1 U7030 ( .A(n5467), .ZN(n5469) );
  INV_X1 U7031 ( .A(n5743), .ZN(n5468) );
  NAND2_X1 U7032 ( .A1(n5885), .A2(n5470), .ZN(n8405) );
  INV_X1 U7033 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5475) );
  XNOR2_X1 U7034 ( .A(n5535), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7035 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  NAND2_X1 U7036 ( .A1(n5474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5476) );
  XNOR2_X1 U7037 ( .A(n5476), .B(n5475), .ZN(n6857) );
  NAND2_X1 U7038 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7039 ( .A1(n6857), .A2(n5480), .ZN(n6590) );
  XNOR2_X1 U7040 ( .A(n5508), .B(n6590), .ZN(n5479) );
  NAND2_X1 U7041 ( .A1(n5479), .A2(n8433), .ZN(n8626) );
  INV_X1 U7042 ( .A(n6857), .ZN(n5747) );
  OR3_X1 U7043 ( .A1(n5508), .A2(n5747), .A3(n8433), .ZN(n8704) );
  NAND2_X1 U7044 ( .A1(n8626), .A2(n8704), .ZN(n9838) );
  NAND2_X1 U7045 ( .A1(n9781), .A2(n9789), .ZN(n6851) );
  NOR2_X1 U7046 ( .A1(n9752), .A2(n6533), .ZN(n6919) );
  INV_X1 U7047 ( .A(n9811), .ZN(n8131) );
  NAND2_X1 U7048 ( .A1(n6920), .A2(n6903), .ZN(n6831) );
  INV_X1 U7049 ( .A(n7157), .ZN(n9825) );
  INV_X1 U7050 ( .A(n7455), .ZN(n7344) );
  NAND2_X1 U7051 ( .A1(n7338), .A2(n7344), .ZN(n7222) );
  INV_X1 U7052 ( .A(n7493), .ZN(n8771) );
  NOR2_X2 U7053 ( .A1(n8628), .A2(n8629), .ZN(n8627) );
  INV_X1 U7054 ( .A(n8511), .ZN(n8747) );
  OR2_X2 U7055 ( .A1(n8508), .A2(n8665), .ZN(n8481) );
  INV_X1 U7056 ( .A(n5508), .ZN(n6986) );
  AOI211_X1 U7057 ( .C1(n7532), .C2(n8423), .A(n9826), .B(n5895), .ZN(n8411)
         );
  INV_X1 U7058 ( .A(n6970), .ZN(n5730) );
  NAND2_X1 U7059 ( .A1(n6570), .A2(n6595), .ZN(n6972) );
  INV_X1 U7060 ( .A(n6595), .ZN(n9776) );
  NAND2_X1 U7061 ( .A1(n5481), .A2(n9776), .ZN(n5729) );
  NAND2_X1 U7062 ( .A1(n5482), .A2(n5729), .ZN(n5610) );
  NAND2_X1 U7063 ( .A1(n5610), .A2(n5483), .ZN(n5615) );
  NAND2_X1 U7064 ( .A1(n9741), .A2(n8131), .ZN(n5731) );
  AND2_X1 U7065 ( .A1(n6912), .A2(n5731), .ZN(n5620) );
  INV_X2 U7066 ( .A(n9746), .ZN(n6910) );
  NAND2_X1 U7067 ( .A1(n6602), .A2(n5484), .ZN(n5487) );
  INV_X1 U7068 ( .A(n5620), .ZN(n5485) );
  NAND2_X1 U7069 ( .A1(n5619), .A2(n9737), .ZN(n5623) );
  INV_X1 U7070 ( .A(n5623), .ZN(n6911) );
  AND2_X1 U7071 ( .A1(n6751), .A2(n5631), .ZN(n5488) );
  NAND2_X1 U7072 ( .A1(n6835), .A2(n5488), .ZN(n5492) );
  INV_X1 U7073 ( .A(n5631), .ZN(n5490) );
  AND2_X1 U7074 ( .A1(n6752), .A2(n5630), .ZN(n5489) );
  INV_X1 U7075 ( .A(n7076), .ZN(n7072) );
  NAND2_X1 U7076 ( .A1(n7073), .A2(n7072), .ZN(n5493) );
  NAND2_X1 U7077 ( .A1(n5493), .A2(n5634), .ZN(n7145) );
  NAND2_X1 U7078 ( .A1(n7145), .A2(n7144), .ZN(n5494) );
  INV_X1 U7079 ( .A(n5650), .ZN(n5495) );
  INV_X1 U7080 ( .A(n7318), .ZN(n7312) );
  NAND2_X1 U7081 ( .A1(n7487), .A2(n7442), .ZN(n5496) );
  INV_X1 U7082 ( .A(n7443), .ZN(n5663) );
  INV_X1 U7083 ( .A(n7448), .ZN(n8766) );
  NAND2_X1 U7084 ( .A1(n8766), .A2(n8279), .ZN(n5497) );
  NAND2_X1 U7085 ( .A1(n8594), .A2(n8599), .ZN(n8557) );
  OR2_X1 U7086 ( .A1(n8590), .A2(n8596), .ZN(n5728) );
  AND2_X1 U7087 ( .A1(n8577), .A2(n5728), .ZN(n8558) );
  OR2_X1 U7088 ( .A1(n8688), .A2(n8249), .ZN(n5676) );
  NAND2_X1 U7089 ( .A1(n8688), .A2(n8249), .ZN(n8537) );
  NAND2_X1 U7090 ( .A1(n5676), .A2(n8537), .ZN(n8563) );
  INV_X1 U7091 ( .A(n8563), .ZN(n8555) );
  AND2_X1 U7092 ( .A1(n8558), .A2(n8555), .ZN(n5498) );
  NAND2_X1 U7093 ( .A1(n8557), .A2(n5498), .ZN(n8536) );
  INV_X1 U7094 ( .A(n8542), .ZN(n5499) );
  INV_X1 U7095 ( .A(n8537), .ZN(n5680) );
  NOR2_X1 U7096 ( .A1(n5499), .A2(n5680), .ZN(n5500) );
  NAND2_X1 U7097 ( .A1(n8590), .A2(n8596), .ZN(n8559) );
  OR2_X1 U7098 ( .A1(n8563), .A2(n8559), .ZN(n8535) );
  AND2_X1 U7099 ( .A1(n5500), .A2(n8535), .ZN(n5501) );
  OR2_X1 U7100 ( .A1(n8676), .A2(n8232), .ZN(n5684) );
  NAND2_X1 U7101 ( .A1(n8676), .A2(n8232), .ZN(n8500) );
  NAND2_X1 U7102 ( .A1(n5684), .A2(n8500), .ZN(n8523) );
  INV_X1 U7103 ( .A(n8523), .ZN(n5502) );
  AND2_X1 U7104 ( .A1(n8519), .A2(n5502), .ZN(n5503) );
  INV_X1 U7105 ( .A(n8498), .ZN(n8501) );
  INV_X1 U7106 ( .A(n8500), .ZN(n5504) );
  NOR2_X1 U7107 ( .A1(n8501), .A2(n5504), .ZN(n5505) );
  INV_X1 U7108 ( .A(n5685), .ZN(n8488) );
  NOR2_X1 U7109 ( .A1(n8487), .A2(n8488), .ZN(n5506) );
  INV_X1 U7110 ( .A(n8470), .ZN(n8467) );
  NAND2_X1 U7111 ( .A1(n8464), .A2(n5694), .ZN(n8447) );
  INV_X1 U7112 ( .A(n8452), .ZN(n5741) );
  NAND2_X1 U7113 ( .A1(n8447), .A2(n5741), .ZN(n5507) );
  NAND2_X1 U7114 ( .A1(n5507), .A2(n5699), .ZN(n8434) );
  NOR2_X1 U7115 ( .A1(n8424), .A2(n8437), .ZN(n5706) );
  INV_X1 U7116 ( .A(n8433), .ZN(n8375) );
  NAND2_X1 U7117 ( .A1(n5508), .A2(n8375), .ZN(n5757) );
  NAND2_X1 U7118 ( .A1(n5747), .A2(n5480), .ZN(n5603) );
  NAND2_X1 U7119 ( .A1(n5757), .A2(n5603), .ZN(n9745) );
  INV_X1 U7120 ( .A(n9745), .ZN(n8566) );
  AOI211_X1 U7121 ( .C1(n5509), .C2(n5743), .A(n8566), .B(n5560), .ZN(n5516)
         );
  OR2_X1 U7122 ( .A1(n8396), .A2(n5510), .ZN(n5515) );
  INV_X1 U7123 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7124 ( .A1(n4279), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7125 ( .A1(n5067), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5511) );
  OAI211_X1 U7126 ( .C1(n5897), .C2(n5446), .A(n5512), .B(n5511), .ZN(n5513)
         );
  INV_X1 U7127 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7128 ( .A1(n6353), .A2(n6359), .ZN(n8619) );
  INV_X1 U7129 ( .A(n6359), .ZN(n6350) );
  OAI22_X1 U7130 ( .A1(n6378), .A2(n8619), .B1(n8437), .B2(n8621), .ZN(n7515)
         );
  OR2_X1 U7131 ( .A1(n5516), .A2(n7515), .ZN(n8404) );
  NOR4_X1 U7132 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5520) );
  NOR4_X1 U7133 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5519) );
  NOR4_X1 U7134 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5518) );
  NOR4_X1 U7135 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5517) );
  NAND4_X1 U7136 ( .A1(n5520), .A2(n5519), .A3(n5518), .A4(n5517), .ZN(n5544)
         );
  NOR2_X1 U7137 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n5524) );
  NOR4_X1 U7138 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5523) );
  NOR4_X1 U7139 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5522) );
  NOR4_X1 U7140 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5521) );
  NAND4_X1 U7141 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n5543)
         );
  NAND2_X1 U7142 ( .A1(n5525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5526) );
  MUX2_X1 U7143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5526), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5528) );
  NAND2_X1 U7144 ( .A1(n5528), .A2(n5527), .ZN(n5547) );
  INV_X1 U7145 ( .A(n5547), .ZN(n7310) );
  OR2_X1 U7146 ( .A1(n5530), .A2(n5529), .ZN(n5532) );
  MUX2_X1 U7147 ( .A(n5532), .B(P2_IR_REG_31__SCAN_IN), .S(n5531), .Z(n5533)
         );
  NAND2_X1 U7148 ( .A1(n5533), .A2(n5525), .ZN(n7375) );
  INV_X1 U7149 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7150 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  NAND2_X1 U7151 ( .A1(n5536), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5545) );
  INV_X1 U7152 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7153 ( .A1(n5545), .A2(n5537), .ZN(n5538) );
  NAND2_X1 U7154 ( .A1(n5538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5540) );
  INV_X1 U7155 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5539) );
  XNOR2_X1 U7156 ( .A(n7179), .B(P2_B_REG_SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7157 ( .A1(n7375), .A2(n5541), .ZN(n5542) );
  OAI21_X1 U7158 ( .B1(n5544), .B2(n5543), .A(n9768), .ZN(n5862) );
  XNOR2_X1 U7159 ( .A(n5545), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5872) );
  AND2_X1 U7160 ( .A1(n6353), .A2(n5878), .ZN(n5873) );
  NOR2_X1 U7161 ( .A1(n9767), .A2(n5873), .ZN(n6587) );
  NAND3_X1 U7162 ( .A1(n5862), .A2(n6587), .A3(n5870), .ZN(n5546) );
  INV_X1 U7163 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9773) );
  AND2_X1 U7164 ( .A1(n7375), .A2(n5547), .ZN(n9775) );
  AOI21_X1 U7165 ( .B1(n9768), .B2(n9773), .A(n9775), .ZN(n5863) );
  AND2_X1 U7166 ( .A1(n7179), .A2(n5547), .ZN(n9770) );
  INV_X1 U7167 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9771) );
  AND2_X2 U7168 ( .A1(n5554), .A2(n5864), .ZN(n9855) );
  MUX2_X1 U7169 ( .A(n5549), .B(n5555), .S(n9855), .Z(n5553) );
  INV_X1 U7170 ( .A(n5878), .ZN(n5550) );
  NAND2_X1 U7171 ( .A1(n7532), .A2(n5551), .ZN(n5552) );
  NAND2_X1 U7172 ( .A1(n5553), .A2(n5552), .ZN(P2_U3548) );
  INV_X1 U7173 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5556) );
  INV_X1 U7174 ( .A(n5864), .ZN(n6589) );
  MUX2_X1 U7175 ( .A(n5556), .B(n5555), .S(n9840), .Z(n5558) );
  NAND2_X1 U7176 ( .A1(n7532), .A2(n6840), .ZN(n5557) );
  NAND2_X1 U7177 ( .A1(n5558), .A2(n5557), .ZN(P2_U3516) );
  INV_X1 U7178 ( .A(n5709), .ZN(n5559) );
  INV_X1 U7179 ( .A(n5887), .ZN(n5571) );
  INV_X1 U7180 ( .A(n5563), .ZN(n5565) );
  NAND2_X1 U7181 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  INV_X1 U7182 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7956) );
  INV_X1 U7183 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5567) );
  MUX2_X1 U7184 ( .A(n7956), .B(n5567), .S(n6156), .Z(n5572) );
  XNOR2_X1 U7185 ( .A(n5572), .B(SI_29_), .ZN(n5568) );
  NAND2_X1 U7186 ( .A1(n7955), .A2(n5576), .ZN(n5570) );
  NAND2_X1 U7187 ( .A1(n5596), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5569) );
  INV_X1 U7188 ( .A(n5727), .ZN(n5710) );
  NAND2_X1 U7189 ( .A1(n8400), .A2(n6378), .ZN(n5726) );
  INV_X1 U7190 ( .A(n5585), .ZN(n5586) );
  INV_X1 U7191 ( .A(n5572), .ZN(n5573) );
  NOR2_X1 U7192 ( .A1(n5573), .A2(SI_29_), .ZN(n5574) );
  MUX2_X1 U7193 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6156), .Z(n5589) );
  NAND2_X1 U7194 ( .A1(n7845), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7195 ( .A1(n5596), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5577) );
  INV_X1 U7196 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U7197 ( .A1(n4279), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7198 ( .A1(n5104), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U7199 ( .C1(n5581), .C2(n9911), .A(n5580), .B(n5579), .ZN(n8271)
         );
  NAND2_X1 U7200 ( .A1(n8726), .A2(n8271), .ZN(n5716) );
  NAND2_X1 U7201 ( .A1(n5067), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7202 ( .A1(n4279), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7203 ( .A1(n5104), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5582) );
  AND3_X1 U7204 ( .A1(n5584), .A2(n5583), .A3(n5582), .ZN(n8385) );
  INV_X1 U7205 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7206 ( .A1(n5588), .A2(SI_30_), .ZN(n5592) );
  NAND2_X1 U7207 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7208 ( .A1(n5592), .A2(n5591), .ZN(n5595) );
  MUX2_X1 U7209 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6156), .Z(n5593) );
  XNOR2_X1 U7210 ( .A(n5593), .B(SI_31_), .ZN(n5594) );
  NAND2_X1 U7211 ( .A1(n8772), .A2(n5576), .ZN(n5598) );
  NAND2_X1 U7212 ( .A1(n5596), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5597) );
  OR2_X1 U7213 ( .A1(n8386), .A2(n8385), .ZN(n5601) );
  INV_X1 U7214 ( .A(n8726), .ZN(n5600) );
  INV_X1 U7215 ( .A(n8271), .ZN(n5599) );
  NAND2_X1 U7216 ( .A1(n5600), .A2(n5599), .ZN(n5712) );
  NAND2_X1 U7217 ( .A1(n8386), .A2(n8385), .ZN(n5715) );
  AOI21_X1 U7218 ( .B1(n6594), .B2(n5603), .A(n5602), .ZN(n5752) );
  INV_X1 U7219 ( .A(n5698), .ZN(n5704) );
  NAND2_X1 U7220 ( .A1(n8375), .A2(n5480), .ZN(n5604) );
  INV_X1 U7221 ( .A(n5605), .ZN(n5674) );
  AND2_X1 U7222 ( .A1(n5607), .A2(n5606), .ZN(n5639) );
  INV_X1 U7223 ( .A(n5639), .ZN(n5608) );
  NAND2_X1 U7224 ( .A1(n5608), .A2(n5644), .ZN(n5609) );
  NAND2_X1 U7225 ( .A1(n5647), .A2(n5609), .ZN(n5638) );
  OAI21_X1 U7226 ( .B1(n5610), .B2(n6936), .A(n6845), .ZN(n5612) );
  INV_X1 U7227 ( .A(n5611), .ZN(n5614) );
  AOI21_X1 U7228 ( .B1(n5612), .B2(n5613), .A(n5614), .ZN(n5618) );
  OAI21_X1 U7229 ( .B1(n5615), .B2(n5614), .A(n5613), .ZN(n5616) );
  INV_X1 U7230 ( .A(n5616), .ZN(n5617) );
  INV_X1 U7231 ( .A(n5721), .ZN(n5719) );
  MUX2_X1 U7232 ( .A(n5618), .B(n5617), .S(n5719), .Z(n5625) );
  AND2_X1 U7233 ( .A1(n5619), .A2(n5732), .ZN(n5621) );
  MUX2_X1 U7234 ( .A(n5621), .B(n5620), .S(n5721), .Z(n5626) );
  NAND2_X1 U7235 ( .A1(n6752), .A2(n5732), .ZN(n5622) );
  AOI21_X1 U7236 ( .B1(n5626), .B2(n5623), .A(n5622), .ZN(n5624) );
  INV_X1 U7237 ( .A(n5626), .ZN(n5629) );
  AND2_X1 U7238 ( .A1(n5627), .A2(n6912), .ZN(n5628) );
  OAI21_X1 U7239 ( .B1(n6752), .B2(n5721), .A(n6754), .ZN(n5633) );
  MUX2_X1 U7240 ( .A(n5631), .B(n5630), .S(n5721), .Z(n5632) );
  INV_X1 U7241 ( .A(n5634), .ZN(n5635) );
  OAI21_X1 U7242 ( .B1(n5640), .B2(n5635), .A(n5639), .ZN(n5636) );
  NAND3_X1 U7243 ( .A1(n5636), .A2(n5650), .A3(n5644), .ZN(n5637) );
  MUX2_X1 U7244 ( .A(n5638), .B(n5637), .S(n5719), .Z(n5657) );
  NAND2_X1 U7245 ( .A1(n5640), .A2(n5639), .ZN(n5641) );
  OAI21_X1 U7246 ( .B1(n5719), .B2(n5642), .A(n5641), .ZN(n5645) );
  NAND3_X1 U7247 ( .A1(n5645), .A2(n5644), .A3(n5643), .ZN(n5646) );
  INV_X1 U7248 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7249 ( .A1(n5651), .A2(n5648), .ZN(n5649) );
  AND2_X1 U7250 ( .A1(n5649), .A2(n5652), .ZN(n5655) );
  NAND2_X1 U7251 ( .A1(n5651), .A2(n5650), .ZN(n5653) );
  NAND2_X1 U7252 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  MUX2_X1 U7253 ( .A(n5655), .B(n5654), .S(n5721), .Z(n5656) );
  MUX2_X1 U7254 ( .A(n5659), .B(n5658), .S(n5721), .Z(n5660) );
  MUX2_X1 U7255 ( .A(n5661), .B(n7442), .S(n5721), .Z(n5662) );
  NAND3_X1 U7256 ( .A1(n5664), .A2(n5663), .A3(n5662), .ZN(n5669) );
  AND2_X1 U7257 ( .A1(n7448), .A2(n5721), .ZN(n5666) );
  NOR2_X1 U7258 ( .A1(n7448), .A2(n5721), .ZN(n5665) );
  MUX2_X1 U7259 ( .A(n5666), .B(n5665), .S(n8279), .Z(n5667) );
  INV_X1 U7260 ( .A(n5667), .ZN(n5668) );
  AOI21_X1 U7261 ( .B1(n5669), .B2(n5668), .A(n8617), .ZN(n5672) );
  OAI21_X1 U7262 ( .B1(n5670), .B2(n5721), .A(n8599), .ZN(n5671) );
  INV_X1 U7263 ( .A(n8559), .ZN(n5675) );
  NAND2_X1 U7264 ( .A1(n8519), .A2(n5676), .ZN(n5682) );
  MUX2_X1 U7265 ( .A(n5679), .B(n5678), .S(n5721), .Z(n5689) );
  INV_X1 U7266 ( .A(n8487), .ZN(n5688) );
  AOI21_X1 U7267 ( .B1(n5681), .B2(n5728), .A(n5680), .ZN(n5683) );
  OAI21_X1 U7268 ( .B1(n5683), .B2(n5682), .A(n4327), .ZN(n5686) );
  NAND4_X1 U7269 ( .A1(n5686), .A2(n5719), .A3(n5685), .A4(n5684), .ZN(n5687)
         );
  NAND2_X1 U7270 ( .A1(n8470), .A2(n5690), .ZN(n5693) );
  NAND2_X1 U7271 ( .A1(n5695), .A2(n5691), .ZN(n5692) );
  MUX2_X1 U7272 ( .A(n5693), .B(n5692), .S(n5721), .Z(n5697) );
  MUX2_X1 U7273 ( .A(n5695), .B(n5694), .S(n5721), .Z(n5696) );
  NAND2_X1 U7274 ( .A1(n5702), .A2(n5700), .ZN(n5701) );
  OAI21_X1 U7275 ( .B1(n8730), .B2(n8273), .A(n5708), .ZN(n5705) );
  MUX2_X1 U7276 ( .A(n5706), .B(n5705), .S(n5721), .Z(n5707) );
  NOR2_X1 U7277 ( .A1(n5710), .A2(n5719), .ZN(n5711) );
  AOI21_X1 U7278 ( .B1(n5719), .B2(n5726), .A(n5711), .ZN(n5713) );
  OAI211_X1 U7279 ( .C1(n5714), .C2(n5713), .A(n5716), .B(n5712), .ZN(n5724)
         );
  INV_X1 U7280 ( .A(n5715), .ZN(n5718) );
  INV_X1 U7281 ( .A(n5716), .ZN(n5717) );
  NOR2_X1 U7282 ( .A1(n5718), .A2(n5717), .ZN(n5745) );
  MUX2_X1 U7283 ( .A(n4301), .B(n5745), .S(n5721), .Z(n5723) );
  INV_X1 U7284 ( .A(n8385), .ZN(n6037) );
  MUX2_X1 U7285 ( .A(n5719), .B(n6037), .S(n8386), .Z(n5720) );
  AOI21_X1 U7286 ( .B1(n8385), .B2(n5721), .A(n5720), .ZN(n5722) );
  INV_X1 U7287 ( .A(n8599), .ZN(n8593) );
  AND2_X1 U7288 ( .A1(n6972), .A2(n5729), .ZN(n9778) );
  NAND4_X1 U7289 ( .A1(n5730), .A2(n5747), .A3(n9778), .A4(n6910), .ZN(n5733)
         );
  NAND2_X1 U7290 ( .A1(n5732), .A2(n5731), .ZN(n6914) );
  NOR4_X1 U7291 ( .A1(n5733), .A2(n9751), .A3(n6844), .A4(n6914), .ZN(n5734)
         );
  INV_X1 U7292 ( .A(n6834), .ZN(n6830) );
  NAND4_X1 U7293 ( .A1(n5734), .A2(n7072), .A3(n6754), .A4(n6830), .ZN(n5735)
         );
  NOR4_X1 U7294 ( .A1(n5735), .A2(n7230), .A3(n7334), .A4(n5188), .ZN(n5736)
         );
  NAND4_X1 U7295 ( .A1(n7485), .A2(n7318), .A3(n7209), .A4(n5736), .ZN(n5737)
         );
  NOR4_X1 U7296 ( .A1(n8593), .A2(n7443), .A3(n8617), .A4(n5737), .ZN(n5738)
         );
  NAND4_X1 U7297 ( .A1(n8542), .A2(n8583), .A3(n8555), .A4(n5738), .ZN(n5739)
         );
  NOR4_X1 U7298 ( .A1(n8487), .A2(n8501), .A3(n8523), .A4(n5739), .ZN(n5740)
         );
  NAND4_X1 U7299 ( .A1(n4625), .A2(n5741), .A3(n8470), .A4(n5740), .ZN(n5742)
         );
  NOR4_X1 U7300 ( .A1(n5888), .A2(n8421), .A3(n5743), .A4(n5742), .ZN(n5744)
         );
  NAND3_X1 U7301 ( .A1(n5745), .A2(n4301), .A3(n5744), .ZN(n5746) );
  XNOR2_X1 U7302 ( .A(n5746), .B(n8433), .ZN(n5748) );
  OAI22_X1 U7303 ( .A1(n5748), .A2(n5480), .B1(n5747), .B2(n5757), .ZN(n5749)
         );
  NAND2_X1 U7304 ( .A1(n5872), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7040) );
  INV_X1 U7305 ( .A(n7040), .ZN(n5751) );
  NOR4_X1 U7306 ( .A1(n9767), .A2(n8621), .A3(n6368), .A4(n5878), .ZN(n5754)
         );
  OAI21_X1 U7307 ( .B1(n7040), .B2(n5508), .A(P2_B_REG_SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7308 ( .A1(n5756), .A2(n5755), .ZN(P2_U3244) );
  NAND2_X1 U7309 ( .A1(n8277), .A2(n6594), .ZN(n5834) );
  INV_X1 U7310 ( .A(n5834), .ZN(n5837) );
  NAND3_X1 U7311 ( .A1(n5757), .A2(n9777), .A3(n6936), .ZN(n5758) );
  XNOR2_X1 U7312 ( .A(n8754), .B(n7527), .ZN(n5835) );
  INV_X1 U7313 ( .A(n5835), .ZN(n5836) );
  NAND2_X1 U7314 ( .A1(n6505), .A2(n6594), .ZN(n5762) );
  XNOR2_X1 U7315 ( .A(n5761), .B(n5762), .ZN(n6514) );
  INV_X1 U7316 ( .A(n6971), .ZN(n5759) );
  NAND2_X1 U7317 ( .A1(n5759), .A2(n6594), .ZN(n6571) );
  NAND2_X1 U7318 ( .A1(n9776), .A2(n5843), .ZN(n5760) );
  AND2_X1 U7319 ( .A1(n6571), .A2(n5760), .ZN(n6515) );
  NAND2_X1 U7320 ( .A1(n6514), .A2(n6515), .ZN(n6508) );
  INV_X1 U7321 ( .A(n5761), .ZN(n5763) );
  NAND2_X1 U7322 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  NAND2_X1 U7323 ( .A1(n6508), .A2(n5764), .ZN(n5765) );
  XNOR2_X1 U7324 ( .A(n9789), .B(n5843), .ZN(n5766) );
  NAND2_X1 U7325 ( .A1(n8289), .A2(n6594), .ZN(n5767) );
  XNOR2_X1 U7326 ( .A(n5766), .B(n5767), .ZN(n6506) );
  INV_X1 U7327 ( .A(n5766), .ZN(n5768) );
  NAND2_X1 U7328 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  INV_X1 U7329 ( .A(n5935), .ZN(n5775) );
  NOR2_X1 U7330 ( .A1(n6847), .A2(n7525), .ZN(n5770) );
  XNOR2_X1 U7331 ( .A(n5093), .B(n5784), .ZN(n6530) );
  NAND2_X1 U7332 ( .A1(n5770), .A2(n6530), .ZN(n5776) );
  INV_X1 U7333 ( .A(n5770), .ZN(n5772) );
  INV_X1 U7334 ( .A(n6530), .ZN(n5771) );
  NAND2_X1 U7335 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U7336 ( .A1(n5776), .A2(n5773), .ZN(n5934) );
  NAND2_X1 U7337 ( .A1(n5775), .A2(n5774), .ZN(n5932) );
  NAND2_X1 U7338 ( .A1(n5095), .A2(n6594), .ZN(n5778) );
  XNOR2_X1 U7339 ( .A(n5778), .B(n8125), .ZN(n6527) );
  NAND2_X1 U7340 ( .A1(n9741), .A2(n6594), .ZN(n5782) );
  XNOR2_X1 U7341 ( .A(n9811), .B(n5784), .ZN(n5781) );
  XNOR2_X1 U7342 ( .A(n5782), .B(n5781), .ZN(n8126) );
  AND2_X1 U7343 ( .A1(n6528), .A2(n8126), .ZN(n5780) );
  INV_X1 U7344 ( .A(n8125), .ZN(n5777) );
  INV_X1 U7345 ( .A(n5781), .ZN(n6581) );
  NAND2_X1 U7346 ( .A1(n5782), .A2(n6581), .ZN(n5783) );
  NAND2_X1 U7347 ( .A1(n6579), .A2(n5783), .ZN(n5785) );
  NAND2_X1 U7348 ( .A1(n8288), .A2(n6594), .ZN(n5788) );
  XNOR2_X1 U7349 ( .A(n6839), .B(n7527), .ZN(n5786) );
  XNOR2_X1 U7350 ( .A(n5788), .B(n5786), .ZN(n6580) );
  INV_X1 U7351 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U7352 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  NOR2_X1 U7353 ( .A1(n7074), .A2(n7525), .ZN(n5790) );
  XNOR2_X1 U7354 ( .A(n6765), .B(n7527), .ZN(n5791) );
  NAND2_X1 U7355 ( .A1(n5790), .A2(n5791), .ZN(n5795) );
  INV_X1 U7356 ( .A(n5790), .ZN(n5792) );
  INV_X1 U7357 ( .A(n5791), .ZN(n6926) );
  NAND2_X1 U7358 ( .A1(n5792), .A2(n6926), .ZN(n5793) );
  NAND2_X1 U7359 ( .A1(n5795), .A2(n5793), .ZN(n5941) );
  INV_X1 U7360 ( .A(n5941), .ZN(n5794) );
  NAND2_X1 U7361 ( .A1(n8286), .A2(n6594), .ZN(n5797) );
  XNOR2_X1 U7362 ( .A(n7233), .B(n7527), .ZN(n5798) );
  XNOR2_X1 U7363 ( .A(n5797), .B(n5798), .ZN(n6927) );
  XNOR2_X1 U7364 ( .A(n7157), .B(n5843), .ZN(n5803) );
  NAND2_X1 U7365 ( .A1(n8285), .A2(n6594), .ZN(n5804) );
  NAND2_X1 U7366 ( .A1(n5803), .A2(n5804), .ZN(n6954) );
  AND2_X1 U7367 ( .A1(n6927), .A2(n6954), .ZN(n5796) );
  NAND2_X1 U7368 ( .A1(n6928), .A2(n5796), .ZN(n5802) );
  INV_X1 U7369 ( .A(n6954), .ZN(n5800) );
  INV_X1 U7370 ( .A(n5797), .ZN(n5799) );
  NAND2_X1 U7371 ( .A1(n5799), .A2(n5798), .ZN(n6955) );
  OR2_X1 U7372 ( .A1(n5800), .A2(n6955), .ZN(n5801) );
  INV_X1 U7373 ( .A(n5803), .ZN(n5806) );
  INV_X1 U7374 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U7375 ( .A1(n5806), .A2(n5805), .ZN(n6953) );
  XNOR2_X1 U7376 ( .A(n7455), .B(n7527), .ZN(n5809) );
  NAND2_X1 U7377 ( .A1(n8284), .A2(n6594), .ZN(n5807) );
  XNOR2_X1 U7378 ( .A(n5809), .B(n5807), .ZN(n6989) );
  INV_X1 U7379 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U7380 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  XNOR2_X1 U7381 ( .A(n7226), .B(n7527), .ZN(n5813) );
  NAND2_X1 U7382 ( .A1(n8283), .A2(n6594), .ZN(n5811) );
  XNOR2_X1 U7383 ( .A(n5813), .B(n5811), .ZN(n7161) );
  NAND2_X1 U7384 ( .A1(n7160), .A2(n7161), .ZN(n5815) );
  INV_X1 U7385 ( .A(n5811), .ZN(n5812) );
  NAND2_X1 U7386 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7387 ( .A1(n5815), .A2(n5814), .ZN(n7168) );
  XNOR2_X1 U7388 ( .A(n7210), .B(n7527), .ZN(n5818) );
  NAND2_X1 U7389 ( .A1(n8282), .A2(n6594), .ZN(n5816) );
  XNOR2_X1 U7390 ( .A(n5818), .B(n5816), .ZN(n7169) );
  NAND2_X1 U7391 ( .A1(n7168), .A2(n7169), .ZN(n5820) );
  INV_X1 U7392 ( .A(n5816), .ZN(n5817) );
  NAND2_X1 U7393 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  XNOR2_X1 U7394 ( .A(n7503), .B(n7527), .ZN(n7301) );
  NAND2_X1 U7395 ( .A1(n8281), .A2(n6594), .ZN(n7300) );
  XNOR2_X1 U7396 ( .A(n7493), .B(n7527), .ZN(n5821) );
  NAND2_X1 U7397 ( .A1(n8280), .A2(n6594), .ZN(n5822) );
  XNOR2_X1 U7398 ( .A(n5821), .B(n5822), .ZN(n7430) );
  INV_X1 U7399 ( .A(n5821), .ZN(n5823) );
  NAND2_X1 U7400 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  XNOR2_X1 U7401 ( .A(n8629), .B(n7527), .ZN(n8195) );
  NOR2_X1 U7402 ( .A1(n8595), .A2(n7525), .ZN(n5827) );
  NOR2_X1 U7403 ( .A1(n8622), .A2(n7525), .ZN(n5826) );
  XNOR2_X1 U7404 ( .A(n7448), .B(n7527), .ZN(n8191) );
  AOI22_X1 U7405 ( .A1(n8195), .A2(n5827), .B1(n5826), .B2(n8191), .ZN(n5831)
         );
  INV_X1 U7406 ( .A(n8191), .ZN(n8193) );
  INV_X1 U7407 ( .A(n5826), .ZN(n8257) );
  INV_X1 U7408 ( .A(n5827), .ZN(n8194) );
  AOI21_X1 U7409 ( .B1(n8193), .B2(n8257), .A(n8194), .ZN(n5829) );
  NAND3_X1 U7410 ( .A1(n8193), .A2(n8257), .A3(n8194), .ZN(n5828) );
  OAI21_X1 U7411 ( .B1(n8195), .B2(n5829), .A(n5828), .ZN(n5830) );
  XNOR2_X1 U7412 ( .A(n8610), .B(n5843), .ZN(n8243) );
  NAND2_X1 U7413 ( .A1(n5315), .A2(n6594), .ZN(n5832) );
  NOR2_X1 U7414 ( .A1(n8243), .A2(n5832), .ZN(n5833) );
  AOI21_X1 U7415 ( .B1(n8243), .B2(n5832), .A(n5833), .ZN(n8205) );
  XNOR2_X1 U7416 ( .A(n5835), .B(n5834), .ZN(n8245) );
  XNOR2_X1 U7417 ( .A(n8574), .B(n7527), .ZN(n5840) );
  INV_X1 U7418 ( .A(n5840), .ZN(n8162) );
  NAND2_X1 U7419 ( .A1(n8539), .A2(n6594), .ZN(n5839) );
  INV_X1 U7420 ( .A(n5839), .ZN(n5838) );
  NAND2_X1 U7421 ( .A1(n8162), .A2(n5838), .ZN(n8164) );
  NOR2_X1 U7422 ( .A1(n8567), .A2(n7525), .ZN(n5842) );
  XNOR2_X1 U7423 ( .A(n8681), .B(n7527), .ZN(n5841) );
  XOR2_X1 U7424 ( .A(n5842), .B(n5841), .Z(n8221) );
  XNOR2_X1 U7425 ( .A(n8676), .B(n5843), .ZN(n5845) );
  NAND2_X1 U7426 ( .A1(n8540), .A2(n6594), .ZN(n5844) );
  XNOR2_X1 U7427 ( .A(n5845), .B(n5844), .ZN(n8173) );
  XNOR2_X1 U7428 ( .A(n8511), .B(n7527), .ZN(n5848) );
  XNOR2_X1 U7429 ( .A(n5847), .B(n5848), .ZN(n8239) );
  INV_X1 U7430 ( .A(n5847), .ZN(n5850) );
  INV_X1 U7431 ( .A(n5848), .ZN(n5849) );
  XNOR2_X1 U7432 ( .A(n8665), .B(n7527), .ZN(n5852) );
  NAND2_X1 U7433 ( .A1(n8505), .A2(n6594), .ZN(n8152) );
  XNOR2_X1 U7434 ( .A(n5855), .B(n5853), .ZN(n8215) );
  NOR2_X1 U7435 ( .A1(n8213), .A2(n7525), .ZN(n8214) );
  INV_X1 U7436 ( .A(n5853), .ZN(n5854) );
  AOI21_X2 U7437 ( .B1(n8215), .B2(n8214), .A(n5856), .ZN(n8180) );
  XNOR2_X1 U7438 ( .A(n8738), .B(n7527), .ZN(n8182) );
  NAND2_X1 U7439 ( .A1(n8275), .A2(n6594), .ZN(n8181) );
  NAND2_X1 U7440 ( .A1(n8180), .A2(n8182), .ZN(n5857) );
  XNOR2_X1 U7441 ( .A(n8443), .B(n7527), .ZN(n8139) );
  NOR2_X1 U7442 ( .A1(n8184), .A2(n7525), .ZN(n5859) );
  NAND2_X1 U7443 ( .A1(n8139), .A2(n5859), .ZN(n7516) );
  OAI21_X1 U7444 ( .B1(n8139), .B2(n5859), .A(n7516), .ZN(n5860) );
  NAND2_X1 U7445 ( .A1(n5861), .A2(n5860), .ZN(n5867) );
  AND2_X1 U7446 ( .A1(n5863), .A2(n5862), .ZN(n6588) );
  NAND2_X1 U7447 ( .A1(n5864), .A2(n6588), .ZN(n5871) );
  INV_X1 U7448 ( .A(n6353), .ZN(n6034) );
  NAND2_X1 U7449 ( .A1(n6034), .A2(n9835), .ZN(n5865) );
  NAND2_X1 U7450 ( .A1(n5867), .A2(n5866), .ZN(n5884) );
  NOR2_X1 U7451 ( .A1(n9777), .A2(n6857), .ZN(n6593) );
  INV_X1 U7452 ( .A(n6593), .ZN(n5868) );
  OR2_X1 U7453 ( .A1(n5879), .A2(n5868), .ZN(n5869) );
  NAND2_X1 U7454 ( .A1(n5871), .A2(n5870), .ZN(n5876) );
  NOR2_X1 U7455 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AND2_X1 U7456 ( .A1(n6351), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U7457 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  AOI22_X1 U7458 ( .A1(n8439), .A2(n8266), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n5881) );
  NOR2_X1 U7459 ( .A1(n8264), .A2(n8619), .ZN(n8198) );
  NOR2_X1 U7460 ( .A1(n8264), .A2(n8621), .ZN(n8199) );
  AOI22_X1 U7461 ( .A1(n8273), .A2(n8198), .B1(n8199), .B2(n8275), .ZN(n5880)
         );
  OAI211_X1 U7462 ( .C1(n8734), .C2(n8270), .A(n5881), .B(n5880), .ZN(n5882)
         );
  INV_X1 U7463 ( .A(n5882), .ZN(n5883) );
  OAI21_X1 U7464 ( .B1(n8272), .B2(n7532), .A(n5885), .ZN(n5886) );
  XNOR2_X1 U7465 ( .A(n5886), .B(n5888), .ZN(n8394) );
  XOR2_X1 U7466 ( .A(n5888), .B(n5887), .Z(n5894) );
  NAND2_X1 U7467 ( .A1(n8272), .A2(n9742), .ZN(n5892) );
  INV_X1 U7468 ( .A(P2_B_REG_SCAN_IN), .ZN(n5889) );
  NOR2_X1 U7469 ( .A1(n6368), .A2(n5889), .ZN(n5890) );
  NOR2_X1 U7470 ( .A1(n8619), .A2(n5890), .ZN(n8383) );
  NAND2_X1 U7471 ( .A1(n5895), .A2(n5902), .ZN(n8382) );
  INV_X1 U7472 ( .A(n9826), .ZN(n8603) );
  OAI211_X1 U7473 ( .C1(n5895), .C2(n5902), .A(n8382), .B(n8603), .ZN(n8397)
         );
  AOI21_X1 U7474 ( .B1(n8394), .B2(n9838), .A(n5896), .ZN(n5905) );
  NOR2_X1 U7475 ( .A1(n9840), .A2(n5897), .ZN(n5898) );
  OAI21_X1 U7476 ( .B1(n5905), .B2(n5900), .A(n5899), .ZN(P2_U3517) );
  NAND2_X1 U7477 ( .A1(n9853), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5901) );
  OAI21_X1 U7478 ( .B1(n5905), .B2(n9853), .A(n5904), .ZN(P2_U3549) );
  NOR2_X1 U7479 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5909) );
  NAND4_X1 U7480 ( .A1(n5909), .A2(n5908), .A3(n6121), .A4(n6336), .ZN(n5914)
         );
  INV_X1 U7481 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5912) );
  INV_X1 U7482 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5911) );
  INV_X1 U7483 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5910) );
  NAND4_X1 U7484 ( .A1(n5912), .A2(n5911), .A3(n6021), .A4(n5910), .ZN(n5913)
         );
  NOR3_X1 U7485 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n5918) );
  NOR2_X1 U7486 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5916) );
  NOR2_X1 U7487 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5915) );
  NAND2_X1 U7488 ( .A1(n5947), .A2(n5919), .ZN(n5920) );
  NAND2_X1 U7489 ( .A1(n5923), .A2(n5955), .ZN(n5921) );
  XNOR2_X1 U7490 ( .A(n5923), .B(n5955), .ZN(n7377) );
  NAND2_X1 U7491 ( .A1(n5924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U7492 ( .A(n5926), .B(n5925), .ZN(n7167) );
  INV_X1 U7493 ( .A(n6199), .ZN(n6127) );
  INV_X1 U7494 ( .A(n5927), .ZN(n5928) );
  NAND2_X1 U7495 ( .A1(n5928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7496 ( .A(n5930), .B(n5929), .ZN(n7042) );
  NAND2_X1 U7497 ( .A1(n6127), .A2(n7042), .ZN(n5979) );
  NOR2_X1 U7498 ( .A1(n5979), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U7499 ( .A(n6351), .ZN(n5931) );
  INV_X1 U7500 ( .A(n6529), .ZN(n5933) );
  AOI211_X1 U7501 ( .C1(n5935), .C2(n5934), .A(n8244), .B(n5933), .ZN(n5939)
         );
  INV_X1 U7502 ( .A(n8289), .ZN(n6516) );
  NOR2_X1 U7503 ( .A1(n8233), .A2(n6516), .ZN(n5938) );
  INV_X1 U7504 ( .A(n8198), .ZN(n8234) );
  OAI22_X1 U7505 ( .A1(n8234), .A2(n6917), .B1(n9797), .B2(n8270), .ZN(n5937)
         );
  INV_X1 U7506 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8295) );
  OAI22_X1 U7507 ( .A1(n8251), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n8295), .ZN(n5936) );
  OR4_X1 U7508 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(P2_U3220)
         );
  INV_X1 U7509 ( .A(n6925), .ZN(n5940) );
  AOI211_X1 U7510 ( .C1(n5942), .C2(n5941), .A(n8244), .B(n5940), .ZN(n5946)
         );
  NOR2_X1 U7511 ( .A1(n8270), .A2(n9820), .ZN(n5945) );
  OAI22_X1 U7512 ( .A1(n7146), .A2(n8234), .B1(n8233), .B2(n6916), .ZN(n5944)
         );
  OAI22_X1 U7513 ( .A1(n8251), .A2(n6762), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6463), .ZN(n5943) );
  OR4_X1 U7514 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(P2_U3215)
         );
  NAND2_X1 U7515 ( .A1(n6016), .A2(n5947), .ZN(n6058) );
  INV_X1 U7516 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6057) );
  INV_X1 U7517 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7518 ( .A1(n6075), .A2(n6103), .ZN(n8068) );
  INV_X1 U7519 ( .A(n7042), .ZN(n5952) );
  OR2_X1 U7520 ( .A1(n8068), .A2(n5952), .ZN(n5953) );
  NAND2_X1 U7521 ( .A1(n5953), .A2(n5979), .ZN(n5965) );
  INV_X1 U7522 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7523 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5957) );
  OR2_X1 U7524 ( .A1(n5965), .A2(n7648), .ZN(n6044) );
  NAND2_X1 U7525 ( .A1(n6044), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7526 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7527 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5962), .ZN(n5959) );
  XNOR2_X1 U7528 ( .A(n5959), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U7529 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5960) );
  NAND2_X1 U7530 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9507) );
  NAND2_X1 U7531 ( .A1(n5986), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U7532 ( .B1(n5986), .B2(P1_REG2_REG_1__SCAN_IN), .A(n5961), .ZN(
        n9492) );
  NOR2_X1 U7533 ( .A1(n9507), .A2(n9492), .ZN(n9491) );
  XNOR2_X1 U7534 ( .A(n9515), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9505) );
  OAI21_X1 U7535 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(n5962), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7536 ( .A(n5963), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7537 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6275), .ZN(n5964) );
  OAI21_X1 U7538 ( .B1(n6275), .B2(P1_REG2_REG_3__SCAN_IN), .A(n5964), .ZN(
        n5968) );
  OR2_X1 U7539 ( .A1(n5965), .A2(P1_U3084), .ZN(n5973) );
  NOR2_X1 U7540 ( .A1(n5973), .A2(n4278), .ZN(n5978) );
  INV_X1 U7541 ( .A(n8123), .ZN(n9512) );
  AND2_X1 U7542 ( .A1(n5978), .A2(n9512), .ZN(n9609) );
  INV_X1 U7543 ( .A(n9609), .ZN(n9578) );
  AOI211_X1 U7544 ( .C1(n5969), .C2(n5968), .A(n6263), .B(n9578), .ZN(n5984)
         );
  INV_X1 U7545 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6133) );
  INV_X1 U7546 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7547 ( .A1(n5986), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5970) );
  OAI21_X1 U7548 ( .B1(n5986), .B2(P1_REG1_REG_1__SCAN_IN), .A(n5970), .ZN(
        n9489) );
  NOR3_X1 U7549 ( .A1(n6133), .A2(n6099), .A3(n9489), .ZN(n9488) );
  AOI21_X1 U7550 ( .B1(n5986), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9488), .ZN(
        n9502) );
  NAND2_X1 U7551 ( .A1(n9515), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5971) );
  OAI21_X1 U7552 ( .B1(n9515), .B2(P1_REG1_REG_2__SCAN_IN), .A(n5971), .ZN(
        n9501) );
  NOR2_X1 U7553 ( .A1(n9502), .A2(n9501), .ZN(n9500) );
  NAND2_X1 U7554 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6275), .ZN(n5972) );
  OAI21_X1 U7555 ( .B1(n6275), .B2(P1_REG1_REG_3__SCAN_IN), .A(n5972), .ZN(
        n5976) );
  NOR2_X1 U7556 ( .A1(n5977), .A2(n5976), .ZN(n6274) );
  INV_X1 U7557 ( .A(n5973), .ZN(n5975) );
  INV_X1 U7558 ( .A(n4278), .ZN(n6042) );
  NOR2_X1 U7559 ( .A1(n8123), .A2(n6042), .ZN(n5974) );
  NAND2_X1 U7560 ( .A1(n5975), .A2(n5974), .ZN(n9536) );
  AOI211_X1 U7561 ( .C1(n5977), .C2(n5976), .A(n6274), .B(n9536), .ZN(n5983)
         );
  INV_X1 U7562 ( .A(n6275), .ZN(n6219) );
  NAND2_X1 U7563 ( .A1(n5978), .A2(n8123), .ZN(n9613) );
  INV_X1 U7564 ( .A(P1_U3083), .ZN(n5980) );
  NAND2_X1 U7565 ( .A1(n5980), .A2(n5979), .ZN(n9605) );
  INV_X1 U7566 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n5981) );
  OAI22_X1 U7567 ( .A1(n6219), .A2(n9613), .B1(n9605), .B2(n5981), .ZN(n5982)
         );
  OR4_X1 U7568 ( .A1(n6234), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(P1_U3244)
         );
  NOR2_X1 U7569 ( .A1(n6156), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8780) );
  AOI22_X1 U7570 ( .A1(n8780), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8297), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n5985) );
  OAI21_X1 U7571 ( .B1(n6214), .B2(n8783), .A(n5985), .ZN(P2_U3355) );
  NAND2_X1 U7572 ( .A1(n6156), .A2(P1_U3084), .ZN(n8121) );
  INV_X1 U7573 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5987) );
  NOR2_X1 U7574 ( .A1(n6156), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9398) );
  INV_X1 U7575 ( .A(n5986), .ZN(n9496) );
  OAI222_X1 U7576 ( .A1(n8121), .A2(n5987), .B1(n9402), .B2(n6159), .C1(
        P1_U3084), .C2(n9496), .ZN(P1_U3352) );
  INV_X1 U7577 ( .A(n8780), .ZN(n7376) );
  INV_X1 U7578 ( .A(n9423), .ZN(n6348) );
  OAI222_X1 U7579 ( .A1(n7376), .A2(n5988), .B1(n8783), .B2(n6180), .C1(
        P2_U3152), .C2(n6348), .ZN(P2_U3356) );
  OAI222_X1 U7580 ( .A1(n7376), .A2(n5033), .B1(n8783), .B2(n6159), .C1(
        P2_U3152), .C2(n6344), .ZN(P2_U3357) );
  INV_X1 U7581 ( .A(n6428), .ZN(n6374) );
  OAI222_X1 U7582 ( .A1(n7376), .A2(n5989), .B1(n8783), .B2(n6300), .C1(
        P2_U3152), .C2(n6374), .ZN(P2_U3354) );
  AOI22_X1 U7583 ( .A1(n8311), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8780), .ZN(n5990) );
  OAI21_X1 U7584 ( .B1(n6475), .B2(n8783), .A(n5990), .ZN(P2_U3353) );
  INV_X1 U7585 ( .A(n8121), .ZN(n6339) );
  INV_X1 U7586 ( .A(n6339), .ZN(n9404) );
  INV_X1 U7587 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7588 ( .A1(n5991), .A2(n6119), .ZN(n5992) );
  XNOR2_X1 U7589 ( .A(n5992), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9523) );
  INV_X1 U7590 ( .A(n9523), .ZN(n6304) );
  OAI222_X1 U7591 ( .A1(n9404), .A2(n6301), .B1(n9402), .B2(n6300), .C1(
        P1_U3084), .C2(n6304), .ZN(P1_U3349) );
  NAND2_X1 U7592 ( .A1(n5993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5994) );
  MUX2_X1 U7593 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5994), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5995) );
  AND2_X1 U7594 ( .A1(n5995), .A2(n5996), .ZN(n6276) );
  INV_X1 U7595 ( .A(n6276), .ZN(n9543) );
  OAI222_X1 U7596 ( .A1(n9404), .A2(n6476), .B1(n9402), .B2(n6475), .C1(
        P1_U3084), .C2(n9543), .ZN(P1_U3348) );
  OAI222_X1 U7597 ( .A1(n9404), .A2(n6216), .B1(n9402), .B2(n6214), .C1(
        P1_U3084), .C2(n6219), .ZN(P1_U3350) );
  INV_X1 U7598 ( .A(n9515), .ZN(n6183) );
  OAI222_X1 U7599 ( .A1(n9404), .A2(n6181), .B1(n9402), .B2(n6180), .C1(
        P1_U3084), .C2(n6183), .ZN(P1_U3351) );
  INV_X1 U7600 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7601 ( .A1(n5996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7602 ( .A(n5997), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6542) );
  INV_X1 U7603 ( .A(n6542), .ZN(n9559) );
  OAI222_X1 U7604 ( .A1(n9404), .A2(n5998), .B1(n9402), .B2(n5999), .C1(
        P1_U3084), .C2(n9559), .ZN(P1_U3347) );
  INV_X1 U7605 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6000) );
  INV_X1 U7606 ( .A(n6437), .ZN(n6445) );
  OAI222_X1 U7607 ( .A1(n7376), .A2(n6000), .B1(n8783), .B2(n5999), .C1(
        P2_U3152), .C2(n6445), .ZN(P2_U3352) );
  AND2_X1 U7608 ( .A1(n7042), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7609 ( .A1(n6199), .A2(n6001), .ZN(n9393) );
  INV_X1 U7610 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7611 ( .A1(n7377), .A2(P1_B_REG_SCAN_IN), .ZN(n6002) );
  MUX2_X1 U7612 ( .A(P1_B_REG_SCAN_IN), .B(n6002), .S(n7167), .Z(n6004) );
  INV_X1 U7613 ( .A(n7386), .ZN(n6003) );
  NAND2_X1 U7614 ( .A1(n6004), .A2(n6003), .ZN(n6076) );
  NAND2_X1 U7615 ( .A1(n6146), .A2(n6076), .ZN(n9650) );
  INV_X1 U7616 ( .A(n9650), .ZN(n9649) );
  NAND2_X1 U7617 ( .A1(n4269), .A2(n7377), .ZN(n6077) );
  OAI21_X1 U7618 ( .B1(n9649), .B2(P1_D_REG_1__SCAN_IN), .A(n6077), .ZN(n6005)
         );
  OAI21_X1 U7619 ( .B1(n6146), .B2(n6006), .A(n6005), .ZN(P1_U3441) );
  INV_X1 U7620 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6009) );
  INV_X1 U7621 ( .A(n6639), .ZN(n6010) );
  OR2_X1 U7622 ( .A1(n6007), .A2(n6119), .ZN(n6008) );
  XNOR2_X1 U7623 ( .A(n6008), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6640) );
  INV_X1 U7624 ( .A(n6640), .ZN(n8938) );
  OAI222_X1 U7625 ( .A1(n9404), .A2(n6009), .B1(n9402), .B2(n6010), .C1(
        P1_U3084), .C2(n8938), .ZN(P1_U3346) );
  INV_X1 U7626 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6011) );
  OAI222_X1 U7627 ( .A1(n7376), .A2(n6011), .B1(n8783), .B2(n6010), .C1(
        P2_U3152), .C2(n6474), .ZN(P2_U3351) );
  INV_X1 U7628 ( .A(n6644), .ZN(n6015) );
  NAND2_X1 U7629 ( .A1(n6012), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U7630 ( .A(n6013), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6645) );
  INV_X1 U7631 ( .A(n6645), .ZN(n6267) );
  OAI222_X1 U7632 ( .A1(n8121), .A2(n6014), .B1(n9402), .B2(n6015), .C1(
        P1_U3084), .C2(n6267), .ZN(P1_U3345) );
  OAI222_X1 U7633 ( .A1(n7376), .A2(n9959), .B1(n8783), .B2(n6015), .C1(
        P2_U3152), .C2(n6458), .ZN(P2_U3350) );
  INV_X1 U7634 ( .A(n6730), .ZN(n6025) );
  NAND2_X1 U7635 ( .A1(n6019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7636 ( .A(n6017), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9572) );
  AOI22_X1 U7637 ( .A1(n9572), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6339), .ZN(n6018) );
  OAI21_X1 U7638 ( .B1(n6025), .B2(n9402), .A(n6018), .ZN(P1_U3344) );
  INV_X1 U7639 ( .A(n6862), .ZN(n6027) );
  NOR2_X1 U7640 ( .A1(n6019), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6050) );
  NOR2_X1 U7641 ( .A1(n6050), .A2(n6119), .ZN(n6020) );
  NAND2_X1 U7642 ( .A1(n6020), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6023) );
  INV_X1 U7643 ( .A(n6020), .ZN(n6022) );
  NAND2_X1 U7644 ( .A1(n6022), .A2(n6021), .ZN(n6029) );
  INV_X1 U7645 ( .A(n6863), .ZN(n9585) );
  OAI222_X1 U7646 ( .A1(n9402), .A2(n6027), .B1(n9585), .B2(P1_U3084), .C1(
        n6024), .C2(n9404), .ZN(P1_U3343) );
  OAI222_X1 U7647 ( .A1(n7376), .A2(n6026), .B1(n8783), .B2(n6025), .C1(n6686), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U7648 ( .A1(n7376), .A2(n9970), .B1(n8783), .B2(n6027), .C1(n6690), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7649 ( .A(n6996), .ZN(n6032) );
  AOI22_X1 U7650 ( .A1(n6818), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8780), .ZN(n6028) );
  OAI21_X1 U7651 ( .B1(n6032), .B2(n8783), .A(n6028), .ZN(P2_U3347) );
  NAND2_X1 U7652 ( .A1(n6029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U7653 ( .A(n6030), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9592) );
  INV_X1 U7654 ( .A(n9592), .ZN(n6400) );
  OAI222_X1 U7655 ( .A1(n9402), .A2(n6032), .B1(n6400), .B2(P1_U3084), .C1(
        n6031), .C2(n9404), .ZN(P1_U3342) );
  OR2_X1 U7656 ( .A1(n7040), .A2(n6354), .ZN(n6033) );
  NAND2_X1 U7657 ( .A1(n9767), .A2(n6033), .ZN(n6036) );
  NAND2_X1 U7658 ( .A1(n6034), .A2(n6354), .ZN(n6035) );
  NAND2_X1 U7659 ( .A1(n6036), .A2(n6035), .ZN(n9731) );
  NOR2_X1 U7660 ( .A1(n9417), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7661 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7662 ( .A1(n6037), .A2(P2_U3966), .ZN(n6038) );
  OAI21_X1 U7663 ( .B1(n6039), .B2(P2_U3966), .A(n6038), .ZN(P2_U3583) );
  INV_X1 U7664 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6048) );
  INV_X1 U7665 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U7666 ( .A1(n6042), .A2(n10011), .ZN(n6040) );
  AOI21_X1 U7667 ( .B1(n9512), .B2(n6040), .A(P1_IR_REG_0__SCAN_IN), .ZN(n9511) );
  NAND3_X1 U7668 ( .A1(n9512), .A2(n6040), .A3(P1_IR_REG_0__SCAN_IN), .ZN(
        n6041) );
  OAI211_X1 U7669 ( .C1(n6042), .C2(P1_REG1_REG_0__SCAN_IN), .A(n6041), .B(
        P1_STATE_REG_SCAN_IN), .ZN(n6043) );
  NOR3_X1 U7670 ( .A1(n6044), .A2(n9511), .A3(n6043), .ZN(n6046) );
  NOR3_X1 U7671 ( .A1(n9536), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6133), .ZN(
        n6045) );
  AOI211_X1 U7672 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6046), .B(
        n6045), .ZN(n6047) );
  OAI21_X1 U7673 ( .B1(n9605), .B2(n6048), .A(n6047), .ZN(P1_U3241) );
  INV_X1 U7674 ( .A(n7180), .ZN(n6054) );
  OAI222_X1 U7675 ( .A1(n7376), .A2(n9928), .B1(n8783), .B2(n6054), .C1(
        P2_U3152), .C2(n6828), .ZN(P2_U3346) );
  NOR2_X1 U7676 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6049) );
  NAND2_X1 U7677 ( .A1(n6050), .A2(n6049), .ZN(n6052) );
  NAND2_X1 U7678 ( .A1(n6052), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6051) );
  MUX2_X1 U7679 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6051), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6053) );
  INV_X1 U7680 ( .A(n7181), .ZN(n6406) );
  OAI222_X1 U7681 ( .A1(n8121), .A2(n6055), .B1(n9402), .B2(n6054), .C1(
        P1_U3084), .C2(n6406), .ZN(P1_U3341) );
  NAND2_X1 U7682 ( .A1(n6058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6060) );
  INV_X1 U7683 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6059) );
  XNOR2_X1 U7684 ( .A(n6060), .B(n6059), .ZN(n8994) );
  AND2_X1 U7685 ( .A1(n6102), .A2(n8994), .ZN(n8110) );
  OR2_X1 U7686 ( .A1(n8068), .A2(n8110), .ZN(n6200) );
  NAND2_X1 U7687 ( .A1(n6200), .A2(n6146), .ZN(n6255) );
  OR2_X1 U7688 ( .A1(n6076), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7689 ( .A1(n4269), .A2(n7167), .ZN(n6061) );
  AND2_X1 U7690 ( .A1(n6062), .A2(n6061), .ZN(n9394) );
  INV_X1 U7691 ( .A(n9394), .ZN(n6073) );
  NOR4_X1 U7692 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6071) );
  NOR4_X1 U7693 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6070) );
  OR4_X1 U7694 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6068) );
  NOR4_X1 U7695 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6066) );
  NOR4_X1 U7696 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6065) );
  NOR4_X1 U7697 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6064) );
  NOR4_X1 U7698 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7699 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6067)
         );
  NOR4_X1 U7700 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6068), .A4(n6067), .ZN(n6069) );
  AND3_X1 U7701 ( .A1(n6071), .A2(n6070), .A3(n6069), .ZN(n6072) );
  OR2_X1 U7702 ( .A1(n6076), .A2(n6072), .ZN(n6138) );
  NAND2_X1 U7703 ( .A1(n6073), .A2(n6138), .ZN(n6074) );
  NOR2_X1 U7704 ( .A1(n6255), .A2(n6074), .ZN(n6284) );
  INV_X1 U7705 ( .A(n8111), .ZN(n6244) );
  OR2_X1 U7706 ( .A1(n9458), .A2(n8994), .ZN(n6080) );
  OR2_X1 U7707 ( .A1(n6076), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6078) );
  AND2_X1 U7708 ( .A1(n6078), .A2(n6077), .ZN(n6283) );
  INV_X1 U7709 ( .A(n6283), .ZN(n6079) );
  AND2_X2 U7710 ( .A1(n6284), .A2(n6257), .ZN(n9709) );
  INV_X1 U7711 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6113) );
  INV_X1 U7712 ( .A(SI_0_), .ZN(n6082) );
  INV_X1 U7713 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U7714 ( .B1(n6156), .B2(n6082), .A(n6081), .ZN(n6084) );
  AND2_X1 U7715 ( .A1(n6084), .A2(n6083), .ZN(n9405) );
  INV_X1 U7716 ( .A(n6290), .ZN(n8071) );
  INV_X1 U7717 ( .A(n6086), .ZN(n6088) );
  NOR3_X1 U7718 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7719 ( .A1(n6088), .A2(n6087), .ZN(n6094) );
  INV_X1 U7720 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6287) );
  OAI22_X1 U7721 ( .A1(n7655), .A2(n6287), .B1(n6227), .B2(n6113), .ZN(n6101)
         );
  OAI22_X1 U7722 ( .A1(n7858), .A2(n6099), .B1(n6230), .B2(n10011), .ZN(n6100)
         );
  OR2_X2 U7723 ( .A1(n6101), .A2(n6100), .ZN(n8937) );
  XNOR2_X1 U7724 ( .A(n8937), .B(n6290), .ZN(n7977) );
  NAND2_X1 U7725 ( .A1(n6075), .A2(n8994), .ZN(n6237) );
  OR2_X1 U7726 ( .A1(n6237), .A2(n6152), .ZN(n6709) );
  NAND2_X1 U7727 ( .A1(n6709), .A2(n6286), .ZN(n6110) );
  INV_X1 U7728 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6785) );
  INV_X1 U7729 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6104) );
  OAI22_X1 U7730 ( .A1(n7655), .A2(n6785), .B1(n6227), .B2(n6104), .ZN(n6105)
         );
  INV_X1 U7731 ( .A(n6105), .ZN(n6109) );
  INV_X1 U7732 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6106) );
  INV_X1 U7733 ( .A(n6107), .ZN(n6108) );
  INV_X1 U7734 ( .A(n6241), .ZN(n8073) );
  OAI22_X1 U7735 ( .A1(n7977), .A2(n6110), .B1(n8073), .B2(n9289), .ZN(n6111)
         );
  INV_X1 U7736 ( .A(n6111), .ZN(n6292) );
  OAI21_X1 U7737 ( .B1(n8071), .B2(n6286), .A(n6292), .ZN(n9375) );
  NAND2_X1 U7738 ( .A1(n9375), .A2(n9709), .ZN(n6112) );
  OAI21_X1 U7739 ( .B1(n9709), .B2(n6113), .A(n6112), .ZN(P1_U3454) );
  INV_X1 U7740 ( .A(n7390), .ZN(n6116) );
  NAND2_X1 U7741 ( .A1(n6118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7742 ( .A(n6114), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7391) );
  AOI22_X1 U7743 ( .A1(n7391), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6339), .ZN(n6115) );
  OAI21_X1 U7744 ( .B1(n6116), .B2(n9402), .A(n6115), .ZN(P1_U3340) );
  OAI222_X1 U7745 ( .A1(n7376), .A2(n6117), .B1(n8783), .B2(n6116), .C1(n7089), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7746 ( .A(n7557), .ZN(n6125) );
  NOR2_X1 U7747 ( .A1(n6118), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6330) );
  NOR2_X1 U7748 ( .A1(n6330), .A2(n6119), .ZN(n6120) );
  NAND2_X1 U7749 ( .A1(n6120), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6123) );
  INV_X1 U7750 ( .A(n6120), .ZN(n6122) );
  NAND2_X1 U7751 ( .A1(n6122), .A2(n6121), .ZN(n6323) );
  AND2_X1 U7752 ( .A1(n6123), .A2(n6323), .ZN(n7558) );
  INV_X1 U7753 ( .A(n7558), .ZN(n7289) );
  OAI222_X1 U7754 ( .A1(n9402), .A2(n6125), .B1(n7289), .B2(P1_U3084), .C1(
        n6124), .C2(n9404), .ZN(P1_U3339) );
  OAI222_X1 U7755 ( .A1(n7376), .A2(n6126), .B1(n8783), .B2(n6125), .C1(n7419), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U7756 ( .A1(n8937), .A2(n6167), .ZN(n6131) );
  NAND2_X1 U7757 ( .A1(n6290), .A2(n6164), .ZN(n6129) );
  NAND2_X1 U7758 ( .A1(n6127), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6128) );
  AND2_X1 U7759 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NOR2_X1 U7760 ( .A1(n6199), .A2(n6133), .ZN(n6134) );
  AOI21_X1 U7761 ( .B1(n4271), .B2(n6290), .A(n6134), .ZN(n6135) );
  INV_X1 U7762 ( .A(n6135), .ZN(n6136) );
  AOI21_X1 U7763 ( .B1(n4270), .B2(n8937), .A(n6136), .ZN(n6137) );
  NAND2_X1 U7764 ( .A1(n6151), .A2(n6137), .ZN(n6154) );
  OAI21_X1 U7765 ( .B1(n6151), .B2(n6137), .A(n6154), .ZN(n9508) );
  AND2_X1 U7766 ( .A1(n9394), .A2(n6138), .ZN(n6253) );
  NAND2_X1 U7767 ( .A1(n6253), .A2(n6283), .ZN(n6143) );
  INV_X1 U7768 ( .A(n6143), .ZN(n6145) );
  AND2_X1 U7769 ( .A1(n8068), .A2(n6146), .ZN(n6139) );
  AND2_X1 U7770 ( .A1(n6139), .A2(n9701), .ZN(n6140) );
  NAND2_X1 U7771 ( .A1(n6145), .A2(n6140), .ZN(n8923) );
  OR2_X1 U7772 ( .A1(n6286), .A2(n8111), .ZN(n6673) );
  INV_X1 U7773 ( .A(n6673), .ZN(n6141) );
  NAND3_X1 U7774 ( .A1(n6143), .A2(n6141), .A3(n6146), .ZN(n6204) );
  INV_X1 U7775 ( .A(n6255), .ZN(n6142) );
  NAND2_X1 U7776 ( .A1(n6143), .A2(n9701), .ZN(n6201) );
  NAND3_X1 U7777 ( .A1(n6204), .A2(n6142), .A3(n6201), .ZN(n8828) );
  AOI22_X1 U7778 ( .A1(n9508), .A2(n8898), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8828), .ZN(n6150) );
  OR2_X1 U7779 ( .A1(n6709), .A2(n9393), .ZN(n8116) );
  NOR2_X1 U7780 ( .A1(n8116), .A2(n6143), .ZN(n6195) );
  NAND2_X1 U7781 ( .A1(n6195), .A2(n8123), .ZN(n8904) );
  NOR2_X1 U7782 ( .A1(n6673), .A2(n9393), .ZN(n6144) );
  NAND2_X1 U7783 ( .A1(n6145), .A2(n6144), .ZN(n6148) );
  INV_X1 U7784 ( .A(n8994), .ZN(n9193) );
  NAND2_X1 U7785 ( .A1(n6146), .A2(n9193), .ZN(n6147) );
  AOI22_X1 U7786 ( .A1(n8918), .A2(n6241), .B1(n6290), .B2(n8894), .ZN(n6149)
         );
  NAND2_X1 U7787 ( .A1(n6150), .A2(n6149), .ZN(P1_U3230) );
  INV_X1 U7788 ( .A(n6151), .ZN(n6153) );
  NAND2_X2 U7789 ( .A1(n6237), .A2(n6152), .ZN(n7799) );
  NAND2_X1 U7790 ( .A1(n6153), .A2(n7799), .ZN(n6155) );
  INV_X1 U7791 ( .A(n6215), .ZN(n6157) );
  NAND2_X1 U7792 ( .A1(n6157), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7793 ( .A1(n6241), .A2(n6167), .ZN(n6165) );
  XNOR2_X1 U7794 ( .A(n6172), .B(n6170), .ZN(n8825) );
  NAND2_X1 U7795 ( .A1(n7801), .A2(n6241), .ZN(n6169) );
  NAND2_X1 U7796 ( .A1(n4256), .A2(n6163), .ZN(n6168) );
  AND2_X1 U7797 ( .A1(n6169), .A2(n6168), .ZN(n8826) );
  NAND2_X1 U7798 ( .A1(n8825), .A2(n8826), .ZN(n8824) );
  INV_X1 U7799 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7800 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7801 ( .A1(n8824), .A2(n6173), .ZN(n6207) );
  INV_X1 U7802 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6175) );
  INV_X1 U7803 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6174) );
  OAI22_X1 U7804 ( .A1(n4272), .A2(n6175), .B1(n6227), .B2(n6174), .ZN(n6179)
         );
  INV_X1 U7805 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6177) );
  INV_X1 U7806 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6176) );
  OAI22_X1 U7807 ( .A1(n4276), .A2(n6177), .B1(n6230), .B2(n6176), .ZN(n6178)
         );
  NAND2_X1 U7808 ( .A1(n9629), .A2(n6167), .ZN(n6186) );
  OR2_X1 U7809 ( .A1(n6213), .A2(n6180), .ZN(n6182) );
  OAI211_X1 U7810 ( .C1(n7569), .C2(n6183), .A(n6182), .B(n4867), .ZN(n6184)
         );
  NAND2_X1 U7811 ( .A1(n9651), .A2(n7793), .ZN(n6185) );
  NAND2_X1 U7812 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  INV_X1 U7813 ( .A(n7799), .ZN(n6222) );
  XNOR2_X1 U7814 ( .A(n6187), .B(n6222), .ZN(n6210) );
  NAND2_X1 U7815 ( .A1(n7801), .A2(n9629), .ZN(n6189) );
  NAND2_X1 U7816 ( .A1(n4256), .A2(n9651), .ZN(n6188) );
  NAND2_X1 U7817 ( .A1(n6189), .A2(n6188), .ZN(n6208) );
  XNOR2_X1 U7818 ( .A(n6210), .B(n6208), .ZN(n6206) );
  XOR2_X1 U7819 ( .A(n4261), .B(n6206), .Z(n6198) );
  INV_X1 U7820 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6190) );
  OAI22_X1 U7821 ( .A1(n4272), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n6227), .B2(
        n6190), .ZN(n6194) );
  INV_X1 U7822 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6192) );
  INV_X1 U7823 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6191) );
  OAI22_X1 U7824 ( .A1(n4276), .A2(n6192), .B1(n6230), .B2(n6191), .ZN(n6193)
         );
  AOI22_X1 U7825 ( .A1(n8918), .A2(n8935), .B1(n9651), .B2(n8894), .ZN(n6197)
         );
  AOI22_X1 U7826 ( .A1(n8901), .A2(n6241), .B1(n8828), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6196) );
  OAI211_X1 U7827 ( .C1(n6198), .C2(n8923), .A(n6197), .B(n6196), .ZN(P1_U3235) );
  AND3_X1 U7828 ( .A1(n6200), .A2(n6199), .A3(n7042), .ZN(n6202) );
  NAND2_X1 U7829 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  NAND2_X1 U7830 ( .A1(n6203), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7831 ( .A1(n6205), .A2(n6204), .ZN(n8907) );
  INV_X1 U7832 ( .A(n8907), .ZN(n8920) );
  NAND2_X1 U7833 ( .A1(n6207), .A2(n6206), .ZN(n6212) );
  INV_X1 U7834 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7835 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7836 ( .A1(n8935), .A2(n4256), .ZN(n6221) );
  OR2_X1 U7837 ( .A1(n6213), .A2(n6214), .ZN(n6218) );
  OR2_X1 U7838 ( .A1(n7957), .A2(n6216), .ZN(n6217) );
  OAI211_X1 U7839 ( .C1(n4274), .C2(n6219), .A(n6218), .B(n6217), .ZN(n6629)
         );
  NAND2_X1 U7840 ( .A1(n6629), .A2(n7793), .ZN(n6220) );
  NAND2_X1 U7841 ( .A1(n6221), .A2(n6220), .ZN(n6223) );
  XNOR2_X1 U7842 ( .A(n6223), .B(n6222), .ZN(n6297) );
  NAND2_X1 U7843 ( .A1(n7801), .A2(n8935), .ZN(n6225) );
  NAND2_X1 U7844 ( .A1(n7824), .A2(n6629), .ZN(n6224) );
  NAND2_X1 U7845 ( .A1(n6225), .A2(n6224), .ZN(n6295) );
  XNOR2_X1 U7846 ( .A(n6294), .B(n6293), .ZN(n6226) );
  NAND2_X1 U7847 ( .A1(n6226), .A2(n8898), .ZN(n6236) );
  INV_X1 U7848 ( .A(n8901), .ZN(n8916) );
  INV_X1 U7849 ( .A(n9629), .ZN(n8076) );
  INV_X1 U7850 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6229) );
  INV_X1 U7851 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6228) );
  OAI22_X1 U7852 ( .A1(n4276), .A2(n6229), .B1(n7848), .B2(n6228), .ZN(n6232)
         );
  XNOR2_X1 U7853 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6778) );
  INV_X1 U7854 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6779) );
  OAI22_X1 U7855 ( .A1(n4272), .A2(n6778), .B1(n7636), .B2(n6779), .ZN(n6231)
         );
  OAI22_X1 U7856 ( .A1(n8916), .A2(n8076), .B1(n6717), .B2(n8904), .ZN(n6233)
         );
  AOI211_X1 U7857 ( .C1(n6629), .C2(n8894), .A(n6234), .B(n6233), .ZN(n6235)
         );
  OAI211_X1 U7858 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8920), .A(n6236), .B(
        n6235), .ZN(P1_U3216) );
  OR2_X1 U7859 ( .A1(n6237), .A2(n6658), .ZN(n6240) );
  OR2_X1 U7860 ( .A1(n6238), .A2(n8062), .ZN(n6239) );
  AND2_X1 U7861 ( .A1(n6240), .A2(n6239), .ZN(n9656) );
  NAND2_X1 U7862 ( .A1(n4448), .A2(n8111), .ZN(n9682) );
  NAND2_X1 U7863 ( .A1(n6243), .A2(n6242), .ZN(n6628) );
  OAI21_X1 U7864 ( .B1(n6242), .B2(n6243), .A(n6628), .ZN(n6793) );
  NAND2_X1 U7865 ( .A1(n6075), .A2(n9193), .ZN(n6246) );
  NAND2_X1 U7866 ( .A1(n6103), .A2(n6244), .ZN(n6245) );
  INV_X1 U7867 ( .A(n9632), .ZN(n9451) );
  NOR2_X1 U7868 ( .A1(n8937), .A2(n8071), .ZN(n6247) );
  OAI21_X1 U7869 ( .B1(n7979), .B2(n6247), .A(n6660), .ZN(n6248) );
  INV_X1 U7870 ( .A(n9289), .ZN(n9628) );
  INV_X1 U7871 ( .A(n9287), .ZN(n9630) );
  AOI222_X1 U7872 ( .A1(n9451), .A2(n6248), .B1(n9629), .B2(n9628), .C1(n8937), 
        .C2(n9630), .ZN(n6784) );
  INV_X1 U7873 ( .A(n9458), .ZN(n9640) );
  NAND2_X1 U7874 ( .A1(n6163), .A2(n6290), .ZN(n6249) );
  NAND3_X1 U7875 ( .A1(n9640), .A2(n7019), .A3(n6249), .ZN(n6786) );
  INV_X1 U7876 ( .A(n6786), .ZN(n6250) );
  AOI21_X1 U7877 ( .B1(n9679), .B2(n6163), .A(n6250), .ZN(n6251) );
  OAI211_X1 U7878 ( .C1(n9373), .C2(n6793), .A(n6784), .B(n6251), .ZN(n6258)
         );
  NAND2_X1 U7879 ( .A1(n6258), .A2(n9709), .ZN(n6252) );
  OAI21_X1 U7880 ( .B1(n9709), .B2(n6104), .A(n6252), .ZN(P1_U3457) );
  INV_X1 U7881 ( .A(n6253), .ZN(n6254) );
  NOR2_X1 U7882 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  AND2_X2 U7883 ( .A1(n6257), .A2(n6256), .ZN(n9721) );
  INV_X1 U7884 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7885 ( .A1(n6258), .A2(n9721), .ZN(n6259) );
  OAI21_X1 U7886 ( .B1(n9721), .B2(n6260), .A(n6259), .ZN(P1_U3524) );
  NOR2_X1 U7887 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6640), .ZN(n6261) );
  AOI21_X1 U7888 ( .B1(n6640), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6261), .ZN(
        n8947) );
  NOR2_X1 U7889 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6276), .ZN(n6262) );
  AOI21_X1 U7890 ( .B1(n6276), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6262), .ZN(
        n9535) );
  AOI21_X1 U7891 ( .B1(n6275), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6263), .ZN(
        n9521) );
  NOR2_X1 U7892 ( .A1(n9523), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6264) );
  AOI21_X1 U7893 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9523), .A(n6264), .ZN(
        n9520) );
  NAND2_X1 U7894 ( .A1(n9521), .A2(n9520), .ZN(n9519) );
  OAI21_X1 U7895 ( .B1(n9523), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9519), .ZN(
        n9534) );
  NAND2_X1 U7896 ( .A1(n9535), .A2(n9534), .ZN(n9533) );
  OAI21_X1 U7897 ( .B1(n6276), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9533), .ZN(
        n9554) );
  INV_X1 U7898 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6265) );
  MUX2_X1 U7899 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6265), .S(n6542), .Z(n6266)
         );
  INV_X1 U7900 ( .A(n6266), .ZN(n9553) );
  NOR2_X1 U7901 ( .A1(n9554), .A2(n9553), .ZN(n9552) );
  INV_X1 U7902 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U7903 ( .A1(n6645), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9943), .B2(
        n6267), .ZN(n6268) );
  OAI21_X1 U7904 ( .B1(n6269), .B2(n6268), .A(n6409), .ZN(n6281) );
  INV_X1 U7905 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6271) );
  INV_X1 U7906 ( .A(n9613), .ZN(n9593) );
  INV_X1 U7907 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6650) );
  NOR2_X1 U7908 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6650), .ZN(n7130) );
  AOI21_X1 U7909 ( .B1(n9593), .B2(n6645), .A(n7130), .ZN(n6270) );
  OAI21_X1 U7910 ( .B1(n9605), .B2(n6271), .A(n6270), .ZN(n6280) );
  INV_X1 U7911 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U7912 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6640), .B1(n8938), .B2(
        n9994), .ZN(n8943) );
  NAND2_X1 U7913 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6276), .ZN(n6272) );
  OAI21_X1 U7914 ( .B1(n6276), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6272), .ZN(
        n9538) );
  NOR2_X1 U7915 ( .A1(n9523), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6273) );
  AOI21_X1 U7916 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9523), .A(n6273), .ZN(
        n9526) );
  AOI21_X1 U7917 ( .B1(n6275), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6274), .ZN(
        n9525) );
  NAND2_X1 U7918 ( .A1(n9526), .A2(n9525), .ZN(n9524) );
  OAI21_X1 U7919 ( .B1(n9523), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9524), .ZN(
        n9539) );
  NOR2_X1 U7920 ( .A1(n9538), .A2(n9539), .ZN(n9537) );
  INV_X1 U7921 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U7922 ( .A1(n6542), .A2(P1_REG1_REG_6__SCAN_IN), .B1(n9714), .B2(
        n9559), .ZN(n9550) );
  NAND2_X1 U7923 ( .A1(n9551), .A2(n9550), .ZN(n9549) );
  OAI21_X1 U7924 ( .B1(n6542), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9549), .ZN(
        n8942) );
  NAND2_X1 U7925 ( .A1(n8943), .A2(n8942), .ZN(n8941) );
  OAI21_X1 U7926 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6640), .A(n8941), .ZN(
        n6278) );
  INV_X1 U7927 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U7928 ( .A(n6649), .B(P1_REG1_REG_8__SCAN_IN), .S(n6645), .Z(n6277)
         );
  NOR2_X1 U7929 ( .A1(n6277), .A2(n6278), .ZN(n6401) );
  AOI211_X1 U7930 ( .C1(n6278), .C2(n6277), .A(n6401), .B(n9536), .ZN(n6279)
         );
  AOI211_X1 U7931 ( .C1(n9609), .C2(n6281), .A(n6280), .B(n6279), .ZN(n6282)
         );
  INV_X1 U7932 ( .A(n6282), .ZN(P1_U3249) );
  NAND2_X1 U7933 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  NAND2_X2 U7934 ( .A1(n6285), .A2(n9635), .ZN(n10029) );
  INV_X2 U7935 ( .A(n10029), .ZN(n9648) );
  OR2_X1 U7936 ( .A1(n6285), .A2(n9193), .ZN(n10037) );
  OAI22_X1 U7937 ( .A1(n10037), .A2(n6286), .B1(n6673), .B2(n6285), .ZN(n6289)
         );
  OAI22_X1 U7938 ( .A1(n10029), .A2(n10011), .B1(n6287), .B2(n9635), .ZN(n6288) );
  AOI21_X1 U7939 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6291) );
  OAI21_X1 U7940 ( .B1(n9648), .B2(n6292), .A(n6291), .ZN(P1_U3291) );
  NAND2_X1 U7941 ( .A1(n6294), .A2(n6293), .ZN(n6299) );
  INV_X1 U7942 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7943 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  NAND2_X1 U7944 ( .A1(n9627), .A2(n7824), .ZN(n6306) );
  OR2_X1 U7945 ( .A1(n6213), .A2(n6300), .ZN(n6303) );
  OR2_X1 U7946 ( .A1(n7957), .A2(n6301), .ZN(n6302) );
  NAND2_X1 U7947 ( .A1(n9666), .A2(n7793), .ZN(n6305) );
  NAND2_X1 U7948 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  XNOR2_X1 U7949 ( .A(n6307), .B(n7822), .ZN(n6482) );
  NAND2_X1 U7950 ( .A1(n7801), .A2(n9627), .ZN(n6309) );
  NAND2_X1 U7951 ( .A1(n7824), .A2(n9666), .ZN(n6308) );
  AND2_X1 U7952 ( .A1(n6309), .A2(n6308), .ZN(n6481) );
  INV_X1 U7953 ( .A(n6481), .ZN(n6483) );
  XNOR2_X1 U7954 ( .A(n6482), .B(n6483), .ZN(n6310) );
  XNOR2_X1 U7955 ( .A(n6487), .B(n6310), .ZN(n6311) );
  NAND2_X1 U7956 ( .A1(n6311), .A2(n8898), .ZN(n6322) );
  AND2_X1 U7957 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9528) );
  INV_X1 U7958 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6313) );
  INV_X1 U7959 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6312) );
  OAI22_X1 U7960 ( .A1(n4276), .A2(n6313), .B1(n7848), .B2(n6312), .ZN(n6319)
         );
  INV_X1 U7961 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7962 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6314) );
  NAND2_X1 U7963 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U7964 ( .A1(n6497), .A2(n6316), .ZN(n6718) );
  INV_X1 U7965 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6317) );
  OAI22_X1 U7966 ( .A1(n4272), .A2(n6718), .B1(n7636), .B2(n6317), .ZN(n6318)
         );
  INV_X1 U7967 ( .A(n8934), .ZN(n6893) );
  OAI22_X1 U7968 ( .A1(n8916), .A2(n6774), .B1(n6893), .B2(n8904), .ZN(n6320)
         );
  AOI211_X1 U7969 ( .C1(n9666), .C2(n8894), .A(n9528), .B(n6320), .ZN(n6321)
         );
  OAI211_X1 U7970 ( .C1(n8920), .C2(n6778), .A(n6322), .B(n6321), .ZN(P1_U3228) );
  INV_X1 U7971 ( .A(n7567), .ZN(n6326) );
  NAND2_X1 U7972 ( .A1(n6323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6325) );
  INV_X1 U7973 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6324) );
  XNOR2_X1 U7974 ( .A(n6325), .B(n6324), .ZN(n8958) );
  OAI222_X1 U7975 ( .A1(n8121), .A2(n7568), .B1(n9402), .B2(n6326), .C1(
        P1_U3084), .C2(n8958), .ZN(P1_U3338) );
  OAI222_X1 U7976 ( .A1(n7376), .A2(n6327), .B1(n8783), .B2(n6326), .C1(
        P2_U3152), .C2(n7464), .ZN(P2_U3343) );
  INV_X1 U7977 ( .A(n7590), .ZN(n6332) );
  INV_X1 U7978 ( .A(n8340), .ZN(n7479) );
  OAI222_X1 U7979 ( .A1(n7376), .A2(n6328), .B1(n8783), .B2(n6332), .C1(n7479), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  NOR2_X1 U7980 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6329) );
  NAND2_X1 U7981 ( .A1(n6330), .A2(n6329), .ZN(n6334) );
  NAND2_X1 U7982 ( .A1(n6334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6331) );
  XNOR2_X1 U7983 ( .A(n6331), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8975) );
  INV_X1 U7984 ( .A(n8975), .ZN(n8965) );
  OAI222_X1 U7985 ( .A1(n8121), .A2(n6333), .B1(n8965), .B2(P1_U3084), .C1(
        n9402), .C2(n6332), .ZN(P1_U3337) );
  INV_X1 U7986 ( .A(n7608), .ZN(n6341) );
  OR2_X1 U7987 ( .A1(n6334), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7988 ( .A1(n6335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7989 ( .A1(n6337), .A2(n6336), .ZN(n6523) );
  OR2_X1 U7990 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  AOI22_X1 U7991 ( .A1(n8987), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6339), .ZN(n6340) );
  OAI21_X1 U7992 ( .B1(n6341), .B2(n9402), .A(n6340), .ZN(P1_U3336) );
  OAI222_X1 U7993 ( .A1(n7376), .A2(n6342), .B1(n8783), .B2(n6341), .C1(n8350), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U7994 ( .A1(n8297), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6349) );
  MUX2_X1 U7995 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6343), .S(n8297), .Z(n8294)
         );
  INV_X1 U7996 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9931) );
  MUX2_X1 U7997 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9931), .S(n9423), .Z(n9426)
         );
  NAND2_X1 U7998 ( .A1(n9410), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6347) );
  INV_X1 U7999 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6345) );
  MUX2_X1 U8000 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6345), .S(n6344), .Z(n6346)
         );
  INV_X1 U8001 ( .A(n6346), .ZN(n9412) );
  NAND3_X1 U8002 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9412), .ZN(n9411) );
  NAND2_X1 U8003 ( .A1(n6347), .A2(n9411), .ZN(n9427) );
  NAND2_X1 U8004 ( .A1(n9426), .A2(n9427), .ZN(n9425) );
  OAI21_X1 U8005 ( .B1(n6348), .B2(n9931), .A(n9425), .ZN(n8293) );
  NAND2_X1 U8006 ( .A1(n8294), .A2(n8293), .ZN(n8292) );
  AND2_X1 U8007 ( .A1(n6349), .A2(n8292), .ZN(n6357) );
  MUX2_X1 U8008 ( .A(n5066), .B(P2_REG2_REG_4__SCAN_IN), .S(n6428), .Z(n6356)
         );
  NOR2_X1 U8009 ( .A1(n6357), .A2(n6356), .ZN(n6427) );
  NAND2_X1 U8010 ( .A1(n6350), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7502) );
  OR2_X1 U8011 ( .A1(n6351), .A2(n7502), .ZN(n6352) );
  OAI211_X1 U8012 ( .C1(n9767), .C2(n6353), .A(n7040), .B(n6352), .ZN(n6355)
         );
  NAND2_X1 U8013 ( .A1(n6355), .A2(n6354), .ZN(n6367) );
  INV_X2 U8014 ( .A(P2_U3966), .ZN(n8291) );
  NAND2_X1 U8015 ( .A1(n6367), .A2(n8291), .ZN(n6358) );
  INV_X1 U8016 ( .A(n6368), .ZN(n7437) );
  NAND2_X1 U8017 ( .A1(n6358), .A2(n7437), .ZN(n9727) );
  OR2_X1 U8018 ( .A1(n9727), .A2(n6359), .ZN(n8370) );
  AOI211_X1 U8019 ( .C1(n6357), .C2(n6356), .A(n6427), .B(n8370), .ZN(n6376)
         );
  AND2_X1 U8020 ( .A1(n6359), .A2(n6358), .ZN(n9424) );
  NAND2_X1 U8021 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6534) );
  INV_X1 U8022 ( .A(n6534), .ZN(n6360) );
  AOI21_X1 U8023 ( .B1(n9417), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6360), .ZN(
        n6373) );
  XNOR2_X1 U8024 ( .A(n6428), .B(n6361), .ZN(n6371) );
  NAND2_X1 U8025 ( .A1(n8297), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8026 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9408) );
  NAND2_X1 U8027 ( .A1(n9410), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6362) );
  OAI21_X1 U8028 ( .B1(n9410), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6362), .ZN(
        n9407) );
  NOR2_X1 U8029 ( .A1(n9408), .A2(n9407), .ZN(n9406) );
  AOI21_X1 U8030 ( .B1(n9410), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9406), .ZN(
        n9421) );
  NAND2_X1 U8031 ( .A1(n9423), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8032 ( .B1(n9423), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6363), .ZN(
        n9420) );
  NOR2_X1 U8033 ( .A1(n9421), .A2(n9420), .ZN(n9419) );
  AOI21_X1 U8034 ( .B1(n9423), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9419), .ZN(
        n8300) );
  OR2_X1 U8035 ( .A1(n8297), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8036 ( .A1(n6364), .A2(n6366), .ZN(n8299) );
  NOR2_X1 U8037 ( .A1(n8300), .A2(n8299), .ZN(n8298) );
  INV_X1 U8038 ( .A(n8298), .ZN(n6365) );
  NAND2_X1 U8039 ( .A1(n6366), .A2(n6365), .ZN(n6370) );
  INV_X1 U8040 ( .A(n6367), .ZN(n6369) );
  NAND2_X1 U8041 ( .A1(n6369), .A2(n6368), .ZN(n9418) );
  NAND2_X1 U8042 ( .A1(n6371), .A2(n6370), .ZN(n6419) );
  OAI211_X1 U8043 ( .C1(n6371), .C2(n6370), .A(n9724), .B(n6419), .ZN(n6372)
         );
  OAI211_X1 U8044 ( .C1(n9726), .C2(n6374), .A(n6373), .B(n6372), .ZN(n6375)
         );
  OR2_X1 U8045 ( .A1(n6376), .A2(n6375), .ZN(P2_U3249) );
  NAND2_X1 U8046 ( .A1(n8291), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6377) );
  OAI21_X1 U8047 ( .B1(n6378), .B2(n8291), .A(n6377), .ZN(P2_U3581) );
  INV_X1 U8048 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7189) );
  INV_X1 U8049 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7575) );
  INV_X1 U8050 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8857) );
  INV_X1 U8051 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10001) );
  INV_X1 U8052 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7693) );
  INV_X1 U8053 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9958) );
  INV_X1 U8054 ( .A(n7757), .ZN(n6390) );
  INV_X1 U8055 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8903) );
  INV_X1 U8056 ( .A(n7811), .ZN(n6392) );
  AND2_X1 U8057 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6391) );
  NAND2_X1 U8058 ( .A1(n6392), .A2(n6391), .ZN(n9074) );
  OR2_X1 U8059 ( .A1(n9074), .A2(n4272), .ZN(n6398) );
  INV_X1 U8060 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8061 ( .A1(n7853), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8062 ( .A1(n7813), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6393) );
  OAI211_X1 U8063 ( .C1(n7852), .C2(n6395), .A(n6394), .B(n6393), .ZN(n6396)
         );
  INV_X1 U8064 ( .A(n6396), .ZN(n6397) );
  INV_X2 U8065 ( .A(P1_U4006), .ZN(n8936) );
  NAND2_X1 U8066 ( .A1(n8936), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6399) );
  OAI21_X1 U8067 ( .B1(n9085), .B2(n8936), .A(n6399), .ZN(P1_U3584) );
  INV_X1 U8068 ( .A(n9536), .ZN(n9620) );
  INV_X1 U8069 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9482) );
  AOI22_X1 U8070 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9592), .B1(n6400), .B2(
        n9482), .ZN(n9596) );
  INV_X1 U8071 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U8072 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6863), .B1(n9585), .B2(
        n6985), .ZN(n9577) );
  NOR2_X1 U8073 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9572), .ZN(n6402) );
  AOI21_X1 U8074 ( .B1(n9572), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6402), .ZN(
        n9564) );
  NAND2_X1 U8075 ( .A1(n9565), .A2(n9564), .ZN(n9563) );
  OAI21_X1 U8076 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9572), .A(n9563), .ZN(
        n9576) );
  NAND2_X1 U8077 ( .A1(n9577), .A2(n9576), .ZN(n9575) );
  OAI21_X1 U8078 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6863), .A(n9575), .ZN(
        n9595) );
  INV_X1 U8079 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7005) );
  MUX2_X1 U8080 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7005), .S(n7181), .Z(n6403)
         );
  NAND2_X1 U8081 ( .A1(n6403), .A2(n6404), .ZN(n6617) );
  OAI21_X1 U8082 ( .B1(n6404), .B2(n6403), .A(n6617), .ZN(n6416) );
  INV_X1 U8083 ( .A(n9605), .ZN(n9619) );
  NAND2_X1 U8084 ( .A1(n9619), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8085 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7366) );
  OAI211_X1 U8086 ( .C1(n9613), .C2(n6406), .A(n6405), .B(n7366), .ZN(n6415)
         );
  NOR2_X1 U8087 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9592), .ZN(n6407) );
  AOI21_X1 U8088 ( .B1(n9592), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6407), .ZN(
        n9599) );
  NAND2_X1 U8089 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9572), .ZN(n6408) );
  OAI21_X1 U8090 ( .B1(n9572), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6408), .ZN(
        n9567) );
  OAI21_X1 U8091 ( .B1(n6645), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6409), .ZN(
        n9568) );
  NOR2_X1 U8092 ( .A1(n9567), .A2(n9568), .ZN(n9566) );
  NAND2_X1 U8093 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6863), .ZN(n6410) );
  OAI21_X1 U8094 ( .B1(n6863), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6410), .ZN(
        n9580) );
  OAI21_X1 U8095 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9592), .A(n9597), .ZN(
        n6413) );
  NAND2_X1 U8096 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7181), .ZN(n6411) );
  OAI21_X1 U8097 ( .B1(n7181), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6411), .ZN(
        n6412) );
  NOR2_X1 U8098 ( .A1(n6412), .A2(n6413), .ZN(n6611) );
  AOI211_X1 U8099 ( .C1(n6413), .C2(n6412), .A(n6611), .B(n9578), .ZN(n6414)
         );
  AOI211_X1 U8100 ( .C1(n9620), .C2(n6416), .A(n6415), .B(n6414), .ZN(n6417)
         );
  INV_X1 U8101 ( .A(n6417), .ZN(P1_U3253) );
  NAND2_X1 U8102 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6576) );
  INV_X1 U8103 ( .A(n6576), .ZN(n6426) );
  NAND2_X1 U8104 ( .A1(n6428), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8105 ( .A1(n6419), .A2(n6418), .ZN(n8314) );
  OR2_X1 U8106 ( .A1(n8311), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8107 ( .A1(n8311), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6420) );
  AND2_X1 U8108 ( .A1(n6421), .A2(n6420), .ZN(n8315) );
  INV_X1 U8109 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6422) );
  MUX2_X1 U8110 ( .A(n6422), .B(P2_REG1_REG_6__SCAN_IN), .S(n6437), .Z(n6423)
         );
  AOI211_X1 U8111 ( .C1(n6424), .C2(n6423), .A(n6436), .B(n9418), .ZN(n6425)
         );
  AOI211_X1 U8112 ( .C1(n9417), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6426), .B(
        n6425), .ZN(n6435) );
  NAND2_X1 U8113 ( .A1(n8311), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6431) );
  AOI21_X1 U8114 ( .B1(n6428), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6427), .ZN(
        n8306) );
  INV_X1 U8115 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6429) );
  MUX2_X1 U8116 ( .A(n6429), .B(P2_REG2_REG_5__SCAN_IN), .S(n8311), .Z(n8307)
         );
  OR2_X1 U8117 ( .A1(n8306), .A2(n8307), .ZN(n6430) );
  NAND2_X1 U8118 ( .A1(n6431), .A2(n6430), .ZN(n6433) );
  MUX2_X1 U8119 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6901), .S(n6437), .Z(n6432)
         );
  NAND2_X1 U8120 ( .A1(n6432), .A2(n6433), .ZN(n6444) );
  OAI211_X1 U8121 ( .C1(n6433), .C2(n6432), .A(n9722), .B(n6444), .ZN(n6434)
         );
  OAI211_X1 U8122 ( .C1(n9726), .C2(n6445), .A(n6435), .B(n6434), .ZN(P2_U3251) );
  AND2_X1 U8123 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6933) );
  NAND2_X1 U8124 ( .A1(n6443), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6438) );
  OAI21_X1 U8125 ( .B1(n6443), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6438), .ZN(
        n6465) );
  NOR2_X1 U8126 ( .A1(n6466), .A2(n6465), .ZN(n6464) );
  INV_X1 U8127 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U8128 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6439), .S(n6458), .Z(n6440)
         );
  NOR2_X1 U8129 ( .A1(n6441), .A2(n6440), .ZN(n6451) );
  AOI211_X1 U8130 ( .C1(n6441), .C2(n6440), .A(n6451), .B(n9418), .ZN(n6442)
         );
  AOI211_X1 U8131 ( .C1(n9417), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6933), .B(
        n6442), .ZN(n6450) );
  MUX2_X1 U8132 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6763), .S(n6443), .Z(n6470)
         );
  OAI21_X1 U8133 ( .B1(n6445), .B2(n6901), .A(n6444), .ZN(n6471) );
  NAND2_X1 U8134 ( .A1(n6470), .A2(n6471), .ZN(n6469) );
  OAI21_X1 U8135 ( .B1(n6474), .B2(n6763), .A(n6469), .ZN(n6448) );
  MUX2_X1 U8136 ( .A(n6446), .B(P2_REG2_REG_8__SCAN_IN), .S(n6458), .Z(n6447)
         );
  NAND2_X1 U8137 ( .A1(n6447), .A2(n6448), .ZN(n6457) );
  OAI211_X1 U8138 ( .C1(n6448), .C2(n6447), .A(n9722), .B(n6457), .ZN(n6449)
         );
  OAI211_X1 U8139 ( .C1(n9726), .C2(n6458), .A(n6450), .B(n6449), .ZN(P2_U3253) );
  NAND2_X1 U8140 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6959) );
  INV_X1 U8141 ( .A(n6959), .ZN(n6456) );
  INV_X1 U8142 ( .A(n6458), .ZN(n6452) );
  MUX2_X1 U8143 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6685), .S(n6686), .Z(n6453)
         );
  NOR2_X1 U8144 ( .A1(n6454), .A2(n6453), .ZN(n6687) );
  AOI211_X1 U8145 ( .C1(n6454), .C2(n6453), .A(n6687), .B(n9418), .ZN(n6455)
         );
  AOI211_X1 U8146 ( .C1(n9417), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6456), .B(
        n6455), .ZN(n6462) );
  OAI21_X1 U8147 ( .B1(n6458), .B2(n6446), .A(n6457), .ZN(n6460) );
  MUX2_X1 U8148 ( .A(n7151), .B(P2_REG2_REG_9__SCAN_IN), .S(n6686), .Z(n6459)
         );
  NAND2_X1 U8149 ( .A1(n6459), .A2(n6460), .ZN(n6682) );
  OAI211_X1 U8150 ( .C1(n6460), .C2(n6459), .A(n9722), .B(n6682), .ZN(n6461)
         );
  OAI211_X1 U8151 ( .C1(n9726), .C2(n6686), .A(n6462), .B(n6461), .ZN(P2_U3254) );
  NOR2_X1 U8152 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6463), .ZN(n6468) );
  AOI211_X1 U8153 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n9418), .ZN(n6467)
         );
  AOI211_X1 U8154 ( .C1(n9417), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6468), .B(
        n6467), .ZN(n6473) );
  OAI211_X1 U8155 ( .C1(n6471), .C2(n6470), .A(n9722), .B(n6469), .ZN(n6472)
         );
  OAI211_X1 U8156 ( .C1(n9726), .C2(n6474), .A(n6473), .B(n6472), .ZN(P2_U3252) );
  NAND2_X1 U8157 ( .A1(n7801), .A2(n8934), .ZN(n6480) );
  OR2_X1 U8158 ( .A1(n6475), .A2(n6213), .ZN(n6478) );
  OR2_X1 U8159 ( .A1(n7957), .A2(n6476), .ZN(n6477) );
  OAI211_X1 U8160 ( .C1(n7569), .C2(n9543), .A(n6478), .B(n6477), .ZN(n6501)
         );
  NAND2_X1 U8161 ( .A1(n7824), .A2(n6501), .ZN(n6479) );
  AND2_X1 U8162 ( .A1(n6480), .A2(n6479), .ZN(n6494) );
  AND2_X1 U8163 ( .A1(n6482), .A2(n6481), .ZN(n6486) );
  INV_X1 U8164 ( .A(n6482), .ZN(n6484) );
  NAND2_X1 U8165 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8166 ( .A1(n8934), .A2(n7824), .ZN(n6490) );
  NAND2_X1 U8167 ( .A1(n6501), .A2(n7808), .ZN(n6489) );
  NAND2_X1 U8168 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  XNOR2_X1 U8169 ( .A(n6491), .B(n7799), .ZN(n6492) );
  OAI21_X1 U8170 ( .B1(n6494), .B2(n4356), .A(n6540), .ZN(n6495) );
  NAND2_X1 U8171 ( .A1(n6495), .A2(n8898), .ZN(n6504) );
  INV_X1 U8172 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6496) );
  OAI22_X1 U8173 ( .A1(n4276), .A2(n9714), .B1(n7848), .B2(n6496), .ZN(n6500)
         );
  INV_X1 U8174 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8175 ( .A1(n6497), .A2(n6561), .ZN(n6498) );
  NAND2_X1 U8176 ( .A1(n6555), .A2(n6498), .ZN(n6562) );
  OAI22_X1 U8177 ( .A1(n4272), .A2(n6562), .B1(n7636), .B2(n6265), .ZN(n6499)
         );
  AND2_X1 U8178 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9541) );
  INV_X1 U8179 ( .A(n8894), .ZN(n8910) );
  OAI22_X1 U8180 ( .A1(n8916), .A2(n6717), .B1(n9675), .B2(n8910), .ZN(n6502)
         );
  AOI211_X1 U8181 ( .C1(n8918), .C2(n8933), .A(n9541), .B(n6502), .ZN(n6503)
         );
  OAI211_X1 U8182 ( .C1(n8920), .C2(n6718), .A(n6504), .B(n6503), .ZN(P1_U3225) );
  NOR2_X1 U8183 ( .A1(n8244), .A2(n7525), .ZN(n8256) );
  AOI22_X1 U8184 ( .A1(n8256), .A2(n8290), .B1(n5866), .B2(n5761), .ZN(n6507)
         );
  NOR2_X1 U8185 ( .A1(n6507), .A2(n6506), .ZN(n6511) );
  OAI22_X1 U8186 ( .A1(n8234), .A2(n6847), .B1(n9789), .B2(n8270), .ZN(n6510)
         );
  NOR2_X1 U8187 ( .A1(n8266), .A2(P2_U3152), .ZN(n6575) );
  INV_X1 U8188 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6852) );
  OAI22_X1 U8189 ( .A1(n8233), .A2(n5042), .B1(n6575), .B2(n6852), .ZN(n6509)
         );
  AOI211_X1 U8190 ( .C1(n6511), .C2(n6508), .A(n6510), .B(n6509), .ZN(n6512)
         );
  OAI21_X1 U8191 ( .B1(n6513), .B2(n8244), .A(n6512), .ZN(P2_U3239) );
  OAI21_X1 U8192 ( .B1(n6515), .B2(n6514), .A(n6508), .ZN(n6520) );
  OAI22_X1 U8193 ( .A1(n8234), .A2(n6516), .B1(n9784), .B2(n8270), .ZN(n6519)
         );
  INV_X1 U8194 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6517) );
  OAI22_X1 U8195 ( .A1(n8233), .A2(n6570), .B1(n6575), .B2(n6517), .ZN(n6518)
         );
  AOI211_X1 U8196 ( .C1(n5866), .C2(n6520), .A(n6519), .B(n6518), .ZN(n6521)
         );
  INV_X1 U8197 ( .A(n6521), .ZN(P2_U3224) );
  INV_X1 U8198 ( .A(n7627), .ZN(n6525) );
  OAI222_X1 U8199 ( .A1(n7376), .A2(n6522), .B1(n8783), .B2(n6525), .C1(
        P2_U3152), .C2(n8357), .ZN(P2_U3340) );
  INV_X1 U8200 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8201 ( .A1(n6523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6524) );
  XNOR2_X1 U8202 ( .A(n6524), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8988) );
  INV_X1 U8203 ( .A(n8988), .ZN(n9614) );
  OAI222_X1 U8204 ( .A1(n8121), .A2(n6526), .B1(n9402), .B2(n6525), .C1(
        P1_U3084), .C2(n9614), .ZN(P1_U3335) );
  NAND2_X1 U8205 ( .A1(n6529), .A2(n6528), .ZN(n8134) );
  OAI21_X1 U8206 ( .B1(n6527), .B2(n6529), .A(n8134), .ZN(n6538) );
  INV_X1 U8207 ( .A(n6527), .ZN(n6531) );
  NAND3_X1 U8208 ( .A1(n8256), .A2(n6531), .A3(n6530), .ZN(n6532) );
  AOI21_X1 U8209 ( .B1(n8233), .B2(n6532), .A(n6847), .ZN(n6537) );
  AOI22_X1 U8210 ( .A1(n8198), .A2(n9741), .B1(n6533), .B2(n8238), .ZN(n6535)
         );
  OAI211_X1 U8211 ( .C1(n9756), .C2(n8251), .A(n6535), .B(n6534), .ZN(n6536)
         );
  AOI211_X1 U8212 ( .C1(n5866), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6539)
         );
  INV_X1 U8213 ( .A(n6539), .ZN(P2_U3232) );
  INV_X2 U8214 ( .A(n6213), .ZN(n6643) );
  AOI22_X1 U8215 ( .A1(n7649), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7648), .B2(
        n6542), .ZN(n6543) );
  NAND2_X1 U8216 ( .A1(n9678), .A2(n7808), .ZN(n6545) );
  NAND2_X1 U8217 ( .A1(n8933), .A2(n7824), .ZN(n6544) );
  NAND2_X1 U8218 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  XNOR2_X1 U8219 ( .A(n6546), .B(n7822), .ZN(n6552) );
  INV_X1 U8220 ( .A(n6552), .ZN(n6550) );
  NAND2_X1 U8221 ( .A1(n7801), .A2(n8933), .ZN(n6548) );
  NAND2_X1 U8222 ( .A1(n9678), .A2(n7824), .ZN(n6547) );
  AND2_X1 U8223 ( .A1(n6548), .A2(n6547), .ZN(n6551) );
  INV_X1 U8224 ( .A(n6551), .ZN(n6549) );
  AND2_X1 U8225 ( .A1(n6552), .A2(n6551), .ZN(n6797) );
  NOR2_X1 U8226 ( .A1(n4357), .A2(n6797), .ZN(n6553) );
  XNOR2_X1 U8227 ( .A(n4264), .B(n6553), .ZN(n6568) );
  INV_X1 U8228 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8229 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  AND2_X1 U8230 ( .A1(n6651), .A2(n6556), .ZN(n6804) );
  NAND2_X1 U8231 ( .A1(n7797), .A2(n6804), .ZN(n6560) );
  NAND2_X1 U8232 ( .A1(n7633), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8233 ( .A1(n7813), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8234 ( .A1(n7853), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6557) );
  NAND4_X1 U8235 ( .A1(n6560), .A2(n6559), .A3(n6558), .A4(n6557), .ZN(n8932)
         );
  NOR2_X1 U8236 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6561), .ZN(n9556) );
  AOI21_X1 U8237 ( .B1(n8918), .B2(n8932), .A(n9556), .ZN(n6566) );
  INV_X1 U8238 ( .A(n6562), .ZN(n6889) );
  NAND2_X1 U8239 ( .A1(n8907), .A2(n6889), .ZN(n6565) );
  NAND2_X1 U8240 ( .A1(n8894), .A2(n9678), .ZN(n6564) );
  NAND2_X1 U8241 ( .A1(n8901), .A2(n8934), .ZN(n6563) );
  NAND4_X1 U8242 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .ZN(n6567)
         );
  AOI21_X1 U8243 ( .B1(n6568), .B2(n8898), .A(n6567), .ZN(n6569) );
  INV_X1 U8244 ( .A(n6569), .ZN(P1_U3237) );
  INV_X1 U8245 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9729) );
  INV_X1 U8246 ( .A(n8256), .ZN(n8242) );
  OAI22_X1 U8247 ( .A1(n8242), .A2(n6570), .B1(n9776), .B2(n8244), .ZN(n6572)
         );
  NAND2_X1 U8248 ( .A1(n6572), .A2(n6571), .ZN(n6574) );
  AOI22_X1 U8249 ( .A1(n8198), .A2(n8290), .B1(n6595), .B2(n8238), .ZN(n6573)
         );
  OAI211_X1 U8250 ( .C1(n6575), .C2(n9729), .A(n6574), .B(n6573), .ZN(P2_U3234) );
  OAI21_X1 U8251 ( .B1(n8251), .B2(n6902), .A(n6576), .ZN(n6578) );
  OAI22_X1 U8252 ( .A1(n8233), .A2(n6837), .B1(n6903), .B2(n8270), .ZN(n6577)
         );
  AOI211_X1 U8253 ( .C1(n8198), .C2(n8287), .A(n6578), .B(n6577), .ZN(n6585)
         );
  INV_X1 U8254 ( .A(n6580), .ZN(n6583) );
  OAI22_X1 U8255 ( .A1(n8242), .A2(n6837), .B1(n6581), .B2(n8244), .ZN(n6582)
         );
  NAND3_X1 U8256 ( .A1(n8137), .A2(n6583), .A3(n6582), .ZN(n6584) );
  OAI211_X1 U8257 ( .C1(n6586), .C2(n8244), .A(n6585), .B(n6584), .ZN(P2_U3241) );
  NAND3_X1 U8258 ( .A1(n6589), .A2(n6588), .A3(n6587), .ZN(n6761) );
  NAND2_X2 U8259 ( .A1(n6761), .A2(n9755), .ZN(n9757) );
  OR2_X1 U8260 ( .A1(n6590), .A2(n8433), .ZN(n6600) );
  NAND2_X1 U8261 ( .A1(n8626), .A2(n6600), .ZN(n6591) );
  INV_X1 U8262 ( .A(n9755), .ZN(n8570) );
  OAI22_X1 U8263 ( .A1(n9778), .A2(n8566), .B1(n5042), .B2(n8619), .ZN(n9780)
         );
  AOI21_X1 U8264 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n8570), .A(n9780), .ZN(
        n6592) );
  MUX2_X1 U8265 ( .A(n5043), .B(n6592), .S(n9757), .Z(n6597) );
  OR2_X1 U8266 ( .A1(n6761), .A2(n6594), .ZN(n7154) );
  INV_X1 U8267 ( .A(n7154), .ZN(n9759) );
  OAI21_X1 U8268 ( .B1(n8609), .B2(n9759), .A(n6595), .ZN(n6596) );
  OAI211_X1 U8269 ( .C1(n9778), .C2(n8584), .A(n6597), .B(n6596), .ZN(P2_U3296) );
  NAND2_X1 U8270 ( .A1(n6598), .A2(n6599), .ZN(n9747) );
  XNOR2_X1 U8271 ( .A(n9747), .B(n6910), .ZN(n9796) );
  INV_X1 U8272 ( .A(n6600), .ZN(n6601) );
  NAND2_X1 U8273 ( .A1(n9757), .A2(n6601), .ZN(n8637) );
  XNOR2_X1 U8274 ( .A(n6602), .B(n6910), .ZN(n6603) );
  NAND2_X1 U8275 ( .A1(n6603), .A2(n9745), .ZN(n6605) );
  INV_X1 U8276 ( .A(n8619), .ZN(n9740) );
  AOI22_X1 U8277 ( .A1(n5095), .A2(n9740), .B1(n9742), .B2(n8289), .ZN(n6604)
         );
  OAI211_X1 U8278 ( .C1(n9796), .C2(n8626), .A(n6605), .B(n6604), .ZN(n9799)
         );
  NAND2_X1 U8279 ( .A1(n9799), .A2(n9757), .ZN(n6610) );
  OAI22_X1 U8280 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n9755), .B1(n6343), .B2(
        n9757), .ZN(n6608) );
  INV_X1 U8281 ( .A(n6851), .ZN(n6606) );
  OAI21_X1 U8282 ( .B1(n6606), .B2(n9797), .A(n9752), .ZN(n9798) );
  NOR2_X1 U8283 ( .A1(n7154), .A2(n9798), .ZN(n6607) );
  AOI211_X1 U8284 ( .C1(n8609), .C2(n5093), .A(n6608), .B(n6607), .ZN(n6609)
         );
  OAI211_X1 U8285 ( .C1(n9796), .C2(n8637), .A(n6610), .B(n6609), .ZN(P2_U3293) );
  INV_X1 U8286 ( .A(n7391), .ZN(n6623) );
  INV_X1 U8287 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6612) );
  MUX2_X1 U8288 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n6612), .S(n7391), .Z(n6613)
         );
  INV_X1 U8289 ( .A(n6613), .ZN(n6614) );
  AOI211_X1 U8290 ( .C1(n6615), .C2(n6614), .A(n7027), .B(n9578), .ZN(n6616)
         );
  AOI21_X1 U8291 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n9619), .A(n6616), .ZN(
        n6622) );
  INV_X1 U8292 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7188) );
  MUX2_X1 U8293 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7188), .S(n7391), .Z(n6619)
         );
  OAI21_X1 U8294 ( .B1(n7181), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6617), .ZN(
        n6618) );
  OAI21_X1 U8295 ( .B1(n6619), .B2(n6618), .A(n7032), .ZN(n6620) );
  AND2_X1 U8296 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7411) );
  AOI21_X1 U8297 ( .B1(n9620), .B2(n6620), .A(n7411), .ZN(n6621) );
  OAI211_X1 U8298 ( .C1(n6623), .C2(n9613), .A(n6622), .B(n6621), .ZN(P1_U3254) );
  INV_X1 U8299 ( .A(n7647), .ZN(n6625) );
  OAI222_X1 U8300 ( .A1(n7376), .A2(n6624), .B1(n8783), .B2(n6625), .C1(
        P2_U3152), .C2(n8433), .ZN(P2_U3339) );
  OAI222_X1 U8301 ( .A1(n8121), .A2(n6626), .B1(n9402), .B2(n6625), .C1(n8994), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  NAND2_X1 U8302 ( .A1(n6241), .A2(n6163), .ZN(n6627) );
  OAI22_X1 U8303 ( .A1(n7023), .A2(n7978), .B1(n9651), .B2(n9629), .ZN(n9624)
         );
  NAND2_X1 U8304 ( .A1(n6774), .A2(n6629), .ZN(n8081) );
  NAND2_X1 U8305 ( .A1(n8935), .A2(n9660), .ZN(n8031) );
  NAND2_X1 U8306 ( .A1(n9624), .A2(n9626), .ZN(n6631) );
  NAND2_X1 U8307 ( .A1(n6774), .A2(n9660), .ZN(n6630) );
  NAND2_X1 U8308 ( .A1(n6631), .A2(n6630), .ZN(n6770) );
  NAND2_X1 U8309 ( .A1(n6717), .A2(n9666), .ZN(n8017) );
  NAND2_X1 U8310 ( .A1(n9627), .A2(n6777), .ZN(n8032) );
  NAND2_X1 U8311 ( .A1(n8017), .A2(n8032), .ZN(n6772) );
  NAND2_X1 U8312 ( .A1(n6717), .A2(n6777), .ZN(n6632) );
  NAND2_X1 U8313 ( .A1(n6893), .A2(n6501), .ZN(n7875) );
  NAND2_X1 U8314 ( .A1(n8934), .A2(n9675), .ZN(n8020) );
  NAND2_X1 U8315 ( .A1(n8934), .A2(n6501), .ZN(n6634) );
  NAND2_X1 U8316 ( .A1(n6723), .A2(n6634), .ZN(n6885) );
  INV_X1 U8317 ( .A(n6885), .ZN(n6636) );
  INV_X1 U8318 ( .A(n8933), .ZN(n6716) );
  INV_X1 U8319 ( .A(n9678), .ZN(n6637) );
  NAND2_X1 U8320 ( .A1(n6637), .A2(n8933), .ZN(n7877) );
  NAND2_X1 U8321 ( .A1(n6637), .A2(n6716), .ZN(n6638) );
  INV_X1 U8322 ( .A(n8932), .ZN(n6894) );
  NAND2_X1 U8323 ( .A1(n6639), .A2(n6643), .ZN(n6642) );
  AOI22_X1 U8324 ( .A1(n7649), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7648), .B2(
        n6640), .ZN(n6641) );
  NAND2_X1 U8325 ( .A1(n6642), .A2(n6641), .ZN(n6803) );
  OR2_X1 U8326 ( .A1(n6894), .A2(n6803), .ZN(n8085) );
  NAND2_X1 U8327 ( .A1(n6803), .A2(n6894), .ZN(n7889) );
  NAND2_X1 U8328 ( .A1(n8085), .A2(n7889), .ZN(n6707) );
  AOI22_X1 U8329 ( .A1(n7649), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7648), .B2(
        n6645), .ZN(n6646) );
  INV_X1 U8330 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6648) );
  OAI22_X1 U8331 ( .A1(n4276), .A2(n6649), .B1(n7848), .B2(n6648), .ZN(n6654)
         );
  NAND2_X1 U8332 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND2_X1 U8333 ( .A1(n6664), .A2(n6652), .ZN(n7132) );
  OAI22_X1 U8334 ( .A1(n4272), .A2(n7132), .B1(n7636), .B2(n9943), .ZN(n6653)
         );
  INV_X1 U8335 ( .A(n8931), .ZN(n6655) );
  NAND2_X1 U8336 ( .A1(n7131), .A2(n6655), .ZN(n7891) );
  NOR2_X1 U8337 ( .A1(n6656), .A2(n6733), .ZN(n6657) );
  OR2_X1 U8338 ( .A1(n6729), .A2(n6657), .ZN(n9693) );
  NAND2_X1 U8339 ( .A1(n6658), .A2(n9193), .ZN(n6659) );
  NOR2_X1 U8340 ( .A1(n9648), .A2(n6659), .ZN(n9645) );
  INV_X1 U8341 ( .A(n9645), .ZN(n6679) );
  NAND2_X1 U8342 ( .A1(n8076), .A2(n9651), .ZN(n8074) );
  NAND2_X1 U8343 ( .A1(n6661), .A2(n8074), .ZN(n9625) );
  INV_X1 U8344 ( .A(n9626), .ZN(n7980) );
  NAND2_X1 U8345 ( .A1(n9625), .A2(n7980), .ZN(n6662) );
  NAND2_X1 U8346 ( .A1(n6771), .A2(n8032), .ZN(n6714) );
  AND2_X1 U8347 ( .A1(n8018), .A2(n8017), .ZN(n8083) );
  NAND2_X1 U8348 ( .A1(n7877), .A2(n8020), .ZN(n7982) );
  NAND2_X1 U8349 ( .A1(n7982), .A2(n7888), .ZN(n8084) );
  INV_X1 U8350 ( .A(n6733), .ZN(n7986) );
  XNOR2_X1 U8351 ( .A(n6734), .B(n7986), .ZN(n6671) );
  NAND2_X1 U8352 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  AND2_X1 U8353 ( .A1(n6736), .A2(n6665), .ZN(n7064) );
  NAND2_X1 U8354 ( .A1(n7797), .A2(n7064), .ZN(n6669) );
  NAND2_X1 U8355 ( .A1(n7633), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U8356 ( .A1(n7813), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8357 ( .A1(n7853), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6666) );
  NAND4_X1 U8358 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n8930)
         );
  OAI22_X1 U8359 ( .A1(n6894), .A2(n9287), .B1(n7121), .B2(n9289), .ZN(n6670)
         );
  AOI21_X1 U8360 ( .B1(n6671), .B2(n9451), .A(n6670), .ZN(n6672) );
  OAI21_X1 U8361 ( .B1(n9693), .B2(n9656), .A(n6672), .ZN(n9696) );
  NAND2_X1 U8362 ( .A1(n9696), .A2(n10029), .ZN(n6678) );
  OAI22_X1 U8363 ( .A1(n10029), .A2(n9943), .B1(n7132), .B2(n9635), .ZN(n6676)
         );
  INV_X1 U8364 ( .A(n7131), .ZN(n9695) );
  NAND2_X1 U8365 ( .A1(n6776), .A2(n9675), .ZN(n6886) );
  INV_X1 U8366 ( .A(n6744), .ZN(n6674) );
  OAI211_X1 U8367 ( .C1(n9695), .C2(n6702), .A(n6674), .B(n9640), .ZN(n9694)
         );
  NOR2_X1 U8368 ( .A1(n9694), .A2(n10037), .ZN(n6675) );
  AOI211_X1 U8369 ( .C1(n10033), .C2(n7131), .A(n6676), .B(n6675), .ZN(n6677)
         );
  OAI211_X1 U8370 ( .C1(n9693), .C2(n6679), .A(n6678), .B(n6677), .ZN(P1_U3283) );
  MUX2_X1 U8371 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7221), .S(n6818), .Z(n6680)
         );
  INV_X1 U8372 ( .A(n6680), .ZN(n6684) );
  MUX2_X1 U8373 ( .A(n6681), .B(P2_REG2_REG_10__SCAN_IN), .S(n6690), .Z(n8321)
         );
  OAI21_X1 U8374 ( .B1(n6686), .B2(n7151), .A(n6682), .ZN(n8322) );
  NAND2_X1 U8375 ( .A1(n8321), .A2(n8322), .ZN(n8320) );
  OAI21_X1 U8376 ( .B1(n6690), .B2(n6681), .A(n8320), .ZN(n6683) );
  NOR2_X1 U8377 ( .A1(n6683), .A2(n6684), .ZN(n6812) );
  AOI21_X1 U8378 ( .B1(n6684), .B2(n6683), .A(n6812), .ZN(n6699) );
  NOR2_X1 U8379 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5215), .ZN(n6696) );
  INV_X1 U8380 ( .A(n6690), .ZN(n8325) );
  OR2_X1 U8381 ( .A1(n6686), .A2(n6685), .ZN(n6689) );
  INV_X1 U8382 ( .A(n6687), .ZN(n6688) );
  INV_X1 U8383 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6691) );
  MUX2_X1 U8384 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6691), .S(n6690), .Z(n8328)
         );
  INV_X1 U8385 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6692) );
  MUX2_X1 U8386 ( .A(n6692), .B(P2_REG1_REG_11__SCAN_IN), .S(n6818), .Z(n6693)
         );
  NOR2_X1 U8387 ( .A1(n6694), .A2(n6693), .ZN(n6817) );
  AOI211_X1 U8388 ( .C1(n6694), .C2(n6693), .A(n6817), .B(n9418), .ZN(n6695)
         );
  AOI211_X1 U8389 ( .C1(n9417), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n6696), .B(
        n6695), .ZN(n6698) );
  NAND2_X1 U8390 ( .A1(n9424), .A2(n6818), .ZN(n6697) );
  OAI211_X1 U8391 ( .C1(n6699), .C2(n8370), .A(n6698), .B(n6697), .ZN(P2_U3256) );
  INV_X1 U8392 ( .A(n6707), .ZN(n7985) );
  OAI21_X1 U8393 ( .B1(n4352), .B2(n7985), .A(n6700), .ZN(n6701) );
  AOI222_X1 U8394 ( .A1(n9451), .A2(n6701), .B1(n8931), .B2(n9628), .C1(n8933), 
        .C2(n9630), .ZN(n9689) );
  INV_X1 U8395 ( .A(n6702), .ZN(n6703) );
  OAI211_X1 U8396 ( .C1(n4504), .C2(n4502), .A(n6703), .B(n9640), .ZN(n9688)
         );
  INV_X1 U8397 ( .A(n9688), .ZN(n6706) );
  INV_X1 U8398 ( .A(n9635), .ZN(n10031) );
  AOI22_X1 U8399 ( .A1(n9648), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6804), .B2(
        n10031), .ZN(n6704) );
  OAI21_X1 U8400 ( .B1(n9638), .B2(n4504), .A(n6704), .ZN(n6705) );
  AOI21_X1 U8401 ( .B1(n6706), .B2(n9644), .A(n6705), .ZN(n6712) );
  XNOR2_X1 U8402 ( .A(n6708), .B(n6707), .ZN(n9691) );
  NAND2_X1 U8403 ( .A1(n6709), .A2(n7799), .ZN(n6710) );
  NAND2_X1 U8404 ( .A1(n9691), .A2(n10041), .ZN(n6711) );
  OAI211_X1 U8405 ( .C1(n9689), .C2(n9648), .A(n6712), .B(n6711), .ZN(P1_U3284) );
  XOR2_X1 U8406 ( .A(n6713), .B(n7872), .Z(n6715) );
  OAI222_X1 U8407 ( .A1(n9287), .A2(n6717), .B1(n9289), .B2(n6716), .C1(n6715), 
        .C2(n9632), .ZN(n9677) );
  INV_X1 U8408 ( .A(n9677), .ZN(n6727) );
  OAI211_X1 U8409 ( .C1(n6776), .C2(n9675), .A(n9640), .B(n6886), .ZN(n9673)
         );
  INV_X1 U8410 ( .A(n9673), .ZN(n6722) );
  NOR2_X1 U8411 ( .A1(n9635), .A2(n6718), .ZN(n6719) );
  AOI21_X1 U8412 ( .B1(n9648), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6719), .ZN(
        n6720) );
  OAI21_X1 U8413 ( .B1(n9638), .B2(n9675), .A(n6720), .ZN(n6721) );
  AOI21_X1 U8414 ( .B1(n9644), .B2(n6722), .A(n6721), .ZN(n6726) );
  NAND2_X1 U8415 ( .A1(n6724), .A2(n6713), .ZN(n9672) );
  NAND3_X1 U8416 ( .A1(n6723), .A2(n9672), .A3(n10041), .ZN(n6725) );
  OAI211_X1 U8417 ( .C1(n6727), .C2(n9648), .A(n6726), .B(n6725), .ZN(P1_U3286) );
  NAND2_X1 U8418 ( .A1(n6730), .A2(n6643), .ZN(n6732) );
  AOI22_X1 U8419 ( .A1(n7649), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7648), .B2(
        n9572), .ZN(n6731) );
  XNOR2_X1 U8420 ( .A(n7063), .B(n7121), .ZN(n7988) );
  XNOR2_X1 U8421 ( .A(n6860), .B(n7988), .ZN(n9706) );
  INV_X1 U8422 ( .A(n9706), .ZN(n6749) );
  XNOR2_X1 U8423 ( .A(n6995), .B(n7988), .ZN(n6735) );
  NAND2_X1 U8424 ( .A1(n6735), .A2(n9451), .ZN(n6743) );
  NAND2_X1 U8425 ( .A1(n6736), .A2(n7117), .ZN(n6737) );
  AND2_X1 U8426 ( .A1(n6870), .A2(n6737), .ZN(n7118) );
  NAND2_X1 U8427 ( .A1(n7797), .A2(n7118), .ZN(n6741) );
  NAND2_X1 U8428 ( .A1(n7633), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8429 ( .A1(n7813), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U8430 ( .A1(n7853), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6738) );
  NAND4_X1 U8431 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n8929)
         );
  AOI22_X1 U8432 ( .A1(n9628), .A2(n8929), .B1(n9630), .B2(n8931), .ZN(n6742)
         );
  NAND2_X1 U8433 ( .A1(n6743), .A2(n6742), .ZN(n9704) );
  OAI211_X1 U8434 ( .C1(n6744), .C2(n9702), .A(n9640), .B(n6877), .ZN(n9700)
         );
  AOI22_X1 U8435 ( .A1(n9648), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7064), .B2(
        n10031), .ZN(n6746) );
  NAND2_X1 U8436 ( .A1(n10033), .A2(n7063), .ZN(n6745) );
  OAI211_X1 U8437 ( .C1(n9700), .C2(n10037), .A(n6746), .B(n6745), .ZN(n6747)
         );
  AOI21_X1 U8438 ( .B1(n9704), .B2(n10029), .A(n6747), .ZN(n6748) );
  OAI21_X1 U8439 ( .B1(n6749), .B2(n9292), .A(n6748), .ZN(P1_U3282) );
  XNOR2_X1 U8440 ( .A(n6750), .B(n6754), .ZN(n9818) );
  INV_X1 U8441 ( .A(n9818), .ZN(n6769) );
  NAND2_X1 U8442 ( .A1(n6835), .A2(n6751), .ZN(n6753) );
  NAND2_X1 U8443 ( .A1(n6753), .A2(n6752), .ZN(n6755) );
  XNOR2_X1 U8444 ( .A(n6755), .B(n6754), .ZN(n6756) );
  NAND2_X1 U8445 ( .A1(n6756), .A2(n9745), .ZN(n6759) );
  OAI22_X1 U8446 ( .A1(n7146), .A2(n8619), .B1(n6916), .B2(n8621), .ZN(n6757)
         );
  INV_X1 U8447 ( .A(n6757), .ZN(n6758) );
  NAND2_X1 U8448 ( .A1(n6759), .A2(n6758), .ZN(n9822) );
  AOI21_X1 U8449 ( .B1(n6831), .B2(n6765), .A(n9826), .ZN(n6760) );
  NAND2_X1 U8450 ( .A1(n6760), .A2(n7081), .ZN(n9819) );
  OR2_X1 U8451 ( .A1(n6761), .A2(n8375), .ZN(n8612) );
  OAI22_X1 U8452 ( .A1(n9757), .A2(n6763), .B1(n6762), .B2(n9755), .ZN(n6764)
         );
  AOI21_X1 U8453 ( .B1(n8609), .B2(n6765), .A(n6764), .ZN(n6766) );
  OAI21_X1 U8454 ( .B1(n9819), .B2(n8612), .A(n6766), .ZN(n6767) );
  AOI21_X1 U8455 ( .B1(n9822), .B2(n9757), .A(n6767), .ZN(n6768) );
  OAI21_X1 U8456 ( .B1(n8584), .B2(n6769), .A(n6768), .ZN(P2_U3289) );
  XOR2_X1 U8457 ( .A(n6770), .B(n6772), .Z(n9668) );
  XNOR2_X1 U8458 ( .A(n6772), .B(n6771), .ZN(n6773) );
  OAI222_X1 U8459 ( .A1(n9289), .A2(n6893), .B1(n9287), .B2(n6774), .C1(n6773), 
        .C2(n9632), .ZN(n9670) );
  NAND2_X1 U8460 ( .A1(n9670), .A2(n10029), .ZN(n6783) );
  INV_X1 U8461 ( .A(n6775), .ZN(n9641) );
  AOI211_X1 U8462 ( .C1(n9666), .C2(n9641), .A(n9458), .B(n6776), .ZN(n9665)
         );
  NOR2_X1 U8463 ( .A1(n9638), .A2(n6777), .ZN(n6781) );
  OAI22_X1 U8464 ( .A1(n10029), .A2(n6779), .B1(n6778), .B2(n9635), .ZN(n6780)
         );
  AOI211_X1 U8465 ( .C1(n9665), .C2(n9644), .A(n6781), .B(n6780), .ZN(n6782)
         );
  OAI211_X1 U8466 ( .C1(n9292), .C2(n9668), .A(n6783), .B(n6782), .ZN(P1_U3287) );
  INV_X1 U8467 ( .A(n6784), .ZN(n6788) );
  OAI22_X1 U8468 ( .A1(n6786), .A2(n9193), .B1(n9635), .B2(n6785), .ZN(n6787)
         );
  OAI21_X1 U8469 ( .B1(n6788), .B2(n6787), .A(n10029), .ZN(n6792) );
  OAI22_X1 U8470 ( .A1(n6789), .A2(n9638), .B1(n10029), .B2(n6106), .ZN(n6790)
         );
  INV_X1 U8471 ( .A(n6790), .ZN(n6791) );
  OAI211_X1 U8472 ( .C1(n9292), .C2(n6793), .A(n6792), .B(n6791), .ZN(P1_U3290) );
  NAND2_X1 U8473 ( .A1(n6803), .A2(n7808), .ZN(n6795) );
  NAND2_X1 U8474 ( .A1(n8932), .A2(n7824), .ZN(n6794) );
  NAND2_X1 U8475 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  XNOR2_X1 U8476 ( .A(n6796), .B(n7799), .ZN(n7044) );
  AOI22_X1 U8477 ( .A1(n6803), .A2(n7824), .B1(n7801), .B2(n8932), .ZN(n7045)
         );
  XNOR2_X1 U8478 ( .A(n7044), .B(n7045), .ZN(n6802) );
  INV_X1 U8479 ( .A(n4357), .ZN(n6798) );
  OAI21_X1 U8480 ( .B1(n6799), .B2(n6797), .A(n6798), .ZN(n6800) );
  INV_X1 U8481 ( .A(n6800), .ZN(n6801) );
  NAND2_X1 U8482 ( .A1(n6801), .A2(n6802), .ZN(n7048) );
  OAI21_X1 U8483 ( .B1(n6802), .B2(n6801), .A(n7048), .ZN(n6810) );
  AND2_X1 U8484 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8940) );
  AOI21_X1 U8485 ( .B1(n8918), .B2(n8931), .A(n8940), .ZN(n6808) );
  NAND2_X1 U8486 ( .A1(n8894), .A2(n6803), .ZN(n6807) );
  NAND2_X1 U8487 ( .A1(n8907), .A2(n6804), .ZN(n6806) );
  NAND2_X1 U8488 ( .A1(n8901), .A2(n8933), .ZN(n6805) );
  NAND4_X1 U8489 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6809)
         );
  AOI21_X1 U8490 ( .B1(n6810), .B2(n8898), .A(n6809), .ZN(n6811) );
  INV_X1 U8491 ( .A(n6811), .ZN(P1_U3211) );
  INV_X1 U8492 ( .A(n7669), .ZN(n6858) );
  OAI222_X1 U8493 ( .A1(n9402), .A2(n6858), .B1(P1_U3084), .B2(n8111), .C1(
        n7670), .C2(n9404), .ZN(P1_U3333) );
  NOR2_X1 U8494 ( .A1(n6818), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U8495 ( .A1(n6813), .A2(n6812), .ZN(n6816) );
  MUX2_X1 U8496 ( .A(n7212), .B(P2_REG2_REG_12__SCAN_IN), .S(n6944), .Z(n6814)
         );
  INV_X1 U8497 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8498 ( .A1(n6815), .A2(n6816), .ZN(n6939) );
  OAI211_X1 U8499 ( .C1(n6816), .C2(n6815), .A(n9722), .B(n6939), .ZN(n6827)
         );
  AOI21_X1 U8500 ( .B1(n6818), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6817), .ZN(
        n6821) );
  MUX2_X1 U8501 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6819), .S(n6944), .Z(n6820)
         );
  NAND2_X1 U8502 ( .A1(n6821), .A2(n6820), .ZN(n6943) );
  OAI21_X1 U8503 ( .B1(n6821), .B2(n6820), .A(n6943), .ZN(n6825) );
  NOR2_X1 U8504 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7172), .ZN(n6824) );
  INV_X1 U8505 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6822) );
  NOR2_X1 U8506 ( .A1(n9731), .A2(n6822), .ZN(n6823) );
  AOI211_X1 U8507 ( .C1(n9724), .C2(n6825), .A(n6824), .B(n6823), .ZN(n6826)
         );
  OAI211_X1 U8508 ( .C1(n9726), .C2(n6828), .A(n6827), .B(n6826), .ZN(P2_U3257) );
  XNOR2_X1 U8509 ( .A(n6829), .B(n6830), .ZN(n6898) );
  INV_X1 U8510 ( .A(n6920), .ZN(n6833) );
  INV_X1 U8511 ( .A(n6831), .ZN(n6832) );
  AOI211_X1 U8512 ( .C1(n6839), .C2(n6833), .A(n9826), .B(n6832), .ZN(n6905)
         );
  XNOR2_X1 U8513 ( .A(n6835), .B(n6834), .ZN(n6836) );
  OAI222_X1 U8514 ( .A1(n8619), .A2(n7074), .B1(n8621), .B2(n6837), .C1(n6836), 
        .C2(n8566), .ZN(n6899) );
  AOI211_X1 U8515 ( .C1(n6898), .C2(n9838), .A(n6905), .B(n6899), .ZN(n6842)
         );
  AOI22_X1 U8516 ( .A1(n5551), .A2(n6839), .B1(n9853), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8517 ( .B1(n6842), .B2(n9853), .A(n6838), .ZN(P2_U3526) );
  INV_X1 U8518 ( .A(n8770), .ZN(n6840) );
  AOI22_X1 U8519 ( .A1(n6840), .A2(n6839), .B1(n5900), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n6841) );
  OAI21_X1 U8520 ( .B1(n6842), .B2(n5900), .A(n6841), .ZN(P2_U3469) );
  XOR2_X1 U8521 ( .A(n6843), .B(n6844), .Z(n9788) );
  XNOR2_X1 U8522 ( .A(n6845), .B(n6844), .ZN(n6849) );
  NAND2_X1 U8523 ( .A1(n8290), .A2(n9742), .ZN(n6846) );
  OAI21_X1 U8524 ( .B1(n6847), .B2(n8619), .A(n6846), .ZN(n6848) );
  AOI21_X1 U8525 ( .B1(n6849), .B2(n9745), .A(n6848), .ZN(n9791) );
  INV_X2 U8526 ( .A(n9757), .ZN(n9766) );
  MUX2_X1 U8527 ( .A(n9791), .B(n9931), .S(n9766), .Z(n6856) );
  OR2_X1 U8528 ( .A1(n9781), .A2(n9789), .ZN(n6850) );
  NAND2_X1 U8529 ( .A1(n6851), .A2(n6850), .ZN(n9790) );
  OAI22_X1 U8530 ( .A1(n7154), .A2(n9790), .B1(n6852), .B2(n9755), .ZN(n6853)
         );
  AOI21_X1 U8531 ( .B1(n8609), .B2(n6854), .A(n6853), .ZN(n6855) );
  OAI211_X1 U8532 ( .C1(n9788), .C2(n8584), .A(n6856), .B(n6855), .ZN(P2_U3294) );
  OAI222_X1 U8533 ( .A1(n7376), .A2(n6859), .B1(n8783), .B2(n6858), .C1(n6857), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8534 ( .A1(n6862), .A2(n6643), .ZN(n6865) );
  AOI22_X1 U8535 ( .A1(n7649), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7648), .B2(
        n6863), .ZN(n6864) );
  INV_X1 U8536 ( .A(n8929), .ZN(n6866) );
  OR2_X1 U8537 ( .A1(n7123), .A2(n6866), .ZN(n7895) );
  NAND2_X1 U8538 ( .A1(n7123), .A2(n6866), .ZN(n7883) );
  NAND2_X1 U8539 ( .A1(n7895), .A2(n7883), .ZN(n7989) );
  OAI21_X1 U8540 ( .B1(n4355), .B2(n7989), .A(n7010), .ZN(n6867) );
  INV_X1 U8541 ( .A(n6867), .ZN(n6967) );
  INV_X1 U8542 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6868) );
  OAI22_X1 U8543 ( .A1(n4277), .A2(n9482), .B1(n7848), .B2(n6868), .ZN(n6873)
         );
  INV_X1 U8544 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8545 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  NAND2_X1 U8546 ( .A1(n7001), .A2(n6871), .ZN(n7284) );
  INV_X1 U8547 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7011) );
  OAI22_X1 U8548 ( .A1(n4272), .A2(n7284), .B1(n7636), .B2(n7011), .ZN(n6872)
         );
  OR2_X1 U8549 ( .A1(n7063), .A2(n7121), .ZN(n7878) );
  INV_X1 U8550 ( .A(n7878), .ZN(n6874) );
  NAND2_X1 U8551 ( .A1(n7063), .A2(n7121), .ZN(n7892) );
  OAI21_X1 U8552 ( .B1(n6995), .B2(n6874), .A(n7892), .ZN(n6875) );
  XNOR2_X1 U8553 ( .A(n6875), .B(n7989), .ZN(n6876) );
  OAI222_X1 U8554 ( .A1(n9289), .A2(n7369), .B1(n9287), .B2(n7121), .C1(n6876), 
        .C2(n9632), .ZN(n6964) );
  INV_X1 U8555 ( .A(n7123), .ZN(n6880) );
  INV_X1 U8556 ( .A(n7012), .ZN(n7013) );
  AOI211_X1 U8557 ( .C1(n7123), .C2(n6877), .A(n9458), .B(n7013), .ZN(n6965)
         );
  NAND2_X1 U8558 ( .A1(n6965), .A2(n9644), .ZN(n6879) );
  AOI22_X1 U8559 ( .A1(n9648), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7118), .B2(
        n10031), .ZN(n6878) );
  OAI211_X1 U8560 ( .C1(n6880), .C2(n9638), .A(n6879), .B(n6878), .ZN(n6881)
         );
  AOI21_X1 U8561 ( .B1(n6964), .B2(n10029), .A(n6881), .ZN(n6882) );
  OAI21_X1 U8562 ( .B1(n6967), .B2(n9292), .A(n6882), .ZN(P1_U3281) );
  INV_X1 U8563 ( .A(n6883), .ZN(n6884) );
  AOI21_X1 U8564 ( .B1(n7874), .B2(n6885), .A(n6884), .ZN(n9683) );
  INV_X1 U8565 ( .A(n9683), .ZN(n9686) );
  AOI21_X1 U8566 ( .B1(n6886), .B2(n9678), .A(n9458), .ZN(n6888) );
  NAND2_X1 U8567 ( .A1(n6888), .A2(n6887), .ZN(n9681) );
  AOI22_X1 U8568 ( .A1(n10033), .A2(n9678), .B1(n10031), .B2(n6889), .ZN(n6890) );
  OAI21_X1 U8569 ( .B1(n10037), .B2(n9681), .A(n6890), .ZN(n6896) );
  INV_X1 U8570 ( .A(n7875), .ZN(n7871) );
  AOI21_X1 U8571 ( .B1(n7872), .B2(n6713), .A(n7871), .ZN(n6891) );
  XNOR2_X1 U8572 ( .A(n6891), .B(n7874), .ZN(n6892) );
  OAI222_X1 U8573 ( .A1(n9289), .A2(n6894), .B1(n9287), .B2(n6893), .C1(n6892), 
        .C2(n9632), .ZN(n9685) );
  MUX2_X1 U8574 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9685), .S(n10029), .Z(n6895)
         );
  AOI211_X1 U8575 ( .C1(n10041), .C2(n9686), .A(n6896), .B(n6895), .ZN(n6897)
         );
  INV_X1 U8576 ( .A(n6897), .ZN(P1_U3285) );
  INV_X1 U8577 ( .A(n6898), .ZN(n6908) );
  INV_X1 U8578 ( .A(n6899), .ZN(n6900) );
  MUX2_X1 U8579 ( .A(n6901), .B(n6900), .S(n9757), .Z(n6907) );
  OAI22_X1 U8580 ( .A1(n9762), .A2(n6903), .B1(n9755), .B2(n6902), .ZN(n6904)
         );
  AOI21_X1 U8581 ( .B1(n6905), .B2(n8634), .A(n6904), .ZN(n6906) );
  OAI211_X1 U8582 ( .C1(n8584), .C2(n6908), .A(n6907), .B(n6906), .ZN(P2_U3290) );
  XOR2_X1 U8583 ( .A(n6914), .B(n6909), .Z(n9816) );
  NAND2_X1 U8584 ( .A1(n6602), .A2(n6910), .ZN(n9738) );
  NAND2_X1 U8585 ( .A1(n9738), .A2(n6911), .ZN(n6913) );
  NAND2_X1 U8586 ( .A1(n6913), .A2(n6912), .ZN(n6915) );
  XNOR2_X1 U8587 ( .A(n6915), .B(n6914), .ZN(n6918) );
  OAI22_X1 U8588 ( .A1(n6917), .A2(n8621), .B1(n6916), .B2(n8619), .ZN(n8128)
         );
  AOI21_X1 U8589 ( .B1(n6918), .B2(n9745), .A(n8128), .ZN(n9814) );
  MUX2_X1 U8590 ( .A(n9814), .B(n6429), .S(n9766), .Z(n6923) );
  INV_X1 U8591 ( .A(n6919), .ZN(n9753) );
  AOI211_X1 U8592 ( .C1(n9811), .C2(n9753), .A(n9826), .B(n6920), .ZN(n9810)
         );
  OAI22_X1 U8593 ( .A1(n9762), .A2(n8131), .B1(n8130), .B2(n9755), .ZN(n6921)
         );
  AOI21_X1 U8594 ( .B1(n9810), .B2(n8634), .A(n6921), .ZN(n6922) );
  OAI211_X1 U8595 ( .C1(n9816), .C2(n8584), .A(n6923), .B(n6922), .ZN(P2_U3291) );
  INV_X1 U8596 ( .A(n7689), .ZN(n6937) );
  OAI222_X1 U8597 ( .A1(n9402), .A2(n6937), .B1(P1_U3084), .B2(n8062), .C1(
        n7690), .C2(n9404), .ZN(P1_U3332) );
  INV_X1 U8598 ( .A(n6927), .ZN(n6924) );
  AOI21_X1 U8599 ( .B1(n6925), .B2(n6924), .A(n8244), .ZN(n6930) );
  NOR3_X1 U8600 ( .A1(n8242), .A2(n6926), .A3(n7074), .ZN(n6929) );
  NAND2_X1 U8601 ( .A1(n6928), .A2(n6927), .ZN(n6956) );
  OAI21_X1 U8602 ( .B1(n6930), .B2(n6929), .A(n6956), .ZN(n6935) );
  INV_X1 U8603 ( .A(n6931), .ZN(n7082) );
  OAI22_X1 U8604 ( .A1(n7332), .A2(n8234), .B1(n8233), .B2(n7074), .ZN(n6932)
         );
  AOI211_X1 U8605 ( .C1(n7082), .C2(n8266), .A(n6933), .B(n6932), .ZN(n6934)
         );
  OAI211_X1 U8606 ( .C1(n7084), .C2(n8270), .A(n6935), .B(n6934), .ZN(P2_U3223) );
  OAI222_X1 U8607 ( .A1(n7376), .A2(n6938), .B1(n8783), .B2(n6937), .C1(n6936), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8608 ( .A1(n6944), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8609 ( .A1(n6940), .A2(n6939), .ZN(n6942) );
  AOI22_X1 U8610 ( .A1(n7094), .A2(n7323), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7089), .ZN(n6941) );
  NOR2_X1 U8611 ( .A1(n6942), .A2(n6941), .ZN(n7088) );
  AOI21_X1 U8612 ( .B1(n6942), .B2(n6941), .A(n7088), .ZN(n6952) );
  AOI22_X1 U8613 ( .A1(n7094), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5253), .B2(
        n7089), .ZN(n6946) );
  OAI21_X1 U8614 ( .B1(n6944), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6943), .ZN(
        n6945) );
  OAI21_X1 U8615 ( .B1(n6946), .B2(n6945), .A(n7093), .ZN(n6950) );
  NOR2_X1 U8616 ( .A1(n6947), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7305) );
  AOI21_X1 U8617 ( .B1(n9417), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7305), .ZN(
        n6948) );
  OAI21_X1 U8618 ( .B1(n9726), .B2(n7089), .A(n6948), .ZN(n6949) );
  AOI21_X1 U8619 ( .B1(n6950), .B2(n9724), .A(n6949), .ZN(n6951) );
  OAI21_X1 U8620 ( .B1(n6952), .B2(n8370), .A(n6951), .ZN(P2_U3258) );
  NAND2_X1 U8621 ( .A1(n6954), .A2(n6953), .ZN(n6958) );
  NAND2_X1 U8622 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  XOR2_X1 U8623 ( .A(n6958), .B(n6957), .Z(n6963) );
  AOI22_X1 U8624 ( .A1(n8199), .A2(n8286), .B1(n8198), .B2(n8284), .ZN(n6960)
         );
  OAI211_X1 U8625 ( .C1(n7150), .C2(n8251), .A(n6960), .B(n6959), .ZN(n6961)
         );
  AOI21_X1 U8626 ( .B1(n7157), .B2(n8238), .A(n6961), .ZN(n6962) );
  OAI21_X1 U8627 ( .B1(n6963), .B2(n8244), .A(n6962), .ZN(P2_U3233) );
  INV_X1 U8628 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6969) );
  AOI211_X1 U8629 ( .C1(n9679), .C2(n7123), .A(n6965), .B(n6964), .ZN(n6966)
         );
  OAI21_X1 U8630 ( .B1(n6967), .B2(n9373), .A(n6966), .ZN(n6983) );
  NAND2_X1 U8631 ( .A1(n6983), .A2(n9709), .ZN(n6968) );
  OAI21_X1 U8632 ( .B1(n9709), .B2(n6969), .A(n6968), .ZN(P1_U3484) );
  XNOR2_X1 U8633 ( .A(n6971), .B(n6970), .ZN(n9787) );
  INV_X1 U8634 ( .A(n6972), .ZN(n6973) );
  NAND2_X1 U8635 ( .A1(n6973), .A2(n6970), .ZN(n6974) );
  NAND3_X1 U8636 ( .A1(n6975), .A2(n9745), .A3(n6974), .ZN(n6977) );
  AOI22_X1 U8637 ( .A1(n9742), .A2(n5481), .B1(n8289), .B2(n9740), .ZN(n6976)
         );
  NAND2_X1 U8638 ( .A1(n6977), .A2(n6976), .ZN(n9785) );
  MUX2_X1 U8639 ( .A(n9785), .B(P2_REG2_REG_1__SCAN_IN), .S(n9766), .Z(n6981)
         );
  NOR2_X1 U8640 ( .A1(n9784), .A2(n9776), .ZN(n9782) );
  NOR3_X1 U8641 ( .A1(n7154), .A2(n9781), .A3(n9782), .ZN(n6978) );
  AOI21_X1 U8642 ( .B1(n8570), .B2(P2_REG3_REG_1__SCAN_IN), .A(n6978), .ZN(
        n6979) );
  OAI21_X1 U8643 ( .B1(n9784), .B2(n9762), .A(n6979), .ZN(n6980) );
  AOI211_X1 U8644 ( .C1(n9764), .C2(n9787), .A(n6981), .B(n6980), .ZN(n6982)
         );
  INV_X1 U8645 ( .A(n6982), .ZN(P2_U3295) );
  NAND2_X1 U8646 ( .A1(n6983), .A2(n9721), .ZN(n6984) );
  OAI21_X1 U8647 ( .B1(n9721), .B2(n6985), .A(n6984), .ZN(P1_U3533) );
  INV_X1 U8648 ( .A(n7711), .ZN(n6987) );
  OAI222_X1 U8649 ( .A1(n8121), .A2(n7712), .B1(n9402), .B2(n6987), .C1(n6132), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U8650 ( .A1(n7376), .A2(n6988), .B1(n8783), .B2(n6987), .C1(
        P2_U3152), .C2(n6986), .ZN(P2_U3336) );
  XNOR2_X1 U8651 ( .A(n6990), .B(n6989), .ZN(n6994) );
  AOI22_X1 U8652 ( .A1(n8199), .A2(n8285), .B1(n8198), .B2(n8283), .ZN(n6991)
         );
  NAND2_X1 U8653 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8323) );
  OAI211_X1 U8654 ( .C1(n7341), .C2(n8251), .A(n6991), .B(n8323), .ZN(n6992)
         );
  AOI21_X1 U8655 ( .B1(n7455), .B2(n8238), .A(n6992), .ZN(n6993) );
  OAI21_X1 U8656 ( .B1(n6994), .B2(n8244), .A(n6993), .ZN(P2_U3219) );
  NAND2_X1 U8657 ( .A1(n7895), .A2(n7878), .ZN(n8037) );
  NAND2_X1 U8658 ( .A1(n7883), .A2(n7892), .ZN(n7879) );
  AND2_X1 U8659 ( .A1(n7879), .A2(n7895), .ZN(n8026) );
  NOR2_X1 U8660 ( .A1(n9042), .A2(n8026), .ZN(n7194) );
  NAND2_X1 U8661 ( .A1(n6996), .A2(n6643), .ZN(n6998) );
  AOI22_X1 U8662 ( .A1(n7649), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7648), .B2(
        n9592), .ZN(n6997) );
  NOR2_X1 U8663 ( .A1(n7286), .A2(n7369), .ZN(n7901) );
  NAND2_X1 U8664 ( .A1(n7286), .A2(n7369), .ZN(n7898) );
  INV_X1 U8665 ( .A(n7898), .ZN(n6999) );
  OR2_X1 U8666 ( .A1(n7901), .A2(n6999), .ZN(n7976) );
  XNOR2_X1 U8667 ( .A(n7194), .B(n7976), .ZN(n7008) );
  INV_X1 U8668 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8669 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U8670 ( .A1(n7190), .A2(n7002), .ZN(n7199) );
  INV_X1 U8671 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7003) );
  OAI22_X1 U8672 ( .A1(n4272), .A2(n7199), .B1(n7848), .B2(n7003), .ZN(n7007)
         );
  INV_X1 U8673 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7004) );
  OAI22_X1 U8674 ( .A1(n4276), .A2(n7005), .B1(n7636), .B2(n7004), .ZN(n7006)
         );
  AOI222_X1 U8675 ( .A1(n9451), .A2(n7008), .B1(n9435), .B2(n9628), .C1(n8929), 
        .C2(n9630), .ZN(n9478) );
  XNOR2_X1 U8676 ( .A(n7184), .B(n7976), .ZN(n9481) );
  NAND2_X1 U8677 ( .A1(n9481), .A2(n10041), .ZN(n7017) );
  OAI22_X1 U8678 ( .A1(n10029), .A2(n7011), .B1(n7284), .B2(n9635), .ZN(n7015)
         );
  INV_X1 U8679 ( .A(n7286), .ZN(n9479) );
  INV_X1 U8680 ( .A(n7197), .ZN(n7198) );
  OAI211_X1 U8681 ( .C1(n9479), .C2(n7013), .A(n7198), .B(n9640), .ZN(n9477)
         );
  NOR2_X1 U8682 ( .A1(n9477), .A2(n10037), .ZN(n7014) );
  AOI211_X1 U8683 ( .C1(n10033), .C2(n7286), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI211_X1 U8684 ( .C1(n9648), .C2(n9478), .A(n7017), .B(n7016), .ZN(P1_U3280) );
  XNOR2_X1 U8685 ( .A(n8078), .B(n7978), .ZN(n7018) );
  AOI222_X1 U8686 ( .A1(n9451), .A2(n7018), .B1(n6241), .B2(n9630), .C1(n8935), 
        .C2(n9628), .ZN(n9653) );
  AOI21_X1 U8687 ( .B1(n9651), .B2(n7019), .A(n9458), .ZN(n7020) );
  NAND2_X1 U8688 ( .A1(n4469), .A2(n7020), .ZN(n9652) );
  NAND2_X1 U8689 ( .A1(n9648), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8690 ( .A1(n10031), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7021) );
  OAI211_X1 U8691 ( .C1(n9652), .C2(n10037), .A(n7022), .B(n7021), .ZN(n7025)
         );
  XOR2_X1 U8692 ( .A(n7023), .B(n7978), .Z(n9655) );
  NOR2_X1 U8693 ( .A1(n9292), .A2(n9655), .ZN(n7024) );
  AOI211_X1 U8694 ( .C1(n10033), .C2(n9651), .A(n7025), .B(n7024), .ZN(n7026)
         );
  OAI21_X1 U8695 ( .B1(n9648), .B2(n9653), .A(n7026), .ZN(P1_U3289) );
  INV_X1 U8696 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7028) );
  NOR2_X1 U8697 ( .A1(n7028), .A2(n7029), .ZN(n7291) );
  AOI211_X1 U8698 ( .C1(n7029), .C2(n7028), .A(n7291), .B(n9578), .ZN(n7030)
         );
  AOI21_X1 U8699 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9619), .A(n7030), .ZN(
        n7038) );
  INV_X1 U8700 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7031) );
  MUX2_X1 U8701 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7031), .S(n7558), .Z(n7034)
         );
  NAND2_X1 U8702 ( .A1(n7034), .A2(n7033), .ZN(n7294) );
  OAI21_X1 U8703 ( .B1(n7034), .B2(n7033), .A(n7294), .ZN(n7036) );
  NAND2_X1 U8704 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8799) );
  INV_X1 U8705 ( .A(n8799), .ZN(n7035) );
  AOI21_X1 U8706 ( .B1(n9620), .B2(n7036), .A(n7035), .ZN(n7037) );
  OAI211_X1 U8707 ( .C1(n7289), .C2(n9613), .A(n7038), .B(n7037), .ZN(P1_U3255) );
  INV_X1 U8708 ( .A(n7730), .ZN(n7041) );
  NAND2_X1 U8709 ( .A1(n8780), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7039) );
  OAI211_X1 U8710 ( .C1(n7041), .C2(n8783), .A(n7040), .B(n7039), .ZN(P2_U3335) );
  NAND2_X1 U8711 ( .A1(n7730), .A2(n9398), .ZN(n7043) );
  OR2_X1 U8712 ( .A1(n7042), .A2(P1_U3084), .ZN(n8117) );
  OAI211_X1 U8713 ( .C1(n7731), .C2(n9404), .A(n7043), .B(n8117), .ZN(P1_U3330) );
  INV_X1 U8714 ( .A(n7044), .ZN(n7046) );
  NAND2_X1 U8715 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  NAND2_X1 U8716 ( .A1(n7131), .A2(n7824), .ZN(n7050) );
  NAND2_X1 U8717 ( .A1(n7801), .A2(n8931), .ZN(n7049) );
  NAND2_X1 U8718 ( .A1(n7050), .A2(n7049), .ZN(n7055) );
  NAND2_X1 U8719 ( .A1(n7054), .A2(n7055), .ZN(n7126) );
  NAND2_X1 U8720 ( .A1(n7131), .A2(n7808), .ZN(n7052) );
  NAND2_X1 U8721 ( .A1(n8931), .A2(n7824), .ZN(n7051) );
  NAND2_X1 U8722 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  XNOR2_X1 U8723 ( .A(n7053), .B(n7822), .ZN(n7129) );
  NAND2_X1 U8724 ( .A1(n7126), .A2(n7129), .ZN(n7058) );
  INV_X1 U8725 ( .A(n7055), .ZN(n7056) );
  NAND2_X1 U8726 ( .A1(n7057), .A2(n7056), .ZN(n7127) );
  NAND2_X1 U8727 ( .A1(n7063), .A2(n7808), .ZN(n7060) );
  NAND2_X1 U8728 ( .A1(n8930), .A2(n7824), .ZN(n7059) );
  NAND2_X1 U8729 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  XNOR2_X1 U8730 ( .A(n7061), .B(n7799), .ZN(n7108) );
  AND2_X1 U8731 ( .A1(n8930), .A2(n7801), .ZN(n7062) );
  AOI21_X1 U8732 ( .B1(n7063), .B2(n7824), .A(n7062), .ZN(n7109) );
  XNOR2_X1 U8733 ( .A(n7108), .B(n7109), .ZN(n7106) );
  XNOR2_X1 U8734 ( .A(n7107), .B(n7106), .ZN(n7070) );
  AND2_X1 U8735 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9570) );
  AOI21_X1 U8736 ( .B1(n8918), .B2(n8929), .A(n9570), .ZN(n7068) );
  NAND2_X1 U8737 ( .A1(n7063), .A2(n8894), .ZN(n7067) );
  NAND2_X1 U8738 ( .A1(n8907), .A2(n7064), .ZN(n7066) );
  NAND2_X1 U8739 ( .A1(n8901), .A2(n8931), .ZN(n7065) );
  NAND4_X1 U8740 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(n7069)
         );
  AOI21_X1 U8741 ( .B1(n7070), .B2(n8898), .A(n7069), .ZN(n7071) );
  INV_X1 U8742 ( .A(n7071), .ZN(P1_U3229) );
  XNOR2_X1 U8743 ( .A(n7073), .B(n7072), .ZN(n7080) );
  OAI22_X1 U8744 ( .A1(n7332), .A2(n8619), .B1(n7074), .B2(n8621), .ZN(n7079)
         );
  OAI21_X1 U8745 ( .B1(n7077), .B2(n7076), .A(n7075), .ZN(n7237) );
  NOR2_X1 U8746 ( .A1(n7237), .A2(n8626), .ZN(n7078) );
  AOI211_X1 U8747 ( .C1(n7080), .C2(n9745), .A(n7079), .B(n7078), .ZN(n7236)
         );
  AOI21_X1 U8748 ( .B1(n7233), .B2(n7081), .A(n7152), .ZN(n7234) );
  AOI22_X1 U8749 ( .A1(n9766), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7082), .B2(
        n8570), .ZN(n7083) );
  OAI21_X1 U8750 ( .B1(n9762), .B2(n7084), .A(n7083), .ZN(n7086) );
  NOR2_X1 U8751 ( .A1(n7237), .A2(n8637), .ZN(n7085) );
  AOI211_X1 U8752 ( .C1(n7234), .C2(n9759), .A(n7086), .B(n7085), .ZN(n7087)
         );
  OAI21_X1 U8753 ( .B1(n7236), .B2(n9766), .A(n7087), .ZN(P2_U3288) );
  AOI21_X1 U8754 ( .B1(n7089), .B2(n7323), .A(n7088), .ZN(n7092) );
  AND2_X1 U8755 ( .A1(n7419), .A2(n7495), .ZN(n7417) );
  INV_X1 U8756 ( .A(n7417), .ZN(n7090) );
  OAI21_X1 U8757 ( .B1(n7495), .B2(n7419), .A(n7090), .ZN(n7091) );
  NOR2_X1 U8758 ( .A1(n7092), .A2(n7091), .ZN(n7416) );
  AOI21_X1 U8759 ( .B1(n7092), .B2(n7091), .A(n7416), .ZN(n7105) );
  NAND2_X1 U8760 ( .A1(n7419), .A2(n7096), .ZN(n7095) );
  OAI21_X1 U8761 ( .B1(n7419), .B2(n7096), .A(n7095), .ZN(n7097) );
  INV_X1 U8762 ( .A(n7097), .ZN(n7098) );
  NAND2_X1 U8763 ( .A1(n7099), .A2(n7098), .ZN(n7420) );
  OAI21_X1 U8764 ( .B1(n7099), .B2(n7098), .A(n7420), .ZN(n7103) );
  NOR2_X1 U8765 ( .A1(n7100), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7432) );
  AOI21_X1 U8766 ( .B1(n9417), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7432), .ZN(
        n7101) );
  OAI21_X1 U8767 ( .B1(n9726), .B2(n7419), .A(n7101), .ZN(n7102) );
  AOI21_X1 U8768 ( .B1(n7103), .B2(n9724), .A(n7102), .ZN(n7104) );
  OAI21_X1 U8769 ( .B1(n7105), .B2(n8370), .A(n7104), .ZN(P2_U3259) );
  INV_X1 U8770 ( .A(n7108), .ZN(n7110) );
  NAND2_X1 U8771 ( .A1(n7110), .A2(n7109), .ZN(n7111) );
  NAND2_X1 U8772 ( .A1(n7123), .A2(n7808), .ZN(n7113) );
  NAND2_X1 U8773 ( .A1(n8929), .A2(n7824), .ZN(n7112) );
  NAND2_X1 U8774 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  XNOR2_X1 U8775 ( .A(n7114), .B(n7822), .ZN(n7271) );
  AND2_X1 U8776 ( .A1(n8929), .A2(n7801), .ZN(n7115) );
  AOI21_X1 U8777 ( .B1(n7123), .B2(n7824), .A(n7115), .ZN(n7272) );
  XNOR2_X1 U8778 ( .A(n7271), .B(n7272), .ZN(n7116) );
  XNOR2_X1 U8779 ( .A(n7276), .B(n7116), .ZN(n7125) );
  NOR2_X1 U8780 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7117), .ZN(n9583) );
  AOI21_X1 U8781 ( .B1(n8918), .B2(n8928), .A(n9583), .ZN(n7120) );
  NAND2_X1 U8782 ( .A1(n8907), .A2(n7118), .ZN(n7119) );
  OAI211_X1 U8783 ( .C1(n7121), .C2(n8916), .A(n7120), .B(n7119), .ZN(n7122)
         );
  AOI21_X1 U8784 ( .B1(n7123), .B2(n8894), .A(n7122), .ZN(n7124) );
  OAI21_X1 U8785 ( .B1(n7125), .B2(n8923), .A(n7124), .ZN(P1_U3215) );
  NAND2_X1 U8786 ( .A1(n7126), .A2(n7127), .ZN(n7128) );
  XOR2_X1 U8787 ( .A(n7129), .B(n7128), .Z(n7139) );
  AOI21_X1 U8788 ( .B1(n8918), .B2(n8930), .A(n7130), .ZN(n7137) );
  NAND2_X1 U8789 ( .A1(n7131), .A2(n8894), .ZN(n7136) );
  INV_X1 U8790 ( .A(n7132), .ZN(n7133) );
  NAND2_X1 U8791 ( .A1(n8907), .A2(n7133), .ZN(n7135) );
  NAND2_X1 U8792 ( .A1(n8901), .A2(n8932), .ZN(n7134) );
  NAND4_X1 U8793 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n7134), .ZN(n7138)
         );
  AOI21_X1 U8794 ( .B1(n7139), .B2(n8898), .A(n7138), .ZN(n7140) );
  INV_X1 U8795 ( .A(n7140), .ZN(P1_U3219) );
  INV_X1 U8796 ( .A(n7141), .ZN(n7142) );
  AOI21_X1 U8797 ( .B1(n7144), .B2(n7143), .A(n7142), .ZN(n9824) );
  XNOR2_X1 U8798 ( .A(n7145), .B(n7144), .ZN(n7148) );
  OAI22_X1 U8799 ( .A1(n7146), .A2(n8621), .B1(n7162), .B2(n8619), .ZN(n7147)
         );
  AOI21_X1 U8800 ( .B1(n7148), .B2(n9745), .A(n7147), .ZN(n7149) );
  OAI21_X1 U8801 ( .B1(n9824), .B2(n8626), .A(n7149), .ZN(n9828) );
  NAND2_X1 U8802 ( .A1(n9828), .A2(n9757), .ZN(n7159) );
  OAI22_X1 U8803 ( .A1(n9757), .A2(n7151), .B1(n7150), .B2(n9755), .ZN(n7156)
         );
  NOR2_X1 U8804 ( .A1(n7152), .A2(n9825), .ZN(n7153) );
  OR2_X1 U8805 ( .A1(n7338), .A2(n7153), .ZN(n9827) );
  NOR2_X1 U8806 ( .A1(n9827), .A2(n7154), .ZN(n7155) );
  AOI211_X1 U8807 ( .C1(n8609), .C2(n7157), .A(n7156), .B(n7155), .ZN(n7158)
         );
  OAI211_X1 U8808 ( .C1(n9824), .C2(n8637), .A(n7159), .B(n7158), .ZN(P2_U3287) );
  XNOR2_X1 U8809 ( .A(n7160), .B(n7161), .ZN(n7166) );
  OAI22_X1 U8810 ( .A1(n8251), .A2(n7220), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5215), .ZN(n7164) );
  OAI22_X1 U8811 ( .A1(n7162), .A2(n8233), .B1(n8234), .B2(n7304), .ZN(n7163)
         );
  AOI211_X1 U8812 ( .C1(n7226), .C2(n8238), .A(n7164), .B(n7163), .ZN(n7165)
         );
  OAI21_X1 U8813 ( .B1(n7166), .B2(n8244), .A(n7165), .ZN(P2_U3238) );
  INV_X1 U8814 ( .A(n7543), .ZN(n7178) );
  OAI222_X1 U8815 ( .A1(n9402), .A2(n7178), .B1(P1_U3084), .B2(n7167), .C1(
        n10002), .C2(n9404), .ZN(P1_U3329) );
  XNOR2_X1 U8816 ( .A(n7168), .B(n7169), .ZN(n7176) );
  NAND2_X1 U8817 ( .A1(n8281), .A2(n9740), .ZN(n7171) );
  NAND2_X1 U8818 ( .A1(n8283), .A2(n9742), .ZN(n7170) );
  AND2_X1 U8819 ( .A1(n7171), .A2(n7170), .ZN(n7206) );
  OAI22_X1 U8820 ( .A1(n8264), .A2(n7206), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7172), .ZN(n7174) );
  NOR2_X1 U8821 ( .A1(n8251), .A2(n7211), .ZN(n7173) );
  AOI211_X1 U8822 ( .C1(n7210), .C2(n8238), .A(n7174), .B(n7173), .ZN(n7175)
         );
  OAI21_X1 U8823 ( .B1(n7176), .B2(n8244), .A(n7175), .ZN(P2_U3226) );
  OAI222_X1 U8824 ( .A1(P2_U3152), .A2(n7179), .B1(n8783), .B2(n7178), .C1(
        n7177), .C2(n7376), .ZN(P2_U3334) );
  NAND2_X1 U8825 ( .A1(n7180), .A2(n6643), .ZN(n7183) );
  AOI22_X1 U8826 ( .A1(n7649), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7648), .B2(
        n7181), .ZN(n7182) );
  INV_X1 U8827 ( .A(n9435), .ZN(n7281) );
  NAND2_X1 U8828 ( .A1(n9472), .A2(n7281), .ZN(n7902) );
  AOI21_X1 U8829 ( .B1(n7992), .B2(n7186), .A(n9010), .ZN(n9476) );
  INV_X1 U8830 ( .A(n9476), .ZN(n9474) );
  INV_X1 U8831 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7187) );
  OAI22_X1 U8832 ( .A1(n7852), .A2(n7188), .B1(n7848), .B2(n7187), .ZN(n7193)
         );
  NAND2_X1 U8833 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  NAND2_X1 U8834 ( .A1(n7404), .A2(n7191), .ZN(n9440) );
  OAI22_X1 U8835 ( .A1(n4272), .A2(n9440), .B1(n7636), .B2(n6612), .ZN(n7192)
         );
  INV_X1 U8836 ( .A(n9454), .ZN(n7900) );
  AOI21_X1 U8837 ( .B1(n7194), .B2(n7898), .A(n7901), .ZN(n7195) );
  XOR2_X1 U8838 ( .A(n7992), .B(n7195), .Z(n7196) );
  OAI222_X1 U8839 ( .A1(n9289), .A2(n7900), .B1(n9287), .B2(n7369), .C1(n9632), 
        .C2(n7196), .ZN(n9470) );
  INV_X1 U8840 ( .A(n9472), .ZN(n7374) );
  AOI211_X1 U8841 ( .C1(n9472), .C2(n7198), .A(n9458), .B(n9443), .ZN(n9471)
         );
  NAND2_X1 U8842 ( .A1(n9471), .A2(n9644), .ZN(n7201) );
  INV_X1 U8843 ( .A(n7199), .ZN(n7371) );
  AOI22_X1 U8844 ( .A1(n9648), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7371), .B2(
        n10031), .ZN(n7200) );
  OAI211_X1 U8845 ( .C1(n7374), .C2(n9638), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U8846 ( .B1(n9470), .B2(n10029), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8847 ( .B1(n9474), .B2(n9292), .A(n7203), .ZN(P1_U3279) );
  OAI211_X1 U8848 ( .C1(n7205), .C2(n7209), .A(n7204), .B(n9745), .ZN(n7207)
         );
  NAND2_X1 U8849 ( .A1(n7207), .A2(n7206), .ZN(n7379) );
  INV_X1 U8850 ( .A(n7379), .ZN(n7217) );
  XNOR2_X1 U8851 ( .A(n7208), .B(n7209), .ZN(n7381) );
  NAND2_X1 U8852 ( .A1(n7381), .A2(n9764), .ZN(n7216) );
  AOI211_X1 U8853 ( .C1(n7210), .C2(n7223), .A(n9826), .B(n4602), .ZN(n7380)
         );
  INV_X1 U8854 ( .A(n7210), .ZN(n7385) );
  NOR2_X1 U8855 ( .A1(n7385), .A2(n9762), .ZN(n7214) );
  OAI22_X1 U8856 ( .A1(n9757), .A2(n7212), .B1(n7211), .B2(n9755), .ZN(n7213)
         );
  AOI211_X1 U8857 ( .C1(n7380), .C2(n8634), .A(n7214), .B(n7213), .ZN(n7215)
         );
  OAI211_X1 U8858 ( .C1(n9766), .C2(n7217), .A(n7216), .B(n7215), .ZN(P2_U3284) );
  XOR2_X1 U8859 ( .A(n7230), .B(n7218), .Z(n7219) );
  AOI222_X1 U8860 ( .A1(n9745), .A2(n7219), .B1(n8282), .B2(n9740), .C1(n8284), 
        .C2(n9742), .ZN(n9834) );
  OAI22_X1 U8861 ( .A1(n9757), .A2(n7221), .B1(n7220), .B2(n9755), .ZN(n7225)
         );
  INV_X1 U8862 ( .A(n7222), .ZN(n7339) );
  INV_X1 U8863 ( .A(n7226), .ZN(n9836) );
  OAI211_X1 U8864 ( .C1(n7339), .C2(n9836), .A(n8603), .B(n7223), .ZN(n9833)
         );
  NOR2_X1 U8865 ( .A1(n9833), .A2(n8612), .ZN(n7224) );
  AOI211_X1 U8866 ( .C1(n8609), .C2(n7226), .A(n7225), .B(n7224), .ZN(n7232)
         );
  NAND2_X1 U8867 ( .A1(n7227), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U8868 ( .A1(n7333), .A2(n7228), .ZN(n7229) );
  XOR2_X1 U8869 ( .A(n7230), .B(n7229), .Z(n9839) );
  NAND2_X1 U8870 ( .A1(n9839), .A2(n9764), .ZN(n7231) );
  OAI211_X1 U8871 ( .C1(n9834), .C2(n9766), .A(n7232), .B(n7231), .ZN(P2_U3285) );
  AOI22_X1 U8872 ( .A1(n7234), .A2(n8603), .B1(n9812), .B2(n7233), .ZN(n7235)
         );
  OAI211_X1 U8873 ( .C1(n8704), .C2(n7237), .A(n7236), .B(n7235), .ZN(n7239)
         );
  NAND2_X1 U8874 ( .A1(n7239), .A2(n9855), .ZN(n7238) );
  OAI21_X1 U8875 ( .B1(n9855), .B2(n6439), .A(n7238), .ZN(P2_U3528) );
  NAND2_X1 U8876 ( .A1(n7239), .A2(n9840), .ZN(n7240) );
  OAI21_X1 U8877 ( .B1(n9840), .B2(n5155), .A(n7240), .ZN(P2_U3475) );
  INV_X1 U8878 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7241) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7241), .ZN(n9863) );
  NOR2_X1 U8881 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7242) );
  AOI21_X1 U8882 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7242), .ZN(n9866) );
  NOR2_X1 U8883 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7243) );
  AOI21_X1 U8884 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7243), .ZN(n9869) );
  NOR2_X1 U8885 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7244) );
  AOI21_X1 U8886 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7244), .ZN(n9872) );
  NOR2_X1 U8887 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7245) );
  AOI21_X1 U8888 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7245), .ZN(n9875) );
  NOR2_X1 U8889 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7251) );
  INV_X1 U8890 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9532) );
  XOR2_X1 U8891 ( .A(n9532), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10063) );
  NAND2_X1 U8892 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7249) );
  XOR2_X1 U8893 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10061) );
  NAND2_X1 U8894 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7247) );
  XNOR2_X1 U8895 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9518), .ZN(n10059) );
  AOI21_X1 U8896 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9856) );
  INV_X1 U8897 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9860) );
  NAND3_X1 U8898 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n9858) );
  OAI21_X1 U8899 ( .B1(n9856), .B2(n9860), .A(n9858), .ZN(n10058) );
  NAND2_X1 U8900 ( .A1(n10059), .A2(n10058), .ZN(n7246) );
  NAND2_X1 U8901 ( .A1(n7247), .A2(n7246), .ZN(n10060) );
  NAND2_X1 U8902 ( .A1(n10061), .A2(n10060), .ZN(n7248) );
  NAND2_X1 U8903 ( .A1(n7249), .A2(n7248), .ZN(n10062) );
  NOR2_X1 U8904 ( .A1(n10063), .A2(n10062), .ZN(n7250) );
  NOR2_X1 U8905 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  NOR2_X1 U8906 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7252), .ZN(n10047) );
  AND2_X1 U8907 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7252), .ZN(n10046) );
  NOR2_X1 U8908 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10046), .ZN(n7253) );
  NOR2_X1 U8909 ( .A1(n10047), .A2(n7253), .ZN(n7254) );
  NAND2_X1 U8910 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7254), .ZN(n7256) );
  XOR2_X1 U8911 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7254), .Z(n10045) );
  NAND2_X1 U8912 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10045), .ZN(n7255) );
  NAND2_X1 U8913 ( .A1(n7256), .A2(n7255), .ZN(n7257) );
  NAND2_X1 U8914 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7257), .ZN(n7259) );
  XOR2_X1 U8915 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7257), .Z(n10057) );
  NAND2_X1 U8916 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10057), .ZN(n7258) );
  NAND2_X1 U8917 ( .A1(n7259), .A2(n7258), .ZN(n7260) );
  NAND2_X1 U8918 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7260), .ZN(n7262) );
  XOR2_X1 U8919 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7260), .Z(n10056) );
  NAND2_X1 U8920 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10056), .ZN(n7261) );
  NAND2_X1 U8921 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  AND2_X1 U8922 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7263), .ZN(n7264) );
  INV_X1 U8923 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10055) );
  XNOR2_X1 U8924 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7263), .ZN(n10054) );
  NOR2_X1 U8925 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  NAND2_X1 U8926 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7265) );
  OAI21_X1 U8927 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7265), .ZN(n9883) );
  AOI21_X1 U8928 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9882), .ZN(n9881) );
  NAND2_X1 U8929 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7266) );
  OAI21_X1 U8930 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n7266), .ZN(n9880) );
  NOR2_X1 U8931 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  AOI21_X1 U8932 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9879), .ZN(n9878) );
  NOR2_X1 U8933 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7267) );
  AOI21_X1 U8934 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7267), .ZN(n9877) );
  NAND2_X1 U8935 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  OAI21_X1 U8936 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9876), .ZN(n9874) );
  NAND2_X1 U8937 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  OAI21_X1 U8938 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9873), .ZN(n9871) );
  NAND2_X1 U8939 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  OAI21_X1 U8940 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9870), .ZN(n9868) );
  NAND2_X1 U8941 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  OAI21_X1 U8942 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9867), .ZN(n9865) );
  NAND2_X1 U8943 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  OAI21_X1 U8944 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9864), .ZN(n9862) );
  NAND2_X1 U8945 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  OAI21_X1 U8946 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9861), .ZN(n10050) );
  NOR2_X1 U8947 ( .A1(n10051), .A2(n10050), .ZN(n7268) );
  NAND2_X1 U8948 ( .A1(n10051), .A2(n10050), .ZN(n10049) );
  OAI21_X1 U8949 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7268), .A(n10049), .ZN(
        n7270) );
  XNOR2_X1 U8950 ( .A(n8379), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7269) );
  XNOR2_X1 U8951 ( .A(n7270), .B(n7269), .ZN(ADD_1071_U4) );
  AND2_X1 U8952 ( .A1(n7271), .A2(n7272), .ZN(n7275) );
  INV_X1 U8953 ( .A(n7271), .ZN(n7274) );
  INV_X1 U8954 ( .A(n7272), .ZN(n7273) );
  NAND2_X1 U8955 ( .A1(n7286), .A2(n7808), .ZN(n7278) );
  NAND2_X1 U8956 ( .A1(n8928), .A2(n7824), .ZN(n7277) );
  NAND2_X1 U8957 ( .A1(n7278), .A2(n7277), .ZN(n7279) );
  XNOR2_X1 U8958 ( .A(n7279), .B(n7799), .ZN(n7359) );
  AND2_X1 U8959 ( .A1(n8928), .A2(n7801), .ZN(n7280) );
  AOI21_X1 U8960 ( .B1(n7286), .B2(n7824), .A(n7280), .ZN(n7357) );
  XNOR2_X1 U8961 ( .A(n7359), .B(n7357), .ZN(n7361) );
  XNOR2_X1 U8962 ( .A(n7362), .B(n7361), .ZN(n7288) );
  AND2_X1 U8963 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9591) );
  NOR2_X1 U8964 ( .A1(n8904), .A2(n7281), .ZN(n7282) );
  AOI211_X1 U8965 ( .C1(n8901), .C2(n8929), .A(n9591), .B(n7282), .ZN(n7283)
         );
  OAI21_X1 U8966 ( .B1(n8920), .B2(n7284), .A(n7283), .ZN(n7285) );
  AOI21_X1 U8967 ( .B1(n7286), .B2(n8894), .A(n7285), .ZN(n7287) );
  OAI21_X1 U8968 ( .B1(n7288), .B2(n8923), .A(n7287), .ZN(P1_U3234) );
  NOR2_X1 U8969 ( .A1(n7290), .A2(n7289), .ZN(n7292) );
  NOR2_X1 U8970 ( .A1(n7292), .A2(n7291), .ZN(n8952) );
  INV_X1 U8971 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9975) );
  AOI211_X1 U8972 ( .C1(n7293), .C2(n9975), .A(n8953), .B(n9578), .ZN(n7299)
         );
  XNOR2_X1 U8973 ( .A(n8958), .B(n8957), .ZN(n7295) );
  INV_X1 U8974 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7574) );
  NOR2_X1 U8975 ( .A1(n7574), .A2(n7295), .ZN(n8959) );
  AOI211_X1 U8976 ( .C1(n7295), .C2(n7574), .A(n8959), .B(n9536), .ZN(n7296)
         );
  AOI21_X1 U8977 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9619), .A(n7296), .ZN(
        n7297) );
  NAND2_X1 U8978 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8915) );
  OAI211_X1 U8979 ( .C1(n9613), .C2(n8958), .A(n7297), .B(n8915), .ZN(n7298)
         );
  OR2_X1 U8980 ( .A1(n7299), .A2(n7298), .ZN(P1_U3256) );
  XNOR2_X1 U8981 ( .A(n7301), .B(n7300), .ZN(n7302) );
  XNOR2_X1 U8982 ( .A(n7303), .B(n7302), .ZN(n7309) );
  INV_X1 U8983 ( .A(n8264), .ZN(n8253) );
  OAI22_X1 U8984 ( .A1(n7304), .A2(n8621), .B1(n7446), .B2(n8619), .ZN(n7316)
         );
  AOI21_X1 U8985 ( .B1(n8253), .B2(n7316), .A(n7305), .ZN(n7306) );
  OAI21_X1 U8986 ( .B1(n7322), .B2(n8251), .A(n7306), .ZN(n7307) );
  AOI21_X1 U8987 ( .B1(n7503), .B2(n8238), .A(n7307), .ZN(n7308) );
  OAI21_X1 U8988 ( .B1(n7309), .B2(n8244), .A(n7308), .ZN(P2_U3236) );
  INV_X1 U8989 ( .A(n7771), .ZN(n7387) );
  AOI22_X1 U8990 ( .A1(n7310), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8780), .ZN(n7311) );
  OAI21_X1 U8991 ( .B1(n7387), .B2(n8783), .A(n7311), .ZN(P2_U3332) );
  NAND2_X1 U8992 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  NAND2_X1 U8993 ( .A1(n7315), .A2(n7314), .ZN(n7317) );
  AOI21_X1 U8994 ( .B1(n7317), .B2(n9745), .A(n7316), .ZN(n7506) );
  NAND2_X1 U8995 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  NAND2_X1 U8996 ( .A1(n7484), .A2(n7320), .ZN(n7504) );
  INV_X1 U8997 ( .A(n7504), .ZN(n7321) );
  NAND2_X1 U8998 ( .A1(n7321), .A2(n9764), .ZN(n7329) );
  OAI22_X1 U8999 ( .A1(n9757), .A2(n7323), .B1(n7322), .B2(n9755), .ZN(n7327)
         );
  AOI21_X1 U9000 ( .B1(n7324), .B2(n7503), .A(n9826), .ZN(n7325) );
  NAND2_X1 U9001 ( .A1(n4294), .A2(n7325), .ZN(n7505) );
  NOR2_X1 U9002 ( .A1(n7505), .A2(n8612), .ZN(n7326) );
  AOI211_X1 U9003 ( .C1(n8609), .C2(n7503), .A(n7327), .B(n7326), .ZN(n7328)
         );
  OAI211_X1 U9004 ( .C1(n9766), .C2(n7506), .A(n7329), .B(n7328), .ZN(P2_U3283) );
  XOR2_X1 U9005 ( .A(n7330), .B(n7334), .Z(n7337) );
  OAI22_X1 U9006 ( .A1(n7332), .A2(n8621), .B1(n7331), .B2(n8619), .ZN(n7336)
         );
  OAI21_X1 U9007 ( .B1(n7227), .B2(n7334), .A(n7333), .ZN(n7459) );
  NOR2_X1 U9008 ( .A1(n7459), .A2(n8626), .ZN(n7335) );
  AOI211_X1 U9009 ( .C1(n7337), .C2(n9745), .A(n7336), .B(n7335), .ZN(n7458)
         );
  INV_X1 U9010 ( .A(n7338), .ZN(n7340) );
  AOI21_X1 U9011 ( .B1(n7455), .B2(n7340), .A(n7339), .ZN(n7456) );
  INV_X1 U9012 ( .A(n7341), .ZN(n7342) );
  AOI22_X1 U9013 ( .A1(n9766), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7342), .B2(
        n8570), .ZN(n7343) );
  OAI21_X1 U9014 ( .B1(n9762), .B2(n7344), .A(n7343), .ZN(n7346) );
  NOR2_X1 U9015 ( .A1(n7459), .A2(n8637), .ZN(n7345) );
  AOI211_X1 U9016 ( .C1(n7456), .C2(n9759), .A(n7346), .B(n7345), .ZN(n7347)
         );
  OAI21_X1 U9017 ( .B1(n7458), .B2(n9766), .A(n7347), .ZN(P2_U3286) );
  NAND2_X1 U9018 ( .A1(n9472), .A2(n7808), .ZN(n7349) );
  NAND2_X1 U9019 ( .A1(n9435), .A2(n7824), .ZN(n7348) );
  NAND2_X1 U9020 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  XNOR2_X1 U9021 ( .A(n7350), .B(n7822), .ZN(n7352) );
  AND2_X1 U9022 ( .A1(n9435), .A2(n7801), .ZN(n7351) );
  AOI21_X1 U9023 ( .B1(n9472), .B2(n7824), .A(n7351), .ZN(n7353) );
  NAND2_X1 U9024 ( .A1(n7352), .A2(n7353), .ZN(n7388) );
  INV_X1 U9025 ( .A(n7352), .ZN(n7355) );
  INV_X1 U9026 ( .A(n7353), .ZN(n7354) );
  NAND2_X1 U9027 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  AND2_X1 U9028 ( .A1(n7388), .A2(n7356), .ZN(n7364) );
  INV_X1 U9029 ( .A(n7357), .ZN(n7358) );
  AND2_X1 U9030 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  NAND2_X1 U9031 ( .A1(n7363), .A2(n7364), .ZN(n7389) );
  OAI21_X1 U9032 ( .B1(n7364), .B2(n4265), .A(n7389), .ZN(n7365) );
  NAND2_X1 U9033 ( .A1(n7365), .A2(n8898), .ZN(n7373) );
  INV_X1 U9034 ( .A(n7366), .ZN(n7367) );
  AOI21_X1 U9035 ( .B1(n8918), .B2(n9454), .A(n7367), .ZN(n7368) );
  OAI21_X1 U9036 ( .B1(n7369), .B2(n8916), .A(n7368), .ZN(n7370) );
  AOI21_X1 U9037 ( .B1(n7371), .B2(n8907), .A(n7370), .ZN(n7372) );
  OAI211_X1 U9038 ( .C1(n7374), .C2(n8910), .A(n7373), .B(n7372), .ZN(P1_U3222) );
  INV_X1 U9039 ( .A(n7752), .ZN(n7378) );
  OAI222_X1 U9040 ( .A1(n7376), .A2(n10016), .B1(n8783), .B2(n7378), .C1(
        P2_U3152), .C2(n7375), .ZN(P2_U3333) );
  OAI222_X1 U9041 ( .A1(n8121), .A2(n7753), .B1(n9402), .B2(n7378), .C1(n7377), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  AOI211_X1 U9042 ( .C1(n7381), .C2(n9838), .A(n7380), .B(n7379), .ZN(n7383)
         );
  MUX2_X1 U9043 ( .A(n6819), .B(n7383), .S(n9855), .Z(n7382) );
  OAI21_X1 U9044 ( .B1(n7385), .B2(n8719), .A(n7382), .ZN(P2_U3532) );
  INV_X1 U9045 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9995) );
  MUX2_X1 U9046 ( .A(n9995), .B(n7383), .S(n9840), .Z(n7384) );
  OAI21_X1 U9047 ( .B1(n7385), .B2(n8770), .A(n7384), .ZN(P2_U3487) );
  NAND2_X1 U9048 ( .A1(n7390), .A2(n6643), .ZN(n7393) );
  AOI22_X1 U9049 ( .A1(n7649), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7648), .B2(
        n7391), .ZN(n7392) );
  NAND2_X1 U9050 ( .A1(n9442), .A2(n7808), .ZN(n7395) );
  NAND2_X1 U9051 ( .A1(n9454), .A2(n7824), .ZN(n7394) );
  NAND2_X1 U9052 ( .A1(n7395), .A2(n7394), .ZN(n7396) );
  XNOR2_X1 U9053 ( .A(n7396), .B(n7822), .ZN(n7398) );
  AND2_X1 U9054 ( .A1(n9454), .A2(n7801), .ZN(n7397) );
  AOI21_X1 U9055 ( .B1(n9442), .B2(n7824), .A(n7397), .ZN(n7399) );
  AND2_X1 U9056 ( .A1(n7398), .A2(n7399), .ZN(n7555) );
  INV_X1 U9057 ( .A(n7398), .ZN(n7401) );
  INV_X1 U9058 ( .A(n7399), .ZN(n7400) );
  NAND2_X1 U9059 ( .A1(n7401), .A2(n7400), .ZN(n7554) );
  NAND2_X1 U9060 ( .A1(n4784), .A2(n7554), .ZN(n7402) );
  XNOR2_X1 U9061 ( .A(n7556), .B(n7402), .ZN(n7415) );
  INV_X1 U9062 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9063 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  AND2_X1 U9064 ( .A1(n7576), .A2(n7405), .ZN(n10032) );
  NAND2_X1 U9065 ( .A1(n7797), .A2(n10032), .ZN(n7409) );
  NAND2_X1 U9066 ( .A1(n7633), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7408) );
  NAND2_X1 U9067 ( .A1(n7813), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U9068 ( .A1(n7853), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7406) );
  NAND4_X1 U9069 ( .A1(n7409), .A2(n7408), .A3(n7407), .A4(n7406), .ZN(n9436)
         );
  NOR2_X1 U9070 ( .A1(n8904), .A2(n9286), .ZN(n7410) );
  AOI211_X1 U9071 ( .C1(n8901), .C2(n9435), .A(n7411), .B(n7410), .ZN(n7412)
         );
  OAI21_X1 U9072 ( .B1(n8920), .B2(n9440), .A(n7412), .ZN(n7413) );
  AOI21_X1 U9073 ( .B1(n9442), .B2(n8894), .A(n7413), .ZN(n7414) );
  OAI21_X1 U9074 ( .B1(n7415), .B2(n8923), .A(n7414), .ZN(P1_U3232) );
  NOR2_X1 U9075 ( .A1(n7417), .A2(n7416), .ZN(n7469) );
  XNOR2_X1 U9076 ( .A(n7470), .B(n7469), .ZN(n7418) );
  NOR2_X1 U9077 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7418), .ZN(n7471) );
  AOI21_X1 U9078 ( .B1(n7418), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7471), .ZN(
        n7428) );
  INV_X1 U9079 ( .A(n7419), .ZN(n7421) );
  XNOR2_X1 U9080 ( .A(n7463), .B(n7464), .ZN(n7422) );
  NOR2_X1 U9081 ( .A1(n8713), .A2(n7422), .ZN(n7465) );
  AOI211_X1 U9082 ( .C1(n7422), .C2(n8713), .A(n7465), .B(n9418), .ZN(n7423)
         );
  INV_X1 U9083 ( .A(n7423), .ZN(n7427) );
  AND2_X1 U9084 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7425) );
  NOR2_X1 U9085 ( .A1(n9726), .A2(n7464), .ZN(n7424) );
  AOI211_X1 U9086 ( .C1(n9417), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7425), .B(
        n7424), .ZN(n7426) );
  OAI211_X1 U9087 ( .C1(n7428), .C2(n8370), .A(n7427), .B(n7426), .ZN(P2_U3260) );
  XOR2_X1 U9088 ( .A(n7429), .B(n7430), .Z(n7436) );
  OAI22_X1 U9089 ( .A1(n8622), .A2(n8619), .B1(n7431), .B2(n8621), .ZN(n7490)
         );
  AOI21_X1 U9090 ( .B1(n8253), .B2(n7490), .A(n7432), .ZN(n7433) );
  OAI21_X1 U9091 ( .B1(n7494), .B2(n8251), .A(n7433), .ZN(n7434) );
  AOI21_X1 U9092 ( .B1(n7493), .B2(n8238), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9093 ( .B1(n7436), .B2(n8244), .A(n7435), .ZN(P2_U3217) );
  INV_X1 U9094 ( .A(n7789), .ZN(n7439) );
  AOI22_X1 U9095 ( .A1(n7437), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8780), .ZN(n7438) );
  OAI21_X1 U9096 ( .B1(n7439), .B2(n8783), .A(n7438), .ZN(P2_U3331) );
  OAI222_X1 U9097 ( .A1(n9402), .A2(n7439), .B1(n4278), .B2(P1_U3084), .C1(
        n7790), .C2(n9404), .ZN(P1_U3326) );
  OAI21_X1 U9098 ( .B1(n7441), .B2(n7443), .A(n7440), .ZN(n8712) );
  INV_X1 U9099 ( .A(n8712), .ZN(n7454) );
  NAND3_X1 U9100 ( .A1(n7487), .A2(n7443), .A3(n7442), .ZN(n7444) );
  AND3_X1 U9101 ( .A1(n7445), .A2(n9745), .A3(n7444), .ZN(n7447) );
  OAI22_X1 U9102 ( .A1(n8595), .A2(n8619), .B1(n7446), .B2(n8621), .ZN(n8261)
         );
  OR2_X1 U9103 ( .A1(n7447), .A2(n8261), .ZN(n8710) );
  AOI211_X1 U9104 ( .C1(n7448), .C2(n7492), .A(n9826), .B(n4597), .ZN(n8711)
         );
  NAND2_X1 U9105 ( .A1(n8711), .A2(n8634), .ZN(n7451) );
  INV_X1 U9106 ( .A(n7449), .ZN(n8267) );
  AOI22_X1 U9107 ( .A1(n9766), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8267), .B2(
        n8570), .ZN(n7450) );
  OAI211_X1 U9108 ( .C1(n8766), .C2(n9762), .A(n7451), .B(n7450), .ZN(n7452)
         );
  AOI21_X1 U9109 ( .B1(n8710), .B2(n9757), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9110 ( .B1(n7454), .B2(n8584), .A(n7453), .ZN(P2_U3281) );
  AOI22_X1 U9111 ( .A1(n7456), .A2(n8603), .B1(n9812), .B2(n7455), .ZN(n7457)
         );
  OAI211_X1 U9112 ( .C1(n8704), .C2(n7459), .A(n7458), .B(n7457), .ZN(n7461)
         );
  NAND2_X1 U9113 ( .A1(n7461), .A2(n9855), .ZN(n7460) );
  OAI21_X1 U9114 ( .B1(n9855), .B2(n6691), .A(n7460), .ZN(P2_U3530) );
  NAND2_X1 U9115 ( .A1(n7461), .A2(n9840), .ZN(n7462) );
  OAI21_X1 U9116 ( .B1(n9840), .B2(n5204), .A(n7462), .ZN(P2_U3481) );
  NOR2_X1 U9117 ( .A1(n7464), .A2(n7463), .ZN(n7466) );
  XNOR2_X1 U9118 ( .A(n8340), .B(n8708), .ZN(n7467) );
  NAND2_X1 U9119 ( .A1(n7467), .A2(n7468), .ZN(n8339) );
  OAI21_X1 U9120 ( .B1(n7468), .B2(n7467), .A(n8339), .ZN(n7481) );
  NOR2_X1 U9121 ( .A1(n7470), .A2(n7469), .ZN(n7472) );
  NOR2_X1 U9122 ( .A1(n7472), .A2(n7471), .ZN(n7475) );
  NAND2_X1 U9123 ( .A1(n8340), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8335) );
  INV_X1 U9124 ( .A(n8335), .ZN(n7473) );
  AOI21_X1 U9125 ( .B1(n8631), .B2(n7479), .A(n7473), .ZN(n7474) );
  NAND2_X1 U9126 ( .A1(n7474), .A2(n7475), .ZN(n8334) );
  OAI211_X1 U9127 ( .C1(n7475), .C2(n7474), .A(n9722), .B(n8334), .ZN(n7478)
         );
  NAND2_X1 U9128 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8200) );
  INV_X1 U9129 ( .A(n8200), .ZN(n7476) );
  AOI21_X1 U9130 ( .B1(n9417), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7476), .ZN(
        n7477) );
  OAI211_X1 U9131 ( .C1(n9726), .C2(n7479), .A(n7478), .B(n7477), .ZN(n7480)
         );
  AOI21_X1 U9132 ( .B1(n9724), .B2(n7481), .A(n7480), .ZN(n7482) );
  INV_X1 U9133 ( .A(n7482), .ZN(P2_U3261) );
  NAND2_X1 U9134 ( .A1(n7484), .A2(n7483), .ZN(n7486) );
  XNOR2_X1 U9135 ( .A(n7486), .B(n7485), .ZN(n8717) );
  INV_X1 U9136 ( .A(n8717), .ZN(n7500) );
  INV_X1 U9137 ( .A(n7487), .ZN(n7488) );
  AOI211_X1 U9138 ( .C1(n5273), .C2(n7489), .A(n8566), .B(n7488), .ZN(n7491)
         );
  OR2_X1 U9139 ( .A1(n7491), .A2(n7490), .ZN(n8715) );
  NAND2_X1 U9140 ( .A1(n8715), .A2(n9757), .ZN(n7499) );
  AOI211_X1 U9141 ( .C1(n7493), .C2(n4294), .A(n9826), .B(n4598), .ZN(n8716)
         );
  NOR2_X1 U9142 ( .A1(n8771), .A2(n9762), .ZN(n7497) );
  OAI22_X1 U9143 ( .A1(n9757), .A2(n7495), .B1(n7494), .B2(n9755), .ZN(n7496)
         );
  AOI211_X1 U9144 ( .C1(n8716), .C2(n8634), .A(n7497), .B(n7496), .ZN(n7498)
         );
  OAI211_X1 U9145 ( .C1(n7500), .C2(n8584), .A(n7499), .B(n7498), .ZN(P2_U3282) );
  INV_X1 U9146 ( .A(n7805), .ZN(n8124) );
  NAND2_X1 U9147 ( .A1(n8780), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7501) );
  OAI211_X1 U9148 ( .C1(n8124), .C2(n8783), .A(n7502), .B(n7501), .ZN(P2_U3330) );
  INV_X1 U9149 ( .A(n7503), .ZN(n7513) );
  INV_X1 U9150 ( .A(n9838), .ZN(n9815) );
  OR2_X1 U9151 ( .A1(n7504), .A2(n9815), .ZN(n7508) );
  AND2_X1 U9152 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  AND2_X1 U9153 ( .A1(n7508), .A2(n7507), .ZN(n7511) );
  MUX2_X1 U9154 ( .A(n7511), .B(n5253), .S(n9853), .Z(n7509) );
  OAI21_X1 U9155 ( .B1(n7513), .B2(n8719), .A(n7509), .ZN(P2_U3533) );
  INV_X1 U9156 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7510) );
  MUX2_X1 U9157 ( .A(n7511), .B(n7510), .S(n5900), .Z(n7512) );
  OAI21_X1 U9158 ( .B1(n7513), .B2(n8770), .A(n7512), .ZN(P2_U3490) );
  INV_X1 U9159 ( .A(n7955), .ZN(n8784) );
  OAI222_X1 U9160 ( .A1(n9402), .A2(n8784), .B1(n7514), .B2(P1_U3084), .C1(
        n7956), .C2(n8121), .ZN(P1_U3324) );
  INV_X1 U9161 ( .A(n7515), .ZN(n7542) );
  INV_X1 U9162 ( .A(n7516), .ZN(n7522) );
  XNOR2_X1 U9163 ( .A(n8424), .B(n7527), .ZN(n7517) );
  NOR2_X1 U9164 ( .A1(n8437), .A2(n7525), .ZN(n7518) );
  NAND2_X1 U9165 ( .A1(n7517), .A2(n7518), .ZN(n7524) );
  INV_X1 U9166 ( .A(n7517), .ZN(n7520) );
  INV_X1 U9167 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9168 ( .A1(n7520), .A2(n7519), .ZN(n7521) );
  NOR2_X1 U9169 ( .A1(n7526), .A2(n7525), .ZN(n7528) );
  XNOR2_X1 U9170 ( .A(n7528), .B(n7527), .ZN(n7530) );
  INV_X1 U9171 ( .A(n7530), .ZN(n7531) );
  NOR3_X1 U9172 ( .A1(n8406), .A2(n8238), .A3(n7531), .ZN(n7529) );
  AOI21_X1 U9173 ( .B1(n8406), .B2(n7531), .A(n7529), .ZN(n7537) );
  NOR3_X1 U9174 ( .A1(n8406), .A2(n7530), .A3(n8238), .ZN(n7534) );
  NOR2_X1 U9175 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  OAI21_X1 U9176 ( .B1(n8406), .B2(n8270), .A(n8244), .ZN(n7535) );
  OAI211_X1 U9177 ( .C1(n7538), .C2(n7537), .A(n7536), .B(n7535), .ZN(n7541)
         );
  INV_X1 U9178 ( .A(n8408), .ZN(n7539) );
  AOI22_X1 U9179 ( .A1(n7539), .A2(n8266), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7540) );
  OAI211_X1 U9180 ( .C1(n7542), .C2(n8264), .A(n7541), .B(n7540), .ZN(P2_U3222) );
  NAND2_X1 U9181 ( .A1(n7543), .A2(n6643), .ZN(n7545) );
  OR2_X1 U9182 ( .A1(n7957), .A2(n10002), .ZN(n7544) );
  NAND2_X1 U9183 ( .A1(n7737), .A2(n9958), .ZN(n7546) );
  NAND2_X1 U9184 ( .A1(n9140), .A2(n7797), .ZN(n7552) );
  INV_X1 U9185 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9186 ( .A1(n7813), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9187 ( .A1(n7853), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7547) );
  OAI211_X1 U9188 ( .C1(n7852), .C2(n7549), .A(n7548), .B(n7547), .ZN(n7550)
         );
  INV_X1 U9189 ( .A(n7550), .ZN(n7551) );
  AOI22_X1 U9190 ( .A1(n9323), .A2(n4256), .B1(n7801), .B2(n9164), .ZN(n7751)
         );
  AOI22_X1 U9191 ( .A1(n9323), .A2(n7793), .B1(n7824), .B2(n9164), .ZN(n7553)
         );
  XNOR2_X1 U9192 ( .A(n7553), .B(n7799), .ZN(n7750) );
  NAND2_X1 U9193 ( .A1(n7557), .A2(n6643), .ZN(n7560) );
  AOI22_X1 U9194 ( .A1(n7558), .A2(n7648), .B1(n7649), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9195 ( .A1(n10034), .A2(n7808), .ZN(n7562) );
  NAND2_X1 U9196 ( .A1(n9436), .A2(n7824), .ZN(n7561) );
  NAND2_X1 U9197 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  XNOR2_X1 U9198 ( .A(n7563), .B(n7799), .ZN(n7566) );
  NAND2_X1 U9199 ( .A1(n10034), .A2(n4256), .ZN(n7565) );
  NAND2_X1 U9200 ( .A1(n9436), .A2(n7801), .ZN(n7564) );
  NAND2_X1 U9201 ( .A1(n7565), .A2(n7564), .ZN(n8798) );
  NAND2_X1 U9202 ( .A1(n7567), .A2(n6643), .ZN(n7572) );
  OAI22_X1 U9203 ( .A1(n8958), .A2(n7569), .B1(n7957), .B2(n7568), .ZN(n7570)
         );
  INV_X1 U9204 ( .A(n7570), .ZN(n7571) );
  NAND2_X1 U9205 ( .A1(n9371), .A2(n7808), .ZN(n7581) );
  INV_X1 U9206 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7573) );
  OAI22_X1 U9207 ( .A1(n7852), .A2(n7574), .B1(n7848), .B2(n7573), .ZN(n7579)
         );
  NAND2_X1 U9208 ( .A1(n7576), .A2(n7575), .ZN(n7577) );
  NAND2_X1 U9209 ( .A1(n7594), .A2(n7577), .ZN(n9280) );
  OAI22_X1 U9210 ( .A1(n4272), .A2(n9280), .B1(n7636), .B2(n9975), .ZN(n7578)
         );
  NAND2_X1 U9211 ( .A1(n9453), .A2(n7824), .ZN(n7580) );
  NAND2_X1 U9212 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  XNOR2_X1 U9213 ( .A(n7582), .B(n7822), .ZN(n7586) );
  NAND2_X1 U9214 ( .A1(n9371), .A2(n4256), .ZN(n7584) );
  NAND2_X1 U9215 ( .A1(n7801), .A2(n9453), .ZN(n7583) );
  NAND2_X1 U9216 ( .A1(n7584), .A2(n7583), .ZN(n8914) );
  NAND2_X1 U9217 ( .A1(n8912), .A2(n8914), .ZN(n7589) );
  INV_X1 U9218 ( .A(n7586), .ZN(n7587) );
  NAND2_X1 U9219 ( .A1(n7588), .A2(n7587), .ZN(n8911) );
  NAND2_X1 U9220 ( .A1(n7589), .A2(n8911), .ZN(n8846) );
  NAND2_X1 U9221 ( .A1(n7590), .A2(n6643), .ZN(n7592) );
  AOI22_X1 U9222 ( .A1(n8975), .A2(n7648), .B1(n7649), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9223 ( .A1(n9365), .A2(n7793), .ZN(n7601) );
  INV_X1 U9224 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9225 ( .A1(n7594), .A2(n7593), .ZN(n7595) );
  AND2_X1 U9226 ( .A1(n7611), .A2(n7595), .ZN(n9270) );
  NAND2_X1 U9227 ( .A1(n9270), .A2(n7797), .ZN(n7599) );
  NAND2_X1 U9228 ( .A1(n7633), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7598) );
  NAND2_X1 U9229 ( .A1(n7813), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U9230 ( .A1(n7853), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7596) );
  NAND4_X1 U9231 ( .A1(n7599), .A2(n7598), .A3(n7597), .A4(n7596), .ZN(n9014)
         );
  NAND2_X1 U9232 ( .A1(n9014), .A2(n7824), .ZN(n7600) );
  NAND2_X1 U9233 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  XNOR2_X1 U9234 ( .A(n7602), .B(n7822), .ZN(n7606) );
  AND2_X1 U9235 ( .A1(n9014), .A2(n7801), .ZN(n7603) );
  AOI21_X1 U9236 ( .B1(n9365), .B2(n7824), .A(n7603), .ZN(n7605) );
  XNOR2_X1 U9237 ( .A(n7606), .B(n7605), .ZN(n8849) );
  NAND2_X1 U9238 ( .A1(n7606), .A2(n7605), .ZN(n7607) );
  NAND2_X1 U9239 ( .A1(n7608), .A2(n6643), .ZN(n7610) );
  AOI22_X1 U9240 ( .A1(n8987), .A2(n7648), .B1(n7649), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9241 ( .A1(n9359), .A2(n7808), .ZN(n7619) );
  NAND2_X1 U9242 ( .A1(n7611), .A2(n8857), .ZN(n7612) );
  NAND2_X1 U9243 ( .A1(n7631), .A2(n7612), .ZN(n9247) );
  NAND2_X1 U9244 ( .A1(n7853), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7613) );
  OAI21_X1 U9245 ( .B1(n9247), .B2(n4272), .A(n7613), .ZN(n7617) );
  INV_X1 U9246 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7615) );
  INV_X1 U9247 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7614) );
  OAI22_X1 U9248 ( .A1(n7852), .A2(n7615), .B1(n7848), .B2(n7614), .ZN(n7616)
         );
  NAND2_X1 U9249 ( .A1(n9015), .A2(n7824), .ZN(n7618) );
  NAND2_X1 U9250 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  XNOR2_X1 U9251 ( .A(n7620), .B(n7799), .ZN(n7622) );
  AND2_X1 U9252 ( .A1(n9015), .A2(n7801), .ZN(n7621) );
  AOI21_X1 U9253 ( .B1(n9359), .B2(n4256), .A(n7621), .ZN(n7623) );
  XNOR2_X1 U9254 ( .A(n7622), .B(n7623), .ZN(n8855) );
  INV_X1 U9255 ( .A(n7622), .ZN(n7624) );
  NAND2_X1 U9256 ( .A1(n7624), .A2(n7623), .ZN(n7625) );
  NAND2_X1 U9257 ( .A1(n7626), .A2(n7625), .ZN(n7642) );
  NAND2_X1 U9258 ( .A1(n7627), .A2(n6643), .ZN(n7629) );
  AOI22_X1 U9259 ( .A1(n8988), .A2(n7648), .B1(n7649), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7628) );
  NAND2_X1 U9260 ( .A1(n9354), .A2(n7808), .ZN(n7638) );
  INV_X1 U9261 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9234) );
  INV_X1 U9262 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U9263 ( .A1(n7631), .A2(n7630), .ZN(n7632) );
  NAND2_X1 U9264 ( .A1(n7653), .A2(n7632), .ZN(n9233) );
  OR2_X1 U9265 ( .A1(n9233), .A2(n4272), .ZN(n7635) );
  AOI22_X1 U9266 ( .A1(n7633), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7813), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n7634) );
  OAI211_X1 U9267 ( .C1(n7636), .C2(n9234), .A(n7635), .B(n7634), .ZN(n9017)
         );
  NAND2_X1 U9268 ( .A1(n9017), .A2(n4256), .ZN(n7637) );
  NAND2_X1 U9269 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  XNOR2_X1 U9270 ( .A(n7639), .B(n7822), .ZN(n7643) );
  NAND2_X1 U9271 ( .A1(n7642), .A2(n7643), .ZN(n8887) );
  NAND2_X1 U9272 ( .A1(n9354), .A2(n4256), .ZN(n7641) );
  NAND2_X1 U9273 ( .A1(n9017), .A2(n7801), .ZN(n7640) );
  NAND2_X1 U9274 ( .A1(n7641), .A2(n7640), .ZN(n8890) );
  NAND2_X1 U9275 ( .A1(n8887), .A2(n8890), .ZN(n7646) );
  INV_X1 U9276 ( .A(n7642), .ZN(n7645) );
  INV_X1 U9277 ( .A(n7643), .ZN(n7644) );
  NAND2_X1 U9278 ( .A1(n7645), .A2(n7644), .ZN(n8888) );
  NAND2_X1 U9279 ( .A1(n7646), .A2(n8888), .ZN(n8817) );
  NAND2_X1 U9280 ( .A1(n7647), .A2(n6643), .ZN(n7651) );
  AOI22_X1 U9281 ( .A1(n7649), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9193), .B2(
        n7648), .ZN(n7650) );
  NAND2_X1 U9282 ( .A1(n9349), .A2(n7793), .ZN(n7662) );
  INV_X1 U9283 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9284 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  NAND2_X1 U9285 ( .A1(n7673), .A2(n7654), .ZN(n9221) );
  OR2_X1 U9286 ( .A1(n9221), .A2(n4272), .ZN(n7660) );
  INV_X1 U9287 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U9288 ( .A1(n7853), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U9289 ( .A1(n7813), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7656) );
  OAI211_X1 U9290 ( .C1(n7852), .C2(n8989), .A(n7657), .B(n7656), .ZN(n7658)
         );
  INV_X1 U9291 ( .A(n7658), .ZN(n7659) );
  NAND2_X1 U9292 ( .A1(n7660), .A2(n7659), .ZN(n9018) );
  NAND2_X1 U9293 ( .A1(n9018), .A2(n7824), .ZN(n7661) );
  NAND2_X1 U9294 ( .A1(n7662), .A2(n7661), .ZN(n7663) );
  XNOR2_X1 U9295 ( .A(n7663), .B(n7822), .ZN(n7667) );
  AND2_X1 U9296 ( .A1(n9018), .A2(n7801), .ZN(n7664) );
  AOI21_X1 U9297 ( .B1(n9349), .B2(n7824), .A(n7664), .ZN(n7666) );
  XNOR2_X1 U9298 ( .A(n7667), .B(n7666), .ZN(n8818) );
  NAND2_X1 U9299 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U9300 ( .A1(n7669), .A2(n6643), .ZN(n7672) );
  OR2_X1 U9301 ( .A1(n7957), .A2(n7670), .ZN(n7671) );
  NAND2_X1 U9302 ( .A1(n9344), .A2(n7793), .ZN(n7681) );
  NAND2_X1 U9303 ( .A1(n7673), .A2(n10001), .ZN(n7674) );
  NAND2_X1 U9304 ( .A1(n7694), .A2(n7674), .ZN(n9208) );
  OR2_X1 U9305 ( .A1(n9208), .A2(n4272), .ZN(n7679) );
  INV_X1 U9306 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U9307 ( .A1(n7813), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U9308 ( .A1(n7853), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7675) );
  OAI211_X1 U9309 ( .C1(n7852), .C2(n9988), .A(n7676), .B(n7675), .ZN(n7677)
         );
  INV_X1 U9310 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9311 ( .A1(n7679), .A2(n7678), .ZN(n9020) );
  NAND2_X1 U9312 ( .A1(n9020), .A2(n4256), .ZN(n7680) );
  NAND2_X1 U9313 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  XNOR2_X1 U9314 ( .A(n7682), .B(n7799), .ZN(n7684) );
  AND2_X1 U9315 ( .A1(n9020), .A2(n7801), .ZN(n7683) );
  AOI21_X1 U9316 ( .B1(n9344), .B2(n4256), .A(n7683), .ZN(n7685) );
  XNOR2_X1 U9317 ( .A(n7684), .B(n7685), .ZN(n8871) );
  INV_X1 U9318 ( .A(n7684), .ZN(n7686) );
  NAND2_X1 U9319 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  NAND2_X1 U9320 ( .A1(n7689), .A2(n6643), .ZN(n7692) );
  OR2_X1 U9321 ( .A1(n7957), .A2(n7690), .ZN(n7691) );
  NAND2_X1 U9322 ( .A1(n9339), .A2(n7793), .ZN(n7703) );
  NAND2_X1 U9323 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  AND2_X1 U9324 ( .A1(n7716), .A2(n7695), .ZN(n9191) );
  NAND2_X1 U9325 ( .A1(n9191), .A2(n7797), .ZN(n7701) );
  INV_X1 U9326 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U9327 ( .A1(n7813), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9328 ( .A1(n7853), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7696) );
  OAI211_X1 U9329 ( .C1(n7852), .C2(n7698), .A(n7697), .B(n7696), .ZN(n7699)
         );
  INV_X1 U9330 ( .A(n7699), .ZN(n7700) );
  NAND2_X1 U9331 ( .A1(n7701), .A2(n7700), .ZN(n9022) );
  NAND2_X1 U9332 ( .A1(n9022), .A2(n4256), .ZN(n7702) );
  NAND2_X1 U9333 ( .A1(n7703), .A2(n7702), .ZN(n7704) );
  XNOR2_X1 U9334 ( .A(n7704), .B(n7799), .ZN(n7706) );
  AND2_X1 U9335 ( .A1(n9022), .A2(n7801), .ZN(n7705) );
  AOI21_X1 U9336 ( .B1(n9339), .B2(n4256), .A(n7705), .ZN(n7707) );
  XNOR2_X1 U9337 ( .A(n7706), .B(n7707), .ZN(n8833) );
  NAND2_X1 U9338 ( .A1(n8832), .A2(n8833), .ZN(n7710) );
  INV_X1 U9339 ( .A(n7706), .ZN(n7708) );
  NAND2_X1 U9340 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  NAND2_X1 U9341 ( .A1(n7711), .A2(n6643), .ZN(n7714) );
  OR2_X1 U9342 ( .A1(n7957), .A2(n7712), .ZN(n7713) );
  INV_X1 U9343 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U9344 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  NAND2_X1 U9345 ( .A1(n7735), .A2(n7717), .ZN(n9177) );
  OR2_X1 U9346 ( .A1(n9177), .A2(n4272), .ZN(n7723) );
  INV_X1 U9347 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9348 ( .A1(n7853), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U9349 ( .A1(n7813), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7718) );
  OAI211_X1 U9350 ( .C1(n7852), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7721)
         );
  INV_X1 U9351 ( .A(n7721), .ZN(n7722) );
  NAND2_X1 U9352 ( .A1(n7723), .A2(n7722), .ZN(n9158) );
  AND2_X1 U9353 ( .A1(n9158), .A2(n7801), .ZN(n7724) );
  AOI21_X1 U9354 ( .B1(n9334), .B2(n4256), .A(n7724), .ZN(n7728) );
  NAND2_X1 U9355 ( .A1(n9334), .A2(n7793), .ZN(n7726) );
  NAND2_X1 U9356 ( .A1(n9158), .A2(n4256), .ZN(n7725) );
  NAND2_X1 U9357 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  XNOR2_X1 U9358 ( .A(n7727), .B(n7799), .ZN(n8881) );
  NAND2_X1 U9359 ( .A1(n8878), .A2(n8881), .ZN(n7729) );
  NAND2_X1 U9360 ( .A1(n7729), .A2(n8879), .ZN(n7749) );
  INV_X1 U9361 ( .A(n7749), .ZN(n7746) );
  NAND2_X1 U9362 ( .A1(n7730), .A2(n6643), .ZN(n7733) );
  OR2_X1 U9363 ( .A1(n7957), .A2(n7731), .ZN(n7732) );
  NAND2_X1 U9364 ( .A1(n9328), .A2(n7808), .ZN(n7744) );
  INV_X1 U9365 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U9366 ( .A1(n7735), .A2(n7734), .ZN(n7736) );
  NAND2_X1 U9367 ( .A1(n7737), .A2(n7736), .ZN(n9154) );
  OR2_X1 U9368 ( .A1(n9154), .A2(n4272), .ZN(n7742) );
  INV_X1 U9369 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U9370 ( .A1(n7813), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U9371 ( .A1(n7853), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7738) );
  OAI211_X1 U9372 ( .C1(n7852), .C2(n10015), .A(n7739), .B(n7738), .ZN(n7740)
         );
  INV_X1 U9373 ( .A(n7740), .ZN(n7741) );
  NAND2_X1 U9374 ( .A1(n7742), .A2(n7741), .ZN(n9146) );
  NAND2_X1 U9375 ( .A1(n9146), .A2(n4256), .ZN(n7743) );
  NAND2_X1 U9376 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  XNOR2_X1 U9377 ( .A(n7745), .B(n7822), .ZN(n7747) );
  INV_X1 U9378 ( .A(n9328), .ZN(n9157) );
  INV_X1 U9379 ( .A(n9146), .ZN(n9173) );
  INV_X1 U9380 ( .A(n7801), .ZN(n7826) );
  OAI22_X1 U9381 ( .A1(n9157), .A2(n7798), .B1(n9173), .B2(n7826), .ZN(n8808)
         );
  AND2_X2 U9382 ( .A1(n7749), .A2(n7748), .ZN(n8807) );
  XOR2_X1 U9383 ( .A(n7751), .B(n7750), .Z(n8865) );
  OR2_X1 U9384 ( .A1(n7957), .A2(n7753), .ZN(n7754) );
  NAND2_X1 U9385 ( .A1(n9319), .A2(n7808), .ZN(n7766) );
  INV_X1 U9386 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9387 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  NAND2_X1 U9388 ( .A1(n7775), .A2(n7758), .ZN(n9130) );
  INV_X1 U9389 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U9390 ( .A1(n7853), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U9391 ( .A1(n7813), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7759) );
  OAI211_X1 U9392 ( .C1(n7852), .C2(n7761), .A(n7760), .B(n7759), .ZN(n7762)
         );
  INV_X1 U9393 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U9394 ( .A1(n9147), .A2(n4256), .ZN(n7765) );
  NAND2_X1 U9395 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  XNOR2_X1 U9396 ( .A(n7767), .B(n7799), .ZN(n7768) );
  AOI22_X1 U9397 ( .A1(n9319), .A2(n7824), .B1(n7801), .B2(n9147), .ZN(n7769)
         );
  XNOR2_X1 U9398 ( .A(n7768), .B(n7769), .ZN(n8840) );
  INV_X1 U9399 ( .A(n7768), .ZN(n7770) );
  OR2_X1 U9400 ( .A1(n7957), .A2(n7772), .ZN(n7773) );
  NAND2_X1 U9401 ( .A1(n9314), .A2(n7808), .ZN(n7784) );
  NAND2_X1 U9402 ( .A1(n7775), .A2(n8903), .ZN(n7776) );
  NAND2_X1 U9403 ( .A1(n9117), .A2(n7797), .ZN(n7782) );
  INV_X1 U9404 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U9405 ( .A1(n7853), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U9406 ( .A1(n7813), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7777) );
  OAI211_X1 U9407 ( .C1(n7852), .C2(n7779), .A(n7778), .B(n7777), .ZN(n7780)
         );
  INV_X1 U9408 ( .A(n7780), .ZN(n7781) );
  NAND2_X1 U9409 ( .A1(n8927), .A2(n4256), .ZN(n7783) );
  NAND2_X1 U9410 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  XNOR2_X1 U9411 ( .A(n7785), .B(n7799), .ZN(n7786) );
  AOI22_X1 U9412 ( .A1(n9314), .A2(n7824), .B1(n7801), .B2(n8927), .ZN(n7787)
         );
  XNOR2_X1 U9413 ( .A(n7786), .B(n7787), .ZN(n8900) );
  INV_X1 U9414 ( .A(n7786), .ZN(n7788) );
  NAND2_X1 U9415 ( .A1(n8899), .A2(n4349), .ZN(n8789) );
  NAND2_X1 U9416 ( .A1(n7789), .A2(n6643), .ZN(n7792) );
  OR2_X1 U9417 ( .A1(n7957), .A2(n7790), .ZN(n7791) );
  XNOR2_X1 U9418 ( .A(n7811), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9102) );
  INV_X1 U9419 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U9420 ( .A1(n7813), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U9421 ( .A1(n7853), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7794) );
  OAI211_X1 U9422 ( .C1(n7852), .C2(n9953), .A(n7795), .B(n7794), .ZN(n7796)
         );
  AOI21_X1 U9423 ( .B1(n9102), .B2(n7797), .A(n7796), .ZN(n9113) );
  OAI22_X1 U9424 ( .A1(n9034), .A2(n6488), .B1(n9113), .B2(n7798), .ZN(n7800)
         );
  XNOR2_X1 U9425 ( .A(n7800), .B(n7799), .ZN(n8787) );
  INV_X1 U9426 ( .A(n8787), .ZN(n7803) );
  AND2_X1 U9427 ( .A1(n8926), .A2(n7801), .ZN(n7802) );
  AOI21_X1 U9428 ( .B1(n9310), .B2(n7824), .A(n7802), .ZN(n8786) );
  INV_X1 U9429 ( .A(n8786), .ZN(n7830) );
  NAND2_X1 U9430 ( .A1(n7803), .A2(n8786), .ZN(n7804) );
  NAND2_X1 U9431 ( .A1(n8789), .A2(n7804), .ZN(n7844) );
  NAND2_X1 U9432 ( .A1(n7805), .A2(n6643), .ZN(n7807) );
  INV_X1 U9433 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8122) );
  OR2_X1 U9434 ( .A1(n7957), .A2(n8122), .ZN(n7806) );
  NAND2_X1 U9435 ( .A1(n9306), .A2(n7808), .ZN(n7821) );
  INV_X1 U9436 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7810) );
  INV_X1 U9437 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7809) );
  OAI21_X1 U9438 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7812) );
  NAND2_X1 U9439 ( .A1(n7812), .A2(n9074), .ZN(n7834) );
  OR2_X1 U9440 ( .A1(n7834), .A2(n4272), .ZN(n7819) );
  INV_X1 U9441 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U9442 ( .A1(n7813), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U9443 ( .A1(n7853), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7814) );
  OAI211_X1 U9444 ( .C1(n7852), .C2(n7816), .A(n7815), .B(n7814), .ZN(n7817)
         );
  INV_X1 U9445 ( .A(n7817), .ZN(n7818) );
  NAND2_X1 U9446 ( .A1(n9038), .A2(n4256), .ZN(n7820) );
  NAND2_X1 U9447 ( .A1(n7821), .A2(n7820), .ZN(n7823) );
  XNOR2_X1 U9448 ( .A(n7823), .B(n7822), .ZN(n7828) );
  NAND2_X1 U9449 ( .A1(n9306), .A2(n4256), .ZN(n7825) );
  OAI21_X1 U9450 ( .B1(n9100), .B2(n7826), .A(n7825), .ZN(n7827) );
  XNOR2_X1 U9451 ( .A(n7828), .B(n7827), .ZN(n7838) );
  INV_X1 U9452 ( .A(n7838), .ZN(n7829) );
  NAND2_X1 U9453 ( .A1(n7829), .A2(n8898), .ZN(n7843) );
  NAND2_X1 U9454 ( .A1(n8787), .A2(n7830), .ZN(n7837) );
  INV_X1 U9455 ( .A(n7837), .ZN(n7831) );
  NOR2_X1 U9456 ( .A1(n7831), .A2(n8923), .ZN(n7832) );
  AND2_X1 U9457 ( .A1(n7838), .A2(n7832), .ZN(n7833) );
  NAND2_X1 U9458 ( .A1(n7844), .A2(n7833), .ZN(n7842) );
  NAND2_X1 U9459 ( .A1(n8926), .A2(n8901), .ZN(n7836) );
  INV_X1 U9460 ( .A(n7834), .ZN(n9089) );
  AOI22_X1 U9461 ( .A1(n9089), .A2(n8907), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7835) );
  OAI211_X1 U9462 ( .C1(n9085), .C2(n8904), .A(n7836), .B(n7835), .ZN(n7840)
         );
  NOR3_X1 U9463 ( .A1(n7838), .A2(n8923), .A3(n7837), .ZN(n7839) );
  AOI211_X1 U9464 ( .C1(n9306), .C2(n8894), .A(n7840), .B(n7839), .ZN(n7841)
         );
  OAI211_X1 U9465 ( .C1(n7844), .C2(n7843), .A(n7842), .B(n7841), .ZN(P1_U3218) );
  NAND2_X1 U9466 ( .A1(n7845), .A2(n6643), .ZN(n7847) );
  INV_X1 U9467 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9403) );
  OR2_X1 U9468 ( .A1(n7957), .A2(n9403), .ZN(n7846) );
  NAND2_X1 U9469 ( .A1(n7847), .A2(n7846), .ZN(n7967) );
  INV_X1 U9470 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U9471 ( .A1(n7853), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7850) );
  INV_X1 U9472 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9921) );
  OR2_X1 U9473 ( .A1(n7848), .A2(n9921), .ZN(n7849) );
  OAI211_X1 U9474 ( .C1(n7852), .C2(n7851), .A(n7850), .B(n7849), .ZN(n8925)
         );
  INV_X1 U9475 ( .A(n8925), .ZN(n9070) );
  INV_X1 U9476 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U9477 ( .A1(n7853), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7856) );
  INV_X1 U9478 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7854) );
  OR2_X1 U9479 ( .A1(n7848), .A2(n7854), .ZN(n7855) );
  OAI211_X1 U9480 ( .C1(n7852), .C2(n7857), .A(n7856), .B(n7855), .ZN(n9002)
         );
  NAND2_X1 U9481 ( .A1(n8107), .A2(n9002), .ZN(n7861) );
  NAND2_X1 U9482 ( .A1(n8772), .A2(n6643), .ZN(n7860) );
  OR2_X1 U9483 ( .A1(n7957), .A2(n6039), .ZN(n7859) );
  NAND2_X1 U9484 ( .A1(n9002), .A2(n8925), .ZN(n7862) );
  NAND2_X1 U9485 ( .A1(n7967), .A2(n7862), .ZN(n8060) );
  OAI211_X1 U9486 ( .C1(n9085), .C2(n4448), .A(n8064), .B(n8060), .ZN(n7863)
         );
  INV_X1 U9487 ( .A(n7863), .ZN(n7966) );
  OR2_X2 U9488 ( .A1(n9319), .A2(n9112), .ZN(n9062) );
  OR2_X1 U9489 ( .A1(n9323), .A2(n9127), .ZN(n7865) );
  OR2_X1 U9490 ( .A1(n9328), .A2(n9173), .ZN(n9059) );
  NAND2_X1 U9491 ( .A1(n7865), .A2(n9059), .ZN(n8011) );
  NAND2_X1 U9492 ( .A1(n9323), .A2(n9127), .ZN(n9061) );
  NAND2_X1 U9493 ( .A1(n8011), .A2(n9061), .ZN(n7864) );
  NAND2_X1 U9494 ( .A1(n9062), .A2(n7864), .ZN(n7867) );
  NAND2_X1 U9495 ( .A1(n9328), .A2(n9173), .ZN(n7969) );
  NAND2_X1 U9496 ( .A1(n9061), .A2(n7969), .ZN(n7934) );
  NAND2_X1 U9497 ( .A1(n7934), .A2(n7865), .ZN(n7866) );
  NAND2_X1 U9498 ( .A1(n7968), .A2(n7866), .ZN(n8051) );
  MUX2_X1 U9499 ( .A(n7867), .B(n8051), .S(n4448), .Z(n7868) );
  INV_X1 U9500 ( .A(n7868), .ZN(n7936) );
  INV_X1 U9501 ( .A(n9017), .ZN(n9254) );
  INV_X1 U9502 ( .A(n9015), .ZN(n9263) );
  OR2_X1 U9503 ( .A1(n9359), .A2(n9263), .ZN(n9050) );
  NAND2_X1 U9504 ( .A1(n7996), .A2(n9050), .ZN(n8009) );
  NAND2_X1 U9505 ( .A1(n9354), .A2(n9254), .ZN(n9051) );
  AND2_X1 U9506 ( .A1(n9359), .A2(n9263), .ZN(n9049) );
  INV_X1 U9507 ( .A(n9049), .ZN(n8023) );
  NAND2_X1 U9508 ( .A1(n9051), .A2(n8023), .ZN(n7869) );
  MUX2_X1 U9509 ( .A(n8009), .B(n7869), .S(n4448), .Z(n7870) );
  AND2_X1 U9510 ( .A1(n7872), .A2(n8020), .ZN(n7873) );
  OAI21_X1 U9511 ( .B1(n7875), .B2(n7964), .A(n7874), .ZN(n7876) );
  AND2_X1 U9512 ( .A1(n8085), .A2(n7877), .ZN(n8022) );
  NAND2_X1 U9513 ( .A1(n7891), .A2(n7889), .ZN(n8028) );
  AOI21_X1 U9514 ( .B1(n7890), .B2(n8022), .A(n8028), .ZN(n7882) );
  NAND2_X1 U9515 ( .A1(n7878), .A2(n8038), .ZN(n7881) );
  INV_X1 U9516 ( .A(n7879), .ZN(n7880) );
  OAI21_X1 U9517 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7884) );
  MUX2_X1 U9518 ( .A(n7884), .B(n7883), .S(n7964), .Z(n7887) );
  INV_X1 U9519 ( .A(n7902), .ZN(n7885) );
  NOR2_X1 U9520 ( .A1(n7885), .A2(n7976), .ZN(n7886) );
  NAND2_X1 U9521 ( .A1(n7887), .A2(n7886), .ZN(n7909) );
  AND2_X1 U9522 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  AOI21_X1 U9523 ( .B1(n7894), .B2(n7893), .A(n8037), .ZN(n7897) );
  NAND2_X1 U9524 ( .A1(n7903), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U9525 ( .A1(n10034), .A2(n9286), .ZN(n8024) );
  NAND2_X1 U9526 ( .A1(n9442), .A2(n7900), .ZN(n9043) );
  NAND2_X1 U9527 ( .A1(n8024), .A2(n9043), .ZN(n7910) );
  NAND2_X1 U9528 ( .A1(n7902), .A2(n7898), .ZN(n8027) );
  AND2_X1 U9529 ( .A1(n8027), .A2(n7903), .ZN(n7899) );
  NOR2_X1 U9530 ( .A1(n7910), .A2(n7899), .ZN(n7906) );
  OR2_X1 U9531 ( .A1(n9442), .A2(n7900), .ZN(n7975) );
  NAND2_X1 U9532 ( .A1(n9044), .A2(n7975), .ZN(n8036) );
  NAND2_X1 U9533 ( .A1(n7902), .A2(n7901), .ZN(n7904) );
  AND2_X1 U9534 ( .A1(n7904), .A2(n7903), .ZN(n9040) );
  INV_X1 U9535 ( .A(n9040), .ZN(n8040) );
  NOR2_X1 U9536 ( .A1(n8036), .A2(n8040), .ZN(n7905) );
  MUX2_X1 U9537 ( .A(n7906), .B(n7905), .S(n7964), .Z(n7907) );
  OAI21_X1 U9538 ( .B1(n7909), .B2(n7908), .A(n7907), .ZN(n7914) );
  INV_X1 U9539 ( .A(n9046), .ZN(n8025) );
  OR2_X1 U9540 ( .A1(n9371), .A2(n9262), .ZN(n9257) );
  NAND2_X1 U9541 ( .A1(n7910), .A2(n9044), .ZN(n7912) );
  NAND2_X1 U9542 ( .A1(n8036), .A2(n8024), .ZN(n7911) );
  MUX2_X1 U9543 ( .A(n7912), .B(n7911), .S(n4448), .Z(n7913) );
  NAND3_X1 U9544 ( .A1(n7914), .A2(n9284), .A3(n7913), .ZN(n7916) );
  INV_X1 U9545 ( .A(n9014), .ZN(n9288) );
  OR2_X1 U9546 ( .A1(n9365), .A2(n9288), .ZN(n8045) );
  NAND2_X1 U9547 ( .A1(n9365), .A2(n9288), .ZN(n9047) );
  MUX2_X1 U9548 ( .A(n9257), .B(n8025), .S(n4448), .Z(n7915) );
  MUX2_X1 U9549 ( .A(n8045), .B(n9047), .S(n7964), .Z(n7917) );
  INV_X1 U9550 ( .A(n9018), .ZN(n9241) );
  OR2_X1 U9551 ( .A1(n9349), .A2(n9241), .ZN(n7974) );
  INV_X1 U9552 ( .A(n9020), .ZN(n9219) );
  NAND2_X1 U9553 ( .A1(n9344), .A2(n9219), .ZN(n7973) );
  NAND2_X1 U9554 ( .A1(n9349), .A2(n9241), .ZN(n9199) );
  NAND2_X1 U9555 ( .A1(n7973), .A2(n9199), .ZN(n9054) );
  INV_X1 U9556 ( .A(n9054), .ZN(n7919) );
  NAND2_X1 U9557 ( .A1(n7920), .A2(n7919), .ZN(n7924) );
  OR2_X1 U9558 ( .A1(n9344), .A2(n9219), .ZN(n9053) );
  AND2_X1 U9559 ( .A1(n9053), .A2(n7974), .ZN(n8006) );
  AND2_X1 U9560 ( .A1(n9199), .A2(n9051), .ZN(n8010) );
  NAND2_X1 U9561 ( .A1(n7921), .A2(n8010), .ZN(n7922) );
  NAND2_X1 U9562 ( .A1(n8006), .A2(n7922), .ZN(n7923) );
  INV_X1 U9563 ( .A(n9022), .ZN(n9204) );
  AND2_X1 U9564 ( .A1(n7972), .A2(n9053), .ZN(n7925) );
  NAND2_X1 U9565 ( .A1(n9339), .A2(n9204), .ZN(n7971) );
  INV_X1 U9566 ( .A(n7971), .ZN(n9056) );
  AOI21_X1 U9567 ( .B1(n7930), .B2(n7925), .A(n9056), .ZN(n7926) );
  NOR2_X1 U9568 ( .A1(n9334), .A2(n9189), .ZN(n9058) );
  NAND2_X1 U9569 ( .A1(n9334), .A2(n9189), .ZN(n9057) );
  OAI21_X1 U9570 ( .B1(n7926), .B2(n9058), .A(n9057), .ZN(n7933) );
  INV_X1 U9571 ( .A(n7972), .ZN(n8007) );
  INV_X1 U9572 ( .A(n7973), .ZN(n7927) );
  NAND2_X1 U9573 ( .A1(n7972), .A2(n7927), .ZN(n7928) );
  AND2_X1 U9574 ( .A1(n7928), .A2(n7971), .ZN(n7929) );
  AND2_X1 U9575 ( .A1(n9057), .A2(n7929), .ZN(n8049) );
  OAI21_X1 U9576 ( .B1(n7930), .B2(n8007), .A(n8049), .ZN(n7931) );
  INV_X1 U9577 ( .A(n9058), .ZN(n8012) );
  NAND2_X1 U9578 ( .A1(n7931), .A2(n8012), .ZN(n7932) );
  NOR2_X1 U9579 ( .A1(n8011), .A2(n7934), .ZN(n7935) );
  INV_X1 U9580 ( .A(n7944), .ZN(n7937) );
  NAND2_X1 U9581 ( .A1(n9096), .A2(n7937), .ZN(n7942) );
  INV_X1 U9582 ( .A(n7968), .ZN(n9063) );
  OAI21_X1 U9583 ( .B1(n9128), .B2(n9063), .A(n9065), .ZN(n7940) );
  NAND2_X1 U9584 ( .A1(n9314), .A2(n9062), .ZN(n7938) );
  NAND2_X1 U9585 ( .A1(n8053), .A2(n7938), .ZN(n7939) );
  MUX2_X1 U9586 ( .A(n7940), .B(n7939), .S(n4448), .Z(n7941) );
  AND2_X1 U9587 ( .A1(n7942), .A2(n7941), .ZN(n7951) );
  NAND2_X1 U9588 ( .A1(n7944), .A2(n7968), .ZN(n7943) );
  AOI21_X1 U9589 ( .B1(n7943), .B2(n9128), .A(n9314), .ZN(n7947) );
  AOI21_X1 U9590 ( .B1(n7945), .B2(n9120), .A(n8927), .ZN(n7946) );
  MUX2_X1 U9591 ( .A(n7947), .B(n7946), .S(n4448), .Z(n7950) );
  NAND2_X1 U9592 ( .A1(n9306), .A2(n9100), .ZN(n8055) );
  MUX2_X1 U9593 ( .A(n9065), .B(n8053), .S(n7964), .Z(n7948) );
  AND2_X1 U9594 ( .A1(n9082), .A2(n7948), .ZN(n7949) );
  OAI21_X1 U9595 ( .B1(n7951), .B2(n7950), .A(n7949), .ZN(n7953) );
  MUX2_X1 U9596 ( .A(n8055), .B(n9066), .S(n7964), .Z(n7952) );
  INV_X1 U9597 ( .A(n7961), .ZN(n7954) );
  NAND2_X1 U9598 ( .A1(n7954), .A2(n9085), .ZN(n7960) );
  NAND2_X1 U9599 ( .A1(n7955), .A2(n6643), .ZN(n7959) );
  OR2_X1 U9600 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  MUX2_X1 U9601 ( .A(n7960), .B(n7964), .S(n9301), .Z(n7965) );
  INV_X1 U9602 ( .A(n9002), .ZN(n7962) );
  AND2_X1 U9603 ( .A1(n7963), .A2(n7962), .ZN(n8108) );
  NOR4_X1 U9604 ( .A1(n4253), .A2(n8104), .A3(n6075), .A4(n8062), .ZN(n8070)
         );
  NOR2_X1 U9605 ( .A1(n9297), .A2(n8925), .ZN(n8105) );
  INV_X1 U9606 ( .A(n8107), .ZN(n8002) );
  NAND2_X1 U9607 ( .A1(n9301), .A2(n9085), .ZN(n8101) );
  INV_X1 U9608 ( .A(n9039), .ZN(n9068) );
  XNOR2_X1 U9609 ( .A(n9323), .B(n9164), .ZN(n9144) );
  INV_X1 U9610 ( .A(n9144), .ZN(n9135) );
  NAND2_X1 U9611 ( .A1(n9059), .A2(n7969), .ZN(n9161) );
  INV_X1 U9612 ( .A(n9057), .ZN(n7970) );
  OR2_X1 U9613 ( .A1(n9058), .A2(n7970), .ZN(n9169) );
  INV_X1 U9614 ( .A(n9169), .ZN(n9170) );
  NAND2_X1 U9615 ( .A1(n9053), .A2(n7973), .ZN(n9202) );
  NAND2_X1 U9616 ( .A1(n7974), .A2(n9199), .ZN(n9216) );
  NAND2_X1 U9617 ( .A1(n7975), .A2(n9043), .ZN(n9434) );
  INV_X1 U9618 ( .A(n9434), .ZN(n7993) );
  INV_X1 U9619 ( .A(n7976), .ZN(n7991) );
  AND2_X1 U9620 ( .A1(n7978), .A2(n7977), .ZN(n7981) );
  NAND4_X1 U9621 ( .A1(n8032), .A2(n7981), .A3(n7980), .A4(n7979), .ZN(n7983)
         );
  NOR2_X1 U9622 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND4_X1 U9623 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n8083), .ZN(n7987)
         );
  NOR3_X1 U9624 ( .A1(n7989), .A2(n7988), .A3(n7987), .ZN(n7990) );
  NAND4_X1 U9625 ( .A1(n7993), .A2(n7992), .A3(n7991), .A4(n7990), .ZN(n7994)
         );
  NOR2_X1 U9626 ( .A1(n7994), .A2(n9448), .ZN(n7995) );
  NAND4_X1 U9627 ( .A1(n9252), .A2(n9264), .A3(n9284), .A4(n7995), .ZN(n7997)
         );
  NOR4_X1 U9628 ( .A1(n9202), .A2(n9216), .A3(n7997), .A4(n9238), .ZN(n7998)
         );
  NAND4_X1 U9629 ( .A1(n4806), .A2(n9170), .A3(n9055), .A4(n7998), .ZN(n7999)
         );
  NOR3_X1 U9630 ( .A1(n9124), .A2(n9135), .A3(n7999), .ZN(n8000) );
  NAND4_X1 U9631 ( .A1(n9082), .A2(n9096), .A3(n8000), .A4(n9109), .ZN(n8001)
         );
  NOR4_X1 U9632 ( .A1(n8105), .A2(n8002), .A3(n9068), .A4(n8001), .ZN(n8003)
         );
  NAND2_X1 U9633 ( .A1(n8003), .A2(n4432), .ZN(n8004) );
  OAI21_X1 U9634 ( .B1(n8004), .B2(n8104), .A(n8062), .ZN(n8067) );
  INV_X1 U9635 ( .A(n8067), .ZN(n8066) );
  INV_X1 U9636 ( .A(n9065), .ZN(n8056) );
  INV_X1 U9637 ( .A(n9062), .ZN(n8005) );
  NOR2_X1 U9638 ( .A1(n9314), .A2(n9128), .ZN(n9064) );
  NOR3_X1 U9639 ( .A1(n8056), .A2(n8005), .A3(n9064), .ZN(n8100) );
  INV_X1 U9640 ( .A(n8006), .ZN(n8008) );
  AOI211_X1 U9641 ( .C1(n8010), .C2(n8009), .A(n8008), .B(n8007), .ZN(n8015)
         );
  INV_X1 U9642 ( .A(n8049), .ZN(n8014) );
  INV_X1 U9643 ( .A(n8011), .ZN(n8013) );
  OAI211_X1 U9644 ( .C1(n8015), .C2(n8014), .A(n8013), .B(n8012), .ZN(n8092)
         );
  INV_X1 U9645 ( .A(n8032), .ZN(n8016) );
  AOI21_X1 U9646 ( .B1(n8017), .B2(n8081), .A(n8016), .ZN(n8021) );
  INV_X1 U9647 ( .A(n8018), .ZN(n8019) );
  AOI21_X1 U9648 ( .B1(n8021), .B2(n8020), .A(n8019), .ZN(n8035) );
  INV_X1 U9649 ( .A(n8022), .ZN(n8034) );
  NAND3_X1 U9650 ( .A1(n9051), .A2(n8023), .A3(n9047), .ZN(n8046) );
  NAND2_X1 U9651 ( .A1(n8025), .A2(n8024), .ZN(n8042) );
  OR2_X1 U9652 ( .A1(n8027), .A2(n8026), .ZN(n9041) );
  INV_X1 U9653 ( .A(n8028), .ZN(n8029) );
  NAND2_X1 U9654 ( .A1(n9043), .A2(n8029), .ZN(n8030) );
  NOR4_X1 U9655 ( .A1(n8046), .A2(n8042), .A3(n9041), .A4(n8030), .ZN(n8091)
         );
  AND2_X1 U9656 ( .A1(n8032), .A2(n8031), .ZN(n8079) );
  NAND4_X1 U9657 ( .A1(n9625), .A2(n8079), .A3(n8085), .A4(n8084), .ZN(n8033)
         );
  OAI211_X1 U9658 ( .C1(n8035), .C2(n8034), .A(n8091), .B(n8033), .ZN(n8050)
         );
  INV_X1 U9659 ( .A(n8036), .ZN(n8044) );
  INV_X1 U9660 ( .A(n8037), .ZN(n8039) );
  AOI21_X1 U9661 ( .B1(n8039), .B2(n8038), .A(n9041), .ZN(n8041) );
  OAI21_X1 U9662 ( .B1(n8041), .B2(n8040), .A(n9043), .ZN(n8043) );
  AOI21_X1 U9663 ( .B1(n8044), .B2(n8043), .A(n8042), .ZN(n8048) );
  NAND2_X1 U9664 ( .A1(n8045), .A2(n9257), .ZN(n9048) );
  INV_X1 U9665 ( .A(n8046), .ZN(n8047) );
  OAI21_X1 U9666 ( .B1(n8048), .B2(n9048), .A(n8047), .ZN(n8088) );
  NAND2_X1 U9667 ( .A1(n8049), .A2(n9199), .ZN(n8095) );
  AOI21_X1 U9668 ( .B1(n8050), .B2(n8088), .A(n8095), .ZN(n8052) );
  INV_X1 U9669 ( .A(n8051), .ZN(n8096) );
  OAI21_X1 U9670 ( .B1(n8092), .B2(n8052), .A(n8096), .ZN(n8058) );
  INV_X1 U9671 ( .A(n8053), .ZN(n8054) );
  AOI21_X1 U9672 ( .B1(n9128), .B2(n9314), .A(n8054), .ZN(n8057) );
  OAI21_X1 U9673 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8098) );
  AOI21_X1 U9674 ( .B1(n8100), .B2(n8058), .A(n8098), .ZN(n8061) );
  NAND2_X1 U9675 ( .A1(n8059), .A2(n9066), .ZN(n8102) );
  OAI211_X1 U9676 ( .C1(n8061), .C2(n8102), .A(n8101), .B(n8060), .ZN(n8063)
         );
  AOI211_X1 U9677 ( .C1(n8064), .C2(n8063), .A(n8062), .B(n8104), .ZN(n8065)
         );
  NOR2_X1 U9678 ( .A1(n8066), .A2(n8065), .ZN(n8069) );
  NAND2_X1 U9679 ( .A1(n8937), .A2(n8071), .ZN(n8072) );
  OAI211_X1 U9680 ( .C1(n8073), .C2(n6163), .A(n6103), .B(n8072), .ZN(n8075)
         );
  NAND2_X1 U9681 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  OAI22_X1 U9682 ( .A1(n8078), .A2(n8077), .B1(n8076), .B2(n9651), .ZN(n8082)
         );
  INV_X1 U9683 ( .A(n8079), .ZN(n8080) );
  AOI21_X1 U9684 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n8087) );
  INV_X1 U9685 ( .A(n8083), .ZN(n8086) );
  OAI211_X1 U9686 ( .C1(n8087), .C2(n8086), .A(n8085), .B(n8084), .ZN(n8090)
         );
  INV_X1 U9687 ( .A(n8088), .ZN(n8089) );
  AOI21_X1 U9688 ( .B1(n8091), .B2(n8090), .A(n8089), .ZN(n8094) );
  INV_X1 U9689 ( .A(n8092), .ZN(n8093) );
  OAI21_X1 U9690 ( .B1(n8095), .B2(n8094), .A(n8093), .ZN(n8097) );
  NAND2_X1 U9691 ( .A1(n8097), .A2(n8096), .ZN(n8099) );
  AOI21_X1 U9692 ( .B1(n8100), .B2(n8099), .A(n8098), .ZN(n8103) );
  OAI21_X1 U9693 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8106) );
  AOI211_X1 U9694 ( .C1(n8107), .C2(n8106), .A(n8105), .B(n8104), .ZN(n8109)
         );
  NOR2_X1 U9695 ( .A1(n8109), .A2(n8108), .ZN(n8115) );
  INV_X1 U9696 ( .A(n8110), .ZN(n8114) );
  NAND3_X1 U9697 ( .A1(n8115), .A2(n9193), .A3(n8111), .ZN(n8113) );
  INV_X1 U9698 ( .A(n8117), .ZN(n8112) );
  OAI211_X1 U9699 ( .C1(n8115), .C2(n8114), .A(n8113), .B(n8112), .ZN(n8120)
         );
  NOR3_X1 U9700 ( .A1(n8116), .A2(n8123), .A3(n4278), .ZN(n8119) );
  OAI21_X1 U9701 ( .B1(n6075), .B2(n8117), .A(P1_B_REG_SCAN_IN), .ZN(n8118) );
  OAI222_X1 U9702 ( .A1(n9402), .A2(n8124), .B1(P1_U3084), .B2(n8123), .C1(
        n8122), .C2(n8121), .ZN(P1_U3325) );
  AOI22_X1 U9703 ( .A1(n8256), .A2(n5095), .B1(n5866), .B2(n8125), .ZN(n8127)
         );
  NOR2_X1 U9704 ( .A1(n8127), .A2(n8126), .ZN(n8135) );
  INV_X1 U9705 ( .A(n8128), .ZN(n8129) );
  OAI22_X1 U9706 ( .A1(n8264), .A2(n8129), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8309), .ZN(n8133) );
  OAI22_X1 U9707 ( .A1(n8131), .A2(n8270), .B1(n8251), .B2(n8130), .ZN(n8132)
         );
  AOI211_X1 U9708 ( .C1(n8135), .C2(n8134), .A(n8133), .B(n8132), .ZN(n8136)
         );
  OAI21_X1 U9709 ( .B1(n8137), .B2(n8244), .A(n8136), .ZN(P2_U3229) );
  NAND3_X1 U9710 ( .A1(n8139), .A2(n8256), .A3(n8274), .ZN(n8140) );
  NAND2_X1 U9711 ( .A1(n8143), .A2(n8142), .ZN(n8148) );
  NOR2_X1 U9712 ( .A1(n8425), .A2(n8251), .ZN(n8146) );
  NOR2_X1 U9713 ( .A1(n8184), .A2(n8621), .ZN(n8144) );
  AOI21_X1 U9714 ( .B1(n8272), .B2(n9740), .A(n8144), .ZN(n8418) );
  NOR2_X1 U9715 ( .A1(n8418), .A2(n8264), .ZN(n8145) );
  AOI211_X1 U9716 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n8146), 
        .B(n8145), .ZN(n8147) );
  OAI211_X1 U9717 ( .C1(n8730), .C2(n8270), .A(n8148), .B(n8147), .ZN(P2_U3216) );
  INV_X1 U9718 ( .A(n8149), .ZN(n8150) );
  NOR2_X1 U9719 ( .A1(n8151), .A2(n8150), .ZN(n8153) );
  NAND3_X1 U9720 ( .A1(n8153), .A2(n5866), .A3(n8152), .ZN(n8160) );
  INV_X1 U9721 ( .A(n8153), .ZN(n8154) );
  NAND3_X1 U9722 ( .A1(n8154), .A2(n8256), .A3(n8505), .ZN(n8159) );
  OAI22_X1 U9723 ( .A1(n8251), .A2(n8483), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8155), .ZN(n8157) );
  OAI22_X1 U9724 ( .A1(n8213), .A2(n8234), .B1(n8233), .B2(n8526), .ZN(n8156)
         );
  AOI211_X1 U9725 ( .C1(n8665), .C2(n8238), .A(n8157), .B(n8156), .ZN(n8158)
         );
  NAND3_X1 U9726 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(P2_U3218) );
  AND2_X1 U9727 ( .A1(n8256), .A2(n8539), .ZN(n8161) );
  AOI22_X1 U9728 ( .A1(n8163), .A2(n5866), .B1(n8162), .B2(n8161), .ZN(n8167)
         );
  NAND3_X1 U9729 ( .A1(n4715), .A2(n5866), .A3(n8164), .ZN(n8166) );
  MUX2_X1 U9730 ( .A(n8167), .B(n8166), .S(n8165), .Z(n8172) );
  INV_X1 U9731 ( .A(n8168), .ZN(n8571) );
  AOI22_X1 U9732 ( .A1(n8266), .A2(n8571), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8171) );
  AOI22_X1 U9733 ( .A1(n8199), .A2(n8277), .B1(n8198), .B2(n8276), .ZN(n8170)
         );
  NAND2_X1 U9734 ( .A1(n8688), .A2(n8238), .ZN(n8169) );
  NAND4_X1 U9735 ( .A1(n8172), .A2(n8171), .A3(n8170), .A4(n8169), .ZN(
        P2_U3221) );
  XNOR2_X1 U9736 ( .A(n8174), .B(n8173), .ZN(n8179) );
  OAI22_X1 U9737 ( .A1(n8251), .A2(n8528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8175), .ZN(n8177) );
  OAI22_X1 U9738 ( .A1(n8526), .A2(n8234), .B1(n8233), .B2(n8567), .ZN(n8176)
         );
  AOI211_X1 U9739 ( .C1(n8676), .C2(n8238), .A(n8177), .B(n8176), .ZN(n8178)
         );
  OAI21_X1 U9740 ( .B1(n8179), .B2(n8244), .A(n8178), .ZN(P2_U3225) );
  XNOR2_X1 U9741 ( .A(n8182), .B(n8181), .ZN(n8183) );
  XNOR2_X1 U9742 ( .A(n8180), .B(n8183), .ZN(n8190) );
  NOR2_X1 U9743 ( .A1(n8251), .A2(n8457), .ZN(n8188) );
  OR2_X1 U9744 ( .A1(n8184), .A2(n8619), .ZN(n8186) );
  OR2_X1 U9745 ( .A1(n8213), .A2(n8621), .ZN(n8185) );
  AND2_X1 U9746 ( .A1(n8186), .A2(n8185), .ZN(n8449) );
  OAI22_X1 U9747 ( .A1(n8449), .A2(n8264), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9997), .ZN(n8187) );
  AOI211_X1 U9748 ( .C1(n8456), .C2(n8238), .A(n8188), .B(n8187), .ZN(n8189)
         );
  OAI21_X1 U9749 ( .B1(n8190), .B2(n8244), .A(n8189), .ZN(P2_U3227) );
  XNOR2_X1 U9750 ( .A(n8192), .B(n8191), .ZN(n8258) );
  AOI22_X1 U9751 ( .A1(n8258), .A2(n8257), .B1(n8193), .B2(n8192), .ZN(n8197)
         );
  XNOR2_X1 U9752 ( .A(n8195), .B(n8194), .ZN(n8196) );
  XNOR2_X1 U9753 ( .A(n8197), .B(n8196), .ZN(n8204) );
  AOI22_X1 U9754 ( .A1(n8199), .A2(n8279), .B1(n8198), .B2(n5315), .ZN(n8201)
         );
  OAI211_X1 U9755 ( .C1(n8630), .C2(n8251), .A(n8201), .B(n8200), .ZN(n8202)
         );
  AOI21_X1 U9756 ( .B1(n8629), .B2(n8238), .A(n8202), .ZN(n8203) );
  OAI21_X1 U9757 ( .B1(n8204), .B2(n8244), .A(n8203), .ZN(P2_U3228) );
  OAI211_X1 U9758 ( .C1(n8206), .C2(n8205), .A(n8246), .B(n5866), .ZN(n8210)
         );
  OAI22_X1 U9759 ( .A1(n8251), .A2(n8606), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8338), .ZN(n8208) );
  OAI22_X1 U9760 ( .A1(n8596), .A2(n8234), .B1(n8233), .B2(n8595), .ZN(n8207)
         );
  AOI211_X1 U9761 ( .C1(n8610), .C2(n8238), .A(n8208), .B(n8207), .ZN(n8209)
         );
  NAND2_X1 U9762 ( .A1(n8210), .A2(n8209), .ZN(P2_U3230) );
  INV_X1 U9763 ( .A(n8474), .ZN(n8212) );
  OAI22_X1 U9764 ( .A1(n8436), .A2(n8619), .B1(n8235), .B2(n8621), .ZN(n8468)
         );
  AOI22_X1 U9765 ( .A1(n8468), .A2(n8253), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8211) );
  OAI21_X1 U9766 ( .B1(n8212), .B2(n8251), .A(n8211), .ZN(n8219) );
  NOR2_X1 U9767 ( .A1(n8242), .A2(n8213), .ZN(n8217) );
  NOR2_X1 U9768 ( .A1(n8214), .A2(n8244), .ZN(n8216) );
  MUX2_X1 U9769 ( .A(n8217), .B(n8216), .S(n8215), .Z(n8218) );
  AOI211_X1 U9770 ( .C1(n8473), .C2(n8238), .A(n8219), .B(n8218), .ZN(n8220)
         );
  INV_X1 U9771 ( .A(n8220), .ZN(P2_U3231) );
  XNOR2_X1 U9772 ( .A(n8222), .B(n8221), .ZN(n8228) );
  INV_X1 U9773 ( .A(n8548), .ZN(n8224) );
  OAI22_X1 U9774 ( .A1(n8251), .A2(n8224), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8223), .ZN(n8226) );
  OAI22_X1 U9775 ( .A1(n8249), .A2(n8233), .B1(n8234), .B2(n8232), .ZN(n8225)
         );
  AOI211_X1 U9776 ( .C1(n8681), .C2(n8238), .A(n8226), .B(n8225), .ZN(n8227)
         );
  OAI21_X1 U9777 ( .B1(n8228), .B2(n8244), .A(n8227), .ZN(P2_U3235) );
  INV_X1 U9778 ( .A(n8512), .ZN(n8231) );
  OAI22_X1 U9779 ( .A1(n8251), .A2(n8231), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8230), .ZN(n8237) );
  OAI22_X1 U9780 ( .A1(n8235), .A2(n8234), .B1(n8233), .B2(n8232), .ZN(n8236)
         );
  AOI211_X1 U9781 ( .C1(n8511), .C2(n8238), .A(n8237), .B(n8236), .ZN(n8241)
         );
  NAND3_X1 U9782 ( .A1(n8239), .A2(n8256), .A3(n8493), .ZN(n8240) );
  OAI211_X1 U9783 ( .C1(n4711), .C2(n8244), .A(n8241), .B(n8240), .ZN(P2_U3237) );
  NOR3_X1 U9784 ( .A1(n8243), .A2(n8620), .A3(n8242), .ZN(n8248) );
  AOI21_X1 U9785 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8247) );
  OAI21_X1 U9786 ( .B1(n8248), .B2(n8247), .A(n4343), .ZN(n8255) );
  OAI22_X1 U9787 ( .A1(n8620), .A2(n8621), .B1(n8249), .B2(n8619), .ZN(n8580)
         );
  NOR2_X1 U9788 ( .A1(n8250), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8355) );
  NOR2_X1 U9789 ( .A1(n8251), .A2(n8585), .ZN(n8252) );
  AOI211_X1 U9790 ( .C1(n8253), .C2(n8580), .A(n8355), .B(n8252), .ZN(n8254)
         );
  OAI211_X1 U9791 ( .C1(n8754), .C2(n8270), .A(n8255), .B(n8254), .ZN(P2_U3240) );
  NAND2_X1 U9792 ( .A1(n8256), .A2(n8279), .ZN(n8260) );
  NAND2_X1 U9793 ( .A1(n5866), .A2(n8257), .ZN(n8259) );
  MUX2_X1 U9794 ( .A(n8260), .B(n8259), .S(n8258), .Z(n8269) );
  INV_X1 U9795 ( .A(n8261), .ZN(n8263) );
  OAI22_X1 U9796 ( .A1(n8264), .A2(n8263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8262), .ZN(n8265) );
  AOI21_X1 U9797 ( .B1(n8267), .B2(n8266), .A(n8265), .ZN(n8268) );
  OAI211_X1 U9798 ( .C1(n8766), .C2(n8270), .A(n8269), .B(n8268), .ZN(P2_U3243) );
  MUX2_X1 U9799 ( .A(n8271), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8291), .Z(
        P2_U3582) );
  MUX2_X1 U9800 ( .A(n8272), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8291), .Z(
        P2_U3580) );
  MUX2_X1 U9801 ( .A(n8273), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8291), .Z(
        P2_U3579) );
  MUX2_X1 U9802 ( .A(n8274), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8291), .Z(
        P2_U3578) );
  MUX2_X1 U9803 ( .A(n8275), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8291), .Z(
        P2_U3577) );
  MUX2_X1 U9804 ( .A(n8492), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8291), .Z(
        P2_U3576) );
  MUX2_X1 U9805 ( .A(n8505), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8291), .Z(
        P2_U3575) );
  MUX2_X1 U9806 ( .A(n8493), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8291), .Z(
        P2_U3574) );
  MUX2_X1 U9807 ( .A(n8540), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8291), .Z(
        P2_U3573) );
  MUX2_X1 U9808 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8276), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9809 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8539), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9810 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8277), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9811 ( .A(n5315), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8291), .Z(
        P2_U3569) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8278), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9813 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8279), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9814 ( .A(n8280), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8291), .Z(
        P2_U3566) );
  MUX2_X1 U9815 ( .A(n8281), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8291), .Z(
        P2_U3565) );
  MUX2_X1 U9816 ( .A(n8282), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8291), .Z(
        P2_U3564) );
  MUX2_X1 U9817 ( .A(n8283), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8291), .Z(
        P2_U3563) );
  MUX2_X1 U9818 ( .A(n8284), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8291), .Z(
        P2_U3562) );
  MUX2_X1 U9819 ( .A(n8285), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8291), .Z(
        P2_U3561) );
  MUX2_X1 U9820 ( .A(n8286), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8291), .Z(
        P2_U3560) );
  MUX2_X1 U9821 ( .A(n8287), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8291), .Z(
        P2_U3559) );
  MUX2_X1 U9822 ( .A(n8288), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8291), .Z(
        P2_U3558) );
  MUX2_X1 U9823 ( .A(n9741), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8291), .Z(
        P2_U3557) );
  MUX2_X1 U9824 ( .A(n5095), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8291), .Z(
        P2_U3556) );
  MUX2_X1 U9825 ( .A(n9743), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8291), .Z(
        P2_U3555) );
  MUX2_X1 U9826 ( .A(n8289), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8291), .Z(
        P2_U3554) );
  MUX2_X1 U9827 ( .A(n8290), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8291), .Z(
        P2_U3553) );
  MUX2_X1 U9828 ( .A(n5481), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8291), .Z(
        P2_U3552) );
  OAI211_X1 U9829 ( .C1(n8294), .C2(n8293), .A(n9722), .B(n8292), .ZN(n8305)
         );
  NOR2_X1 U9830 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8295), .ZN(n8296) );
  AOI21_X1 U9831 ( .B1(n9417), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8296), .ZN(
        n8304) );
  NAND2_X1 U9832 ( .A1(n9424), .A2(n8297), .ZN(n8303) );
  AOI21_X1 U9833 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8301) );
  NAND2_X1 U9834 ( .A1(n9724), .A2(n8301), .ZN(n8302) );
  NAND4_X1 U9835 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(
        P2_U3248) );
  XOR2_X1 U9836 ( .A(n8307), .B(n8306), .Z(n8308) );
  NAND2_X1 U9837 ( .A1(n9722), .A2(n8308), .ZN(n8319) );
  NOR2_X1 U9838 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8309), .ZN(n8310) );
  AOI21_X1 U9839 ( .B1(n9417), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8310), .ZN(
        n8318) );
  NAND2_X1 U9840 ( .A1(n9424), .A2(n8311), .ZN(n8317) );
  INV_X1 U9841 ( .A(n8312), .ZN(n8313) );
  OAI211_X1 U9842 ( .C1(n8315), .C2(n8314), .A(n9724), .B(n8313), .ZN(n8316)
         );
  NAND4_X1 U9843 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(
        P2_U3250) );
  OAI211_X1 U9844 ( .C1(n8322), .C2(n8321), .A(n9722), .B(n8320), .ZN(n8333)
         );
  INV_X1 U9845 ( .A(n8323), .ZN(n8324) );
  AOI21_X1 U9846 ( .B1(n9417), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8324), .ZN(
        n8332) );
  NAND2_X1 U9847 ( .A1(n9424), .A2(n8325), .ZN(n8331) );
  AOI21_X1 U9848 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n8329) );
  NAND2_X1 U9849 ( .A1(n9724), .A2(n8329), .ZN(n8330) );
  NAND4_X1 U9850 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .ZN(
        P2_U3255) );
  NAND2_X1 U9851 ( .A1(n8335), .A2(n8334), .ZN(n8337) );
  XNOR2_X1 U9852 ( .A(n8350), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U9853 ( .A1(n8336), .A2(n8337), .ZN(n8348) );
  OAI211_X1 U9854 ( .C1(n8337), .C2(n8336), .A(n9722), .B(n8348), .ZN(n8347)
         );
  NOR2_X1 U9855 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8338), .ZN(n8345) );
  OAI21_X1 U9856 ( .B1(n8340), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8339), .ZN(
        n8343) );
  XNOR2_X1 U9857 ( .A(n8350), .B(n8341), .ZN(n8342) );
  NOR2_X1 U9858 ( .A1(n8342), .A2(n8343), .ZN(n8351) );
  AOI211_X1 U9859 ( .C1(n8343), .C2(n8342), .A(n8351), .B(n9418), .ZN(n8344)
         );
  AOI211_X1 U9860 ( .C1(n9417), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8345), .B(
        n8344), .ZN(n8346) );
  OAI211_X1 U9861 ( .C1(n9726), .C2(n8350), .A(n8347), .B(n8346), .ZN(P2_U3262) );
  OAI21_X1 U9862 ( .B1(n8607), .B2(n8350), .A(n8348), .ZN(n8362) );
  XNOR2_X1 U9863 ( .A(n8368), .B(n8362), .ZN(n8349) );
  NOR2_X1 U9864 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8349), .ZN(n8364) );
  AOI21_X1 U9865 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8349), .A(n8364), .ZN(
        n8361) );
  INV_X1 U9866 ( .A(n8350), .ZN(n8352) );
  AOI22_X1 U9867 ( .A1(n8368), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8695), .B2(
        n8357), .ZN(n8353) );
  NAND2_X1 U9868 ( .A1(n8354), .A2(n8353), .ZN(n8367) );
  OAI21_X1 U9869 ( .B1(n8354), .B2(n8353), .A(n8367), .ZN(n8359) );
  AOI21_X1 U9870 ( .B1(n9417), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8355), .ZN(
        n8356) );
  OAI21_X1 U9871 ( .B1(n9726), .B2(n8357), .A(n8356), .ZN(n8358) );
  AOI21_X1 U9872 ( .B1(n8359), .B2(n9724), .A(n8358), .ZN(n8360) );
  OAI21_X1 U9873 ( .B1(n8361), .B2(n8370), .A(n8360), .ZN(P2_U3263) );
  NOR2_X1 U9874 ( .A1(n8368), .A2(n8362), .ZN(n8363) );
  NOR2_X1 U9875 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  XOR2_X1 U9876 ( .A(n8366), .B(n8365), .Z(n8371) );
  OAI21_X1 U9877 ( .B1(n8368), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8367), .ZN(
        n8369) );
  OAI22_X1 U9878 ( .A1(n8371), .A2(n8370), .B1(n8372), .B2(n9418), .ZN(n8377)
         );
  NAND2_X1 U9879 ( .A1(n8371), .A2(n9722), .ZN(n8374) );
  AOI21_X1 U9880 ( .B1(n8372), .B2(n9724), .A(n9424), .ZN(n8373) );
  NAND2_X1 U9881 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  MUX2_X1 U9882 ( .A(n8377), .B(n8376), .S(n8375), .Z(n8381) );
  NAND2_X1 U9883 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8378) );
  OAI21_X1 U9884 ( .B1(n9731), .B2(n8379), .A(n8378), .ZN(n8380) );
  INV_X1 U9885 ( .A(n8382), .ZN(n8390) );
  NAND2_X1 U9886 ( .A1(n8726), .A2(n8390), .ZN(n8389) );
  INV_X1 U9887 ( .A(n8383), .ZN(n8384) );
  OR2_X1 U9888 ( .A1(n8385), .A2(n8384), .ZN(n8641) );
  NOR2_X1 U9889 ( .A1(n9766), .A2(n8641), .ZN(n8392) );
  INV_X1 U9890 ( .A(n8386), .ZN(n8722) );
  NOR2_X1 U9891 ( .A1(n8722), .A2(n9762), .ZN(n8387) );
  AOI211_X1 U9892 ( .C1(n9766), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8392), .B(
        n8387), .ZN(n8388) );
  OAI21_X1 U9893 ( .B1(n8638), .B2(n8612), .A(n8388), .ZN(P2_U3265) );
  OAI211_X1 U9894 ( .C1(n8726), .C2(n8390), .A(n8603), .B(n8389), .ZN(n8642)
         );
  NOR2_X1 U9895 ( .A1(n8726), .A2(n9762), .ZN(n8391) );
  AOI211_X1 U9896 ( .C1(n9766), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8392), .B(
        n8391), .ZN(n8393) );
  OAI21_X1 U9897 ( .B1(n8612), .B2(n8642), .A(n8393), .ZN(P2_U3266) );
  NAND2_X1 U9898 ( .A1(n8394), .A2(n9764), .ZN(n8402) );
  INV_X1 U9899 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8395) );
  OAI22_X1 U9900 ( .A1(n8396), .A2(n9755), .B1(n8395), .B2(n9757), .ZN(n8399)
         );
  NOR2_X1 U9901 ( .A1(n8397), .A2(n8612), .ZN(n8398) );
  AOI211_X1 U9902 ( .C1(n8609), .C2(n8400), .A(n8399), .B(n8398), .ZN(n8401)
         );
  OAI211_X1 U9903 ( .C1(n8403), .C2(n9766), .A(n8402), .B(n8401), .ZN(P2_U3267) );
  INV_X1 U9904 ( .A(n8404), .ZN(n8414) );
  NAND2_X1 U9905 ( .A1(n8405), .A2(n9764), .ZN(n8413) );
  NOR2_X1 U9906 ( .A1(n8406), .A2(n9762), .ZN(n8410) );
  OAI22_X1 U9907 ( .A1(n8408), .A2(n9755), .B1(n8407), .B2(n9757), .ZN(n8409)
         );
  AOI211_X1 U9908 ( .C1(n8411), .C2(n8634), .A(n8410), .B(n8409), .ZN(n8412)
         );
  OAI211_X1 U9909 ( .C1(n8414), .C2(n9766), .A(n8413), .B(n8412), .ZN(P2_U3268) );
  NAND2_X1 U9910 ( .A1(n8415), .A2(n8421), .ZN(n8416) );
  NAND2_X1 U9911 ( .A1(n8416), .A2(n9745), .ZN(n8417) );
  OR2_X1 U9912 ( .A1(n4334), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U9913 ( .A1(n8419), .A2(n8418), .ZN(n8644) );
  INV_X1 U9914 ( .A(n8644), .ZN(n8431) );
  OAI21_X1 U9915 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8646) );
  NAND2_X1 U9916 ( .A1(n8646), .A2(n9764), .ZN(n8430) );
  AOI211_X1 U9917 ( .C1(n8424), .C2(n4287), .A(n9826), .B(n4606), .ZN(n8645)
         );
  INV_X1 U9918 ( .A(n8425), .ZN(n8426) );
  AOI22_X1 U9919 ( .A1(n8426), .A2(n8570), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9766), .ZN(n8427) );
  OAI21_X1 U9920 ( .B1(n8730), .B2(n9762), .A(n8427), .ZN(n8428) );
  AOI21_X1 U9921 ( .B1(n8645), .B2(n8634), .A(n8428), .ZN(n8429) );
  OAI211_X1 U9922 ( .C1(n9766), .C2(n8431), .A(n8430), .B(n8429), .ZN(P2_U3269) );
  OR2_X1 U9923 ( .A1(n8454), .A2(n8734), .ZN(n8432) );
  AND2_X1 U9924 ( .A1(n8650), .A2(n8433), .ZN(n8438) );
  XNOR2_X1 U9925 ( .A(n8434), .B(n4625), .ZN(n8435) );
  OAI222_X1 U9926 ( .A1(n8619), .A2(n8437), .B1(n8621), .B2(n8436), .C1(n8566), 
        .C2(n8435), .ZN(n8649) );
  AOI211_X1 U9927 ( .C1(n8570), .C2(n8439), .A(n8438), .B(n8649), .ZN(n8446)
         );
  OAI21_X1 U9928 ( .B1(n8442), .B2(n8441), .A(n8440), .ZN(n8651) );
  NAND2_X1 U9929 ( .A1(n8651), .A2(n9764), .ZN(n8445) );
  AOI22_X1 U9930 ( .A1(n8443), .A2(n8609), .B1(n9766), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8444) );
  OAI211_X1 U9931 ( .C1(n9766), .C2(n8446), .A(n8445), .B(n8444), .ZN(P2_U3270) );
  XNOR2_X1 U9932 ( .A(n8447), .B(n8452), .ZN(n8448) );
  NAND2_X1 U9933 ( .A1(n8448), .A2(n9745), .ZN(n8450) );
  NAND2_X1 U9934 ( .A1(n8450), .A2(n8449), .ZN(n8654) );
  INV_X1 U9935 ( .A(n8654), .ZN(n8463) );
  OAI21_X1 U9936 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8656) );
  NAND2_X1 U9937 ( .A1(n8656), .A2(n9764), .ZN(n8462) );
  INV_X1 U9938 ( .A(n8472), .ZN(n8455) );
  AOI211_X1 U9939 ( .C1(n8456), .C2(n8455), .A(n9826), .B(n8454), .ZN(n8655)
         );
  INV_X1 U9940 ( .A(n8457), .ZN(n8458) );
  AOI22_X1 U9941 ( .A1(n9766), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8458), .B2(
        n8570), .ZN(n8459) );
  OAI21_X1 U9942 ( .B1(n8738), .B2(n9762), .A(n8459), .ZN(n8460) );
  AOI21_X1 U9943 ( .B1(n8655), .B2(n8634), .A(n8460), .ZN(n8461) );
  OAI211_X1 U9944 ( .C1(n9766), .C2(n8463), .A(n8462), .B(n8461), .ZN(P2_U3271) );
  INV_X1 U9945 ( .A(n8464), .ZN(n8465) );
  AOI211_X1 U9946 ( .C1(n8467), .C2(n8466), .A(n8566), .B(n8465), .ZN(n8469)
         );
  OR2_X1 U9947 ( .A1(n8469), .A2(n8468), .ZN(n8659) );
  INV_X1 U9948 ( .A(n8659), .ZN(n8479) );
  XNOR2_X1 U9949 ( .A(n8471), .B(n8470), .ZN(n8661) );
  NAND2_X1 U9950 ( .A1(n8661), .A2(n9764), .ZN(n8478) );
  AOI211_X1 U9951 ( .C1(n8473), .C2(n8481), .A(n9826), .B(n8472), .ZN(n8660)
         );
  INV_X1 U9952 ( .A(n8473), .ZN(n8742) );
  AOI22_X1 U9953 ( .A1(n9766), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8474), .B2(
        n8570), .ZN(n8475) );
  OAI21_X1 U9954 ( .B1(n8742), .B2(n9762), .A(n8475), .ZN(n8476) );
  AOI21_X1 U9955 ( .B1(n8660), .B2(n8634), .A(n8476), .ZN(n8477) );
  OAI211_X1 U9956 ( .C1(n9766), .C2(n8479), .A(n8478), .B(n8477), .ZN(P2_U3272) );
  OAI21_X1 U9957 ( .B1(n4649), .B2(n8487), .A(n8480), .ZN(n8668) );
  INV_X1 U9958 ( .A(n8481), .ZN(n8482) );
  AOI211_X1 U9959 ( .C1(n8665), .C2(n8508), .A(n9826), .B(n8482), .ZN(n8664)
         );
  INV_X1 U9960 ( .A(n8483), .ZN(n8484) );
  AOI22_X1 U9961 ( .A1(n9766), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8484), .B2(
        n8570), .ZN(n8485) );
  OAI21_X1 U9962 ( .B1(n8486), .B2(n9762), .A(n8485), .ZN(n8496) );
  INV_X1 U9963 ( .A(n8503), .ZN(n8489) );
  OAI21_X1 U9964 ( .B1(n8489), .B2(n8488), .A(n8487), .ZN(n8491) );
  NAND2_X1 U9965 ( .A1(n8491), .A2(n8490), .ZN(n8494) );
  AOI222_X1 U9966 ( .A1(n9745), .A2(n8494), .B1(n8493), .B2(n9742), .C1(n8492), 
        .C2(n9740), .ZN(n8667) );
  NOR2_X1 U9967 ( .A1(n8667), .A2(n9766), .ZN(n8495) );
  AOI211_X1 U9968 ( .C1(n8664), .C2(n8634), .A(n8496), .B(n8495), .ZN(n8497)
         );
  OAI21_X1 U9969 ( .B1(n8668), .B2(n8584), .A(n8497), .ZN(P2_U3273) );
  XNOR2_X1 U9970 ( .A(n8499), .B(n8498), .ZN(n8671) );
  INV_X1 U9971 ( .A(n8671), .ZN(n8517) );
  NAND2_X1 U9972 ( .A1(n8521), .A2(n8500), .ZN(n8502) );
  NAND2_X1 U9973 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  NAND3_X1 U9974 ( .A1(n8504), .A2(n9745), .A3(n8503), .ZN(n8507) );
  AOI22_X1 U9975 ( .A1(n8505), .A2(n9740), .B1(n9742), .B2(n8540), .ZN(n8506)
         );
  NAND2_X1 U9976 ( .A1(n8507), .A2(n8506), .ZN(n8669) );
  INV_X1 U9977 ( .A(n8527), .ZN(n8510) );
  INV_X1 U9978 ( .A(n8508), .ZN(n8509) );
  AOI211_X1 U9979 ( .C1(n8511), .C2(n8510), .A(n9826), .B(n8509), .ZN(n8670)
         );
  NAND2_X1 U9980 ( .A1(n8670), .A2(n8634), .ZN(n8514) );
  AOI22_X1 U9981 ( .A1(n9766), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8512), .B2(
        n8570), .ZN(n8513) );
  OAI211_X1 U9982 ( .C1(n8747), .C2(n9762), .A(n8514), .B(n8513), .ZN(n8515)
         );
  AOI21_X1 U9983 ( .B1(n8669), .B2(n9757), .A(n8515), .ZN(n8516) );
  OAI21_X1 U9984 ( .B1(n8517), .B2(n8584), .A(n8516), .ZN(P2_U3274) );
  XOR2_X1 U9985 ( .A(n8523), .B(n8518), .Z(n8678) );
  NAND2_X1 U9986 ( .A1(n8520), .A2(n8519), .ZN(n8524) );
  INV_X1 U9987 ( .A(n8521), .ZN(n8522) );
  AOI21_X1 U9988 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8525) );
  OAI222_X1 U9989 ( .A1(n8621), .A2(n8567), .B1(n8619), .B2(n8526), .C1(n8566), 
        .C2(n8525), .ZN(n8674) );
  AOI211_X1 U9990 ( .C1(n8676), .C2(n4594), .A(n9826), .B(n8527), .ZN(n8675)
         );
  NAND2_X1 U9991 ( .A1(n8675), .A2(n8634), .ZN(n8531) );
  INV_X1 U9992 ( .A(n8528), .ZN(n8529) );
  AOI22_X1 U9993 ( .A1(n9766), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8529), .B2(
        n8570), .ZN(n8530) );
  OAI211_X1 U9994 ( .C1(n8532), .C2(n9762), .A(n8531), .B(n8530), .ZN(n8533)
         );
  AOI21_X1 U9995 ( .B1(n8674), .B2(n9757), .A(n8533), .ZN(n8534) );
  OAI21_X1 U9996 ( .B1(n8678), .B2(n8584), .A(n8534), .ZN(P2_U3275) );
  AND2_X1 U9997 ( .A1(n8536), .A2(n8535), .ZN(n8561) );
  NAND2_X1 U9998 ( .A1(n8561), .A2(n8537), .ZN(n8538) );
  XNOR2_X1 U9999 ( .A(n8538), .B(n8542), .ZN(n8541) );
  AOI222_X1 U10000 ( .A1(n9745), .A2(n8541), .B1(n8540), .B2(n9740), .C1(n8539), .C2(n9742), .ZN(n8683) );
  INV_X1 U10001 ( .A(n8685), .ZN(n8544) );
  NAND2_X1 U10002 ( .A1(n8543), .A2(n8542), .ZN(n8679) );
  NAND3_X1 U10003 ( .A1(n8544), .A2(n9764), .A3(n8679), .ZN(n8554) );
  NAND2_X1 U10004 ( .A1(n8568), .A2(n8681), .ZN(n8545) );
  NAND2_X1 U10005 ( .A1(n8545), .A2(n8603), .ZN(n8546) );
  NOR2_X1 U10006 ( .A1(n8547), .A2(n8546), .ZN(n8680) );
  INV_X1 U10007 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10008 ( .A1(n8681), .A2(n8609), .ZN(n8550) );
  NAND2_X1 U10009 ( .A1(n8570), .A2(n8548), .ZN(n8549) );
  OAI211_X1 U10010 ( .C1(n9757), .C2(n8551), .A(n8550), .B(n8549), .ZN(n8552)
         );
  AOI21_X1 U10011 ( .B1(n8680), .B2(n8634), .A(n8552), .ZN(n8553) );
  OAI211_X1 U10012 ( .C1(n9766), .C2(n8683), .A(n8554), .B(n8553), .ZN(
        P2_U3276) );
  XNOR2_X1 U10013 ( .A(n8556), .B(n8555), .ZN(n8690) );
  NAND2_X1 U10014 ( .A1(n8557), .A2(n8558), .ZN(n8560) );
  AND2_X1 U10015 ( .A1(n8560), .A2(n8559), .ZN(n8564) );
  INV_X1 U10016 ( .A(n8561), .ZN(n8562) );
  AOI21_X1 U10017 ( .B1(n8564), .B2(n8563), .A(n8562), .ZN(n8565) );
  OAI222_X1 U10018 ( .A1(n8619), .A2(n8567), .B1(n8621), .B2(n8596), .C1(n8566), .C2(n8565), .ZN(n8686) );
  INV_X1 U10019 ( .A(n8568), .ZN(n8569) );
  AOI211_X1 U10020 ( .C1(n8688), .C2(n8587), .A(n9826), .B(n8569), .ZN(n8687)
         );
  NAND2_X1 U10021 ( .A1(n8687), .A2(n8634), .ZN(n8573) );
  AOI22_X1 U10022 ( .A1(n9766), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8571), .B2(
        n8570), .ZN(n8572) );
  OAI211_X1 U10023 ( .C1(n8574), .C2(n9762), .A(n8573), .B(n8572), .ZN(n8575)
         );
  AOI21_X1 U10024 ( .B1(n8686), .B2(n9757), .A(n8575), .ZN(n8576) );
  OAI21_X1 U10025 ( .B1(n8690), .B2(n8584), .A(n8576), .ZN(P2_U3277) );
  NAND2_X1 U10026 ( .A1(n8557), .A2(n8577), .ZN(n8579) );
  INV_X1 U10027 ( .A(n8583), .ZN(n8578) );
  XNOR2_X1 U10028 ( .A(n8579), .B(n8578), .ZN(n8581) );
  AOI21_X1 U10029 ( .B1(n8581), .B2(n9745), .A(n8580), .ZN(n8692) );
  XOR2_X1 U10030 ( .A(n8583), .B(n8582), .Z(n8693) );
  OR2_X1 U10031 ( .A1(n8693), .A2(n8584), .ZN(n8592) );
  OAI22_X1 U10032 ( .A1(n9757), .A2(n8586), .B1(n8585), .B2(n9755), .ZN(n8589)
         );
  OAI211_X1 U10033 ( .C1(n8605), .C2(n8754), .A(n8603), .B(n8587), .ZN(n8691)
         );
  NOR2_X1 U10034 ( .A1(n8691), .A2(n8612), .ZN(n8588) );
  AOI211_X1 U10035 ( .C1(n8609), .C2(n8590), .A(n8589), .B(n8588), .ZN(n8591)
         );
  OAI211_X1 U10036 ( .C1(n9766), .C2(n8692), .A(n8592), .B(n8591), .ZN(
        P2_U3278) );
  XNOR2_X1 U10037 ( .A(n8594), .B(n8593), .ZN(n8598) );
  OAI22_X1 U10038 ( .A1(n8596), .A2(n8619), .B1(n8595), .B2(n8621), .ZN(n8597)
         );
  AOI21_X1 U10039 ( .B1(n8598), .B2(n9745), .A(n8597), .ZN(n8699) );
  AND2_X1 U10040 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  OR2_X1 U10041 ( .A1(n8602), .A2(n8601), .ZN(n8697) );
  OAI21_X1 U10042 ( .B1(n8627), .B2(n8758), .A(n8603), .ZN(n8604) );
  OR2_X1 U10043 ( .A1(n8605), .A2(n8604), .ZN(n8698) );
  OAI22_X1 U10044 ( .A1(n9757), .A2(n8607), .B1(n8606), .B2(n9755), .ZN(n8608)
         );
  AOI21_X1 U10045 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8611) );
  OAI21_X1 U10046 ( .B1(n8698), .B2(n8612), .A(n8611), .ZN(n8613) );
  AOI21_X1 U10047 ( .B1(n8697), .B2(n9764), .A(n8613), .ZN(n8614) );
  OAI21_X1 U10048 ( .B1(n9766), .B2(n8699), .A(n8614), .ZN(P2_U3279) );
  OAI21_X1 U10049 ( .B1(n8616), .B2(n8617), .A(n8615), .ZN(n8703) );
  XNOR2_X1 U10050 ( .A(n8618), .B(n8617), .ZN(n8624) );
  OAI22_X1 U10051 ( .A1(n8622), .A2(n8621), .B1(n8620), .B2(n8619), .ZN(n8623)
         );
  AOI21_X1 U10052 ( .B1(n8624), .B2(n9745), .A(n8623), .ZN(n8625) );
  OAI21_X1 U10053 ( .B1(n8703), .B2(n8626), .A(n8625), .ZN(n8705) );
  NAND2_X1 U10054 ( .A1(n8705), .A2(n9757), .ZN(n8636) );
  AOI211_X1 U10055 ( .C1(n8629), .C2(n8628), .A(n9826), .B(n8627), .ZN(n8706)
         );
  INV_X1 U10056 ( .A(n8629), .ZN(n8762) );
  NOR2_X1 U10057 ( .A1(n8762), .A2(n9762), .ZN(n8633) );
  OAI22_X1 U10058 ( .A1(n9757), .A2(n8631), .B1(n8630), .B2(n9755), .ZN(n8632)
         );
  AOI211_X1 U10059 ( .C1(n8706), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8635)
         );
  OAI211_X1 U10060 ( .C1(n8703), .C2(n8637), .A(n8636), .B(n8635), .ZN(
        P2_U3280) );
  INV_X1 U10061 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8639) );
  MUX2_X1 U10062 ( .A(n8639), .B(n8720), .S(n9855), .Z(n8640) );
  OAI21_X1 U10063 ( .B1(n8722), .B2(n8719), .A(n8640), .ZN(P2_U3551) );
  MUX2_X1 U10064 ( .A(n9911), .B(n8723), .S(n9855), .Z(n8643) );
  OAI21_X1 U10065 ( .B1(n8726), .B2(n8719), .A(n8643), .ZN(P2_U3550) );
  INV_X1 U10066 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8647) );
  AOI211_X1 U10067 ( .C1(n8646), .C2(n9838), .A(n8645), .B(n8644), .ZN(n8727)
         );
  MUX2_X1 U10068 ( .A(n8647), .B(n8727), .S(n9855), .Z(n8648) );
  OAI21_X1 U10069 ( .B1(n8730), .B2(n8719), .A(n8648), .ZN(P2_U3547) );
  INV_X1 U10070 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8652) );
  AOI211_X1 U10071 ( .C1(n8651), .C2(n9838), .A(n8650), .B(n8649), .ZN(n8731)
         );
  MUX2_X1 U10072 ( .A(n8652), .B(n8731), .S(n9855), .Z(n8653) );
  OAI21_X1 U10073 ( .B1(n8734), .B2(n8719), .A(n8653), .ZN(P2_U3546) );
  INV_X1 U10074 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8657) );
  AOI211_X1 U10075 ( .C1(n8656), .C2(n9838), .A(n8655), .B(n8654), .ZN(n8735)
         );
  MUX2_X1 U10076 ( .A(n8657), .B(n8735), .S(n9855), .Z(n8658) );
  OAI21_X1 U10077 ( .B1(n8738), .B2(n8719), .A(n8658), .ZN(P2_U3545) );
  INV_X1 U10078 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8662) );
  AOI211_X1 U10079 ( .C1(n8661), .C2(n9838), .A(n8660), .B(n8659), .ZN(n8739)
         );
  MUX2_X1 U10080 ( .A(n8662), .B(n8739), .S(n9855), .Z(n8663) );
  OAI21_X1 U10081 ( .B1(n8742), .B2(n8719), .A(n8663), .ZN(P2_U3544) );
  AOI21_X1 U10082 ( .B1(n9812), .B2(n8665), .A(n8664), .ZN(n8666) );
  OAI211_X1 U10083 ( .C1(n8668), .C2(n9815), .A(n8667), .B(n8666), .ZN(n8743)
         );
  MUX2_X1 U10084 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8743), .S(n9855), .Z(
        P2_U3543) );
  INV_X1 U10085 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8672) );
  AOI211_X1 U10086 ( .C1(n8671), .C2(n9838), .A(n8670), .B(n8669), .ZN(n8744)
         );
  MUX2_X1 U10087 ( .A(n8672), .B(n8744), .S(n9855), .Z(n8673) );
  OAI21_X1 U10088 ( .B1(n8747), .B2(n8719), .A(n8673), .ZN(P2_U3542) );
  AOI211_X1 U10089 ( .C1(n9812), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8677)
         );
  OAI21_X1 U10090 ( .B1(n8678), .B2(n9815), .A(n8677), .ZN(n8748) );
  MUX2_X1 U10091 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8748), .S(n9855), .Z(
        P2_U3541) );
  NAND2_X1 U10092 ( .A1(n8679), .A2(n9838), .ZN(n8684) );
  AOI21_X1 U10093 ( .B1(n9812), .B2(n8681), .A(n8680), .ZN(n8682) );
  OAI211_X1 U10094 ( .C1(n8685), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8749)
         );
  MUX2_X1 U10095 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8749), .S(n9855), .Z(
        P2_U3540) );
  AOI211_X1 U10096 ( .C1(n9812), .C2(n8688), .A(n8687), .B(n8686), .ZN(n8689)
         );
  OAI21_X1 U10097 ( .B1(n9815), .B2(n8690), .A(n8689), .ZN(n8750) );
  MUX2_X1 U10098 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8750), .S(n9855), .Z(
        P2_U3539) );
  OAI211_X1 U10099 ( .C1(n8693), .C2(n9815), .A(n8692), .B(n8691), .ZN(n8694)
         );
  INV_X1 U10100 ( .A(n8694), .ZN(n8751) );
  MUX2_X1 U10101 ( .A(n8695), .B(n8751), .S(n9855), .Z(n8696) );
  OAI21_X1 U10102 ( .B1(n8754), .B2(n8719), .A(n8696), .ZN(P2_U3538) );
  NAND2_X1 U10103 ( .A1(n8697), .A2(n9838), .ZN(n8700) );
  NAND3_X1 U10104 ( .A1(n8700), .A2(n8699), .A3(n8698), .ZN(n8755) );
  MUX2_X1 U10105 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8755), .S(n9855), .Z(n8701) );
  INV_X1 U10106 ( .A(n8701), .ZN(n8702) );
  OAI21_X1 U10107 ( .B1(n8758), .B2(n8719), .A(n8702), .ZN(P2_U3537) );
  INV_X1 U10108 ( .A(n8703), .ZN(n8707) );
  INV_X1 U10109 ( .A(n8704), .ZN(n9831) );
  AOI211_X1 U10110 ( .C1(n8707), .C2(n9831), .A(n8706), .B(n8705), .ZN(n8759)
         );
  MUX2_X1 U10111 ( .A(n8708), .B(n8759), .S(n9855), .Z(n8709) );
  OAI21_X1 U10112 ( .B1(n8762), .B2(n8719), .A(n8709), .ZN(P2_U3536) );
  AOI211_X1 U10113 ( .C1(n9838), .C2(n8712), .A(n8711), .B(n8710), .ZN(n8763)
         );
  MUX2_X1 U10114 ( .A(n8713), .B(n8763), .S(n9855), .Z(n8714) );
  OAI21_X1 U10115 ( .B1(n8766), .B2(n8719), .A(n8714), .ZN(P2_U3535) );
  AOI211_X1 U10116 ( .C1(n8717), .C2(n9838), .A(n8716), .B(n8715), .ZN(n8767)
         );
  MUX2_X1 U10117 ( .A(n7096), .B(n8767), .S(n9855), .Z(n8718) );
  OAI21_X1 U10118 ( .B1(n8771), .B2(n8719), .A(n8718), .ZN(P2_U3534) );
  INV_X1 U10119 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8721) );
  INV_X1 U10120 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U10121 ( .A(n8724), .B(n8723), .S(n9840), .Z(n8725) );
  OAI21_X1 U10122 ( .B1(n8726), .B2(n8770), .A(n8725), .ZN(P2_U3518) );
  MUX2_X1 U10123 ( .A(n8728), .B(n8727), .S(n9840), .Z(n8729) );
  OAI21_X1 U10124 ( .B1(n8730), .B2(n8770), .A(n8729), .ZN(P2_U3515) );
  MUX2_X1 U10125 ( .A(n8732), .B(n8731), .S(n9840), .Z(n8733) );
  OAI21_X1 U10126 ( .B1(n8734), .B2(n8770), .A(n8733), .ZN(P2_U3514) );
  MUX2_X1 U10127 ( .A(n8736), .B(n8735), .S(n9840), .Z(n8737) );
  OAI21_X1 U10128 ( .B1(n8738), .B2(n8770), .A(n8737), .ZN(P2_U3513) );
  MUX2_X1 U10129 ( .A(n8740), .B(n8739), .S(n9840), .Z(n8741) );
  OAI21_X1 U10130 ( .B1(n8742), .B2(n8770), .A(n8741), .ZN(P2_U3512) );
  MUX2_X1 U10131 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8743), .S(n9840), .Z(
        P2_U3511) );
  INV_X1 U10132 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8745) );
  MUX2_X1 U10133 ( .A(n8745), .B(n8744), .S(n9840), .Z(n8746) );
  OAI21_X1 U10134 ( .B1(n8747), .B2(n8770), .A(n8746), .ZN(P2_U3510) );
  MUX2_X1 U10135 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8748), .S(n9840), .Z(
        P2_U3509) );
  MUX2_X1 U10136 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8749), .S(n9840), .Z(
        P2_U3508) );
  MUX2_X1 U10137 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8750), .S(n9840), .Z(
        P2_U3507) );
  INV_X1 U10138 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8752) );
  MUX2_X1 U10139 ( .A(n8752), .B(n8751), .S(n9840), .Z(n8753) );
  OAI21_X1 U10140 ( .B1(n8754), .B2(n8770), .A(n8753), .ZN(P2_U3505) );
  MUX2_X1 U10141 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8755), .S(n9840), .Z(n8756) );
  INV_X1 U10142 ( .A(n8756), .ZN(n8757) );
  OAI21_X1 U10143 ( .B1(n8758), .B2(n8770), .A(n8757), .ZN(P2_U3502) );
  INV_X1 U10144 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8760) );
  MUX2_X1 U10145 ( .A(n8760), .B(n8759), .S(n9840), .Z(n8761) );
  OAI21_X1 U10146 ( .B1(n8762), .B2(n8770), .A(n8761), .ZN(P2_U3499) );
  MUX2_X1 U10147 ( .A(n8764), .B(n8763), .S(n9840), .Z(n8765) );
  OAI21_X1 U10148 ( .B1(n8766), .B2(n8770), .A(n8765), .ZN(P2_U3496) );
  INV_X1 U10149 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8768) );
  MUX2_X1 U10150 ( .A(n8768), .B(n8767), .S(n9840), .Z(n8769) );
  OAI21_X1 U10151 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(P2_U3493) );
  INV_X1 U10152 ( .A(n8772), .ZN(n8777) );
  INV_X1 U10153 ( .A(n8773), .ZN(n8774) );
  NOR4_X1 U10154 ( .A1(n8774), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5529), .A4(
        P2_U3152), .ZN(n8775) );
  AOI21_X1 U10155 ( .B1(n8780), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8775), .ZN(
        n8776) );
  OAI21_X1 U10156 ( .B1(n8777), .B2(n8783), .A(n8776), .ZN(P2_U3327) );
  INV_X1 U10157 ( .A(n7845), .ZN(n9401) );
  AOI22_X1 U10158 ( .A1(n8778), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8780), .ZN(n8779) );
  OAI21_X1 U10159 ( .B1(n9401), .B2(n8783), .A(n8779), .ZN(P2_U3328) );
  AOI22_X1 U10160 ( .A1(n8781), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8780), .ZN(n8782) );
  OAI21_X1 U10161 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(P2_U3329) );
  MUX2_X1 U10162 ( .A(n8785), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10163 ( .A(n8787), .B(n8786), .ZN(n8788) );
  XNOR2_X1 U10164 ( .A(n8789), .B(n8788), .ZN(n8794) );
  AOI22_X1 U10165 ( .A1(n8927), .A2(n8901), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8791) );
  NAND2_X1 U10166 ( .A1(n9102), .A2(n8907), .ZN(n8790) );
  OAI211_X1 U10167 ( .C1(n9100), .C2(n8904), .A(n8791), .B(n8790), .ZN(n8792)
         );
  AOI21_X1 U10168 ( .B1(n9310), .B2(n8894), .A(n8792), .ZN(n8793) );
  OAI21_X1 U10169 ( .B1(n8794), .B2(n8923), .A(n8793), .ZN(P1_U3212) );
  NAND2_X1 U10170 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  XOR2_X1 U10171 ( .A(n8798), .B(n8797), .Z(n8804) );
  NAND2_X1 U10172 ( .A1(n8901), .A2(n9454), .ZN(n8800) );
  OAI211_X1 U10173 ( .C1(n9262), .C2(n8904), .A(n8800), .B(n8799), .ZN(n8802)
         );
  INV_X1 U10174 ( .A(n10034), .ZN(n9462) );
  NOR2_X1 U10175 ( .A1(n9462), .A2(n8910), .ZN(n8801) );
  AOI211_X1 U10176 ( .C1(n10032), .C2(n8907), .A(n8802), .B(n8801), .ZN(n8803)
         );
  OAI21_X1 U10177 ( .B1(n8804), .B2(n8923), .A(n8803), .ZN(P1_U3213) );
  INV_X1 U10178 ( .A(n8805), .ZN(n8806) );
  NOR2_X1 U10179 ( .A1(n8807), .A2(n8806), .ZN(n8809) );
  XNOR2_X1 U10180 ( .A(n8809), .B(n8808), .ZN(n8814) );
  NAND2_X1 U10181 ( .A1(n9164), .A2(n8918), .ZN(n8811) );
  AOI22_X1 U10182 ( .A1(n9158), .A2(n8901), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8810) );
  OAI211_X1 U10183 ( .C1(n8920), .C2(n9154), .A(n8811), .B(n8810), .ZN(n8812)
         );
  AOI21_X1 U10184 ( .B1(n9328), .B2(n8894), .A(n8812), .ZN(n8813) );
  OAI21_X1 U10185 ( .B1(n8814), .B2(n8923), .A(n8813), .ZN(P1_U3214) );
  INV_X1 U10186 ( .A(n8815), .ZN(n8816) );
  AOI21_X1 U10187 ( .B1(n8818), .B2(n4262), .A(n8816), .ZN(n8823) );
  AOI22_X1 U10188 ( .A1(n8918), .A2(n9020), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8820) );
  NAND2_X1 U10189 ( .A1(n8901), .A2(n9017), .ZN(n8819) );
  OAI211_X1 U10190 ( .C1(n8920), .C2(n9221), .A(n8820), .B(n8819), .ZN(n8821)
         );
  AOI21_X1 U10191 ( .B1(n9349), .B2(n8894), .A(n8821), .ZN(n8822) );
  OAI21_X1 U10192 ( .B1(n8823), .B2(n8923), .A(n8822), .ZN(P1_U3217) );
  OAI21_X1 U10193 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(n8827) );
  NAND2_X1 U10194 ( .A1(n8827), .A2(n8898), .ZN(n8831) );
  AOI22_X1 U10195 ( .A1(n8918), .A2(n9629), .B1(n6163), .B2(n8894), .ZN(n8830)
         );
  AOI22_X1 U10196 ( .A1(n8901), .A2(n8937), .B1(n8828), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8829) );
  NAND3_X1 U10197 ( .A1(n8831), .A2(n8830), .A3(n8829), .ZN(P1_U3220) );
  XOR2_X1 U10198 ( .A(n8833), .B(n8832), .Z(n8838) );
  AOI22_X1 U10199 ( .A1(n9158), .A2(n8918), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8835) );
  NAND2_X1 U10200 ( .A1(n8907), .A2(n9191), .ZN(n8834) );
  OAI211_X1 U10201 ( .C1(n9219), .C2(n8916), .A(n8835), .B(n8834), .ZN(n8836)
         );
  AOI21_X1 U10202 ( .B1(n9339), .B2(n8894), .A(n8836), .ZN(n8837) );
  OAI21_X1 U10203 ( .B1(n8838), .B2(n8923), .A(n8837), .ZN(P1_U3221) );
  XOR2_X1 U10204 ( .A(n8840), .B(n8839), .Z(n8845) );
  NAND2_X1 U10205 ( .A1(n8927), .A2(n8918), .ZN(n8842) );
  AOI22_X1 U10206 ( .A1(n9164), .A2(n8901), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8841) );
  OAI211_X1 U10207 ( .C1(n8920), .C2(n9130), .A(n8842), .B(n8841), .ZN(n8843)
         );
  AOI21_X1 U10208 ( .B1(n9319), .B2(n8894), .A(n8843), .ZN(n8844) );
  OAI21_X1 U10209 ( .B1(n8845), .B2(n8923), .A(n8844), .ZN(P1_U3223) );
  INV_X1 U10210 ( .A(n8847), .ZN(n8848) );
  AOI21_X1 U10211 ( .B1(n8849), .B2(n4263), .A(n8848), .ZN(n8854) );
  AOI22_X1 U10212 ( .A1(n8918), .A2(n9015), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8851) );
  NAND2_X1 U10213 ( .A1(n8907), .A2(n9270), .ZN(n8850) );
  OAI211_X1 U10214 ( .C1(n9262), .C2(n8916), .A(n8851), .B(n8850), .ZN(n8852)
         );
  AOI21_X1 U10215 ( .B1(n9365), .B2(n8894), .A(n8852), .ZN(n8853) );
  OAI21_X1 U10216 ( .B1(n8854), .B2(n8923), .A(n8853), .ZN(P1_U3224) );
  XOR2_X1 U10217 ( .A(n8856), .B(n8855), .Z(n8862) );
  OAI22_X1 U10218 ( .A1(n8904), .A2(n9254), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8857), .ZN(n8858) );
  AOI21_X1 U10219 ( .B1(n8901), .B2(n9014), .A(n8858), .ZN(n8859) );
  OAI21_X1 U10220 ( .B1(n8920), .B2(n9247), .A(n8859), .ZN(n8860) );
  AOI21_X1 U10221 ( .B1(n9359), .B2(n8894), .A(n8860), .ZN(n8861) );
  OAI21_X1 U10222 ( .B1(n8862), .B2(n8923), .A(n8861), .ZN(P1_U3226) );
  OAI21_X1 U10223 ( .B1(n8865), .B2(n4267), .A(n8864), .ZN(n8866) );
  NAND2_X1 U10224 ( .A1(n8866), .A2(n8898), .ZN(n8870) );
  AOI22_X1 U10225 ( .A1(n9146), .A2(n8901), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8867) );
  OAI21_X1 U10226 ( .B1(n9112), .B2(n8904), .A(n8867), .ZN(n8868) );
  AOI21_X1 U10227 ( .B1(n9140), .B2(n8907), .A(n8868), .ZN(n8869) );
  OAI211_X1 U10228 ( .C1(n9142), .C2(n8910), .A(n8870), .B(n8869), .ZN(
        P1_U3227) );
  XOR2_X1 U10229 ( .A(n8872), .B(n8871), .Z(n8877) );
  OAI22_X1 U10230 ( .A1(n9204), .A2(n8904), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10001), .ZN(n8873) );
  AOI21_X1 U10231 ( .B1(n8901), .B2(n9018), .A(n8873), .ZN(n8874) );
  OAI21_X1 U10232 ( .B1(n8920), .B2(n9208), .A(n8874), .ZN(n8875) );
  AOI21_X1 U10233 ( .B1(n9344), .B2(n8894), .A(n8875), .ZN(n8876) );
  OAI21_X1 U10234 ( .B1(n8877), .B2(n8923), .A(n8876), .ZN(P1_U3231) );
  NAND2_X1 U10235 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  XOR2_X1 U10236 ( .A(n8881), .B(n8880), .Z(n8886) );
  NAND2_X1 U10237 ( .A1(n9146), .A2(n8918), .ZN(n8883) );
  AOI22_X1 U10238 ( .A1(n9022), .A2(n8901), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8882) );
  OAI211_X1 U10239 ( .C1(n8920), .C2(n9177), .A(n8883), .B(n8882), .ZN(n8884)
         );
  AOI21_X1 U10240 ( .B1(n9334), .B2(n8894), .A(n8884), .ZN(n8885) );
  OAI21_X1 U10241 ( .B1(n8886), .B2(n8923), .A(n8885), .ZN(P1_U3233) );
  NAND2_X1 U10242 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  XOR2_X1 U10243 ( .A(n8890), .B(n8889), .Z(n8896) );
  NAND2_X1 U10244 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9611) );
  OAI21_X1 U10245 ( .B1(n9241), .B2(n8904), .A(n9611), .ZN(n8891) );
  AOI21_X1 U10246 ( .B1(n8901), .B2(n9015), .A(n8891), .ZN(n8892) );
  OAI21_X1 U10247 ( .B1(n8920), .B2(n9233), .A(n8892), .ZN(n8893) );
  AOI21_X1 U10248 ( .B1(n9354), .B2(n8894), .A(n8893), .ZN(n8895) );
  OAI21_X1 U10249 ( .B1(n8896), .B2(n8923), .A(n8895), .ZN(P1_U3236) );
  OAI211_X1 U10250 ( .C1(n8897), .C2(n8900), .A(n8899), .B(n8898), .ZN(n8909)
         );
  NAND2_X1 U10251 ( .A1(n9147), .A2(n8901), .ZN(n8902) );
  OAI21_X1 U10252 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8903), .A(n8902), .ZN(
        n8906) );
  NOR2_X1 U10253 ( .A1(n9113), .A2(n8904), .ZN(n8905) );
  AOI211_X1 U10254 ( .C1(n9117), .C2(n8907), .A(n8906), .B(n8905), .ZN(n8908)
         );
  OAI211_X1 U10255 ( .C1(n9120), .C2(n8910), .A(n8909), .B(n8908), .ZN(
        P1_U3238) );
  NAND2_X1 U10256 ( .A1(n8911), .A2(n8912), .ZN(n8913) );
  XOR2_X1 U10257 ( .A(n8914), .B(n8913), .Z(n8924) );
  OAI21_X1 U10258 ( .B1(n8916), .B2(n9286), .A(n8915), .ZN(n8917) );
  AOI21_X1 U10259 ( .B1(n8918), .B2(n9014), .A(n8917), .ZN(n8919) );
  OAI21_X1 U10260 ( .B1(n8920), .B2(n9280), .A(n8919), .ZN(n8921) );
  AOI21_X1 U10261 ( .B1(n9371), .B2(n8894), .A(n8921), .ZN(n8922) );
  OAI21_X1 U10262 ( .B1(n8924), .B2(n8923), .A(n8922), .ZN(P1_U3239) );
  MUX2_X1 U10263 ( .A(n9002), .B(P1_DATAO_REG_31__SCAN_IN), .S(n8936), .Z(
        P1_U3586) );
  MUX2_X1 U10264 ( .A(n8925), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8936), .Z(
        P1_U3585) );
  MUX2_X1 U10265 ( .A(n9038), .B(P1_DATAO_REG_28__SCAN_IN), .S(n8936), .Z(
        P1_U3583) );
  MUX2_X1 U10266 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8926), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10267 ( .A(n8927), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8936), .Z(
        P1_U3581) );
  MUX2_X1 U10268 ( .A(n9147), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8936), .Z(
        P1_U3580) );
  MUX2_X1 U10269 ( .A(n9164), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8936), .Z(
        P1_U3579) );
  MUX2_X1 U10270 ( .A(n9146), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8936), .Z(
        P1_U3578) );
  MUX2_X1 U10271 ( .A(n9158), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8936), .Z(
        P1_U3577) );
  MUX2_X1 U10272 ( .A(n9022), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8936), .Z(
        P1_U3576) );
  MUX2_X1 U10273 ( .A(n9020), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8936), .Z(
        P1_U3575) );
  MUX2_X1 U10274 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9018), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10275 ( .A(n9017), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8936), .Z(
        P1_U3573) );
  MUX2_X1 U10276 ( .A(n9015), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8936), .Z(
        P1_U3572) );
  MUX2_X1 U10277 ( .A(n9014), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8936), .Z(
        P1_U3571) );
  MUX2_X1 U10278 ( .A(n9453), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8936), .Z(
        P1_U3570) );
  MUX2_X1 U10279 ( .A(n9436), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8936), .Z(
        P1_U3569) );
  MUX2_X1 U10280 ( .A(n9454), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8936), .Z(
        P1_U3568) );
  MUX2_X1 U10281 ( .A(n9435), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8936), .Z(
        P1_U3567) );
  MUX2_X1 U10282 ( .A(n8928), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8936), .Z(
        P1_U3566) );
  MUX2_X1 U10283 ( .A(n8929), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8936), .Z(
        P1_U3565) );
  MUX2_X1 U10284 ( .A(n8930), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8936), .Z(
        P1_U3564) );
  MUX2_X1 U10285 ( .A(n8931), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8936), .Z(
        P1_U3563) );
  MUX2_X1 U10286 ( .A(n8932), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8936), .Z(
        P1_U3562) );
  MUX2_X1 U10287 ( .A(n8933), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8936), .Z(
        P1_U3561) );
  MUX2_X1 U10288 ( .A(n8934), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8936), .Z(
        P1_U3560) );
  MUX2_X1 U10289 ( .A(n9627), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8936), .Z(
        P1_U3559) );
  MUX2_X1 U10290 ( .A(n8935), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8936), .Z(
        P1_U3558) );
  MUX2_X1 U10291 ( .A(n9629), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8936), .Z(
        P1_U3557) );
  MUX2_X1 U10292 ( .A(n6241), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8936), .Z(
        P1_U3556) );
  MUX2_X1 U10293 ( .A(n8937), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8936), .Z(
        P1_U3555) );
  NOR2_X1 U10294 ( .A1(n9613), .A2(n8938), .ZN(n8939) );
  AOI211_X1 U10295 ( .C1(n9619), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n8940), .B(
        n8939), .ZN(n8951) );
  OAI21_X1 U10296 ( .B1(n8943), .B2(n8942), .A(n8941), .ZN(n8944) );
  NAND2_X1 U10297 ( .A1(n8944), .A2(n9620), .ZN(n8950) );
  OAI21_X1 U10298 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  NAND2_X1 U10299 ( .A1(n8948), .A2(n9609), .ZN(n8949) );
  NAND3_X1 U10300 ( .A1(n8951), .A2(n8950), .A3(n8949), .ZN(P1_U3248) );
  NOR2_X1 U10301 ( .A1(n8952), .A2(n8958), .ZN(n8954) );
  INV_X1 U10302 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8955) );
  MUX2_X1 U10303 ( .A(n8955), .B(P1_REG2_REG_16__SCAN_IN), .S(n8975), .Z(n8956) );
  AOI211_X1 U10304 ( .C1(n4344), .C2(n8956), .A(n8969), .B(n9578), .ZN(n8968)
         );
  NOR2_X1 U10305 ( .A1(n8958), .A2(n8957), .ZN(n8960) );
  XNOR2_X1 U10306 ( .A(n8975), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8961) );
  NOR2_X1 U10307 ( .A1(n8962), .A2(n8961), .ZN(n8974) );
  AOI211_X1 U10308 ( .C1(n8962), .C2(n8961), .A(n8974), .B(n9536), .ZN(n8967)
         );
  NAND2_X1 U10309 ( .A1(n9619), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U10310 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n8963) );
  OAI211_X1 U10311 ( .C1(n9613), .C2(n8965), .A(n8964), .B(n8963), .ZN(n8966)
         );
  OR3_X1 U10312 ( .A1(n8968), .A2(n8967), .A3(n8966), .ZN(P1_U3257) );
  AOI21_X1 U10313 ( .B1(n8975), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8969), .ZN(
        n8972) );
  NAND2_X1 U10314 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8987), .ZN(n8970) );
  OAI21_X1 U10315 ( .B1(n8987), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8970), .ZN(
        n8971) );
  NOR2_X1 U10316 ( .A1(n8972), .A2(n8971), .ZN(n8982) );
  AOI211_X1 U10317 ( .C1(n8972), .C2(n8971), .A(n8982), .B(n9578), .ZN(n8973)
         );
  AOI21_X1 U10318 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n9619), .A(n8973), .ZN(
        n8981) );
  AND2_X1 U10319 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8979) );
  XNOR2_X1 U10320 ( .A(n8987), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8976) );
  NOR2_X1 U10321 ( .A1(n8977), .A2(n8976), .ZN(n8986) );
  AOI211_X1 U10322 ( .C1(n8977), .C2(n8976), .A(n8986), .B(n9536), .ZN(n8978)
         );
  AOI211_X1 U10323 ( .C1(n9593), .C2(n8987), .A(n8979), .B(n8978), .ZN(n8980)
         );
  NAND2_X1 U10324 ( .A1(n8981), .A2(n8980), .ZN(P1_U3258) );
  OR2_X1 U10325 ( .A1(n8988), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U10326 ( .A1(n8988), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U10327 ( .A1(n8984), .A2(n8983), .ZN(n9608) );
  INV_X1 U10328 ( .A(n8993), .ZN(n8991) );
  INV_X1 U10329 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8985) );
  AOI22_X1 U10330 ( .A1(n8988), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8985), .B2(
        n9614), .ZN(n9618) );
  AOI21_X1 U10331 ( .B1(n8987), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8986), .ZN(
        n9617) );
  NAND2_X1 U10332 ( .A1(n9618), .A2(n9617), .ZN(n9616) );
  OAI21_X1 U10333 ( .B1(n8992), .B2(n9536), .A(n9613), .ZN(n8990) );
  AOI21_X1 U10334 ( .B1(n8991), .B2(n9609), .A(n8990), .ZN(n8996) );
  AOI22_X1 U10335 ( .A1(n8993), .A2(n9609), .B1(n9620), .B2(n8992), .ZN(n8995)
         );
  MUX2_X1 U10336 ( .A(n8996), .B(n8995), .S(n8994), .Z(n8998) );
  NAND2_X1 U10337 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n8997) );
  OAI211_X1 U10338 ( .C1(n4812), .C2(n9605), .A(n8998), .B(n8997), .ZN(
        P1_U3260) );
  INV_X1 U10339 ( .A(n9442), .ZN(n9465) );
  NAND2_X1 U10340 ( .A1(n9443), .A2(n9465), .ZN(n9459) );
  INV_X1 U10341 ( .A(n9365), .ZN(n9272) );
  INV_X1 U10342 ( .A(n9354), .ZN(n9232) );
  INV_X1 U10343 ( .A(n9344), .ZN(n9212) );
  NAND2_X1 U10344 ( .A1(n9220), .A2(n9212), .ZN(n9205) );
  NOR2_X2 U10345 ( .A1(n9137), .A2(n9319), .ZN(n9129) );
  NAND2_X1 U10346 ( .A1(n9297), .A2(n9073), .ZN(n9005) );
  XNOR2_X1 U10347 ( .A(n9294), .B(n9005), .ZN(n8999) );
  NAND2_X1 U10348 ( .A1(n8999), .A2(n9640), .ZN(n9293) );
  INV_X1 U10349 ( .A(P1_B_REG_SCAN_IN), .ZN(n9000) );
  NOR2_X1 U10350 ( .A1(n4278), .A2(n9000), .ZN(n9069) );
  INV_X1 U10351 ( .A(n9069), .ZN(n9001) );
  NAND3_X1 U10352 ( .A1(n9628), .A2(n9002), .A3(n9001), .ZN(n9295) );
  NOR2_X1 U10353 ( .A1(n9648), .A2(n9295), .ZN(n9007) );
  NOR2_X1 U10354 ( .A1(n9294), .A2(n9638), .ZN(n9003) );
  AOI211_X1 U10355 ( .C1(n9648), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9007), .B(
        n9003), .ZN(n9004) );
  OAI21_X1 U10356 ( .B1(n9293), .B2(n10037), .A(n9004), .ZN(P1_U3261) );
  OAI211_X1 U10357 ( .C1(n9297), .C2(n9073), .A(n9640), .B(n9005), .ZN(n9296)
         );
  NOR2_X1 U10358 ( .A1(n9297), .A2(n9638), .ZN(n9006) );
  AOI211_X1 U10359 ( .C1(n9648), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9007), .B(
        n9006), .ZN(n9008) );
  OAI21_X1 U10360 ( .B1(n10037), .B2(n9296), .A(n9008), .ZN(P1_U3262) );
  INV_X1 U10361 ( .A(n9371), .ZN(n9279) );
  NOR2_X1 U10362 ( .A1(n9279), .A2(n9262), .ZN(n9013) );
  NOR2_X1 U10363 ( .A1(n9359), .A2(n9015), .ZN(n9016) );
  INV_X1 U10364 ( .A(n9359), .ZN(n9246) );
  NOR2_X1 U10365 ( .A1(n9349), .A2(n9018), .ZN(n9019) );
  INV_X1 U10366 ( .A(n9349), .ZN(n9225) );
  NOR2_X1 U10367 ( .A1(n9212), .A2(n9219), .ZN(n9021) );
  NAND2_X1 U10368 ( .A1(n9181), .A2(n9189), .ZN(n9024) );
  NOR2_X1 U10369 ( .A1(n9328), .A2(n9146), .ZN(n9027) );
  NAND2_X1 U10370 ( .A1(n9328), .A2(n9146), .ZN(n9026) );
  NOR2_X1 U10371 ( .A1(n9142), .A2(n9127), .ZN(n9028) );
  NAND2_X1 U10372 ( .A1(n9030), .A2(n9029), .ZN(n9108) );
  NAND2_X1 U10373 ( .A1(n9108), .A2(n9031), .ZN(n9033) );
  NAND2_X1 U10374 ( .A1(n9120), .A2(n9128), .ZN(n9032) );
  NAND2_X1 U10375 ( .A1(n9033), .A2(n9032), .ZN(n9095) );
  NAND2_X1 U10376 ( .A1(n9095), .A2(n9097), .ZN(n9036) );
  NAND2_X1 U10377 ( .A1(n9034), .A2(n9113), .ZN(n9035) );
  INV_X1 U10378 ( .A(n9082), .ZN(n9037) );
  INV_X1 U10379 ( .A(n9298), .ZN(n9080) );
  INV_X1 U10380 ( .A(n9043), .ZN(n9449) );
  INV_X1 U10381 ( .A(n9044), .ZN(n9045) );
  NOR2_X1 U10382 ( .A1(n9239), .A2(n9238), .ZN(n9237) );
  INV_X1 U10383 ( .A(n9051), .ZN(n9052) );
  NOR2_X1 U10384 ( .A1(n9237), .A2(n9052), .ZN(n9217) );
  INV_X1 U10385 ( .A(n9055), .ZN(n9187) );
  INV_X1 U10386 ( .A(n9059), .ZN(n9060) );
  INV_X1 U10387 ( .A(n9066), .ZN(n9067) );
  NOR3_X1 U10388 ( .A1(n9070), .A2(n9069), .A3(n9289), .ZN(n9071) );
  AOI21_X1 U10389 ( .B1(n9038), .B2(n9630), .A(n9071), .ZN(n9072) );
  AOI211_X1 U10390 ( .C1(n9301), .C2(n9086), .A(n9458), .B(n9073), .ZN(n9300)
         );
  NAND2_X1 U10391 ( .A1(n9300), .A2(n9644), .ZN(n9077) );
  INV_X1 U10392 ( .A(n9074), .ZN(n9075) );
  AOI22_X1 U10393 ( .A1(n9075), .A2(n10031), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n9648), .ZN(n9076) );
  OAI211_X1 U10394 ( .C1(n4495), .C2(n9638), .A(n9077), .B(n9076), .ZN(n9078)
         );
  AOI21_X1 U10395 ( .B1(n9299), .B2(n10029), .A(n9078), .ZN(n9079) );
  OAI21_X1 U10396 ( .B1(n9080), .B2(n9292), .A(n9079), .ZN(P1_U3355) );
  XNOR2_X1 U10397 ( .A(n9083), .B(n9082), .ZN(n9084) );
  INV_X1 U10398 ( .A(n9101), .ZN(n9088) );
  INV_X1 U10399 ( .A(n9086), .ZN(n9087) );
  AOI211_X1 U10400 ( .C1(n9306), .C2(n9088), .A(n9458), .B(n9087), .ZN(n9305)
         );
  NAND2_X1 U10401 ( .A1(n9305), .A2(n9644), .ZN(n9091) );
  AOI22_X1 U10402 ( .A1(n9089), .A2(n10031), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n9648), .ZN(n9090) );
  OAI211_X1 U10403 ( .C1(n9092), .C2(n9638), .A(n9091), .B(n9090), .ZN(n9093)
         );
  AOI21_X1 U10404 ( .B1(n9304), .B2(n10029), .A(n9093), .ZN(n9094) );
  OAI21_X1 U10405 ( .B1(n9307), .B2(n9292), .A(n9094), .ZN(P1_U3263) );
  XNOR2_X1 U10406 ( .A(n9095), .B(n9096), .ZN(n9311) );
  AOI22_X1 U10407 ( .A1(n9310), .A2(n10033), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9648), .ZN(n9107) );
  XNOR2_X1 U10408 ( .A(n9098), .B(n9097), .ZN(n9099) );
  AOI211_X1 U10409 ( .C1(n9310), .C2(n9114), .A(n9458), .B(n9101), .ZN(n9309)
         );
  INV_X1 U10410 ( .A(n9309), .ZN(n9104) );
  INV_X1 U10411 ( .A(n9102), .ZN(n9103) );
  OAI22_X1 U10412 ( .A1(n9104), .A2(n9193), .B1(n9635), .B2(n9103), .ZN(n9105)
         );
  OAI21_X1 U10413 ( .B1(n9308), .B2(n9105), .A(n10029), .ZN(n9106) );
  OAI211_X1 U10414 ( .C1(n9311), .C2(n9292), .A(n9107), .B(n9106), .ZN(
        P1_U3264) );
  XNOR2_X1 U10415 ( .A(n9108), .B(n9109), .ZN(n9316) );
  XNOR2_X1 U10416 ( .A(n9110), .B(n9109), .ZN(n9111) );
  OAI222_X1 U10417 ( .A1(n9289), .A2(n9113), .B1(n9287), .B2(n9112), .C1(n9111), .C2(n9632), .ZN(n9312) );
  INV_X1 U10418 ( .A(n9129), .ZN(n9116) );
  INV_X1 U10419 ( .A(n9114), .ZN(n9115) );
  AOI211_X1 U10420 ( .C1(n9314), .C2(n9116), .A(n9458), .B(n9115), .ZN(n9313)
         );
  NAND2_X1 U10421 ( .A1(n9313), .A2(n9644), .ZN(n9119) );
  AOI22_X1 U10422 ( .A1(n9117), .A2(n10031), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9648), .ZN(n9118) );
  OAI211_X1 U10423 ( .C1(n9120), .C2(n9638), .A(n9119), .B(n9118), .ZN(n9121)
         );
  AOI21_X1 U10424 ( .B1(n9312), .B2(n10029), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10425 ( .B1(n9316), .B2(n9292), .A(n9122), .ZN(P1_U3265) );
  XOR2_X1 U10426 ( .A(n9124), .B(n9123), .Z(n9321) );
  AOI22_X1 U10427 ( .A1(n9319), .A2(n10033), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9648), .ZN(n9134) );
  XNOR2_X1 U10428 ( .A(n9125), .B(n9124), .ZN(n9126) );
  OAI222_X1 U10429 ( .A1(n9289), .A2(n9128), .B1(n9287), .B2(n9127), .C1(n9126), .C2(n9632), .ZN(n9317) );
  AOI211_X1 U10430 ( .C1(n9319), .C2(n9137), .A(n9458), .B(n9129), .ZN(n9318)
         );
  INV_X1 U10431 ( .A(n9318), .ZN(n9131) );
  OAI22_X1 U10432 ( .A1(n9131), .A2(n9193), .B1(n9635), .B2(n9130), .ZN(n9132)
         );
  OAI21_X1 U10433 ( .B1(n9317), .B2(n9132), .A(n10029), .ZN(n9133) );
  OAI211_X1 U10434 ( .C1(n9321), .C2(n9292), .A(n9134), .B(n9133), .ZN(
        P1_U3266) );
  XNOR2_X1 U10435 ( .A(n9136), .B(n9135), .ZN(n9326) );
  INV_X1 U10436 ( .A(n9153), .ZN(n9139) );
  INV_X1 U10437 ( .A(n9137), .ZN(n9138) );
  AOI211_X1 U10438 ( .C1(n9323), .C2(n9139), .A(n9458), .B(n9138), .ZN(n9322)
         );
  AOI22_X1 U10439 ( .A1(n9140), .A2(n10031), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9648), .ZN(n9141) );
  OAI21_X1 U10440 ( .B1(n9142), .B2(n9638), .A(n9141), .ZN(n9150) );
  OAI21_X1 U10441 ( .B1(n9145), .B2(n9144), .A(n9143), .ZN(n9148) );
  AOI222_X1 U10442 ( .A1(n9451), .A2(n9148), .B1(n9147), .B2(n9628), .C1(n9146), .C2(n9630), .ZN(n9325) );
  NOR2_X1 U10443 ( .A1(n9325), .A2(n9648), .ZN(n9149) );
  AOI211_X1 U10444 ( .C1(n9322), .C2(n9644), .A(n9150), .B(n9149), .ZN(n9151)
         );
  OAI21_X1 U10445 ( .B1(n9326), .B2(n9292), .A(n9151), .ZN(P1_U3267) );
  XNOR2_X1 U10446 ( .A(n9152), .B(n4806), .ZN(n9331) );
  AOI211_X1 U10447 ( .C1(n9328), .C2(n9174), .A(n9458), .B(n9153), .ZN(n9327)
         );
  INV_X1 U10448 ( .A(n9154), .ZN(n9155) );
  AOI22_X1 U10449 ( .A1(n9155), .A2(n10031), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9648), .ZN(n9156) );
  OAI21_X1 U10450 ( .B1(n9157), .B2(n9638), .A(n9156), .ZN(n9166) );
  AND2_X1 U10451 ( .A1(n9158), .A2(n9630), .ZN(n9163) );
  AOI211_X1 U10452 ( .C1(n9161), .C2(n9160), .A(n9632), .B(n9159), .ZN(n9162)
         );
  AOI211_X1 U10453 ( .C1(n9628), .C2(n9164), .A(n9163), .B(n9162), .ZN(n9330)
         );
  NOR2_X1 U10454 ( .A1(n9330), .A2(n9648), .ZN(n9165) );
  AOI211_X1 U10455 ( .C1(n9327), .C2(n9644), .A(n9166), .B(n9165), .ZN(n9167)
         );
  OAI21_X1 U10456 ( .B1(n9331), .B2(n9292), .A(n9167), .ZN(P1_U3268) );
  XNOR2_X1 U10457 ( .A(n9168), .B(n9169), .ZN(n9336) );
  XNOR2_X1 U10458 ( .A(n9171), .B(n9170), .ZN(n9172) );
  OAI222_X1 U10459 ( .A1(n9289), .A2(n9173), .B1(n9287), .B2(n9204), .C1(n9172), .C2(n9632), .ZN(n9332) );
  INV_X1 U10460 ( .A(n9190), .ZN(n9176) );
  INV_X1 U10461 ( .A(n9174), .ZN(n9175) );
  AOI211_X1 U10462 ( .C1(n9334), .C2(n9176), .A(n9458), .B(n9175), .ZN(n9333)
         );
  NAND2_X1 U10463 ( .A1(n9333), .A2(n9644), .ZN(n9180) );
  INV_X1 U10464 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U10465 ( .A1(n9178), .A2(n10031), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9648), .ZN(n9179) );
  OAI211_X1 U10466 ( .C1(n9181), .C2(n9638), .A(n9180), .B(n9179), .ZN(n9182)
         );
  AOI21_X1 U10467 ( .B1(n9332), .B2(n10029), .A(n9182), .ZN(n9183) );
  OAI21_X1 U10468 ( .B1(n9336), .B2(n9292), .A(n9183), .ZN(P1_U3269) );
  OAI21_X1 U10469 ( .B1(n4312), .B2(n9187), .A(n9184), .ZN(n9341) );
  AOI22_X1 U10470 ( .A1(n9339), .A2(n10033), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n9648), .ZN(n9197) );
  AOI21_X1 U10471 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9188) );
  OAI222_X1 U10472 ( .A1(n9289), .A2(n9189), .B1(n9287), .B2(n9219), .C1(n9632), .C2(n9188), .ZN(n9337) );
  AOI211_X1 U10473 ( .C1(n9339), .C2(n9205), .A(n9458), .B(n9190), .ZN(n9338)
         );
  INV_X1 U10474 ( .A(n9338), .ZN(n9194) );
  INV_X1 U10475 ( .A(n9191), .ZN(n9192) );
  OAI22_X1 U10476 ( .A1(n9194), .A2(n9193), .B1(n9635), .B2(n9192), .ZN(n9195)
         );
  OAI21_X1 U10477 ( .B1(n9337), .B2(n9195), .A(n10029), .ZN(n9196) );
  OAI211_X1 U10478 ( .C1(n9341), .C2(n9292), .A(n9197), .B(n9196), .ZN(
        P1_U3270) );
  XNOR2_X1 U10479 ( .A(n9198), .B(n9202), .ZN(n9346) );
  INV_X1 U10480 ( .A(n9199), .ZN(n9200) );
  NOR2_X1 U10481 ( .A1(n4494), .A2(n9200), .ZN(n9201) );
  XOR2_X1 U10482 ( .A(n9202), .B(n9201), .Z(n9203) );
  OAI222_X1 U10483 ( .A1(n9289), .A2(n9204), .B1(n9287), .B2(n9241), .C1(n9203), .C2(n9632), .ZN(n9342) );
  INV_X1 U10484 ( .A(n9220), .ZN(n9207) );
  INV_X1 U10485 ( .A(n9205), .ZN(n9206) );
  AOI211_X1 U10486 ( .C1(n9344), .C2(n9207), .A(n9458), .B(n9206), .ZN(n9343)
         );
  NAND2_X1 U10487 ( .A1(n9343), .A2(n9644), .ZN(n9211) );
  INV_X1 U10488 ( .A(n9208), .ZN(n9209) );
  AOI22_X1 U10489 ( .A1(n9648), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9209), .B2(
        n10031), .ZN(n9210) );
  OAI211_X1 U10490 ( .C1(n9212), .C2(n9638), .A(n9211), .B(n9210), .ZN(n9213)
         );
  AOI21_X1 U10491 ( .B1(n9342), .B2(n10029), .A(n9213), .ZN(n9214) );
  OAI21_X1 U10492 ( .B1(n9346), .B2(n9292), .A(n9214), .ZN(P1_U3271) );
  XOR2_X1 U10493 ( .A(n9216), .B(n9215), .Z(n9351) );
  AOI21_X1 U10494 ( .B1(n9217), .B2(n9216), .A(n4494), .ZN(n9218) );
  OAI222_X1 U10495 ( .A1(n9289), .A2(n9219), .B1(n9287), .B2(n9254), .C1(n9632), .C2(n9218), .ZN(n9347) );
  AOI211_X1 U10496 ( .C1(n9349), .C2(n9229), .A(n9458), .B(n9220), .ZN(n9348)
         );
  NAND2_X1 U10497 ( .A1(n9348), .A2(n9644), .ZN(n9224) );
  INV_X1 U10498 ( .A(n9221), .ZN(n9222) );
  AOI22_X1 U10499 ( .A1(n9648), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9222), .B2(
        n10031), .ZN(n9223) );
  OAI211_X1 U10500 ( .C1(n9225), .C2(n9638), .A(n9224), .B(n9223), .ZN(n9226)
         );
  AOI21_X1 U10501 ( .B1(n9347), .B2(n10029), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10502 ( .B1(n9351), .B2(n9292), .A(n9227), .ZN(P1_U3272) );
  XNOR2_X1 U10503 ( .A(n9228), .B(n9238), .ZN(n9356) );
  INV_X1 U10504 ( .A(n9245), .ZN(n9231) );
  INV_X1 U10505 ( .A(n9229), .ZN(n9230) );
  AOI211_X1 U10506 ( .C1(n9354), .C2(n9231), .A(n9458), .B(n9230), .ZN(n9353)
         );
  NOR2_X1 U10507 ( .A1(n9232), .A2(n9638), .ZN(n9236) );
  OAI22_X1 U10508 ( .A1(n10029), .A2(n9234), .B1(n9233), .B2(n9635), .ZN(n9235) );
  AOI211_X1 U10509 ( .C1(n9353), .C2(n9644), .A(n9236), .B(n9235), .ZN(n9243)
         );
  AOI21_X1 U10510 ( .B1(n9239), .B2(n9238), .A(n9237), .ZN(n9240) );
  OAI222_X1 U10511 ( .A1(n9289), .A2(n9241), .B1(n9287), .B2(n9263), .C1(n9632), .C2(n9240), .ZN(n9352) );
  NAND2_X1 U10512 ( .A1(n9352), .A2(n10029), .ZN(n9242) );
  OAI211_X1 U10513 ( .C1(n9356), .C2(n9292), .A(n9243), .B(n9242), .ZN(
        P1_U3273) );
  XNOR2_X1 U10514 ( .A(n9244), .B(n9252), .ZN(n9361) );
  AOI211_X1 U10515 ( .C1(n9359), .C2(n9267), .A(n9458), .B(n9245), .ZN(n9358)
         );
  NOR2_X1 U10516 ( .A1(n9246), .A2(n9638), .ZN(n9250) );
  INV_X1 U10517 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9248) );
  OAI22_X1 U10518 ( .A1(n10029), .A2(n9248), .B1(n9247), .B2(n9635), .ZN(n9249) );
  AOI211_X1 U10519 ( .C1(n9358), .C2(n9644), .A(n9250), .B(n9249), .ZN(n9256)
         );
  XOR2_X1 U10520 ( .A(n9252), .B(n9251), .Z(n9253) );
  OAI222_X1 U10521 ( .A1(n9289), .A2(n9254), .B1(n9287), .B2(n9288), .C1(n9253), .C2(n9632), .ZN(n9357) );
  NAND2_X1 U10522 ( .A1(n9357), .A2(n10029), .ZN(n9255) );
  OAI211_X1 U10523 ( .C1(n9361), .C2(n9292), .A(n9256), .B(n9255), .ZN(
        P1_U3274) );
  INV_X1 U10524 ( .A(n9257), .ZN(n9258) );
  NOR2_X1 U10525 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  XOR2_X1 U10526 ( .A(n9264), .B(n9260), .Z(n9261) );
  OAI222_X1 U10527 ( .A1(n9289), .A2(n9263), .B1(n9287), .B2(n9262), .C1(n9632), .C2(n9261), .ZN(n9363) );
  INV_X1 U10528 ( .A(n9363), .ZN(n9276) );
  INV_X1 U10529 ( .A(n9368), .ZN(n9266) );
  NAND2_X1 U10530 ( .A1(n9265), .A2(n9264), .ZN(n9362) );
  NAND3_X1 U10531 ( .A1(n9266), .A2(n10041), .A3(n9362), .ZN(n9275) );
  INV_X1 U10532 ( .A(n9278), .ZN(n9269) );
  INV_X1 U10533 ( .A(n9267), .ZN(n9268) );
  AOI211_X1 U10534 ( .C1(n9365), .C2(n9269), .A(n9458), .B(n9268), .ZN(n9364)
         );
  AOI22_X1 U10535 ( .A1(n9648), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9270), .B2(
        n10031), .ZN(n9271) );
  OAI21_X1 U10536 ( .B1(n9272), .B2(n9638), .A(n9271), .ZN(n9273) );
  AOI21_X1 U10537 ( .B1(n9364), .B2(n9644), .A(n9273), .ZN(n9274) );
  OAI211_X1 U10538 ( .C1(n9648), .C2(n9276), .A(n9275), .B(n9274), .ZN(
        P1_U3275) );
  XOR2_X1 U10539 ( .A(n9277), .B(n9284), .Z(n9374) );
  AOI211_X1 U10540 ( .C1(n9371), .C2(n9460), .A(n9458), .B(n9278), .ZN(n9370)
         );
  NOR2_X1 U10541 ( .A1(n9279), .A2(n9638), .ZN(n9282) );
  OAI22_X1 U10542 ( .A1(n10029), .A2(n9975), .B1(n9280), .B2(n9635), .ZN(n9281) );
  AOI211_X1 U10543 ( .C1(n9370), .C2(n9644), .A(n9282), .B(n9281), .ZN(n9291)
         );
  XOR2_X1 U10544 ( .A(n9284), .B(n9283), .Z(n9285) );
  OAI222_X1 U10545 ( .A1(n9289), .A2(n9288), .B1(n9287), .B2(n9286), .C1(n9632), .C2(n9285), .ZN(n9369) );
  NAND2_X1 U10546 ( .A1(n9369), .A2(n10029), .ZN(n9290) );
  OAI211_X1 U10547 ( .C1(n9374), .C2(n9292), .A(n9291), .B(n9290), .ZN(
        P1_U3276) );
  OAI211_X1 U10548 ( .C1(n9294), .C2(n9701), .A(n9293), .B(n9295), .ZN(n9376)
         );
  MUX2_X1 U10549 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9376), .S(n9721), .Z(
        P1_U3554) );
  OAI211_X1 U10550 ( .C1(n9297), .C2(n9701), .A(n9296), .B(n9295), .ZN(n9377)
         );
  MUX2_X1 U10551 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9377), .S(n9721), .Z(
        P1_U3553) );
  NAND2_X1 U10552 ( .A1(n9298), .A2(n9705), .ZN(n9303) );
  NAND2_X1 U10553 ( .A1(n9303), .A2(n9302), .ZN(n9378) );
  MUX2_X1 U10554 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9378), .S(n9721), .Z(
        P1_U3552) );
  MUX2_X1 U10555 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9380), .S(n9721), .Z(
        P1_U3550) );
  AOI211_X1 U10556 ( .C1(n9679), .C2(n9314), .A(n9313), .B(n9312), .ZN(n9315)
         );
  OAI21_X1 U10557 ( .B1(n9316), .B2(n9373), .A(n9315), .ZN(n9381) );
  MUX2_X1 U10558 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9381), .S(n9721), .Z(
        P1_U3549) );
  AOI211_X1 U10559 ( .C1(n9679), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9320)
         );
  OAI21_X1 U10560 ( .B1(n9321), .B2(n9373), .A(n9320), .ZN(n9382) );
  MUX2_X1 U10561 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9382), .S(n9721), .Z(
        P1_U3548) );
  AOI21_X1 U10562 ( .B1(n9679), .B2(n9323), .A(n9322), .ZN(n9324) );
  OAI211_X1 U10563 ( .C1(n9326), .C2(n9373), .A(n9325), .B(n9324), .ZN(n9383)
         );
  MUX2_X1 U10564 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9383), .S(n9721), .Z(
        P1_U3547) );
  AOI21_X1 U10565 ( .B1(n9679), .B2(n9328), .A(n9327), .ZN(n9329) );
  OAI211_X1 U10566 ( .C1(n9331), .C2(n9373), .A(n9330), .B(n9329), .ZN(n9384)
         );
  MUX2_X1 U10567 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9384), .S(n9721), .Z(
        P1_U3546) );
  AOI211_X1 U10568 ( .C1(n9679), .C2(n9334), .A(n9333), .B(n9332), .ZN(n9335)
         );
  OAI21_X1 U10569 ( .B1(n9336), .B2(n9373), .A(n9335), .ZN(n9385) );
  MUX2_X1 U10570 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9385), .S(n9721), .Z(
        P1_U3545) );
  AOI211_X1 U10571 ( .C1(n9679), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  OAI21_X1 U10572 ( .B1(n9341), .B2(n9373), .A(n9340), .ZN(n9386) );
  MUX2_X1 U10573 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9386), .S(n9721), .Z(
        P1_U3544) );
  AOI211_X1 U10574 ( .C1(n9679), .C2(n9344), .A(n9343), .B(n9342), .ZN(n9345)
         );
  OAI21_X1 U10575 ( .B1(n9346), .B2(n9373), .A(n9345), .ZN(n9387) );
  MUX2_X1 U10576 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9387), .S(n9721), .Z(
        P1_U3543) );
  AOI211_X1 U10577 ( .C1(n9679), .C2(n9349), .A(n9348), .B(n9347), .ZN(n9350)
         );
  OAI21_X1 U10578 ( .B1(n9351), .B2(n9373), .A(n9350), .ZN(n9388) );
  MUX2_X1 U10579 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9388), .S(n9721), .Z(
        P1_U3542) );
  AOI211_X1 U10580 ( .C1(n9679), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9355)
         );
  OAI21_X1 U10581 ( .B1(n9356), .B2(n9373), .A(n9355), .ZN(n9389) );
  MUX2_X1 U10582 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9389), .S(n9721), .Z(
        P1_U3541) );
  AOI211_X1 U10583 ( .C1(n9679), .C2(n9359), .A(n9358), .B(n9357), .ZN(n9360)
         );
  OAI21_X1 U10584 ( .B1(n9361), .B2(n9373), .A(n9360), .ZN(n9390) );
  MUX2_X1 U10585 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9390), .S(n9721), .Z(
        P1_U3540) );
  NAND2_X1 U10586 ( .A1(n9362), .A2(n9705), .ZN(n9367) );
  AOI211_X1 U10587 ( .C1(n9679), .C2(n9365), .A(n9364), .B(n9363), .ZN(n9366)
         );
  OAI21_X1 U10588 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9391) );
  MUX2_X1 U10589 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9391), .S(n9721), .Z(
        P1_U3539) );
  AOI211_X1 U10590 ( .C1(n9679), .C2(n9371), .A(n9370), .B(n9369), .ZN(n9372)
         );
  OAI21_X1 U10591 ( .B1(n9374), .B2(n9373), .A(n9372), .ZN(n9392) );
  MUX2_X1 U10592 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9392), .S(n9721), .Z(
        P1_U3538) );
  MUX2_X1 U10593 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9375), .S(n9721), .Z(
        P1_U3523) );
  MUX2_X1 U10594 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9376), .S(n9709), .Z(
        P1_U3522) );
  MUX2_X1 U10595 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9377), .S(n9709), .Z(
        P1_U3521) );
  MUX2_X1 U10596 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9378), .S(n9709), .Z(
        P1_U3520) );
  MUX2_X1 U10597 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9381), .S(n9709), .Z(
        P1_U3517) );
  MUX2_X1 U10598 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9382), .S(n9709), .Z(
        P1_U3516) );
  MUX2_X1 U10599 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9383), .S(n9709), .Z(
        P1_U3515) );
  MUX2_X1 U10600 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9384), .S(n9709), .Z(
        P1_U3514) );
  MUX2_X1 U10601 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9385), .S(n9709), .Z(
        P1_U3513) );
  MUX2_X1 U10602 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9386), .S(n9709), .Z(
        P1_U3512) );
  MUX2_X1 U10603 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9387), .S(n9709), .Z(
        P1_U3511) );
  MUX2_X1 U10604 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9388), .S(n9709), .Z(
        P1_U3510) );
  MUX2_X1 U10605 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9389), .S(n9709), .Z(
        P1_U3508) );
  MUX2_X1 U10606 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9390), .S(n9709), .Z(
        P1_U3505) );
  MUX2_X1 U10607 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9391), .S(n9709), .Z(
        P1_U3502) );
  MUX2_X1 U10608 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9392), .S(n9709), .Z(
        P1_U3499) );
  MUX2_X1 U10609 ( .A(n9394), .B(P1_D_REG_0__SCAN_IN), .S(n9393), .Z(P1_U3440)
         );
  INV_X1 U10610 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9395) );
  NAND3_X1 U10611 ( .A1(n9395), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9396) );
  OAI22_X1 U10612 ( .A1(n6094), .A2(n9396), .B1(n6039), .B2(n9404), .ZN(n9397)
         );
  AOI21_X1 U10613 ( .B1(n8772), .B2(n9398), .A(n9397), .ZN(n9399) );
  INV_X1 U10614 ( .A(n9399), .ZN(P1_U3322) );
  OAI222_X1 U10615 ( .A1(n9404), .A2(n9403), .B1(n9402), .B2(n9401), .C1(
        P1_U3084), .C2(n6098), .ZN(P1_U3323) );
  MUX2_X1 U10616 ( .A(n9405), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10617 ( .A1(n9417), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9416) );
  AOI211_X1 U10618 ( .C1(n9408), .C2(n9407), .A(n9406), .B(n9418), .ZN(n9409)
         );
  AOI21_X1 U10619 ( .B1(n9424), .B2(n9410), .A(n9409), .ZN(n9415) );
  INV_X1 U10620 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9735) );
  NOR2_X1 U10621 ( .A1(n9735), .A2(n5043), .ZN(n9413) );
  OAI211_X1 U10622 ( .C1(n9413), .C2(n9412), .A(n9722), .B(n9411), .ZN(n9414)
         );
  NAND3_X1 U10623 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(P2_U3246) );
  AOI22_X1 U10624 ( .A1(n9417), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9430) );
  AOI211_X1 U10625 ( .C1(n9421), .C2(n9420), .A(n9419), .B(n9418), .ZN(n9422)
         );
  AOI21_X1 U10626 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9429) );
  OAI211_X1 U10627 ( .C1(n9427), .C2(n9426), .A(n9722), .B(n9425), .ZN(n9428)
         );
  NAND3_X1 U10628 ( .A1(n9430), .A2(n9429), .A3(n9428), .ZN(P2_U3247) );
  OAI21_X1 U10629 ( .B1(n9432), .B2(n9434), .A(n9431), .ZN(n9469) );
  INV_X1 U10630 ( .A(n9656), .ZN(n9687) );
  AOI21_X1 U10631 ( .B1(n9434), .B2(n9433), .A(n9450), .ZN(n9438) );
  AOI22_X1 U10632 ( .A1(n9628), .A2(n9436), .B1(n9630), .B2(n9435), .ZN(n9437)
         );
  OAI21_X1 U10633 ( .B1(n9438), .B2(n9632), .A(n9437), .ZN(n9439) );
  AOI21_X1 U10634 ( .B1(n9469), .B2(n9687), .A(n9439), .ZN(n9466) );
  INV_X1 U10635 ( .A(n9440), .ZN(n9441) );
  AOI222_X1 U10636 ( .A1(n9442), .A2(n10033), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9648), .C1(n10031), .C2(n9441), .ZN(n9446) );
  OAI211_X1 U10637 ( .C1(n9443), .C2(n9465), .A(n9640), .B(n9459), .ZN(n9464)
         );
  INV_X1 U10638 ( .A(n9464), .ZN(n9444) );
  AOI22_X1 U10639 ( .A1(n9469), .A2(n9645), .B1(n9644), .B2(n9444), .ZN(n9445)
         );
  OAI211_X1 U10640 ( .C1(n9648), .C2(n9466), .A(n9446), .B(n9445), .ZN(
        P1_U3278) );
  XNOR2_X1 U10641 ( .A(n9447), .B(n9448), .ZN(n10042) );
  OAI21_X1 U10642 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(n9452) );
  NAND2_X1 U10643 ( .A1(n9452), .A2(n9451), .ZN(n9456) );
  AOI22_X1 U10644 ( .A1(n9630), .A2(n9454), .B1(n9628), .B2(n9453), .ZN(n9455)
         );
  OAI21_X1 U10645 ( .B1(n9457), .B2(n9456), .A(n9455), .ZN(n10030) );
  AOI21_X1 U10646 ( .B1(n9459), .B2(n10034), .A(n9458), .ZN(n9461) );
  NAND2_X1 U10647 ( .A1(n9461), .A2(n9460), .ZN(n10038) );
  OAI21_X1 U10648 ( .B1(n9462), .B2(n9701), .A(n10038), .ZN(n9463) );
  AOI211_X1 U10649 ( .C1(n10042), .C2(n9705), .A(n10030), .B(n9463), .ZN(n9484) );
  AOI22_X1 U10650 ( .A1(n9721), .A2(n9484), .B1(n7031), .B2(n9718), .ZN(
        P1_U3537) );
  INV_X1 U10651 ( .A(n9682), .ZN(n9699) );
  OAI21_X1 U10652 ( .B1(n9465), .B2(n9701), .A(n9464), .ZN(n9468) );
  INV_X1 U10653 ( .A(n9466), .ZN(n9467) );
  AOI211_X1 U10654 ( .C1(n9699), .C2(n9469), .A(n9468), .B(n9467), .ZN(n9485)
         );
  AOI22_X1 U10655 ( .A1(n9721), .A2(n9485), .B1(n7188), .B2(n9718), .ZN(
        P1_U3536) );
  AOI211_X1 U10656 ( .C1(n9679), .C2(n9472), .A(n9471), .B(n9470), .ZN(n9473)
         );
  OAI21_X1 U10657 ( .B1(n9474), .B2(n9682), .A(n9473), .ZN(n9475) );
  AOI21_X1 U10658 ( .B1(n9476), .B2(n9687), .A(n9475), .ZN(n9486) );
  AOI22_X1 U10659 ( .A1(n9721), .A2(n9486), .B1(n7005), .B2(n9718), .ZN(
        P1_U3535) );
  OAI211_X1 U10660 ( .C1(n9479), .C2(n9701), .A(n9478), .B(n9477), .ZN(n9480)
         );
  AOI21_X1 U10661 ( .B1(n9481), .B2(n9705), .A(n9480), .ZN(n9487) );
  AOI22_X1 U10662 ( .A1(n9721), .A2(n9487), .B1(n9482), .B2(n9718), .ZN(
        P1_U3534) );
  INV_X1 U10663 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9483) );
  AOI22_X1 U10664 ( .A1(n9709), .A2(n9484), .B1(n9483), .B2(n9707), .ZN(
        P1_U3496) );
  AOI22_X1 U10665 ( .A1(n9709), .A2(n9485), .B1(n7187), .B2(n9707), .ZN(
        P1_U3493) );
  AOI22_X1 U10666 ( .A1(n9709), .A2(n9486), .B1(n7003), .B2(n9707), .ZN(
        P1_U3490) );
  AOI22_X1 U10667 ( .A1(n9709), .A2(n9487), .B1(n6868), .B2(n9707), .ZN(
        P1_U3487) );
  XNOR2_X1 U10668 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10669 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U10670 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9490) );
  AOI211_X1 U10671 ( .C1(n9490), .C2(n9489), .A(n9488), .B(n9536), .ZN(n9494)
         );
  AOI211_X1 U10672 ( .C1(n9507), .C2(n9492), .A(n9491), .B(n9578), .ZN(n9493)
         );
  AOI211_X1 U10673 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9494), 
        .B(n9493), .ZN(n9499) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9495) );
  OAI22_X1 U10675 ( .A1(n9496), .A2(n9613), .B1(n9605), .B2(n9495), .ZN(n9497)
         );
  INV_X1 U10676 ( .A(n9497), .ZN(n9498) );
  NAND2_X1 U10677 ( .A1(n9499), .A2(n9498), .ZN(P1_U3242) );
  AOI211_X1 U10678 ( .C1(n9502), .C2(n9501), .A(n9500), .B(n9536), .ZN(n9503)
         );
  AOI21_X1 U10679 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9503), 
        .ZN(n9517) );
  AOI211_X1 U10680 ( .C1(n9506), .C2(n9505), .A(n9504), .B(n9578), .ZN(n9514)
         );
  INV_X1 U10681 ( .A(n9507), .ZN(n9510) );
  INV_X1 U10682 ( .A(n9508), .ZN(n9509) );
  MUX2_X1 U10683 ( .A(n9510), .B(n9509), .S(n4278), .Z(n9513) );
  AOI211_X1 U10684 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n8936), .ZN(n9527)
         );
  AOI211_X1 U10685 ( .C1(n9593), .C2(n9515), .A(n9514), .B(n9527), .ZN(n9516)
         );
  OAI211_X1 U10686 ( .C1(n9605), .C2(n9518), .A(n9517), .B(n9516), .ZN(
        P1_U3243) );
  OAI21_X1 U10687 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  AOI22_X1 U10688 ( .A1(n9593), .A2(n9523), .B1(n9609), .B2(n9522), .ZN(n9531)
         );
  OAI21_X1 U10689 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9529) );
  AOI211_X1 U10690 ( .C1(n9620), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9530)
         );
  OAI211_X1 U10691 ( .C1(n9605), .C2(n9532), .A(n9531), .B(n9530), .ZN(
        P1_U3245) );
  OAI21_X1 U10692 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9542) );
  AOI211_X1 U10693 ( .C1(n9539), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9540)
         );
  AOI211_X1 U10694 ( .C1(n9609), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9548)
         );
  INV_X1 U10695 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9545) );
  OR2_X1 U10696 ( .A1(n9613), .A2(n9543), .ZN(n9544) );
  OAI21_X1 U10697 ( .B1(n9605), .B2(n9545), .A(n9544), .ZN(n9546) );
  INV_X1 U10698 ( .A(n9546), .ZN(n9547) );
  NAND2_X1 U10699 ( .A1(n9548), .A2(n9547), .ZN(P1_U3246) );
  OAI21_X1 U10700 ( .B1(n9551), .B2(n9550), .A(n9549), .ZN(n9557) );
  AOI211_X1 U10701 ( .C1(n9554), .C2(n9553), .A(n9552), .B(n9578), .ZN(n9555)
         );
  AOI211_X1 U10702 ( .C1(n9620), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9562)
         );
  INV_X1 U10703 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9558) );
  OAI22_X1 U10704 ( .A1(n9559), .A2(n9613), .B1(n9605), .B2(n9558), .ZN(n9560)
         );
  INV_X1 U10705 ( .A(n9560), .ZN(n9561) );
  NAND2_X1 U10706 ( .A1(n9562), .A2(n9561), .ZN(P1_U3247) );
  OAI21_X1 U10707 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9571) );
  AOI211_X1 U10708 ( .C1(n9568), .C2(n9567), .A(n9566), .B(n9578), .ZN(n9569)
         );
  AOI211_X1 U10709 ( .C1(n9571), .C2(n9620), .A(n9570), .B(n9569), .ZN(n9574)
         );
  AOI22_X1 U10710 ( .A1(n9619), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9593), .B2(
        n9572), .ZN(n9573) );
  NAND2_X1 U10711 ( .A1(n9574), .A2(n9573), .ZN(P1_U3250) );
  OAI21_X1 U10712 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9584) );
  AOI211_X1 U10713 ( .C1(n9581), .C2(n9580), .A(n9579), .B(n9578), .ZN(n9582)
         );
  AOI211_X1 U10714 ( .C1(n9584), .C2(n9620), .A(n9583), .B(n9582), .ZN(n9590)
         );
  INV_X1 U10715 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9587) );
  OR2_X1 U10716 ( .A1(n9613), .A2(n9585), .ZN(n9586) );
  OAI21_X1 U10717 ( .B1(n9605), .B2(n9587), .A(n9586), .ZN(n9588) );
  INV_X1 U10718 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U10719 ( .A1(n9590), .A2(n9589), .ZN(P1_U3251) );
  INV_X1 U10720 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9604) );
  AOI21_X1 U10721 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9603) );
  OAI21_X1 U10722 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9601) );
  OAI21_X1 U10723 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9600) );
  AOI22_X1 U10724 ( .A1(n9601), .A2(n9620), .B1(n9600), .B2(n9609), .ZN(n9602)
         );
  OAI211_X1 U10725 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(
        P1_U3252) );
  AOI21_X1 U10726 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9610) );
  NAND2_X1 U10727 ( .A1(n9610), .A2(n9609), .ZN(n9612) );
  OAI211_X1 U10728 ( .C1(n9614), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9615)
         );
  INV_X1 U10729 ( .A(n9615), .ZN(n9623) );
  OAI21_X1 U10730 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9621) );
  AOI22_X1 U10731 ( .A1(n9621), .A2(n9620), .B1(n9619), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U10732 ( .A1(n9623), .A2(n9622), .ZN(P1_U3259) );
  XNOR2_X1 U10733 ( .A(n9626), .B(n9624), .ZN(n9664) );
  XNOR2_X1 U10734 ( .A(n9626), .B(n9625), .ZN(n9633) );
  AOI22_X1 U10735 ( .A1(n9630), .A2(n9629), .B1(n9628), .B2(n9627), .ZN(n9631)
         );
  OAI21_X1 U10736 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9634) );
  AOI21_X1 U10737 ( .B1(n9687), .B2(n9664), .A(n9634), .ZN(n9661) );
  NOR2_X1 U10738 ( .A1(n9635), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9636) );
  AOI21_X1 U10739 ( .B1(n9648), .B2(P1_REG2_REG_3__SCAN_IN), .A(n9636), .ZN(
        n9637) );
  OAI21_X1 U10740 ( .B1(n9638), .B2(n9660), .A(n9637), .ZN(n9639) );
  INV_X1 U10741 ( .A(n9639), .ZN(n9647) );
  OAI211_X1 U10742 ( .C1(n9660), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9659)
         );
  INV_X1 U10743 ( .A(n9659), .ZN(n9643) );
  AOI22_X1 U10744 ( .A1(n9664), .A2(n9645), .B1(n9644), .B2(n9643), .ZN(n9646)
         );
  OAI211_X1 U10745 ( .C1(n9648), .C2(n9661), .A(n9647), .B(n9646), .ZN(
        P1_U3288) );
  AND2_X1 U10746 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9650), .ZN(P1_U3292) );
  AND2_X1 U10747 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9650), .ZN(P1_U3293) );
  AND2_X1 U10748 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9650), .ZN(P1_U3294) );
  AND2_X1 U10749 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9650), .ZN(P1_U3295) );
  AND2_X1 U10750 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9650), .ZN(P1_U3296) );
  AND2_X1 U10751 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9650), .ZN(P1_U3297) );
  AND2_X1 U10752 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9650), .ZN(P1_U3298) );
  AND2_X1 U10753 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9650), .ZN(P1_U3299) );
  AND2_X1 U10754 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9650), .ZN(P1_U3300) );
  AND2_X1 U10755 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9650), .ZN(P1_U3301) );
  INV_X1 U10756 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U10757 ( .A1(n9649), .A2(n9940), .ZN(P1_U3302) );
  AND2_X1 U10758 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9650), .ZN(P1_U3303) );
  AND2_X1 U10759 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9650), .ZN(P1_U3304) );
  AND2_X1 U10760 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9650), .ZN(P1_U3305) );
  AND2_X1 U10761 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9650), .ZN(P1_U3306) );
  AND2_X1 U10762 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9650), .ZN(P1_U3307) );
  AND2_X1 U10763 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9650), .ZN(P1_U3308) );
  AND2_X1 U10764 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9650), .ZN(P1_U3309) );
  INV_X1 U10765 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U10766 ( .A1(n9649), .A2(n10013), .ZN(P1_U3310) );
  AND2_X1 U10767 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9650), .ZN(P1_U3311) );
  AND2_X1 U10768 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9650), .ZN(P1_U3312) );
  AND2_X1 U10769 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9650), .ZN(P1_U3313) );
  AND2_X1 U10770 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9650), .ZN(P1_U3314) );
  AND2_X1 U10771 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9650), .ZN(P1_U3315) );
  AND2_X1 U10772 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9650), .ZN(P1_U3316) );
  AND2_X1 U10773 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9650), .ZN(P1_U3317) );
  AND2_X1 U10774 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9650), .ZN(P1_U3318) );
  AND2_X1 U10775 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9650), .ZN(P1_U3319) );
  INV_X1 U10776 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U10777 ( .A1(n9649), .A2(n9956), .ZN(P1_U3320) );
  AND2_X1 U10778 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9650), .ZN(P1_U3321) );
  INV_X1 U10779 ( .A(n9651), .ZN(n9654) );
  OAI211_X1 U10780 ( .C1(n9654), .C2(n9701), .A(n9653), .B(n9652), .ZN(n9658)
         );
  AOI21_X1 U10781 ( .B1(n9656), .B2(n9682), .A(n9655), .ZN(n9657) );
  NOR2_X1 U10782 ( .A1(n9658), .A2(n9657), .ZN(n9710) );
  AOI22_X1 U10783 ( .A1(n9709), .A2(n9710), .B1(n6174), .B2(n9707), .ZN(
        P1_U3460) );
  OAI21_X1 U10784 ( .B1(n9660), .B2(n9701), .A(n9659), .ZN(n9663) );
  INV_X1 U10785 ( .A(n9661), .ZN(n9662) );
  AOI211_X1 U10786 ( .C1(n9699), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9711)
         );
  AOI22_X1 U10787 ( .A1(n9709), .A2(n9711), .B1(n6190), .B2(n9707), .ZN(
        P1_U3463) );
  INV_X1 U10788 ( .A(n9668), .ZN(n9671) );
  AOI21_X1 U10789 ( .B1(n9679), .B2(n9666), .A(n9665), .ZN(n9667) );
  OAI21_X1 U10790 ( .B1(n9668), .B2(n9682), .A(n9667), .ZN(n9669) );
  AOI211_X1 U10791 ( .C1(n9687), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9712)
         );
  AOI22_X1 U10792 ( .A1(n9709), .A2(n9712), .B1(n6228), .B2(n9707), .ZN(
        P1_U3466) );
  NAND3_X1 U10793 ( .A1(n6723), .A2(n9672), .A3(n9705), .ZN(n9674) );
  OAI211_X1 U10794 ( .C1(n9675), .C2(n9701), .A(n9674), .B(n9673), .ZN(n9676)
         );
  NOR2_X1 U10795 ( .A1(n9677), .A2(n9676), .ZN(n9713) );
  AOI22_X1 U10796 ( .A1(n9709), .A2(n9713), .B1(n6312), .B2(n9707), .ZN(
        P1_U3469) );
  NAND2_X1 U10797 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  OAI211_X1 U10798 ( .C1(n9683), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9684)
         );
  AOI211_X1 U10799 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9715)
         );
  AOI22_X1 U10800 ( .A1(n9709), .A2(n9715), .B1(n6496), .B2(n9707), .ZN(
        P1_U3472) );
  OAI211_X1 U10801 ( .C1(n4504), .C2(n9701), .A(n9689), .B(n9688), .ZN(n9690)
         );
  AOI21_X1 U10802 ( .B1(n9705), .B2(n9691), .A(n9690), .ZN(n9716) );
  INV_X1 U10803 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9692) );
  AOI22_X1 U10804 ( .A1(n9709), .A2(n9716), .B1(n9692), .B2(n9707), .ZN(
        P1_U3475) );
  INV_X1 U10805 ( .A(n9693), .ZN(n9698) );
  OAI21_X1 U10806 ( .B1(n9695), .B2(n9701), .A(n9694), .ZN(n9697) );
  AOI211_X1 U10807 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9717)
         );
  AOI22_X1 U10808 ( .A1(n9709), .A2(n9717), .B1(n6648), .B2(n9707), .ZN(
        P1_U3478) );
  OAI21_X1 U10809 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9703) );
  AOI211_X1 U10810 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9720)
         );
  INV_X1 U10811 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U10812 ( .A1(n9709), .A2(n9720), .B1(n9708), .B2(n9707), .ZN(
        P1_U3481) );
  AOI22_X1 U10813 ( .A1(n9721), .A2(n9710), .B1(n6177), .B2(n9718), .ZN(
        P1_U3525) );
  AOI22_X1 U10814 ( .A1(n9721), .A2(n9711), .B1(n6192), .B2(n9718), .ZN(
        P1_U3526) );
  AOI22_X1 U10815 ( .A1(n9721), .A2(n9712), .B1(n6229), .B2(n9718), .ZN(
        P1_U3527) );
  AOI22_X1 U10816 ( .A1(n9721), .A2(n9713), .B1(n6313), .B2(n9718), .ZN(
        P1_U3528) );
  AOI22_X1 U10817 ( .A1(n9721), .A2(n9715), .B1(n9714), .B2(n9718), .ZN(
        P1_U3529) );
  AOI22_X1 U10818 ( .A1(n9721), .A2(n9716), .B1(n9994), .B2(n9718), .ZN(
        P1_U3530) );
  AOI22_X1 U10819 ( .A1(n9721), .A2(n9717), .B1(n6649), .B2(n9718), .ZN(
        P1_U3531) );
  INV_X1 U10820 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10821 ( .A1(n9721), .A2(n9720), .B1(n9719), .B2(n9718), .ZN(
        P1_U3532) );
  AOI22_X1 U10822 ( .A1(n9722), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9724), .ZN(n9736) );
  INV_X1 U10823 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U10824 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  OAI211_X1 U10825 ( .C1(n9727), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9726), .B(
        n9725), .ZN(n9728) );
  INV_X1 U10826 ( .A(n9728), .ZN(n9734) );
  INV_X1 U10827 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9730) );
  OAI22_X1 U10828 ( .A1(n9731), .A2(n9730), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9729), .ZN(n9732) );
  INV_X1 U10829 ( .A(n9732), .ZN(n9733) );
  OAI221_X1 U10830 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9736), .C1(n9735), .C2(
        n9734), .A(n9733), .ZN(P2_U3245) );
  NAND2_X1 U10831 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  XOR2_X1 U10832 ( .A(n9751), .B(n9739), .Z(n9744) );
  AOI222_X1 U10833 ( .A1(n9745), .A2(n9744), .B1(n9743), .B2(n9742), .C1(n9741), .C2(n9740), .ZN(n9805) );
  NAND2_X1 U10834 ( .A1(n9747), .A2(n9746), .ZN(n9749) );
  NAND2_X1 U10835 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  XNOR2_X1 U10836 ( .A(n9751), .B(n9750), .ZN(n9808) );
  INV_X1 U10837 ( .A(n9752), .ZN(n9754) );
  OAI21_X1 U10838 ( .B1(n9803), .B2(n9754), .A(n9753), .ZN(n9804) );
  INV_X1 U10839 ( .A(n9804), .ZN(n9760) );
  OAI22_X1 U10840 ( .A1(n9757), .A2(n5066), .B1(n9756), .B2(n9755), .ZN(n9758)
         );
  AOI21_X1 U10841 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9761) );
  OAI21_X1 U10842 ( .B1(n9803), .B2(n9762), .A(n9761), .ZN(n9763) );
  AOI21_X1 U10843 ( .B1(n9764), .B2(n9808), .A(n9763), .ZN(n9765) );
  OAI21_X1 U10844 ( .B1(n9766), .B2(n9805), .A(n9765), .ZN(P2_U3292) );
  NOR2_X1 U10845 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  AND2_X1 U10846 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9772), .ZN(P2_U3297) );
  AND2_X1 U10847 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9772), .ZN(P2_U3298) );
  AND2_X1 U10848 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9772), .ZN(P2_U3299) );
  AND2_X1 U10849 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9772), .ZN(P2_U3300) );
  AND2_X1 U10850 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9772), .ZN(P2_U3301) );
  AND2_X1 U10851 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9772), .ZN(P2_U3302) );
  AND2_X1 U10852 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9772), .ZN(P2_U3303) );
  AND2_X1 U10853 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9772), .ZN(P2_U3304) );
  AND2_X1 U10854 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9772), .ZN(P2_U3305) );
  AND2_X1 U10855 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9772), .ZN(P2_U3306) );
  AND2_X1 U10856 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9772), .ZN(P2_U3307) );
  INV_X1 U10857 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U10858 ( .A1(n9769), .A2(n9922), .ZN(P2_U3308) );
  AND2_X1 U10859 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9772), .ZN(P2_U3309) );
  AND2_X1 U10860 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9772), .ZN(P2_U3310) );
  INV_X1 U10861 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U10862 ( .A1(n9769), .A2(n9912), .ZN(P2_U3311) );
  AND2_X1 U10863 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9772), .ZN(P2_U3312) );
  AND2_X1 U10864 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9772), .ZN(P2_U3313) );
  AND2_X1 U10865 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9772), .ZN(P2_U3314) );
  AND2_X1 U10866 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9772), .ZN(P2_U3315) );
  AND2_X1 U10867 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9772), .ZN(P2_U3316) );
  AND2_X1 U10868 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9772), .ZN(P2_U3317) );
  AND2_X1 U10869 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9772), .ZN(P2_U3318) );
  AND2_X1 U10870 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9772), .ZN(P2_U3319) );
  AND2_X1 U10871 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9772), .ZN(P2_U3320) );
  INV_X1 U10872 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U10873 ( .A1(n9769), .A2(n9939), .ZN(P2_U3321) );
  AND2_X1 U10874 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9772), .ZN(P2_U3322) );
  AND2_X1 U10875 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9772), .ZN(P2_U3323) );
  AND2_X1 U10876 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9772), .ZN(P2_U3324) );
  AND2_X1 U10877 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9772), .ZN(P2_U3325) );
  AND2_X1 U10878 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9772), .ZN(P2_U3326) );
  AOI22_X1 U10879 ( .A1(n9771), .A2(n9772), .B1(n9770), .B2(n9774), .ZN(
        P2_U3437) );
  AOI22_X1 U10880 ( .A1(n9775), .A2(n9774), .B1(n9773), .B2(n9772), .ZN(
        P2_U3438) );
  OAI22_X1 U10881 ( .A1(n9778), .A2(n9815), .B1(n9777), .B2(n9776), .ZN(n9779)
         );
  NOR2_X1 U10882 ( .A1(n9780), .A2(n9779), .ZN(n9841) );
  INV_X1 U10883 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U10884 ( .A1(n9840), .A2(n9841), .B1(n9955), .B2(n5900), .ZN(
        P2_U3451) );
  OR3_X1 U10885 ( .A1(n9782), .A2(n9781), .A3(n9826), .ZN(n9783) );
  OAI21_X1 U10886 ( .B1(n9784), .B2(n9835), .A(n9783), .ZN(n9786) );
  AOI211_X1 U10887 ( .C1(n9838), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9843)
         );
  INV_X1 U10888 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10889 ( .A1(n9840), .A2(n9843), .B1(n9909), .B2(n5900), .ZN(
        P2_U3454) );
  INV_X1 U10890 ( .A(n9788), .ZN(n9794) );
  OAI22_X1 U10891 ( .A1(n9790), .A2(n9826), .B1(n9789), .B2(n9835), .ZN(n9793)
         );
  INV_X1 U10892 ( .A(n9791), .ZN(n9792) );
  AOI211_X1 U10893 ( .C1(n9838), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9845)
         );
  INV_X1 U10894 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U10895 ( .A1(n9840), .A2(n9845), .B1(n9795), .B2(n5900), .ZN(
        P2_U3457) );
  INV_X1 U10896 ( .A(n9796), .ZN(n9801) );
  OAI22_X1 U10897 ( .A1(n9798), .A2(n9826), .B1(n9797), .B2(n9835), .ZN(n9800)
         );
  AOI211_X1 U10898 ( .C1(n9831), .C2(n9801), .A(n9800), .B(n9799), .ZN(n9846)
         );
  INV_X1 U10899 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9802) );
  AOI22_X1 U10900 ( .A1(n9840), .A2(n9846), .B1(n9802), .B2(n5900), .ZN(
        P2_U3460) );
  OAI22_X1 U10901 ( .A1(n9804), .A2(n9826), .B1(n9803), .B2(n9835), .ZN(n9807)
         );
  INV_X1 U10902 ( .A(n9805), .ZN(n9806) );
  AOI211_X1 U10903 ( .C1(n9838), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9847)
         );
  INV_X1 U10904 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10905 ( .A1(n9840), .A2(n9847), .B1(n9809), .B2(n5900), .ZN(
        P2_U3463) );
  AOI21_X1 U10906 ( .B1(n9812), .B2(n9811), .A(n9810), .ZN(n9813) );
  OAI211_X1 U10907 ( .C1(n9816), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9817)
         );
  INV_X1 U10908 ( .A(n9817), .ZN(n9849) );
  AOI22_X1 U10909 ( .A1(n9840), .A2(n9849), .B1(n5105), .B2(n5900), .ZN(
        P2_U3466) );
  AND2_X1 U10910 ( .A1(n9818), .A2(n9838), .ZN(n9823) );
  OAI21_X1 U10911 ( .B1(n9820), .B2(n9835), .A(n9819), .ZN(n9821) );
  NOR3_X1 U10912 ( .A1(n9823), .A2(n9822), .A3(n9821), .ZN(n9851) );
  AOI22_X1 U10913 ( .A1(n9840), .A2(n9851), .B1(n5139), .B2(n5900), .ZN(
        P2_U3472) );
  INV_X1 U10914 ( .A(n9824), .ZN(n9830) );
  OAI22_X1 U10915 ( .A1(n9827), .A2(n9826), .B1(n9825), .B2(n9835), .ZN(n9829)
         );
  AOI211_X1 U10916 ( .C1(n9831), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9852)
         );
  INV_X1 U10917 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10918 ( .A1(n9840), .A2(n9852), .B1(n9832), .B2(n5900), .ZN(
        P2_U3478) );
  OAI211_X1 U10919 ( .C1(n9836), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9837)
         );
  AOI21_X1 U10920 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(n9854) );
  AOI22_X1 U10921 ( .A1(n9840), .A2(n9854), .B1(n5219), .B2(n5900), .ZN(
        P2_U3484) );
  AOI22_X1 U10922 ( .A1(n9855), .A2(n9841), .B1(n9723), .B2(n9853), .ZN(
        P2_U3520) );
  INV_X1 U10923 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10924 ( .A1(n9855), .A2(n9843), .B1(n9842), .B2(n9853), .ZN(
        P2_U3521) );
  INV_X1 U10925 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U10926 ( .A1(n9855), .A2(n9845), .B1(n9844), .B2(n9853), .ZN(
        P2_U3522) );
  AOI22_X1 U10927 ( .A1(n9855), .A2(n9846), .B1(n5082), .B2(n9853), .ZN(
        P2_U3523) );
  AOI22_X1 U10928 ( .A1(n9855), .A2(n9847), .B1(n6361), .B2(n9853), .ZN(
        P2_U3524) );
  INV_X1 U10929 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10930 ( .A1(n9855), .A2(n9849), .B1(n9848), .B2(n9853), .ZN(
        P2_U3525) );
  INV_X1 U10931 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10932 ( .A1(n9855), .A2(n9851), .B1(n9850), .B2(n9853), .ZN(
        P2_U3527) );
  AOI22_X1 U10933 ( .A1(n9855), .A2(n9852), .B1(n6685), .B2(n9853), .ZN(
        P2_U3529) );
  AOI22_X1 U10934 ( .A1(n9855), .A2(n9854), .B1(n6692), .B2(n9853), .ZN(
        P2_U3531) );
  INV_X1 U10935 ( .A(n9856), .ZN(n9857) );
  NAND2_X1 U10936 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  XOR2_X1 U10937 ( .A(n9860), .B(n9859), .Z(ADD_1071_U5) );
  XOR2_X1 U10938 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10939 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(ADD_1071_U56) );
  OAI21_X1 U10940 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(ADD_1071_U57) );
  OAI21_X1 U10941 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(ADD_1071_U58) );
  OAI21_X1 U10942 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(ADD_1071_U59) );
  OAI21_X1 U10943 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(ADD_1071_U60) );
  OAI21_X1 U10944 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(ADD_1071_U61) );
  AOI21_X1 U10945 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(ADD_1071_U62) );
  AOI21_X1 U10946 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(ADD_1071_U63) );
  NAND4_X1 U10947 ( .A1(keyinput20), .A2(keyinput44), .A3(keyinput16), .A4(
        keyinput35), .ZN(n9888) );
  NAND4_X1 U10948 ( .A1(keyinput43), .A2(keyinput39), .A3(keyinput62), .A4(
        keyinput63), .ZN(n9887) );
  NAND4_X1 U10949 ( .A1(keyinput55), .A2(keyinput10), .A3(keyinput11), .A4(
        keyinput6), .ZN(n9886) );
  NAND4_X1 U10950 ( .A1(keyinput30), .A2(keyinput27), .A3(keyinput19), .A4(
        keyinput23), .ZN(n9885) );
  NOR4_X1 U10951 ( .A1(n9888), .A2(n9887), .A3(n9886), .A4(n9885), .ZN(n10028)
         );
  NAND3_X1 U10952 ( .A1(keyinput49), .A2(keyinput22), .A3(keyinput56), .ZN(
        n9906) );
  NOR2_X1 U10953 ( .A1(keyinput4), .A2(keyinput7), .ZN(n9892) );
  NAND3_X1 U10954 ( .A1(keyinput51), .A2(keyinput14), .A3(keyinput54), .ZN(
        n9890) );
  NAND3_X1 U10955 ( .A1(keyinput18), .A2(keyinput40), .A3(keyinput41), .ZN(
        n9889) );
  NOR4_X1 U10956 ( .A1(keyinput50), .A2(keyinput37), .A3(n9890), .A4(n9889), 
        .ZN(n9891) );
  NAND4_X1 U10957 ( .A1(keyinput26), .A2(keyinput34), .A3(n9892), .A4(n9891), 
        .ZN(n9905) );
  NAND3_X1 U10958 ( .A1(keyinput60), .A2(keyinput52), .A3(keyinput61), .ZN(
        n9903) );
  NOR2_X1 U10959 ( .A1(keyinput8), .A2(keyinput3), .ZN(n9896) );
  NAND3_X1 U10960 ( .A1(keyinput15), .A2(keyinput48), .A3(keyinput2), .ZN(
        n9894) );
  NAND3_X1 U10961 ( .A1(keyinput29), .A2(keyinput21), .A3(keyinput25), .ZN(
        n9893) );
  NOR4_X1 U10962 ( .A1(keyinput59), .A2(keyinput45), .A3(n9894), .A4(n9893), 
        .ZN(n9895) );
  NAND4_X1 U10963 ( .A1(keyinput24), .A2(keyinput0), .A3(n9896), .A4(n9895), 
        .ZN(n9902) );
  NOR4_X1 U10964 ( .A1(keyinput9), .A2(keyinput5), .A3(keyinput1), .A4(
        keyinput33), .ZN(n9900) );
  NOR4_X1 U10965 ( .A1(keyinput53), .A2(keyinput28), .A3(keyinput32), .A4(
        keyinput42), .ZN(n9899) );
  NOR4_X1 U10966 ( .A1(keyinput46), .A2(keyinput47), .A3(keyinput38), .A4(
        keyinput31), .ZN(n9898) );
  AND4_X1 U10967 ( .A1(keyinput13), .A2(keyinput17), .A3(keyinput12), .A4(
        keyinput57), .ZN(n9897) );
  NAND4_X1 U10968 ( .A1(n9900), .A2(n9899), .A3(n9898), .A4(n9897), .ZN(n9901)
         );
  OR4_X1 U10969 ( .A1(keyinput58), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(
        n9904) );
  NOR4_X1 U10970 ( .A1(keyinput36), .A2(n9906), .A3(n9905), .A4(n9904), .ZN(
        n10027) );
  INV_X1 U10971 ( .A(keyinput36), .ZN(n9908) );
  AOI22_X1 U10972 ( .A1(n9909), .A2(keyinput49), .B1(P1_ADDR_REG_6__SCAN_IN), 
        .B2(n9908), .ZN(n9907) );
  OAI221_X1 U10973 ( .B1(n9909), .B2(keyinput49), .C1(n9908), .C2(
        P1_ADDR_REG_6__SCAN_IN), .A(n9907), .ZN(n9919) );
  AOI22_X1 U10974 ( .A1(n9912), .A2(keyinput4), .B1(keyinput26), .B2(n9911), 
        .ZN(n9910) );
  OAI221_X1 U10975 ( .B1(n9912), .B2(keyinput4), .C1(n9911), .C2(keyinput26), 
        .A(n9910), .ZN(n9918) );
  XNOR2_X1 U10976 ( .A(P1_B_REG_SCAN_IN), .B(keyinput56), .ZN(n9916) );
  XNOR2_X1 U10977 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput22), .ZN(n9915) );
  XNOR2_X1 U10978 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput7), .ZN(n9914) );
  XNOR2_X1 U10979 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput34), .ZN(n9913) );
  NAND4_X1 U10980 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n9917)
         );
  NOR3_X1 U10981 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(n9967) );
  AOI22_X1 U10982 ( .A1(n9922), .A2(keyinput51), .B1(keyinput14), .B2(n9921), 
        .ZN(n9920) );
  OAI221_X1 U10983 ( .B1(n9922), .B2(keyinput51), .C1(n9921), .C2(keyinput14), 
        .A(n9920), .ZN(n9935) );
  INV_X1 U10984 ( .A(SI_26_), .ZN(n9925) );
  INV_X1 U10985 ( .A(keyinput50), .ZN(n9924) );
  AOI22_X1 U10986 ( .A1(n9925), .A2(keyinput54), .B1(P2_ADDR_REG_0__SCAN_IN), 
        .B2(n9924), .ZN(n9923) );
  OAI221_X1 U10987 ( .B1(n9925), .B2(keyinput54), .C1(n9924), .C2(
        P2_ADDR_REG_0__SCAN_IN), .A(n9923), .ZN(n9934) );
  INV_X1 U10988 ( .A(keyinput18), .ZN(n9927) );
  AOI22_X1 U10989 ( .A1(n9928), .A2(keyinput37), .B1(P2_ADDR_REG_6__SCAN_IN), 
        .B2(n9927), .ZN(n9926) );
  OAI221_X1 U10990 ( .B1(n9928), .B2(keyinput37), .C1(n9927), .C2(
        P2_ADDR_REG_6__SCAN_IN), .A(n9926), .ZN(n9933) );
  INV_X1 U10991 ( .A(keyinput40), .ZN(n9930) );
  AOI22_X1 U10992 ( .A1(n9931), .A2(keyinput41), .B1(P2_ADDR_REG_1__SCAN_IN), 
        .B2(n9930), .ZN(n9929) );
  OAI221_X1 U10993 ( .B1(n9931), .B2(keyinput41), .C1(n9930), .C2(
        P2_ADDR_REG_1__SCAN_IN), .A(n9929), .ZN(n9932) );
  NOR4_X1 U10994 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(n9966)
         );
  AOI22_X1 U10995 ( .A1(n6763), .A2(keyinput52), .B1(n9937), .B2(keyinput61), 
        .ZN(n9936) );
  OAI221_X1 U10996 ( .B1(n6763), .B2(keyinput52), .C1(n9937), .C2(keyinput61), 
        .A(n9936), .ZN(n9949) );
  AOI22_X1 U10997 ( .A1(n9940), .A2(keyinput0), .B1(keyinput3), .B2(n9939), 
        .ZN(n9938) );
  OAI221_X1 U10998 ( .B1(n9940), .B2(keyinput0), .C1(n9939), .C2(keyinput3), 
        .A(n9938), .ZN(n9948) );
  INV_X1 U10999 ( .A(SI_6_), .ZN(n9942) );
  AOI22_X1 U11000 ( .A1(n9943), .A2(keyinput8), .B1(n9942), .B2(keyinput24), 
        .ZN(n9941) );
  OAI221_X1 U11001 ( .B1(n9943), .B2(keyinput8), .C1(n9942), .C2(keyinput24), 
        .A(n9941), .ZN(n9947) );
  XNOR2_X1 U11002 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput60), .ZN(n9945) );
  XNOR2_X1 U11003 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput58), .ZN(n9944) );
  NAND2_X1 U11004 ( .A1(n9945), .A2(n9944), .ZN(n9946) );
  NOR4_X1 U11005 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n9965)
         );
  INV_X1 U11006 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11007 ( .A1(n9951), .A2(keyinput15), .B1(keyinput48), .B2(n6681), 
        .ZN(n9950) );
  OAI221_X1 U11008 ( .B1(n9951), .B2(keyinput15), .C1(n6681), .C2(keyinput48), 
        .A(n9950), .ZN(n9963) );
  AOI22_X1 U11009 ( .A1(n9953), .A2(keyinput59), .B1(keyinput2), .B2(n5129), 
        .ZN(n9952) );
  OAI221_X1 U11010 ( .B1(n9953), .B2(keyinput59), .C1(n5129), .C2(keyinput2), 
        .A(n9952), .ZN(n9962) );
  AOI22_X1 U11011 ( .A1(n9956), .A2(keyinput45), .B1(keyinput29), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11012 ( .B1(n9956), .B2(keyinput45), .C1(n9955), .C2(keyinput29), 
        .A(n9954), .ZN(n9961) );
  AOI22_X1 U11013 ( .A1(n9959), .A2(keyinput21), .B1(keyinput25), .B2(n9958), 
        .ZN(n9957) );
  OAI221_X1 U11014 ( .B1(n9959), .B2(keyinput21), .C1(n9958), .C2(keyinput25), 
        .A(n9957), .ZN(n9960) );
  NOR4_X1 U11015 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9964)
         );
  NAND4_X1 U11016 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n10026) );
  AOI22_X1 U11017 ( .A1(n7151), .A2(keyinput20), .B1(n4879), .B2(keyinput39), 
        .ZN(n9968) );
  OAI221_X1 U11018 ( .B1(n7151), .B2(keyinput20), .C1(n4879), .C2(keyinput39), 
        .A(n9968), .ZN(n9980) );
  AOI22_X1 U11019 ( .A1(n9970), .A2(keyinput1), .B1(keyinput32), .B2(n5043), 
        .ZN(n9969) );
  OAI221_X1 U11020 ( .B1(n9970), .B2(keyinput1), .C1(n5043), .C2(keyinput32), 
        .A(n9969), .ZN(n9979) );
  INV_X1 U11021 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9973) );
  INV_X1 U11022 ( .A(keyinput5), .ZN(n9972) );
  AOI22_X1 U11023 ( .A1(n9973), .A2(keyinput33), .B1(P1_ADDR_REG_1__SCAN_IN), 
        .B2(n9972), .ZN(n9971) );
  OAI221_X1 U11024 ( .B1(n9973), .B2(keyinput33), .C1(n9972), .C2(
        P1_ADDR_REG_1__SCAN_IN), .A(n9971), .ZN(n9978) );
  INV_X1 U11025 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11026 ( .A1(n9976), .A2(keyinput47), .B1(n9975), .B2(keyinput27), 
        .ZN(n9974) );
  OAI221_X1 U11027 ( .B1(n9976), .B2(keyinput47), .C1(n9975), .C2(keyinput27), 
        .A(n9974), .ZN(n9977) );
  NOR4_X1 U11028 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n10024)
         );
  AOI22_X1 U11029 ( .A1(n8407), .A2(keyinput9), .B1(n8955), .B2(keyinput31), 
        .ZN(n9981) );
  OAI221_X1 U11030 ( .B1(n8407), .B2(keyinput9), .C1(n8955), .C2(keyinput31), 
        .A(n9981), .ZN(n9986) );
  AOI22_X1 U11031 ( .A1(n5564), .A2(keyinput35), .B1(P1_U3084), .B2(keyinput62), .ZN(n9982) );
  OAI221_X1 U11032 ( .B1(n5564), .B2(keyinput35), .C1(P1_U3084), .C2(
        keyinput62), .A(n9982), .ZN(n9985) );
  XNOR2_X1 U11033 ( .A(n9983), .B(keyinput23), .ZN(n9984) );
  OR3_X1 U11034 ( .A1(n9986), .A2(n9985), .A3(n9984), .ZN(n9992) );
  AOI22_X1 U11035 ( .A1(n7652), .A2(keyinput13), .B1(keyinput19), .B2(n9988), 
        .ZN(n9987) );
  OAI221_X1 U11036 ( .B1(n7652), .B2(keyinput13), .C1(n9988), .C2(keyinput19), 
        .A(n9987), .ZN(n9991) );
  INV_X1 U11037 ( .A(keyinput44), .ZN(n9989) );
  XNOR2_X1 U11038 ( .A(n9989), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n9990) );
  NOR3_X1 U11039 ( .A1(n9992), .A2(n9991), .A3(n9990), .ZN(n10023) );
  AOI22_X1 U11040 ( .A1(n9995), .A2(keyinput57), .B1(n9994), .B2(keyinput6), 
        .ZN(n9993) );
  OAI221_X1 U11041 ( .B1(n9995), .B2(keyinput57), .C1(n9994), .C2(keyinput6), 
        .A(n9993), .ZN(n10006) );
  AOI22_X1 U11042 ( .A1(n5118), .A2(keyinput38), .B1(n9997), .B2(keyinput10), 
        .ZN(n9996) );
  OAI221_X1 U11043 ( .B1(n5118), .B2(keyinput38), .C1(n9997), .C2(keyinput10), 
        .A(n9996), .ZN(n10005) );
  INV_X1 U11044 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9999) );
  AOI22_X1 U11045 ( .A1(n5105), .A2(keyinput43), .B1(n9999), .B2(keyinput55), 
        .ZN(n9998) );
  OAI221_X1 U11046 ( .B1(n5105), .B2(keyinput43), .C1(n9999), .C2(keyinput55), 
        .A(n9998), .ZN(n10004) );
  AOI22_X1 U11047 ( .A1(n10002), .A2(keyinput28), .B1(keyinput30), .B2(n10001), 
        .ZN(n10000) );
  OAI221_X1 U11048 ( .B1(n10002), .B2(keyinput28), .C1(n10001), .C2(keyinput30), .A(n10000), .ZN(n10003) );
  NOR4_X1 U11049 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10022) );
  INV_X1 U11050 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U11051 ( .A1(n10009), .A2(keyinput46), .B1(n10008), .B2(keyinput17), 
        .ZN(n10007) );
  OAI221_X1 U11052 ( .B1(n10009), .B2(keyinput46), .C1(n10008), .C2(keyinput17), .A(n10007), .ZN(n10020) );
  AOI22_X1 U11053 ( .A1(n10011), .A2(keyinput53), .B1(keyinput11), .B2(n6685), 
        .ZN(n10010) );
  OAI221_X1 U11054 ( .B1(n10011), .B2(keyinput53), .C1(n6685), .C2(keyinput11), 
        .A(n10010), .ZN(n10019) );
  AOI22_X1 U11055 ( .A1(n7005), .A2(keyinput42), .B1(n10013), .B2(keyinput12), 
        .ZN(n10012) );
  OAI221_X1 U11056 ( .B1(n7005), .B2(keyinput42), .C1(n10013), .C2(keyinput12), 
        .A(n10012), .ZN(n10018) );
  AOI22_X1 U11057 ( .A1(n10016), .A2(keyinput16), .B1(keyinput63), .B2(n10015), 
        .ZN(n10014) );
  OAI221_X1 U11058 ( .B1(n10016), .B2(keyinput16), .C1(n10015), .C2(keyinput63), .A(n10014), .ZN(n10017) );
  NOR4_X1 U11059 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10021) );
  NAND4_X1 U11060 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10025) );
  AOI211_X1 U11061 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10044) );
  AND2_X1 U11062 ( .A1(n10030), .A2(n10029), .ZN(n10040) );
  AOI22_X1 U11063 ( .A1(n9648), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10032), 
        .B2(n10031), .ZN(n10036) );
  NAND2_X1 U11064 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  OAI211_X1 U11065 ( .C1(n10038), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10039) );
  AOI211_X1 U11066 ( .C1(n10042), .C2(n10041), .A(n10040), .B(n10039), .ZN(
        n10043) );
  XNOR2_X1 U11067 ( .A(n10044), .B(n10043), .ZN(P1_U3277) );
  XOR2_X1 U11068 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10045), .Z(ADD_1071_U50) );
  NOR2_X1 U11069 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  XOR2_X1 U11070 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10048), .Z(ADD_1071_U51) );
  OAI21_X1 U11071 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(n10052) );
  XNOR2_X1 U11072 ( .A(n10052), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11073 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U47) );
  XOR2_X1 U11074 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10056), .Z(ADD_1071_U48) );
  XOR2_X1 U11075 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10057), .Z(ADD_1071_U49) );
  XOR2_X1 U11076 ( .A(n10059), .B(n10058), .Z(ADD_1071_U54) );
  XOR2_X1 U11077 ( .A(n10061), .B(n10060), .Z(ADD_1071_U53) );
  XNOR2_X1 U11078 ( .A(n10063), .B(n10062), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5072 ( .A(n5051), .Z(n6354) );
  CLKBUF_X1 U5277 ( .A(n6215), .Z(n7957) );
endmodule

