

module b14_C_SARLock_k_64_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665;

  NAND2_X1 U2265 ( .A1(n4046), .A2(n2452), .ZN(n4034) );
  CLKBUF_X2 U2266 ( .A(n2294), .Z(n3588) );
  OR2_X1 U2267 ( .A1(n2266), .A2(n2659), .ZN(n2270) );
  AOI21_X1 U2269 ( .B1(n4034), .B2(n2467), .A(n2466), .ZN(n4008) );
  BUF_X1 U2270 ( .A(n2286), .Z(n3590) );
  XNOR2_X1 U2271 ( .A(n3841), .B(n3842), .ZN(n4127) );
  NOR2_X2 U2272 ( .A1(n2271), .A2(IR_REG_27__SCAN_IN), .ZN(n2564) );
  NOR2_X2 U2273 ( .A1(n2743), .A2(n2742), .ZN(n2741) );
  AND2_X1 U2274 ( .A1(n4468), .A2(n2269), .ZN(n2294) );
  NAND4_X1 U2275 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .ZN(n3756)
         );
  CLKBUF_X2 U2276 ( .A(n2295), .Z(n2318) );
  INV_X4 U2277 ( .A(n3457), .ZN(n3413) );
  NAND2_X1 U2278 ( .A1(n2562), .A2(n4470), .ZN(n2845) );
  INV_X2 U2279 ( .A(IR_REG_31__SCAN_IN), .ZN(n2659) );
  OR2_X1 U2280 ( .A1(n3877), .A2(n2253), .ZN(n2235) );
  NAND2_X1 U2281 ( .A1(n2492), .A2(n2491), .ZN(n3967) );
  NOR2_X1 U2282 ( .A1(n4559), .A2(REG1_REG_16__SCAN_IN), .ZN(n4560) );
  XNOR2_X1 U2283 ( .A(n3812), .B(n3811), .ZN(n4559) );
  NAND2_X1 U2284 ( .A1(n4548), .A2(n3810), .ZN(n3812) );
  NAND2_X1 U2285 ( .A1(n4539), .A2(n3809), .ZN(n4549) );
  NAND2_X1 U2286 ( .A1(n4505), .A2(n3043), .ZN(n4515) );
  NOR2_X1 U2287 ( .A1(n4124), .A2(n3465), .ZN(n3296) );
  AND2_X1 U2288 ( .A1(n3678), .A2(n3675), .ZN(n3636) );
  NOR2_X1 U2289 ( .A1(n2697), .A2(n2209), .ZN(n2768) );
  NAND2_X1 U2290 ( .A1(n3755), .A2(n3025), .ZN(n3684) );
  INV_X1 U2291 ( .A(n2916), .ZN(n3755) );
  NAND2_X2 U2292 ( .A1(n2288), .A2(n2287), .ZN(n2291) );
  AND4_X1 U2293 ( .A1(n2312), .A2(n2311), .A3(n2310), .A4(n2309), .ZN(n2916)
         );
  AND3_X1 U2294 ( .A1(n2285), .A2(n2284), .A3(n2283), .ZN(n2288) );
  AND2_X2 U2295 ( .A1(n2843), .A2(n4588), .ZN(n4607) );
  AND2_X1 U2296 ( .A1(n2760), .A2(n2211), .ZN(n2743) );
  NAND2_X1 U2297 ( .A1(n2267), .A2(n2660), .ZN(n2268) );
  XNOR2_X1 U2298 ( .A(n2270), .B(n2263), .ZN(n2269) );
  MUX2_X1 U2299 ( .A(IR_REG_31__SCAN_IN), .B(n2265), .S(IR_REG_29__SCAN_IN), 
        .Z(n2267) );
  NAND2_X2 U2300 ( .A1(n2708), .A2(n2845), .ZN(n3456) );
  NAND2_X2 U2301 ( .A1(n2845), .A2(n2781), .ZN(n3457) );
  NAND2_X1 U2302 ( .A1(n2121), .A2(n2123), .ZN(n4479) );
  AND2_X1 U2303 ( .A1(n2228), .A2(n2261), .ZN(n2161) );
  AND4_X1 U2304 ( .A1(n2145), .A2(n2144), .A3(n2143), .A4(n2142), .ZN(n2228)
         );
  AND4_X1 U2305 ( .A1(n2260), .A2(n2259), .A3(n2258), .A4(n2557), .ZN(n2261)
         );
  NOR2_X1 U2306 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2289)
         );
  NOR2_X1 U2307 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2260)
         );
  NOR2_X1 U2308 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2259)
         );
  NOR2_X1 U2309 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2258)
         );
  INV_X1 U2310 ( .A(IR_REG_20__SCAN_IN), .ZN(n2557) );
  NOR2_X1 U2311 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2145)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2144)
         );
  NOR2_X1 U2313 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2143)
         );
  NOR2_X1 U2314 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2142)
         );
  NOR2_X1 U2315 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2087)
         );
  NOR2_X1 U2316 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2248)
         );
  AOI211_X1 U2317 ( .C1(n4127), .C2(n4651), .A(n4126), .B(n4125), .ZN(n4264)
         );
  OAI21_X2 U2318 ( .B1(n3895), .B2(n2250), .A(n2530), .ZN(n3877) );
  OAI21_X2 U2319 ( .B1(n3942), .B2(n2238), .A(n2236), .ZN(n3895) );
  OAI21_X2 U2320 ( .B1(n3967), .B2(n2502), .A(n2501), .ZN(n3955) );
  NAND2_X1 U2321 ( .A1(n4515), .A2(n4516), .ZN(n4514) );
  NOR2_X1 U2322 ( .A1(n2198), .A2(n2197), .ZN(n2196) );
  NOR2_X1 U2323 ( .A1(n3340), .A2(n3428), .ZN(n2197) );
  INV_X1 U2324 ( .A(n3336), .ZN(n2198) );
  OR2_X2 U2325 ( .A1(n3076), .A2(n3456), .ZN(n3459) );
  OAI22_X1 U2326 ( .A1(n2768), .A2(n2698), .B1(n4663), .B2(n2770), .ZN(n2208)
         );
  AND2_X1 U2327 ( .A1(n2656), .A2(n2272), .ZN(n2274) );
  AND2_X1 U2328 ( .A1(n2179), .A2(n2175), .ZN(n2174) );
  INV_X1 U2329 ( .A(n3462), .ZN(n2175) );
  INV_X1 U2330 ( .A(n2845), .ZN(n2085) );
  INV_X1 U2331 ( .A(n2295), .ZN(n2571) );
  NAND2_X1 U2332 ( .A1(n2675), .A2(n2676), .ZN(n3772) );
  XNOR2_X1 U2333 ( .A(n2134), .B(n2687), .ZN(n3787) );
  XNOR2_X1 U2334 ( .A(n2208), .B(n3055), .ZN(n3040) );
  NAND2_X1 U2335 ( .A1(n4514), .A2(n3044), .ZN(n3045) );
  NOR2_X1 U2336 ( .A1(n3724), .A2(n3842), .ZN(n2163) );
  NAND2_X1 U2337 ( .A1(n2562), .A2(n2844), .ZN(n4640) );
  NAND2_X1 U2338 ( .A1(n3065), .A2(n4525), .ZN(n3796) );
  NOR2_X1 U2339 ( .A1(n4536), .A2(n2426), .ZN(n4535) );
  NOR2_X1 U2340 ( .A1(n4621), .A2(REG1_REG_17__SCAN_IN), .ZN(n2207) );
  NAND2_X1 U2341 ( .A1(n4582), .A2(n4583), .ZN(n4580) );
  NAND2_X1 U2342 ( .A1(n2262), .A2(n2244), .ZN(n2243) );
  INV_X1 U2343 ( .A(IR_REG_22__SCAN_IN), .ZN(n2262) );
  INV_X1 U2344 ( .A(n3445), .ZN(n2191) );
  NOR2_X1 U2345 ( .A1(n2024), .A2(n3445), .ZN(n2189) );
  INV_X1 U2346 ( .A(n2196), .ZN(n2083) );
  AND2_X1 U2347 ( .A1(n2195), .A2(n2081), .ZN(n2080) );
  NAND2_X1 U2348 ( .A1(n2196), .A2(n2082), .ZN(n2081) );
  NAND2_X1 U2349 ( .A1(n2249), .A2(n2043), .ZN(n2233) );
  AND2_X1 U2350 ( .A1(n3970), .A2(n2596), .ZN(n3711) );
  NOR2_X1 U2351 ( .A1(n3603), .A2(n2158), .ZN(n2157) );
  NAND2_X1 U2352 ( .A1(n2378), .A2(n2227), .ZN(n2226) );
  NAND2_X1 U2353 ( .A1(n3684), .A2(n3681), .ZN(n3022) );
  NAND2_X1 U2354 ( .A1(n2291), .A2(n2831), .ZN(n3678) );
  NAND2_X1 U2355 ( .A1(n2800), .A2(n3636), .ZN(n2799) );
  NOR2_X1 U2356 ( .A1(n3943), .A2(n4161), .ZN(n2102) );
  NOR2_X1 U2357 ( .A1(n4018), .A2(n3361), .ZN(n3977) );
  AND2_X1 U2358 ( .A1(n3175), .A2(n3208), .ZN(n2100) );
  INV_X1 U2359 ( .A(n2242), .ZN(n2086) );
  INV_X1 U2360 ( .A(IR_REG_23__SCAN_IN), .ZN(n2621) );
  NOR2_X2 U2361 ( .A1(n2071), .A2(n2301), .ZN(n2162) );
  INV_X1 U2362 ( .A(IR_REG_13__SCAN_IN), .ZN(n2257) );
  OR2_X1 U2363 ( .A1(n2473), .A2(IR_REG_17__SCAN_IN), .ZN(n2486) );
  INV_X1 U2364 ( .A(IR_REG_14__SCAN_IN), .ZN(n2460) );
  AND2_X1 U2365 ( .A1(n3544), .A2(n3382), .ZN(n2066) );
  XNOR2_X1 U2366 ( .A(n2870), .B(n3457), .ZN(n2913) );
  OAI21_X1 U2367 ( .B1(n3353), .B2(n2193), .A(n2057), .ZN(n2192) );
  INV_X1 U2368 ( .A(n3552), .ZN(n2193) );
  NAND2_X1 U2369 ( .A1(n2182), .A2(n3562), .ZN(n2181) );
  NAND2_X1 U2370 ( .A1(n2028), .A2(n2056), .ZN(n2178) );
  INV_X1 U2371 ( .A(n2178), .ZN(n2177) );
  AOI21_X1 U2372 ( .B1(n2712), .B2(n2957), .A(n2709), .ZN(n2784) );
  INV_X1 U2373 ( .A(n4162), .ZN(n3477) );
  NAND2_X1 U2374 ( .A1(n2077), .A2(n2076), .ZN(n2079) );
  INV_X1 U2375 ( .A(n3509), .ZN(n2076) );
  NAND2_X1 U2376 ( .A1(n3507), .A2(n3510), .ZN(n2077) );
  OR2_X1 U2377 ( .A1(n2519), .A2(n4429), .ZN(n2526) );
  AOI21_X1 U2378 ( .B1(n3436), .B2(n3402), .A(n3401), .ZN(n3509) );
  OAI21_X1 U2379 ( .B1(n3459), .B2(n2575), .A(n2714), .ZN(n2785) );
  NOR2_X1 U2380 ( .A1(n2494), .A2(n4346), .ZN(n2504) );
  OR2_X1 U2381 ( .A1(n3475), .A2(n2255), .ZN(n2067) );
  INV_X1 U2382 ( .A(n3170), .ZN(n2070) );
  NOR2_X1 U2383 ( .A1(n2526), .A2(n4347), .ZN(n2538) );
  NOR2_X1 U2384 ( .A1(n2424), .A2(n4371), .ZN(n2443) );
  NAND2_X1 U2385 ( .A1(n3312), .A2(n2150), .ZN(n2152) );
  NOR2_X1 U2386 ( .A1(n2268), .A2(n2151), .ZN(n2150) );
  INV_X1 U2387 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2151) );
  OR2_X1 U2388 ( .A1(n2269), .A2(n2148), .ZN(n2147) );
  INV_X1 U2389 ( .A(IR_REG_1__SCAN_IN), .ZN(n2124) );
  INV_X1 U2390 ( .A(IR_REG_0__SCAN_IN), .ZN(n2112) );
  NAND2_X1 U2391 ( .A1(n2120), .A2(n2674), .ZN(n2119) );
  INV_X1 U2392 ( .A(n2123), .ZN(n2120) );
  XNOR2_X1 U2393 ( .A(n2690), .B(n2763), .ZN(n2757) );
  AOI21_X1 U2394 ( .B1(n3787), .B2(REG2_REG_3__SCAN_IN), .A(n2038), .ZN(n2677)
         );
  NAND2_X1 U2395 ( .A1(n2757), .A2(REG1_REG_4__SCAN_IN), .ZN(n2760) );
  NOR2_X1 U2396 ( .A1(n2772), .A2(n2980), .ZN(n2107) );
  NOR2_X1 U2397 ( .A1(n2772), .A2(n2106), .ZN(n2105) );
  NAND2_X1 U2398 ( .A1(n2033), .A2(n2061), .ZN(n4494) );
  NAND2_X1 U2399 ( .A1(n3040), .A2(REG1_REG_8__SCAN_IN), .ZN(n2061) );
  NAND2_X1 U2400 ( .A1(n4531), .A2(n3046), .ZN(n3050) );
  NAND2_X1 U2401 ( .A1(n4564), .A2(n2141), .ZN(n2140) );
  OR2_X1 U2402 ( .A1(n4621), .A2(REG2_REG_17__SCAN_IN), .ZN(n2141) );
  OR2_X1 U2403 ( .A1(n2548), .A2(n3464), .ZN(n3835) );
  AND2_X1 U2404 ( .A1(n4059), .A2(n3839), .ZN(n2096) );
  INV_X1 U2405 ( .A(n2252), .ZN(n2234) );
  NAND2_X1 U2406 ( .A1(n2601), .A2(n2026), .ZN(n2164) );
  AOI21_X1 U2407 ( .B1(n2239), .B2(n2237), .A(n2049), .ZN(n2236) );
  INV_X1 U2408 ( .A(n2239), .ZN(n2238) );
  INV_X1 U2409 ( .A(n2518), .ZN(n2237) );
  AND4_X1 U2410 ( .A1(n2448), .A2(n2447), .A3(n2446), .A4(n2445), .ZN(n4031)
         );
  AOI21_X1 U2411 ( .B1(n2223), .B2(n2222), .A(n2046), .ZN(n2221) );
  INV_X1 U2412 ( .A(n3217), .ZN(n2225) );
  AOI21_X1 U2413 ( .B1(n2170), .B2(n2168), .A(n2167), .ZN(n2166) );
  INV_X1 U2414 ( .A(n2170), .ZN(n2169) );
  INV_X1 U2415 ( .A(n3704), .ZN(n2167) );
  AOI21_X1 U2416 ( .B1(n2219), .B2(n2364), .A(n2037), .ZN(n2217) );
  OAI21_X1 U2417 ( .B1(n3070), .B2(n2583), .A(n3693), .ZN(n3137) );
  OAI21_X1 U2418 ( .B1(n3023), .B2(n2580), .A(n3684), .ZN(n2941) );
  OAI21_X1 U2419 ( .B1(n2486), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2488) );
  INV_X1 U2420 ( .A(IR_REG_19__SCAN_IN), .ZN(n2487) );
  INV_X1 U2421 ( .A(n3022), .ZN(n3638) );
  NAND2_X1 U2422 ( .A1(n2708), .A2(n4617), .ZN(n2838) );
  NAND2_X1 U2423 ( .A1(n2575), .A2(n2797), .ZN(n3671) );
  NAND2_X1 U2424 ( .A1(n3887), .A2(n2029), .ZN(n3309) );
  NOR2_X1 U2425 ( .A1(n3925), .A2(n4141), .ZN(n3900) );
  INV_X1 U2426 ( .A(n3746), .ZN(n4145) );
  INV_X1 U2427 ( .A(n4047), .ZN(n4212) );
  NOR2_X1 U2428 ( .A1(n4103), .A2(n3276), .ZN(n3236) );
  NAND2_X1 U2429 ( .A1(n3628), .A2(n2606), .ZN(n4047) );
  AND2_X1 U2430 ( .A1(n2617), .A2(n2664), .ZN(n2662) );
  NAND2_X1 U2431 ( .A1(n2622), .A2(n2621), .ZN(n2620) );
  OAI21_X1 U2432 ( .B1(n2622), .B2(n2621), .A(n2620), .ZN(n2877) );
  INV_X1 U2433 ( .A(IR_REG_15__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U2434 ( .A1(n2659), .A2(IR_REG_1__SCAN_IN), .ZN(n2123) );
  NAND2_X1 U2435 ( .A1(n2110), .A2(n2111), .ZN(n2121) );
  NAND2_X1 U2436 ( .A1(n2112), .A2(n2124), .ZN(n2110) );
  NAND2_X1 U2437 ( .A1(n2122), .A2(IR_REG_0__SCAN_IN), .ZN(n2111) );
  NAND2_X1 U2438 ( .A1(n2067), .A2(n2066), .ZN(n3542) );
  INV_X1 U2439 ( .A(n3747), .ZN(n3921) );
  NAND2_X1 U2440 ( .A1(n2931), .A2(n2930), .ZN(n2952) );
  NAND2_X1 U2441 ( .A1(n2790), .A2(n2734), .ZN(n3576) );
  INV_X1 U2442 ( .A(n4171), .ZN(n3547) );
  OR2_X1 U2443 ( .A1(n2819), .A2(n2818), .ZN(n2084) );
  NAND2_X1 U2444 ( .A1(n2825), .A2(n2873), .ZN(n2826) );
  OR2_X1 U2445 ( .A1(n2824), .A2(n2823), .ZN(n2825) );
  NAND2_X1 U2446 ( .A1(n2790), .A2(n2789), .ZN(n3567) );
  OAI211_X1 U2447 ( .C1(n3868), .C2(n2571), .A(n2541), .B(n2540), .ZN(n4122)
         );
  NAND4_X1 U2448 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n4236)
         );
  NAND3_X1 U2449 ( .A1(n2126), .A2(n2128), .A3(n2125), .ZN(n4536) );
  AND2_X1 U2450 ( .A1(n2129), .A2(n2132), .ZN(n2128) );
  OR2_X1 U2451 ( .A1(n3796), .A2(n2130), .ZN(n2126) );
  NAND2_X1 U2452 ( .A1(n2139), .A2(n4526), .ZN(n2138) );
  NAND2_X1 U2453 ( .A1(n2140), .A2(n4577), .ZN(n2139) );
  NOR2_X1 U2454 ( .A1(n2140), .A2(n4577), .ZN(n4576) );
  XNOR2_X1 U2455 ( .A(n2062), .B(n3817), .ZN(n3822) );
  NAND2_X1 U2456 ( .A1(n4580), .A2(n2060), .ZN(n2062) );
  AND2_X1 U2457 ( .A1(n2572), .A2(n3657), .ZN(n2844) );
  INV_X2 U2458 ( .A(n4656), .ZN(n4658) );
  INV_X1 U2459 ( .A(n3268), .ZN(n2082) );
  AOI21_X1 U2460 ( .B1(n2196), .B2(n3337), .A(n2052), .ZN(n2195) );
  AND2_X1 U2461 ( .A1(n2780), .A2(n2901), .ZN(n2276) );
  INV_X1 U2462 ( .A(n2184), .ZN(n2182) );
  INV_X1 U2463 ( .A(n3456), .ZN(n3410) );
  NAND2_X1 U2464 ( .A1(n3772), .A2(n2135), .ZN(n2134) );
  NAND2_X1 U2465 ( .A1(n3767), .A2(REG2_REG_2__SCAN_IN), .ZN(n2135) );
  AOI21_X1 U2466 ( .B1(n3941), .B2(n2518), .A(n2047), .ZN(n2239) );
  INV_X1 U2467 ( .A(n2157), .ZN(n2155) );
  INV_X1 U2468 ( .A(n2254), .ZN(n2222) );
  INV_X1 U2469 ( .A(n3697), .ZN(n2168) );
  INV_X1 U2470 ( .A(n4092), .ZN(n2401) );
  AOI21_X1 U2471 ( .B1(n3637), .B2(n2355), .A(n2216), .ZN(n2215) );
  INV_X1 U2472 ( .A(n2364), .ZN(n2216) );
  OAI21_X1 U2473 ( .B1(n3671), .B2(n2574), .A(n2576), .ZN(n2800) );
  NOR2_X1 U2474 ( .A1(n4121), .A2(n4130), .ZN(n2104) );
  NAND2_X1 U2475 ( .A1(n2884), .A2(n2946), .ZN(n2091) );
  NAND2_X1 U2476 ( .A1(n2088), .A2(n2087), .ZN(n2242) );
  INV_X1 U2477 ( .A(n2243), .ZN(n2088) );
  NOR2_X1 U2478 ( .A1(n2386), .A2(IR_REG_9__SCAN_IN), .ZN(n2396) );
  INV_X1 U2479 ( .A(IR_REG_6__SCAN_IN), .ZN(n2348) );
  INV_X1 U2480 ( .A(IR_REG_2__SCAN_IN), .ZN(n2256) );
  NOR2_X1 U2481 ( .A1(n2247), .A2(n2201), .ZN(n2200) );
  INV_X1 U2482 ( .A(n2951), .ZN(n2201) );
  NAND2_X1 U2483 ( .A1(n3087), .A2(n2956), .ZN(n2204) );
  INV_X1 U2484 ( .A(n3086), .ZN(n3087) );
  NAND2_X1 U2485 ( .A1(n2200), .A2(n2074), .ZN(n2073) );
  INV_X1 U2486 ( .A(n2930), .ZN(n2074) );
  NOR2_X1 U2487 ( .A1(n3563), .A2(n2185), .ZN(n2184) );
  INV_X1 U2488 ( .A(n3483), .ZN(n2185) );
  INV_X1 U2489 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U2490 ( .A1(n2368), .A2(n2367), .ZN(n2380) );
  AND2_X1 U2491 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2319) );
  INV_X1 U2492 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4347) );
  AOI21_X1 U2493 ( .B1(n2189), .B2(n2192), .A(n2048), .ZN(n2188) );
  NAND2_X1 U2494 ( .A1(n2192), .A2(n2191), .ZN(n2190) );
  OR2_X1 U2495 ( .A1(n2480), .A2(n2479), .ZN(n2494) );
  NAND2_X1 U2496 ( .A1(n2512), .A2(REG3_REG_22__SCAN_IN), .ZN(n2519) );
  AND2_X1 U2497 ( .A1(n2504), .A2(REG3_REG_21__SCAN_IN), .ZN(n2512) );
  OAI22_X1 U2498 ( .A1(n2820), .A2(n3415), .B1(n2831), .B2(n3456), .ZN(n2821)
         );
  AOI21_X1 U2499 ( .B1(n2291), .B2(n3417), .A(n2822), .ZN(n2823) );
  NAND2_X1 U2500 ( .A1(n3499), .A2(n3498), .ZN(n3354) );
  NOR2_X1 U2501 ( .A1(n3499), .A2(n3498), .ZN(n3353) );
  AND2_X1 U2502 ( .A1(n2332), .A2(REG3_REG_6__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U2503 ( .A1(n2079), .A2(n2056), .ZN(n2186) );
  AND3_X1 U2504 ( .A1(n3593), .A2(n3592), .A3(n3591), .ZN(n3626) );
  XNOR2_X1 U2505 ( .A(n4479), .B(n2684), .ZN(n3762) );
  NAND2_X1 U2506 ( .A1(n3762), .A2(n3761), .ZN(n3760) );
  AND2_X1 U2507 ( .A1(n2109), .A2(n2108), .ZN(n3056) );
  NAND2_X1 U2508 ( .A1(n4474), .A2(REG2_REG_7__SCAN_IN), .ZN(n2108) );
  XNOR2_X1 U2509 ( .A(n3056), .B(n3055), .ZN(n3057) );
  NAND2_X1 U2510 ( .A1(n4506), .A2(REG1_REG_10__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U2511 ( .A1(n3050), .A2(n2210), .ZN(n3805) );
  AND2_X1 U2512 ( .A1(n3048), .A2(n2053), .ZN(n2210) );
  AND2_X1 U2513 ( .A1(n3794), .A2(n3807), .ZN(n2131) );
  OR2_X1 U2514 ( .A1(n3795), .A2(n3807), .ZN(n2130) );
  NAND2_X1 U2515 ( .A1(n2131), .A2(n3795), .ZN(n2129) );
  OR2_X1 U2516 ( .A1(n3807), .A2(n3794), .ZN(n2132) );
  NAND2_X1 U2517 ( .A1(n3805), .A2(n2053), .ZN(n3808) );
  OAI21_X1 U2518 ( .B1(n3877), .B2(n2051), .A(n2231), .ZN(n3297) );
  INV_X1 U2519 ( .A(n2232), .ZN(n2231) );
  OAI21_X1 U2520 ( .B1(n2042), .B2(n2233), .A(n2246), .ZN(n2232) );
  OR2_X1 U2521 ( .A1(n3613), .A2(n3618), .ZN(n3635) );
  INV_X1 U2522 ( .A(n4142), .ZN(n3906) );
  AND2_X1 U2523 ( .A1(n3917), .A2(n2597), .ZN(n3941) );
  OAI21_X1 U2524 ( .B1(n4048), .B2(n2156), .A(n2153), .ZN(n3953) );
  AOI21_X1 U2525 ( .B1(n2155), .B2(n3711), .A(n2154), .ZN(n2153) );
  INV_X1 U2526 ( .A(n3711), .ZN(n2156) );
  INV_X1 U2527 ( .A(n3605), .ZN(n2154) );
  NAND2_X1 U2528 ( .A1(n4048), .A2(n2157), .ZN(n3971) );
  NAND2_X1 U2529 ( .A1(n4048), .A2(n3596), .ZN(n4027) );
  AND2_X1 U2530 ( .A1(n3988), .A2(n3987), .ZN(n4035) );
  NOR3_X1 U2531 ( .A1(n4070), .A2(n4060), .A3(n4199), .ZN(n4052) );
  OR2_X1 U2532 ( .A1(n4069), .A2(n4068), .ZN(n4066) );
  AND2_X1 U2533 ( .A1(n3218), .A2(n3220), .ZN(n4092) );
  NAND2_X1 U2534 ( .A1(n3137), .A2(n3696), .ZN(n2584) );
  NAND2_X1 U2535 ( .A1(n2582), .A2(n3690), .ZN(n3070) );
  OAI21_X1 U2536 ( .B1(n2941), .B2(n2940), .A(n3688), .ZN(n2976) );
  NAND2_X1 U2537 ( .A1(n2579), .A2(n3680), .ZN(n3023) );
  AND2_X1 U2538 ( .A1(n3680), .A2(n3677), .ZN(n3639) );
  INV_X1 U2539 ( .A(n4640), .ZN(n3076) );
  NAND2_X1 U2540 ( .A1(n2637), .A2(n2668), .ZN(n2840) );
  AND2_X1 U2541 ( .A1(n3887), .A2(n2103), .ZN(n4112) );
  AND2_X1 U2542 ( .A1(n2029), .A2(n3616), .ZN(n2103) );
  NAND2_X1 U2543 ( .A1(n3887), .A2(n2104), .ZN(n3846) );
  AND2_X1 U2544 ( .A1(n3887), .A2(n3866), .ZN(n3864) );
  NAND2_X1 U2545 ( .A1(n2525), .A2(DATAI_25_), .ZN(n3889) );
  AND2_X1 U2546 ( .A1(n3900), .A2(n3889), .ZN(n3887) );
  NAND2_X1 U2547 ( .A1(n2525), .A2(DATAI_24_), .ZN(n3902) );
  NAND2_X1 U2548 ( .A1(n2601), .A2(n3632), .ZN(n3898) );
  NAND2_X1 U2549 ( .A1(n3957), .A2(n2030), .ZN(n3925) );
  INV_X1 U2550 ( .A(n3937), .ZN(n3943) );
  NAND2_X1 U2551 ( .A1(n3957), .A2(n2102), .ZN(n3945) );
  NAND2_X1 U2552 ( .A1(n3957), .A2(n3962), .ZN(n3958) );
  NOR2_X1 U2553 ( .A1(n3587), .A2(n2500), .ZN(n4170) );
  AND4_X1 U2554 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n4191)
         );
  NOR2_X1 U2555 ( .A1(n4070), .A2(n4199), .ZN(n4071) );
  INV_X1 U2556 ( .A(n2639), .ZN(n4208) );
  AND4_X1 U2557 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n4220)
         );
  NAND2_X1 U2558 ( .A1(n3133), .A2(n2045), .ZN(n4103) );
  NAND2_X1 U2559 ( .A1(n3133), .A2(n2100), .ZN(n4101) );
  INV_X1 U2560 ( .A(n3160), .ZN(n3175) );
  NOR2_X1 U2561 ( .A1(n3075), .A2(n3074), .ZN(n3135) );
  AND2_X1 U2562 ( .A1(n3135), .A2(n3138), .ZN(n3133) );
  NAND2_X1 U2563 ( .A1(n2090), .A2(n2089), .ZN(n3075) );
  AND3_X1 U2564 ( .A1(n2859), .A2(n3025), .A3(n2581), .ZN(n2089) );
  INV_X1 U2565 ( .A(n2091), .ZN(n2090) );
  AND2_X1 U2566 ( .A1(n4471), .A2(n2844), .ZN(n4200) );
  INV_X1 U2567 ( .A(n4651), .ZN(n4227) );
  NOR2_X1 U2568 ( .A1(n2092), .A2(n2867), .ZN(n3018) );
  NAND2_X1 U2569 ( .A1(n4093), .A2(n4641), .ZN(n4651) );
  OAI21_X1 U2570 ( .B1(n2315), .B2(n2280), .A(n2279), .ZN(n2797) );
  NAND2_X1 U2571 ( .A1(n2315), .A2(IR_REG_0__SCAN_IN), .ZN(n2279) );
  INV_X1 U2572 ( .A(n4648), .ZN(n4641) );
  XNOR2_X1 U2573 ( .A(n2559), .B(n2244), .ZN(n3657) );
  NAND2_X1 U2574 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2206) );
  AND3_X1 U2575 ( .A1(n2461), .A2(n2460), .A3(n2459), .ZN(n2462) );
  AND2_X1 U2576 ( .A1(n2407), .A2(n2400), .ZN(n3054) );
  OR3_X1 U2577 ( .A1(n2374), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2386) );
  INV_X1 U2578 ( .A(IR_REG_7__SCAN_IN), .ZN(n2350) );
  INV_X1 U2579 ( .A(IR_REG_3__SCAN_IN), .ZN(n2302) );
  AND4_X1 U2580 ( .A1(n2359), .A2(n2358), .A3(n2357), .A4(n2356), .ZN(n3152)
         );
  OAI21_X1 U2581 ( .B1(n2931), .B2(n2075), .A(n2072), .ZN(n3090) );
  INV_X1 U2582 ( .A(n2200), .ZN(n2075) );
  AND2_X1 U2583 ( .A1(n2073), .A2(n2202), .ZN(n2072) );
  NAND2_X1 U2584 ( .A1(n2204), .A2(n2203), .ZN(n2202) );
  NAND2_X1 U2585 ( .A1(n3090), .A2(n3089), .ZN(n3114) );
  NAND2_X1 U2586 ( .A1(n2078), .A2(n3562), .ZN(n3455) );
  NAND2_X1 U2587 ( .A1(n2186), .A2(n2184), .ZN(n2078) );
  AND2_X1 U2588 ( .A1(n2199), .A2(n3336), .ZN(n3430) );
  OR2_X1 U2589 ( .A1(n3338), .A2(n3337), .ZN(n2199) );
  AND2_X1 U2590 ( .A1(n3395), .A2(n2064), .ZN(n2063) );
  NAND2_X1 U2591 ( .A1(n3475), .A2(n2066), .ZN(n2065) );
  NAND2_X1 U2592 ( .A1(n2066), .A2(n2255), .ZN(n2064) );
  NAND2_X1 U2593 ( .A1(n3204), .A2(n3203), .ZN(n3258) );
  NAND2_X1 U2594 ( .A1(n2874), .A2(n2873), .ZN(n2875) );
  NAND2_X1 U2595 ( .A1(n2187), .A2(n2192), .ZN(n3444) );
  NAND2_X1 U2596 ( .A1(n2194), .A2(n2024), .ZN(n2187) );
  NAND2_X1 U2597 ( .A1(n2177), .A2(n3462), .ZN(n2176) );
  AOI22_X1 U2598 ( .A1(n2174), .A2(n2178), .B1(n2180), .B2(n3462), .ZN(n2173)
         );
  AND4_X1 U2599 ( .A1(n2347), .A2(n2346), .A3(n2345), .A4(n2344), .ZN(n3139)
         );
  INV_X1 U2600 ( .A(n2901), .ZN(n2896) );
  AND4_X1 U2601 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(n4239)
         );
  INV_X1 U2602 ( .A(n4195), .ZN(n4209) );
  OR2_X1 U2603 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  INV_X1 U2604 ( .A(n4172), .ZN(n3555) );
  INV_X1 U2605 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4346) );
  AND2_X1 U2606 ( .A1(n2067), .A2(n3382), .ZN(n3543) );
  AND2_X1 U2607 ( .A1(n2790), .A2(n2722), .ZN(n3545) );
  OAI21_X1 U2608 ( .B1(n2070), .B2(n2069), .A(n2068), .ZN(n3267) );
  AOI21_X1 U2609 ( .B1(n3203), .B2(n3173), .A(n2044), .ZN(n2068) );
  INV_X1 U2610 ( .A(n3203), .ZN(n2069) );
  AOI21_X1 U2611 ( .B1(n2194), .B2(n3354), .A(n3353), .ZN(n3554) );
  AND4_X1 U2612 ( .A1(n2324), .A2(n2323), .A3(n2322), .A4(n2321), .ZN(n2992)
         );
  NAND2_X1 U2613 ( .A1(n2952), .A2(n2951), .ZN(n2205) );
  OR2_X1 U2614 ( .A1(n2543), .A2(n2539), .ZN(n3868) );
  NAND2_X1 U2615 ( .A1(n2186), .A2(n3483), .ZN(n3565) );
  NAND2_X1 U2616 ( .A1(n2881), .A2(n2880), .ZN(n3580) );
  AND2_X1 U2617 ( .A1(n2957), .A2(n2727), .ZN(n3736) );
  INV_X1 U2618 ( .A(n3626), .ZN(n3828) );
  OAI211_X1 U2619 ( .C1(n3849), .C2(n2571), .A(n2546), .B(n2545), .ZN(n4131)
         );
  NAND2_X1 U2620 ( .A1(n2536), .A2(n2535), .ZN(n3746) );
  OAI211_X1 U2621 ( .C1(n3905), .C2(n2571), .A(n2529), .B(n2528), .ZN(n3747)
         );
  NAND4_X1 U2622 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n4162)
         );
  NAND4_X1 U2623 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n4171)
         );
  NAND4_X1 U2624 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n3997)
         );
  INV_X1 U2625 ( .A(n4000), .ZN(n4029) );
  INV_X1 U2626 ( .A(n4191), .ZN(n3748) );
  INV_X1 U2627 ( .A(n4031), .ZN(n4201) );
  INV_X1 U2628 ( .A(n4239), .ZN(n3749) );
  INV_X1 U2629 ( .A(n3139), .ZN(n3752) );
  OR2_X1 U2630 ( .A1(n2286), .A2(n3786), .ZN(n2300) );
  OR2_X1 U2631 ( .A1(n2286), .A2(n2673), .ZN(n2287) );
  AND2_X1 U2632 ( .A1(n2147), .A2(n2152), .ZN(n2146) );
  OR2_X1 U2633 ( .A1(n2708), .A2(n2665), .ZN(n3757) );
  OAI22_X1 U2634 ( .A1(n2122), .A2(n2112), .B1(n2124), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2114) );
  NAND2_X1 U2635 ( .A1(n2121), .A2(n2117), .ZN(n2116) );
  AOI22_X1 U2636 ( .A1(n2756), .A2(REG2_REG_4__SCAN_IN), .B1(n4477), .B2(n2678), .ZN(n2739) );
  NAND2_X1 U2637 ( .A1(n2690), .A2(n4477), .ZN(n2211) );
  NOR2_X1 U2638 ( .A1(n2696), .A2(n2106), .ZN(n2209) );
  AOI21_X1 U2639 ( .B1(n2702), .B2(REG2_REG_6__SCAN_IN), .A(n2058), .ZN(n2773)
         );
  XNOR2_X1 U2640 ( .A(n3808), .B(n2133), .ZN(n4540) );
  NAND2_X1 U2641 ( .A1(n4540), .A2(REG1_REG_14__SCAN_IN), .ZN(n4539) );
  NOR2_X1 U2642 ( .A1(n4535), .A2(n3798), .ZN(n4545) );
  OR2_X1 U2643 ( .A1(n3796), .A2(n3795), .ZN(n2127) );
  NAND2_X1 U2644 ( .A1(n3836), .A2(n4599), .ZN(n2099) );
  OAI21_X1 U2645 ( .B1(n3840), .B2(n4084), .A(n2095), .ZN(n2094) );
  NOR2_X1 U2646 ( .A1(n3838), .A2(n2096), .ZN(n2095) );
  NAND2_X1 U2647 ( .A1(n2230), .A2(n2249), .ZN(n3841) );
  NAND2_X1 U2648 ( .A1(n2235), .A2(n2042), .ZN(n2230) );
  NAND2_X1 U2649 ( .A1(n2164), .A2(n2603), .ZN(n3843) );
  INV_X1 U2650 ( .A(n4170), .ZN(n3981) );
  NAND2_X1 U2651 ( .A1(n2225), .A2(n2254), .ZN(n2224) );
  INV_X1 U2652 ( .A(n4084), .ZN(n4036) );
  NAND2_X1 U2653 ( .A1(n2556), .A2(n2489), .ZN(n3820) );
  OR2_X1 U2654 ( .A1(n2838), .A2(n2732), .ZN(n4588) );
  AND2_X1 U2655 ( .A1(n4020), .A2(n3076), .ZN(n4601) );
  INV_X1 U2656 ( .A(n4601), .ZN(n4106) );
  INV_X1 U2657 ( .A(n2797), .ZN(n2897) );
  AND2_X1 U2658 ( .A1(n3671), .A2(n3673), .ZN(n3633) );
  AND2_X1 U2659 ( .A1(n4591), .A2(n3820), .ZN(n4020) );
  AND2_X1 U2660 ( .A1(n4591), .A2(n4200), .ZN(n4059) );
  OR2_X1 U2661 ( .A1(n2644), .A2(n2840), .ZN(n4662) );
  NOR2_X1 U2662 ( .A1(n4656), .A2(n4640), .ZN(n4460) );
  NAND2_X1 U2663 ( .A1(n2663), .A2(n2729), .ZN(n4614) );
  XNOR2_X1 U2664 ( .A(n2616), .B(IR_REG_26__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U2665 ( .A1(n2031), .A2(IR_REG_31__SCAN_IN), .ZN(n2616) );
  XNOR2_X1 U2666 ( .A(n2611), .B(n2610), .ZN(n2653) );
  NAND2_X1 U2667 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2611) );
  XNOR2_X1 U2668 ( .A(n2560), .B(IR_REG_22__SCAN_IN), .ZN(n3739) );
  INV_X1 U2669 ( .A(n3657), .ZN(n4470) );
  AND2_X1 U2670 ( .A1(n2449), .A2(n2440), .ZN(n4625) );
  NAND2_X1 U2671 ( .A1(n2084), .A2(n2817), .ZN(n2829) );
  INV_X1 U2672 ( .A(n2136), .ZN(n4585) );
  OAI21_X1 U2673 ( .B1(n4576), .B2(n2138), .A(n2137), .ZN(n2136) );
  OAI21_X1 U2674 ( .B1(n2097), .B2(n4607), .A(n2093), .ZN(U3354) );
  AOI21_X1 U2675 ( .B1(n4261), .B2(n4601), .A(n2098), .ZN(n2097) );
  INV_X1 U2676 ( .A(n2094), .ZN(n2093) );
  NAND2_X1 U2677 ( .A1(n3837), .A2(n2099), .ZN(n2098) );
  OR2_X1 U2678 ( .A1(n3315), .A2(n4466), .ZN(n2642) );
  NAND2_X2 U2679 ( .A1(n2085), .A2(n2708), .ZN(n3421) );
  INV_X1 U2680 ( .A(n2355), .ZN(n2219) );
  NAND2_X1 U2681 ( .A1(n3750), .A2(n3160), .ZN(n2022) );
  AND2_X1 U2682 ( .A1(n2827), .A2(n2817), .ZN(n2023) );
  AND2_X1 U2683 ( .A1(n2057), .A2(n3354), .ZN(n2024) );
  NAND2_X1 U2684 ( .A1(n2070), .A2(n3171), .ZN(n3204) );
  NAND2_X1 U2685 ( .A1(n2224), .A2(n2223), .ZN(n3284) );
  AND2_X1 U2686 ( .A1(n3630), .A2(n3632), .ZN(n2025) );
  AND2_X1 U2687 ( .A1(n2165), .A2(n2025), .ZN(n2026) );
  OR2_X1 U2688 ( .A1(n4199), .A2(n4028), .ZN(n2027) );
  NOR2_X1 U2689 ( .A1(n3454), .A2(n2183), .ZN(n2028) );
  NAND2_X1 U2690 ( .A1(n2354), .A2(n2353), .ZN(n3081) );
  AND2_X1 U2691 ( .A1(n2104), .A2(n3465), .ZN(n2029) );
  AND2_X1 U2692 ( .A1(n2102), .A2(n3926), .ZN(n2030) );
  NAND2_X1 U2693 ( .A1(n2292), .A2(n2577), .ZN(n2806) );
  MUX2_X1 U2694 ( .A(n2274), .B(n2273), .S(IR_REG_27__SCAN_IN), .Z(n2315) );
  INV_X1 U2695 ( .A(n2315), .ZN(n2525) );
  INV_X1 U2696 ( .A(n3421), .ZN(n2871) );
  NAND3_X1 U2697 ( .A1(n2664), .A2(n2619), .A3(n4469), .ZN(n2708) );
  INV_X2 U2698 ( .A(n2525), .ZN(n3587) );
  NAND3_X1 U2699 ( .A1(n2161), .A2(n2162), .A3(n2160), .ZN(n2031) );
  XNOR2_X1 U2700 ( .A(n2206), .B(n2557), .ZN(n2562) );
  OR2_X1 U2701 ( .A1(n3174), .A2(n3208), .ZN(n2032) );
  NAND2_X1 U2702 ( .A1(n2208), .A2(n3039), .ZN(n2033) );
  INV_X1 U2703 ( .A(n2079), .ZN(n3482) );
  AND2_X1 U2704 ( .A1(n3940), .A2(n2518), .ZN(n2034) );
  AND2_X1 U2705 ( .A1(n2313), .A2(n2304), .ZN(n4478) );
  NAND3_X1 U2706 ( .A1(n2278), .A2(n2277), .A3(n2146), .ZN(n2712) );
  XNOR2_X1 U2707 ( .A(n3297), .B(n3635), .ZN(n3314) );
  OR2_X1 U2708 ( .A1(n2558), .A2(IR_REG_21__SCAN_IN), .ZN(n2035) );
  NAND2_X1 U2709 ( .A1(n4236), .A2(n3328), .ZN(n2036) );
  NAND2_X1 U2710 ( .A1(n2161), .A2(n2162), .ZN(n2558) );
  NAND2_X1 U2711 ( .A1(n2065), .A2(n2063), .ZN(n3436) );
  OR2_X1 U2712 ( .A1(n2558), .A2(n2242), .ZN(n2612) );
  AND2_X1 U2713 ( .A1(n3751), .A2(n3117), .ZN(n2037) );
  AND2_X1 U2714 ( .A1(n2134), .A2(n4478), .ZN(n2038) );
  INV_X1 U2715 ( .A(n3637), .ZN(n2353) );
  AND2_X1 U2716 ( .A1(n3691), .A2(n3693), .ZN(n3637) );
  INV_X1 U2717 ( .A(n2291), .ZN(n2820) );
  OR2_X1 U2718 ( .A1(n4096), .A2(n3197), .ZN(n2039) );
  AND2_X1 U2719 ( .A1(n2235), .A2(n2252), .ZN(n2040) );
  AND2_X1 U2720 ( .A1(n2401), .A2(n2032), .ZN(n2041) );
  AND2_X1 U2721 ( .A1(n2036), .A2(n3285), .ZN(n2223) );
  INV_X1 U2722 ( .A(n2118), .ZN(n2117) );
  NAND2_X1 U2723 ( .A1(n2123), .A2(REG2_REG_1__SCAN_IN), .ZN(n2118) );
  INV_X1 U2724 ( .A(n4475), .ZN(n2106) );
  NAND2_X1 U2725 ( .A1(n3269), .A2(n3268), .ZN(n3338) );
  INV_X1 U2726 ( .A(n3501), .ZN(n2194) );
  AND2_X1 U2727 ( .A1(n2162), .A2(n2228), .ZN(n2463) );
  NOR2_X1 U2728 ( .A1(n3344), .A2(n3343), .ZN(n3490) );
  NOR2_X1 U2729 ( .A1(n2234), .A2(n2542), .ZN(n2042) );
  INV_X1 U2730 ( .A(n3701), .ZN(n2171) );
  INV_X1 U2731 ( .A(IR_REG_21__SCAN_IN), .ZN(n2244) );
  INV_X1 U2732 ( .A(n4100), .ZN(n4088) );
  OR2_X1 U2733 ( .A1(n4131), .A2(n4121), .ZN(n2043) );
  AND3_X1 U2734 ( .A1(n2228), .A2(n2229), .A3(n2248), .ZN(n2421) );
  NAND2_X1 U2735 ( .A1(n2226), .A2(n2032), .ZN(n4089) );
  AND2_X1 U2736 ( .A1(n2224), .A2(n2036), .ZN(n3283) );
  AND2_X1 U2737 ( .A1(n3257), .A2(n3256), .ZN(n2044) );
  AND2_X1 U2738 ( .A1(n2100), .A2(n4088), .ZN(n2045) );
  AND2_X1 U2739 ( .A1(n4220), .A2(n4208), .ZN(n2046) );
  NOR2_X1 U2740 ( .A1(n4142), .A2(n3386), .ZN(n2047) );
  NOR2_X1 U2741 ( .A1(n3366), .A2(n3365), .ZN(n2048) );
  NOR2_X1 U2742 ( .A1(n3906), .A2(n3926), .ZN(n2049) );
  XOR2_X1 U2743 ( .A(n3339), .B(n3457), .Z(n2050) );
  INV_X1 U2744 ( .A(n2050), .ZN(n3340) );
  OR2_X1 U2745 ( .A1(n2233), .A2(n2253), .ZN(n2051) );
  OR2_X1 U2746 ( .A1(n3942), .A2(n3941), .ZN(n3940) );
  AND2_X1 U2747 ( .A1(n3340), .A2(n3428), .ZN(n2052) );
  INV_X1 U2748 ( .A(n2180), .ZN(n2179) );
  OAI21_X1 U2749 ( .B1(n3454), .B2(n2181), .A(n2245), .ZN(n2180) );
  INV_X1 U2750 ( .A(n3720), .ZN(n2165) );
  INV_X1 U2751 ( .A(n4060), .ZN(n4190) );
  NAND2_X1 U2752 ( .A1(n3133), .A2(n3175), .ZN(n3101) );
  INV_X1 U2753 ( .A(n3596), .ZN(n2158) );
  NOR2_X1 U2754 ( .A1(n3286), .A2(n2639), .ZN(n2640) );
  OR2_X1 U2755 ( .A1(n3806), .A2(n4229), .ZN(n2053) );
  INV_X1 U2756 ( .A(n3562), .ZN(n2183) );
  NAND2_X1 U2757 ( .A1(n2205), .A2(n2956), .ZN(n3085) );
  NAND2_X1 U2758 ( .A1(n3081), .A2(n2355), .ZN(n3136) );
  NAND2_X1 U2759 ( .A1(n2218), .A2(n2217), .ZN(n3100) );
  OR3_X1 U2760 ( .A1(n4070), .A2(n2027), .A3(n4060), .ZN(n2054) );
  NOR3_X1 U2761 ( .A1(n4070), .A2(n2027), .A3(n2055), .ZN(n2101) );
  OR2_X1 U2762 ( .A1(n4060), .A2(n4017), .ZN(n2055) );
  NAND2_X1 U2763 ( .A1(n3409), .A2(n3408), .ZN(n2056) );
  NAND2_X1 U2764 ( .A1(n3360), .A2(n3359), .ZN(n2057) );
  AND2_X1 U2765 ( .A1(n3977), .A2(n3981), .ZN(n3957) );
  NAND2_X1 U2766 ( .A1(n2806), .A2(n2293), .ZN(n2852) );
  AND2_X1 U2767 ( .A1(n2701), .A2(n4475), .ZN(n2058) );
  NAND2_X1 U2768 ( .A1(n2525), .A2(DATAI_21_), .ZN(n3962) );
  INV_X1 U2769 ( .A(n4121), .ZN(n3847) );
  NOR2_X1 U2770 ( .A1(n3587), .A2(n2547), .ZN(n4121) );
  INV_X1 U2771 ( .A(n4526), .ZN(n4575) );
  AND2_X1 U2772 ( .A1(n2681), .A2(n3737), .ZN(n4526) );
  INV_X1 U2773 ( .A(n2867), .ZN(n2884) );
  INV_X1 U2774 ( .A(n3926), .ZN(n3386) );
  NAND2_X1 U2775 ( .A1(n2525), .A2(DATAI_23_), .ZN(n3926) );
  OR2_X1 U2776 ( .A1(n2091), .A2(n2092), .ZN(n2059) );
  INV_X1 U2777 ( .A(IR_REG_25__SCAN_IN), .ZN(n2241) );
  OR2_X1 U2778 ( .A1(n4620), .A2(n3815), .ZN(n2060) );
  AOI21_X1 U2779 ( .B1(n4579), .B2(ADDR_REG_18__SCAN_IN), .A(n4578), .ZN(n2137) );
  NAND2_X1 U2780 ( .A1(n4494), .A2(n4495), .ZN(n4493) );
  NOR2_X1 U2781 ( .A1(n4560), .A2(n3813), .ZN(n4569) );
  NOR2_X1 U2782 ( .A1(n4570), .A2(n2207), .ZN(n4582) );
  INV_X1 U2783 ( .A(n2301), .ZN(n2229) );
  NAND2_X1 U2784 ( .A1(n2463), .A2(n2462), .ZN(n2473) );
  NAND2_X1 U2785 ( .A1(n2248), .A2(n2257), .ZN(n2071) );
  OAI21_X1 U2786 ( .B1(n3269), .B2(n2083), .A(n2080), .ZN(n3344) );
  NAND2_X1 U2787 ( .A1(n2023), .A2(n2084), .ZN(n2874) );
  NAND2_X1 U2788 ( .A1(n2086), .A2(n2241), .ZN(n2240) );
  NAND2_X1 U2789 ( .A1(n2859), .A2(n3025), .ZN(n2092) );
  NAND2_X1 U2790 ( .A1(n2884), .A2(n2859), .ZN(n3019) );
  INV_X1 U2791 ( .A(n2101), .ZN(n4018) );
  AOI22_X1 U2792 ( .A1(n2702), .A2(n2107), .B1(n2701), .B2(n2105), .ZN(n2109)
         );
  INV_X1 U2793 ( .A(n2109), .ZN(n2771) );
  NAND3_X1 U2794 ( .A1(n2115), .A2(n2113), .A3(n3759), .ZN(n3768) );
  NAND3_X1 U2795 ( .A1(n2114), .A2(REG2_REG_1__SCAN_IN), .A3(n2119), .ZN(n2113) );
  NAND3_X1 U2796 ( .A1(n2118), .A2(n2119), .A3(n2121), .ZN(n2115) );
  OAI211_X1 U2797 ( .C1(n2121), .C2(REG2_REG_1__SCAN_IN), .A(n2116), .B(n2119), 
        .ZN(n3758) );
  NAND2_X1 U2798 ( .A1(n2124), .A2(IR_REG_31__SCAN_IN), .ZN(n2122) );
  NAND2_X1 U2799 ( .A1(n3796), .A2(n2131), .ZN(n2125) );
  NAND2_X1 U2800 ( .A1(n2127), .A2(n3794), .ZN(n3797) );
  INV_X1 U2801 ( .A(n3807), .ZN(n2133) );
  XNOR2_X2 U2802 ( .A(n2290), .B(IR_REG_2__SCAN_IN), .ZN(n3767) );
  AND2_X2 U2803 ( .A1(n4468), .A2(n3312), .ZN(n2295) );
  INV_X1 U2804 ( .A(n2268), .ZN(n4468) );
  NAND2_X1 U2805 ( .A1(n2268), .A2(REG2_REG_0__SCAN_IN), .ZN(n2148) );
  NAND2_X1 U2806 ( .A1(n2149), .A2(n2268), .ZN(n2286) );
  INV_X1 U2807 ( .A(n2269), .ZN(n2149) );
  NOR2_X1 U2808 ( .A1(n2240), .A2(IR_REG_26__SCAN_IN), .ZN(n2159) );
  NAND3_X1 U2809 ( .A1(n2161), .A2(n2159), .A3(n2162), .ZN(n2271) );
  INV_X1 U2810 ( .A(n2240), .ZN(n2160) );
  INV_X1 U2811 ( .A(n3636), .ZN(n2577) );
  NAND2_X1 U2812 ( .A1(n2164), .A2(n2163), .ZN(n3845) );
  NAND2_X1 U2813 ( .A1(n2601), .A2(n2025), .ZN(n3880) );
  OAI21_X1 U2814 ( .B1(n3098), .B2(n2169), .A(n2166), .ZN(n4086) );
  OAI21_X1 U2815 ( .B1(n3098), .B2(n3097), .A(n3697), .ZN(n3123) );
  AOI21_X1 U2816 ( .B1(n3097), .B2(n3697), .A(n2171), .ZN(n2170) );
  NAND2_X1 U2817 ( .A1(n3482), .A2(n2174), .ZN(n2172) );
  OAI211_X1 U2818 ( .C1(n3482), .C2(n2176), .A(n2173), .B(n2172), .ZN(n3463)
         );
  OAI21_X1 U2819 ( .B1(n2194), .B2(n2190), .A(n2188), .ZN(n3518) );
  INV_X1 U2820 ( .A(n2247), .ZN(n2203) );
  INV_X2 U2821 ( .A(n3459), .ZN(n3417) );
  NAND2_X1 U2822 ( .A1(n2212), .A2(n2305), .ZN(n2213) );
  INV_X1 U2823 ( .A(n2293), .ZN(n2212) );
  NAND3_X1 U2824 ( .A1(n2214), .A2(n2306), .A3(n2213), .ZN(n3027) );
  NAND3_X1 U2825 ( .A1(n2292), .A2(n2305), .A3(n2577), .ZN(n2214) );
  NAND2_X1 U2826 ( .A1(n2354), .A2(n2215), .ZN(n2218) );
  NAND2_X1 U2827 ( .A1(n3217), .A2(n2223), .ZN(n2220) );
  NAND2_X1 U2828 ( .A1(n2220), .A2(n2221), .ZN(n4065) );
  NAND2_X1 U2829 ( .A1(n2226), .A2(n2041), .ZN(n4090) );
  NAND2_X1 U2830 ( .A1(n2378), .A2(n2377), .ZN(n3129) );
  AND2_X1 U2831 ( .A1(n2377), .A2(n2039), .ZN(n2227) );
  NAND2_X1 U2832 ( .A1(n2229), .A2(n2248), .ZN(n2325) );
  NOR2_X1 U2833 ( .A1(n2558), .A2(n2243), .ZN(n2609) );
  NAND2_X1 U2834 ( .A1(n2294), .A2(REG1_REG_0__SCAN_IN), .ZN(n2278) );
  NAND2_X1 U2835 ( .A1(n3344), .A2(n3343), .ZN(n3489) );
  OAI22_X1 U2836 ( .A1(n2783), .A2(n3415), .B1(n2896), .B2(n3456), .ZN(n2782)
         );
  AND4_X1 U2837 ( .A1(n2275), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n2783)
         );
  INV_X1 U2838 ( .A(n3940), .ZN(n4155) );
  NAND2_X1 U2839 ( .A1(n2296), .A2(REG0_REG_1__SCAN_IN), .ZN(n2780) );
  AND2_X2 U2840 ( .A1(n2269), .A2(n2268), .ZN(n2296) );
  OR2_X1 U2841 ( .A1(n3453), .A2(n3452), .ZN(n2245) );
  OR2_X1 U2842 ( .A1(n3869), .A2(n3847), .ZN(n2246) );
  AND2_X1 U2843 ( .A1(n2964), .A2(n2963), .ZN(n2247) );
  OR2_X1 U2844 ( .A1(n4122), .A2(n4130), .ZN(n2249) );
  AND2_X1 U2845 ( .A1(n3747), .A2(n4141), .ZN(n2250) );
  AND2_X1 U2846 ( .A1(n4209), .A2(n4080), .ZN(n2251) );
  OR2_X1 U2847 ( .A1(n4145), .A2(n3889), .ZN(n2252) );
  AND2_X1 U2848 ( .A1(n4145), .A2(n3889), .ZN(n2253) );
  OR2_X1 U2849 ( .A1(n4236), .A2(n3328), .ZN(n2254) );
  NOR2_X1 U2850 ( .A1(n3587), .A2(n2555), .ZN(n3295) );
  AND2_X1 U2851 ( .A1(n3473), .A2(n3472), .ZN(n2255) );
  NOR2_X1 U2852 ( .A1(n3850), .A2(n3866), .ZN(n2542) );
  NAND2_X1 U2853 ( .A1(n3921), .A2(n3902), .ZN(n2530) );
  NAND2_X1 U2854 ( .A1(n3381), .A2(n3380), .ZN(n3382) );
  INV_X1 U2855 ( .A(IR_REG_30__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2856 ( .A1(n4172), .A2(n3361), .ZN(n2490) );
  OR2_X1 U2857 ( .A1(n3753), .A2(n2990), .ZN(n2339) );
  NAND2_X1 U2858 ( .A1(n4162), .A2(n3943), .ZN(n2518) );
  OAI21_X1 U2859 ( .B1(n2975), .B2(n2340), .A(n2339), .ZN(n3082) );
  INV_X1 U2860 ( .A(IR_REG_28__SCAN_IN), .ZN(n2272) );
  AND2_X1 U2861 ( .A1(n3437), .A2(n3438), .ZN(n3395) );
  AND2_X1 U2862 ( .A1(n2443), .A2(n2442), .ZN(n2453) );
  INV_X1 U2863 ( .A(n4219), .ZN(n4235) );
  AND2_X1 U2864 ( .A1(n3739), .A2(n4470), .ZN(n2719) );
  AND2_X1 U2865 ( .A1(n2319), .A2(REG3_REG_5__SCAN_IN), .ZN(n2332) );
  OR2_X1 U2866 ( .A1(n2415), .A2(n2412), .ZN(n2424) );
  OR2_X1 U2867 ( .A1(n2388), .A2(n3260), .ZN(n2415) );
  NAND2_X1 U2868 ( .A1(n2453), .A2(REG3_REG_17__SCAN_IN), .ZN(n2480) );
  INV_X1 U2869 ( .A(n4131), .ZN(n3869) );
  AND3_X1 U2870 ( .A1(n2717), .A2(n2842), .A3(n2839), .ZN(n2790) );
  AND2_X1 U2871 ( .A1(n2538), .A2(n2537), .ZN(n2543) );
  INV_X1 U2872 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3260) );
  INV_X1 U2873 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4371) );
  INV_X1 U2874 ( .A(n3666), .ZN(n3842) );
  INV_X1 U2875 ( .A(n4049), .ZN(n2451) );
  INV_X1 U2876 ( .A(n4200), .ZN(n4232) );
  INV_X1 U2877 ( .A(n3902), .ZN(n4141) );
  AND2_X1 U2878 ( .A1(n3710), .A2(n3596), .ZN(n4049) );
  INV_X1 U2879 ( .A(n3328), .ZN(n4218) );
  NAND2_X1 U2880 ( .A1(n2750), .A2(n2719), .ZN(n4238) );
  NAND2_X1 U2881 ( .A1(n2788), .A2(n2719), .ZN(n4219) );
  INV_X1 U2882 ( .A(DATAI_0_), .ZN(n2280) );
  INV_X1 U2883 ( .A(IR_REG_24__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U2884 ( .A1(n2341), .A2(REG3_REG_7__SCAN_IN), .ZN(n2368) );
  AND2_X1 U2885 ( .A1(n3835), .A2(n2549), .ZN(n3469) );
  INV_X1 U2886 ( .A(n3567), .ZN(n3579) );
  AND2_X1 U2887 ( .A1(n2554), .A2(n2553), .ZN(n4124) );
  AND4_X1 U2888 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n4000)
         );
  NOR2_X1 U2889 ( .A1(n3587), .A2(n2670), .ZN(n2680) );
  INV_X1 U2890 ( .A(n3616), .ZN(n3839) );
  INV_X1 U2891 ( .A(n4238), .ZN(n4224) );
  INV_X1 U2892 ( .A(n4607), .ZN(n4591) );
  NOR2_X1 U2893 ( .A1(n4662), .A2(n4640), .ZN(n4246) );
  NAND2_X1 U2894 ( .A1(n2525), .A2(DATAI_26_), .ZN(n3866) );
  INV_X1 U2895 ( .A(n3361), .ZN(n4002) );
  INV_X1 U2896 ( .A(n4199), .ZN(n4080) );
  AND2_X1 U2897 ( .A1(n2562), .A2(n2563), .ZN(n4648) );
  INV_X1 U2898 ( .A(n2838), .ZN(n2729) );
  INV_X1 U2899 ( .A(n3545), .ZN(n3583) );
  NAND4_X1 U2900 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n4142)
         );
  INV_X1 U2901 ( .A(n4220), .ZN(n4074) );
  NAND2_X1 U2902 ( .A1(n2681), .A2(n2788), .ZN(n4586) );
  NAND2_X1 U2903 ( .A1(n3102), .A2(n2974), .ZN(n4084) );
  OR2_X1 U2904 ( .A1(n3315), .A2(n4251), .ZN(n2647) );
  INV_X1 U2905 ( .A(n4246), .ZN(n4251) );
  INV_X2 U2906 ( .A(n4662), .ZN(n4665) );
  INV_X1 U2907 ( .A(n4460), .ZN(n4466) );
  OR2_X1 U2908 ( .A1(n2644), .A2(n2717), .ZN(n4656) );
  INV_X1 U2909 ( .A(n4614), .ZN(n4616) );
  INV_X1 U2910 ( .A(D_REG_0__SCAN_IN), .ZN(n4373) );
  AND2_X1 U2911 ( .A1(n2877), .A2(STATE_REG_SCAN_IN), .ZN(n4617) );
  INV_X1 U2912 ( .A(n3054), .ZN(n4631) );
  AND2_X1 U2913 ( .A1(n2360), .A2(n2352), .ZN(n4474) );
  INV_X1 U2914 ( .A(n3757), .ZN(U4043) );
  NAND2_X1 U2915 ( .A1(n2289), .A2(n2256), .ZN(n2301) );
  NAND2_X1 U2916 ( .A1(n2564), .A2(n2272), .ZN(n2264) );
  NOR2_X2 U2917 ( .A1(n2264), .A2(IR_REG_29__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2918 ( .A1(n2264), .A2(IR_REG_31__SCAN_IN), .ZN(n2265) );
  INV_X1 U2919 ( .A(n2266), .ZN(n2660) );
  INV_X1 U2920 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2674) );
  OR2_X1 U2921 ( .A1(n2286), .A2(n2674), .ZN(n2275) );
  NAND2_X1 U2922 ( .A1(n2294), .A2(REG1_REG_1__SCAN_IN), .ZN(n2778) );
  XNOR2_X1 U2923 ( .A(n2270), .B(IR_REG_30__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U2924 ( .A1(n2295), .A2(REG3_REG_1__SCAN_IN), .ZN(n2779) );
  NAND4_X1 U2925 ( .A1(n2275), .A2(n2778), .A3(n2780), .A4(n2779), .ZN(n2281)
         );
  NAND2_X1 U2926 ( .A1(n2271), .A2(IR_REG_31__SCAN_IN), .ZN(n2656) );
  NOR2_X1 U2927 ( .A1(n2656), .A2(n2272), .ZN(n2273) );
  MUX2_X1 U2928 ( .A(DATAI_1_), .B(n4479), .S(n2315), .Z(n2901) );
  NAND2_X1 U2929 ( .A1(n2281), .A2(n2896), .ZN(n3672) );
  NAND4_X1 U2930 ( .A1(n2275), .A2(n2779), .A3(n2276), .A4(n2778), .ZN(n2576)
         );
  NAND2_X1 U2931 ( .A1(n3672), .A2(n2576), .ZN(n2574) );
  INV_X1 U2932 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U2933 ( .A1(n2296), .A2(REG0_REG_0__SCAN_IN), .ZN(n2277) );
  AND2_X1 U2934 ( .A1(n2712), .A2(n2797), .ZN(n2899) );
  NAND2_X1 U2935 ( .A1(n2574), .A2(n2899), .ZN(n2898) );
  NAND2_X1 U2936 ( .A1(n2281), .A2(n2901), .ZN(n2282) );
  NAND2_X1 U2937 ( .A1(n2898), .A2(n2282), .ZN(n2807) );
  INV_X1 U2938 ( .A(n2807), .ZN(n2292) );
  NAND2_X1 U2939 ( .A1(n2294), .A2(REG1_REG_2__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2940 ( .A1(n2296), .A2(REG0_REG_2__SCAN_IN), .ZN(n2284) );
  NAND2_X1 U2941 ( .A1(n2295), .A2(REG3_REG_2__SCAN_IN), .ZN(n2283) );
  INV_X1 U2942 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2673) );
  OR2_X1 U2943 ( .A1(n2289), .A2(n2659), .ZN(n2290) );
  MUX2_X1 U2944 ( .A(DATAI_2_), .B(n3767), .S(n2315), .Z(n2812) );
  INV_X1 U2945 ( .A(n2812), .ZN(n2831) );
  NAND2_X1 U2946 ( .A1(n2820), .A2(n2812), .ZN(n3675) );
  NAND2_X1 U2947 ( .A1(n2820), .A2(n2831), .ZN(n2293) );
  INV_X1 U2948 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U2949 ( .A1(n2294), .A2(REG1_REG_3__SCAN_IN), .ZN(n2299) );
  INV_X1 U2950 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U2951 ( .A1(n2318), .A2(n2882), .ZN(n2298) );
  NAND2_X1 U2952 ( .A1(n2296), .A2(REG0_REG_3__SCAN_IN), .ZN(n2297) );
  NAND2_X1 U2953 ( .A1(n2301), .A2(IR_REG_31__SCAN_IN), .ZN(n2303) );
  NAND2_X1 U2954 ( .A1(n2303), .A2(n2302), .ZN(n2313) );
  OR2_X1 U2955 ( .A1(n2303), .A2(n2302), .ZN(n2304) );
  MUX2_X1 U2956 ( .A(DATAI_3_), .B(n4478), .S(n3587), .Z(n2867) );
  NAND2_X1 U2957 ( .A1(n3756), .A2(n2867), .ZN(n2305) );
  INV_X1 U2958 ( .A(n3756), .ZN(n2578) );
  NAND2_X1 U2959 ( .A1(n2578), .A2(n2884), .ZN(n2306) );
  INV_X1 U2960 ( .A(n3027), .ZN(n2316) );
  NAND2_X1 U2961 ( .A1(n2294), .A2(REG1_REG_4__SCAN_IN), .ZN(n2312) );
  NOR2_X1 U2962 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2307) );
  NOR2_X1 U2963 ( .A1(n2319), .A2(n2307), .ZN(n2912) );
  NAND2_X1 U2964 ( .A1(n2318), .A2(n2912), .ZN(n2311) );
  NAND2_X1 U2965 ( .A1(n2296), .A2(REG0_REG_4__SCAN_IN), .ZN(n2310) );
  INV_X1 U2966 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2308) );
  OR2_X1 U2967 ( .A1(n2286), .A2(n2308), .ZN(n2309) );
  NAND2_X1 U2968 ( .A1(n2313), .A2(IR_REG_31__SCAN_IN), .ZN(n2314) );
  XNOR2_X1 U2969 ( .A(n2314), .B(IR_REG_4__SCAN_IN), .ZN(n4477) );
  MUX2_X1 U2970 ( .A(DATAI_4_), .B(n4477), .S(n3587), .Z(n3020) );
  INV_X1 U2971 ( .A(n3020), .ZN(n3025) );
  NAND2_X1 U2972 ( .A1(n2916), .A2(n3020), .ZN(n3681) );
  NAND2_X1 U2973 ( .A1(n2316), .A2(n3022), .ZN(n3026) );
  NAND2_X1 U2974 ( .A1(n3755), .A2(n3020), .ZN(n2317) );
  NAND2_X1 U2975 ( .A1(n3026), .A2(n2317), .ZN(n2939) );
  NAND2_X1 U2976 ( .A1(n3588), .A2(REG1_REG_5__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2977 ( .A1(n3589), .A2(REG0_REG_5__SCAN_IN), .ZN(n2323) );
  NOR2_X1 U2978 ( .A1(n2319), .A2(REG3_REG_5__SCAN_IN), .ZN(n2320) );
  NOR2_X1 U2979 ( .A1(n2332), .A2(n2320), .ZN(n3005) );
  NAND2_X1 U2980 ( .A1(n2318), .A2(n3005), .ZN(n2322) );
  OR2_X1 U2981 ( .A1(n3590), .A2(n3007), .ZN(n2321) );
  INV_X1 U2982 ( .A(DATAI_5_), .ZN(n2328) );
  NAND2_X1 U2983 ( .A1(n2325), .A2(IR_REG_31__SCAN_IN), .ZN(n2327) );
  INV_X1 U2984 ( .A(IR_REG_5__SCAN_IN), .ZN(n2326) );
  XNOR2_X1 U2985 ( .A(n2327), .B(n2326), .ZN(n2745) );
  MUX2_X1 U2986 ( .A(n2328), .B(n2745), .S(n3587), .Z(n2946) );
  NAND2_X1 U2987 ( .A1(n2992), .A2(n2946), .ZN(n2329) );
  NAND2_X1 U2988 ( .A1(n2939), .A2(n2329), .ZN(n2331) );
  INV_X1 U2989 ( .A(n2992), .ZN(n3754) );
  INV_X1 U2990 ( .A(n2946), .ZN(n3009) );
  NAND2_X1 U2991 ( .A1(n3754), .A2(n3009), .ZN(n2330) );
  NAND2_X1 U2992 ( .A1(n2331), .A2(n2330), .ZN(n2975) );
  INV_X1 U2993 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2980) );
  OR2_X1 U2994 ( .A1(n3590), .A2(n2980), .ZN(n2337) );
  NAND2_X1 U2995 ( .A1(n3588), .A2(REG1_REG_6__SCAN_IN), .ZN(n2336) );
  NOR2_X1 U2996 ( .A1(n2332), .A2(REG3_REG_6__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2997 ( .A1(n2341), .A2(n2333), .ZN(n2978) );
  NAND2_X1 U2998 ( .A1(n2318), .A2(n2978), .ZN(n2335) );
  NAND2_X1 U2999 ( .A1(n3589), .A2(REG0_REG_6__SCAN_IN), .ZN(n2334) );
  NAND4_X1 U3000 ( .A1(n2337), .A2(n2336), .A3(n2335), .A4(n2334), .ZN(n3753)
         );
  NOR2_X1 U3001 ( .A1(n2325), .A2(IR_REG_5__SCAN_IN), .ZN(n2349) );
  OR2_X1 U3002 ( .A1(n2349), .A2(n2659), .ZN(n2338) );
  XNOR2_X1 U3003 ( .A(n2338), .B(IR_REG_6__SCAN_IN), .ZN(n4475) );
  MUX2_X1 U3004 ( .A(DATAI_6_), .B(n4475), .S(n3587), .Z(n2990) );
  AND2_X1 U3005 ( .A1(n3753), .A2(n2990), .ZN(n2340) );
  INV_X1 U3006 ( .A(n3082), .ZN(n2354) );
  NAND2_X1 U3007 ( .A1(n3588), .A2(REG1_REG_7__SCAN_IN), .ZN(n2347) );
  OAI21_X1 U3008 ( .B1(n2341), .B2(REG3_REG_7__SCAN_IN), .A(n2368), .ZN(n3096)
         );
  INV_X1 U3009 ( .A(n3096), .ZN(n2342) );
  NAND2_X1 U3010 ( .A1(n2318), .A2(n2342), .ZN(n2346) );
  NAND2_X1 U3011 ( .A1(n3589), .A2(REG0_REG_7__SCAN_IN), .ZN(n2345) );
  INV_X1 U3012 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2343) );
  OR2_X1 U3013 ( .A1(n3590), .A2(n2343), .ZN(n2344) );
  NAND2_X1 U3014 ( .A1(n2349), .A2(n2348), .ZN(n2374) );
  NAND2_X1 U3015 ( .A1(n2374), .A2(IR_REG_31__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3016 ( .A1(n2351), .A2(n2350), .ZN(n2360) );
  OR2_X1 U3017 ( .A1(n2351), .A2(n2350), .ZN(n2352) );
  MUX2_X1 U3018 ( .A(DATAI_7_), .B(n4474), .S(n3587), .Z(n3074) );
  NAND2_X1 U3019 ( .A1(n3139), .A2(n3074), .ZN(n3691) );
  INV_X1 U3020 ( .A(n3074), .ZN(n3091) );
  NAND2_X1 U3021 ( .A1(n3752), .A2(n3091), .ZN(n3693) );
  NAND2_X1 U3022 ( .A1(n3752), .A2(n3074), .ZN(n2355) );
  NAND2_X1 U3023 ( .A1(n3588), .A2(REG1_REG_8__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3024 ( .A1(n3589), .A2(REG0_REG_8__SCAN_IN), .ZN(n2358) );
  XNOR2_X1 U3025 ( .A(n2368), .B(REG3_REG_8__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U3026 ( .A1(n2318), .A2(n4587), .ZN(n2357) );
  INV_X1 U3027 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4590) );
  OR2_X1 U3028 ( .A1(n3590), .A2(n4590), .ZN(n2356) );
  INV_X1 U3029 ( .A(DATAI_8_), .ZN(n2363) );
  NAND2_X1 U3030 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  INV_X1 U3031 ( .A(IR_REG_8__SCAN_IN), .ZN(n2361) );
  XNOR2_X1 U3032 ( .A(n2362), .B(n2361), .ZN(n3055) );
  MUX2_X1 U3033 ( .A(n2363), .B(n3055), .S(n3587), .Z(n3138) );
  NAND2_X1 U3034 ( .A1(n3152), .A2(n3138), .ZN(n2364) );
  INV_X1 U3035 ( .A(n3152), .ZN(n3751) );
  INV_X1 U3036 ( .A(n3138), .ZN(n3117) );
  INV_X1 U3037 ( .A(n3100), .ZN(n2376) );
  INV_X1 U3038 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2365) );
  OR2_X1 U3039 ( .A1(n3590), .A2(n2365), .ZN(n2373) );
  NAND2_X1 U3040 ( .A1(n3588), .A2(REG1_REG_9__SCAN_IN), .ZN(n2372) );
  INV_X1 U3041 ( .A(n2368), .ZN(n2366) );
  AOI21_X1 U3042 ( .B1(n2366), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3043 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2367) );
  OR2_X1 U3044 ( .A1(n2369), .A2(n2380), .ZN(n3103) );
  INV_X1 U3045 ( .A(n3103), .ZN(n3177) );
  NAND2_X1 U3046 ( .A1(n2318), .A2(n3177), .ZN(n2371) );
  NAND2_X1 U3047 ( .A1(n3589), .A2(REG0_REG_9__SCAN_IN), .ZN(n2370) );
  NAND4_X1 U3048 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2370), .ZN(n3750)
         );
  NAND2_X1 U3049 ( .A1(n2386), .A2(IR_REG_31__SCAN_IN), .ZN(n2375) );
  XNOR2_X1 U3050 ( .A(n2375), .B(IR_REG_9__SCAN_IN), .ZN(n4634) );
  MUX2_X1 U3051 ( .A(DATAI_9_), .B(n4634), .S(n3587), .Z(n3160) );
  NAND2_X1 U3052 ( .A1(n2376), .A2(n2022), .ZN(n2378) );
  INV_X1 U3053 ( .A(n3750), .ZN(n2585) );
  NAND2_X1 U3054 ( .A1(n2585), .A2(n3175), .ZN(n2377) );
  INV_X1 U3055 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2379) );
  OR2_X1 U3056 ( .A1(n3590), .A2(n2379), .ZN(n2385) );
  NAND2_X1 U3057 ( .A1(n3588), .A2(REG1_REG_10__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U3058 ( .A1(n3589), .A2(REG0_REG_10__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3059 ( .A1(n2380), .A2(REG3_REG_10__SCAN_IN), .ZN(n2388) );
  OR2_X1 U3060 ( .A1(n2380), .A2(REG3_REG_10__SCAN_IN), .ZN(n2381) );
  AND2_X1 U3061 ( .A1(n2388), .A2(n2381), .ZN(n3194) );
  NAND2_X1 U3062 ( .A1(n2318), .A2(n3194), .ZN(n2382) );
  NAND4_X1 U3063 ( .A1(n2385), .A2(n2384), .A3(n2383), .A4(n2382), .ZN(n4096)
         );
  OR2_X1 U3064 ( .A1(n2396), .A2(n2659), .ZN(n2387) );
  XNOR2_X1 U3065 ( .A(n2387), .B(IR_REG_10__SCAN_IN), .ZN(n3059) );
  MUX2_X1 U3066 ( .A(DATAI_10_), .B(n3059), .S(n3587), .Z(n3197) );
  INV_X1 U3067 ( .A(n4096), .ZN(n3174) );
  INV_X1 U3068 ( .A(n3197), .ZN(n3208) );
  NAND2_X1 U3069 ( .A1(n3588), .A2(REG1_REG_11__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3070 ( .A1(n3589), .A2(REG0_REG_11__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3071 ( .A1(n2388), .A2(n3260), .ZN(n2389) );
  AND2_X1 U3072 ( .A1(n2415), .A2(n2389), .ZN(n4104) );
  NAND2_X1 U3073 ( .A1(n2318), .A2(n4104), .ZN(n2392) );
  INV_X1 U3074 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2390) );
  OR2_X1 U3075 ( .A1(n3590), .A2(n2390), .ZN(n2391) );
  INV_X1 U3076 ( .A(IR_REG_10__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3077 ( .A1(n2396), .A2(n2395), .ZN(n2397) );
  NAND2_X1 U3078 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  INV_X1 U3079 ( .A(IR_REG_11__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U3080 ( .A1(n2399), .A2(n2398), .ZN(n2407) );
  OR2_X1 U3081 ( .A1(n2399), .A2(n2398), .ZN(n2400) );
  MUX2_X1 U3082 ( .A(DATAI_11_), .B(n3054), .S(n3587), .Z(n4100) );
  NAND2_X1 U3083 ( .A1(n4239), .A2(n4100), .ZN(n3218) );
  NAND2_X1 U3084 ( .A1(n3749), .A2(n4088), .ZN(n3220) );
  NAND2_X1 U3085 ( .A1(n4239), .A2(n4088), .ZN(n2402) );
  NAND2_X1 U3086 ( .A1(n4090), .A2(n2402), .ZN(n3232) );
  INV_X1 U3087 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3238) );
  OR2_X1 U3088 ( .A1(n3590), .A2(n3238), .ZN(n2406) );
  NAND2_X1 U3089 ( .A1(n3588), .A2(REG1_REG_12__SCAN_IN), .ZN(n2405) );
  XNOR2_X1 U3090 ( .A(n2415), .B(REG3_REG_12__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U3091 ( .A1(n2318), .A2(n3280), .ZN(n2404) );
  NAND2_X1 U3092 ( .A1(n3589), .A2(REG0_REG_12__SCAN_IN), .ZN(n2403) );
  NAND4_X1 U3093 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(n4223)
         );
  NAND2_X1 U3094 ( .A1(n2407), .A2(IR_REG_31__SCAN_IN), .ZN(n2408) );
  XNOR2_X1 U3095 ( .A(n2408), .B(IR_REG_12__SCAN_IN), .ZN(n3063) );
  MUX2_X1 U3096 ( .A(DATAI_12_), .B(n3063), .S(n3587), .Z(n3276) );
  NAND2_X1 U3097 ( .A1(n4223), .A2(n3276), .ZN(n2409) );
  NAND2_X1 U3098 ( .A1(n3232), .A2(n2409), .ZN(n2411) );
  INV_X1 U3099 ( .A(n4223), .ZN(n3261) );
  INV_X1 U3100 ( .A(n3276), .ZN(n4233) );
  NAND2_X1 U3101 ( .A1(n3261), .A2(n4233), .ZN(n2410) );
  NAND2_X1 U3102 ( .A1(n2411), .A2(n2410), .ZN(n3217) );
  INV_X1 U3103 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4398) );
  OR2_X1 U3104 ( .A1(n3590), .A2(n4398), .ZN(n2420) );
  NAND2_X1 U3105 ( .A1(n3588), .A2(REG1_REG_13__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3106 ( .A1(n3589), .A2(REG0_REG_13__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3107 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2412) );
  INV_X1 U3108 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2414) );
  INV_X1 U3109 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2413) );
  OAI21_X1 U3110 ( .B1(n2415), .B2(n2414), .A(n2413), .ZN(n2416) );
  AND2_X1 U3111 ( .A1(n2424), .A2(n2416), .ZN(n3538) );
  NAND2_X1 U3112 ( .A1(n2318), .A2(n3538), .ZN(n2417) );
  NOR2_X1 U3113 ( .A1(n2421), .A2(n2659), .ZN(n2422) );
  MUX2_X1 U3114 ( .A(n2659), .B(n2422), .S(IR_REG_13__SCAN_IN), .Z(n2423) );
  OR2_X1 U3115 ( .A1(n2423), .A2(n2463), .ZN(n3806) );
  INV_X1 U3116 ( .A(n3806), .ZN(n4473) );
  MUX2_X1 U3117 ( .A(DATAI_13_), .B(n4473), .S(n3587), .Z(n3328) );
  NAND2_X1 U3118 ( .A1(n3588), .A2(REG1_REG_14__SCAN_IN), .ZN(n2430) );
  AND2_X1 U3119 ( .A1(n2424), .A2(n4371), .ZN(n2425) );
  NOR2_X1 U3120 ( .A1(n2443), .A2(n2425), .ZN(n3432) );
  NAND2_X1 U3121 ( .A1(n2318), .A2(n3432), .ZN(n2429) );
  NAND2_X1 U3122 ( .A1(n3589), .A2(REG0_REG_14__SCAN_IN), .ZN(n2428) );
  INV_X1 U3123 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2426) );
  OR2_X1 U3124 ( .A1(n3590), .A2(n2426), .ZN(n2427) );
  OR2_X1 U3125 ( .A1(n2463), .A2(n2659), .ZN(n2431) );
  XNOR2_X1 U3126 ( .A(n2431), .B(IR_REG_14__SCAN_IN), .ZN(n3807) );
  MUX2_X1 U3127 ( .A(DATAI_14_), .B(n3807), .S(n3587), .Z(n2639) );
  NAND2_X1 U3128 ( .A1(n4220), .A2(n2639), .ZN(n3594) );
  NAND2_X1 U3129 ( .A1(n4074), .A2(n4208), .ZN(n3602) );
  NAND2_X1 U3130 ( .A1(n3594), .A2(n3602), .ZN(n3285) );
  INV_X1 U3131 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2432) );
  OR2_X1 U3132 ( .A1(n3590), .A2(n2432), .ZN(n2437) );
  NAND2_X1 U3133 ( .A1(n3588), .A2(REG1_REG_15__SCAN_IN), .ZN(n2436) );
  INV_X1 U3134 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2433) );
  XNOR2_X1 U3135 ( .A(n2443), .B(n2433), .ZN(n4076) );
  NAND2_X1 U3136 ( .A1(n2318), .A2(n4076), .ZN(n2435) );
  NAND2_X1 U3137 ( .A1(n3589), .A2(REG0_REG_15__SCAN_IN), .ZN(n2434) );
  NAND4_X1 U3138 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2434), .ZN(n4195)
         );
  NAND2_X1 U3139 ( .A1(n2463), .A2(n2460), .ZN(n2438) );
  NAND2_X1 U3140 ( .A1(n2438), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3141 ( .A1(n2439), .A2(n2461), .ZN(n2449) );
  OR2_X1 U3142 ( .A1(n2439), .A2(n2461), .ZN(n2440) );
  MUX2_X1 U3143 ( .A(DATAI_15_), .B(n4625), .S(n3587), .Z(n4199) );
  NAND2_X1 U3144 ( .A1(n4195), .A2(n4199), .ZN(n2441) );
  AOI21_X1 U3145 ( .B1(n4065), .B2(n2441), .A(n2251), .ZN(n4045) );
  NAND2_X1 U3146 ( .A1(n3588), .A2(REG1_REG_16__SCAN_IN), .ZN(n2448) );
  AND2_X1 U3147 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2442) );
  AOI21_X1 U31480 ( .B1(n2443), .B2(REG3_REG_15__SCAN_IN), .A(
        REG3_REG_16__SCAN_IN), .ZN(n2444) );
  OR2_X1 U31490 ( .A1(n2453), .A2(n2444), .ZN(n4053) );
  INV_X1 U3150 ( .A(n4053), .ZN(n3495) );
  NAND2_X1 U3151 ( .A1(n2318), .A2(n3495), .ZN(n2447) );
  NAND2_X1 U3152 ( .A1(n3589), .A2(REG0_REG_16__SCAN_IN), .ZN(n2446) );
  INV_X1 U3153 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4054) );
  OR2_X1 U3154 ( .A1(n3590), .A2(n4054), .ZN(n2445) );
  NAND2_X1 U3155 ( .A1(n2449), .A2(IR_REG_31__SCAN_IN), .ZN(n2450) );
  XNOR2_X1 U3156 ( .A(n2450), .B(IR_REG_16__SCAN_IN), .ZN(n3811) );
  MUX2_X1 U3157 ( .A(DATAI_16_), .B(n3811), .S(n3587), .Z(n4060) );
  NAND2_X1 U3158 ( .A1(n4031), .A2(n4060), .ZN(n3710) );
  NAND2_X1 U3159 ( .A1(n4201), .A2(n4190), .ZN(n3596) );
  NAND2_X1 U3160 ( .A1(n4045), .A2(n2451), .ZN(n4046) );
  NAND2_X1 U3161 ( .A1(n4201), .A2(n4060), .ZN(n2452) );
  NAND2_X1 U3162 ( .A1(n3588), .A2(REG1_REG_17__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3163 ( .A1(n3589), .A2(REG0_REG_17__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3164 ( .A1(n2453), .A2(REG3_REG_17__SCAN_IN), .ZN(n2454) );
  AND2_X1 U3165 ( .A1(n2454), .A2(n2480), .ZN(n4038) );
  NAND2_X1 U3166 ( .A1(n2295), .A2(n4038), .ZN(n2456) );
  INV_X1 U3167 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4040) );
  OR2_X1 U3168 ( .A1(n3590), .A2(n4040), .ZN(n2455) );
  INV_X1 U3169 ( .A(DATAI_17_), .ZN(n2465) );
  INV_X1 U3170 ( .A(IR_REG_16__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3171 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  XNOR2_X1 U3172 ( .A(n2464), .B(IR_REG_17__SCAN_IN), .ZN(n4621) );
  INV_X1 U3173 ( .A(n4621), .ZN(n4573) );
  MUX2_X1 U3174 ( .A(n2465), .B(n4573), .S(n3587), .Z(n4037) );
  NAND2_X1 U3175 ( .A1(n4191), .A2(n4037), .ZN(n2467) );
  INV_X1 U3176 ( .A(n4037), .ZN(n4028) );
  AND2_X1 U3177 ( .A1(n3748), .A2(n4028), .ZN(n2466) );
  NAND2_X1 U3178 ( .A1(n3588), .A2(REG1_REG_18__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3179 ( .A1(n3589), .A2(REG0_REG_18__SCAN_IN), .ZN(n2471) );
  XNOR2_X1 U3180 ( .A(n2480), .B(REG3_REG_18__SCAN_IN), .ZN(n4021) );
  NAND2_X1 U3181 ( .A1(n2295), .A2(n4021), .ZN(n2470) );
  INV_X1 U3182 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2468) );
  OR2_X1 U3183 ( .A1(n3590), .A2(n2468), .ZN(n2469) );
  NAND2_X1 U3184 ( .A1(n2486), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  XNOR2_X1 U3185 ( .A(n2474), .B(IR_REG_18__SCAN_IN), .ZN(n3804) );
  MUX2_X1 U3186 ( .A(DATAI_18_), .B(n3804), .S(n3587), .Z(n4017) );
  NAND2_X1 U3187 ( .A1(n4000), .A2(n4017), .ZN(n3990) );
  INV_X1 U3188 ( .A(n4017), .ZN(n3556) );
  NAND2_X1 U3189 ( .A1(n4029), .A2(n3556), .ZN(n3991) );
  NAND2_X1 U3190 ( .A1(n3990), .A2(n3991), .ZN(n4010) );
  NAND2_X1 U3191 ( .A1(n4008), .A2(n4010), .ZN(n4009) );
  NAND2_X1 U3192 ( .A1(n4000), .A2(n3556), .ZN(n2475) );
  NAND2_X1 U3193 ( .A1(n4009), .A2(n2475), .ZN(n3986) );
  INV_X1 U3194 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2476) );
  OR2_X1 U3195 ( .A1(n3590), .A2(n2476), .ZN(n2485) );
  NAND2_X1 U3196 ( .A1(n3588), .A2(REG1_REG_19__SCAN_IN), .ZN(n2484) );
  INV_X1 U3197 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2478) );
  INV_X1 U3198 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2477) );
  OAI21_X1 U3199 ( .B1(n2480), .B2(n2478), .A(n2477), .ZN(n2481) );
  NAND2_X1 U3200 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2479) );
  AND2_X1 U3201 ( .A1(n2481), .A2(n2494), .ZN(n4003) );
  NAND2_X1 U3202 ( .A1(n2295), .A2(n4003), .ZN(n2483) );
  NAND2_X1 U3203 ( .A1(n3589), .A2(REG0_REG_19__SCAN_IN), .ZN(n2482) );
  NAND4_X1 U3204 ( .A1(n2485), .A2(n2484), .A3(n2483), .A4(n2482), .ZN(n4172)
         );
  NAND2_X1 U3205 ( .A1(n2488), .A2(n2487), .ZN(n2556) );
  OR2_X1 U3206 ( .A1(n2488), .A2(n2487), .ZN(n2489) );
  INV_X1 U3207 ( .A(n3820), .ZN(n4472) );
  MUX2_X1 U3208 ( .A(DATAI_19_), .B(n4472), .S(n3587), .Z(n3361) );
  NAND2_X1 U3209 ( .A1(n3986), .A2(n2490), .ZN(n2492) );
  NAND2_X1 U32100 ( .A1(n3555), .A2(n4002), .ZN(n2491) );
  INV_X1 U32110 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2493) );
  OR2_X1 U32120 ( .A1(n3590), .A2(n2493), .ZN(n2499) );
  NAND2_X1 U32130 ( .A1(n3588), .A2(REG1_REG_20__SCAN_IN), .ZN(n2498) );
  AND2_X1 U32140 ( .A1(n2494), .A2(n4346), .ZN(n2495) );
  NOR2_X1 U32150 ( .A1(n2504), .A2(n2495), .ZN(n3978) );
  NAND2_X1 U32160 ( .A1(n2318), .A2(n3978), .ZN(n2497) );
  NAND2_X1 U32170 ( .A1(n2296), .A2(REG0_REG_20__SCAN_IN), .ZN(n2496) );
  INV_X1 U32180 ( .A(DATAI_20_), .ZN(n2500) );
  NOR2_X1 U32190 ( .A1(n3997), .A2(n4170), .ZN(n2502) );
  NAND2_X1 U32200 ( .A1(n3997), .A2(n4170), .ZN(n2501) );
  INV_X1 U32210 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2503) );
  OR2_X1 U32220 ( .A1(n3590), .A2(n2503), .ZN(n2509) );
  NAND2_X1 U32230 ( .A1(n3588), .A2(REG1_REG_21__SCAN_IN), .ZN(n2508) );
  NOR2_X1 U32240 ( .A1(n2504), .A2(REG3_REG_21__SCAN_IN), .ZN(n2505) );
  NOR2_X1 U32250 ( .A1(n2512), .A2(n2505), .ZN(n3959) );
  NAND2_X1 U32260 ( .A1(n2295), .A2(n3959), .ZN(n2507) );
  NAND2_X1 U32270 ( .A1(n2296), .A2(REG0_REG_21__SCAN_IN), .ZN(n2506) );
  INV_X1 U32280 ( .A(n3962), .ZN(n4161) );
  AND2_X1 U32290 ( .A1(n4171), .A2(n4161), .ZN(n2511) );
  NAND2_X1 U32300 ( .A1(n3547), .A2(n3962), .ZN(n2510) );
  OAI21_X2 U32310 ( .B1(n3955), .B2(n2511), .A(n2510), .ZN(n3942) );
  INV_X1 U32320 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3948) );
  OR2_X1 U32330 ( .A1(n3590), .A2(n3948), .ZN(n2517) );
  NAND2_X1 U32340 ( .A1(n3588), .A2(REG1_REG_22__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32350 ( .A1(n3589), .A2(REG0_REG_22__SCAN_IN), .ZN(n2515) );
  OR2_X1 U32360 ( .A1(n2512), .A2(REG3_REG_22__SCAN_IN), .ZN(n2513) );
  AND2_X1 U32370 ( .A1(n2513), .A2(n2519), .ZN(n3946) );
  NAND2_X1 U32380 ( .A1(n2318), .A2(n3946), .ZN(n2514) );
  NAND2_X1 U32390 ( .A1(n2525), .A2(DATAI_22_), .ZN(n3937) );
  NAND2_X1 U32400 ( .A1(n3477), .A2(n3943), .ZN(n3917) );
  NAND2_X1 U32410 ( .A1(n4162), .A2(n3937), .ZN(n2597) );
  OR2_X1 U32420 ( .A1(n3590), .A2(n4389), .ZN(n2524) );
  NAND2_X1 U32430 ( .A1(n2519), .A2(n4429), .ZN(n2520) );
  AND2_X1 U32440 ( .A1(n2526), .A2(n2520), .ZN(n3928) );
  NAND2_X1 U32450 ( .A1(n3928), .A2(n2295), .ZN(n2523) );
  NAND2_X1 U32460 ( .A1(n3588), .A2(REG1_REG_23__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32470 ( .A1(n2296), .A2(REG0_REG_23__SCAN_IN), .ZN(n2521) );
  AND2_X1 U32480 ( .A1(n2526), .A2(n4347), .ZN(n2527) );
  OR2_X1 U32490 ( .A1(n2527), .A2(n2538), .ZN(n3905) );
  INV_X1 U32500 ( .A(n3590), .ZN(n2568) );
  AOI22_X1 U32510 ( .A1(n2568), .A2(REG2_REG_24__SCAN_IN), .B1(n2296), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32520 ( .A1(n3588), .A2(REG1_REG_24__SCAN_IN), .ZN(n2528) );
  INV_X1 U32530 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4336) );
  XNOR2_X1 U32540 ( .A(n2538), .B(n4336), .ZN(n3890) );
  NAND2_X1 U32550 ( .A1(n3890), .A2(n2295), .ZN(n2536) );
  INV_X1 U32560 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32570 ( .A1(n3588), .A2(REG1_REG_25__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32580 ( .A1(n3589), .A2(REG0_REG_25__SCAN_IN), .ZN(n2531) );
  OAI211_X1 U32590 ( .C1(n2533), .C2(n3590), .A(n2532), .B(n2531), .ZN(n2534)
         );
  INV_X1 U32600 ( .A(n2534), .ZN(n2535) );
  AND2_X1 U32610 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2537) );
  AOI21_X1 U32620 ( .B1(n2538), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2539) );
  AOI22_X1 U32630 ( .A1(n3588), .A2(REG1_REG_26__SCAN_IN), .B1(n3589), .B2(
        REG0_REG_26__SCAN_IN), .ZN(n2541) );
  INV_X1 U32640 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3867) );
  OR2_X1 U32650 ( .A1(n3590), .A2(n3867), .ZN(n2540) );
  INV_X1 U32660 ( .A(n4122), .ZN(n3850) );
  INV_X1 U32670 ( .A(n3866), .ZN(n4130) );
  NAND2_X1 U32680 ( .A1(n2543), .A2(REG3_REG_27__SCAN_IN), .ZN(n2548) );
  OR2_X1 U32690 ( .A1(n2543), .A2(REG3_REG_27__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32700 ( .A1(n2548), .A2(n2544), .ZN(n3849) );
  AOI22_X1 U32710 ( .A1(n3588), .A2(REG1_REG_27__SCAN_IN), .B1(n2296), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2546) );
  INV_X1 U32720 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3848) );
  OR2_X1 U32730 ( .A1(n3590), .A2(n3848), .ZN(n2545) );
  INV_X1 U32740 ( .A(DATAI_27_), .ZN(n2547) );
  INV_X1 U32750 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U32760 ( .A1(n2548), .A2(n3464), .ZN(n2549) );
  NAND2_X1 U32770 ( .A1(n3469), .A2(n2295), .ZN(n2554) );
  INV_X1 U32780 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U32790 ( .A1(n3589), .A2(REG0_REG_28__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32800 ( .A1(n3588), .A2(REG1_REG_28__SCAN_IN), .ZN(n2550) );
  OAI211_X1 U32810 ( .C1(n3590), .C2(n3316), .A(n2551), .B(n2550), .ZN(n2552)
         );
  INV_X1 U32820 ( .A(n2552), .ZN(n2553) );
  INV_X1 U32830 ( .A(DATAI_28_), .ZN(n2555) );
  AND2_X1 U32840 ( .A1(n4124), .A2(n3295), .ZN(n3613) );
  NOR2_X1 U32850 ( .A1(n4124), .A2(n3295), .ZN(n3618) );
  NAND2_X1 U32860 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32870 ( .A1(n2035), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  XNOR2_X1 U32880 ( .A(n2845), .B(n3739), .ZN(n2561) );
  NAND2_X1 U32890 ( .A1(n2561), .A2(n3820), .ZN(n4093) );
  NOR2_X1 U32900 ( .A1(n3820), .A2(n3739), .ZN(n2563) );
  NOR2_X1 U32910 ( .A1(n2564), .A2(n2659), .ZN(n2565) );
  MUX2_X1 U32920 ( .A(n2659), .B(n2565), .S(IR_REG_28__SCAN_IN), .Z(n2566) );
  INV_X1 U32930 ( .A(n2566), .ZN(n2567) );
  NAND2_X1 U32940 ( .A1(n2567), .A2(n2264), .ZN(n2788) );
  INV_X1 U32950 ( .A(n2788), .ZN(n2750) );
  AOI22_X1 U32960 ( .A1(REG1_REG_29__SCAN_IN), .A2(n3588), .B1(n2568), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U32970 ( .A1(n3589), .A2(REG0_REG_29__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U32980 ( .C1(n3835), .C2(n2571), .A(n2570), .B(n2569), .ZN(n3744)
         );
  INV_X1 U32990 ( .A(n3744), .ZN(n3466) );
  INV_X1 U33000 ( .A(n2562), .ZN(n4471) );
  INV_X1 U33010 ( .A(n3739), .ZN(n2572) );
  INV_X1 U33020 ( .A(n3295), .ZN(n3465) );
  OAI22_X1 U33030 ( .A1(n3466), .A2(n4219), .B1(n4232), .B2(n3465), .ZN(n2573)
         );
  AOI21_X1 U33040 ( .B1(n4224), .B2(n4131), .A(n2573), .ZN(n2608) );
  INV_X1 U33050 ( .A(n2712), .ZN(n2575) );
  NAND2_X1 U33060 ( .A1(n2799), .A2(n3675), .ZN(n2853) );
  NAND2_X1 U33070 ( .A1(n2578), .A2(n2867), .ZN(n3680) );
  NAND2_X1 U33080 ( .A1(n3756), .A2(n2884), .ZN(n3677) );
  NAND2_X1 U33090 ( .A1(n2853), .A2(n3639), .ZN(n2579) );
  INV_X1 U33100 ( .A(n3681), .ZN(n2580) );
  AND2_X1 U33110 ( .A1(n3754), .A2(n2946), .ZN(n2940) );
  NAND2_X1 U33120 ( .A1(n2992), .A2(n3009), .ZN(n3688) );
  INV_X1 U33130 ( .A(n2990), .ZN(n2581) );
  NAND2_X1 U33140 ( .A1(n3753), .A2(n2581), .ZN(n3686) );
  NAND2_X1 U33150 ( .A1(n2976), .A2(n3686), .ZN(n2582) );
  INV_X1 U33160 ( .A(n3753), .ZN(n2933) );
  NAND2_X1 U33170 ( .A1(n2933), .A2(n2990), .ZN(n3690) );
  INV_X1 U33180 ( .A(n3691), .ZN(n2583) );
  NAND2_X1 U33190 ( .A1(n3152), .A2(n3117), .ZN(n3696) );
  NAND2_X1 U33200 ( .A1(n3751), .A2(n3138), .ZN(n3692) );
  NAND2_X1 U33210 ( .A1(n2584), .A2(n3692), .ZN(n3098) );
  AND2_X1 U33220 ( .A1(n3750), .A2(n3175), .ZN(n3097) );
  NAND2_X1 U33230 ( .A1(n2585), .A2(n3160), .ZN(n3697) );
  NAND2_X1 U33240 ( .A1(n4096), .A2(n3208), .ZN(n3701) );
  NAND2_X1 U33250 ( .A1(n3174), .A2(n3197), .ZN(n3704) );
  NAND2_X1 U33260 ( .A1(n4223), .A2(n4233), .ZN(n3233) );
  NAND2_X1 U33270 ( .A1(n4236), .A2(n4218), .ZN(n3214) );
  NAND2_X1 U33280 ( .A1(n3233), .A2(n3214), .ZN(n2587) );
  INV_X1 U33290 ( .A(n3220), .ZN(n2586) );
  NOR2_X1 U33300 ( .A1(n2587), .A2(n2586), .ZN(n3702) );
  NAND2_X1 U33310 ( .A1(n4086), .A2(n3702), .ZN(n2590) );
  NAND2_X1 U33320 ( .A1(n3261), .A2(n3276), .ZN(n3234) );
  NAND2_X1 U33330 ( .A1(n3218), .A2(n3234), .ZN(n2589) );
  INV_X1 U33340 ( .A(n2587), .ZN(n2588) );
  NOR2_X1 U33350 ( .A1(n4236), .A2(n4218), .ZN(n3215) );
  AOI21_X1 U33360 ( .B1(n2589), .B2(n2588), .A(n3215), .ZN(n3706) );
  NAND2_X1 U33370 ( .A1(n2590), .A2(n3706), .ZN(n3595) );
  INV_X1 U33380 ( .A(n3285), .ZN(n3662) );
  NAND2_X1 U33390 ( .A1(n3595), .A2(n3662), .ZN(n2591) );
  NAND2_X1 U33400 ( .A1(n2591), .A2(n3594), .ZN(n4069) );
  NAND2_X1 U33410 ( .A1(n4209), .A2(n4199), .ZN(n3598) );
  NAND2_X1 U33420 ( .A1(n4195), .A2(n4080), .ZN(n3601) );
  NAND2_X1 U33430 ( .A1(n3598), .A2(n3601), .ZN(n4068) );
  NAND2_X1 U33440 ( .A1(n4066), .A2(n3601), .ZN(n4050) );
  NAND2_X1 U33450 ( .A1(n4050), .A2(n4049), .ZN(n4048) );
  NAND2_X1 U33460 ( .A1(n4172), .A2(n4002), .ZN(n2592) );
  AND2_X1 U33470 ( .A1(n3991), .A2(n2592), .ZN(n2594) );
  NAND2_X1 U33480 ( .A1(n3748), .A2(n4037), .ZN(n3987) );
  NAND2_X1 U33490 ( .A1(n2594), .A2(n3987), .ZN(n3603) );
  NAND2_X1 U33500 ( .A1(n4191), .A2(n4028), .ZN(n3988) );
  NAND2_X1 U33510 ( .A1(n3990), .A2(n3988), .ZN(n2595) );
  NOR2_X1 U33520 ( .A1(n4172), .A2(n4002), .ZN(n2593) );
  AOI21_X1 U3353 ( .B1(n2595), .B2(n2594), .A(n2593), .ZN(n3970) );
  INV_X1 U33540 ( .A(n3997), .ZN(n4165) );
  NAND2_X1 U3355 ( .A1(n4165), .A2(n4170), .ZN(n2596) );
  NAND2_X1 U3356 ( .A1(n3997), .A2(n3981), .ZN(n3605) );
  NAND2_X1 U3357 ( .A1(n3547), .A2(n4161), .ZN(n3915) );
  AND2_X1 U3358 ( .A1(n3915), .A2(n3917), .ZN(n3717) );
  NAND2_X1 U3359 ( .A1(n3953), .A2(n3717), .ZN(n2600) );
  NAND2_X1 U3360 ( .A1(n4142), .A2(n3926), .ZN(n3631) );
  AND2_X1 U3361 ( .A1(n2597), .A2(n3631), .ZN(n3722) );
  AND2_X1 U3362 ( .A1(n4171), .A2(n3962), .ZN(n3914) );
  NAND2_X1 U3363 ( .A1(n3917), .A2(n3914), .ZN(n2598) );
  NAND2_X1 U3364 ( .A1(n3722), .A2(n2598), .ZN(n3611) );
  INV_X1 U3365 ( .A(n3611), .ZN(n2599) );
  NAND2_X1 U3366 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  NOR2_X1 U3367 ( .A1(n4142), .A2(n3926), .ZN(n3608) );
  INV_X1 U3368 ( .A(n3608), .ZN(n3632) );
  OR2_X1 U3369 ( .A1(n3747), .A2(n3902), .ZN(n3630) );
  INV_X1 U3370 ( .A(n3630), .ZN(n3609) );
  OR2_X1 U3371 ( .A1(n4122), .A2(n3866), .ZN(n2602) );
  OR2_X1 U3372 ( .A1(n3746), .A2(n3889), .ZN(n3859) );
  NAND2_X1 U3373 ( .A1(n2602), .A2(n3859), .ZN(n3720) );
  NAND2_X1 U3374 ( .A1(n3746), .A2(n3889), .ZN(n3644) );
  NAND2_X1 U3375 ( .A1(n3747), .A2(n3902), .ZN(n3879) );
  AND2_X1 U3376 ( .A1(n3644), .A2(n3879), .ZN(n3858) );
  NAND2_X1 U3377 ( .A1(n4122), .A2(n3866), .ZN(n3619) );
  OAI21_X1 U3378 ( .B1(n3720), .B2(n3858), .A(n3619), .ZN(n3724) );
  INV_X1 U3379 ( .A(n3724), .ZN(n2603) );
  XNOR2_X1 U3380 ( .A(n4131), .B(n4121), .ZN(n3666) );
  NOR2_X1 U3381 ( .A1(n4131), .A2(n3847), .ZN(n3612) );
  INV_X1 U3382 ( .A(n3612), .ZN(n2604) );
  NAND2_X1 U3383 ( .A1(n3845), .A2(n2604), .ZN(n3300) );
  INV_X1 U3384 ( .A(n3635), .ZN(n2605) );
  XNOR2_X1 U3385 ( .A(n3300), .B(n2605), .ZN(n2607) );
  NAND2_X1 U3386 ( .A1(n4471), .A2(n4470), .ZN(n3628) );
  NAND2_X1 U3387 ( .A1(n4472), .A2(n3739), .ZN(n2606) );
  NAND2_X1 U3388 ( .A1(n2607), .A2(n4047), .ZN(n3320) );
  OAI211_X1 U3389 ( .C1(n3314), .C2(n4227), .A(n2608), .B(n3320), .ZN(n2645)
         );
  OR2_X1 U3390 ( .A1(n2609), .A2(n2659), .ZN(n2622) );
  NAND2_X1 U3391 ( .A1(n2612), .A2(IR_REG_31__SCAN_IN), .ZN(n2613) );
  MUX2_X1 U3392 ( .A(IR_REG_31__SCAN_IN), .B(n2613), .S(IR_REG_25__SCAN_IN), 
        .Z(n2614) );
  NAND2_X1 U3393 ( .A1(n2614), .A2(n2031), .ZN(n2618) );
  NAND2_X1 U3394 ( .A1(n2653), .A2(n2618), .ZN(n2615) );
  MUX2_X1 U3395 ( .A(n2653), .B(n2615), .S(B_REG_SCAN_IN), .Z(n2617) );
  INV_X1 U3396 ( .A(D_REG_1__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3397 ( .A1(n2662), .A2(n2667), .ZN(n2839) );
  INV_X1 U3398 ( .A(n2664), .ZN(n2636) );
  NAND2_X1 U3399 ( .A1(n2636), .A2(n2618), .ZN(n2715) );
  NAND2_X1 U3400 ( .A1(n2839), .A2(n2715), .ZN(n2635) );
  INV_X1 U3401 ( .A(n2653), .ZN(n2619) );
  INV_X1 U3402 ( .A(n2618), .ZN(n4469) );
  NAND2_X1 U3403 ( .A1(n4648), .A2(n3657), .ZN(n2732) );
  NAND2_X1 U3404 ( .A1(n2562), .A2(n3820), .ZN(n2718) );
  NAND2_X1 U3405 ( .A1(n2718), .A2(n2719), .ZN(n2836) );
  NAND2_X1 U3406 ( .A1(n2732), .A2(n2836), .ZN(n2623) );
  NOR2_X1 U3407 ( .A1(n2838), .A2(n2623), .ZN(n2634) );
  NOR4_X1 U3408 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2627) );
  NOR4_X1 U3409 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2626) );
  NOR4_X1 U3410 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2625) );
  NOR4_X1 U3411 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2624) );
  NAND4_X1 U3412 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n2633)
         );
  NOR2_X1 U3413 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_9__SCAN_IN), .ZN(n2631) );
  NOR4_X1 U3414 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2630) );
  NOR4_X1 U3415 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2629) );
  NOR4_X1 U3416 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2628) );
  NAND4_X1 U3417 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n2632)
         );
  OAI21_X1 U3418 ( .B1(n2633), .B2(n2632), .A(n2662), .ZN(n2716) );
  NAND3_X1 U3419 ( .A1(n2635), .A2(n2634), .A3(n2716), .ZN(n2644) );
  NAND2_X1 U3420 ( .A1(n2662), .A2(n4373), .ZN(n2637) );
  NAND2_X1 U3421 ( .A1(n2636), .A2(n2653), .ZN(n2668) );
  INV_X1 U3422 ( .A(n2840), .ZN(n2717) );
  MUX2_X1 U3423 ( .A(REG0_REG_28__SCAN_IN), .B(n2645), .S(n4658), .Z(n2638) );
  INV_X1 U3424 ( .A(n2638), .ZN(n2643) );
  NAND2_X1 U3425 ( .A1(n2896), .A2(n2897), .ZN(n2895) );
  NOR2_X1 U3426 ( .A1(n2895), .A2(n2812), .ZN(n2859) );
  NAND2_X1 U3427 ( .A1(n3236), .A2(n4218), .ZN(n3286) );
  INV_X1 U3428 ( .A(n2640), .ZN(n4070) );
  INV_X1 U3429 ( .A(n3846), .ZN(n2641) );
  OAI21_X1 U3430 ( .B1(n2641), .B2(n3465), .A(n3309), .ZN(n3315) );
  NAND2_X1 U3431 ( .A1(n2643), .A2(n2642), .ZN(U3514) );
  MUX2_X1 U3432 ( .A(REG1_REG_28__SCAN_IN), .B(n2645), .S(n4665), .Z(n2646) );
  INV_X1 U3433 ( .A(n2646), .ZN(n2648) );
  NAND2_X1 U3434 ( .A1(n2648), .A2(n2647), .ZN(U3546) );
  INV_X1 U3435 ( .A(n4617), .ZN(n2665) );
  INV_X2 U3436 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3437 ( .A(n3767), .ZN(n3778) );
  INV_X1 U3438 ( .A(DATAI_2_), .ZN(n2649) );
  MUX2_X1 U3439 ( .A(n3778), .B(n2649), .S(U3149), .Z(n2650) );
  INV_X1 U3440 ( .A(n2650), .ZN(U3350) );
  MUX2_X1 U3441 ( .A(n2363), .B(n3055), .S(STATE_REG_SCAN_IN), .Z(n2651) );
  INV_X1 U3442 ( .A(n2651), .ZN(U3344) );
  INV_X1 U3443 ( .A(DATAI_22_), .ZN(n4368) );
  NAND2_X1 U3444 ( .A1(n3739), .A2(STATE_REG_SCAN_IN), .ZN(n2652) );
  OAI21_X1 U3445 ( .B1(STATE_REG_SCAN_IN), .B2(n4368), .A(n2652), .ZN(U3330)
         );
  INV_X1 U3446 ( .A(DATAI_24_), .ZN(n4426) );
  MUX2_X1 U3447 ( .A(n4426), .B(n2653), .S(STATE_REG_SCAN_IN), .Z(n2654) );
  INV_X1 U3448 ( .A(n2654), .ZN(U3328) );
  INV_X1 U3449 ( .A(DATAI_26_), .ZN(n4388) );
  NAND2_X1 U3450 ( .A1(n2664), .A2(STATE_REG_SCAN_IN), .ZN(n2655) );
  OAI21_X1 U3451 ( .B1(STATE_REG_SCAN_IN), .B2(n4388), .A(n2655), .ZN(U3326)
         );
  XNOR2_X1 U3452 ( .A(n2656), .B(IR_REG_27__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U3453 ( .A1(n4483), .A2(STATE_REG_SCAN_IN), .ZN(n2657) );
  OAI21_X1 U3454 ( .B1(STATE_REG_SCAN_IN), .B2(n2547), .A(n2657), .ZN(U3325)
         );
  NAND2_X1 U3455 ( .A1(n2750), .A2(STATE_REG_SCAN_IN), .ZN(n2658) );
  OAI21_X1 U3456 ( .B1(STATE_REG_SCAN_IN), .B2(n2555), .A(n2658), .ZN(U3324)
         );
  INV_X1 U3457 ( .A(DATAI_31_), .ZN(n3585) );
  OR4_X1 U34580 ( .A1(n2660), .A2(IR_REG_30__SCAN_IN), .A3(n2659), .A4(U3149), 
        .ZN(n2661) );
  OAI21_X1 U34590 ( .B1(STATE_REG_SCAN_IN), .B2(n3585), .A(n2661), .ZN(U3321)
         );
  INV_X1 U3460 ( .A(n2662), .ZN(n2663) );
  NOR3_X1 U3461 ( .A1(n2665), .A2(n2664), .A3(n4469), .ZN(n2666) );
  AOI21_X1 U3462 ( .B1(n4614), .B2(n2667), .A(n2666), .ZN(U3459) );
  INV_X1 U3463 ( .A(n2668), .ZN(n2669) );
  AOI22_X1 U3464 ( .A1(n4614), .A2(n4373), .B1(n2669), .B2(n4617), .ZN(U3458)
         );
  AND2_X1 U3465 ( .A1(n2877), .A2(n2719), .ZN(n2670) );
  OR2_X1 U3466 ( .A1(n2877), .A2(U3149), .ZN(n3741) );
  NAND2_X1 U34670 ( .A1(n2838), .A2(n3741), .ZN(n2679) );
  INV_X1 U3468 ( .A(n2679), .ZN(n2671) );
  NOR2_X2 U34690 ( .A1(n2680), .A2(n2671), .ZN(n4579) );
  NOR2_X1 U3470 ( .A1(n4579), .A2(U4043), .ZN(U3148) );
  INV_X1 U34710 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U3472 ( .A1(n4172), .A2(U4043), .ZN(n2672) );
  OAI21_X1 U34730 ( .B1(U4043), .B2(n4350), .A(n2672), .ZN(U3569) );
  INV_X1 U3474 ( .A(n2745), .ZN(n4476) );
  MUX2_X1 U34750 ( .A(REG2_REG_2__SCAN_IN), .B(n2673), .S(n3767), .Z(n2676) );
  AND2_X1 U3476 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3759)
         );
  NAND2_X1 U34770 ( .A1(n4479), .A2(REG2_REG_1__SCAN_IN), .ZN(n3769) );
  NAND2_X1 U3478 ( .A1(n3768), .A2(n3769), .ZN(n2675) );
  XNOR2_X1 U34790 ( .A(n2677), .B(n4477), .ZN(n2756) );
  INV_X1 U3480 ( .A(n2677), .ZN(n2678) );
  INV_X1 U34810 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3007) );
  MUX2_X1 U3482 ( .A(REG2_REG_5__SCAN_IN), .B(n3007), .S(n2745), .Z(n2738) );
  NOR2_X1 U34830 ( .A1(n2739), .A2(n2738), .ZN(n2737) );
  AOI21_X1 U3484 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4476), .A(n2737), .ZN(n2700)
         );
  XNOR2_X1 U34850 ( .A(n2700), .B(n4475), .ZN(n2702) );
  XNOR2_X1 U3486 ( .A(n2702), .B(REG2_REG_6__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U34870 ( .A1(n2680), .A2(n2679), .ZN(n4492) );
  INV_X1 U3488 ( .A(n4492), .ZN(n2681) );
  INV_X1 U34890 ( .A(n4483), .ZN(n2749) );
  NOR2_X1 U3490 ( .A1(n2788), .A2(n2749), .ZN(n3737) );
  INV_X1 U34910 ( .A(n4586), .ZN(n3783) );
  NAND2_X1 U3492 ( .A1(n4579), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U34930 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n2968) );
  NAND2_X1 U3494 ( .A1(n2682), .A2(n2968), .ZN(n2693) );
  INV_X1 U34950 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2683) );
  MUX2_X1 U3496 ( .A(REG1_REG_2__SCAN_IN), .B(n2683), .S(n3767), .Z(n3775) );
  INV_X1 U34970 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2684) );
  AND2_X1 U3498 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3761)
         );
  NAND2_X1 U34990 ( .A1(n4479), .A2(REG1_REG_1__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3500 ( .A1(n3760), .A2(n2685), .ZN(n3774) );
  NAND2_X1 U35010 ( .A1(n3775), .A2(n3774), .ZN(n3773) );
  NAND2_X1 U3502 ( .A1(n3767), .A2(REG1_REG_2__SCAN_IN), .ZN(n2686) );
  NAND2_X1 U35030 ( .A1(n3773), .A2(n2686), .ZN(n2688) );
  INV_X1 U3504 ( .A(n4478), .ZN(n2687) );
  XNOR2_X1 U35050 ( .A(n2688), .B(n2687), .ZN(n3785) );
  NAND2_X1 U35060 ( .A1(n3785), .A2(REG1_REG_3__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U35070 ( .A1(n2688), .A2(n4478), .ZN(n2689) );
  NAND2_X1 U35080 ( .A1(n3784), .A2(n2689), .ZN(n2690) );
  INV_X1 U35090 ( .A(n4477), .ZN(n2763) );
  MUX2_X1 U35100 ( .A(REG1_REG_5__SCAN_IN), .B(n4399), .S(n2745), .Z(n2742) );
  AOI21_X1 U35110 ( .B1(REG1_REG_5__SCAN_IN), .B2(n4476), .A(n2741), .ZN(n2696) );
  XOR2_X1 U35120 ( .A(n4475), .B(n2696), .Z(n2691) );
  INV_X1 U35130 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2997) );
  NOR2_X2 U35140 ( .A1(n4492), .A2(n4483), .ZN(n4581) );
  INV_X1 U35150 ( .A(n4581), .ZN(n2740) );
  NOR2_X1 U35160 ( .A1(n2691), .A2(n2997), .ZN(n2697) );
  AOI211_X1 U35170 ( .C1(n2691), .C2(n2997), .A(n2740), .B(n2697), .ZN(n2692)
         );
  AOI211_X1 U35180 ( .C1(n3783), .C2(n4475), .A(n2693), .B(n2692), .ZN(n2694)
         );
  OAI21_X1 U35190 ( .B1(n2695), .B2(n4575), .A(n2694), .ZN(U3246) );
  NOR2_X1 U35200 ( .A1(n4474), .A2(REG1_REG_7__SCAN_IN), .ZN(n2698) );
  INV_X1 U35210 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4663) );
  INV_X1 U35220 ( .A(n4474), .ZN(n2770) );
  XOR2_X1 U35230 ( .A(REG1_REG_8__SCAN_IN), .B(n3040), .Z(n2699) );
  NAND2_X1 U35240 ( .A1(n2699), .A2(n4581), .ZN(n2707) );
  INV_X1 U35250 ( .A(n2700), .ZN(n2701) );
  MUX2_X1 U35260 ( .A(n2343), .B(REG2_REG_7__SCAN_IN), .S(n4474), .Z(n2772) );
  XNOR2_X1 U35270 ( .A(REG2_REG_8__SCAN_IN), .B(n3057), .ZN(n2703) );
  NAND2_X1 U35280 ( .A1(n4526), .A2(n2703), .ZN(n2704) );
  NAND2_X1 U35290 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3118) );
  NAND2_X1 U35300 ( .A1(n2704), .A2(n3118), .ZN(n2705) );
  AOI21_X1 U35310 ( .B1(n4579), .B2(ADDR_REG_8__SCAN_IN), .A(n2705), .ZN(n2706) );
  OAI211_X1 U35320 ( .C1(n4586), .C2(n3055), .A(n2707), .B(n2706), .ZN(U3248)
         );
  INV_X1 U35330 ( .A(n3421), .ZN(n2957) );
  NOR2_X1 U35340 ( .A1(n2897), .A2(n3456), .ZN(n2709) );
  INV_X1 U35350 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2710) );
  OR2_X1 U35360 ( .A1(n2708), .A2(n2710), .ZN(n2711) );
  NAND2_X1 U35370 ( .A1(n2784), .A2(n2711), .ZN(n2786) );
  INV_X1 U35380 ( .A(n2708), .ZN(n2713) );
  AOI22_X1 U35390 ( .A1(n2797), .A2(n2957), .B1(IR_REG_0__SCAN_IN), .B2(n2713), 
        .ZN(n2714) );
  XNOR2_X1 U35400 ( .A(n2786), .B(n2785), .ZN(n2751) );
  AND2_X1 U35410 ( .A1(n2716), .A2(n2715), .ZN(n2842) );
  NAND2_X1 U35420 ( .A1(n2718), .A2(n2844), .ZN(n2721) );
  INV_X1 U35430 ( .A(n2719), .ZN(n2720) );
  NAND2_X1 U35440 ( .A1(n2721), .A2(n2720), .ZN(n2723) );
  NOR2_X1 U35450 ( .A1(n2838), .A2(n2723), .ZN(n2722) );
  INV_X1 U35460 ( .A(n2790), .ZN(n2728) );
  NAND2_X1 U35470 ( .A1(n2723), .A2(n4232), .ZN(n2724) );
  NAND2_X1 U35480 ( .A1(n2728), .A2(n2724), .ZN(n2725) );
  NAND2_X1 U35490 ( .A1(n2725), .A2(n2836), .ZN(n2879) );
  INV_X1 U35500 ( .A(n2879), .ZN(n2730) );
  NAND2_X1 U35510 ( .A1(n3820), .A2(n3739), .ZN(n2781) );
  INV_X1 U35520 ( .A(n2781), .ZN(n2726) );
  AND2_X1 U35530 ( .A1(n4617), .A2(n2726), .ZN(n2727) );
  NAND2_X1 U35540 ( .A1(n2728), .A2(n3736), .ZN(n2880) );
  NAND3_X1 U35550 ( .A1(n2730), .A2(n2729), .A3(n2880), .ZN(n2833) );
  NOR2_X1 U35560 ( .A1(n2838), .A2(n4232), .ZN(n2731) );
  NAND2_X1 U35570 ( .A1(n2790), .A2(n2731), .ZN(n2733) );
  AND2_X2 U35580 ( .A1(n2733), .A2(n4588), .ZN(n3577) );
  INV_X1 U35590 ( .A(n2281), .ZN(n2803) );
  AND2_X1 U35600 ( .A1(n2788), .A2(n3736), .ZN(n2734) );
  OAI22_X1 U35610 ( .A1(n3577), .A2(n2897), .B1(n2803), .B2(n3576), .ZN(n2735)
         );
  AOI21_X1 U35620 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2833), .A(n2735), .ZN(n2736) );
  OAI21_X1 U35630 ( .B1(n2751), .B2(n3583), .A(n2736), .ZN(U3229) );
  AOI211_X1 U35640 ( .C1(n2739), .C2(n2738), .A(n2737), .B(n4575), .ZN(n2748)
         );
  AOI211_X1 U35650 ( .C1(n2743), .C2(n2742), .A(n2741), .B(n2740), .ZN(n2747)
         );
  AND2_X1 U35660 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2935) );
  AOI21_X1 U35670 ( .B1(n4579), .B2(ADDR_REG_5__SCAN_IN), .A(n2935), .ZN(n2744) );
  OAI21_X1 U35680 ( .B1(n4586), .B2(n2745), .A(n2744), .ZN(n2746) );
  OR3_X1 U35690 ( .A1(n2748), .A2(n2747), .A3(n2746), .ZN(U3245) );
  NAND3_X1 U35700 ( .A1(n2751), .A2(n2750), .A3(n2749), .ZN(n2755) );
  AOI21_X1 U35710 ( .B1(n3737), .B2(n3759), .A(n3757), .ZN(n2754) );
  AND2_X1 U35720 ( .A1(n4483), .A2(n2752), .ZN(n2753) );
  OR2_X1 U35730 ( .A1(n2788), .A2(n2753), .ZN(n4484) );
  NAND2_X1 U35740 ( .A1(n4484), .A2(n2112), .ZN(n4487) );
  NAND3_X1 U35750 ( .A1(n2755), .A2(n2754), .A3(n4487), .ZN(n3782) );
  XOR2_X1 U35760 ( .A(REG2_REG_4__SCAN_IN), .B(n2756), .Z(n2765) );
  INV_X1 U35770 ( .A(n2757), .ZN(n2758) );
  INV_X1 U35780 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U35790 ( .A1(n2758), .A2(n4660), .ZN(n2759) );
  NAND3_X1 U35800 ( .A1(n4581), .A2(n2760), .A3(n2759), .ZN(n2762) );
  AND2_X1 U35810 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2924) );
  AOI21_X1 U3582 ( .B1(n4579), .B2(ADDR_REG_4__SCAN_IN), .A(n2924), .ZN(n2761)
         );
  OAI211_X1 U3583 ( .C1(n4586), .C2(n2763), .A(n2762), .B(n2761), .ZN(n2764)
         );
  AOI21_X1 U3584 ( .B1(n4526), .B2(n2765), .A(n2764), .ZN(n2766) );
  NAND2_X1 U3585 ( .A1(n3782), .A2(n2766), .ZN(U3244) );
  MUX2_X1 U3586 ( .A(REG1_REG_7__SCAN_IN), .B(n4663), .S(n4474), .Z(n2767) );
  XNOR2_X1 U3587 ( .A(n2768), .B(n2767), .ZN(n2776) );
  INV_X1 U3588 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4424) );
  NOR2_X1 U3589 ( .A1(STATE_REG_SCAN_IN), .A2(n4424), .ZN(n3093) );
  AOI21_X1 U3590 ( .B1(n4579), .B2(ADDR_REG_7__SCAN_IN), .A(n3093), .ZN(n2769)
         );
  OAI21_X1 U3591 ( .B1(n4586), .B2(n2770), .A(n2769), .ZN(n2775) );
  AOI211_X1 U3592 ( .C1(n2773), .C2(n2772), .A(n4575), .B(n2771), .ZN(n2774)
         );
  AOI211_X1 U3593 ( .C1(n4581), .C2(n2776), .A(n2775), .B(n2774), .ZN(n2777)
         );
  INV_X1 U3594 ( .A(n2777), .ZN(U3247) );
  XNOR2_X1 U3595 ( .A(n2782), .B(n3457), .ZN(n2815) );
  INV_X2 U3596 ( .A(n2871), .ZN(n3415) );
  OAI22_X1 U3597 ( .A1(n2783), .A2(n3459), .B1(n2896), .B2(n3415), .ZN(n2816)
         );
  XNOR2_X1 U3598 ( .A(n2815), .B(n2816), .ZN(n2819) );
  AOI22_X1 U3599 ( .A1(n2786), .A2(n2785), .B1(n3413), .B2(n2784), .ZN(n2818)
         );
  XNOR2_X1 U3600 ( .A(n2819), .B(n2818), .ZN(n2794) );
  INV_X1 U3601 ( .A(n3576), .ZN(n3275) );
  INV_X1 U3602 ( .A(n3736), .ZN(n2787) );
  NOR2_X1 U3603 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  AOI22_X1 U3604 ( .A1(n2291), .A2(n3275), .B1(n3579), .B2(n2712), .ZN(n2791)
         );
  OAI21_X1 U3605 ( .B1(n3577), .B2(n2896), .A(n2791), .ZN(n2792) );
  AOI21_X1 U3606 ( .B1(REG3_REG_1__SCAN_IN), .B2(n2833), .A(n2792), .ZN(n2793)
         );
  OAI21_X1 U3607 ( .B1(n2794), .B2(n3583), .A(n2793), .ZN(U3219) );
  NAND2_X1 U3608 ( .A1(n2712), .A2(n2897), .ZN(n3673) );
  NOR2_X1 U3609 ( .A1(n3633), .A2(n4641), .ZN(n2796) );
  INV_X1 U3610 ( .A(n4093), .ZN(n3968) );
  NOR2_X1 U3611 ( .A1(n3968), .A2(n4047), .ZN(n2795) );
  OAI22_X1 U3612 ( .A1(n3633), .A2(n2795), .B1(n2803), .B2(n4219), .ZN(n2849)
         );
  AOI211_X1 U3613 ( .C1(n2844), .C2(n2797), .A(n2796), .B(n2849), .ZN(n4638)
         );
  NAND2_X1 U3614 ( .A1(n4662), .A2(REG1_REG_0__SCAN_IN), .ZN(n2798) );
  OAI21_X1 U3615 ( .B1(n4638), .B2(n4662), .A(n2798), .ZN(U3518) );
  OAI21_X1 U3616 ( .B1(n3636), .B2(n2800), .A(n2799), .ZN(n2805) );
  NAND2_X1 U3617 ( .A1(n2812), .A2(n4200), .ZN(n2802) );
  NAND2_X1 U3618 ( .A1(n3756), .A2(n4235), .ZN(n2801) );
  OAI211_X1 U3619 ( .C1(n2803), .C2(n4238), .A(n2802), .B(n2801), .ZN(n2804)
         );
  AOI21_X1 U3620 ( .B1(n2805), .B2(n4047), .A(n2804), .ZN(n2810) );
  NAND2_X1 U3621 ( .A1(n2807), .A2(n3636), .ZN(n2808) );
  NAND2_X1 U3622 ( .A1(n2806), .A2(n2808), .ZN(n4603) );
  NAND2_X1 U3623 ( .A1(n4603), .A2(n3968), .ZN(n2809) );
  AND2_X1 U3624 ( .A1(n2810), .A2(n2809), .ZN(n4606) );
  NAND2_X1 U3625 ( .A1(n4603), .A2(n4648), .ZN(n2811) );
  NAND2_X1 U3626 ( .A1(n4606), .A2(n2811), .ZN(n2864) );
  INV_X1 U3627 ( .A(n2864), .ZN(n2814) );
  AOI21_X1 U3628 ( .B1(n2812), .B2(n2895), .A(n2859), .ZN(n4600) );
  AOI22_X1 U3629 ( .A1(n4600), .A2(n4460), .B1(REG0_REG_2__SCAN_IN), .B2(n4656), .ZN(n2813) );
  OAI21_X1 U3630 ( .B1(n2814), .B2(n4656), .A(n2813), .ZN(U3471) );
  NAND2_X1 U3631 ( .A1(n2815), .A2(n2816), .ZN(n2817) );
  XNOR2_X1 U3632 ( .A(n2821), .B(n3413), .ZN(n2824) );
  NOR2_X1 U3633 ( .A1(n2831), .A2(n3415), .ZN(n2822) );
  NAND2_X1 U3634 ( .A1(n2824), .A2(n2823), .ZN(n2873) );
  INV_X1 U3635 ( .A(n2826), .ZN(n2827) );
  INV_X1 U3636 ( .A(n2874), .ZN(n2828) );
  AOI21_X1 U3637 ( .B1(n2829), .B2(n2826), .A(n2828), .ZN(n2835) );
  AOI22_X1 U3638 ( .A1(n2281), .A2(n3579), .B1(n3275), .B2(n3756), .ZN(n2830)
         );
  OAI21_X1 U3639 ( .B1(n3577), .B2(n2831), .A(n2830), .ZN(n2832) );
  AOI21_X1 U3640 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2833), .A(n2832), .ZN(n2834)
         );
  OAI21_X1 U3641 ( .B1(n2835), .B2(n3583), .A(n2834), .ZN(U3234) );
  INV_X1 U3642 ( .A(n2836), .ZN(n2837) );
  NOR2_X1 U3643 ( .A1(n2838), .A2(n2837), .ZN(n2841) );
  NAND4_X1 U3644 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), .ZN(n2843)
         );
  AOI21_X1 U3645 ( .B1(n4020), .B2(n2844), .A(n4059), .ZN(n2851) );
  OR2_X1 U3646 ( .A1(n2845), .A2(n3820), .ZN(n2973) );
  INV_X1 U3647 ( .A(n2973), .ZN(n2846) );
  NAND2_X1 U3648 ( .A1(n3102), .A2(n2846), .ZN(n3985) );
  INV_X1 U3649 ( .A(n4588), .ZN(n4599) );
  AOI22_X1 U3650 ( .A1(n4607), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4599), .ZN(n2847) );
  OAI21_X1 U3651 ( .B1(n3633), .B2(n3985), .A(n2847), .ZN(n2848) );
  AOI21_X1 U3652 ( .B1(n2849), .B2(n3102), .A(n2848), .ZN(n2850) );
  OAI21_X1 U3653 ( .B1(n2851), .B2(n2897), .A(n2850), .ZN(U3290) );
  XNOR2_X1 U3654 ( .A(n2852), .B(n3639), .ZN(n2894) );
  INV_X1 U3655 ( .A(n2894), .ZN(n2858) );
  XNOR2_X1 U3656 ( .A(n2853), .B(n3639), .ZN(n2856) );
  AOI22_X1 U3657 ( .A1(n2291), .A2(n4224), .B1(n4200), .B2(n2867), .ZN(n2854)
         );
  OAI21_X1 U3658 ( .B1(n2916), .B2(n4219), .A(n2854), .ZN(n2855) );
  AOI21_X1 U3659 ( .B1(n2856), .B2(n4047), .A(n2855), .ZN(n2857) );
  OAI21_X1 U3660 ( .B1(n2894), .B2(n4093), .A(n2857), .ZN(n2889) );
  AOI21_X1 U3661 ( .B1(n4648), .B2(n2858), .A(n2889), .ZN(n2863) );
  OAI21_X1 U3662 ( .B1(n2859), .B2(n2884), .A(n3019), .ZN(n2860) );
  INV_X1 U3663 ( .A(n2860), .ZN(n2891) );
  AOI22_X1 U3664 ( .A1(n2891), .A2(n4460), .B1(REG0_REG_3__SCAN_IN), .B2(n4656), .ZN(n2861) );
  OAI21_X1 U3665 ( .B1(n2863), .B2(n4656), .A(n2861), .ZN(U3473) );
  AOI22_X1 U3666 ( .A1(n2891), .A2(n4246), .B1(REG1_REG_3__SCAN_IN), .B2(n4662), .ZN(n2862) );
  OAI21_X1 U3667 ( .B1(n2863), .B2(n4662), .A(n2862), .ZN(U3521) );
  MUX2_X1 U3668 ( .A(REG1_REG_2__SCAN_IN), .B(n2864), .S(n4665), .Z(n2865) );
  AOI21_X1 U3669 ( .B1(n4246), .B2(n4600), .A(n2865), .ZN(n2866) );
  INV_X1 U3670 ( .A(n2866), .ZN(U3520) );
  NAND2_X1 U3671 ( .A1(n3756), .A2(n2957), .ZN(n2869) );
  NAND2_X1 U3672 ( .A1(n2867), .A2(n3410), .ZN(n2868) );
  NAND2_X1 U3673 ( .A1(n2869), .A2(n2868), .ZN(n2870) );
  NOR2_X1 U3674 ( .A1(n2884), .A2(n3415), .ZN(n2872) );
  AOI21_X1 U3675 ( .B1(n3756), .B2(n3417), .A(n2872), .ZN(n2914) );
  XNOR2_X1 U3676 ( .A(n2913), .B(n2914), .ZN(n2876) );
  NAND2_X1 U3677 ( .A1(n2875), .A2(n2876), .ZN(n2920) );
  OAI21_X1 U3678 ( .B1(n2876), .B2(n2875), .A(n2920), .ZN(n2887) );
  NAND2_X1 U3679 ( .A1(n2708), .A2(n2877), .ZN(n2878) );
  OAI21_X1 U3680 ( .B1(n2879), .B2(n2878), .A(STATE_REG_SCAN_IN), .ZN(n2881)
         );
  MUX2_X1 U3681 ( .A(U3149), .B(n3580), .S(n2882), .Z(n2886) );
  AOI22_X1 U3682 ( .A1(n3579), .A2(n2291), .B1(n3755), .B2(n3275), .ZN(n2883)
         );
  OAI21_X1 U3683 ( .B1(n3577), .B2(n2884), .A(n2883), .ZN(n2885) );
  AOI211_X1 U3684 ( .C1(n2887), .C2(n3545), .A(n2886), .B(n2885), .ZN(n2888)
         );
  INV_X1 U3685 ( .A(n2888), .ZN(U3215) );
  NAND2_X1 U3686 ( .A1(n2889), .A2(n4591), .ZN(n2893) );
  OAI22_X1 U3687 ( .A1(n4591), .A2(n3786), .B1(REG3_REG_3__SCAN_IN), .B2(n4588), .ZN(n2890) );
  AOI21_X1 U3688 ( .B1(n2891), .B2(n4601), .A(n2890), .ZN(n2892) );
  OAI211_X1 U3689 ( .C1(n2894), .C2(n3985), .A(n2893), .B(n2892), .ZN(U3287)
         );
  OAI21_X1 U3690 ( .B1(n2897), .B2(n2896), .A(n2895), .ZN(n4639) );
  OR2_X1 U3691 ( .A1(n2574), .A2(n2899), .ZN(n2900) );
  NAND2_X1 U3692 ( .A1(n2898), .A2(n2900), .ZN(n4642) );
  NAND2_X1 U3693 ( .A1(n2901), .A2(n4200), .ZN(n2903) );
  NAND2_X1 U3694 ( .A1(n2712), .A2(n4224), .ZN(n2902) );
  OAI211_X1 U3695 ( .C1(n2820), .C2(n4219), .A(n2903), .B(n2902), .ZN(n2904)
         );
  INV_X1 U3696 ( .A(n2904), .ZN(n2907) );
  XNOR2_X1 U3697 ( .A(n2574), .B(n3671), .ZN(n2905) );
  NAND2_X1 U3698 ( .A1(n2905), .A2(n4047), .ZN(n2906) );
  OAI211_X1 U3699 ( .C1(n4642), .C2(n4093), .A(n2907), .B(n2906), .ZN(n4644)
         );
  MUX2_X1 U3700 ( .A(n4644), .B(REG2_REG_1__SCAN_IN), .S(n4607), .Z(n2908) );
  INV_X1 U3701 ( .A(n2908), .ZN(n2911) );
  INV_X1 U3702 ( .A(n4642), .ZN(n2909) );
  INV_X1 U3703 ( .A(n3985), .ZN(n4602) );
  AOI22_X1 U3704 ( .A1(n2909), .A2(n4602), .B1(REG3_REG_1__SCAN_IN), .B2(n4599), .ZN(n2910) );
  OAI211_X1 U3705 ( .C1(n4106), .C2(n4639), .A(n2911), .B(n2910), .ZN(U3289)
         );
  INV_X1 U3706 ( .A(n3580), .ZN(n3213) );
  INV_X1 U3707 ( .A(n2912), .ZN(n3021) );
  INV_X1 U3708 ( .A(n2913), .ZN(n2915) );
  NAND2_X1 U3709 ( .A1(n2915), .A2(n2914), .ZN(n2918) );
  AND2_X1 U3710 ( .A1(n2920), .A2(n2918), .ZN(n2922) );
  OAI22_X1 U3711 ( .A1(n2916), .A2(n3415), .B1(n3456), .B2(n3025), .ZN(n2917)
         );
  XNOR2_X1 U3712 ( .A(n2917), .B(n3413), .ZN(n2927) );
  OAI22_X1 U3713 ( .A1(n2916), .A2(n3459), .B1(n3415), .B2(n3025), .ZN(n2928)
         );
  XNOR2_X1 U3714 ( .A(n2927), .B(n2928), .ZN(n2921) );
  AND2_X1 U3715 ( .A1(n2921), .A2(n2918), .ZN(n2919) );
  NAND2_X1 U3716 ( .A1(n2920), .A2(n2919), .ZN(n2931) );
  OAI211_X1 U3717 ( .C1(n2922), .C2(n2921), .A(n3545), .B(n2931), .ZN(n2926)
         );
  OAI22_X1 U3718 ( .A1(n3577), .A2(n3025), .B1(n2992), .B2(n3576), .ZN(n2923)
         );
  AOI211_X1 U3719 ( .C1(n3579), .C2(n3756), .A(n2924), .B(n2923), .ZN(n2925)
         );
  OAI211_X1 U3720 ( .C1(n3213), .C2(n3021), .A(n2926), .B(n2925), .ZN(U3227)
         );
  INV_X1 U3721 ( .A(n2927), .ZN(n2929) );
  NAND2_X1 U3722 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  OAI22_X1 U3723 ( .A1(n2992), .A2(n3415), .B1(n2946), .B2(n3456), .ZN(n2932)
         );
  XNOR2_X1 U3724 ( .A(n2932), .B(n3413), .ZN(n2953) );
  OAI22_X1 U3725 ( .A1(n2992), .A2(n3459), .B1(n2946), .B2(n3421), .ZN(n2954)
         );
  XNOR2_X1 U3726 ( .A(n2953), .B(n2954), .ZN(n2951) );
  XNOR2_X1 U3727 ( .A(n2952), .B(n2951), .ZN(n2938) );
  OAI22_X1 U3728 ( .A1(n3577), .A2(n2946), .B1(n2933), .B2(n3576), .ZN(n2934)
         );
  AOI211_X1 U3729 ( .C1(n3579), .C2(n3755), .A(n2935), .B(n2934), .ZN(n2937)
         );
  NAND2_X1 U3730 ( .A1(n3580), .A2(n3005), .ZN(n2936) );
  OAI211_X1 U3731 ( .C1(n2938), .C2(n3583), .A(n2937), .B(n2936), .ZN(U3224)
         );
  INV_X1 U3732 ( .A(n2940), .ZN(n3683) );
  NAND2_X1 U3733 ( .A1(n3683), .A2(n3688), .ZN(n3647) );
  XOR2_X1 U3734 ( .A(n2939), .B(n3647), .Z(n3016) );
  XNOR2_X1 U3735 ( .A(n2941), .B(n3647), .ZN(n2942) );
  NAND2_X1 U3736 ( .A1(n2942), .A2(n4047), .ZN(n3013) );
  NOR2_X1 U3737 ( .A1(n2946), .A2(n4232), .ZN(n2943) );
  AOI21_X1 U3738 ( .B1(n3753), .B2(n4235), .A(n2943), .ZN(n2944) );
  OAI211_X1 U3739 ( .C1(n2916), .C2(n4238), .A(n3013), .B(n2944), .ZN(n2945)
         );
  AOI21_X1 U3740 ( .B1(n3016), .B2(n4651), .A(n2945), .ZN(n2988) );
  NAND2_X1 U3741 ( .A1(n4656), .A2(REG0_REG_5__SCAN_IN), .ZN(n2950) );
  OR2_X1 U3742 ( .A1(n3018), .A2(n2946), .ZN(n2947) );
  NAND2_X1 U3743 ( .A1(n2059), .A2(n2947), .ZN(n3012) );
  INV_X1 U3744 ( .A(n3012), .ZN(n2948) );
  NAND2_X1 U3745 ( .A1(n2948), .A2(n4460), .ZN(n2949) );
  OAI211_X1 U3746 ( .C1(n2988), .C2(n4656), .A(n2950), .B(n2949), .ZN(U3477)
         );
  INV_X1 U3747 ( .A(n2953), .ZN(n2955) );
  NAND2_X1 U3748 ( .A1(n2955), .A2(n2954), .ZN(n2956) );
  NAND2_X1 U3749 ( .A1(n3753), .A2(n2957), .ZN(n2959) );
  NAND2_X1 U3750 ( .A1(n2990), .A2(n3410), .ZN(n2958) );
  NAND2_X1 U3751 ( .A1(n2959), .A2(n2958), .ZN(n2960) );
  XNOR2_X1 U3752 ( .A(n2960), .B(n3457), .ZN(n2966) );
  INV_X1 U3753 ( .A(n2966), .ZN(n2964) );
  NAND2_X1 U3754 ( .A1(n3753), .A2(n3417), .ZN(n2962) );
  NAND2_X1 U3755 ( .A1(n2990), .A2(n2957), .ZN(n2961) );
  NAND2_X1 U3756 ( .A1(n2962), .A2(n2961), .ZN(n2965) );
  INV_X1 U3757 ( .A(n2965), .ZN(n2963) );
  AND2_X1 U3758 ( .A1(n2966), .A2(n2965), .ZN(n3086) );
  NOR2_X1 U3759 ( .A1(n2247), .A2(n3086), .ZN(n2967) );
  XNOR2_X1 U3760 ( .A(n3085), .B(n2967), .ZN(n2972) );
  INV_X1 U3761 ( .A(n3577), .ZN(n3277) );
  AOI22_X1 U3762 ( .A1(n3277), .A2(n2990), .B1(n3752), .B2(n3275), .ZN(n2969)
         );
  OAI211_X1 U3763 ( .C1(n2992), .C2(n3567), .A(n2969), .B(n2968), .ZN(n2970)
         );
  AOI21_X1 U3764 ( .B1(n2978), .B2(n3580), .A(n2970), .ZN(n2971) );
  OAI21_X1 U3765 ( .B1(n2972), .B2(n3583), .A(n2971), .ZN(U3236) );
  NAND2_X1 U3766 ( .A1(n4093), .A2(n2973), .ZN(n2974) );
  NAND2_X1 U3767 ( .A1(n3690), .A2(n3686), .ZN(n3648) );
  XNOR2_X1 U3768 ( .A(n2975), .B(n3648), .ZN(n2996) );
  XOR2_X1 U3769 ( .A(n3648), .B(n2976), .Z(n2994) );
  NAND2_X1 U3770 ( .A1(n3102), .A2(n4047), .ZN(n3294) );
  INV_X1 U3771 ( .A(n3294), .ZN(n2986) );
  NAND2_X1 U3772 ( .A1(n2059), .A2(n2990), .ZN(n2977) );
  NAND2_X1 U3773 ( .A1(n3075), .A2(n2977), .ZN(n3001) );
  INV_X1 U3774 ( .A(n2978), .ZN(n2979) );
  OAI22_X1 U3775 ( .A1(n4591), .A2(n2980), .B1(n2979), .B2(n4588), .ZN(n2981)
         );
  AOI21_X1 U3776 ( .B1(n2990), .B2(n4059), .A(n2981), .ZN(n2984) );
  AND2_X1 U3777 ( .A1(n4591), .A2(n4235), .ZN(n4073) );
  INV_X1 U3778 ( .A(n4073), .ZN(n4056) );
  NAND2_X1 U3779 ( .A1(n3102), .A2(n4224), .ZN(n4055) );
  OAI22_X1 U3780 ( .A1(n4056), .A2(n3139), .B1(n2992), .B2(n4055), .ZN(n2982)
         );
  INV_X1 U3781 ( .A(n2982), .ZN(n2983) );
  OAI211_X1 U3782 ( .C1(n3001), .C2(n4106), .A(n2984), .B(n2983), .ZN(n2985)
         );
  AOI21_X1 U3783 ( .B1(n2994), .B2(n2986), .A(n2985), .ZN(n2987) );
  OAI21_X1 U3784 ( .B1(n4084), .B2(n2996), .A(n2987), .ZN(U3284) );
  MUX2_X1 U3785 ( .A(n2988), .B(n4399), .S(n4662), .Z(n2989) );
  OAI21_X1 U3786 ( .B1(n4251), .B2(n3012), .A(n2989), .ZN(U3523) );
  AOI22_X1 U3787 ( .A1(n3752), .A2(n4235), .B1(n4200), .B2(n2990), .ZN(n2991)
         );
  OAI21_X1 U3788 ( .B1(n2992), .B2(n4238), .A(n2991), .ZN(n2993) );
  AOI21_X1 U3789 ( .B1(n2994), .B2(n4047), .A(n2993), .ZN(n2995) );
  OAI21_X1 U3790 ( .B1(n4227), .B2(n2996), .A(n2995), .ZN(n3003) );
  OAI22_X1 U3791 ( .A1(n3001), .A2(n4251), .B1(n4665), .B2(n2997), .ZN(n2998)
         );
  AOI21_X1 U3792 ( .B1(n3003), .B2(n4665), .A(n2998), .ZN(n2999) );
  INV_X1 U3793 ( .A(n2999), .ZN(U3524) );
  INV_X1 U3794 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3000) );
  OAI22_X1 U3795 ( .A1(n3001), .A2(n4466), .B1(n4658), .B2(n3000), .ZN(n3002)
         );
  AOI21_X1 U3796 ( .B1(n3003), .B2(n4658), .A(n3002), .ZN(n3004) );
  INV_X1 U3797 ( .A(n3004), .ZN(U3479) );
  INV_X1 U3798 ( .A(n3005), .ZN(n3006) );
  OAI22_X1 U3799 ( .A1(n4591), .A2(n3007), .B1(n3006), .B2(n4588), .ZN(n3008)
         );
  AOI21_X1 U3800 ( .B1(n3009), .B2(n4059), .A(n3008), .ZN(n3011) );
  INV_X1 U3801 ( .A(n4055), .ZN(n4075) );
  AOI22_X1 U3802 ( .A1(n3755), .A2(n4075), .B1(n4073), .B2(n3753), .ZN(n3010)
         );
  OAI211_X1 U3803 ( .C1(n3012), .C2(n4106), .A(n3011), .B(n3010), .ZN(n3015)
         );
  NOR2_X1 U3804 ( .A1(n3013), .A2(n4607), .ZN(n3014) );
  AOI211_X1 U3805 ( .C1(n3016), .C2(n4036), .A(n3015), .B(n3014), .ZN(n3017)
         );
  INV_X1 U3806 ( .A(n3017), .ZN(U3285) );
  AOI211_X1 U3807 ( .C1(n3020), .C2(n3019), .A(n4640), .B(n3018), .ZN(n4647)
         );
  NOR2_X1 U3808 ( .A1(n4588), .A2(n3021), .ZN(n3033) );
  XOR2_X1 U3809 ( .A(n3638), .B(n3023), .Z(n3032) );
  NAND2_X1 U3810 ( .A1(n3756), .A2(n4224), .ZN(n3024) );
  OAI21_X1 U3811 ( .B1(n4232), .B2(n3025), .A(n3024), .ZN(n3030) );
  NAND2_X1 U3812 ( .A1(n3027), .A2(n3638), .ZN(n3028) );
  NAND2_X1 U3813 ( .A1(n3026), .A2(n3028), .ZN(n3034) );
  NOR2_X1 U3814 ( .A1(n3034), .A2(n4093), .ZN(n3029) );
  AOI211_X1 U3815 ( .C1(n4235), .C2(n3754), .A(n3030), .B(n3029), .ZN(n3031)
         );
  OAI21_X1 U3816 ( .B1(n4212), .B2(n3032), .A(n3031), .ZN(n4646) );
  AOI211_X1 U3817 ( .C1(n4647), .C2(n3820), .A(n3033), .B(n4646), .ZN(n3036)
         );
  INV_X1 U3818 ( .A(n3034), .ZN(n4649) );
  AOI22_X1 U3819 ( .A1(n4649), .A2(n4602), .B1(REG2_REG_4__SCAN_IN), .B2(n4607), .ZN(n3035) );
  OAI21_X1 U3820 ( .B1(n3036), .B2(n4607), .A(n3035), .ZN(U3286) );
  NAND2_X1 U3821 ( .A1(n3054), .A2(REG1_REG_11__SCAN_IN), .ZN(n3044) );
  INV_X1 U3822 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3037) );
  AOI22_X1 U3823 ( .A1(n3054), .A2(REG1_REG_11__SCAN_IN), .B1(n3037), .B2(
        n4631), .ZN(n4516) );
  NAND2_X1 U3824 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4634), .ZN(n3041) );
  INV_X1 U3825 ( .A(n4634), .ZN(n4501) );
  INV_X1 U3826 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3038) );
  AOI22_X1 U3827 ( .A1(REG1_REG_9__SCAN_IN), .A2(n4634), .B1(n4501), .B2(n3038), .ZN(n4495) );
  INV_X1 U3828 ( .A(n3055), .ZN(n3039) );
  NAND2_X1 U3829 ( .A1(n3041), .A2(n4493), .ZN(n3042) );
  NAND2_X1 U3830 ( .A1(n3059), .A2(n3042), .ZN(n3043) );
  INV_X1 U3831 ( .A(n3059), .ZN(n4633) );
  XNOR2_X1 U3832 ( .A(n3042), .B(n4633), .ZN(n4506) );
  NAND2_X1 U3833 ( .A1(n3063), .A2(n3045), .ZN(n3046) );
  INV_X1 U3834 ( .A(n3063), .ZN(n4629) );
  XNOR2_X1 U3835 ( .A(n3045), .B(n4629), .ZN(n4532) );
  NAND2_X1 U3836 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4532), .ZN(n4531) );
  NAND2_X1 U3837 ( .A1(n3806), .A2(REG1_REG_13__SCAN_IN), .ZN(n3047) );
  OAI21_X1 U3838 ( .B1(n3806), .B2(REG1_REG_13__SCAN_IN), .A(n3047), .ZN(n3049) );
  INV_X1 U3839 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4229) );
  NAND2_X1 U3840 ( .A1(n3806), .A2(n4229), .ZN(n3048) );
  OAI211_X1 U3841 ( .C1(n3050), .C2(n3049), .A(n3805), .B(n4581), .ZN(n3052)
         );
  AND2_X1 U3842 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3537) );
  AOI21_X1 U3843 ( .B1(n4579), .B2(ADDR_REG_13__SCAN_IN), .A(n3537), .ZN(n3051) );
  OAI211_X1 U3844 ( .C1(n4586), .C2(n3806), .A(n3052), .B(n3051), .ZN(n3069)
         );
  NOR2_X1 U3845 ( .A1(n3806), .A2(n4398), .ZN(n3795) );
  NAND2_X1 U3846 ( .A1(n3806), .A2(n4398), .ZN(n3794) );
  INV_X1 U3847 ( .A(n3794), .ZN(n3053) );
  NOR2_X1 U3848 ( .A1(n3795), .A2(n3053), .ZN(n3067) );
  NAND2_X1 U3849 ( .A1(n3054), .A2(REG2_REG_11__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U3850 ( .A1(n3054), .A2(REG2_REG_11__SCAN_IN), .B1(n2390), .B2(
        n4631), .ZN(n4519) );
  NAND2_X1 U3851 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4634), .ZN(n3058) );
  AOI22_X1 U3852 ( .A1(REG2_REG_9__SCAN_IN), .A2(n4634), .B1(n4501), .B2(n2365), .ZN(n4498) );
  OAI22_X1 U3853 ( .A1(n3057), .A2(n4590), .B1(n3056), .B2(n3055), .ZN(n4497)
         );
  NAND2_X1 U3854 ( .A1(n4498), .A2(n4497), .ZN(n4496) );
  NAND2_X1 U3855 ( .A1(n3058), .A2(n4496), .ZN(n3060) );
  NAND2_X1 U3856 ( .A1(n3059), .A2(n3060), .ZN(n3061) );
  XNOR2_X1 U3857 ( .A(n3060), .B(n4633), .ZN(n4508) );
  NAND2_X1 U3858 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U3859 ( .A1(n3061), .A2(n4507), .ZN(n4518) );
  NAND2_X1 U3860 ( .A1(n4519), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U3861 ( .A1(n3062), .A2(n4517), .ZN(n3064) );
  NAND2_X1 U3862 ( .A1(n3063), .A2(n3064), .ZN(n3065) );
  XNOR2_X1 U3863 ( .A(n3064), .B(n4629), .ZN(n4527) );
  NAND2_X1 U3864 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4527), .ZN(n4525) );
  OAI21_X1 U3865 ( .B1(n3067), .B2(n3796), .A(n4526), .ZN(n3066) );
  AOI21_X1 U3866 ( .B1(n3067), .B2(n3796), .A(n3066), .ZN(n3068) );
  OR2_X1 U3867 ( .A1(n3069), .A2(n3068), .ZN(U3253) );
  OAI22_X1 U3868 ( .A1(n3152), .A2(n4219), .B1(n3091), .B2(n4232), .ZN(n3073)
         );
  XOR2_X1 U3869 ( .A(n3637), .B(n3070), .Z(n3071) );
  NOR2_X1 U3870 ( .A1(n3071), .A2(n4212), .ZN(n3072) );
  AOI211_X1 U3871 ( .C1(n4224), .C2(n3753), .A(n3073), .B(n3072), .ZN(n4655)
         );
  NAND2_X1 U3872 ( .A1(n3075), .A2(n3074), .ZN(n3077) );
  NAND2_X1 U3873 ( .A1(n3077), .A2(n3076), .ZN(n3078) );
  OR2_X1 U3874 ( .A1(n3135), .A2(n3078), .ZN(n4654) );
  INV_X1 U3875 ( .A(n4654), .ZN(n3080) );
  OAI22_X1 U3876 ( .A1(n4591), .A2(n2343), .B1(n3096), .B2(n4588), .ZN(n3079)
         );
  AOI21_X1 U3877 ( .B1(n3080), .B2(n4020), .A(n3079), .ZN(n3084) );
  NAND2_X1 U3878 ( .A1(n3082), .A2(n3637), .ZN(n4652) );
  NAND3_X1 U3879 ( .A1(n3081), .A2(n4652), .A3(n4036), .ZN(n3083) );
  OAI211_X1 U3880 ( .C1(n4655), .C2(n4607), .A(n3084), .B(n3083), .ZN(U3283)
         );
  OAI22_X1 U3881 ( .A1(n3139), .A2(n3415), .B1(n3456), .B2(n3091), .ZN(n3088)
         );
  XNOR2_X1 U3882 ( .A(n3088), .B(n3413), .ZN(n3110) );
  OAI22_X1 U3883 ( .A1(n3139), .A2(n3459), .B1(n3415), .B2(n3091), .ZN(n3111)
         );
  XNOR2_X1 U3884 ( .A(n3110), .B(n3111), .ZN(n3089) );
  OAI211_X1 U3885 ( .C1(n3090), .C2(n3089), .A(n3114), .B(n3545), .ZN(n3095)
         );
  OAI22_X1 U3886 ( .A1(n3577), .A2(n3091), .B1(n3152), .B2(n3576), .ZN(n3092)
         );
  AOI211_X1 U3887 ( .C1(n3579), .C2(n3753), .A(n3093), .B(n3092), .ZN(n3094)
         );
  OAI211_X1 U3888 ( .C1(n3213), .C2(n3096), .A(n3095), .B(n3094), .ZN(U3210)
         );
  INV_X1 U3889 ( .A(n3097), .ZN(n3699) );
  NAND2_X1 U3890 ( .A1(n3699), .A2(n3697), .ZN(n3646) );
  XNOR2_X1 U3891 ( .A(n3098), .B(n3646), .ZN(n3099) );
  NAND2_X1 U3892 ( .A1(n3099), .A2(n4047), .ZN(n3151) );
  XOR2_X1 U3893 ( .A(n3100), .B(n3646), .Z(n3154) );
  NAND2_X1 U3894 ( .A1(n3154), .A2(n4036), .ZN(n3109) );
  OAI21_X1 U3895 ( .B1(n3133), .B2(n3175), .A(n3101), .ZN(n3159) );
  INV_X1 U3896 ( .A(n3159), .ZN(n3107) );
  INV_X1 U3897 ( .A(n4607), .ZN(n3102) );
  OAI22_X1 U3898 ( .A1(n3103), .A2(n4588), .B1(n2365), .B2(n3102), .ZN(n3106)
         );
  AOI22_X1 U3899 ( .A1(n4059), .A2(n3160), .B1(n4073), .B2(n4096), .ZN(n3104)
         );
  OAI21_X1 U3900 ( .B1(n3152), .B2(n4055), .A(n3104), .ZN(n3105) );
  AOI211_X1 U3901 ( .C1(n3107), .C2(n4601), .A(n3106), .B(n3105), .ZN(n3108)
         );
  OAI211_X1 U3902 ( .C1(n4607), .C2(n3151), .A(n3109), .B(n3108), .ZN(U3281)
         );
  INV_X1 U3903 ( .A(n3110), .ZN(n3112) );
  NAND2_X1 U3904 ( .A1(n3112), .A2(n3111), .ZN(n3113) );
  NAND2_X1 U3905 ( .A1(n3114), .A2(n3113), .ZN(n3167) );
  OAI22_X1 U3906 ( .A1(n3152), .A2(n3459), .B1(n3138), .B2(n3415), .ZN(n3166)
         );
  OAI22_X1 U3907 ( .A1(n3152), .A2(n3421), .B1(n3138), .B2(n3456), .ZN(n3115)
         );
  XNOR2_X1 U3908 ( .A(n3115), .B(n3457), .ZN(n3165) );
  XOR2_X1 U3909 ( .A(n3166), .B(n3165), .Z(n3116) );
  XNOR2_X1 U3910 ( .A(n3167), .B(n3116), .ZN(n3122) );
  AOI22_X1 U3911 ( .A1(n3277), .A2(n3117), .B1(n3275), .B2(n3750), .ZN(n3119)
         );
  OAI211_X1 U3912 ( .C1(n3139), .C2(n3567), .A(n3119), .B(n3118), .ZN(n3120)
         );
  AOI21_X1 U3913 ( .B1(n4587), .B2(n3580), .A(n3120), .ZN(n3121) );
  OAI21_X1 U3914 ( .B1(n3122), .B2(n3583), .A(n3121), .ZN(U3218) );
  AND2_X1 U3915 ( .A1(n3704), .A2(n3701), .ZN(n3654) );
  XNOR2_X1 U3916 ( .A(n3123), .B(n3654), .ZN(n3184) );
  INV_X1 U3917 ( .A(n3184), .ZN(n3132) );
  INV_X1 U3918 ( .A(n4101), .ZN(n3124) );
  AOI21_X1 U3919 ( .B1(n3197), .B2(n3101), .A(n3124), .ZN(n3192) );
  INV_X1 U3920 ( .A(n4059), .ZN(n4079) );
  AOI22_X1 U3921 ( .A1(n3749), .A2(n4073), .B1(n4075), .B2(n3750), .ZN(n3126)
         );
  AOI22_X1 U3922 ( .A1(n4607), .A2(REG2_REG_10__SCAN_IN), .B1(n3194), .B2(
        n4599), .ZN(n3125) );
  OAI211_X1 U3923 ( .C1(n3208), .C2(n4079), .A(n3126), .B(n3125), .ZN(n3127)
         );
  AOI21_X1 U3924 ( .B1(n3192), .B2(n4601), .A(n3127), .ZN(n3131) );
  INV_X1 U3925 ( .A(n3654), .ZN(n3128) );
  XNOR2_X1 U3926 ( .A(n3129), .B(n3128), .ZN(n3185) );
  NAND2_X1 U3927 ( .A1(n3185), .A2(n4036), .ZN(n3130) );
  OAI211_X1 U3928 ( .C1(n3132), .C2(n3294), .A(n3131), .B(n3130), .ZN(U3280)
         );
  INV_X1 U3929 ( .A(n3133), .ZN(n3134) );
  OAI21_X1 U3930 ( .B1(n3135), .B2(n3138), .A(n3134), .ZN(n4593) );
  INV_X1 U3931 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4386) );
  XNOR2_X1 U3932 ( .A(n3152), .B(n3138), .ZN(n3650) );
  XNOR2_X1 U3933 ( .A(n3136), .B(n3650), .ZN(n4595) );
  XNOR2_X1 U3934 ( .A(n3137), .B(n3650), .ZN(n3142) );
  OAI22_X1 U3935 ( .A1(n3139), .A2(n4238), .B1(n4232), .B2(n3138), .ZN(n3140)
         );
  AOI21_X1 U3936 ( .B1(n4235), .B2(n3750), .A(n3140), .ZN(n3141) );
  OAI21_X1 U3937 ( .B1(n3142), .B2(n4212), .A(n3141), .ZN(n3143) );
  AOI21_X1 U3938 ( .B1(n3968), .B2(n4595), .A(n3143), .ZN(n4598) );
  INV_X1 U3939 ( .A(n4598), .ZN(n3144) );
  AOI21_X1 U3940 ( .B1(n4648), .B2(n4595), .A(n3144), .ZN(n3146) );
  MUX2_X1 U3941 ( .A(n4386), .B(n3146), .S(n4665), .Z(n3145) );
  OAI21_X1 U3942 ( .B1(n4593), .B2(n4251), .A(n3145), .ZN(U3526) );
  INV_X1 U3943 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3147) );
  MUX2_X1 U3944 ( .A(n3147), .B(n3146), .S(n4658), .Z(n3148) );
  OAI21_X1 U3945 ( .B1(n4593), .B2(n4466), .A(n3148), .ZN(U3483) );
  NOR2_X1 U3946 ( .A1(n3175), .A2(n4232), .ZN(n3149) );
  AOI21_X1 U3947 ( .B1(n4096), .B2(n4235), .A(n3149), .ZN(n3150) );
  OAI211_X1 U3948 ( .C1(n3152), .C2(n4238), .A(n3151), .B(n3150), .ZN(n3153)
         );
  AOI21_X1 U3949 ( .B1(n3154), .B2(n4651), .A(n3153), .ZN(n3156) );
  MUX2_X1 U3950 ( .A(n3038), .B(n3156), .S(n4665), .Z(n3155) );
  OAI21_X1 U3951 ( .B1(n4251), .B2(n3159), .A(n3155), .ZN(U3527) );
  INV_X1 U3952 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3157) );
  MUX2_X1 U3953 ( .A(n3157), .B(n3156), .S(n4658), .Z(n3158) );
  OAI21_X1 U3954 ( .B1(n3159), .B2(n4466), .A(n3158), .ZN(U3485) );
  NAND2_X1 U3955 ( .A1(n3750), .A2(n2957), .ZN(n3162) );
  NAND2_X1 U3956 ( .A1(n3160), .A2(n3410), .ZN(n3161) );
  NAND2_X1 U3957 ( .A1(n3162), .A2(n3161), .ZN(n3163) );
  XNOR2_X1 U3958 ( .A(n3163), .B(n3413), .ZN(n3196) );
  NOR2_X1 U3959 ( .A1(n3175), .A2(n3415), .ZN(n3164) );
  AOI21_X1 U3960 ( .B1(n3750), .B2(n3417), .A(n3164), .ZN(n3195) );
  XNOR2_X1 U3961 ( .A(n3196), .B(n3195), .ZN(n3173) );
  OAI21_X1 U3962 ( .B1(n3167), .B2(n3166), .A(n3165), .ZN(n3169) );
  NAND2_X1 U3963 ( .A1(n3167), .A2(n3166), .ZN(n3168) );
  NAND2_X1 U3964 ( .A1(n3169), .A2(n3168), .ZN(n3170) );
  INV_X1 U3965 ( .A(n3173), .ZN(n3171) );
  INV_X1 U3966 ( .A(n3204), .ZN(n3172) );
  AOI21_X1 U3967 ( .B1(n3173), .B2(n3170), .A(n3172), .ZN(n3180) );
  AND2_X1 U3968 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4503) );
  OAI22_X1 U3969 ( .A1(n3577), .A2(n3175), .B1(n3174), .B2(n3576), .ZN(n3176)
         );
  AOI211_X1 U3970 ( .C1(n3579), .C2(n3751), .A(n4503), .B(n3176), .ZN(n3179)
         );
  NAND2_X1 U3971 ( .A1(n3580), .A2(n3177), .ZN(n3178) );
  OAI211_X1 U3972 ( .C1(n3180), .C2(n3583), .A(n3179), .B(n3178), .ZN(U3228)
         );
  NAND2_X1 U3973 ( .A1(n3197), .A2(n4200), .ZN(n3182) );
  NAND2_X1 U3974 ( .A1(n3750), .A2(n4224), .ZN(n3181) );
  OAI211_X1 U3975 ( .C1(n4239), .C2(n4219), .A(n3182), .B(n3181), .ZN(n3183)
         );
  AOI21_X1 U3976 ( .B1(n3184), .B2(n4047), .A(n3183), .ZN(n3187) );
  NAND2_X1 U3977 ( .A1(n3185), .A2(n4651), .ZN(n3186) );
  NAND2_X1 U3978 ( .A1(n3187), .A2(n3186), .ZN(n3190) );
  MUX2_X1 U3979 ( .A(n3190), .B(REG1_REG_10__SCAN_IN), .S(n4662), .Z(n3188) );
  AOI21_X1 U3980 ( .B1(n4246), .B2(n3192), .A(n3188), .ZN(n3189) );
  INV_X1 U3981 ( .A(n3189), .ZN(U3528) );
  MUX2_X1 U3982 ( .A(n3190), .B(REG0_REG_10__SCAN_IN), .S(n4656), .Z(n3191) );
  AOI21_X1 U3983 ( .B1(n3192), .B2(n4460), .A(n3191), .ZN(n3193) );
  INV_X1 U3984 ( .A(n3193), .ZN(U3487) );
  INV_X1 U3985 ( .A(n3194), .ZN(n3212) );
  NAND2_X1 U3986 ( .A1(n3196), .A2(n3195), .ZN(n3202) );
  AND2_X1 U3987 ( .A1(n3204), .A2(n3202), .ZN(n3206) );
  NAND2_X1 U3988 ( .A1(n4096), .A2(n2957), .ZN(n3199) );
  NAND2_X1 U3989 ( .A1(n3197), .A2(n3410), .ZN(n3198) );
  NAND2_X1 U3990 ( .A1(n3199), .A2(n3198), .ZN(n3200) );
  XNOR2_X1 U3991 ( .A(n3200), .B(n3457), .ZN(n3257) );
  NOR2_X1 U3992 ( .A1(n3208), .A2(n3415), .ZN(n3201) );
  AOI21_X1 U3993 ( .B1(n4096), .B2(n3417), .A(n3201), .ZN(n3255) );
  XNOR2_X1 U3994 ( .A(n3257), .B(n3255), .ZN(n3205) );
  AND2_X1 U3995 ( .A1(n3205), .A2(n3202), .ZN(n3203) );
  OAI211_X1 U3996 ( .C1(n3206), .C2(n3205), .A(n3545), .B(n3258), .ZN(n3211)
         );
  INV_X1 U3997 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3207) );
  NOR2_X1 U3998 ( .A1(STATE_REG_SCAN_IN), .A2(n3207), .ZN(n4512) );
  OAI22_X1 U3999 ( .A1(n3577), .A2(n3208), .B1(n4239), .B2(n3576), .ZN(n3209)
         );
  AOI211_X1 U4000 ( .C1(n3579), .C2(n3750), .A(n4512), .B(n3209), .ZN(n3210)
         );
  OAI211_X1 U4001 ( .C1(n3213), .C2(n3212), .A(n3211), .B(n3210), .ZN(U3214)
         );
  INV_X1 U4002 ( .A(n3214), .ZN(n3216) );
  OR2_X1 U4003 ( .A1(n3216), .A2(n3215), .ZN(n3661) );
  XOR2_X1 U4004 ( .A(n3661), .B(n3217), .Z(n4226) );
  INV_X1 U4005 ( .A(n3218), .ZN(n3219) );
  OR2_X1 U4006 ( .A1(n4086), .A2(n3219), .ZN(n3221) );
  NAND2_X1 U4007 ( .A1(n3221), .A2(n3220), .ZN(n3244) );
  INV_X1 U4008 ( .A(n3233), .ZN(n3222) );
  AOI21_X1 U4009 ( .B1(n3244), .B2(n3234), .A(n3222), .ZN(n3223) );
  XNOR2_X1 U4010 ( .A(n3223), .B(n3661), .ZN(n3224) );
  NOR2_X1 U4011 ( .A1(n3224), .A2(n4212), .ZN(n4221) );
  OR2_X1 U4012 ( .A1(n3236), .A2(n4218), .ZN(n3225) );
  NAND2_X1 U4013 ( .A1(n3286), .A2(n3225), .ZN(n4457) );
  INV_X1 U4014 ( .A(n3538), .ZN(n3226) );
  OAI22_X1 U4015 ( .A1(n4591), .A2(n4398), .B1(n3226), .B2(n4588), .ZN(n3227)
         );
  AOI21_X1 U4016 ( .B1(n4075), .B2(n4223), .A(n3227), .ZN(n3229) );
  AOI22_X1 U4017 ( .A1(n4074), .A2(n4073), .B1(n4059), .B2(n3328), .ZN(n3228)
         );
  OAI211_X1 U4018 ( .C1(n4457), .C2(n4106), .A(n3229), .B(n3228), .ZN(n3230)
         );
  AOI21_X1 U4019 ( .B1(n4221), .B2(n4591), .A(n3230), .ZN(n3231) );
  OAI21_X1 U4020 ( .B1(n4226), .B2(n4084), .A(n3231), .ZN(U3277) );
  AND2_X1 U4021 ( .A1(n3234), .A2(n3233), .ZN(n3655) );
  INV_X1 U4022 ( .A(n3655), .ZN(n3243) );
  XNOR2_X1 U4023 ( .A(n3232), .B(n3243), .ZN(n4231) );
  AND2_X1 U4024 ( .A1(n4103), .A2(n3276), .ZN(n3235) );
  NOR2_X1 U4025 ( .A1(n3236), .A2(n3235), .ZN(n4461) );
  NAND2_X1 U4026 ( .A1(n4461), .A2(n4601), .ZN(n3242) );
  INV_X1 U4027 ( .A(n3280), .ZN(n3237) );
  OAI22_X1 U4028 ( .A1(n4591), .A2(n3238), .B1(n3237), .B2(n4588), .ZN(n3239)
         );
  AOI21_X1 U4029 ( .B1(n3276), .B2(n4059), .A(n3239), .ZN(n3241) );
  AOI22_X1 U4030 ( .A1(n3749), .A2(n4075), .B1(n4073), .B2(n4236), .ZN(n3240)
         );
  NAND3_X1 U4031 ( .A1(n3242), .A2(n3241), .A3(n3240), .ZN(n3247) );
  XNOR2_X1 U4032 ( .A(n3244), .B(n3243), .ZN(n3245) );
  NAND2_X1 U4033 ( .A1(n3245), .A2(n4047), .ZN(n4242) );
  NOR2_X1 U4034 ( .A1(n4242), .A2(n4607), .ZN(n3246) );
  AOI211_X1 U4035 ( .C1(n4036), .C2(n4231), .A(n3247), .B(n3246), .ZN(n3248)
         );
  INV_X1 U4036 ( .A(n3248), .ZN(U3278) );
  OAI22_X1 U4037 ( .A1(n4239), .A2(n3421), .B1(n4088), .B2(n3456), .ZN(n3249)
         );
  XNOR2_X1 U4038 ( .A(n3249), .B(n3413), .ZN(n3254) );
  INV_X1 U4039 ( .A(n3254), .ZN(n3252) );
  NOR2_X1 U4040 ( .A1(n4088), .A2(n3415), .ZN(n3250) );
  AOI21_X1 U4041 ( .B1(n3749), .B2(n3417), .A(n3250), .ZN(n3253) );
  INV_X1 U4042 ( .A(n3253), .ZN(n3251) );
  NAND2_X1 U40430 ( .A1(n3252), .A2(n3251), .ZN(n3268) );
  NAND2_X1 U4044 ( .A1(n3254), .A2(n3253), .ZN(n3266) );
  NAND2_X1 U4045 ( .A1(n3268), .A2(n3266), .ZN(n3259) );
  INV_X1 U4046 ( .A(n3255), .ZN(n3256) );
  XOR2_X1 U4047 ( .A(n3259), .B(n3267), .Z(n3265) );
  NOR2_X1 U4048 ( .A1(STATE_REG_SCAN_IN), .A2(n3260), .ZN(n4523) );
  OAI22_X1 U4049 ( .A1(n3577), .A2(n4088), .B1(n3261), .B2(n3576), .ZN(n3262)
         );
  AOI211_X1 U4050 ( .C1(n3579), .C2(n4096), .A(n4523), .B(n3262), .ZN(n3264)
         );
  NAND2_X1 U4051 ( .A1(n3580), .A2(n4104), .ZN(n3263) );
  OAI211_X1 U4052 ( .C1(n3265), .C2(n3583), .A(n3264), .B(n3263), .ZN(U3233)
         );
  NAND2_X1 U4053 ( .A1(n3267), .A2(n3266), .ZN(n3269) );
  NAND2_X1 U4054 ( .A1(n4223), .A2(n2957), .ZN(n3271) );
  NAND2_X1 U4055 ( .A1(n3276), .A2(n3410), .ZN(n3270) );
  NAND2_X1 U4056 ( .A1(n3271), .A2(n3270), .ZN(n3272) );
  XNOR2_X1 U4057 ( .A(n3272), .B(n3413), .ZN(n3530) );
  INV_X1 U4058 ( .A(n3530), .ZN(n3529) );
  NOR2_X1 U4059 ( .A1(n4233), .A2(n3415), .ZN(n3273) );
  AOI21_X1 U4060 ( .B1(n4223), .B2(n3417), .A(n3273), .ZN(n3532) );
  XNOR2_X1 U4061 ( .A(n3529), .B(n3532), .ZN(n3274) );
  XNOR2_X1 U4062 ( .A(n3338), .B(n3274), .ZN(n3282) );
  AOI22_X1 U4063 ( .A1(n3277), .A2(n3276), .B1(n3275), .B2(n4236), .ZN(n3278)
         );
  NAND2_X1 U4064 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4528) );
  OAI211_X1 U4065 ( .C1(n4239), .C2(n3567), .A(n3278), .B(n4528), .ZN(n3279)
         );
  AOI21_X1 U4066 ( .B1(n3280), .B2(n3580), .A(n3279), .ZN(n3281) );
  OAI21_X1 U4067 ( .B1(n3282), .B2(n3583), .A(n3281), .ZN(U3221) );
  XNOR2_X1 U4068 ( .A(n3595), .B(n3285), .ZN(n4213) );
  OAI21_X1 U4069 ( .B1(n3283), .B2(n3285), .A(n3284), .ZN(n4215) );
  NAND2_X1 U4070 ( .A1(n4215), .A2(n4036), .ZN(n3293) );
  INV_X1 U4071 ( .A(n3286), .ZN(n3287) );
  OAI21_X1 U4072 ( .B1(n3287), .B2(n4208), .A(n4070), .ZN(n4453) );
  INV_X1 U4073 ( .A(n4453), .ZN(n3291) );
  AOI22_X1 U4074 ( .A1(n4075), .A2(n4236), .B1(n4073), .B2(n4195), .ZN(n3289)
         );
  AOI22_X1 U4075 ( .A1(n4607), .A2(REG2_REG_14__SCAN_IN), .B1(n3432), .B2(
        n4599), .ZN(n3288) );
  OAI211_X1 U4076 ( .C1(n4208), .C2(n4079), .A(n3289), .B(n3288), .ZN(n3290)
         );
  AOI21_X1 U4077 ( .B1(n3291), .B2(n4601), .A(n3290), .ZN(n3292) );
  OAI211_X1 U4078 ( .C1(n4213), .C2(n3294), .A(n3293), .B(n3292), .ZN(U3276)
         );
  INV_X1 U4079 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3308) );
  INV_X1 U4080 ( .A(n4124), .ZN(n3745) );
  AOI21_X1 U4081 ( .B1(n3297), .B2(n3635), .A(n3296), .ZN(n3298) );
  NAND2_X1 U4082 ( .A1(n2525), .A2(DATAI_29_), .ZN(n3616) );
  XNOR2_X1 U4083 ( .A(n3744), .B(n3616), .ZN(n3665) );
  XNOR2_X1 U4084 ( .A(n3298), .B(n3665), .ZN(n3833) );
  INV_X1 U4085 ( .A(n3618), .ZN(n3299) );
  AOI21_X1 U4086 ( .B1(n3300), .B2(n3299), .A(n3613), .ZN(n3301) );
  XNOR2_X1 U4087 ( .A(n3301), .B(n3665), .ZN(n3305) );
  AOI21_X1 U4088 ( .B1(n4483), .B2(B_REG_SCAN_IN), .A(n4219), .ZN(n3827) );
  INV_X1 U4089 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4090 ( .A1(n3588), .A2(REG1_REG_30__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U4091 ( .A1(n3589), .A2(REG0_REG_30__SCAN_IN), .ZN(n3302) );
  OAI211_X1 U4092 ( .C1(n3590), .C2(n3304), .A(n3303), .B(n3302), .ZN(n3743)
         );
  AOI22_X1 U4093 ( .A1(n3305), .A2(n4047), .B1(n3827), .B2(n3743), .ZN(n3837)
         );
  NAND2_X1 U4094 ( .A1(n3839), .A2(n4200), .ZN(n3306) );
  OAI211_X1 U4095 ( .C1(n4124), .C2(n4238), .A(n3837), .B(n3306), .ZN(n3307)
         );
  AOI21_X1 U4096 ( .B1(n3833), .B2(n4651), .A(n3307), .ZN(n4259) );
  MUX2_X1 U4097 ( .A(n3308), .B(n4259), .S(n4665), .Z(n3311) );
  AOI21_X1 U4098 ( .B1(n3839), .B2(n3309), .A(n4112), .ZN(n4261) );
  NAND2_X1 U4099 ( .A1(n4261), .A2(n4246), .ZN(n3310) );
  NAND2_X1 U4100 ( .A1(n3311), .A2(n3310), .ZN(U3547) );
  INV_X1 U4101 ( .A(DATAI_30_), .ZN(n3586) );
  NAND2_X1 U4102 ( .A1(n3312), .A2(STATE_REG_SCAN_IN), .ZN(n3313) );
  OAI21_X1 U4103 ( .B1(STATE_REG_SCAN_IN), .B2(n3586), .A(n3313), .ZN(U3322)
         );
  INV_X1 U4104 ( .A(n3315), .ZN(n3323) );
  AOI22_X1 U4105 ( .A1(n4073), .A2(n3744), .B1(n4131), .B2(n4075), .ZN(n3319)
         );
  NOR2_X1 U4106 ( .A1(n3102), .A2(n3316), .ZN(n3317) );
  AOI21_X1 U4107 ( .B1(n3469), .B2(n4599), .A(n3317), .ZN(n3318) );
  OAI211_X1 U4108 ( .C1(n3465), .C2(n4079), .A(n3319), .B(n3318), .ZN(n3322)
         );
  NOR2_X1 U4109 ( .A1(n3320), .A2(n4607), .ZN(n3321) );
  AOI211_X1 U4110 ( .C1(n4601), .C2(n3323), .A(n3322), .B(n3321), .ZN(n3324)
         );
  OAI21_X1 U4111 ( .B1(n3314), .B2(n4084), .A(n3324), .ZN(U3262) );
  NAND2_X1 U4112 ( .A1(n4236), .A2(n2957), .ZN(n3326) );
  NAND2_X1 U4113 ( .A1(n3328), .A2(n3410), .ZN(n3325) );
  NAND2_X1 U4114 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  XNOR2_X1 U4115 ( .A(n3327), .B(n3457), .ZN(n3331) );
  NAND2_X1 U4116 ( .A1(n4236), .A2(n3417), .ZN(n3330) );
  NAND2_X1 U4117 ( .A1(n3328), .A2(n2957), .ZN(n3329) );
  NAND2_X1 U4118 ( .A1(n3330), .A2(n3329), .ZN(n3332) );
  NAND2_X1 U4119 ( .A1(n3331), .A2(n3332), .ZN(n3528) );
  OAI21_X1 U4120 ( .B1(n3530), .B2(n3532), .A(n3528), .ZN(n3337) );
  NAND3_X1 U4121 ( .A1(n3528), .A2(n3532), .A3(n3530), .ZN(n3335) );
  INV_X1 U4122 ( .A(n3331), .ZN(n3334) );
  INV_X1 U4123 ( .A(n3332), .ZN(n3333) );
  NAND2_X1 U4124 ( .A1(n3334), .A2(n3333), .ZN(n3527) );
  AND2_X1 U4125 ( .A1(n3335), .A2(n3527), .ZN(n3336) );
  OAI22_X1 U4126 ( .A1(n4220), .A2(n3421), .B1(n3456), .B2(n4208), .ZN(n3339)
         );
  OAI22_X1 U4127 ( .A1(n4220), .A2(n3459), .B1(n3415), .B2(n4208), .ZN(n3428)
         );
  OAI22_X1 U4128 ( .A1(n4209), .A2(n3421), .B1(n3456), .B2(n4080), .ZN(n3341)
         );
  XNOR2_X1 U4129 ( .A(n3341), .B(n3457), .ZN(n3343) );
  NOR2_X1 U4130 ( .A1(n4080), .A2(n3415), .ZN(n3342) );
  AOI21_X1 U4131 ( .B1(n4195), .B2(n3417), .A(n3342), .ZN(n3574) );
  NOR2_X1 U4132 ( .A1(n3490), .A2(n3574), .ZN(n3350) );
  OAI22_X1 U4133 ( .A1(n4031), .A2(n3459), .B1(n4190), .B2(n3421), .ZN(n3346)
         );
  OAI22_X1 U4134 ( .A1(n4031), .A2(n3421), .B1(n4190), .B2(n3456), .ZN(n3345)
         );
  XNOR2_X1 U4135 ( .A(n3345), .B(n3457), .ZN(n3347) );
  XOR2_X1 U4136 ( .A(n3346), .B(n3347), .Z(n3491) );
  NAND2_X1 U4137 ( .A1(n3489), .A2(n3491), .ZN(n3349) );
  OAI21_X1 U4138 ( .B1(n3350), .B2(n3349), .A(n3348), .ZN(n3501) );
  OAI22_X1 U4139 ( .A1(n4191), .A2(n3421), .B1(n4037), .B2(n3456), .ZN(n3351)
         );
  XOR2_X1 U4140 ( .A(n3457), .B(n3351), .Z(n3499) );
  NOR2_X1 U4141 ( .A1(n4037), .A2(n3415), .ZN(n3352) );
  AOI21_X1 U4142 ( .B1(n3748), .B2(n3417), .A(n3352), .ZN(n3498) );
  OAI22_X1 U4143 ( .A1(n4000), .A2(n3421), .B1(n3456), .B2(n3556), .ZN(n3355)
         );
  XNOR2_X1 U4144 ( .A(n3355), .B(n3413), .ZN(n3360) );
  INV_X1 U4145 ( .A(n3360), .ZN(n3358) );
  NOR2_X1 U4146 ( .A1(n3556), .A2(n3415), .ZN(n3356) );
  AOI21_X1 U4147 ( .B1(n4029), .B2(n3417), .A(n3356), .ZN(n3359) );
  INV_X1 U4148 ( .A(n3359), .ZN(n3357) );
  NAND2_X1 U4149 ( .A1(n3358), .A2(n3357), .ZN(n3552) );
  NAND2_X1 U4150 ( .A1(n4172), .A2(n2957), .ZN(n3363) );
  NAND2_X1 U4151 ( .A1(n3361), .A2(n3410), .ZN(n3362) );
  NAND2_X1 U4152 ( .A1(n3363), .A2(n3362), .ZN(n3364) );
  XNOR2_X1 U4153 ( .A(n3364), .B(n3457), .ZN(n3366) );
  OAI22_X1 U4154 ( .A1(n3555), .A2(n3459), .B1(n3415), .B2(n4002), .ZN(n3365)
         );
  XNOR2_X1 U4155 ( .A(n3366), .B(n3365), .ZN(n3445) );
  NAND2_X1 U4156 ( .A1(n3997), .A2(n2957), .ZN(n3368) );
  NAND2_X1 U4157 ( .A1(n4170), .A2(n3410), .ZN(n3367) );
  NAND2_X1 U4158 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  XNOR2_X1 U4159 ( .A(n3369), .B(n3457), .ZN(n3372) );
  NAND2_X1 U4160 ( .A1(n3997), .A2(n3417), .ZN(n3371) );
  NAND2_X1 U4161 ( .A1(n4170), .A2(n2871), .ZN(n3370) );
  NAND2_X1 U4162 ( .A1(n3371), .A2(n3370), .ZN(n3373) );
  NAND2_X1 U4163 ( .A1(n3372), .A2(n3373), .ZN(n3519) );
  NAND2_X1 U4164 ( .A1(n3518), .A2(n3519), .ZN(n3517) );
  INV_X1 U4165 ( .A(n3372), .ZN(n3375) );
  INV_X1 U4166 ( .A(n3373), .ZN(n3374) );
  NAND2_X1 U4167 ( .A1(n3375), .A2(n3374), .ZN(n3521) );
  NAND2_X1 U4168 ( .A1(n3517), .A2(n3521), .ZN(n3475) );
  NAND2_X1 U4169 ( .A1(n4171), .A2(n2957), .ZN(n3377) );
  NAND2_X1 U4170 ( .A1(n4161), .A2(n3410), .ZN(n3376) );
  NAND2_X1 U4171 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  XNOR2_X1 U4172 ( .A(n3378), .B(n3413), .ZN(n3473) );
  NOR2_X1 U4173 ( .A1(n3962), .A2(n3421), .ZN(n3379) );
  AOI21_X1 U4174 ( .B1(n4171), .B2(n3417), .A(n3379), .ZN(n3472) );
  INV_X1 U4175 ( .A(n3473), .ZN(n3381) );
  INV_X1 U4176 ( .A(n3472), .ZN(n3380) );
  OAI22_X1 U4177 ( .A1(n3477), .A2(n3459), .B1(n3415), .B2(n3937), .ZN(n3392)
         );
  NAND2_X1 U4178 ( .A1(n4162), .A2(n2957), .ZN(n3384) );
  NAND2_X1 U4179 ( .A1(n3943), .A2(n3410), .ZN(n3383) );
  NAND2_X1 U4180 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  XNOR2_X1 U4181 ( .A(n3385), .B(n3457), .ZN(n3391) );
  XOR2_X1 U4182 ( .A(n3392), .B(n3391), .Z(n3544) );
  NAND2_X1 U4183 ( .A1(n4142), .A2(n2957), .ZN(n3388) );
  NAND2_X1 U4184 ( .A1(n3386), .A2(n3410), .ZN(n3387) );
  NAND2_X1 U4185 ( .A1(n3388), .A2(n3387), .ZN(n3389) );
  XNOR2_X1 U4186 ( .A(n3389), .B(n3457), .ZN(n3399) );
  NOR2_X1 U4187 ( .A1(n3926), .A2(n3415), .ZN(n3390) );
  AOI21_X1 U4188 ( .B1(n4142), .B2(n3417), .A(n3390), .ZN(n3397) );
  XNOR2_X1 U4189 ( .A(n3399), .B(n3397), .ZN(n3437) );
  INV_X1 U4190 ( .A(n3391), .ZN(n3394) );
  INV_X1 U4191 ( .A(n3392), .ZN(n3393) );
  NAND2_X1 U4192 ( .A1(n3394), .A2(n3393), .ZN(n3438) );
  NOR2_X1 U4193 ( .A1(n3902), .A2(n3415), .ZN(n3396) );
  AOI21_X1 U4194 ( .B1(n3747), .B2(n3417), .A(n3396), .ZN(n3401) );
  INV_X1 U4195 ( .A(n3397), .ZN(n3398) );
  NAND2_X1 U4196 ( .A1(n3399), .A2(n3398), .ZN(n3402) );
  NAND3_X1 U4197 ( .A1(n3436), .A2(n3401), .A3(n3402), .ZN(n3507) );
  OAI22_X1 U4198 ( .A1(n3921), .A2(n3421), .B1(n3456), .B2(n3902), .ZN(n3400)
         );
  XNOR2_X1 U4199 ( .A(n3400), .B(n3457), .ZN(n3510) );
  NAND2_X1 U4200 ( .A1(n3746), .A2(n2957), .ZN(n3405) );
  INV_X1 U4201 ( .A(n3889), .ZN(n3403) );
  NAND2_X1 U4202 ( .A1(n3403), .A2(n3410), .ZN(n3404) );
  NAND2_X1 U4203 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  XNOR2_X1 U4204 ( .A(n3406), .B(n3413), .ZN(n3409) );
  NOR2_X1 U4205 ( .A1(n3889), .A2(n3415), .ZN(n3407) );
  AOI21_X1 U4206 ( .B1(n3746), .B2(n3417), .A(n3407), .ZN(n3408) );
  OR2_X1 U4207 ( .A1(n3409), .A2(n3408), .ZN(n3483) );
  NAND2_X1 U4208 ( .A1(n4122), .A2(n2871), .ZN(n3412) );
  NAND2_X1 U4209 ( .A1(n4130), .A2(n3410), .ZN(n3411) );
  NAND2_X1 U4210 ( .A1(n3412), .A2(n3411), .ZN(n3414) );
  XNOR2_X1 U4211 ( .A(n3414), .B(n3413), .ZN(n3419) );
  NOR2_X1 U4212 ( .A1(n3866), .A2(n3415), .ZN(n3416) );
  AOI21_X1 U4213 ( .B1(n4122), .B2(n3417), .A(n3416), .ZN(n3418) );
  NOR2_X1 U4214 ( .A1(n3419), .A2(n3418), .ZN(n3563) );
  NAND2_X1 U4215 ( .A1(n3419), .A2(n3418), .ZN(n3562) );
  OAI22_X1 U4216 ( .A1(n3869), .A2(n3421), .B1(n3847), .B2(n3456), .ZN(n3420)
         );
  XNOR2_X1 U4217 ( .A(n3420), .B(n3457), .ZN(n3450) );
  OAI22_X1 U4218 ( .A1(n3869), .A2(n3459), .B1(n3847), .B2(n3421), .ZN(n3451)
         );
  XNOR2_X1 U4219 ( .A(n3450), .B(n3451), .ZN(n3454) );
  XNOR2_X1 U4220 ( .A(n3455), .B(n3454), .ZN(n3427) );
  INV_X1 U4221 ( .A(n3849), .ZN(n3425) );
  INV_X1 U4222 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U4223 ( .A1(n4122), .A2(n3579), .ZN(n3422) );
  OAI21_X1 U4224 ( .B1(STATE_REG_SCAN_IN), .B2(n4374), .A(n3422), .ZN(n3424)
         );
  OAI22_X1 U4225 ( .A1(n4124), .A2(n3576), .B1(n3577), .B2(n3847), .ZN(n3423)
         );
  AOI211_X1 U4226 ( .C1(n3425), .C2(n3580), .A(n3424), .B(n3423), .ZN(n3426)
         );
  OAI21_X1 U4227 ( .B1(n3427), .B2(n3583), .A(n3426), .ZN(U3211) );
  XNOR2_X1 U4228 ( .A(n2050), .B(n3428), .ZN(n3429) );
  XNOR2_X1 U4229 ( .A(n3430), .B(n3429), .ZN(n3435) );
  NOR2_X1 U4230 ( .A1(STATE_REG_SCAN_IN), .A2(n4371), .ZN(n4538) );
  OAI22_X1 U4231 ( .A1(n3577), .A2(n4208), .B1(n4209), .B2(n3576), .ZN(n3431)
         );
  AOI211_X1 U4232 ( .C1(n3579), .C2(n4236), .A(n4538), .B(n3431), .ZN(n3434)
         );
  NAND2_X1 U4233 ( .A1(n3580), .A2(n3432), .ZN(n3433) );
  OAI211_X1 U4234 ( .C1(n3435), .C2(n3583), .A(n3434), .B(n3433), .ZN(U3212)
         );
  NAND2_X1 U4235 ( .A1(n3436), .A2(n3545), .ZN(n3443) );
  AOI21_X1 U4236 ( .B1(n3542), .B2(n3438), .A(n3437), .ZN(n3442) );
  OAI22_X1 U4237 ( .A1(n3477), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n4429), 
        .ZN(n3440) );
  OAI22_X1 U4238 ( .A1(n3921), .A2(n3576), .B1(n3577), .B2(n3926), .ZN(n3439)
         );
  AOI211_X1 U4239 ( .C1(n3928), .C2(n3580), .A(n3440), .B(n3439), .ZN(n3441)
         );
  OAI21_X1 U4240 ( .B1(n3443), .B2(n3442), .A(n3441), .ZN(U3213) );
  XOR2_X1 U4241 ( .A(n3445), .B(n3444), .Z(n3449) );
  NAND2_X1 U4242 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3819) );
  OAI21_X1 U4243 ( .B1(n4000), .B2(n3567), .A(n3819), .ZN(n3447) );
  OAI22_X1 U4244 ( .A1(n3577), .A2(n4002), .B1(n4165), .B2(n3576), .ZN(n3446)
         );
  AOI211_X1 U4245 ( .C1(n4003), .C2(n3580), .A(n3447), .B(n3446), .ZN(n3448)
         );
  OAI21_X1 U4246 ( .B1(n3449), .B2(n3583), .A(n3448), .ZN(U3216) );
  INV_X1 U4247 ( .A(n3450), .ZN(n3453) );
  INV_X1 U4248 ( .A(n3451), .ZN(n3452) );
  OAI22_X1 U4249 ( .A1(n4124), .A2(n3421), .B1(n3456), .B2(n3465), .ZN(n3458)
         );
  XNOR2_X1 U4250 ( .A(n3458), .B(n3457), .ZN(n3461) );
  OAI22_X1 U4251 ( .A1(n4124), .A2(n3459), .B1(n3415), .B2(n3465), .ZN(n3460)
         );
  XNOR2_X1 U4252 ( .A(n3461), .B(n3460), .ZN(n3462) );
  NAND2_X1 U4253 ( .A1(n3463), .A2(n3545), .ZN(n3471) );
  OAI22_X1 U4254 ( .A1(n3869), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n3464), 
        .ZN(n3468) );
  OAI22_X1 U4255 ( .A1(n3466), .A2(n3576), .B1(n3577), .B2(n3465), .ZN(n3467)
         );
  AOI211_X1 U4256 ( .C1(n3469), .C2(n3580), .A(n3468), .B(n3467), .ZN(n3470)
         );
  NAND2_X1 U4257 ( .A1(n3471), .A2(n3470), .ZN(U3217) );
  XNOR2_X1 U4258 ( .A(n3473), .B(n3472), .ZN(n3474) );
  XNOR2_X1 U4259 ( .A(n3475), .B(n3474), .ZN(n3481) );
  INV_X1 U4260 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3476) );
  OAI22_X1 U4261 ( .A1(n4165), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n3476), 
        .ZN(n3479) );
  OAI22_X1 U4262 ( .A1(n3577), .A2(n3962), .B1(n3477), .B2(n3576), .ZN(n3478)
         );
  AOI211_X1 U4263 ( .C1(n3959), .C2(n3580), .A(n3479), .B(n3478), .ZN(n3480)
         );
  OAI21_X1 U4264 ( .B1(n3481), .B2(n3583), .A(n3480), .ZN(U3220) );
  NAND2_X1 U4265 ( .A1(n2056), .A2(n3483), .ZN(n3484) );
  XNOR2_X1 U4266 ( .A(n3482), .B(n3484), .ZN(n3488) );
  OAI22_X1 U4267 ( .A1(n3921), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n4336), 
        .ZN(n3486) );
  OAI22_X1 U4268 ( .A1(n3850), .A2(n3576), .B1(n3577), .B2(n3889), .ZN(n3485)
         );
  AOI211_X1 U4269 ( .C1(n3890), .C2(n3580), .A(n3486), .B(n3485), .ZN(n3487)
         );
  OAI21_X1 U4270 ( .B1(n3488), .B2(n3583), .A(n3487), .ZN(U3222) );
  AOI21_X1 U4271 ( .B1(n3574), .B2(n3489), .A(n3490), .ZN(n3492) );
  XNOR2_X1 U4272 ( .A(n3492), .B(n3491), .ZN(n3497) );
  NAND2_X1 U4273 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4554) );
  OAI21_X1 U4274 ( .B1(n4209), .B2(n3567), .A(n4554), .ZN(n3494) );
  OAI22_X1 U4275 ( .A1(n3577), .A2(n4190), .B1(n4191), .B2(n3576), .ZN(n3493)
         );
  AOI211_X1 U4276 ( .C1(n3495), .C2(n3580), .A(n3494), .B(n3493), .ZN(n3496)
         );
  OAI21_X1 U4277 ( .B1(n3497), .B2(n3583), .A(n3496), .ZN(U3223) );
  XNOR2_X1 U4278 ( .A(n3499), .B(n3498), .ZN(n3500) );
  XNOR2_X1 U4279 ( .A(n3501), .B(n3500), .ZN(n3506) );
  INV_X1 U4280 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3502) );
  NOR2_X1 U4281 ( .A1(STATE_REG_SCAN_IN), .A2(n3502), .ZN(n4567) );
  OAI22_X1 U4282 ( .A1(n3577), .A2(n4037), .B1(n4000), .B2(n3576), .ZN(n3503)
         );
  AOI211_X1 U4283 ( .C1(n3579), .C2(n4201), .A(n4567), .B(n3503), .ZN(n3505)
         );
  NAND2_X1 U4284 ( .A1(n3580), .A2(n4038), .ZN(n3504) );
  OAI211_X1 U4285 ( .C1(n3506), .C2(n3583), .A(n3505), .B(n3504), .ZN(U3225)
         );
  INV_X1 U4286 ( .A(n3507), .ZN(n3508) );
  NOR2_X1 U4287 ( .A1(n3509), .A2(n3508), .ZN(n3511) );
  XNOR2_X1 U4288 ( .A(n3511), .B(n3510), .ZN(n3516) );
  INV_X1 U4289 ( .A(n3905), .ZN(n3514) );
  OAI22_X1 U4290 ( .A1(n3906), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n4347), 
        .ZN(n3513) );
  OAI22_X1 U4291 ( .A1(n4145), .A2(n3576), .B1(n3577), .B2(n3902), .ZN(n3512)
         );
  AOI211_X1 U4292 ( .C1(n3514), .C2(n3580), .A(n3513), .B(n3512), .ZN(n3515)
         );
  OAI21_X1 U4293 ( .B1(n3516), .B2(n3583), .A(n3515), .ZN(U3226) );
  INV_X1 U4294 ( .A(n3517), .ZN(n3522) );
  AOI21_X1 U4295 ( .B1(n3521), .B2(n3519), .A(n3518), .ZN(n3520) );
  AOI21_X1 U4296 ( .B1(n3522), .B2(n3521), .A(n3520), .ZN(n3526) );
  OAI22_X1 U4297 ( .A1(n3555), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n4346), 
        .ZN(n3524) );
  OAI22_X1 U4298 ( .A1(n3577), .A2(n3981), .B1(n3547), .B2(n3576), .ZN(n3523)
         );
  AOI211_X1 U4299 ( .C1(n3978), .C2(n3580), .A(n3524), .B(n3523), .ZN(n3525)
         );
  OAI21_X1 U4300 ( .B1(n3526), .B2(n3583), .A(n3525), .ZN(U3230) );
  NAND2_X1 U4301 ( .A1(n3528), .A2(n3527), .ZN(n3535) );
  NOR2_X1 U4302 ( .A1(n3338), .A2(n3529), .ZN(n3533) );
  INV_X1 U4303 ( .A(n3338), .ZN(n3531) );
  OAI22_X1 U4304 ( .A1(n3533), .A2(n3532), .B1(n3531), .B2(n3530), .ZN(n3534)
         );
  XOR2_X1 U4305 ( .A(n3535), .B(n3534), .Z(n3541) );
  OAI22_X1 U4306 ( .A1(n3577), .A2(n4218), .B1(n4220), .B2(n3576), .ZN(n3536)
         );
  AOI211_X1 U4307 ( .C1(n3579), .C2(n4223), .A(n3537), .B(n3536), .ZN(n3540)
         );
  NAND2_X1 U4308 ( .A1(n3580), .A2(n3538), .ZN(n3539) );
  OAI211_X1 U4309 ( .C1(n3541), .C2(n3583), .A(n3540), .B(n3539), .ZN(U3231)
         );
  OAI21_X1 U4310 ( .B1(n3544), .B2(n3543), .A(n3542), .ZN(n3546) );
  NAND2_X1 U4311 ( .A1(n3546), .A2(n3545), .ZN(n3551) );
  INV_X1 U4312 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4338) );
  OAI22_X1 U4313 ( .A1(n3547), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n4338), 
        .ZN(n3549) );
  OAI22_X1 U4314 ( .A1(n3577), .A2(n3937), .B1(n3906), .B2(n3576), .ZN(n3548)
         );
  AOI211_X1 U4315 ( .C1(n3946), .C2(n3580), .A(n3549), .B(n3548), .ZN(n3550)
         );
  NAND2_X1 U4316 ( .A1(n3551), .A2(n3550), .ZN(U3232) );
  NAND2_X1 U4317 ( .A1(n2057), .A2(n3552), .ZN(n3553) );
  XNOR2_X1 U4318 ( .A(n3554), .B(n3553), .ZN(n3561) );
  OAI22_X1 U4319 ( .A1(n3577), .A2(n3556), .B1(n3555), .B2(n3576), .ZN(n3558)
         );
  NAND2_X1 U4320 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U4321 ( .B1(n4191), .B2(n3567), .A(n4574), .ZN(n3557) );
  NOR2_X1 U4322 ( .A1(n3558), .A2(n3557), .ZN(n3560) );
  NAND2_X1 U4323 ( .A1(n3580), .A2(n4021), .ZN(n3559) );
  OAI211_X1 U4324 ( .C1(n3561), .C2(n3583), .A(n3560), .B(n3559), .ZN(U3235)
         );
  NOR2_X1 U4325 ( .A1(n3563), .A2(n2183), .ZN(n3564) );
  XNOR2_X1 U4326 ( .A(n3565), .B(n3564), .ZN(n3572) );
  INV_X1 U4327 ( .A(n3868), .ZN(n3570) );
  INV_X1 U4328 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3566) );
  OAI22_X1 U4329 ( .A1(n4145), .A2(n3567), .B1(STATE_REG_SCAN_IN), .B2(n3566), 
        .ZN(n3569) );
  OAI22_X1 U4330 ( .A1(n3869), .A2(n3576), .B1(n3577), .B2(n3866), .ZN(n3568)
         );
  AOI211_X1 U4331 ( .C1(n3570), .C2(n3580), .A(n3569), .B(n3568), .ZN(n3571)
         );
  OAI21_X1 U4332 ( .B1(n3572), .B2(n3583), .A(n3571), .ZN(U3237) );
  INV_X1 U4333 ( .A(n3490), .ZN(n3573) );
  NAND2_X1 U4334 ( .A1(n3573), .A2(n3489), .ZN(n3575) );
  XNOR2_X1 U4335 ( .A(n3575), .B(n3574), .ZN(n3584) );
  NOR2_X1 U4336 ( .A1(STATE_REG_SCAN_IN), .A2(n2433), .ZN(n4547) );
  OAI22_X1 U4337 ( .A1(n3577), .A2(n4080), .B1(n4031), .B2(n3576), .ZN(n3578)
         );
  AOI211_X1 U4338 ( .C1(n3579), .C2(n4074), .A(n4547), .B(n3578), .ZN(n3582)
         );
  NAND2_X1 U4339 ( .A1(n3580), .A2(n4076), .ZN(n3581) );
  OAI211_X1 U4340 ( .C1(n3584), .C2(n3583), .A(n3582), .B(n3581), .ZN(U3238)
         );
  NOR2_X1 U4341 ( .A1(n3587), .A2(n3585), .ZN(n3826) );
  NOR2_X1 U4342 ( .A1(n3587), .A2(n3586), .ZN(n4118) );
  INV_X1 U4343 ( .A(n4118), .ZN(n3825) );
  NAND2_X1 U4344 ( .A1(n3743), .A2(n3825), .ZN(n3645) );
  NAND2_X1 U4345 ( .A1(n3588), .A2(REG1_REG_31__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4346 ( .A1(n3589), .A2(REG0_REG_31__SCAN_IN), .ZN(n3592) );
  INV_X1 U4347 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3830) );
  OR2_X1 U4348 ( .A1(n3590), .A2(n3830), .ZN(n3591) );
  NAND2_X1 U4349 ( .A1(n3645), .A2(n3828), .ZN(n3629) );
  INV_X1 U4350 ( .A(n3710), .ZN(n3599) );
  NAND2_X1 U4351 ( .A1(n3594), .A2(n3598), .ZN(n3708) );
  NOR3_X1 U4352 ( .A1(n3595), .A2(n3599), .A3(n3708), .ZN(n3597) );
  OAI21_X1 U4353 ( .B1(n3597), .B2(n2158), .A(n3711), .ZN(n3607) );
  INV_X1 U4354 ( .A(n3598), .ZN(n3600) );
  AOI211_X1 U4355 ( .C1(n3602), .C2(n3601), .A(n3600), .B(n3599), .ZN(n3604)
         );
  OAI21_X1 U4356 ( .B1(n3604), .B2(n3603), .A(n3711), .ZN(n3606) );
  AND2_X1 U4357 ( .A1(n3606), .A2(n3605), .ZN(n3714) );
  NAND2_X1 U4358 ( .A1(n3607), .A2(n3714), .ZN(n3610) );
  NOR2_X1 U4359 ( .A1(n3609), .A2(n3608), .ZN(n3718) );
  OAI221_X1 U4360 ( .B1(n3611), .B2(n3717), .C1(n3611), .C2(n3610), .A(n3718), 
        .ZN(n3615) );
  OR2_X1 U4361 ( .A1(n3613), .A2(n3612), .ZN(n3621) );
  INV_X1 U4362 ( .A(n3826), .ZN(n3829) );
  NAND2_X1 U4363 ( .A1(n3828), .A2(n3829), .ZN(n3727) );
  OAI21_X1 U4364 ( .B1(n3743), .B2(n3825), .A(n3727), .ZN(n3659) );
  INV_X1 U4365 ( .A(n3659), .ZN(n3614) );
  OAI21_X1 U4366 ( .B1(n3744), .B2(n3616), .A(n3614), .ZN(n3620) );
  AOI211_X1 U4367 ( .C1(n3858), .C2(n3615), .A(n3621), .B(n3620), .ZN(n3624)
         );
  AND2_X1 U4368 ( .A1(n3744), .A2(n3616), .ZN(n3617) );
  OR2_X1 U4369 ( .A1(n3618), .A2(n3617), .ZN(n3723) );
  INV_X1 U4370 ( .A(n3723), .ZN(n3622) );
  NAND3_X1 U4371 ( .A1(n3666), .A2(n3622), .A3(n3619), .ZN(n3623) );
  AOI21_X1 U4372 ( .B1(n3622), .B2(n3621), .A(n3620), .ZN(n3729) );
  AOI22_X1 U4373 ( .A1(n3624), .A2(n2165), .B1(n3623), .B2(n3729), .ZN(n3625)
         );
  AOI21_X1 U4374 ( .B1(n3626), .B2(n4118), .A(n3625), .ZN(n3627) );
  AOI211_X1 U4375 ( .C1(n3826), .C2(n3629), .A(n3628), .B(n3627), .ZN(n3734)
         );
  NAND2_X1 U4376 ( .A1(n3630), .A2(n3879), .ZN(n3896) );
  NAND2_X1 U4377 ( .A1(n3632), .A2(n3631), .ZN(n3920) );
  NAND4_X1 U4378 ( .A1(n3941), .A2(n4049), .A3(n3633), .A4(n4035), .ZN(n3634)
         );
  NOR4_X1 U4379 ( .A1(n3635), .A2(n3896), .A3(n3920), .A4(n3634), .ZN(n3643)
         );
  AND4_X1 U4380 ( .A1(n3638), .A2(n3637), .A3(n4092), .A4(n3636), .ZN(n3642)
         );
  INV_X1 U4381 ( .A(n3639), .ZN(n3640) );
  INV_X1 U4382 ( .A(n3914), .ZN(n3713) );
  NAND2_X1 U4383 ( .A1(n3713), .A2(n3915), .ZN(n3956) );
  NOR4_X1 U4384 ( .A1(n3640), .A2(n3956), .A3(n2574), .A4(n4068), .ZN(n3641)
         );
  NAND3_X1 U4385 ( .A1(n3643), .A2(n3642), .A3(n3641), .ZN(n3670) );
  XNOR2_X1 U4386 ( .A(n4172), .B(n4002), .ZN(n3993) );
  NAND2_X1 U4387 ( .A1(n3859), .A2(n3644), .ZN(n3881) );
  INV_X1 U4388 ( .A(n3881), .ZN(n3664) );
  OAI21_X1 U4389 ( .B1(n3828), .B2(n3829), .A(n3645), .ZN(n3728) );
  INV_X1 U4390 ( .A(n3646), .ZN(n3652) );
  INV_X1 U4391 ( .A(n3647), .ZN(n3651) );
  INV_X1 U4392 ( .A(n3648), .ZN(n3649) );
  AND4_X1 U4393 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3653)
         );
  AND3_X1 U4394 ( .A1(n3655), .A2(n3654), .A3(n3653), .ZN(n3656) );
  NAND2_X1 U4395 ( .A1(n3657), .A2(n3656), .ZN(n3658) );
  OR2_X1 U4396 ( .A1(n3728), .A2(n3658), .ZN(n3660) );
  NOR3_X1 U4397 ( .A1(n3661), .A2(n3660), .A3(n3659), .ZN(n3663) );
  INV_X1 U4398 ( .A(n4010), .ZN(n4012) );
  NAND4_X1 U4399 ( .A1(n3664), .A2(n3663), .A3(n4012), .A4(n3662), .ZN(n3669)
         );
  INV_X1 U4400 ( .A(n3665), .ZN(n3667) );
  XNOR2_X1 U4401 ( .A(n4122), .B(n3866), .ZN(n3857) );
  INV_X1 U4402 ( .A(n3857), .ZN(n3861) );
  XNOR2_X1 U4403 ( .A(n3997), .B(n4170), .ZN(n3972) );
  NAND4_X1 U4404 ( .A1(n3667), .A2(n3666), .A3(n3861), .A4(n3972), .ZN(n3668)
         );
  NOR4_X1 U4405 ( .A1(n3670), .A2(n3993), .A3(n3669), .A4(n3668), .ZN(n3732)
         );
  NOR2_X1 U4406 ( .A1(n3869), .A2(n4121), .ZN(n3726) );
  INV_X1 U4407 ( .A(n3671), .ZN(n3674) );
  OAI211_X1 U4408 ( .C1(n3674), .C2(n4470), .A(n3673), .B(n3672), .ZN(n3676)
         );
  NAND3_X1 U4409 ( .A1(n3676), .A2(n3675), .A3(n2576), .ZN(n3679) );
  NAND3_X1 U4410 ( .A1(n3679), .A2(n3678), .A3(n3677), .ZN(n3682) );
  NAND3_X1 U4411 ( .A1(n3682), .A2(n3681), .A3(n3680), .ZN(n3685) );
  NAND3_X1 U4412 ( .A1(n3685), .A2(n3684), .A3(n3683), .ZN(n3689) );
  INV_X1 U4413 ( .A(n3686), .ZN(n3687) );
  AOI21_X1 U4414 ( .B1(n3689), .B2(n3688), .A(n3687), .ZN(n3695) );
  NAND2_X1 U4415 ( .A1(n3691), .A2(n3690), .ZN(n3694) );
  OAI211_X1 U4416 ( .C1(n3695), .C2(n3694), .A(n3693), .B(n3692), .ZN(n3698)
         );
  NAND3_X1 U4417 ( .A1(n3698), .A2(n3697), .A3(n3696), .ZN(n3700) );
  NAND2_X1 U4418 ( .A1(n3700), .A2(n3699), .ZN(n3705) );
  INV_X1 U4419 ( .A(n3702), .ZN(n3703) );
  AOI211_X1 U4420 ( .C1(n3705), .C2(n3704), .A(n2171), .B(n3703), .ZN(n3709)
         );
  INV_X1 U4421 ( .A(n3706), .ZN(n3707) );
  NOR3_X1 U4422 ( .A1(n3709), .A2(n3708), .A3(n3707), .ZN(n3712) );
  OAI211_X1 U4423 ( .C1(n3712), .C2(n2158), .A(n3711), .B(n3710), .ZN(n3715)
         );
  NAND3_X1 U4424 ( .A1(n3715), .A2(n3714), .A3(n3713), .ZN(n3716) );
  NAND2_X1 U4425 ( .A1(n3717), .A2(n3716), .ZN(n3721) );
  INV_X1 U4426 ( .A(n3718), .ZN(n3719) );
  AOI211_X1 U4427 ( .C1(n3722), .C2(n3721), .A(n3720), .B(n3719), .ZN(n3725)
         );
  OR4_X1 U4428 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3730) );
  AOI22_X1 U4429 ( .A1(n3730), .A2(n3729), .B1(n3728), .B2(n3727), .ZN(n3731)
         );
  MUX2_X1 U4430 ( .A(n3732), .B(n3731), .S(n2562), .Z(n3733) );
  NOR2_X1 U4431 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  XNOR2_X1 U4432 ( .A(n3735), .B(n3820), .ZN(n3742) );
  NAND2_X1 U4433 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  OAI211_X1 U4434 ( .C1(n3739), .C2(n3741), .A(n3738), .B(B_REG_SCAN_IN), .ZN(
        n3740) );
  OAI21_X1 U4435 ( .B1(n3742), .B2(n3741), .A(n3740), .ZN(U3239) );
  MUX2_X1 U4436 ( .A(n3828), .B(DATAO_REG_31__SCAN_IN), .S(n3757), .Z(U3581)
         );
  MUX2_X1 U4437 ( .A(n3743), .B(DATAO_REG_30__SCAN_IN), .S(n3757), .Z(U3580)
         );
  MUX2_X1 U4438 ( .A(n3744), .B(DATAO_REG_29__SCAN_IN), .S(n3757), .Z(U3579)
         );
  MUX2_X1 U4439 ( .A(DATAO_REG_28__SCAN_IN), .B(n3745), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4440 ( .A(n4131), .B(DATAO_REG_27__SCAN_IN), .S(n3757), .Z(U3577)
         );
  MUX2_X1 U4441 ( .A(n4122), .B(DATAO_REG_26__SCAN_IN), .S(n3757), .Z(U3576)
         );
  MUX2_X1 U4442 ( .A(n3746), .B(DATAO_REG_25__SCAN_IN), .S(n3757), .Z(U3575)
         );
  MUX2_X1 U4443 ( .A(n3747), .B(DATAO_REG_24__SCAN_IN), .S(n3757), .Z(U3574)
         );
  MUX2_X1 U4444 ( .A(n4142), .B(DATAO_REG_23__SCAN_IN), .S(n3757), .Z(U3573)
         );
  MUX2_X1 U4445 ( .A(n4162), .B(DATAO_REG_22__SCAN_IN), .S(n3757), .Z(U3572)
         );
  MUX2_X1 U4446 ( .A(n4171), .B(DATAO_REG_21__SCAN_IN), .S(n3757), .Z(U3571)
         );
  MUX2_X1 U4447 ( .A(n3997), .B(DATAO_REG_20__SCAN_IN), .S(n3757), .Z(U3570)
         );
  MUX2_X1 U4448 ( .A(DATAO_REG_18__SCAN_IN), .B(n4029), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4449 ( .A(DATAO_REG_17__SCAN_IN), .B(n3748), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4450 ( .A(DATAO_REG_16__SCAN_IN), .B(n4201), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4451 ( .A(n4195), .B(DATAO_REG_15__SCAN_IN), .S(n3757), .Z(U3565)
         );
  MUX2_X1 U4452 ( .A(DATAO_REG_14__SCAN_IN), .B(n4074), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4453 ( .A(n4236), .B(DATAO_REG_13__SCAN_IN), .S(n3757), .Z(U3563)
         );
  MUX2_X1 U4454 ( .A(n4223), .B(DATAO_REG_12__SCAN_IN), .S(n3757), .Z(U3562)
         );
  MUX2_X1 U4455 ( .A(DATAO_REG_11__SCAN_IN), .B(n3749), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4456 ( .A(n4096), .B(DATAO_REG_10__SCAN_IN), .S(n3757), .Z(U3560)
         );
  MUX2_X1 U4457 ( .A(n3750), .B(DATAO_REG_9__SCAN_IN), .S(n3757), .Z(U3559) );
  MUX2_X1 U4458 ( .A(DATAO_REG_8__SCAN_IN), .B(n3751), .S(U4043), .Z(U3558) );
  MUX2_X1 U4459 ( .A(DATAO_REG_7__SCAN_IN), .B(n3752), .S(U4043), .Z(U3557) );
  MUX2_X1 U4460 ( .A(n3753), .B(DATAO_REG_6__SCAN_IN), .S(n3757), .Z(U3556) );
  MUX2_X1 U4461 ( .A(DATAO_REG_5__SCAN_IN), .B(n3754), .S(U4043), .Z(U3555) );
  MUX2_X1 U4462 ( .A(DATAO_REG_4__SCAN_IN), .B(n3755), .S(U4043), .Z(U3554) );
  MUX2_X1 U4463 ( .A(n3756), .B(DATAO_REG_3__SCAN_IN), .S(n3757), .Z(U3553) );
  MUX2_X1 U4464 ( .A(DATAO_REG_2__SCAN_IN), .B(n2291), .S(U4043), .Z(U3552) );
  MUX2_X1 U4465 ( .A(DATAO_REG_1__SCAN_IN), .B(n2281), .S(U4043), .Z(U3551) );
  MUX2_X1 U4466 ( .A(n2712), .B(DATAO_REG_0__SCAN_IN), .S(n3757), .Z(U3550) );
  NAND2_X1 U4467 ( .A1(n3783), .A2(n4479), .ZN(n3766) );
  OAI211_X1 U4468 ( .C1(n3759), .C2(n3758), .A(n4526), .B(n3768), .ZN(n3765)
         );
  AOI22_X1 U4469 ( .A1(n4579), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3764) );
  OAI211_X1 U4470 ( .C1(n3762), .C2(n3761), .A(n4581), .B(n3760), .ZN(n3763)
         );
  NAND4_X1 U4471 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(U3241)
         );
  AOI22_X1 U4472 ( .A1(n4579), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3781) );
  MUX2_X1 U4473 ( .A(n2673), .B(REG2_REG_2__SCAN_IN), .S(n3767), .Z(n3770) );
  NAND3_X1 U4474 ( .A1(n3770), .A2(n3769), .A3(n3768), .ZN(n3771) );
  NAND3_X1 U4475 ( .A1(n4526), .A2(n3772), .A3(n3771), .ZN(n3777) );
  OAI211_X1 U4476 ( .C1(n3775), .C2(n3774), .A(n4581), .B(n3773), .ZN(n3776)
         );
  AND2_X1 U4477 ( .A1(n3777), .A2(n3776), .ZN(n3780) );
  OR2_X1 U4478 ( .A1(n4586), .A2(n3778), .ZN(n3779) );
  NAND4_X1 U4479 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(U3242)
         );
  NAND2_X1 U4480 ( .A1(n3783), .A2(n4478), .ZN(n3792) );
  AOI22_X1 U4481 ( .A1(n4579), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3791) );
  OAI211_X1 U4482 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3785), .A(n4581), .B(n3784), 
        .ZN(n3790) );
  XNOR2_X1 U4483 ( .A(n3787), .B(n3786), .ZN(n3788) );
  NAND2_X1 U4484 ( .A1(n4526), .A2(n3788), .ZN(n3789) );
  NAND4_X1 U4485 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(U3243)
         );
  MUX2_X1 U4486 ( .A(n2476), .B(REG2_REG_19__SCAN_IN), .S(n3820), .Z(n3803) );
  INV_X1 U4487 ( .A(n3804), .ZN(n4620) );
  AOI22_X1 U4488 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4620), .B1(n3804), .B2(
        n2468), .ZN(n4577) );
  NOR2_X1 U4489 ( .A1(n4621), .A2(REG2_REG_17__SCAN_IN), .ZN(n3793) );
  AOI21_X1 U4490 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4621), .A(n3793), .ZN(n4565) );
  NOR2_X1 U4491 ( .A1(n2133), .A2(n3797), .ZN(n3798) );
  NAND2_X1 U4492 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4625), .ZN(n3799) );
  OAI21_X1 U4493 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4625), .A(n3799), .ZN(n4544) );
  NOR2_X1 U4494 ( .A1(n4545), .A2(n4544), .ZN(n4543) );
  AOI21_X1 U4495 ( .B1(n4625), .B2(REG2_REG_15__SCAN_IN), .A(n4543), .ZN(n3800) );
  INV_X1 U4496 ( .A(n3811), .ZN(n4624) );
  NAND2_X1 U4497 ( .A1(n3800), .A2(n4624), .ZN(n3801) );
  XNOR2_X1 U4498 ( .A(n3800), .B(n3811), .ZN(n4556) );
  NAND2_X1 U4499 ( .A1(n4556), .A2(n4054), .ZN(n4555) );
  NAND2_X1 U4500 ( .A1(n3801), .A2(n4555), .ZN(n4563) );
  NAND2_X1 U4501 ( .A1(n4565), .A2(n4563), .ZN(n4564) );
  AOI21_X1 U4502 ( .B1(n3804), .B2(REG2_REG_18__SCAN_IN), .A(n4576), .ZN(n3802) );
  XOR2_X1 U4503 ( .A(n3803), .B(n3802), .Z(n3824) );
  INV_X1 U4504 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4505 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3804), .B1(n4620), .B2(
        n3815), .ZN(n4583) );
  INV_X1 U4506 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U4507 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4625), .ZN(n3810) );
  INV_X1 U4508 ( .A(n4625), .ZN(n4553) );
  AOI22_X1 U4509 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4625), .B1(n4553), .B2(
        n4206), .ZN(n4550) );
  NAND2_X1 U4510 ( .A1(n3807), .A2(n3808), .ZN(n3809) );
  NAND2_X1 U4511 ( .A1(n4550), .A2(n4549), .ZN(n4548) );
  NOR2_X1 U4512 ( .A1(n3811), .A2(n3812), .ZN(n3813) );
  AOI22_X1 U4513 ( .A1(n4621), .A2(n3814), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4573), .ZN(n4568) );
  NOR2_X1 U4514 ( .A1(n4569), .A2(n4568), .ZN(n4570) );
  INV_X1 U4515 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3816) );
  MUX2_X1 U4516 ( .A(REG1_REG_19__SCAN_IN), .B(n3816), .S(n3820), .Z(n3817) );
  NAND2_X1 U4517 ( .A1(n4579), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3818) );
  OAI211_X1 U4518 ( .C1(n4586), .C2(n3820), .A(n3819), .B(n3818), .ZN(n3821)
         );
  AOI21_X1 U4519 ( .B1(n3822), .B2(n4581), .A(n3821), .ZN(n3823) );
  OAI21_X1 U4520 ( .B1(n3824), .B2(n4575), .A(n3823), .ZN(U3259) );
  NAND2_X1 U4521 ( .A1(n4112), .A2(n3825), .ZN(n4113) );
  XNOR2_X1 U4522 ( .A(n4113), .B(n3826), .ZN(n4255) );
  NAND2_X1 U4523 ( .A1(n3828), .A2(n3827), .ZN(n4116) );
  OAI21_X1 U4524 ( .B1(n3829), .B2(n4232), .A(n4116), .ZN(n4252) );
  NOR2_X1 U4525 ( .A1(n4591), .A2(n3830), .ZN(n3831) );
  AOI21_X1 U4526 ( .B1(n4252), .B2(n4591), .A(n3831), .ZN(n3832) );
  OAI21_X1 U4527 ( .B1(n4255), .B2(n4106), .A(n3832), .ZN(U3260) );
  INV_X1 U4528 ( .A(n3833), .ZN(n3840) );
  INV_X1 U4529 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3834) );
  OAI22_X1 U4530 ( .A1(n4124), .A2(n4055), .B1(n3834), .B2(n4591), .ZN(n3838)
         );
  INV_X1 U4531 ( .A(n3835), .ZN(n3836) );
  INV_X1 U4532 ( .A(n4127), .ZN(n3856) );
  NAND2_X1 U4533 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  AOI21_X1 U4534 ( .B1(n3845), .B2(n3844), .A(n4212), .ZN(n4126) );
  OAI21_X1 U4535 ( .B1(n3864), .B2(n3847), .A(n3846), .ZN(n4267) );
  OAI22_X1 U4536 ( .A1(n3849), .A2(n4588), .B1(n3848), .B2(n4591), .ZN(n3852)
         );
  OAI22_X1 U4537 ( .A1(n4124), .A2(n4056), .B1(n3850), .B2(n4055), .ZN(n3851)
         );
  AOI211_X1 U4538 ( .C1(n4121), .C2(n4059), .A(n3852), .B(n3851), .ZN(n3853)
         );
  OAI21_X1 U4539 ( .B1(n4267), .B2(n4106), .A(n3853), .ZN(n3854) );
  AOI21_X1 U4540 ( .B1(n4126), .B2(n4591), .A(n3854), .ZN(n3855) );
  OAI21_X1 U4541 ( .B1(n3856), .B2(n4084), .A(n3855), .ZN(U3263) );
  XNOR2_X1 U4542 ( .A(n2040), .B(n3857), .ZN(n4135) );
  INV_X1 U4543 ( .A(n4135), .ZN(n3876) );
  NAND2_X1 U4544 ( .A1(n3880), .A2(n3858), .ZN(n3860) );
  NAND2_X1 U4545 ( .A1(n3860), .A2(n3859), .ZN(n3862) );
  XNOR2_X1 U4546 ( .A(n3862), .B(n3861), .ZN(n3863) );
  NAND2_X1 U4547 ( .A1(n3863), .A2(n4047), .ZN(n4133) );
  INV_X1 U4548 ( .A(n4133), .ZN(n3874) );
  INV_X1 U4549 ( .A(n3864), .ZN(n3865) );
  OAI21_X1 U4550 ( .B1(n3887), .B2(n3866), .A(n3865), .ZN(n4271) );
  OAI22_X1 U4551 ( .A1(n3868), .A2(n4588), .B1(n3867), .B2(n4591), .ZN(n3871)
         );
  OAI22_X1 U4552 ( .A1(n3869), .A2(n4056), .B1(n4145), .B2(n4055), .ZN(n3870)
         );
  AOI211_X1 U4553 ( .C1(n4130), .C2(n4059), .A(n3871), .B(n3870), .ZN(n3872)
         );
  OAI21_X1 U4554 ( .B1(n4271), .B2(n4106), .A(n3872), .ZN(n3873) );
  AOI21_X1 U4555 ( .B1(n3874), .B2(n4591), .A(n3873), .ZN(n3875) );
  OAI21_X1 U4556 ( .B1(n3876), .B2(n4084), .A(n3875), .ZN(U3264) );
  INV_X1 U4557 ( .A(n3877), .ZN(n3878) );
  XOR2_X1 U4558 ( .A(n3881), .B(n3878), .Z(n4138) );
  INV_X1 U4559 ( .A(n4138), .ZN(n3894) );
  NAND2_X1 U4560 ( .A1(n3880), .A2(n3879), .ZN(n3882) );
  XNOR2_X1 U4561 ( .A(n3882), .B(n3881), .ZN(n3883) );
  NAND2_X1 U4562 ( .A1(n3883), .A2(n4047), .ZN(n3886) );
  NOR2_X1 U4563 ( .A1(n3889), .A2(n4232), .ZN(n3884) );
  AOI21_X1 U4564 ( .B1(n4122), .B2(n4235), .A(n3884), .ZN(n3885) );
  OAI211_X1 U4565 ( .C1(n3921), .C2(n4238), .A(n3886), .B(n3885), .ZN(n4137)
         );
  INV_X1 U4566 ( .A(n3887), .ZN(n3888) );
  OAI21_X1 U4567 ( .B1(n3900), .B2(n3889), .A(n3888), .ZN(n4275) );
  AOI22_X1 U4568 ( .A1(n3890), .A2(n4599), .B1(n4607), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n3891) );
  OAI21_X1 U4569 ( .B1(n4275), .B2(n4106), .A(n3891), .ZN(n3892) );
  AOI21_X1 U4570 ( .B1(n4137), .B2(n3102), .A(n3892), .ZN(n3893) );
  OAI21_X1 U4571 ( .B1(n3894), .B2(n4084), .A(n3893), .ZN(U3265) );
  XOR2_X1 U4572 ( .A(n3896), .B(n3895), .Z(n4147) );
  INV_X1 U4573 ( .A(n4147), .ZN(n3913) );
  INV_X1 U4574 ( .A(n3896), .ZN(n3897) );
  XNOR2_X1 U4575 ( .A(n3898), .B(n3897), .ZN(n3899) );
  NAND2_X1 U4576 ( .A1(n3899), .A2(n4047), .ZN(n4144) );
  INV_X1 U4577 ( .A(n4144), .ZN(n3911) );
  INV_X1 U4578 ( .A(n3925), .ZN(n3903) );
  INV_X1 U4579 ( .A(n3900), .ZN(n3901) );
  OAI21_X1 U4580 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(n4279) );
  INV_X1 U4581 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3904) );
  OAI22_X1 U4582 ( .A1(n3905), .A2(n4588), .B1(n4591), .B2(n3904), .ZN(n3908)
         );
  OAI22_X1 U4583 ( .A1(n4145), .A2(n4056), .B1(n3906), .B2(n4055), .ZN(n3907)
         );
  AOI211_X1 U4584 ( .C1(n4141), .C2(n4059), .A(n3908), .B(n3907), .ZN(n3909)
         );
  OAI21_X1 U4585 ( .B1(n4279), .B2(n4106), .A(n3909), .ZN(n3910) );
  AOI21_X1 U4586 ( .B1(n3911), .B2(n3102), .A(n3910), .ZN(n3912) );
  OAI21_X1 U4587 ( .B1(n3913), .B2(n4084), .A(n3912), .ZN(U3266) );
  XNOR2_X1 U4588 ( .A(n2034), .B(n3920), .ZN(n4151) );
  INV_X1 U4589 ( .A(n4151), .ZN(n3933) );
  OR2_X1 U4590 ( .A1(n3953), .A2(n3914), .ZN(n3916) );
  NAND2_X1 U4591 ( .A1(n3916), .A2(n3915), .ZN(n3934) );
  INV_X1 U4592 ( .A(n3917), .ZN(n3918) );
  AOI21_X1 U4593 ( .B1(n3934), .B2(n3941), .A(n3918), .ZN(n3919) );
  XOR2_X1 U4594 ( .A(n3920), .B(n3919), .Z(n3924) );
  OAI22_X1 U4595 ( .A1(n3921), .A2(n4219), .B1(n4232), .B2(n3926), .ZN(n3922)
         );
  AOI21_X1 U4596 ( .B1(n4224), .B2(n4162), .A(n3922), .ZN(n3923) );
  OAI21_X1 U4597 ( .B1(n3924), .B2(n4212), .A(n3923), .ZN(n4150) );
  INV_X1 U4598 ( .A(n3945), .ZN(n3927) );
  OAI21_X1 U4599 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n4283) );
  NOR2_X1 U4600 ( .A1(n4283), .A2(n4106), .ZN(n3931) );
  INV_X1 U4601 ( .A(n3928), .ZN(n3929) );
  OAI22_X1 U4602 ( .A1(n3102), .A2(n4389), .B1(n3929), .B2(n4588), .ZN(n3930)
         );
  AOI211_X1 U4603 ( .C1(n4150), .C2(n4591), .A(n3931), .B(n3930), .ZN(n3932)
         );
  OAI21_X1 U4604 ( .B1(n3933), .B2(n4084), .A(n3932), .ZN(U3267) );
  XNOR2_X1 U4605 ( .A(n3934), .B(n3941), .ZN(n3939) );
  NAND2_X1 U4606 ( .A1(n4171), .A2(n4224), .ZN(n3936) );
  NAND2_X1 U4607 ( .A1(n4142), .A2(n4235), .ZN(n3935) );
  OAI211_X1 U4608 ( .C1(n4232), .C2(n3937), .A(n3936), .B(n3935), .ZN(n3938)
         );
  AOI21_X1 U4609 ( .B1(n3939), .B2(n4047), .A(n3938), .ZN(n4157) );
  NAND2_X1 U4610 ( .A1(n3942), .A2(n3941), .ZN(n4154) );
  NAND3_X1 U4611 ( .A1(n3940), .A2(n4036), .A3(n4154), .ZN(n3952) );
  NAND2_X1 U4612 ( .A1(n3958), .A2(n3943), .ZN(n3944) );
  NAND2_X1 U4613 ( .A1(n3945), .A2(n3944), .ZN(n4287) );
  INV_X1 U4614 ( .A(n4287), .ZN(n3950) );
  INV_X1 U4615 ( .A(n3946), .ZN(n3947) );
  OAI22_X1 U4616 ( .A1(n3102), .A2(n3948), .B1(n3947), .B2(n4588), .ZN(n3949)
         );
  AOI21_X1 U4617 ( .B1(n3950), .B2(n4601), .A(n3949), .ZN(n3951) );
  OAI211_X1 U4618 ( .C1(n4607), .C2(n4157), .A(n3952), .B(n3951), .ZN(U3268)
         );
  XNOR2_X1 U4619 ( .A(n3953), .B(n3956), .ZN(n3954) );
  NAND2_X1 U4620 ( .A1(n3954), .A2(n4047), .ZN(n4164) );
  XOR2_X1 U4621 ( .A(n3956), .B(n3955), .Z(n4167) );
  NAND2_X1 U4622 ( .A1(n4167), .A2(n4036), .ZN(n3966) );
  OAI21_X1 U4623 ( .B1(n3957), .B2(n3962), .A(n3958), .ZN(n4291) );
  INV_X1 U4624 ( .A(n4291), .ZN(n3964) );
  AOI22_X1 U4625 ( .A1(n4075), .A2(n3997), .B1(n4073), .B2(n4162), .ZN(n3961)
         );
  AOI22_X1 U4626 ( .A1(n4607), .A2(REG2_REG_21__SCAN_IN), .B1(n3959), .B2(
        n4599), .ZN(n3960) );
  OAI211_X1 U4627 ( .C1(n3962), .C2(n4079), .A(n3961), .B(n3960), .ZN(n3963)
         );
  AOI21_X1 U4628 ( .B1(n3964), .B2(n4601), .A(n3963), .ZN(n3965) );
  OAI211_X1 U4629 ( .C1(n4607), .C2(n4164), .A(n3966), .B(n3965), .ZN(U3269)
         );
  XNOR2_X1 U4630 ( .A(n3967), .B(n3972), .ZN(n4175) );
  INV_X1 U4631 ( .A(n4175), .ZN(n3969) );
  NAND2_X1 U4632 ( .A1(n3969), .A2(n3968), .ZN(n3976) );
  NAND2_X1 U4633 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  XNOR2_X1 U4634 ( .A(n3973), .B(n3972), .ZN(n3974) );
  NAND2_X1 U4635 ( .A1(n3974), .A2(n4047), .ZN(n3975) );
  NAND2_X1 U4636 ( .A1(n3976), .A2(n3975), .ZN(n4177) );
  NAND2_X1 U4637 ( .A1(n4177), .A2(n3102), .ZN(n3984) );
  INV_X1 U4638 ( .A(n3977), .ZN(n4001) );
  AOI21_X1 U4639 ( .B1(n4170), .B2(n4001), .A(n3957), .ZN(n4294) );
  AOI22_X1 U4640 ( .A1(n4075), .A2(n4172), .B1(n4073), .B2(n4171), .ZN(n3980)
         );
  AOI22_X1 U4641 ( .A1(n4607), .A2(REG2_REG_20__SCAN_IN), .B1(n3978), .B2(
        n4599), .ZN(n3979) );
  OAI211_X1 U4642 ( .C1(n3981), .C2(n4079), .A(n3980), .B(n3979), .ZN(n3982)
         );
  AOI21_X1 U4643 ( .B1(n4294), .B2(n4601), .A(n3982), .ZN(n3983) );
  OAI211_X1 U4644 ( .C1(n4175), .C2(n3985), .A(n3984), .B(n3983), .ZN(U3270)
         );
  XNOR2_X1 U4645 ( .A(n3986), .B(n3993), .ZN(n4181) );
  INV_X1 U4646 ( .A(n4181), .ZN(n4007) );
  INV_X1 U4647 ( .A(n3987), .ZN(n3989) );
  OAI21_X1 U4648 ( .B1(n4027), .B2(n3989), .A(n3988), .ZN(n4013) );
  INV_X1 U4649 ( .A(n3990), .ZN(n3992) );
  OAI21_X1 U4650 ( .B1(n4013), .B2(n3992), .A(n3991), .ZN(n3994) );
  XNOR2_X1 U4651 ( .A(n3994), .B(n3993), .ZN(n3995) );
  NAND2_X1 U4652 ( .A1(n3995), .A2(n4047), .ZN(n3999) );
  NOR2_X1 U4653 ( .A1(n4002), .A2(n4232), .ZN(n3996) );
  AOI21_X1 U4654 ( .B1(n3997), .B2(n4235), .A(n3996), .ZN(n3998) );
  OAI211_X1 U4655 ( .C1(n4000), .C2(n4238), .A(n3999), .B(n3998), .ZN(n4180)
         );
  OAI21_X1 U4656 ( .B1(n2101), .B2(n4002), .A(n4001), .ZN(n4299) );
  AOI22_X1 U4657 ( .A1(n4607), .A2(REG2_REG_19__SCAN_IN), .B1(n4003), .B2(
        n4599), .ZN(n4004) );
  OAI21_X1 U4658 ( .B1(n4299), .B2(n4106), .A(n4004), .ZN(n4005) );
  AOI21_X1 U4659 ( .B1(n4180), .B2(n4591), .A(n4005), .ZN(n4006) );
  OAI21_X1 U4660 ( .B1(n4007), .B2(n4084), .A(n4006), .ZN(U3271) );
  OAI21_X1 U4661 ( .B1(n4008), .B2(n4010), .A(n4009), .ZN(n4011) );
  INV_X1 U4662 ( .A(n4011), .ZN(n4185) );
  XNOR2_X1 U4663 ( .A(n4013), .B(n4012), .ZN(n4016) );
  AOI22_X1 U4664 ( .A1(n4172), .A2(n4235), .B1(n4017), .B2(n4200), .ZN(n4014)
         );
  OAI21_X1 U4665 ( .B1(n4191), .B2(n4238), .A(n4014), .ZN(n4015) );
  AOI21_X1 U4666 ( .B1(n4016), .B2(n4047), .A(n4015), .ZN(n4184) );
  INV_X1 U4667 ( .A(n4184), .ZN(n4025) );
  AOI21_X1 U4668 ( .B1(n2054), .B2(n4017), .A(n4640), .ZN(n4019) );
  NAND2_X1 U4669 ( .A1(n4019), .A2(n4018), .ZN(n4183) );
  INV_X1 U4670 ( .A(n4020), .ZN(n4023) );
  AOI22_X1 U4671 ( .A1(n4607), .A2(REG2_REG_18__SCAN_IN), .B1(n4021), .B2(
        n4599), .ZN(n4022) );
  OAI21_X1 U4672 ( .B1(n4183), .B2(n4023), .A(n4022), .ZN(n4024) );
  AOI21_X1 U4673 ( .B1(n4025), .B2(n3102), .A(n4024), .ZN(n4026) );
  OAI21_X1 U4674 ( .B1(n4185), .B2(n4084), .A(n4026), .ZN(U3272) );
  XOR2_X1 U4675 ( .A(n4035), .B(n4027), .Z(n4033) );
  AOI22_X1 U4676 ( .A1(n4029), .A2(n4235), .B1(n4200), .B2(n4028), .ZN(n4030)
         );
  OAI21_X1 U4677 ( .B1(n4031), .B2(n4238), .A(n4030), .ZN(n4032) );
  AOI21_X1 U4678 ( .B1(n4033), .B2(n4047), .A(n4032), .ZN(n4187) );
  XNOR2_X1 U4679 ( .A(n4034), .B(n4035), .ZN(n4186) );
  NAND2_X1 U4680 ( .A1(n4186), .A2(n4036), .ZN(n4044) );
  OAI21_X1 U4681 ( .B1(n4052), .B2(n4037), .A(n2054), .ZN(n4189) );
  INV_X1 U4682 ( .A(n4189), .ZN(n4042) );
  INV_X1 U4683 ( .A(n4038), .ZN(n4039) );
  OAI22_X1 U4684 ( .A1(n3102), .A2(n4040), .B1(n4039), .B2(n4588), .ZN(n4041)
         );
  AOI21_X1 U4685 ( .B1(n4042), .B2(n4601), .A(n4041), .ZN(n4043) );
  OAI211_X1 U4686 ( .C1(n4607), .C2(n4187), .A(n4044), .B(n4043), .ZN(U3273)
         );
  OAI21_X1 U4687 ( .B1(n4045), .B2(n2451), .A(n4046), .ZN(n4198) );
  OAI211_X1 U4688 ( .C1(n4050), .C2(n4049), .A(n4048), .B(n4047), .ZN(n4196)
         );
  INV_X1 U4689 ( .A(n4196), .ZN(n4063) );
  NOR2_X1 U4690 ( .A1(n4071), .A2(n4190), .ZN(n4051) );
  OR2_X1 U4691 ( .A1(n4052), .A2(n4051), .ZN(n4192) );
  OAI22_X1 U4692 ( .A1(n3102), .A2(n4054), .B1(n4053), .B2(n4588), .ZN(n4058)
         );
  OAI22_X1 U4693 ( .A1(n4056), .A2(n4191), .B1(n4209), .B2(n4055), .ZN(n4057)
         );
  AOI211_X1 U4694 ( .C1(n4060), .C2(n4059), .A(n4058), .B(n4057), .ZN(n4061)
         );
  OAI21_X1 U4695 ( .B1(n4192), .B2(n4106), .A(n4061), .ZN(n4062) );
  AOI21_X1 U4696 ( .B1(n4063), .B2(n3102), .A(n4062), .ZN(n4064) );
  OAI21_X1 U4697 ( .B1(n4198), .B2(n4084), .A(n4064), .ZN(U3274) );
  XNOR2_X1 U4698 ( .A(n4065), .B(n4068), .ZN(n4205) );
  INV_X1 U4699 ( .A(n4205), .ZN(n4085) );
  INV_X1 U4700 ( .A(n4066), .ZN(n4067) );
  AOI211_X1 U4701 ( .C1(n4069), .C2(n4068), .A(n4212), .B(n4067), .ZN(n4203)
         );
  INV_X1 U4702 ( .A(n4071), .ZN(n4072) );
  OAI21_X1 U4703 ( .B1(n2640), .B2(n4080), .A(n4072), .ZN(n4449) );
  NOR2_X1 U4704 ( .A1(n4449), .A2(n4106), .ZN(n4082) );
  AOI22_X1 U4705 ( .A1(n4075), .A2(n4074), .B1(n4201), .B2(n4073), .ZN(n4078)
         );
  AOI22_X1 U4706 ( .A1(n4607), .A2(REG2_REG_15__SCAN_IN), .B1(n4076), .B2(
        n4599), .ZN(n4077) );
  OAI211_X1 U4707 ( .C1(n4080), .C2(n4079), .A(n4078), .B(n4077), .ZN(n4081)
         );
  AOI211_X1 U4708 ( .C1(n4203), .C2(n4591), .A(n4082), .B(n4081), .ZN(n4083)
         );
  OAI21_X1 U4709 ( .B1(n4085), .B2(n4084), .A(n4083), .ZN(U3275) );
  XOR2_X1 U4710 ( .A(n4092), .B(n4086), .Z(n4098) );
  NAND2_X1 U4711 ( .A1(n4223), .A2(n4235), .ZN(n4087) );
  OAI21_X1 U4712 ( .B1(n4232), .B2(n4088), .A(n4087), .ZN(n4095) );
  INV_X1 U4713 ( .A(n4090), .ZN(n4091) );
  AOI21_X1 U4714 ( .B1(n4092), .B2(n4089), .A(n4091), .ZN(n4099) );
  NOR2_X1 U4715 ( .A1(n4099), .A2(n4093), .ZN(n4094) );
  AOI211_X1 U4716 ( .C1(n4224), .C2(n4096), .A(n4095), .B(n4094), .ZN(n4097)
         );
  OAI21_X1 U4717 ( .B1(n4212), .B2(n4098), .A(n4097), .ZN(n4248) );
  INV_X1 U4718 ( .A(n4248), .ZN(n4109) );
  INV_X1 U4719 ( .A(n4099), .ZN(n4249) );
  NAND2_X1 U4720 ( .A1(n4101), .A2(n4100), .ZN(n4102) );
  NAND2_X1 U4721 ( .A1(n4103), .A2(n4102), .ZN(n4467) );
  AOI22_X1 U4722 ( .A1(n4607), .A2(REG2_REG_11__SCAN_IN), .B1(n4104), .B2(
        n4599), .ZN(n4105) );
  OAI21_X1 U4723 ( .B1(n4467), .B2(n4106), .A(n4105), .ZN(n4107) );
  AOI21_X1 U4724 ( .B1(n4249), .B2(n4602), .A(n4107), .ZN(n4108) );
  OAI21_X1 U4725 ( .B1(n4109), .B2(n4607), .A(n4108), .ZN(U3279) );
  NAND2_X1 U4726 ( .A1(n4252), .A2(n4665), .ZN(n4111) );
  NAND2_X1 U4727 ( .A1(n4662), .A2(REG1_REG_31__SCAN_IN), .ZN(n4110) );
  OAI211_X1 U4728 ( .C1(n4255), .C2(n4251), .A(n4111), .B(n4110), .ZN(U3549)
         );
  INV_X1 U4729 ( .A(n4112), .ZN(n4115) );
  INV_X1 U4730 ( .A(n4113), .ZN(n4114) );
  AOI21_X1 U4731 ( .B1(n4118), .B2(n4115), .A(n4114), .ZN(n4480) );
  INV_X1 U4732 ( .A(n4480), .ZN(n4258) );
  INV_X1 U4733 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4119) );
  INV_X1 U4734 ( .A(n4116), .ZN(n4117) );
  AOI21_X1 U4735 ( .B1(n4118), .B2(n4200), .A(n4117), .ZN(n4482) );
  MUX2_X1 U4736 ( .A(n4119), .B(n4482), .S(n4665), .Z(n4120) );
  OAI21_X1 U4737 ( .B1(n4258), .B2(n4251), .A(n4120), .ZN(U3548) );
  INV_X1 U4738 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U4739 ( .A1(n4122), .A2(n4224), .B1(n4121), .B2(n4200), .ZN(n4123)
         );
  OAI21_X1 U4740 ( .B1(n4124), .B2(n4219), .A(n4123), .ZN(n4125) );
  MUX2_X1 U4741 ( .A(n4128), .B(n4264), .S(n4665), .Z(n4129) );
  OAI21_X1 U4742 ( .B1(n4251), .B2(n4267), .A(n4129), .ZN(U3545) );
  INV_X1 U4743 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4744 ( .A1(n4131), .A2(n4235), .B1(n4200), .B2(n4130), .ZN(n4132)
         );
  OAI211_X1 U4745 ( .C1(n4145), .C2(n4238), .A(n4133), .B(n4132), .ZN(n4134)
         );
  AOI21_X1 U4746 ( .B1(n4135), .B2(n4651), .A(n4134), .ZN(n4268) );
  MUX2_X1 U4747 ( .A(n4428), .B(n4268), .S(n4665), .Z(n4136) );
  OAI21_X1 U4748 ( .B1(n4251), .B2(n4271), .A(n4136), .ZN(U3544) );
  INV_X1 U4749 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4139) );
  AOI21_X1 U4750 ( .B1(n4138), .B2(n4651), .A(n4137), .ZN(n4272) );
  MUX2_X1 U4751 ( .A(n4139), .B(n4272), .S(n4665), .Z(n4140) );
  OAI21_X1 U4752 ( .B1(n4251), .B2(n4275), .A(n4140), .ZN(U3543) );
  INV_X1 U4753 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4754 ( .A1(n4142), .A2(n4224), .B1(n4141), .B2(n4200), .ZN(n4143)
         );
  OAI211_X1 U4755 ( .C1(n4145), .C2(n4219), .A(n4144), .B(n4143), .ZN(n4146)
         );
  AOI21_X1 U4756 ( .B1(n4147), .B2(n4651), .A(n4146), .ZN(n4276) );
  MUX2_X1 U4757 ( .A(n4148), .B(n4276), .S(n4665), .Z(n4149) );
  OAI21_X1 U4758 ( .B1(n4251), .B2(n4279), .A(n4149), .ZN(U3542) );
  INV_X1 U4759 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4152) );
  AOI21_X1 U4760 ( .B1(n4151), .B2(n4651), .A(n4150), .ZN(n4280) );
  MUX2_X1 U4761 ( .A(n4152), .B(n4280), .S(n4665), .Z(n4153) );
  OAI21_X1 U4762 ( .B1(n4251), .B2(n4283), .A(n4153), .ZN(U3541) );
  NAND2_X1 U4763 ( .A1(n4154), .A2(n4651), .ZN(n4156) );
  OR2_X1 U4764 ( .A1(n4156), .A2(n4155), .ZN(n4158) );
  NAND2_X1 U4765 ( .A1(n4158), .A2(n4157), .ZN(n4284) );
  MUX2_X1 U4766 ( .A(REG1_REG_22__SCAN_IN), .B(n4284), .S(n4665), .Z(n4159) );
  INV_X1 U4767 ( .A(n4159), .ZN(n4160) );
  OAI21_X1 U4768 ( .B1(n4251), .B2(n4287), .A(n4160), .ZN(U3540) );
  INV_X1 U4769 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4770 ( .A1(n4162), .A2(n4235), .B1(n4200), .B2(n4161), .ZN(n4163)
         );
  OAI211_X1 U4771 ( .C1(n4165), .C2(n4238), .A(n4164), .B(n4163), .ZN(n4166)
         );
  AOI21_X1 U4772 ( .B1(n4167), .B2(n4651), .A(n4166), .ZN(n4288) );
  MUX2_X1 U4773 ( .A(n4168), .B(n4288), .S(n4665), .Z(n4169) );
  OAI21_X1 U4774 ( .B1(n4251), .B2(n4291), .A(n4169), .ZN(U3539) );
  AOI22_X1 U4775 ( .A1(n4171), .A2(n4235), .B1(n4200), .B2(n4170), .ZN(n4174)
         );
  NAND2_X1 U4776 ( .A1(n4172), .A2(n4224), .ZN(n4173) );
  OAI211_X1 U4777 ( .C1(n4175), .C2(n4641), .A(n4174), .B(n4173), .ZN(n4176)
         );
  OR2_X1 U4778 ( .A1(n4177), .A2(n4176), .ZN(n4292) );
  MUX2_X1 U4779 ( .A(REG1_REG_20__SCAN_IN), .B(n4292), .S(n4665), .Z(n4178) );
  AOI21_X1 U4780 ( .B1(n4246), .B2(n4294), .A(n4178), .ZN(n4179) );
  INV_X1 U4781 ( .A(n4179), .ZN(U3538) );
  AOI21_X1 U4782 ( .B1(n4181), .B2(n4651), .A(n4180), .ZN(n4296) );
  MUX2_X1 U4783 ( .A(n3816), .B(n4296), .S(n4665), .Z(n4182) );
  OAI21_X1 U4784 ( .B1(n4251), .B2(n4299), .A(n4182), .ZN(U3537) );
  OAI211_X1 U4785 ( .C1(n4185), .C2(n4227), .A(n4184), .B(n4183), .ZN(n4300)
         );
  MUX2_X1 U4786 ( .A(REG1_REG_18__SCAN_IN), .B(n4300), .S(n4665), .Z(U3536) );
  NAND2_X1 U4787 ( .A1(n4186), .A2(n4651), .ZN(n4188) );
  OAI211_X1 U4788 ( .C1(n4640), .C2(n4189), .A(n4188), .B(n4187), .ZN(n4301)
         );
  MUX2_X1 U4789 ( .A(n4301), .B(REG1_REG_17__SCAN_IN), .S(n4662), .Z(U3535) );
  OAI22_X1 U4790 ( .A1(n4191), .A2(n4219), .B1(n4190), .B2(n4232), .ZN(n4194)
         );
  NOR2_X1 U4791 ( .A1(n4192), .A2(n4640), .ZN(n4193) );
  AOI211_X1 U4792 ( .C1(n4224), .C2(n4195), .A(n4194), .B(n4193), .ZN(n4197)
         );
  OAI211_X1 U4793 ( .C1(n4198), .C2(n4227), .A(n4197), .B(n4196), .ZN(n4446)
         );
  MUX2_X1 U4794 ( .A(REG1_REG_16__SCAN_IN), .B(n4446), .S(n4665), .Z(U3534) );
  INV_X1 U4795 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U4796 ( .A1(n4201), .A2(n4235), .B1(n4200), .B2(n4199), .ZN(n4202)
         );
  OAI21_X1 U4797 ( .B1(n4220), .B2(n4238), .A(n4202), .ZN(n4204) );
  AOI211_X1 U4798 ( .C1(n4651), .C2(n4205), .A(n4204), .B(n4203), .ZN(n4447)
         );
  MUX2_X1 U4799 ( .A(n4206), .B(n4447), .S(n4665), .Z(n4207) );
  OAI21_X1 U4800 ( .B1(n4251), .B2(n4449), .A(n4207), .ZN(U3533) );
  OAI22_X1 U4801 ( .A1(n4209), .A2(n4219), .B1(n4208), .B2(n4232), .ZN(n4210)
         );
  AOI21_X1 U4802 ( .B1(n4224), .B2(n4236), .A(n4210), .ZN(n4211) );
  OAI21_X1 U4803 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n4214) );
  AOI21_X1 U4804 ( .B1(n4215), .B2(n4651), .A(n4214), .ZN(n4451) );
  INV_X1 U4805 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4216) );
  MUX2_X1 U4806 ( .A(n4451), .B(n4216), .S(n4662), .Z(n4217) );
  OAI21_X1 U4807 ( .B1(n4251), .B2(n4453), .A(n4217), .ZN(U3532) );
  OAI22_X1 U4808 ( .A1(n4220), .A2(n4219), .B1(n4232), .B2(n4218), .ZN(n4222)
         );
  AOI211_X1 U4809 ( .C1(n4224), .C2(n4223), .A(n4222), .B(n4221), .ZN(n4225)
         );
  OAI21_X1 U4810 ( .B1(n4227), .B2(n4226), .A(n4225), .ZN(n4228) );
  INV_X1 U4811 ( .A(n4228), .ZN(n4454) );
  MUX2_X1 U4812 ( .A(n4229), .B(n4454), .S(n4665), .Z(n4230) );
  OAI21_X1 U4813 ( .B1(n4251), .B2(n4457), .A(n4230), .ZN(U3531) );
  NAND2_X1 U4814 ( .A1(n4231), .A2(n4651), .ZN(n4244) );
  NOR2_X1 U4815 ( .A1(n4233), .A2(n4232), .ZN(n4234) );
  AOI21_X1 U4816 ( .B1(n4236), .B2(n4235), .A(n4234), .ZN(n4237) );
  OAI21_X1 U4817 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(n4240) );
  INV_X1 U4818 ( .A(n4240), .ZN(n4241) );
  AND2_X1 U4819 ( .A1(n4242), .A2(n4241), .ZN(n4243) );
  NAND2_X1 U4820 ( .A1(n4244), .A2(n4243), .ZN(n4458) );
  MUX2_X1 U4821 ( .A(n4458), .B(REG1_REG_12__SCAN_IN), .S(n4662), .Z(n4245) );
  AOI21_X1 U4822 ( .B1(n4246), .B2(n4461), .A(n4245), .ZN(n4247) );
  INV_X1 U4823 ( .A(n4247), .ZN(U3530) );
  AOI21_X1 U4824 ( .B1(n4648), .B2(n4249), .A(n4248), .ZN(n4463) );
  MUX2_X1 U4825 ( .A(n3037), .B(n4463), .S(n4665), .Z(n4250) );
  OAI21_X1 U4826 ( .B1(n4251), .B2(n4467), .A(n4250), .ZN(U3529) );
  NAND2_X1 U4827 ( .A1(n4252), .A2(n4658), .ZN(n4254) );
  NAND2_X1 U4828 ( .A1(n4656), .A2(REG0_REG_31__SCAN_IN), .ZN(n4253) );
  OAI211_X1 U4829 ( .C1(n4255), .C2(n4466), .A(n4254), .B(n4253), .ZN(U3517)
         );
  INV_X1 U4830 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4256) );
  MUX2_X1 U4831 ( .A(n4256), .B(n4482), .S(n4658), .Z(n4257) );
  OAI21_X1 U4832 ( .B1(n4258), .B2(n4466), .A(n4257), .ZN(U3516) );
  INV_X1 U4833 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4260) );
  MUX2_X1 U4834 ( .A(n4260), .B(n4259), .S(n4658), .Z(n4263) );
  NAND2_X1 U4835 ( .A1(n4261), .A2(n4460), .ZN(n4262) );
  NAND2_X1 U4836 ( .A1(n4263), .A2(n4262), .ZN(U3515) );
  INV_X1 U4837 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4265) );
  MUX2_X1 U4838 ( .A(n4265), .B(n4264), .S(n4658), .Z(n4266) );
  OAI21_X1 U4839 ( .B1(n4267), .B2(n4466), .A(n4266), .ZN(U3513) );
  INV_X1 U4840 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4269) );
  MUX2_X1 U4841 ( .A(n4269), .B(n4268), .S(n4658), .Z(n4270) );
  OAI21_X1 U4842 ( .B1(n4271), .B2(n4466), .A(n4270), .ZN(U3512) );
  INV_X1 U4843 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4273) );
  MUX2_X1 U4844 ( .A(n4273), .B(n4272), .S(n4658), .Z(n4274) );
  OAI21_X1 U4845 ( .B1(n4275), .B2(n4466), .A(n4274), .ZN(U3511) );
  INV_X1 U4846 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4277) );
  MUX2_X1 U4847 ( .A(n4277), .B(n4276), .S(n4658), .Z(n4278) );
  OAI21_X1 U4848 ( .B1(n4279), .B2(n4466), .A(n4278), .ZN(U3510) );
  INV_X1 U4849 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4281) );
  MUX2_X1 U4850 ( .A(n4281), .B(n4280), .S(n4658), .Z(n4282) );
  OAI21_X1 U4851 ( .B1(n4283), .B2(n4466), .A(n4282), .ZN(U3509) );
  MUX2_X1 U4852 ( .A(REG0_REG_22__SCAN_IN), .B(n4284), .S(n4658), .Z(n4285) );
  INV_X1 U4853 ( .A(n4285), .ZN(n4286) );
  OAI21_X1 U4854 ( .B1(n4287), .B2(n4466), .A(n4286), .ZN(U3508) );
  INV_X1 U4855 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4289) );
  MUX2_X1 U4856 ( .A(n4289), .B(n4288), .S(n4658), .Z(n4290) );
  OAI21_X1 U4857 ( .B1(n4291), .B2(n4466), .A(n4290), .ZN(U3507) );
  MUX2_X1 U4858 ( .A(REG0_REG_20__SCAN_IN), .B(n4292), .S(n4658), .Z(n4293) );
  AOI21_X1 U4859 ( .B1(n4294), .B2(n4460), .A(n4293), .ZN(n4295) );
  INV_X1 U4860 ( .A(n4295), .ZN(U3506) );
  INV_X1 U4861 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4297) );
  MUX2_X1 U4862 ( .A(n4297), .B(n4296), .S(n4658), .Z(n4298) );
  OAI21_X1 U4863 ( .B1(n4299), .B2(n4466), .A(n4298), .ZN(U3505) );
  MUX2_X1 U4864 ( .A(REG0_REG_18__SCAN_IN), .B(n4300), .S(n4658), .Z(U3503) );
  MUX2_X1 U4865 ( .A(n4301), .B(REG0_REG_17__SCAN_IN), .S(n4656), .Z(n4445) );
  NOR4_X1 U4866 ( .A1(keyinput7), .A2(keyinput56), .A3(keyinput25), .A4(
        keyinput0), .ZN(n4307) );
  INV_X1 U4867 ( .A(keyinput62), .ZN(n4302) );
  NOR3_X1 U4868 ( .A1(keyinput52), .A2(keyinput11), .A3(n4302), .ZN(n4306) );
  NAND3_X1 U4869 ( .A1(keyinput48), .A2(keyinput57), .A3(keyinput22), .ZN(
        n4304) );
  NAND3_X1 U4870 ( .A1(keyinput27), .A2(keyinput18), .A3(keyinput6), .ZN(n4303) );
  NOR4_X1 U4871 ( .A1(keyinput63), .A2(keyinput38), .A3(n4304), .A4(n4303), 
        .ZN(n4305) );
  NAND4_X1 U4872 ( .A1(n4307), .A2(keyinput33), .A3(n4306), .A4(n4305), .ZN(
        n4315) );
  NAND3_X1 U4873 ( .A1(keyinput53), .A2(keyinput45), .A3(keyinput24), .ZN(
        n4314) );
  NAND2_X1 U4874 ( .A1(keyinput43), .A2(keyinput8), .ZN(n4308) );
  NOR3_X1 U4875 ( .A1(keyinput14), .A2(keyinput55), .A3(n4308), .ZN(n4312) );
  NOR3_X1 U4876 ( .A1(keyinput32), .A2(keyinput41), .A3(keyinput2), .ZN(n4311)
         );
  NAND2_X1 U4877 ( .A1(keyinput40), .A2(keyinput50), .ZN(n4309) );
  NOR3_X1 U4878 ( .A1(keyinput46), .A2(keyinput39), .A3(n4309), .ZN(n4310) );
  NAND4_X1 U4879 ( .A1(n4312), .A2(keyinput3), .A3(n4311), .A4(n4310), .ZN(
        n4313) );
  NOR4_X1 U4880 ( .A1(keyinput37), .A2(n4315), .A3(n4314), .A4(n4313), .ZN(
        n4331) );
  NOR3_X1 U4881 ( .A1(keyinput34), .A2(keyinput20), .A3(keyinput21), .ZN(n4321) );
  NAND2_X1 U4882 ( .A1(keyinput28), .A2(keyinput5), .ZN(n4316) );
  NOR3_X1 U4883 ( .A1(keyinput29), .A2(keyinput30), .A3(n4316), .ZN(n4320) );
  INV_X1 U4884 ( .A(keyinput13), .ZN(n4318) );
  NAND4_X1 U4885 ( .A1(keyinput10), .A2(keyinput61), .A3(keyinput54), .A4(
        keyinput16), .ZN(n4317) );
  NOR4_X1 U4886 ( .A1(keyinput51), .A2(keyinput12), .A3(n4318), .A4(n4317), 
        .ZN(n4319) );
  NAND4_X1 U4887 ( .A1(keyinput35), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(
        n4329) );
  NAND3_X1 U4888 ( .A1(keyinput15), .A2(keyinput58), .A3(keyinput19), .ZN(
        n4328) );
  NOR3_X1 U4889 ( .A1(keyinput60), .A2(keyinput1), .A3(keyinput47), .ZN(n4326)
         );
  INV_X1 U4890 ( .A(keyinput31), .ZN(n4322) );
  NOR4_X1 U4891 ( .A1(keyinput44), .A2(keyinput26), .A3(keyinput36), .A4(n4322), .ZN(n4325) );
  INV_X1 U4892 ( .A(keyinput4), .ZN(n4323) );
  NOR4_X1 U4893 ( .A1(keyinput49), .A2(keyinput59), .A3(keyinput42), .A4(n4323), .ZN(n4324) );
  NAND4_X1 U4894 ( .A1(keyinput17), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(
        n4327) );
  NOR4_X1 U4895 ( .A1(keyinput23), .A2(n4329), .A3(n4328), .A4(n4327), .ZN(
        n4330) );
  AOI21_X1 U4896 ( .B1(n4331), .B2(n4330), .A(keyinput9), .ZN(n4443) );
  INV_X1 U4897 ( .A(keyinput61), .ZN(n4334) );
  INV_X1 U4898 ( .A(keyinput54), .ZN(n4333) );
  AOI22_X1 U4899 ( .A1(n4334), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n4333), .ZN(n4332) );
  OAI221_X1 U4900 ( .B1(n4334), .B2(DATAO_REG_6__SCAN_IN), .C1(n4333), .C2(
        DATAO_REG_1__SCAN_IN), .A(n4332), .ZN(n4344) );
  AOI22_X1 U4901 ( .A1(n4336), .A2(keyinput13), .B1(keyinput10), .B2(n2533), 
        .ZN(n4335) );
  OAI221_X1 U4902 ( .B1(n4336), .B2(keyinput13), .C1(n2533), .C2(keyinput10), 
        .A(n4335), .ZN(n4343) );
  AOI22_X1 U4903 ( .A1(n4338), .A2(keyinput20), .B1(keyinput35), .B2(n3904), 
        .ZN(n4337) );
  OAI221_X1 U4904 ( .B1(n4338), .B2(keyinput20), .C1(n3904), .C2(keyinput35), 
        .A(n4337), .ZN(n4342) );
  INV_X1 U4905 ( .A(keyinput52), .ZN(n4340) );
  AOI22_X1 U4906 ( .A1(n4289), .A2(keyinput11), .B1(DATAO_REG_17__SCAN_IN), 
        .B2(n4340), .ZN(n4339) );
  OAI221_X1 U4907 ( .B1(n4289), .B2(keyinput11), .C1(n4340), .C2(
        DATAO_REG_17__SCAN_IN), .A(n4339), .ZN(n4341) );
  OR4_X1 U4908 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(n4352) );
  OAI22_X1 U4909 ( .A1(n4347), .A2(keyinput16), .B1(n4346), .B2(keyinput34), 
        .ZN(n4345) );
  AOI221_X1 U4910 ( .B1(n4347), .B2(keyinput16), .C1(keyinput34), .C2(n4346), 
        .A(n4345), .ZN(n4349) );
  XOR2_X1 U4911 ( .A(n2476), .B(keyinput51), .Z(n4348) );
  OAI211_X1 U4912 ( .C1(keyinput9), .C2(n4350), .A(n4349), .B(n4348), .ZN(
        n4351) );
  NOR2_X1 U4913 ( .A1(n4352), .A2(n4351), .ZN(n4441) );
  INV_X1 U4914 ( .A(keyinput22), .ZN(n4354) );
  OAI22_X1 U4915 ( .A1(n2112), .A2(keyinput57), .B1(n4354), .B2(
        ADDR_REG_2__SCAN_IN), .ZN(n4353) );
  AOI221_X1 U4916 ( .B1(n2112), .B2(keyinput57), .C1(ADDR_REG_2__SCAN_IN), 
        .C2(n4354), .A(n4353), .ZN(n4365) );
  INV_X1 U4917 ( .A(keyinput63), .ZN(n4356) );
  OAI22_X1 U4918 ( .A1(n2980), .A2(keyinput27), .B1(n4356), .B2(
        ADDR_REG_5__SCAN_IN), .ZN(n4355) );
  AOI221_X1 U4919 ( .B1(n2980), .B2(keyinput27), .C1(ADDR_REG_5__SCAN_IN), 
        .C2(n4356), .A(n4355), .ZN(n4364) );
  INV_X1 U4920 ( .A(keyinput18), .ZN(n4359) );
  INV_X1 U4921 ( .A(keyinput38), .ZN(n4358) );
  OAI22_X1 U4922 ( .A1(n4359), .A2(ADDR_REG_10__SCAN_IN), .B1(n4358), .B2(
        ADDR_REG_11__SCAN_IN), .ZN(n4357) );
  AOI221_X1 U4923 ( .B1(n4359), .B2(ADDR_REG_10__SCAN_IN), .C1(
        ADDR_REG_11__SCAN_IN), .C2(n4358), .A(n4357), .ZN(n4363) );
  INV_X1 U4924 ( .A(keyinput6), .ZN(n4361) );
  OAI22_X1 U4925 ( .A1(n4229), .A2(keyinput7), .B1(n4361), .B2(
        REG2_REG_12__SCAN_IN), .ZN(n4360) );
  AOI221_X1 U4926 ( .B1(n4229), .B2(keyinput7), .C1(REG2_REG_12__SCAN_IN), 
        .C2(n4361), .A(n4360), .ZN(n4362) );
  NAND4_X1 U4927 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4381)
         );
  INV_X1 U4928 ( .A(D_REG_8__SCAN_IN), .ZN(n4612) );
  INV_X1 U4929 ( .A(D_REG_2__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U4930 ( .A1(n4612), .A2(keyinput14), .B1(keyinput43), .B2(n4615), 
        .ZN(n4366) );
  OAI221_X1 U4931 ( .B1(n4612), .B2(keyinput14), .C1(n4615), .C2(keyinput43), 
        .A(n4366), .ZN(n4380) );
  INV_X1 U4932 ( .A(DATAI_18_), .ZN(n4619) );
  AOI22_X1 U4933 ( .A1(n4368), .A2(keyinput30), .B1(keyinput48), .B2(n4619), 
        .ZN(n4367) );
  OAI221_X1 U4934 ( .B1(n4368), .B2(keyinput30), .C1(n4619), .C2(keyinput48), 
        .A(n4367), .ZN(n4379) );
  AOI22_X1 U4935 ( .A1(n2343), .A2(keyinput0), .B1(n2426), .B2(keyinput33), 
        .ZN(n4369) );
  OAI221_X1 U4936 ( .B1(n2343), .B2(keyinput0), .C1(n2426), .C2(keyinput33), 
        .A(n4369), .ZN(n4377) );
  AOI22_X1 U4937 ( .A1(n4371), .A2(keyinput12), .B1(n2241), .B2(keyinput40), 
        .ZN(n4370) );
  OAI221_X1 U4938 ( .B1(n4371), .B2(keyinput12), .C1(n2241), .C2(keyinput40), 
        .A(n4370), .ZN(n4376) );
  AOI22_X1 U4939 ( .A1(n4374), .A2(keyinput3), .B1(n4373), .B2(keyinput50), 
        .ZN(n4372) );
  OAI221_X1 U4940 ( .B1(n4374), .B2(keyinput3), .C1(n4373), .C2(keyinput50), 
        .A(n4372), .ZN(n4375) );
  OR3_X1 U4941 ( .A1(n4377), .A2(n4376), .A3(n4375), .ZN(n4378) );
  NOR4_X1 U4942 ( .A1(n4381), .A2(n4380), .A3(n4379), .A4(n4378), .ZN(n4440)
         );
  INV_X1 U4943 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4384) );
  INV_X1 U4944 ( .A(DATAI_4_), .ZN(n4383) );
  OAI22_X1 U4945 ( .A1(n4384), .A2(keyinput31), .B1(n4383), .B2(keyinput36), 
        .ZN(n4382) );
  AOI221_X1 U4946 ( .B1(n4384), .B2(keyinput31), .C1(keyinput36), .C2(n4383), 
        .A(n4382), .ZN(n4439) );
  AOI22_X1 U4947 ( .A1(n2328), .A2(keyinput59), .B1(n4386), .B2(keyinput42), 
        .ZN(n4385) );
  OAI221_X1 U4948 ( .B1(n2328), .B2(keyinput59), .C1(n4386), .C2(keyinput42), 
        .A(n4385), .ZN(n4391) );
  INV_X1 U4949 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4950 ( .A1(n4389), .A2(keyinput21), .B1(n4388), .B2(keyinput29), 
        .ZN(n4387) );
  OAI221_X1 U4951 ( .B1(n4389), .B2(keyinput21), .C1(n4388), .C2(keyinput29), 
        .A(n4387), .ZN(n4390) );
  NOR2_X1 U4952 ( .A1(n4391), .A2(n4390), .ZN(n4417) );
  AOI22_X1 U4953 ( .A1(n4265), .A2(keyinput19), .B1(n3308), .B2(keyinput60), 
        .ZN(n4392) );
  OAI221_X1 U4954 ( .B1(n4265), .B2(keyinput19), .C1(n3308), .C2(keyinput60), 
        .A(n4392), .ZN(n4396) );
  INV_X1 U4955 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U4956 ( .A1(n4394), .A2(keyinput62), .B1(n4281), .B2(keyinput15), 
        .ZN(n4393) );
  OAI221_X1 U4957 ( .B1(n4394), .B2(keyinput62), .C1(n4281), .C2(keyinput15), 
        .A(n4393), .ZN(n4395) );
  NOR2_X1 U4958 ( .A1(n4396), .A2(n4395), .ZN(n4416) );
  INV_X1 U4959 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4960 ( .A1(n4399), .A2(keyinput56), .B1(n4398), .B2(keyinput25), 
        .ZN(n4397) );
  OAI221_X1 U4961 ( .B1(n4399), .B2(keyinput56), .C1(n4398), .C2(keyinput25), 
        .A(n4397), .ZN(n4405) );
  XNOR2_X1 U4962 ( .A(IR_REG_1__SCAN_IN), .B(keyinput26), .ZN(n4403) );
  XNOR2_X1 U4963 ( .A(IR_REG_23__SCAN_IN), .B(keyinput39), .ZN(n4402) );
  XNOR2_X1 U4964 ( .A(IR_REG_13__SCAN_IN), .B(keyinput44), .ZN(n4401) );
  XNOR2_X1 U4965 ( .A(REG0_REG_12__SCAN_IN), .B(keyinput17), .ZN(n4400) );
  NAND4_X1 U4966 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(n4404)
         );
  NOR2_X1 U4967 ( .A1(n4405), .A2(n4404), .ZN(n4415) );
  INV_X1 U4968 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U4969 ( .A1(n2363), .A2(keyinput4), .B1(n4407), .B2(keyinput53), 
        .ZN(n4406) );
  OAI221_X1 U4970 ( .B1(n2363), .B2(keyinput4), .C1(n4407), .C2(keyinput53), 
        .A(n4406), .ZN(n4413) );
  XNOR2_X1 U4971 ( .A(keyinput49), .B(REG0_REG_4__SCAN_IN), .ZN(n4411) );
  XNOR2_X1 U4972 ( .A(IR_REG_29__SCAN_IN), .B(keyinput45), .ZN(n4410) );
  XNOR2_X1 U4973 ( .A(keyinput46), .B(DATAI_29_), .ZN(n4409) );
  XNOR2_X1 U4974 ( .A(keyinput37), .B(REG3_REG_15__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4975 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4412)
         );
  NOR2_X1 U4976 ( .A1(n4413), .A2(n4412), .ZN(n4414) );
  NAND4_X1 U4977 ( .A1(n4417), .A2(n4416), .A3(n4415), .A4(n4414), .ZN(n4437)
         );
  INV_X1 U4978 ( .A(D_REG_31__SCAN_IN), .ZN(n4608) );
  INV_X1 U4979 ( .A(D_REG_6__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U4980 ( .A1(n4608), .A2(keyinput55), .B1(keyinput32), .B2(n4613), 
        .ZN(n4418) );
  OAI221_X1 U4981 ( .B1(n4608), .B2(keyinput55), .C1(n4613), .C2(keyinput32), 
        .A(n4418), .ZN(n4436) );
  INV_X1 U4982 ( .A(D_REG_27__SCAN_IN), .ZN(n4609) );
  INV_X1 U4983 ( .A(D_REG_9__SCAN_IN), .ZN(n4611) );
  AOI22_X1 U4984 ( .A1(n4609), .A2(keyinput24), .B1(keyinput8), .B2(n4611), 
        .ZN(n4419) );
  OAI221_X1 U4985 ( .B1(n4609), .B2(keyinput24), .C1(n4611), .C2(keyinput8), 
        .A(n4419), .ZN(n4435) );
  INV_X1 U4986 ( .A(IR_REG_12__SCAN_IN), .ZN(n4422) );
  INV_X1 U4987 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U4988 ( .A1(n4422), .A2(keyinput1), .B1(keyinput47), .B2(n4421), 
        .ZN(n4420) );
  OAI221_X1 U4989 ( .B1(n4422), .B2(keyinput1), .C1(n4421), .C2(keyinput47), 
        .A(n4420), .ZN(n4433) );
  INV_X1 U4990 ( .A(D_REG_16__SCAN_IN), .ZN(n4610) );
  AOI22_X1 U4991 ( .A1(n4610), .A2(keyinput41), .B1(keyinput2), .B2(n4424), 
        .ZN(n4423) );
  OAI221_X1 U4992 ( .B1(n4610), .B2(keyinput41), .C1(n4424), .C2(keyinput2), 
        .A(n4423), .ZN(n4432) );
  INV_X1 U4993 ( .A(DATAI_23_), .ZN(n4618) );
  AOI22_X1 U4994 ( .A1(n4426), .A2(keyinput5), .B1(n4618), .B2(keyinput28), 
        .ZN(n4425) );
  OAI221_X1 U4995 ( .B1(n4426), .B2(keyinput5), .C1(n4618), .C2(keyinput28), 
        .A(n4425), .ZN(n4431) );
  AOI22_X1 U4996 ( .A1(n4429), .A2(keyinput58), .B1(keyinput23), .B2(n4428), 
        .ZN(n4427) );
  OAI221_X1 U4997 ( .B1(n4429), .B2(keyinput58), .C1(n4428), .C2(keyinput23), 
        .A(n4427), .ZN(n4430) );
  OR4_X1 U4998 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4434) );
  NOR4_X1 U4999 ( .A1(n4437), .A2(n4436), .A3(n4435), .A4(n4434), .ZN(n4438)
         );
  AND4_X1 U5000 ( .A1(n4441), .A2(n4440), .A3(n4439), .A4(n4438), .ZN(n4442)
         );
  OAI21_X1 U5001 ( .B1(DATAO_REG_19__SCAN_IN), .B2(n4443), .A(n4442), .ZN(
        n4444) );
  XNOR2_X1 U5002 ( .A(n4445), .B(n4444), .ZN(U3501) );
  MUX2_X1 U5003 ( .A(REG0_REG_16__SCAN_IN), .B(n4446), .S(n4658), .Z(U3499) );
  MUX2_X1 U5004 ( .A(n4407), .B(n4447), .S(n4658), .Z(n4448) );
  OAI21_X1 U5005 ( .B1(n4449), .B2(n4466), .A(n4448), .ZN(U3497) );
  INV_X1 U5006 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U5007 ( .A(n4451), .B(n4450), .S(n4656), .Z(n4452) );
  OAI21_X1 U5008 ( .B1(n4453), .B2(n4466), .A(n4452), .ZN(U3495) );
  INV_X1 U5009 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4455) );
  MUX2_X1 U5010 ( .A(n4455), .B(n4454), .S(n4658), .Z(n4456) );
  OAI21_X1 U5011 ( .B1(n4457), .B2(n4466), .A(n4456), .ZN(U3493) );
  MUX2_X1 U5012 ( .A(n4458), .B(REG0_REG_12__SCAN_IN), .S(n4656), .Z(n4459) );
  AOI21_X1 U5013 ( .B1(n4461), .B2(n4460), .A(n4459), .ZN(n4462) );
  INV_X1 U5014 ( .A(n4462), .ZN(U3491) );
  INV_X1 U5015 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U5016 ( .A(n4464), .B(n4463), .S(n4658), .Z(n4465) );
  OAI21_X1 U5017 ( .B1(n4467), .B2(n4466), .A(n4465), .ZN(U3489) );
  MUX2_X1 U5018 ( .A(n4468), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5019 ( .A(DATAI_25_), .B(n4469), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5020 ( .A(DATAI_21_), .B(n4470), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5021 ( .A(DATAI_20_), .B(n4471), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5022 ( .A(n4472), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5023 ( .A(n4473), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5024 ( .A(n4474), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5025 ( .A(n4475), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5026 ( .A(n4476), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5027 ( .A(DATAI_4_), .B(n4477), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5028 ( .A(n4478), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5029 ( .A(n4479), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5030 ( .A1(n4480), .A2(n4601), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4607), .ZN(n4481) );
  OAI21_X1 U5031 ( .B1(n4607), .B2(n4482), .A(n4481), .ZN(U3261) );
  NOR2_X1 U5032 ( .A1(n4483), .A2(REG1_REG_0__SCAN_IN), .ZN(n4485) );
  NOR2_X1 U5033 ( .A1(n4484), .A2(n4485), .ZN(n4486) );
  MUX2_X1 U5034 ( .A(n4486), .B(n4485), .S(n2112), .Z(n4489) );
  INV_X1 U5035 ( .A(n4487), .ZN(n4488) );
  OR2_X1 U5036 ( .A1(n4489), .A2(n4488), .ZN(n4491) );
  AOI22_X1 U5037 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4579), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4490) );
  OAI21_X1 U5038 ( .B1(n4492), .B2(n4491), .A(n4490), .ZN(U3240) );
  OAI211_X1 U5039 ( .C1(n4495), .C2(n4494), .A(n4581), .B(n4493), .ZN(n4500)
         );
  OAI211_X1 U5040 ( .C1(n4498), .C2(n4497), .A(n4526), .B(n4496), .ZN(n4499)
         );
  OAI211_X1 U5041 ( .C1(n4586), .C2(n4501), .A(n4500), .B(n4499), .ZN(n4502)
         );
  AOI211_X1 U5042 ( .C1(n4579), .C2(ADDR_REG_9__SCAN_IN), .A(n4503), .B(n4502), 
        .ZN(n4504) );
  INV_X1 U5043 ( .A(n4504), .ZN(U3249) );
  OAI211_X1 U5044 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4506), .A(n4581), .B(n4505), .ZN(n4510) );
  OAI211_X1 U5045 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4508), .A(n4526), .B(n4507), .ZN(n4509) );
  OAI211_X1 U5046 ( .C1(n4586), .C2(n4633), .A(n4510), .B(n4509), .ZN(n4511)
         );
  AOI211_X1 U5047 ( .C1(n4579), .C2(ADDR_REG_10__SCAN_IN), .A(n4512), .B(n4511), .ZN(n4513) );
  INV_X1 U5048 ( .A(n4513), .ZN(U3250) );
  OAI211_X1 U5049 ( .C1(n4516), .C2(n4515), .A(n4581), .B(n4514), .ZN(n4521)
         );
  OAI211_X1 U5050 ( .C1(n4519), .C2(n4518), .A(n4526), .B(n4517), .ZN(n4520)
         );
  OAI211_X1 U5051 ( .C1(n4586), .C2(n4631), .A(n4521), .B(n4520), .ZN(n4522)
         );
  AOI211_X1 U5052 ( .C1(n4579), .C2(ADDR_REG_11__SCAN_IN), .A(n4523), .B(n4522), .ZN(n4524) );
  INV_X1 U5053 ( .A(n4524), .ZN(U3251) );
  OAI211_X1 U5054 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4527), .A(n4526), .B(n4525), .ZN(n4529) );
  NAND2_X1 U5055 ( .A1(n4529), .A2(n4528), .ZN(n4530) );
  AOI21_X1 U5056 ( .B1(n4579), .B2(ADDR_REG_12__SCAN_IN), .A(n4530), .ZN(n4534) );
  OAI211_X1 U5057 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4532), .A(n4581), .B(n4531), .ZN(n4533) );
  OAI211_X1 U5058 ( .C1(n4586), .C2(n4629), .A(n4534), .B(n4533), .ZN(U3252)
         );
  AOI211_X1 U5059 ( .C1(n2426), .C2(n4536), .A(n4535), .B(n4575), .ZN(n4537)
         );
  AOI211_X1 U5060 ( .C1(n4579), .C2(ADDR_REG_14__SCAN_IN), .A(n4538), .B(n4537), .ZN(n4542) );
  OAI211_X1 U5061 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4540), .A(n4581), .B(n4539), .ZN(n4541) );
  OAI211_X1 U5062 ( .C1(n4586), .C2(n2133), .A(n4542), .B(n4541), .ZN(U3254)
         );
  AOI211_X1 U5063 ( .C1(n4545), .C2(n4544), .A(n4543), .B(n4575), .ZN(n4546)
         );
  AOI211_X1 U5064 ( .C1(n4579), .C2(ADDR_REG_15__SCAN_IN), .A(n4547), .B(n4546), .ZN(n4552) );
  OAI211_X1 U5065 ( .C1(n4550), .C2(n4549), .A(n4581), .B(n4548), .ZN(n4551)
         );
  OAI211_X1 U5066 ( .C1(n4586), .C2(n4553), .A(n4552), .B(n4551), .ZN(U3255)
         );
  INV_X1 U5067 ( .A(n4554), .ZN(n4558) );
  AOI221_X1 U5068 ( .B1(n4556), .B2(n4555), .C1(n4054), .C2(n4555), .A(n4575), 
        .ZN(n4557) );
  AOI211_X1 U5069 ( .C1(n4579), .C2(ADDR_REG_16__SCAN_IN), .A(n4558), .B(n4557), .ZN(n4562) );
  OAI221_X1 U5070 ( .B1(n4560), .B2(REG1_REG_16__SCAN_IN), .C1(n4560), .C2(
        n4559), .A(n4581), .ZN(n4561) );
  OAI211_X1 U5071 ( .C1(n4586), .C2(n4624), .A(n4562), .B(n4561), .ZN(U3256)
         );
  AOI221_X1 U5072 ( .B1(n4565), .B2(n4564), .C1(n4563), .C2(n4564), .A(n4575), 
        .ZN(n4566) );
  AOI211_X1 U5073 ( .C1(n4579), .C2(ADDR_REG_17__SCAN_IN), .A(n4567), .B(n4566), .ZN(n4572) );
  OAI221_X1 U5074 ( .B1(n4570), .B2(n4569), .C1(n4570), .C2(n4568), .A(n4581), 
        .ZN(n4571) );
  OAI211_X1 U5075 ( .C1(n4586), .C2(n4573), .A(n4572), .B(n4571), .ZN(U3257)
         );
  INV_X1 U5076 ( .A(n4574), .ZN(n4578) );
  OAI211_X1 U5077 ( .C1(n4583), .C2(n4582), .A(n4581), .B(n4580), .ZN(n4584)
         );
  OAI211_X1 U5078 ( .C1(n4586), .C2(n4620), .A(n4585), .B(n4584), .ZN(U3258)
         );
  INV_X1 U5079 ( .A(n4587), .ZN(n4589) );
  OAI22_X1 U5080 ( .A1(n4591), .A2(n4590), .B1(n4589), .B2(n4588), .ZN(n4592)
         );
  INV_X1 U5081 ( .A(n4592), .ZN(n4597) );
  INV_X1 U5082 ( .A(n4593), .ZN(n4594) );
  AOI22_X1 U5083 ( .A1(n4595), .A2(n4602), .B1(n4601), .B2(n4594), .ZN(n4596)
         );
  OAI211_X1 U5084 ( .C1(n4607), .C2(n4598), .A(n4597), .B(n4596), .ZN(U3282)
         );
  AOI22_X1 U5085 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4599), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4607), .ZN(n4605) );
  AOI22_X1 U5086 ( .A1(n4603), .A2(n4602), .B1(n4601), .B2(n4600), .ZN(n4604)
         );
  OAI211_X1 U5087 ( .C1(n4607), .C2(n4606), .A(n4605), .B(n4604), .ZN(U3288)
         );
  NOR2_X1 U5088 ( .A1(n4616), .A2(n4608), .ZN(U3291) );
  AND2_X1 U5089 ( .A1(D_REG_30__SCAN_IN), .A2(n4614), .ZN(U3292) );
  AND2_X1 U5090 ( .A1(D_REG_29__SCAN_IN), .A2(n4614), .ZN(U3293) );
  AND2_X1 U5091 ( .A1(D_REG_28__SCAN_IN), .A2(n4614), .ZN(U3294) );
  NOR2_X1 U5092 ( .A1(n4616), .A2(n4609), .ZN(U3295) );
  AND2_X1 U5093 ( .A1(D_REG_26__SCAN_IN), .A2(n4614), .ZN(U3296) );
  AND2_X1 U5094 ( .A1(D_REG_25__SCAN_IN), .A2(n4614), .ZN(U3297) );
  AND2_X1 U5095 ( .A1(D_REG_24__SCAN_IN), .A2(n4614), .ZN(U3298) );
  AND2_X1 U5096 ( .A1(D_REG_23__SCAN_IN), .A2(n4614), .ZN(U3299) );
  AND2_X1 U5097 ( .A1(D_REG_22__SCAN_IN), .A2(n4614), .ZN(U3300) );
  AND2_X1 U5098 ( .A1(D_REG_21__SCAN_IN), .A2(n4614), .ZN(U3301) );
  AND2_X1 U5099 ( .A1(D_REG_20__SCAN_IN), .A2(n4614), .ZN(U3302) );
  AND2_X1 U5100 ( .A1(D_REG_19__SCAN_IN), .A2(n4614), .ZN(U3303) );
  AND2_X1 U5101 ( .A1(D_REG_18__SCAN_IN), .A2(n4614), .ZN(U3304) );
  AND2_X1 U5102 ( .A1(D_REG_17__SCAN_IN), .A2(n4614), .ZN(U3305) );
  NOR2_X1 U5103 ( .A1(n4616), .A2(n4610), .ZN(U3306) );
  AND2_X1 U5104 ( .A1(D_REG_15__SCAN_IN), .A2(n4614), .ZN(U3307) );
  AND2_X1 U5105 ( .A1(D_REG_14__SCAN_IN), .A2(n4614), .ZN(U3308) );
  AND2_X1 U5106 ( .A1(D_REG_13__SCAN_IN), .A2(n4614), .ZN(U3309) );
  AND2_X1 U5107 ( .A1(D_REG_12__SCAN_IN), .A2(n4614), .ZN(U3310) );
  AND2_X1 U5108 ( .A1(D_REG_11__SCAN_IN), .A2(n4614), .ZN(U3311) );
  AND2_X1 U5109 ( .A1(D_REG_10__SCAN_IN), .A2(n4614), .ZN(U3312) );
  NOR2_X1 U5110 ( .A1(n4616), .A2(n4611), .ZN(U3313) );
  NOR2_X1 U5111 ( .A1(n4616), .A2(n4612), .ZN(U3314) );
  AND2_X1 U5112 ( .A1(D_REG_7__SCAN_IN), .A2(n4614), .ZN(U3315) );
  NOR2_X1 U5113 ( .A1(n4616), .A2(n4613), .ZN(U3316) );
  AND2_X1 U5114 ( .A1(D_REG_5__SCAN_IN), .A2(n4614), .ZN(U3317) );
  AND2_X1 U5115 ( .A1(D_REG_4__SCAN_IN), .A2(n4614), .ZN(U3318) );
  AND2_X1 U5116 ( .A1(D_REG_3__SCAN_IN), .A2(n4614), .ZN(U3319) );
  NOR2_X1 U5117 ( .A1(n4616), .A2(n4615), .ZN(U3320) );
  AOI21_X1 U5118 ( .B1(U3149), .B2(n4618), .A(n4617), .ZN(U3329) );
  AOI22_X1 U5119 ( .A1(STATE_REG_SCAN_IN), .A2(n4620), .B1(n4619), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5120 ( .A1(U3149), .A2(n4621), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4622) );
  INV_X1 U5121 ( .A(n4622), .ZN(U3335) );
  INV_X1 U5122 ( .A(DATAI_16_), .ZN(n4623) );
  AOI22_X1 U5123 ( .A1(STATE_REG_SCAN_IN), .A2(n4624), .B1(n4623), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5124 ( .A1(U3149), .A2(n4625), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4626) );
  INV_X1 U5125 ( .A(n4626), .ZN(U3337) );
  INV_X1 U5126 ( .A(DATAI_14_), .ZN(n4627) );
  AOI22_X1 U5127 ( .A1(STATE_REG_SCAN_IN), .A2(n2133), .B1(n4627), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5128 ( .A(DATAI_12_), .ZN(n4628) );
  AOI22_X1 U5129 ( .A1(STATE_REG_SCAN_IN), .A2(n4629), .B1(n4628), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5130 ( .A(DATAI_11_), .ZN(n4630) );
  AOI22_X1 U5131 ( .A1(STATE_REG_SCAN_IN), .A2(n4631), .B1(n4630), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5132 ( .A(DATAI_10_), .ZN(n4632) );
  AOI22_X1 U5133 ( .A1(STATE_REG_SCAN_IN), .A2(n4633), .B1(n4632), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5134 ( .A1(U3149), .A2(n4634), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4635) );
  INV_X1 U5135 ( .A(n4635), .ZN(U3343) );
  OAI22_X1 U5136 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4636) );
  INV_X1 U5137 ( .A(n4636), .ZN(U3352) );
  INV_X1 U5138 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U5139 ( .A1(n4658), .A2(n4638), .B1(n4637), .B2(n4656), .ZN(U3467)
         );
  OAI22_X1 U5140 ( .A1(n4642), .A2(n4641), .B1(n4640), .B2(n4639), .ZN(n4643)
         );
  NOR2_X1 U5141 ( .A1(n4644), .A2(n4643), .ZN(n4659) );
  INV_X1 U5142 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U5143 ( .A1(n4658), .A2(n4659), .B1(n4645), .B2(n4656), .ZN(U3469)
         );
  AOI211_X1 U5144 ( .C1(n4649), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4661)
         );
  INV_X1 U5145 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U5146 ( .A1(n4658), .A2(n4661), .B1(n4650), .B2(n4656), .ZN(U3475)
         );
  NAND3_X1 U5147 ( .A1(n3081), .A2(n4652), .A3(n4651), .ZN(n4653) );
  AND3_X1 U5148 ( .A1(n4655), .A2(n4654), .A3(n4653), .ZN(n4664) );
  INV_X1 U5149 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5150 ( .A1(n4658), .A2(n4664), .B1(n4657), .B2(n4656), .ZN(U3481)
         );
  AOI22_X1 U5151 ( .A1(n4665), .A2(n4659), .B1(n2684), .B2(n4662), .ZN(U3519)
         );
  AOI22_X1 U5152 ( .A1(n4665), .A2(n4661), .B1(n4660), .B2(n4662), .ZN(U3522)
         );
  AOI22_X1 U5153 ( .A1(n4665), .A2(n4664), .B1(n4663), .B2(n4662), .ZN(U3525)
         );
  CLKBUF_X1 U2268 ( .A(n2296), .Z(n3589) );
endmodule

