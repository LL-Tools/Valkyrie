

module b20_C_SARLock_k_64_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101;

  INV_X4 U4793 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X2 U4794 ( .A(n7034), .ZN(n9854) );
  NAND2_X1 U4795 ( .A1(n5572), .A2(n7684), .ZN(n6313) );
  NAND2_X1 U4796 ( .A1(n8387), .A2(n8342), .ZN(n8310) );
  INV_X1 U4797 ( .A(n5865), .ZN(n5968) );
  INV_X1 U4798 ( .A(n6034), .ZN(n6050) );
  INV_X1 U4799 ( .A(n5865), .ZN(n6052) );
  NOR2_X1 U4800 ( .A1(n4932), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U4801 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4913) );
  OAI21_X1 U4802 ( .B1(n6729), .B2(P2_D_REG_0__SCAN_IN), .A(n6757), .ZN(n6987)
         );
  INV_X1 U4803 ( .A(n8310), .ZN(n8326) );
  NAND2_X1 U4804 ( .A1(n5128), .A2(n9477), .ZN(n5129) );
  INV_X1 U4805 ( .A(n5184), .ZN(n5420) );
  INV_X1 U4806 ( .A(n7456), .ZN(n7131) );
  INV_X1 U4807 ( .A(n6963), .ZN(n9573) );
  AND4_X1 U4808 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n7033)
         );
  NAND2_X1 U4809 ( .A1(n6668), .A2(n6667), .ZN(n6729) );
  NAND2_X1 U4810 ( .A1(n5266), .A2(n5265), .ZN(n9608) );
  AND2_X1 U4811 ( .A1(n5076), .A2(n5101), .ZN(n6316) );
  XNOR2_X1 U4812 ( .A(n5242), .B(n5241), .ZN(n6759) );
  AND3_X1 U4813 ( .A1(n5244), .A2(n4912), .A3(n4911), .ZN(n4286) );
  NAND2_X2 U4814 ( .A1(n7642), .A2(n6117), .ZN(n7829) );
  NAND2_X2 U4815 ( .A1(n4585), .A2(n4583), .ZN(n7642) );
  OAI21_X2 U4816 ( .B1(n7641), .B2(n4459), .A(n4457), .ZN(n7816) );
  NAND2_X2 U4817 ( .A1(n9224), .A2(n6221), .ZN(n9204) );
  NAND2_X2 U4818 ( .A1(n5592), .A2(n4359), .ZN(n9224) );
  NAND2_X2 U4819 ( .A1(n9310), .A2(n6146), .ZN(n9297) );
  NAND2_X2 U4820 ( .A1(n4400), .A2(n9309), .ZN(n9310) );
  OAI211_X2 U4821 ( .C1(n6351), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n4876), .B(
        n4875), .ZN(n6992) );
  NAND2_X2 U4822 ( .A1(n6990), .A2(n6989), .ZN(n7112) );
  OAI222_X1 U4823 ( .A1(n9450), .A2(n8114), .B1(P1_U3086), .B2(n5605), .C1(
        n9452), .C2(n8907), .ZN(P1_U3327) );
  AND2_X4 U4824 ( .A1(n4779), .A2(n4778), .ZN(n6722) );
  INV_X1 U4825 ( .A(n6330), .ZN(n8902) );
  INV_X1 U4826 ( .A(n4910), .ZN(n5430) );
  CLKBUF_X1 U4827 ( .A(n5168), .Z(n4287) );
  BUF_X4 U4828 ( .A(n5168), .Z(n4288) );
  AND2_X2 U4829 ( .A1(n4727), .A2(n9548), .ZN(n9535) );
  OR2_X1 U4830 ( .A1(n9234), .A2(n5491), .ZN(n5493) );
  OAI21_X1 U4831 ( .B1(n9249), .B2(n5475), .A(n4461), .ZN(n9234) );
  AND2_X1 U4832 ( .A1(n8422), .A2(n8145), .ZN(n8485) );
  OAI21_X1 U4833 ( .B1(n8410), .B2(n8134), .A(n8136), .ZN(n8475) );
  NOR2_X2 U4834 ( .A1(n7941), .A2(n7942), .ZN(n5964) );
  AND2_X1 U4835 ( .A1(n5956), .A2(n4313), .ZN(n7942) );
  NAND2_X1 U4836 ( .A1(n7370), .A2(n7371), .ZN(n7529) );
  NAND2_X2 U4837 ( .A1(n8208), .A2(n8236), .ZN(n8357) );
  NAND2_X1 U4838 ( .A1(n4699), .A2(n5580), .ZN(n7317) );
  INV_X1 U4839 ( .A(n9039), .ZN(n5274) );
  INV_X1 U4840 ( .A(n9040), .ZN(n5260) );
  NOR2_X1 U4841 ( .A1(n8529), .A2(n7437), .ZN(n4332) );
  INV_X4 U4842 ( .A(n7795), .ZN(n8161) );
  INV_X1 U4843 ( .A(n5611), .ZN(n5151) );
  CLKBUF_X2 U4845 ( .A(n6615), .Z(n4293) );
  NAND2_X2 U4846 ( .A1(n6034), .A2(n6031), .ZN(n4290) );
  INV_X1 U4847 ( .A(n5854), .ZN(n5865) );
  OR2_X1 U4848 ( .A1(n8317), .A2(n6736), .ZN(n6359) );
  NAND2_X2 U4849 ( .A1(n6034), .A2(n6031), .ZN(n5856) );
  XNOR2_X1 U4850 ( .A(n5182), .B(n5183), .ZN(n6736) );
  CLKBUF_X2 U4851 ( .A(n6351), .Z(n8316) );
  CLKBUF_X1 U4852 ( .A(n9464), .Z(n4294) );
  CLKBUF_X2 U4853 ( .A(n6356), .Z(n4298) );
  CLKBUF_X1 U4854 ( .A(n5117), .Z(n9445) );
  AND2_X1 U4855 ( .A1(n6330), .A2(n6329), .ZN(n6356) );
  NAND2_X2 U4856 ( .A1(n8384), .A2(n6847), .ZN(n6661) );
  INV_X1 U4857 ( .A(n6328), .ZN(n6329) );
  XNOR2_X1 U4858 ( .A(n6327), .B(n6326), .ZN(n6328) );
  XNOR2_X1 U4859 ( .A(n5658), .B(n6323), .ZN(n8384) );
  MUX2_X1 U4860 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5660), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5661) );
  INV_X8 U4861 ( .A(n6722), .ZN(n6717) );
  AND2_X1 U4862 ( .A1(n8603), .A2(n8602), .ZN(n8818) );
  NAND2_X1 U4863 ( .A1(n4718), .A2(n4716), .ZN(n4715) );
  OR2_X1 U4864 ( .A1(n4724), .A2(n6187), .ZN(n4718) );
  AND2_X1 U4865 ( .A1(n8595), .A2(n8594), .ZN(n8819) );
  OR2_X1 U4866 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  OR2_X1 U4867 ( .A1(n8591), .A2(n8590), .ZN(n8595) );
  AND2_X1 U4868 ( .A1(n8628), .A2(n8629), .ZN(n8630) );
  NAND2_X1 U4869 ( .A1(n4405), .A2(n4406), .ZN(n6009) );
  XNOR2_X1 U4870 ( .A(n8333), .B(n4676), .ZN(n8578) );
  INV_X1 U4871 ( .A(n4549), .ZN(n8627) );
  NAND2_X1 U4872 ( .A1(n9264), .A2(n5462), .ZN(n9249) );
  NAND2_X1 U4873 ( .A1(n8485), .A2(n8484), .ZN(n8483) );
  NAND2_X1 U4874 ( .A1(n4768), .A2(n4343), .ZN(n9264) );
  NAND2_X1 U4875 ( .A1(n9291), .A2(n4772), .ZN(n4768) );
  OAI21_X1 U4876 ( .B1(n8672), .B2(n4377), .A(n6539), .ZN(n8662) );
  NAND2_X1 U4877 ( .A1(n4450), .A2(n4449), .ZN(n9291) );
  OR2_X1 U4878 ( .A1(n8730), .A2(n4577), .ZN(n4574) );
  NAND2_X1 U4879 ( .A1(n6086), .A2(n6743), .ZN(n9398) );
  OR2_X1 U4880 ( .A1(n7999), .A2(n4572), .ZN(n4567) );
  AOI21_X1 U4881 ( .B1(n7916), .B2(n4331), .A(n4882), .ZN(n8010) );
  NAND2_X1 U4882 ( .A1(n5515), .A2(n5514), .ZN(n9348) );
  OAI21_X1 U4883 ( .B1(n7420), .B2(n4346), .A(n4622), .ZN(n4621) );
  INV_X1 U4884 ( .A(n7921), .ZN(n8249) );
  NAND2_X1 U4885 ( .A1(n6454), .A2(n6453), .ZN(n8038) );
  INV_X1 U4886 ( .A(n7536), .ZN(n4596) );
  NAND4_X1 U4887 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n9039)
         );
  NAND4_X1 U4888 ( .A1(n5259), .A2(n5258), .A3(n5257), .A4(n5256), .ZN(n9040)
         );
  CLKBUF_X1 U4889 ( .A(n5844), .Z(n9047) );
  NAND2_X1 U4890 ( .A1(n4443), .A2(n4440), .ZN(n5277) );
  AND2_X2 U4891 ( .A1(n9441), .A2(n6061), .ZN(n9542) );
  OAI21_X1 U4892 ( .B1(n6743), .B2(n4726), .A(n4725), .ZN(n9548) );
  NAND4_X2 U4893 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n5844)
         );
  NAND4_X1 U4894 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n6192)
         );
  NAND4_X1 U4895 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n5855)
         );
  INV_X2 U4896 ( .A(n7118), .ZN(n9863) );
  OAI211_X1 U4897 ( .C1(n6743), .C2(n9497), .A(n5145), .B(n5144), .ZN(n5611)
         );
  BUF_X2 U4898 ( .A(n5192), .Z(n6087) );
  INV_X2 U4899 ( .A(n5143), .ZN(n6182) );
  AND2_X1 U4900 ( .A1(n5120), .A2(n5119), .ZN(n5192) );
  AND2_X1 U4901 ( .A1(n5121), .A2(n8109), .ZN(n4910) );
  AND3_X1 U4902 ( .A1(n6355), .A2(n6354), .A3(n6353), .ZN(n7224) );
  NAND4_X1 U4903 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n8532)
         );
  NAND4_X2 U4904 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n9842)
         );
  AND4_X1 U4905 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n7147)
         );
  AND2_X1 U4906 ( .A1(n5834), .A2(n6313), .ZN(n5835) );
  INV_X2 U4907 ( .A(n8317), .ZN(n8307) );
  AND2_X1 U4908 ( .A1(n6356), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6342) );
  OR2_X2 U4909 ( .A1(n5106), .A2(n5105), .ZN(n6714) );
  NAND2_X1 U4910 ( .A1(n9445), .A2(n5118), .ZN(n8109) );
  BUF_X2 U4911 ( .A(n6356), .Z(n4297) );
  NAND2_X1 U4912 ( .A1(n5117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U4913 ( .A1(n5104), .A2(n5103), .ZN(n5105) );
  INV_X2 U4914 ( .A(n6661), .ZN(n6499) );
  AND2_X2 U4915 ( .A1(n6330), .A2(n6328), .ZN(n6346) );
  XNOR2_X1 U4916 ( .A(n5089), .B(n5088), .ZN(n5833) );
  XNOR2_X1 U4917 ( .A(n5636), .B(n5635), .ZN(n8117) );
  NAND2_X1 U4918 ( .A1(n5646), .A2(n5645), .ZN(n8172) );
  XNOR2_X1 U4919 ( .A(n6324), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U4920 ( .A1(n5087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U4921 ( .A(n5067), .B(n5066), .ZN(n5106) );
  INV_X1 U4922 ( .A(n7992), .ZN(n5103) );
  XNOR2_X1 U4923 ( .A(n5082), .B(n5081), .ZN(n7684) );
  OAI21_X1 U4924 ( .B1(n5073), .B2(n5065), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5067) );
  OR2_X1 U4925 ( .A1(n8894), .A2(n5694), .ZN(n6324) );
  OR2_X1 U4926 ( .A1(n5077), .A2(n5176), .ZN(n5078) );
  NAND2_X1 U4927 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  CLKBUF_X1 U4928 ( .A(n5060), .Z(n5069) );
  NAND2_X1 U4929 ( .A1(n5085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5412) );
  AND2_X1 U4930 ( .A1(n5079), .A2(n5081), .ZN(n5077) );
  AOI21_X1 U4931 ( .B1(n5059), .B2(P1_IR_REG_25__SCAN_IN), .A(n4426), .ZN(
        n4425) );
  NOR2_X1 U4932 ( .A1(n5083), .A2(n5062), .ZN(n5079) );
  XNOR2_X1 U4933 ( .A(n4944), .B(SI_2_), .ZN(n5142) );
  NAND2_X1 U4934 ( .A1(n5696), .A2(n5695), .ZN(n6727) );
  XNOR2_X1 U4935 ( .A(n4481), .B(n5710), .ZN(n7026) );
  NOR2_X1 U4936 ( .A1(n5666), .A2(n5630), .ZN(n5631) );
  AND2_X1 U4937 ( .A1(n4360), .A2(n6611), .ZN(n4895) );
  NOR2_X1 U4938 ( .A1(n5706), .A2(n4874), .ZN(n5663) );
  NAND3_X1 U4939 ( .A1(n5693), .A2(n4873), .A3(n4748), .ZN(n5706) );
  INV_X1 U4940 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5081) );
  INV_X1 U4941 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U4942 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4914) );
  INV_X1 U4943 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5114) );
  INV_X4 U4944 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4945 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6611) );
  NOR2_X1 U4946 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5064) );
  INV_X1 U4947 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5668) );
  NOR2_X1 U4948 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4605) );
  NOR2_X1 U4949 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4872) );
  INV_X1 U4950 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5710) );
  NOR2_X1 U4951 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4603) );
  NOR2_X1 U4952 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4604) );
  OAI21_X2 U4953 ( .B1(n7431), .B2(n4332), .A(n6621), .ZN(n7420) );
  NAND2_X2 U4954 ( .A1(n5139), .A2(n6722), .ZN(n5184) );
  NAND2_X1 U4955 ( .A1(n5061), .A2(n4919), .ZN(n5083) );
  NAND2_X1 U4956 ( .A1(n6034), .A2(n6031), .ZN(n4289) );
  INV_X1 U4957 ( .A(n5139), .ZN(n5128) );
  NAND2_X1 U4958 ( .A1(n5139), .A2(n6717), .ZN(n4292) );
  NAND2_X1 U4959 ( .A1(n5139), .A2(n6717), .ZN(n5143) );
  NAND4_X2 U4960 ( .A1(n4286), .A2(n5174), .A3(n4914), .A4(n4913), .ZN(n5243)
         );
  AOI21_X1 U4961 ( .B1(n5844), .B2(n5848), .A(n5849), .ZN(n5851) );
  OAI21_X2 U4962 ( .B1(n7090), .B2(n4713), .A(n4711), .ZN(n6099) );
  NAND2_X2 U4963 ( .A1(n4931), .A2(n5115), .ZN(n5605) );
  XNOR2_X1 U4964 ( .A(n4934), .B(n4933), .ZN(n9464) );
  AOI21_X2 U4965 ( .B1(n9297), .B2(n9298), .A(n6285), .ZN(n9280) );
  AND2_X1 U4966 ( .A1(n8902), .A2(n6328), .ZN(n4295) );
  INV_X1 U4967 ( .A(n4295), .ZN(n4296) );
  AND2_X4 U4968 ( .A1(n8902), .A2(n6328), .ZN(n6376) );
  NAND2_X1 U4969 ( .A1(n8262), .A2(n8265), .ZN(n8263) );
  NAND2_X1 U4970 ( .A1(n4679), .A2(n8275), .ZN(n4678) );
  NAND2_X1 U4971 ( .A1(n8272), .A2(n8729), .ZN(n4679) );
  INV_X1 U4972 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5627) );
  OAI21_X1 U4973 ( .B1(n4304), .B2(n4625), .A(n4328), .ZN(n4624) );
  INV_X1 U4974 ( .A(n6622), .ZN(n4625) );
  INV_X1 U4975 ( .A(n5659), .ZN(n5657) );
  NAND2_X1 U4976 ( .A1(n4723), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U4977 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  OR2_X1 U4978 ( .A1(n4724), .A2(n9401), .ZN(n4723) );
  AND2_X1 U4979 ( .A1(n9401), .A2(n6307), .ZN(n4722) );
  NAND2_X2 U4980 ( .A1(n5605), .A2(n9464), .ZN(n5139) );
  NAND2_X1 U4981 ( .A1(n9209), .A2(n4533), .ZN(n9128) );
  NOR2_X1 U4982 ( .A1(n9140), .A2(n4534), .ZN(n4533) );
  INV_X1 U4983 ( .A(n4535), .ZN(n4534) );
  AOI21_X1 U4984 ( .B1(n8204), .B2(n4334), .A(n4311), .ZN(n4677) );
  AND2_X1 U4985 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U4986 ( .A1(n7528), .A2(n6122), .ZN(n4706) );
  AND2_X1 U4987 ( .A1(n6125), .A2(n6124), .ZN(n4707) );
  NAND2_X1 U4988 ( .A1(n8263), .A2(n8326), .ZN(n8271) );
  NAND2_X1 U4989 ( .A1(n8174), .A2(n8326), .ZN(n4794) );
  NAND2_X1 U4990 ( .A1(n4795), .A2(n8310), .ZN(n4791) );
  NAND2_X1 U4991 ( .A1(n4678), .A2(n4342), .ZN(n4792) );
  OAI211_X1 U4992 ( .C1(n6147), .C2(n4904), .A(n6149), .B(n6146), .ZN(n6144)
         );
  NOR2_X1 U4993 ( .A1(n6217), .A2(n6307), .ZN(n4518) );
  NAND2_X1 U4994 ( .A1(n4444), .A2(n4445), .ZN(n4798) );
  NAND2_X1 U4995 ( .A1(n4383), .A2(n5006), .ZN(n4445) );
  NAND2_X1 U4996 ( .A1(n4985), .A2(n4984), .ZN(n4997) );
  INV_X1 U4997 ( .A(SI_14_), .ZN(n4984) );
  OR2_X1 U4998 ( .A1(n8305), .A2(n4675), .ZN(n8312) );
  NAND2_X1 U4999 ( .A1(n4676), .A2(n8304), .ZN(n4675) );
  AOI21_X1 U5000 ( .B1(n4672), .B2(n8619), .A(n4666), .ZN(n4665) );
  OR2_X1 U5001 ( .A1(n4667), .A2(n8329), .ZN(n4666) );
  NAND2_X1 U5002 ( .A1(n8330), .A2(n8310), .ZN(n4667) );
  AOI21_X1 U5003 ( .B1(n8203), .B2(n8226), .A(n4566), .ZN(n4565) );
  INV_X1 U5004 ( .A(n8348), .ZN(n4566) );
  OR2_X1 U5005 ( .A1(n6729), .A2(n6680), .ZN(n6699) );
  AND2_X1 U5006 ( .A1(n6669), .A2(n6754), .ZN(n7045) );
  OR2_X1 U5007 ( .A1(n8881), .A2(n8746), .ZN(n8178) );
  INV_X1 U5008 ( .A(n8255), .ZN(n4573) );
  OR2_X1 U5009 ( .A1(n8888), .A2(n8457), .ZN(n8267) );
  OR2_X1 U5010 ( .A1(n8099), .A2(n8748), .ZN(n8261) );
  OR2_X1 U5011 ( .A1(n8211), .A2(n8209), .ZN(n8208) );
  INV_X1 U5012 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U5013 ( .A1(n8916), .A2(n4411), .ZN(n4404) );
  AND2_X1 U5014 ( .A1(n4408), .A2(n4403), .ZN(n4402) );
  NAND2_X1 U5015 ( .A1(n8917), .A2(n4411), .ZN(n4403) );
  NOR2_X1 U5016 ( .A1(n8924), .A2(n4409), .ZN(n4408) );
  INV_X1 U5017 ( .A(n8965), .ZN(n4409) );
  NOR2_X1 U5018 ( .A1(n4831), .A2(n5900), .ZN(n4830) );
  OR2_X1 U5019 ( .A1(n4837), .A2(n4832), .ZN(n4831) );
  INV_X1 U5020 ( .A(n7127), .ZN(n4832) );
  NAND2_X1 U5021 ( .A1(n4840), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5022 ( .A1(n4836), .A2(n7166), .ZN(n4833) );
  INV_X1 U5023 ( .A(n7178), .ZN(n4839) );
  NAND2_X1 U5024 ( .A1(n7063), .A2(n5880), .ZN(n5887) );
  INV_X1 U5025 ( .A(n8109), .ZN(n5120) );
  INV_X1 U5026 ( .A(n5431), .ZN(n4773) );
  NOR2_X1 U5027 ( .A1(n9317), .A2(n9380), .ZN(n9283) );
  NOR2_X1 U5028 ( .A1(n8946), .A2(n7835), .ZN(n4543) );
  NAND2_X1 U5029 ( .A1(n9580), .A2(n4462), .ZN(n4785) );
  NAND2_X1 U5030 ( .A1(n7323), .A2(n9044), .ZN(n6263) );
  INV_X1 U5031 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5032 ( .B1(n4764), .B2(n4763), .A(n5523), .ZN(n4762) );
  NAND2_X1 U5033 ( .A1(n5535), .A2(n5536), .ZN(n5548) );
  INV_X1 U5034 ( .A(n5060), .ZN(n4926) );
  AND2_X1 U5035 ( .A1(n5039), .A2(n5038), .ZN(n5512) );
  OAI21_X1 U5036 ( .B1(n4798), .B2(n4797), .A(n4796), .ZN(n5448) );
  AOI21_X1 U5037 ( .B1(n4800), .B2(n4804), .A(n4805), .ZN(n4796) );
  NOR2_X1 U5038 ( .A1(n4800), .A2(n4807), .ZN(n4797) );
  OAI21_X1 U5039 ( .B1(n5017), .B2(n4806), .A(n4382), .ZN(n4805) );
  INV_X1 U5040 ( .A(n4798), .ZN(n5411) );
  NOR2_X1 U5041 ( .A1(n4822), .A2(n4442), .ZN(n4441) );
  NOR2_X1 U5042 ( .A1(n5291), .A2(n4828), .ZN(n4827) );
  INV_X1 U5043 ( .A(n4979), .ZN(n4828) );
  NAND2_X1 U5044 ( .A1(n4589), .A2(n4812), .ZN(n5263) );
  AOI21_X1 U5045 ( .B1(n4813), .B2(n4815), .A(n4350), .ZN(n4812) );
  NAND2_X1 U5046 ( .A1(n4964), .A2(SI_7_), .ZN(n4968) );
  AND2_X1 U5047 ( .A1(n6661), .A2(n6722), .ZN(n4608) );
  NOR2_X1 U5048 ( .A1(n8443), .A2(n4878), .ZN(n4877) );
  INV_X1 U5049 ( .A(n8123), .ZN(n4878) );
  NAND2_X1 U5050 ( .A1(n5648), .A2(n5647), .ZN(n6698) );
  NAND2_X1 U5051 ( .A1(n8628), .A2(n6645), .ZN(n8615) );
  NAND2_X1 U5052 ( .A1(n6530), .A2(n8279), .ZN(n8672) );
  NAND2_X1 U5053 ( .A1(n8742), .A2(n6633), .ZN(n8733) );
  INV_X1 U5054 ( .A(n4624), .ZN(n4622) );
  INV_X2 U5055 ( .A(n8316), .ZN(n6500) );
  NAND2_X2 U5056 ( .A1(n6682), .A2(n6651), .ZN(n9844) );
  NAND2_X1 U5057 ( .A1(n5633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5643) );
  INV_X1 U5058 ( .A(n6087), .ZN(n5557) );
  OR2_X1 U5059 ( .A1(n5315), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5350) );
  NOR2_X1 U5060 ( .A1(n9401), .A2(n9128), .ZN(n9131) );
  AOI21_X1 U5061 ( .B1(n4306), .B2(n4453), .A(n4373), .ZN(n4449) );
  NOR2_X1 U5062 ( .A1(n9620), .A2(n5833), .ZN(n6061) );
  AND2_X1 U5063 ( .A1(n5072), .A2(n9443), .ZN(n7311) );
  OR2_X1 U5064 ( .A1(n6313), .A2(n5833), .ZN(n9513) );
  NAND2_X1 U5065 ( .A1(n7880), .A2(n7723), .ZN(n6842) );
  NAND2_X1 U5066 ( .A1(n5600), .A2(n5599), .ZN(n9541) );
  OR2_X1 U5067 ( .A1(n5075), .A2(n5074), .ZN(n5076) );
  NAND2_X1 U5068 ( .A1(n5330), .A2(n4993), .ZN(n5333) );
  AND2_X1 U5069 ( .A1(n8157), .A2(n8618), .ZN(n8158) );
  INV_X1 U5070 ( .A(n7559), .ZN(n8382) );
  OR2_X1 U5071 ( .A1(n6852), .A2(n6847), .ZN(n9817) );
  OR2_X1 U5072 ( .A1(n4504), .A2(n4301), .ZN(n4500) );
  NAND2_X1 U5073 ( .A1(n4715), .A2(n4501), .ZN(n4498) );
  OAI21_X1 U5074 ( .B1(n5143), .B2(n8112), .A(n5057), .ZN(n9140) );
  NAND2_X1 U5075 ( .A1(n8185), .A2(n8184), .ZN(n8188) );
  NAND2_X1 U5076 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5077 ( .A1(n8254), .A2(n4340), .ZN(n4662) );
  NOR2_X1 U5078 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  INV_X1 U5079 ( .A(n8359), .ZN(n4659) );
  INV_X1 U5080 ( .A(n4660), .ZN(n4657) );
  AOI21_X1 U5081 ( .B1(n4703), .B2(n4704), .A(n4584), .ZN(n4702) );
  NAND2_X1 U5082 ( .A1(n4487), .A2(n6117), .ZN(n4486) );
  OAI21_X1 U5083 ( .B1(n6116), .B2(n6272), .A(n6276), .ZN(n4487) );
  NAND2_X1 U5084 ( .A1(n6119), .A2(n6118), .ZN(n4485) );
  INV_X1 U5085 ( .A(n6140), .ZN(n6119) );
  NAND2_X1 U5086 ( .A1(n4793), .A2(n8279), .ZN(n4787) );
  AND2_X1 U5087 ( .A1(n8277), .A2(n8326), .ZN(n4793) );
  OR2_X1 U5088 ( .A1(n6225), .A2(n6096), .ZN(n4521) );
  AOI21_X1 U5089 ( .B1(n4352), .B2(n4511), .A(n4518), .ZN(n4510) );
  OAI21_X1 U5090 ( .B1(n6173), .B2(n6176), .A(n6172), .ZN(n4496) );
  INV_X1 U5091 ( .A(n4810), .ZN(n4803) );
  NAND2_X1 U5092 ( .A1(n4680), .A2(n8298), .ZN(n8301) );
  OAI21_X1 U5093 ( .B1(n8295), .B2(n8294), .A(n4683), .ZN(n4682) );
  OR2_X1 U5094 ( .A1(n6691), .A2(n8600), .ZN(n8306) );
  INV_X1 U5095 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4896) );
  NOR2_X1 U5096 ( .A1(n5900), .A2(n4837), .ZN(n4836) );
  AND2_X1 U5097 ( .A1(n8946), .A2(n5396), .ZN(n6280) );
  NOR2_X1 U5098 ( .A1(n5212), .A2(n4592), .ZN(n4591) );
  INV_X1 U5099 ( .A(n4958), .ZN(n4592) );
  NAND2_X1 U5100 ( .A1(n8312), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U5101 ( .A1(n4676), .A2(n4674), .ZN(n4673) );
  INV_X1 U5102 ( .A(n8311), .ZN(n4674) );
  NAND2_X1 U5103 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  NOR2_X1 U5104 ( .A1(n8332), .A2(n8310), .ZN(n4671) );
  NAND2_X1 U5105 ( .A1(n4634), .A2(n4633), .ZN(n9675) );
  NOR2_X1 U5106 ( .A1(n4737), .A2(n6734), .ZN(n4738) );
  OAI21_X1 U5107 ( .B1(n5708), .B2(n4737), .A(n4735), .ZN(n9728) );
  AND2_X1 U5108 ( .A1(n4736), .A2(n6734), .ZN(n4735) );
  NAND2_X1 U5109 ( .A1(n4480), .A2(n5709), .ZN(n4736) );
  INV_X1 U5110 ( .A(n7008), .ZN(n4480) );
  NAND2_X1 U5111 ( .A1(n9732), .A2(n4471), .ZN(n5726) );
  NOR2_X1 U5112 ( .A1(n7195), .A2(n4472), .ZN(n4471) );
  INV_X1 U5113 ( .A(n5721), .ZN(n4472) );
  NAND2_X1 U5114 ( .A1(n5726), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5115 ( .A1(n4476), .A2(n4314), .ZN(n4740) );
  AND2_X1 U5116 ( .A1(n6534), .A2(n6533), .ZN(n6543) );
  NOR2_X1 U5117 ( .A1(n6525), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6534) );
  NOR2_X1 U5118 ( .A1(n6475), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U5119 ( .B1(n8654), .B2(n4546), .A(n4545), .ZN(n8333) );
  NAND2_X1 U5120 ( .A1(n4324), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5121 ( .A1(n4548), .A2(n4324), .ZN(n4545) );
  INV_X1 U5122 ( .A(n4553), .ZN(n4547) );
  OR2_X1 U5123 ( .A1(n8826), .A2(n8599), .ZN(n8302) );
  OR2_X1 U5124 ( .A1(n8837), .A2(n8468), .ZN(n8296) );
  NOR2_X1 U5125 ( .A1(n4620), .A2(n4616), .ZN(n4615) );
  OR2_X1 U5126 ( .A1(n8848), .A2(n8487), .ZN(n8338) );
  OR2_X1 U5127 ( .A1(n8864), .A2(n8693), .ZN(n8277) );
  CLKBUF_X1 U5128 ( .A(n5663), .Z(n5664) );
  OR2_X1 U5129 ( .A1(n5717), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5723) );
  OR2_X1 U5130 ( .A1(n5960), .A2(n7944), .ZN(n4845) );
  AOI21_X1 U5131 ( .B1(n4303), .B2(n4423), .A(n4355), .ZN(n4420) );
  OR2_X1 U5132 ( .A1(n9401), .A2(n6307), .ZN(n6186) );
  NAND2_X1 U5133 ( .A1(n4488), .A2(n6178), .ZN(n4724) );
  NAND2_X1 U5134 ( .A1(n4491), .A2(n6096), .ZN(n4490) );
  INV_X1 U5135 ( .A(n9401), .ZN(n6187) );
  NOR2_X1 U5136 ( .A1(n9178), .A2(n4538), .ZN(n4537) );
  INV_X1 U5137 ( .A(n9413), .ZN(n4538) );
  INV_X1 U5138 ( .A(n6236), .ZN(n6171) );
  OR2_X1 U5139 ( .A1(n9354), .A2(n5593), .ZN(n6221) );
  OR2_X1 U5140 ( .A1(n9427), .A2(n5460), .ZN(n6155) );
  NOR2_X1 U5141 ( .A1(n9377), .A2(n9427), .ZN(n4528) );
  OR2_X1 U5142 ( .A1(n9437), .A2(n9031), .ZN(n6146) );
  OR2_X1 U5143 ( .A1(n8946), .A2(n5396), .ZN(n6135) );
  NOR2_X1 U5144 ( .A1(n7643), .A2(n7644), .ZN(n6117) );
  NAND2_X1 U5145 ( .A1(n7467), .A2(n7466), .ZN(n4585) );
  NAND2_X1 U5146 ( .A1(n4596), .A2(n9037), .ZN(n6125) );
  NOR2_X1 U5147 ( .A1(n4755), .A2(n4752), .ZN(n4751) );
  INV_X1 U5148 ( .A(n7510), .ZN(n4755) );
  INV_X1 U5149 ( .A(n5261), .ZN(n4754) );
  AOI21_X1 U5150 ( .B1(n4714), .B2(n6261), .A(n4712), .ZN(n4711) );
  NAND2_X1 U5151 ( .A1(n4347), .A2(n4766), .ZN(n4763) );
  NAND2_X1 U5152 ( .A1(n6080), .A2(n6079), .ZN(n6181) );
  OR2_X1 U5153 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NAND2_X1 U5154 ( .A1(n5045), .A2(n5044), .ZN(n5535) );
  NAND2_X1 U5155 ( .A1(n4429), .A2(n4427), .ZN(n5045) );
  AOI21_X1 U5156 ( .B1(n4430), .B2(n4433), .A(n4428), .ZN(n4427) );
  INV_X1 U5157 ( .A(n5446), .ZN(n5019) );
  INV_X1 U5158 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4915) );
  OR2_X1 U5159 ( .A1(n4988), .A2(n4995), .ZN(n4989) );
  OAI21_X1 U5160 ( .B1(n4443), .B2(n4821), .A(n4438), .ZN(n4990) );
  AND2_X1 U5161 ( .A1(n4968), .A2(n4967), .ZN(n5222) );
  AND2_X1 U5162 ( .A1(n7362), .A2(n7360), .ZN(n4881) );
  INV_X1 U5163 ( .A(n8666), .ZN(n8436) );
  NOR2_X1 U5164 ( .A1(n4894), .A2(n8149), .ZN(n4893) );
  INV_X1 U5165 ( .A(n8148), .ZN(n4894) );
  XNOR2_X1 U5166 ( .A(n6995), .B(n7112), .ZN(n7029) );
  NAND2_X1 U5167 ( .A1(n4606), .A2(n4608), .ZN(n6336) );
  INV_X1 U5168 ( .A(n6726), .ZN(n4606) );
  NAND2_X1 U5169 ( .A1(n8007), .A2(n4884), .ZN(n4883) );
  INV_X1 U5170 ( .A(n7983), .ZN(n4884) );
  NOR2_X1 U5171 ( .A1(n7919), .A2(n4886), .ZN(n4885) );
  INV_X1 U5172 ( .A(n7915), .ZN(n4886) );
  AND2_X1 U5173 ( .A1(n8323), .A2(n8322), .ZN(n8572) );
  AND3_X1 U5174 ( .A1(n6529), .A2(n6528), .A3(n6527), .ZN(n8143) );
  AND4_X1 U5175 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n8457)
         );
  XNOR2_X1 U5176 ( .A(n7026), .B(n5707), .ZN(n7008) );
  AOI21_X1 U5177 ( .B1(n7026), .B2(n5789), .A(n7003), .ZN(n9716) );
  NAND2_X1 U5178 ( .A1(n9765), .A2(n5760), .ZN(n5761) );
  OAI21_X1 U5179 ( .B1(n7582), .B2(n4473), .A(n4474), .ZN(n4476) );
  AOI21_X1 U5180 ( .B1(n5732), .B2(n4475), .A(n7731), .ZN(n4474) );
  INV_X1 U5181 ( .A(n5732), .ZN(n4473) );
  NAND2_X1 U5182 ( .A1(n7582), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U5183 ( .B1(n7580), .B2(n4640), .A(n4638), .ZN(n4642) );
  INV_X1 U5184 ( .A(n5762), .ZN(n4640) );
  AOI21_X1 U5185 ( .B1(n5762), .B2(n4639), .A(n7728), .ZN(n4638) );
  XNOR2_X1 U5186 ( .A(n4740), .B(n8073), .ZN(n8069) );
  OR2_X1 U5187 ( .A1(n8053), .A2(n5737), .ZN(n4734) );
  AND2_X1 U5188 ( .A1(n4734), .A2(n4733), .ZN(n9774) );
  INV_X1 U5189 ( .A(n9775), .ZN(n4733) );
  NOR2_X1 U5190 ( .A1(n5742), .A2(n9811), .ZN(n8565) );
  OR2_X1 U5191 ( .A1(n6551), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U5192 ( .A1(n4311), .A2(n4564), .ZN(n4562) );
  INV_X1 U5193 ( .A(n8226), .ZN(n4564) );
  NAND2_X1 U5194 ( .A1(n4563), .A2(n4565), .ZN(n7430) );
  NAND2_X1 U5195 ( .A1(n7294), .A2(n8226), .ZN(n4563) );
  AND2_X1 U5196 ( .A1(n8231), .A2(n7418), .ZN(n8348) );
  INV_X1 U5197 ( .A(n8648), .ZN(n8618) );
  OR2_X1 U5198 ( .A1(n8832), .A2(n8618), .ZN(n8608) );
  AND2_X1 U5199 ( .A1(n4333), .A2(n6642), .ZN(n4650) );
  AND2_X1 U5200 ( .A1(n8296), .A2(n8297), .ZN(n8638) );
  OR2_X1 U5201 ( .A1(n8843), .A2(n8436), .ZN(n8335) );
  NAND2_X1 U5202 ( .A1(n8673), .A2(n8675), .ZN(n4617) );
  AND2_X1 U5203 ( .A1(n6639), .A2(n6638), .ZN(n4651) );
  AOI21_X1 U5204 ( .B1(n4578), .B2(n4576), .A(n8274), .ZN(n4575) );
  OR2_X1 U5205 ( .A1(n8875), .A2(n8413), .ZN(n8709) );
  AND2_X1 U5206 ( .A1(n6632), .A2(n6630), .ZN(n4649) );
  AOI21_X1 U5207 ( .B1(n4571), .B2(n8256), .A(n4569), .ZN(n4568) );
  INV_X1 U5208 ( .A(n8264), .ZN(n4569) );
  AND2_X1 U5209 ( .A1(n8267), .A2(n8265), .ZN(n8757) );
  INV_X1 U5210 ( .A(n8073), .ZN(n6424) );
  INV_X1 U5211 ( .A(n4559), .ZN(n4558) );
  OAI21_X1 U5212 ( .B1(n6411), .B2(n4299), .A(n8229), .ZN(n4559) );
  OR2_X1 U5213 ( .A1(n9889), .A2(n7820), .ZN(n8225) );
  AND2_X1 U5214 ( .A1(n4325), .A2(n4631), .ZN(n4626) );
  NOR2_X1 U5215 ( .A1(n4628), .A2(n4339), .ZN(n4627) );
  INV_X1 U5216 ( .A(n4321), .ZN(n4628) );
  INV_X1 U5217 ( .A(n8745), .ZN(n9841) );
  OR2_X1 U5218 ( .A1(n6687), .A2(n8387), .ZN(n9885) );
  NOR2_X1 U5219 ( .A1(n6941), .A2(n6946), .ZN(n6935) );
  NOR2_X1 U5220 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4684) );
  NAND2_X1 U5221 ( .A1(n5643), .A2(n5634), .ZN(n5645) );
  XNOR2_X1 U5222 ( .A(n5654), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8342) );
  INV_X1 U5223 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4873) );
  INV_X1 U5224 ( .A(n5955), .ZN(n4844) );
  NAND2_X1 U5225 ( .A1(n5956), .A2(n5955), .ZN(n4847) );
  INV_X1 U5226 ( .A(n4407), .ZN(n4406) );
  NAND2_X1 U5227 ( .A1(n4404), .A2(n4402), .ZN(n4405) );
  OAI21_X1 U5228 ( .B1(n8924), .B2(n4410), .A(n6004), .ZN(n4407) );
  NAND2_X1 U5229 ( .A1(n5983), .A2(n5984), .ZN(n4863) );
  NAND2_X1 U5230 ( .A1(n7399), .A2(n5915), .ZN(n7744) );
  AOI21_X1 U5231 ( .B1(n4856), .B2(n4302), .A(n4379), .ZN(n4855) );
  NOR2_X1 U5232 ( .A1(n4857), .A2(n8957), .ZN(n4856) );
  NOR2_X1 U5233 ( .A1(n4302), .A2(n8910), .ZN(n4857) );
  INV_X1 U5234 ( .A(n5888), .ZN(n5889) );
  INV_X1 U5235 ( .A(n5887), .ZN(n4401) );
  NAND2_X1 U5236 ( .A1(n9006), .A2(n4416), .ZN(n4415) );
  NOR2_X1 U5237 ( .A1(n4417), .A2(n4418), .ZN(n4416) );
  INV_X1 U5238 ( .A(n9005), .ZN(n4418) );
  NAND2_X1 U5239 ( .A1(n4413), .A2(n8941), .ZN(n4412) );
  INV_X1 U5240 ( .A(n5967), .ZN(n4413) );
  AOI22_X1 U5241 ( .A1(n9580), .A2(n6052), .B1(n5848), .B2(n9044), .ZN(n7059)
         );
  XNOR2_X1 U5242 ( .A(n5875), .B(n6050), .ZN(n7060) );
  NAND2_X1 U5243 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U5244 ( .A1(n4290), .A2(n9580), .ZN(n5873) );
  NAND3_X1 U5245 ( .A1(n5838), .A2(n5837), .A3(n5839), .ZN(n6865) );
  INV_X1 U5246 ( .A(n5980), .ZN(n4862) );
  NAND2_X1 U5247 ( .A1(n7124), .A2(n7127), .ZN(n7164) );
  NOR2_X1 U5248 ( .A1(n4503), .A2(n4502), .ZN(n6312) );
  NAND2_X1 U5249 ( .A1(n4719), .A2(n6308), .ZN(n4503) );
  AND4_X1 U5250 ( .A1(n5211), .A2(n5210), .A3(n4484), .A4(n4483), .ZN(n5219)
         );
  NAND2_X1 U5251 ( .A1(n6088), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5252 ( .A1(n6087), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U5253 ( .A1(n4454), .A2(n4366), .ZN(n9158) );
  NOR2_X1 U5254 ( .A1(n9173), .A2(n4456), .ZN(n4455) );
  NAND2_X1 U5255 ( .A1(n9209), .A2(n9413), .ZN(n9192) );
  NOR2_X1 U5256 ( .A1(n5511), .A2(n4765), .ZN(n4764) );
  INV_X1 U5257 ( .A(n5492), .ZN(n4765) );
  NAND2_X1 U5258 ( .A1(n4767), .A2(n5593), .ZN(n4766) );
  OR2_X1 U5259 ( .A1(n6008), .A2(n9028), .ZN(n4461) );
  OR2_X1 U5260 ( .A1(n9377), .A2(n8919), .ZN(n6154) );
  INV_X1 U5261 ( .A(n4770), .ZN(n4769) );
  OAI21_X1 U5262 ( .B1(n4367), .B2(n4771), .A(n4776), .ZN(n4770) );
  OR2_X1 U5263 ( .A1(n9377), .A2(n8926), .ZN(n4776) );
  AND2_X1 U5264 ( .A1(n6155), .A2(n6159), .ZN(n9261) );
  NAND2_X1 U5265 ( .A1(n9280), .A2(n9279), .ZN(n9278) );
  NOR2_X1 U5266 ( .A1(n4544), .A2(n4540), .ZN(n4539) );
  INV_X1 U5267 ( .A(n9437), .ZN(n4544) );
  INV_X1 U5268 ( .A(n4541), .ZN(n4540) );
  NAND2_X1 U5269 ( .A1(n4319), .A2(n5397), .ZN(n7937) );
  AND2_X1 U5270 ( .A1(n4458), .A2(n5379), .ZN(n4457) );
  OR2_X1 U5271 ( .A1(n4459), .A2(n5360), .ZN(n4458) );
  OR2_X1 U5272 ( .A1(n8120), .A2(n5143), .ZN(n5337) );
  NAND2_X1 U5273 ( .A1(n6126), .A2(n6125), .ZN(n7525) );
  NOR2_X1 U5274 ( .A1(n4523), .A2(n7450), .ZN(n9515) );
  INV_X1 U5275 ( .A(n4785), .ZN(n5581) );
  INV_X1 U5276 ( .A(n5578), .ZN(n4700) );
  OR2_X1 U5277 ( .A1(n9549), .A2(n9548), .ZN(n9552) );
  INV_X1 U5278 ( .A(n9541), .ZN(n9506) );
  AND2_X1 U5279 ( .A1(n6043), .A2(n5107), .ZN(n7312) );
  INV_X1 U5280 ( .A(n9548), .ZN(n6841) );
  NAND2_X1 U5281 ( .A1(n5071), .A2(n5104), .ZN(n9442) );
  XNOR2_X1 U5282 ( .A(n6181), .B(n6180), .ZN(n8898) );
  AND2_X1 U5283 ( .A1(n4871), .A2(n4925), .ZN(n4870) );
  AND2_X1 U5284 ( .A1(n4928), .A2(n4933), .ZN(n4871) );
  XNOR2_X1 U5285 ( .A(n5535), .B(n5536), .ZN(n8103) );
  XNOR2_X1 U5286 ( .A(n5524), .B(n5525), .ZN(n8084) );
  OAI21_X1 U5287 ( .B1(n5476), .B2(n4433), .A(n4430), .ZN(n5524) );
  AND2_X1 U5288 ( .A1(n4436), .A2(n5495), .ZN(n5513) );
  NAND2_X1 U5289 ( .A1(n5476), .A2(n5035), .ZN(n4436) );
  XNOR2_X1 U5290 ( .A(n5498), .B(n5497), .ZN(n7979) );
  INV_X1 U5291 ( .A(n4799), .ZN(n5434) );
  NAND2_X1 U5292 ( .A1(n4447), .A2(n4829), .ZN(n5399) );
  XNOR2_X1 U5293 ( .A(n5383), .B(n5382), .ZN(n7151) );
  NAND2_X1 U5294 ( .A1(n4443), .A2(n4441), .ZN(n4437) );
  NOR2_X1 U5295 ( .A1(n5308), .A2(n4826), .ZN(n4823) );
  INV_X1 U5296 ( .A(n4442), .ZN(n4440) );
  NAND2_X1 U5297 ( .A1(n4952), .A2(n4951), .ZN(n5182) );
  AND2_X1 U5298 ( .A1(n5179), .A2(n5178), .ZN(n5216) );
  XNOR2_X1 U5299 ( .A(n4941), .B(SI_1_), .ZN(n5127) );
  NAND2_X1 U5300 ( .A1(n5137), .A2(n4939), .ZN(n5126) );
  NAND2_X1 U5301 ( .A1(n8133), .A2(n8132), .ZN(n8410) );
  OR2_X1 U5302 ( .A1(n8159), .A2(n8599), .ZN(n8160) );
  AND4_X1 U5303 ( .A1(n6432), .A2(n6431), .A3(n6430), .A4(n6429), .ZN(n8209)
         );
  AND4_X1 U5304 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n8748)
         );
  AND2_X1 U5305 ( .A1(n6442), .A2(n6441), .ZN(n7921) );
  AND4_X1 U5306 ( .A1(n6487), .A2(n6486), .A3(n6485), .A4(n6484), .ZN(n8746)
         );
  INV_X1 U5307 ( .A(n7879), .ZN(n8387) );
  INV_X1 U5308 ( .A(n8143), .ZN(n8703) );
  NAND2_X1 U5309 ( .A1(n7580), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7579) );
  OR2_X1 U5310 ( .A1(P2_U3150), .A2(n5827), .ZN(n9737) );
  NOR2_X1 U5311 ( .A1(n8565), .A2(n8564), .ZN(n8563) );
  NAND2_X1 U5312 ( .A1(n8566), .A2(n8567), .ZN(n4745) );
  INV_X1 U5313 ( .A(n4397), .ZN(n4396) );
  NOR2_X1 U5314 ( .A1(n4654), .A2(n9817), .ZN(n4468) );
  XNOR2_X1 U5315 ( .A(n5776), .B(n5775), .ZN(n4654) );
  NAND2_X1 U5316 ( .A1(n6522), .A2(n6521), .ZN(n8792) );
  AND2_X1 U5317 ( .A1(n6434), .A2(n6433), .ZN(n7958) );
  NAND2_X1 U5318 ( .A1(n7042), .A2(n6614), .ZN(n9832) );
  XNOR2_X1 U5319 ( .A(n5669), .B(n5668), .ZN(n7559) );
  NOR2_X1 U5320 ( .A1(n4869), .A2(n8988), .ZN(n4867) );
  AND2_X1 U5321 ( .A1(n8990), .A2(n6038), .ZN(n6706) );
  NAND2_X1 U5322 ( .A1(n5318), .A2(n5317), .ZN(n7663) );
  OR2_X1 U5323 ( .A1(n6919), .A2(n5143), .ZN(n5318) );
  NAND2_X1 U5324 ( .A1(n4851), .A2(n4849), .ZN(n8990) );
  NOR2_X1 U5325 ( .A1(n4853), .A2(n4850), .ZN(n4849) );
  INV_X1 U5326 ( .A(n8991), .ZN(n4850) );
  NOR2_X1 U5327 ( .A1(n6060), .A2(n6047), .ZN(n9007) );
  NAND2_X1 U5328 ( .A1(n5490), .A2(n5489), .ZN(n9027) );
  AND2_X1 U5329 ( .A1(n4695), .A2(n4694), .ZN(n6774) );
  NAND2_X1 U5330 ( .A1(n6813), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4694) );
  OAI21_X1 U5331 ( .B1(n9117), .B2(n9486), .A(n4693), .ZN(n4692) );
  AOI21_X1 U5332 ( .B1(n9118), .B2(n9492), .A(n9478), .ZN(n4693) );
  OAI21_X1 U5333 ( .B1(n9122), .B2(n4782), .A(n9121), .ZN(n4691) );
  OR2_X1 U5334 ( .A1(n9131), .A2(n9130), .ZN(n9331) );
  AND2_X1 U5335 ( .A1(n9154), .A2(n9153), .ZN(n9335) );
  NAND2_X1 U5336 ( .A1(n5534), .A2(n5533), .ZN(n9170) );
  NAND2_X1 U5337 ( .A1(n5202), .A2(n5201), .ZN(n7456) );
  NAND2_X1 U5338 ( .A1(n9404), .A2(n9428), .ZN(n4600) );
  NAND2_X1 U5339 ( .A1(n4601), .A2(n9335), .ZN(n9403) );
  INV_X1 U5340 ( .A(n4602), .ZN(n4601) );
  OAI21_X1 U5341 ( .B1(n9336), .B2(n9583), .A(n9334), .ZN(n4602) );
  AOI211_X1 U5342 ( .C1(n9339), .C2(n9635), .A(n9338), .B(n9337), .ZN(n9406)
         );
  NAND2_X1 U5343 ( .A1(n5056), .A2(n6080), .ZN(n8112) );
  NAND2_X1 U5344 ( .A1(n4657), .A2(n4344), .ZN(n4656) );
  AOI21_X1 U5345 ( .B1(n4705), .B2(n5586), .A(n4351), .ZN(n4703) );
  INV_X1 U5346 ( .A(n4705), .ZN(n4704) );
  NAND2_X1 U5347 ( .A1(n6110), .A2(n6109), .ZN(n6120) );
  AOI21_X1 U5348 ( .B1(n4486), .B2(n4307), .A(n4485), .ZN(n6139) );
  OAI21_X1 U5349 ( .B1(n4520), .B2(n4515), .A(n9248), .ZN(n4514) );
  INV_X1 U5350 ( .A(n4519), .ZN(n4515) );
  NAND2_X1 U5351 ( .A1(n6230), .A2(n6096), .ZN(n4520) );
  NAND2_X1 U5352 ( .A1(n4788), .A2(n4787), .ZN(n4789) );
  NOR2_X1 U5353 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  INV_X1 U5354 ( .A(n4521), .ZN(n4513) );
  INV_X1 U5355 ( .A(n4514), .ZN(n4511) );
  AOI21_X1 U5356 ( .B1(n4521), .B2(n6156), .A(n4517), .ZN(n4516) );
  AND2_X1 U5357 ( .A1(n6161), .A2(n6160), .ZN(n6217) );
  NOR2_X1 U5358 ( .A1(n8289), .A2(n8326), .ZN(n4683) );
  AOI21_X1 U5359 ( .B1(n4731), .B2(n4730), .A(n6169), .ZN(n6177) );
  NOR2_X1 U5360 ( .A1(n9220), .A2(n6165), .ZN(n4730) );
  INV_X1 U5361 ( .A(n6166), .ZN(n4731) );
  INV_X1 U5362 ( .A(n4829), .ZN(n4446) );
  NAND2_X1 U5363 ( .A1(n4448), .A2(n4968), .ZN(n4814) );
  INV_X1 U5364 ( .A(n5241), .ZN(n4448) );
  AOI21_X1 U5365 ( .B1(n5817), .B2(n9810), .A(n5816), .ZN(n5819) );
  INV_X1 U5366 ( .A(n7944), .ZN(n4846) );
  OR2_X1 U5367 ( .A1(n7657), .A2(n4423), .ZN(n4422) );
  INV_X1 U5368 ( .A(n5946), .ZN(n4423) );
  INV_X1 U5369 ( .A(n7177), .ZN(n4840) );
  OAI21_X1 U5370 ( .B1(n4492), .B2(n6242), .A(n9149), .ZN(n4491) );
  AOI21_X1 U5371 ( .B1(n4729), .B2(n4728), .A(n6240), .ZN(n4492) );
  NOR2_X1 U5372 ( .A1(n6176), .A2(n6236), .ZN(n4728) );
  NAND2_X1 U5373 ( .A1(n6177), .A2(n6224), .ZN(n4729) );
  NAND2_X1 U5374 ( .A1(n4495), .A2(n4494), .ZN(n4493) );
  NOR2_X1 U5375 ( .A1(n6174), .A2(n6096), .ZN(n4494) );
  NAND2_X1 U5376 ( .A1(n4496), .A2(n6175), .ZN(n4495) );
  INV_X1 U5377 ( .A(n6188), .ZN(n4721) );
  NOR2_X1 U5378 ( .A1(n6008), .A2(n4527), .ZN(n4526) );
  INV_X1 U5379 ( .A(n4528), .ZN(n4527) );
  NOR2_X1 U5380 ( .A1(n5951), .A2(n4530), .ZN(n4529) );
  INV_X1 U5381 ( .A(n4531), .ZN(n4530) );
  INV_X1 U5382 ( .A(n5525), .ZN(n4428) );
  NOR2_X1 U5383 ( .A1(n5034), .A2(n4435), .ZN(n4434) );
  INV_X1 U5384 ( .A(n5512), .ZN(n4435) );
  OR2_X1 U5385 ( .A1(n5418), .A2(SI_20_), .ZN(n5017) );
  NAND2_X1 U5386 ( .A1(n5011), .A2(n5010), .ZN(n4806) );
  NOR2_X1 U5387 ( .A1(n5017), .A2(n4811), .ZN(n4807) );
  INV_X1 U5388 ( .A(n4801), .ZN(n4800) );
  OAI21_X1 U5389 ( .B1(n4808), .B2(n4802), .A(n5016), .ZN(n4801) );
  NAND2_X1 U5390 ( .A1(n4803), .A2(SI_20_), .ZN(n4802) );
  OR2_X1 U5391 ( .A1(n4808), .A2(n10036), .ZN(n4804) );
  NAND2_X1 U5392 ( .A1(n5013), .A2(n5012), .ZN(n5018) );
  INV_X1 U5393 ( .A(SI_19_), .ZN(n5012) );
  INV_X1 U5394 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5007) );
  INV_X1 U5395 ( .A(SI_17_), .ZN(n5002) );
  INV_X1 U5396 ( .A(n4439), .ZN(n4438) );
  OAI21_X1 U5397 ( .B1(n4821), .B2(n4441), .A(n4986), .ZN(n4439) );
  INV_X1 U5398 ( .A(n4823), .ZN(n4822) );
  NOR2_X1 U5399 ( .A1(n4814), .A2(n4588), .ZN(n4587) );
  INV_X1 U5400 ( .A(n4963), .ZN(n4588) );
  INV_X1 U5401 ( .A(n4814), .ZN(n4815) );
  INV_X1 U5402 ( .A(n5222), .ZN(n4813) );
  INV_X1 U5403 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4912) );
  INV_X1 U5404 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4911) );
  OR2_X1 U5405 ( .A1(n6987), .A2(n6986), .ZN(n6990) );
  NAND2_X1 U5406 ( .A1(n9675), .A2(n5749), .ZN(n9693) );
  NAND2_X1 U5407 ( .A1(n5720), .A2(n9727), .ZN(n9732) );
  AOI21_X1 U5408 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6918), .A(n8016), .ZN(
        n5766) );
  AOI21_X1 U5409 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6918), .A(n8022), .ZN(
        n5736) );
  NOR2_X1 U5410 ( .A1(n9774), .A2(n4732), .ZN(n5739) );
  AND2_X1 U5411 ( .A1(n9790), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4732) );
  AOI21_X1 U5412 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9806), .A(n9791), .ZN(
        n5741) );
  NOR2_X1 U5413 ( .A1(n5819), .A2(n5818), .ZN(n8554) );
  NOR2_X1 U5414 ( .A1(n6443), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6456) );
  AND2_X1 U5415 ( .A1(n6405), .A2(n6404), .ZN(n6417) );
  NAND2_X1 U5416 ( .A1(n8216), .A2(n8199), .ZN(n8343) );
  NOR2_X1 U5417 ( .A1(n8335), .A2(n4552), .ZN(n4551) );
  INV_X1 U5418 ( .A(n8297), .ZN(n4552) );
  NAND2_X1 U5419 ( .A1(n8336), .A2(n8297), .ZN(n4553) );
  OR2_X1 U5420 ( .A1(n8792), .A2(n8143), .ZN(n8279) );
  NAND2_X1 U5421 ( .A1(n8792), .A2(n8143), .ZN(n8278) );
  INV_X1 U5422 ( .A(n4578), .ZN(n4577) );
  AND2_X1 U5423 ( .A1(n8175), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U5424 ( .A1(n4580), .A2(n6488), .ZN(n4579) );
  INV_X1 U5425 ( .A(n4580), .ZN(n4576) );
  NOR2_X1 U5426 ( .A1(n8339), .A2(n4581), .ZN(n4580) );
  INV_X1 U5427 ( .A(n8176), .ZN(n4581) );
  INV_X1 U5428 ( .A(n8757), .ZN(n6632) );
  NAND2_X1 U5429 ( .A1(n4556), .A2(n4554), .ZN(n7908) );
  AOI21_X1 U5430 ( .B1(n4305), .B2(n4299), .A(n4555), .ZN(n4554) );
  INV_X1 U5431 ( .A(n8208), .ZN(n4555) );
  OR2_X1 U5432 ( .A1(n6700), .A2(n6681), .ZN(n6941) );
  NOR2_X1 U5433 ( .A1(n6685), .A2(n7045), .ZN(n6947) );
  NAND2_X1 U5434 ( .A1(n5637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5650) );
  INV_X1 U5435 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5649) );
  INV_X1 U5436 ( .A(n6313), .ZN(n5832) );
  INV_X1 U5437 ( .A(n5856), .ZN(n6033) );
  OR4_X1 U5438 ( .A1(n6300), .A2(n6216), .A3(n6245), .A4(n6215), .ZN(n6253) );
  OR2_X1 U5439 ( .A1(n9140), .A2(n5570), .ZN(n6244) );
  INV_X1 U5440 ( .A(n5533), .ZN(n4456) );
  NOR2_X1 U5441 ( .A1(n9404), .A2(n4536), .ZN(n4535) );
  INV_X1 U5442 ( .A(n4537), .ZN(n4536) );
  AOI21_X1 U5443 ( .B1(n9173), .B2(n6176), .A(n6242), .ZN(n4586) );
  AND2_X1 U5444 ( .A1(n9283), .A2(n4524), .ZN(n9215) );
  AND2_X1 U5445 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U5446 ( .A1(n5408), .A2(n4452), .ZN(n4451) );
  INV_X1 U5447 ( .A(n5397), .ZN(n4452) );
  INV_X1 U5448 ( .A(n5408), .ZN(n4453) );
  AND2_X1 U5449 ( .A1(n4543), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5450 ( .A1(n4460), .A2(n5378), .ZN(n4459) );
  NAND2_X1 U5451 ( .A1(n5361), .A2(n5360), .ZN(n4460) );
  NOR2_X1 U5452 ( .A1(n7663), .A2(n7536), .ZN(n4531) );
  NAND2_X1 U5453 ( .A1(n4785), .A2(n6263), .ZN(n4786) );
  NAND2_X1 U5454 ( .A1(n9283), .A2(n4526), .ZN(n9251) );
  INV_X1 U5455 ( .A(n7834), .ZN(n7650) );
  NAND2_X1 U5456 ( .A1(n7535), .A2(n4529), .ZN(n7651) );
  NOR2_X1 U5457 ( .A1(n7511), .A2(n9608), .ZN(n7513) );
  OR3_X1 U5458 ( .A1(n6046), .A2(n6741), .A3(P1_U3086), .ZN(n6740) );
  INV_X1 U5459 ( .A(n5549), .ZN(n5053) );
  AND2_X1 U5460 ( .A1(n5547), .A2(n5049), .ZN(n5536) );
  AOI21_X1 U5461 ( .B1(n4434), .B2(n4432), .A(n4431), .ZN(n4430) );
  INV_X1 U5462 ( .A(n5039), .ZN(n4431) );
  INV_X1 U5463 ( .A(n5035), .ZN(n4432) );
  INV_X1 U5464 ( .A(n4434), .ZN(n4433) );
  INV_X1 U5465 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U5466 ( .A1(n5073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5075) );
  INV_X1 U5467 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U5468 ( .A1(n5075), .A2(n5074), .ZN(n5101) );
  NOR2_X1 U5469 ( .A1(n5418), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U5470 ( .A1(n4809), .A2(n5018), .ZN(n4808) );
  NAND2_X1 U5471 ( .A1(n4810), .A2(n5011), .ZN(n4809) );
  INV_X1 U5472 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U5473 ( .A1(n5381), .A2(SI_16_), .ZN(n4829) );
  AND2_X1 U5474 ( .A1(n4999), .A2(n4998), .ZN(n5000) );
  OR2_X1 U5475 ( .A1(SI_15_), .A2(n4997), .ZN(n4998) );
  AND2_X1 U5476 ( .A1(n4995), .A2(n4994), .ZN(n4996) );
  OR2_X1 U5477 ( .A1(n5350), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U5478 ( .A1(n4978), .A2(n4320), .ZN(n4442) );
  OR2_X1 U5479 ( .A1(n5183), .A2(n4818), .ZN(n4816) );
  OAI21_X1 U5480 ( .B1(n6717), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4948), .ZN(
        n4949) );
  NAND2_X1 U5481 ( .A1(n6717), .A2(n6718), .ZN(n4948) );
  NOR2_X2 U5482 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5174) );
  NAND2_X1 U5483 ( .A1(n6722), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U5484 ( .A1(n6717), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4936) );
  INV_X1 U5485 ( .A(n6731), .ZN(n4607) );
  AND2_X1 U5486 ( .A1(n7792), .A2(n4889), .ZN(n4888) );
  NAND2_X1 U5487 ( .A1(n7766), .A2(n7787), .ZN(n4889) );
  OR2_X1 U5488 ( .A1(n7105), .A2(n7138), .ZN(n7228) );
  INV_X1 U5489 ( .A(n8528), .ZN(n7760) );
  OR2_X1 U5490 ( .A1(n7764), .A2(n7766), .ZN(n7788) );
  INV_X1 U5491 ( .A(n8475), .ZN(n8141) );
  NAND2_X1 U5492 ( .A1(n7916), .A2(n4885), .ZN(n7984) );
  NAND2_X1 U5493 ( .A1(n7788), .A2(n7787), .ZN(n7865) );
  XNOR2_X1 U5494 ( .A(n9854), .B(n7112), .ZN(n7105) );
  NAND2_X1 U5495 ( .A1(n8441), .A2(n8126), .ZN(n8493) );
  OAI21_X1 U5496 ( .B1(n8464), .B2(n8432), .A(n8431), .ZN(n8430) );
  NAND2_X1 U5497 ( .A1(n8313), .A2(n4322), .ZN(n8325) );
  OR2_X1 U5498 ( .A1(n4668), .A2(n4665), .ZN(n8313) );
  AOI21_X1 U5499 ( .B1(n4672), .B2(n8823), .A(n4669), .ZN(n4668) );
  AND2_X1 U5500 ( .A1(n6567), .A2(n6566), .ZN(n8468) );
  INV_X1 U5501 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U5502 ( .A1(n4634), .A2(n5749), .ZN(n9673) );
  OAI21_X1 U5503 ( .B1(n6847), .B2(P2_REG2_REG_1__SCAN_IN), .A(n4395), .ZN(
        n5785) );
  NAND2_X1 U5504 ( .A1(n6847), .A2(n9676), .ZN(n4395) );
  OR2_X1 U5505 ( .A1(n5751), .A2(n6896), .ZN(n4636) );
  NAND3_X1 U5506 ( .A1(n4636), .A2(n7017), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n7019) );
  OR2_X1 U5507 ( .A1(n6887), .A2(n9895), .ZN(n7012) );
  AND2_X1 U5508 ( .A1(n4739), .A2(n9728), .ZN(n4466) );
  XNOR2_X1 U5509 ( .A(n5754), .B(n9710), .ZN(n9720) );
  OR2_X1 U5510 ( .A1(n5723), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U5511 ( .A1(n4741), .A2(n9751), .ZN(n9756) );
  NAND2_X1 U5512 ( .A1(n4742), .A2(n9752), .ZN(n9754) );
  INV_X1 U5513 ( .A(n4743), .ZN(n4742) );
  OAI21_X1 U5514 ( .B1(n7191), .B2(n4613), .A(n4610), .ZN(n9765) );
  INV_X1 U5515 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4612) );
  INV_X1 U5516 ( .A(n4740), .ZN(n5733) );
  AND2_X1 U5517 ( .A1(n4642), .A2(n4641), .ZN(n5763) );
  NAND2_X1 U5518 ( .A1(n7734), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5519 ( .B1(n8049), .B2(n4647), .A(n4646), .ZN(n9777) );
  NAND2_X1 U5520 ( .A1(n4648), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U5521 ( .A1(n5767), .A2(n4648), .ZN(n4646) );
  INV_X1 U5522 ( .A(n9778), .ZN(n4648) );
  NOR2_X1 U5523 ( .A1(n8049), .A2(n8048), .ZN(n8047) );
  AOI21_X1 U5524 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9790), .A(n9777), .ZN(
        n5769) );
  XNOR2_X1 U5525 ( .A(n5739), .B(n8538), .ZN(n8543) );
  OAI21_X1 U5526 ( .B1(n8534), .B2(n4644), .A(n4643), .ZN(n9793) );
  NAND2_X1 U5527 ( .A1(n4645), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U5528 ( .A1(n5770), .A2(n4645), .ZN(n4643) );
  INV_X1 U5529 ( .A(n9794), .ZN(n4645) );
  OAI21_X1 U5530 ( .B1(n8543), .B2(n4478), .A(n4477), .ZN(n9791) );
  NAND2_X1 U5531 ( .A1(n4479), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U5532 ( .A1(n5740), .A2(n4479), .ZN(n4477) );
  INV_X1 U5533 ( .A(n9792), .ZN(n4479) );
  NOR2_X1 U5534 ( .A1(n8543), .A2(n8544), .ZN(n8542) );
  XNOR2_X1 U5535 ( .A(n9810), .B(n5741), .ZN(n9812) );
  NOR2_X1 U5536 ( .A1(n9813), .A2(n9812), .ZN(n9811) );
  AOI21_X1 U5537 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9806), .A(n9793), .ZN(
        n5771) );
  OAI21_X1 U5538 ( .B1(n9737), .B2(n8562), .A(n8561), .ZN(n4397) );
  NAND2_X1 U5539 ( .A1(n8559), .A2(n4391), .ZN(n4398) );
  OR2_X1 U5540 ( .A1(n6593), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U5541 ( .A1(n6543), .A2(n6542), .ZN(n6551) );
  AND4_X1 U5542 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n8693)
         );
  NAND2_X1 U5543 ( .A1(n6504), .A2(n6503), .ZN(n6515) );
  NAND2_X1 U5544 ( .A1(n4629), .A2(n4321), .ZN(n7689) );
  NAND2_X1 U5545 ( .A1(n4630), .A2(n4325), .ZN(n4629) );
  OR2_X1 U5546 ( .A1(n6377), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6385) );
  INV_X1 U5547 ( .A(n8344), .ZN(n9838) );
  OR2_X1 U5548 ( .A1(n8532), .A2(n7055), .ZN(n8181) );
  NAND2_X1 U5549 ( .A1(n6698), .A2(n6950), .ZN(n6946) );
  OR2_X1 U5550 ( .A1(n7048), .A2(n7047), .ZN(n7051) );
  OR2_X1 U5551 ( .A1(n8572), .A2(n8571), .ZN(n8812) );
  NAND2_X1 U5552 ( .A1(n6604), .A2(n6603), .ZN(n6691) );
  OR2_X1 U5553 ( .A1(n8112), .A2(n8317), .ZN(n6604) );
  OR2_X1 U5554 ( .A1(n6601), .A2(n8610), .ZN(n8589) );
  AND2_X1 U5555 ( .A1(n6589), .A2(n6588), .ZN(n8599) );
  AND2_X1 U5556 ( .A1(n8302), .A2(n8303), .ZN(n8616) );
  OR2_X1 U5557 ( .A1(n4907), .A2(n8643), .ZN(n8629) );
  AND2_X1 U5558 ( .A1(n8608), .A2(n8609), .ZN(n8631) );
  AOI21_X1 U5559 ( .B1(n8674), .B2(n4619), .A(n8283), .ZN(n4618) );
  INV_X1 U5560 ( .A(n8675), .ZN(n4619) );
  OR2_X1 U5561 ( .A1(n8730), .A2(n6488), .ZN(n4582) );
  NAND2_X1 U5562 ( .A1(n4582), .A2(n4580), .ZN(n8719) );
  INV_X1 U5563 ( .A(n9890), .ZN(n9873) );
  XNOR2_X1 U5564 ( .A(n5650), .B(n5649), .ZN(n5826) );
  AND2_X1 U5565 ( .A1(n5642), .A2(n5659), .ZN(n6667) );
  OR2_X1 U5566 ( .A1(n5689), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5683) );
  AND2_X1 U5567 ( .A1(n5718), .A2(n5723), .ZN(n9726) );
  INV_X1 U5568 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5714) );
  MUX2_X1 U5569 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5698), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5700) );
  NAND2_X1 U5570 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5698) );
  INV_X1 U5571 ( .A(n5904), .ZN(n4424) );
  OR2_X1 U5572 ( .A1(n5268), .A2(n6977), .ZN(n5282) );
  OR2_X1 U5573 ( .A1(n5990), .A2(n5989), .ZN(n4411) );
  NAND2_X1 U5574 ( .A1(n5319), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5338) );
  INV_X1 U5575 ( .A(n5321), .ZN(n5319) );
  XNOR2_X1 U5576 ( .A(n6009), .B(n6010), .ZN(n8973) );
  OR2_X1 U5577 ( .A1(n5467), .A2(n8976), .ZN(n5484) );
  NAND2_X1 U5578 ( .A1(n5451), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5467) );
  INV_X1 U5579 ( .A(n5453), .ZN(n5451) );
  OAI21_X1 U5580 ( .B1(n4855), .B2(n4854), .A(n4381), .ZN(n4853) );
  INV_X1 U5581 ( .A(n8934), .ZN(n4854) );
  INV_X1 U5582 ( .A(n8995), .ZN(n8983) );
  NAND2_X1 U5583 ( .A1(n5371), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5392) );
  INV_X1 U5584 ( .A(n5372), .ZN(n5371) );
  NOR2_X1 U5585 ( .A1(n4717), .A2(n9398), .ZN(n4716) );
  NAND2_X1 U5586 ( .A1(n6186), .A2(n9020), .ZN(n4717) );
  NOR2_X1 U5587 ( .A1(n4301), .A2(n4310), .ZN(n4501) );
  NOR2_X1 U5588 ( .A1(n4506), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U5589 ( .A1(n4507), .A2(n9119), .ZN(n4505) );
  INV_X1 U5590 ( .A(n6253), .ZN(n4506) );
  NAND2_X1 U5591 ( .A1(n7880), .A2(n5572), .ZN(n4507) );
  INV_X1 U5592 ( .A(n4719), .ZN(n4497) );
  NAND2_X1 U5593 ( .A1(n4687), .A2(n4686), .ZN(n6876) );
  NAND2_X1 U5594 ( .A1(n6776), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4686) );
  INV_X1 U5595 ( .A(n6791), .ZN(n4687) );
  OR2_X1 U5596 ( .A1(n6810), .A2(n6809), .ZN(n4695) );
  NOR2_X1 U5597 ( .A1(n6972), .A2(n4685), .ZN(n6974) );
  AND2_X1 U5598 ( .A1(n6973), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U5599 ( .A1(n6974), .A2(n6975), .ZN(n7073) );
  OR2_X1 U5600 ( .A1(n7277), .A2(n7276), .ZN(n7274) );
  AND2_X1 U5601 ( .A1(n7274), .A2(n7244), .ZN(n7247) );
  NOR2_X1 U5602 ( .A1(n7883), .A2(n4688), .ZN(n9056) );
  AND2_X1 U5603 ( .A1(n7884), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4688) );
  AND2_X1 U5604 ( .A1(n6744), .A2(n6743), .ZN(n6769) );
  AND2_X1 U5605 ( .A1(n5607), .A2(n6869), .ZN(n8982) );
  INV_X1 U5606 ( .A(n9158), .ZN(n9155) );
  NAND2_X1 U5607 ( .A1(n9209), .A2(n4535), .ZN(n9162) );
  INV_X1 U5608 ( .A(n9148), .ZN(n9150) );
  OR2_X1 U5609 ( .A1(n9404), .A2(n5561), .ZN(n9149) );
  NAND2_X1 U5610 ( .A1(n4761), .A2(n4763), .ZN(n4759) );
  NOR2_X1 U5611 ( .A1(n9348), .A2(n9216), .ZN(n9209) );
  NAND2_X1 U5612 ( .A1(n9215), .A2(n4767), .ZN(n9216) );
  AOI21_X1 U5613 ( .B1(n4594), .B2(n9276), .A(n4517), .ZN(n4593) );
  NAND2_X1 U5614 ( .A1(n9283), .A2(n5612), .ZN(n9284) );
  NAND2_X1 U5615 ( .A1(n5424), .A2(n5423), .ZN(n5437) );
  INV_X1 U5616 ( .A(n5426), .ZN(n5424) );
  INV_X1 U5617 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10064) );
  AND2_X1 U5618 ( .A1(n6153), .A2(n6149), .ZN(n9298) );
  INV_X1 U5619 ( .A(n6208), .ZN(n7936) );
  NAND2_X1 U5620 ( .A1(n7650), .A2(n4543), .ZN(n7932) );
  AND2_X1 U5621 ( .A1(n6135), .A2(n6118), .ZN(n7815) );
  AND2_X1 U5622 ( .A1(n5951), .A2(n5575), .ZN(n7644) );
  OAI21_X1 U5623 ( .B1(n7550), .B2(n5344), .A(n5345), .ZN(n7641) );
  OR2_X1 U5624 ( .A1(n5338), .A2(n7707), .ZN(n5354) );
  OR2_X1 U5625 ( .A1(n5354), .A2(n7949), .ZN(n5372) );
  NAND2_X1 U5626 ( .A1(n4585), .A2(n6128), .ZN(n7543) );
  NOR2_X1 U5627 ( .A1(n7551), .A2(n4584), .ZN(n4583) );
  AND2_X1 U5628 ( .A1(n6128), .A2(n6127), .ZN(n7466) );
  NAND2_X1 U5629 ( .A1(n7535), .A2(n4596), .ZN(n7534) );
  INV_X1 U5630 ( .A(n7525), .ZN(n7527) );
  NAND2_X1 U5631 ( .A1(n7529), .A2(n5587), .ZN(n7526) );
  AOI21_X1 U5632 ( .B1(n4754), .B2(n7510), .A(n4345), .ZN(n4753) );
  NAND2_X1 U5633 ( .A1(n4708), .A2(n4508), .ZN(n9505) );
  AOI21_X1 U5634 ( .B1(n4711), .B2(n4713), .A(n4709), .ZN(n4508) );
  INV_X1 U5635 ( .A(n6098), .ZN(n4709) );
  AND2_X1 U5636 ( .A1(n7567), .A2(n7131), .ZN(n4522) );
  INV_X1 U5637 ( .A(n4786), .ZN(n7316) );
  OR2_X1 U5638 ( .A1(n5184), .A2(n6721), .ZN(n5144) );
  OR2_X1 U5639 ( .A1(n5143), .A2(n6726), .ZN(n5145) );
  NAND2_X1 U5640 ( .A1(n9534), .A2(n5577), .ZN(n7562) );
  NAND2_X1 U5641 ( .A1(n4758), .A2(n4761), .ZN(n9191) );
  OR2_X1 U5642 ( .A1(n5493), .A2(n4763), .ZN(n4758) );
  INV_X1 U5643 ( .A(n9620), .ZN(n9551) );
  INV_X1 U5644 ( .A(n7663), .ZN(n9626) );
  INV_X1 U5645 ( .A(n9635), .ZN(n9583) );
  NAND2_X1 U5646 ( .A1(n4291), .A2(n6766), .ZN(n4784) );
  OR2_X1 U5647 ( .A1(n6842), .A2(n5111), .ZN(n9632) );
  AND2_X1 U5648 ( .A1(n5108), .A2(n7312), .ZN(n5621) );
  NAND2_X1 U5649 ( .A1(n9537), .A2(n9644), .ZN(n9635) );
  INV_X1 U5650 ( .A(n6740), .ZN(n9441) );
  XNOR2_X1 U5651 ( .A(n5552), .B(n5551), .ZN(n8113) );
  INV_X1 U5652 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4925) );
  INV_X1 U5653 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U5654 ( .A1(n5077), .A2(n5063), .ZN(n5073) );
  AND2_X1 U5655 ( .A1(n5494), .A2(n5030), .ZN(n5477) );
  INV_X1 U5656 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U5657 ( .A1(n5225), .A2(n4968), .ZN(n5242) );
  NAND2_X1 U5658 ( .A1(n7361), .A2(n4881), .ZN(n7411) );
  AND4_X1 U5659 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n7995)
         );
  NAND2_X1 U5660 ( .A1(n7984), .A2(n7983), .ZN(n8008) );
  AND2_X1 U5661 ( .A1(n4891), .A2(n4892), .ZN(n8401) );
  INV_X1 U5662 ( .A(n8527), .ZN(n7820) );
  AOI21_X1 U5663 ( .B1(n4881), .B2(n7338), .A(n4336), .ZN(n4879) );
  INV_X1 U5664 ( .A(n4881), .ZN(n4880) );
  NAND2_X1 U5665 ( .A1(n8124), .A2(n8123), .ZN(n8442) );
  NAND2_X1 U5666 ( .A1(n7916), .A2(n7915), .ZN(n7918) );
  AND4_X1 U5667 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n8244)
         );
  NAND2_X1 U5668 ( .A1(n6938), .A2(n9834), .ZN(n8501) );
  NAND2_X1 U5669 ( .A1(n4883), .A2(n4341), .ZN(n4882) );
  NAND2_X1 U5670 ( .A1(n7117), .A2(n8390), .ZN(n8514) );
  INV_X1 U5671 ( .A(n8599), .ZN(n8632) );
  NAND2_X1 U5672 ( .A1(n6577), .A2(n6576), .ZN(n8648) );
  NAND2_X1 U5673 ( .A1(n6558), .A2(n6557), .ZN(n8666) );
  INV_X1 U5674 ( .A(n8479), .ZN(n8723) );
  INV_X1 U5675 ( .A(n8748), .ZN(n8521) );
  INV_X1 U5676 ( .A(n7995), .ZN(n8523) );
  INV_X1 U5677 ( .A(n8244), .ZN(n8524) );
  OR2_X1 U5678 ( .A1(n6698), .A2(n5651), .ZN(n8557) );
  NAND2_X1 U5679 ( .A1(n5784), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U5680 ( .A1(n4635), .A2(n7016), .ZN(n7021) );
  NAND2_X1 U5681 ( .A1(n7019), .A2(n7017), .ZN(n4635) );
  AND2_X1 U5682 ( .A1(n7581), .A2(n5732), .ZN(n7732) );
  AND2_X1 U5683 ( .A1(n7579), .A2(n5762), .ZN(n7729) );
  INV_X1 U5684 ( .A(n4734), .ZN(n9776) );
  XNOR2_X1 U5685 ( .A(n5769), .B(n8538), .ZN(n8534) );
  NOR2_X1 U5686 ( .A1(n8534), .A2(n10033), .ZN(n8533) );
  OAI21_X1 U5687 ( .B1(n7294), .B2(n8203), .A(n8226), .ZN(n7428) );
  INV_X1 U5688 ( .A(n8581), .ZN(n8756) );
  INV_X1 U5689 ( .A(n9834), .ZN(n8755) );
  NAND2_X1 U5690 ( .A1(n6661), .A2(n4335), .ZN(n4876) );
  NAND2_X1 U5691 ( .A1(n8752), .A2(n7157), .ZN(n8741) );
  INV_X1 U5692 ( .A(n6939), .ZN(n7055) );
  AND3_X2 U5693 ( .A1(n7048), .A2(n6701), .A3(n6700), .ZN(n9904) );
  AND2_X1 U5694 ( .A1(n8309), .A2(n8308), .ZN(n8817) );
  NOR2_X1 U5695 ( .A1(n8578), .A2(n9885), .ZN(n6665) );
  NAND2_X1 U5696 ( .A1(n6580), .A2(n6579), .ZN(n8826) );
  NAND2_X1 U5697 ( .A1(n6570), .A2(n6569), .ZN(n8832) );
  NAND2_X1 U5698 ( .A1(n6560), .A2(n6559), .ZN(n8837) );
  OAI21_X1 U5699 ( .B1(n8654), .B2(n8289), .A(n8335), .ZN(n8639) );
  NAND2_X1 U5700 ( .A1(n6550), .A2(n6549), .ZN(n8843) );
  NAND2_X1 U5701 ( .A1(n6541), .A2(n6540), .ZN(n8848) );
  NAND2_X1 U5702 ( .A1(n6532), .A2(n6531), .ZN(n8854) );
  NAND2_X1 U5703 ( .A1(n4617), .A2(n8674), .ZN(n8677) );
  NAND2_X1 U5704 ( .A1(n6513), .A2(n6512), .ZN(n8864) );
  NAND2_X1 U5705 ( .A1(n6502), .A2(n6501), .ZN(n8869) );
  NAND2_X1 U5706 ( .A1(n6490), .A2(n6489), .ZN(n8875) );
  NAND2_X1 U5707 ( .A1(n6483), .A2(n6482), .ZN(n8881) );
  AND2_X1 U5708 ( .A1(n8737), .A2(n8736), .ZN(n8879) );
  NAND2_X1 U5709 ( .A1(n6473), .A2(n6472), .ZN(n8888) );
  AND2_X1 U5710 ( .A1(n8751), .A2(n8750), .ZN(n8886) );
  NAND2_X1 U5711 ( .A1(n4567), .A2(n4568), .ZN(n8758) );
  NAND2_X1 U5712 ( .A1(n6464), .A2(n6463), .ZN(n8099) );
  NAND2_X1 U5713 ( .A1(n4570), .A2(n7994), .ZN(n8089) );
  OR2_X1 U5714 ( .A1(n7999), .A2(n8255), .ZN(n4570) );
  NAND2_X1 U5715 ( .A1(n4557), .A2(n4558), .ZN(n7775) );
  OR2_X1 U5716 ( .A1(n6412), .A2(n4299), .ZN(n4557) );
  NAND2_X1 U5717 ( .A1(n6415), .A2(n6414), .ZN(n8207) );
  INV_X1 U5718 ( .A(n8822), .ZN(n8889) );
  NAND2_X1 U5719 ( .A1(n4623), .A2(n4304), .ZN(n7698) );
  NAND2_X1 U5720 ( .A1(n4630), .A2(n4626), .ZN(n4623) );
  OR2_X1 U5721 ( .A1(n9893), .A2(n9873), .ZN(n8822) );
  INV_X2 U5722 ( .A(n9893), .ZN(n9891) );
  AND2_X1 U5723 ( .A1(n5826), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6950) );
  INV_X1 U5724 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6326) );
  INV_X1 U5725 ( .A(n6667), .ZN(n8086) );
  INV_X1 U5726 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U5727 ( .A1(n5645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5636) );
  INV_X1 U5728 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9961) );
  INV_X1 U5729 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7902) );
  INV_X1 U5730 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7878) );
  XNOR2_X1 U5731 ( .A(n5652), .B(n5632), .ZN(n7879) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10021) );
  XNOR2_X1 U5733 ( .A(n6612), .B(n6611), .ZN(n7682) );
  INV_X1 U5734 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7558) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7349) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7289) );
  INV_X1 U5737 ( .A(n6471), .ZN(n9806) );
  OR2_X1 U5738 ( .A1(n5691), .A2(n5690), .ZN(n8073) );
  INV_X1 U5739 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U5740 ( .A1(n5706), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4481) );
  NAND2_X1 U5741 ( .A1(n4749), .A2(n4747), .ZN(n5696) );
  NAND2_X1 U5742 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4748), .ZN(n4747) );
  OAI21_X1 U5743 ( .B1(n5693), .B2(n5694), .A(P2_IR_REG_2__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5744 ( .A1(n5700), .A2(n5699), .ZN(n6724) );
  INV_X1 U5745 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7949) );
  AND2_X1 U5746 ( .A1(n4847), .A2(n5960), .ZN(n7946) );
  NAND2_X1 U5747 ( .A1(n4859), .A2(n4858), .ZN(n8916) );
  NAND2_X1 U5748 ( .A1(n4861), .A2(n4863), .ZN(n4858) );
  AND2_X1 U5749 ( .A1(n4384), .A2(n4316), .ZN(n4414) );
  AND2_X1 U5750 ( .A1(n7476), .A2(n5906), .ZN(n7400) );
  AOI21_X1 U5751 ( .B1(n8964), .B2(n8965), .A(n4901), .ZN(n8925) );
  NAND2_X1 U5752 ( .A1(n4852), .A2(n4855), .ZN(n8933) );
  NAND2_X1 U5753 ( .A1(n8909), .A2(n4856), .ZN(n4852) );
  NAND2_X1 U5754 ( .A1(n4371), .A2(n8950), .ZN(n8949) );
  AOI21_X1 U5755 ( .B1(n8909), .B2(n8910), .A(n4302), .ZN(n8956) );
  INV_X1 U5756 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U5757 ( .A1(n7656), .A2(n7657), .ZN(n4421) );
  NAND2_X1 U5758 ( .A1(n4841), .A2(n7164), .ZN(n7169) );
  OR2_X1 U5759 ( .A1(n6065), .A2(P1_U3086), .ZN(n8998) );
  AND2_X1 U5760 ( .A1(n4851), .A2(n4848), .ZN(n8992) );
  INV_X1 U5761 ( .A(n4853), .ZN(n4848) );
  INV_X1 U5762 ( .A(n9001), .ZN(n9011) );
  INV_X1 U5763 ( .A(n8998), .ZN(n9013) );
  OR2_X1 U5764 ( .A1(n8959), .A2(n5563), .ZN(n5510) );
  INV_X1 U5765 ( .A(n5219), .ZN(n9042) );
  NAND4_X1 U5766 ( .A1(n5196), .A2(n5195), .A3(n5194), .A4(n5193), .ZN(n9043)
         );
  NAND4_X1 U5767 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n9045)
         );
  INV_X1 U5768 ( .A(P1_U3973), .ZN(n9046) );
  NAND2_X1 U5769 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4697) );
  NOR2_X1 U5770 ( .A1(n9487), .A2(n4326), .ZN(n6793) );
  NOR2_X1 U5771 ( .A1(n6793), .A2(n6792), .ZN(n6791) );
  AND2_X1 U5772 ( .A1(n6875), .A2(n4696), .ZN(n6810) );
  NAND2_X1 U5773 ( .A1(n6766), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4696) );
  INV_X1 U5774 ( .A(n4695), .ZN(n6808) );
  NOR2_X1 U5775 ( .A1(n6902), .A2(n4370), .ZN(n6905) );
  NOR2_X1 U5776 ( .A1(n6905), .A2(n6904), .ZN(n6972) );
  AND2_X1 U5777 ( .A1(n5316), .A2(n5350), .ZN(n7386) );
  NOR2_X1 U5778 ( .A1(n7666), .A2(n4689), .ZN(n7670) );
  AND2_X1 U5779 ( .A1(n7667), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5780 ( .A1(n7670), .A2(n7669), .ZN(n7883) );
  XNOR2_X1 U5781 ( .A(n9056), .B(n9055), .ZN(n7885) );
  NOR2_X1 U5782 ( .A1(n9472), .A2(n6869), .ZN(n9478) );
  OR2_X1 U5783 ( .A1(n9102), .A2(n9101), .ZN(n9113) );
  NOR2_X1 U5784 ( .A1(n9123), .A2(n9620), .ZN(n9327) );
  NAND2_X1 U5785 ( .A1(n4760), .A2(n4766), .ZN(n9199) );
  NAND2_X1 U5786 ( .A1(n5493), .A2(n4764), .ZN(n4760) );
  NAND2_X1 U5787 ( .A1(n5592), .A2(n6218), .ZN(n9221) );
  NAND2_X1 U5788 ( .A1(n5493), .A2(n5492), .ZN(n9214) );
  AND2_X1 U5789 ( .A1(n9278), .A2(n6154), .ZN(n9258) );
  NAND2_X1 U5790 ( .A1(n4768), .A2(n4769), .ZN(n9262) );
  NAND2_X1 U5791 ( .A1(n4774), .A2(n5431), .ZN(n9277) );
  NAND2_X1 U5792 ( .A1(n4775), .A2(n4367), .ZN(n4774) );
  INV_X1 U5793 ( .A(n9291), .ZN(n4775) );
  NAND2_X1 U5794 ( .A1(n5422), .A2(n5421), .ZN(n9380) );
  NAND2_X1 U5795 ( .A1(n7937), .A2(n5408), .ZN(n4777) );
  NAND2_X1 U5796 ( .A1(n5387), .A2(n5386), .ZN(n8946) );
  NAND2_X1 U5797 ( .A1(n4756), .A2(n5261), .ZN(n7509) );
  NAND2_X1 U5798 ( .A1(n7491), .A2(n7492), .ZN(n4756) );
  INV_X1 U5799 ( .A(n9542), .ZN(n9294) );
  OR2_X1 U5800 ( .A1(n9543), .A2(n7315), .ZN(n9325) );
  OR2_X1 U5801 ( .A1(n9543), .A2(n7321), .ZN(n9545) );
  INV_X1 U5802 ( .A(n9272), .ZN(n9554) );
  NAND2_X1 U5803 ( .A1(n6743), .A2(n9453), .ZN(n4725) );
  INV_X1 U5804 ( .A(n9545), .ZN(n9296) );
  AND2_X2 U5805 ( .A1(n5621), .A2(n6044), .ZN(n10083) );
  NAND2_X1 U5806 ( .A1(n6185), .A2(n6184), .ZN(n9401) );
  INV_X1 U5807 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4599) );
  AND2_X1 U5808 ( .A1(n5527), .A2(n5526), .ZN(n9413) );
  NAND2_X1 U5809 ( .A1(n5450), .A2(n5449), .ZN(n9427) );
  AND2_X1 U5810 ( .A1(n5414), .A2(n5413), .ZN(n9437) );
  AND2_X2 U5811 ( .A1(n5621), .A2(n7313), .ZN(n9650) );
  AND2_X1 U5812 ( .A1(n9442), .A2(n9441), .ZN(n9558) );
  NAND2_X1 U5813 ( .A1(n4928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4929) );
  INV_X1 U5814 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U5815 ( .A1(n5069), .A2(n4425), .ZN(n7992) );
  AND2_X1 U5816 ( .A1(n5176), .A2(n4923), .ZN(n4426) );
  INV_X1 U5817 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7980) );
  INV_X1 U5818 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7882) );
  INV_X1 U5819 ( .A(n6316), .ZN(n7880) );
  INV_X1 U5820 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7721) );
  INV_X1 U5821 ( .A(n5572), .ZN(n7723) );
  INV_X1 U5822 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7288) );
  INV_X1 U5823 ( .A(n9049), .ZN(n9055) );
  INV_X1 U5824 ( .A(n5330), .ZN(n5332) );
  NAND2_X1 U5825 ( .A1(n4824), .A2(n4823), .ZN(n5310) );
  NAND2_X1 U5826 ( .A1(n4824), .A2(n4825), .ZN(n5309) );
  NAND2_X1 U5827 ( .A1(n4819), .A2(n4955), .ZN(n5199) );
  XNOR2_X1 U5828 ( .A(n5200), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6813) );
  INV_X2 U5829 ( .A(n8557), .ZN(P2_U3893) );
  NAND2_X1 U5830 ( .A1(n9809), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6854) );
  AOI21_X1 U5831 ( .B1(n4746), .B2(n9758), .A(n4744), .ZN(n8568) );
  OR2_X1 U5832 ( .A1(n4329), .A2(n8563), .ZN(n4746) );
  NAND2_X1 U5833 ( .A1(n4470), .A2(n9758), .ZN(n4469) );
  NOR2_X1 U5834 ( .A1(n4653), .A2(n4468), .ZN(n4467) );
  XNOR2_X1 U5835 ( .A(n5747), .B(n5820), .ZN(n4470) );
  NAND2_X1 U5836 ( .A1(n4869), .A2(n9007), .ZN(n4868) );
  AND2_X1 U5837 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  OAI21_X1 U5838 ( .B1(n9120), .B2(n9119), .A(n4690), .ZN(P1_U3262) );
  AOI21_X1 U5839 ( .B1(n4692), .B2(n9119), .A(n4691), .ZN(n4690) );
  AND2_X1 U5840 ( .A1(n9140), .A2(n9373), .ZN(n5620) );
  NAND2_X1 U5841 ( .A1(n4465), .A2(n4463), .ZN(P1_U3550) );
  AOI21_X1 U5842 ( .B1(n9404), .B2(n9373), .A(n4464), .ZN(n4463) );
  NAND2_X1 U5843 ( .A1(n9403), .A2(n10083), .ZN(n4465) );
  NOR2_X1 U5844 ( .A1(n10083), .A2(n9984), .ZN(n4464) );
  NAND2_X1 U5845 ( .A1(n9178), .A2(n9373), .ZN(n4393) );
  AOI21_X1 U5846 ( .B1(n9403), .B2(n9650), .A(n4597), .ZN(n9405) );
  NAND2_X1 U5847 ( .A1(n4600), .A2(n4598), .ZN(n4597) );
  OR2_X1 U5848 ( .A1(n9650), .A2(n4599), .ZN(n4598) );
  OAI21_X1 U5849 ( .B1(n9451), .B2(n9452), .A(n4864), .ZN(P1_U3325) );
  INV_X1 U5850 ( .A(n4865), .ZN(n4864) );
  INV_X2 U5851 ( .A(n6031), .ZN(n5848) );
  NAND2_X1 U5852 ( .A1(n8206), .A2(n8225), .ZN(n4299) );
  OR2_X1 U5853 ( .A1(n5197), .A2(n4957), .ZN(n4300) );
  AND2_X1 U5854 ( .A1(n6255), .A2(n5833), .ZN(n4301) );
  INV_X1 U5855 ( .A(n6346), .ZN(n6474) );
  INV_X1 U5856 ( .A(n6474), .ZN(n6553) );
  AND2_X1 U5857 ( .A1(n6018), .A2(n6017), .ZN(n4302) );
  NAND2_X1 U5858 ( .A1(n8483), .A2(n4893), .ZN(n4892) );
  AND2_X1 U5859 ( .A1(n4422), .A2(n7706), .ZN(n4303) );
  INV_X1 U5860 ( .A(n7338), .ZN(n7335) );
  OR2_X1 U5861 ( .A1(n4627), .A2(n4906), .ZN(n4304) );
  INV_X1 U5862 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6323) );
  OR2_X1 U5863 ( .A1(n9398), .A2(n9019), .ZN(n6308) );
  AND2_X1 U5864 ( .A1(n4558), .A2(n8236), .ZN(n4305) );
  AND2_X1 U5865 ( .A1(n4353), .A2(n4451), .ZN(n4306) );
  NAND2_X1 U5866 ( .A1(n7450), .A2(n5219), .ZN(n6197) );
  INV_X1 U5867 ( .A(n6197), .ZN(n4712) );
  INV_X1 U5868 ( .A(n6159), .ZN(n4517) );
  NAND2_X1 U5869 ( .A1(n9626), .A2(n7545), .ZN(n6128) );
  INV_X1 U5870 ( .A(n6128), .ZN(n4584) );
  NAND2_X1 U5871 ( .A1(n5172), .A2(n4323), .ZN(n9044) );
  INV_X1 U5872 ( .A(n9044), .ZN(n4462) );
  OR2_X1 U5873 ( .A1(n9413), .A2(n9024), .ZN(n6288) );
  AND2_X1 U5874 ( .A1(n4898), .A2(n7828), .ZN(n4307) );
  AND2_X1 U5875 ( .A1(n4833), .A2(n4838), .ZN(n4308) );
  AND2_X1 U5876 ( .A1(n4652), .A2(n6638), .ZN(n4309) );
  NAND2_X1 U5877 ( .A1(n6308), .A2(n5572), .ZN(n4310) );
  NAND2_X1 U5878 ( .A1(n8224), .A2(n7418), .ZN(n4311) );
  BUF_X1 U5879 ( .A(n5139), .Z(n6743) );
  AND2_X1 U5880 ( .A1(n4955), .A2(n4951), .ZN(n4312) );
  NOR2_X1 U5881 ( .A1(n5960), .A2(n4844), .ZN(n4313) );
  INV_X1 U5882 ( .A(n5582), .ZN(n4714) );
  INV_X1 U5883 ( .A(n7420), .ZN(n4630) );
  NAND2_X1 U5884 ( .A1(n6412), .A2(n6411), .ZN(n7686) );
  OR2_X1 U5885 ( .A1(n6413), .A2(n5781), .ZN(n4314) );
  INV_X1 U5886 ( .A(n5495), .ZN(n5034) );
  INV_X1 U5887 ( .A(n8688), .ZN(n4616) );
  OR2_X1 U5888 ( .A1(n5381), .A2(SI_16_), .ZN(n4315) );
  NAND2_X1 U5889 ( .A1(n5974), .A2(n5973), .ZN(n4316) );
  AND2_X1 U5890 ( .A1(n4529), .A2(n4532), .ZN(n4317) );
  AND2_X1 U5891 ( .A1(n4368), .A2(n7567), .ZN(n4318) );
  INV_X2 U5892 ( .A(n5267), .ZN(n5601) );
  OR2_X1 U5893 ( .A1(n7816), .A2(n7815), .ZN(n4319) );
  AND2_X1 U5894 ( .A1(n6714), .A2(n5832), .ZN(n5854) );
  NAND2_X1 U5895 ( .A1(n5693), .A2(n4748), .ZN(n5695) );
  NAND3_X1 U5896 ( .A1(n6345), .A2(n6344), .A3(n6343), .ZN(n6615) );
  OR2_X1 U5897 ( .A1(n4973), .A2(SI_9_), .ZN(n4320) );
  NAND2_X1 U5898 ( .A1(n6643), .A2(n6642), .ZN(n8640) );
  OR2_X1 U5899 ( .A1(n9883), .A2(n8528), .ZN(n4321) );
  OR2_X1 U5900 ( .A1(n8312), .A2(n8311), .ZN(n4322) );
  AND3_X1 U5901 ( .A1(n5171), .A2(n5170), .A3(n5169), .ZN(n4323) );
  INV_X1 U5902 ( .A(n4821), .ZN(n4820) );
  OAI21_X1 U5903 ( .B1(n4827), .B2(n4822), .A(n4982), .ZN(n4821) );
  NAND2_X1 U5904 ( .A1(n5263), .A2(n5262), .ZN(n4443) );
  NAND2_X1 U5905 ( .A1(n6640), .A2(n8688), .ZN(n8673) );
  NAND2_X1 U5906 ( .A1(n7026), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5709) );
  INV_X1 U5907 ( .A(n5709), .ZN(n4737) );
  OAI21_X1 U5908 ( .B1(n8916), .B2(n8917), .A(n4411), .ZN(n8964) );
  OR2_X1 U5909 ( .A1(n6602), .A2(n8592), .ZN(n4324) );
  NAND2_X1 U5910 ( .A1(n9883), .A2(n8528), .ZN(n4325) );
  INV_X1 U5911 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4748) );
  AND2_X1 U5912 ( .A1(n6777), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U5913 ( .A1(n6661), .A2(n6717), .ZN(n6351) );
  XOR2_X1 U5914 ( .A(n5127), .B(n5126), .Z(n4327) );
  NAND2_X1 U5915 ( .A1(n5298), .A2(n5297), .ZN(n7536) );
  OR2_X1 U5916 ( .A1(n8207), .A2(n8526), .ZN(n4328) );
  AOI21_X1 U5917 ( .B1(n8430), .B2(n8506), .A(n8507), .ZN(n8505) );
  AND2_X1 U5918 ( .A1(n8565), .A2(n8564), .ZN(n4329) );
  OR3_X1 U5919 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4330) );
  AND2_X1 U5920 ( .A1(n5631), .A2(n5664), .ZN(n6609) );
  AND2_X1 U5921 ( .A1(n4885), .A2(n8007), .ZN(n4331) );
  NOR2_X1 U5922 ( .A1(n8641), .A2(n4907), .ZN(n4333) );
  INV_X1 U5923 ( .A(n4710), .ZN(n7442) );
  AND2_X1 U5924 ( .A1(n8348), .A2(n8222), .ZN(n4334) );
  AND2_X1 U5925 ( .A1(n4327), .A2(n6722), .ZN(n4335) );
  AND2_X1 U5926 ( .A1(n7410), .A2(n7422), .ZN(n4336) );
  NOR2_X1 U5927 ( .A1(n8542), .A2(n5740), .ZN(n4337) );
  NOR2_X1 U5928 ( .A1(n8533), .A2(n5770), .ZN(n4338) );
  AND2_X1 U5929 ( .A1(n5724), .A2(n5729), .ZN(n6391) );
  INV_X1 U5930 ( .A(n6391), .ZN(n7195) );
  NOR2_X1 U5931 ( .A1(n9889), .A2(n8527), .ZN(n4339) );
  NAND2_X1 U5932 ( .A1(n5641), .A2(n5640), .ZN(n5659) );
  AND2_X1 U5933 ( .A1(n8251), .A2(n8250), .ZN(n4340) );
  NAND2_X1 U5934 ( .A1(n8006), .A2(n8005), .ZN(n4341) );
  AND2_X1 U5935 ( .A1(n8276), .A2(n8273), .ZN(n4342) );
  AND2_X1 U5936 ( .A1(n4769), .A2(n5461), .ZN(n4343) );
  OR2_X1 U5937 ( .A1(n9640), .A2(n5574), .ZN(n7828) );
  NAND2_X1 U5938 ( .A1(n8254), .A2(n8248), .ZN(n4344) );
  OR2_X1 U5939 ( .A1(n8255), .A2(n8256), .ZN(n8341) );
  INV_X1 U5940 ( .A(n8341), .ZN(n4661) );
  NOR2_X1 U5941 ( .A1(n9608), .A2(n9039), .ZN(n4345) );
  NAND2_X1 U5942 ( .A1(n4626), .A2(n6622), .ZN(n4346) );
  OR2_X1 U5943 ( .A1(n9348), .A2(n9025), .ZN(n4347) );
  INV_X1 U5944 ( .A(n4826), .ZN(n4825) );
  NOR2_X1 U5945 ( .A1(n4980), .A2(SI_11_), .ZN(n4826) );
  NAND2_X1 U5946 ( .A1(n6609), .A2(n6611), .ZN(n5653) );
  NAND2_X1 U5947 ( .A1(n4443), .A2(n4320), .ZN(n4348) );
  INV_X1 U5948 ( .A(n4906), .ZN(n4631) );
  AND2_X1 U5949 ( .A1(n4908), .A2(n8208), .ZN(n4349) );
  NAND2_X1 U5950 ( .A1(n8972), .A2(n6012), .ZN(n8909) );
  AND2_X1 U5951 ( .A1(n4971), .A2(n4970), .ZN(n4350) );
  NAND2_X1 U5952 ( .A1(n6127), .A2(n6126), .ZN(n4351) );
  INV_X1 U5953 ( .A(n4595), .ZN(n4594) );
  NAND2_X1 U5954 ( .A1(n9261), .A2(n6154), .ZN(n4595) );
  NAND2_X1 U5955 ( .A1(n4516), .A2(n4519), .ZN(n4352) );
  AND2_X1 U5956 ( .A1(n4905), .A2(n5409), .ZN(n4353) );
  AND2_X1 U5957 ( .A1(n5185), .A2(n4784), .ZN(n4354) );
  NAND2_X1 U5958 ( .A1(n5955), .A2(n4846), .ZN(n4355) );
  INV_X1 U5959 ( .A(n6179), .ZN(n4489) );
  OR2_X1 U5960 ( .A1(n9172), .A2(n9173), .ZN(n4356) );
  NOR3_X1 U5961 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4357) );
  AND2_X1 U5962 ( .A1(n9190), .A2(n4759), .ZN(n4358) );
  AND2_X1 U5963 ( .A1(n5594), .A2(n6218), .ZN(n4359) );
  AND2_X1 U5964 ( .A1(n5632), .A2(n4896), .ZN(n4360) );
  AND2_X1 U5965 ( .A1(n6626), .A2(n6625), .ZN(n4361) );
  NAND2_X1 U5966 ( .A1(n6850), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4362) );
  AND2_X1 U5967 ( .A1(n6146), .A2(n6148), .ZN(n9309) );
  OR2_X1 U5968 ( .A1(n5653), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4363) );
  INV_X1 U5969 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4933) );
  AND2_X1 U5970 ( .A1(n4398), .A2(n4396), .ZN(n4364) );
  INV_X1 U5971 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U5972 ( .A1(n4437), .A2(n4820), .ZN(n5330) );
  INV_X1 U5973 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4698) );
  XNOR2_X1 U5974 ( .A(n5078), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5572) );
  AND2_X1 U5975 ( .A1(n7650), .A2(n9018), .ZN(n4365) );
  OR2_X1 U5976 ( .A1(n9023), .A2(n9178), .ZN(n4366) );
  INV_X1 U5977 ( .A(n9477), .ZN(n6778) );
  XNOR2_X1 U5978 ( .A(n4697), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9477) );
  OR2_X1 U5979 ( .A1(n9380), .A2(n9030), .ZN(n4367) );
  AND2_X1 U5980 ( .A1(n7323), .A2(n9573), .ZN(n4368) );
  AND2_X1 U5981 ( .A1(n7650), .A2(n4541), .ZN(n4369) );
  INV_X1 U5982 ( .A(n6413), .ZN(n7734) );
  AND2_X1 U5983 ( .A1(n6906), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U5984 ( .A1(n4777), .A2(n5409), .ZN(n9308) );
  OAI21_X1 U5985 ( .B1(n7641), .B2(n5361), .A(n5360), .ZN(n7832) );
  NAND2_X1 U5986 ( .A1(n5329), .A2(n5328), .ZN(n7550) );
  NAND2_X1 U5987 ( .A1(n4421), .A2(n5946), .ZN(n7705) );
  AND3_X1 U5988 ( .A1(n4415), .A2(n4316), .A3(n4412), .ZN(n4371) );
  AND2_X1 U5989 ( .A1(n9283), .A2(n4528), .ZN(n4372) );
  INV_X1 U5990 ( .A(n5010), .ZN(n4811) );
  AND2_X1 U5991 ( .A1(n9437), .A2(n8918), .ZN(n4373) );
  NAND2_X1 U5992 ( .A1(n5500), .A2(n5499), .ZN(n9354) );
  INV_X1 U5993 ( .A(n9354), .ZN(n4767) );
  NAND2_X1 U5994 ( .A1(n5466), .A2(n5465), .ZN(n6008) );
  INV_X1 U5995 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U5996 ( .A1(n6631), .A2(n6630), .ZN(n8743) );
  INV_X1 U5997 ( .A(n8369), .ZN(n4670) );
  NAND2_X1 U5998 ( .A1(n5554), .A2(n5553), .ZN(n9404) );
  NOR2_X1 U5999 ( .A1(n8047), .A2(n5767), .ZN(n4374) );
  AND2_X1 U6000 ( .A1(n4582), .A2(n8176), .ZN(n4375) );
  INV_X1 U6001 ( .A(n7835), .ZN(n9018) );
  NAND2_X1 U6002 ( .A1(n5370), .A2(n5369), .ZN(n7835) );
  AND2_X1 U6003 ( .A1(n8282), .A2(n8287), .ZN(n8674) );
  INV_X1 U6004 ( .A(n8674), .ZN(n4620) );
  AND2_X1 U6005 ( .A1(n4637), .A2(n6625), .ZN(n4376) );
  NOR2_X1 U6006 ( .A1(n8854), .A2(n8694), .ZN(n4377) );
  NAND2_X1 U6007 ( .A1(n6592), .A2(n6591), .ZN(n8770) );
  INV_X1 U6008 ( .A(n4772), .ZN(n4771) );
  NOR2_X1 U6009 ( .A1(n5445), .A2(n4773), .ZN(n4772) );
  INV_X1 U6010 ( .A(n5951), .ZN(n9633) );
  NAND2_X1 U6011 ( .A1(n5337), .A2(n5336), .ZN(n5951) );
  AND2_X1 U6012 ( .A1(n8949), .A2(n4860), .ZN(n4378) );
  NAND2_X1 U6013 ( .A1(n4354), .A2(n5186), .ZN(n9580) );
  INV_X1 U6014 ( .A(n9580), .ZN(n7323) );
  AND2_X1 U6015 ( .A1(n8277), .A2(n8684), .ZN(n8702) );
  NOR2_X1 U6016 ( .A1(n6024), .A2(n6023), .ZN(n4379) );
  XNOR2_X1 U6017 ( .A(n6055), .B(n6057), .ZN(n4380) );
  INV_X1 U6018 ( .A(n4380), .ZN(n4869) );
  NAND2_X1 U6019 ( .A1(n6030), .A2(n6029), .ZN(n4381) );
  OR2_X1 U6020 ( .A1(SI_20_), .A2(n5018), .ZN(n4382) );
  INV_X1 U6021 ( .A(n4901), .ZN(n4410) );
  OR2_X1 U6022 ( .A1(n5398), .A2(n4446), .ZN(n4383) );
  INV_X1 U6023 ( .A(n4861), .ZN(n4860) );
  NAND2_X1 U6024 ( .A1(n8306), .A2(n8330), .ZN(n8368) );
  INV_X1 U6025 ( .A(n8368), .ZN(n4676) );
  AND2_X1 U6026 ( .A1(n4863), .A2(n8950), .ZN(n4384) );
  AND2_X1 U6027 ( .A1(n4856), .A2(n8934), .ZN(n4385) );
  AND2_X1 U6028 ( .A1(n4568), .A2(n8265), .ZN(n4386) );
  AND2_X1 U6029 ( .A1(n8278), .A2(n8684), .ZN(n4387) );
  INV_X1 U6030 ( .A(n4572), .ZN(n4571) );
  OAI21_X1 U6031 ( .B1(n4573), .B2(n8256), .A(n8261), .ZN(n4572) );
  NOR2_X1 U6032 ( .A1(n6568), .A2(n4551), .ZN(n4550) );
  INV_X1 U6033 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U6034 ( .A1(n5481), .A2(n5480), .ZN(n9235) );
  INV_X1 U6035 ( .A(n9235), .ZN(n4525) );
  NAND2_X1 U6036 ( .A1(n5402), .A2(n5401), .ZN(n7933) );
  INV_X1 U6037 ( .A(n7933), .ZN(n4542) );
  INV_X1 U6038 ( .A(n5833), .ZN(n9119) );
  INV_X1 U6039 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4726) );
  XNOR2_X1 U6040 ( .A(n5070), .B(n4925), .ZN(n8088) );
  INV_X1 U6041 ( .A(n8088), .ZN(n5104) );
  INV_X1 U6042 ( .A(n7492), .ZN(n4752) );
  AND2_X1 U6043 ( .A1(n7535), .A2(n4531), .ZN(n4388) );
  NAND2_X1 U6044 ( .A1(n7264), .A2(n7256), .ZN(n7292) );
  NAND2_X1 U6045 ( .A1(n7169), .A2(n5894), .ZN(n7176) );
  INV_X1 U6046 ( .A(n6261), .ZN(n4713) );
  NAND2_X1 U6047 ( .A1(n5436), .A2(n5435), .ZN(n9377) );
  NAND2_X1 U6048 ( .A1(n7061), .A2(n5878), .ZN(n7063) );
  NAND4_X1 U6049 ( .A1(n4835), .A2(n4308), .A3(n4834), .A4(n4424), .ZN(n7476)
         );
  NAND2_X1 U6050 ( .A1(n4401), .A2(n5889), .ZN(n7124) );
  NOR2_X1 U6051 ( .A1(n7230), .A2(n7225), .ZN(n4389) );
  NAND2_X1 U6052 ( .A1(n7336), .A2(n7335), .ZN(n7361) );
  INV_X1 U6053 ( .A(SI_20_), .ZN(n10036) );
  NAND2_X1 U6054 ( .A1(n4368), .A2(n4522), .ZN(n4523) );
  NAND2_X1 U6055 ( .A1(n5538), .A2(n5537), .ZN(n9178) );
  AND2_X1 U6056 ( .A1(n7361), .A2(n7360), .ZN(n4390) );
  NOR2_X1 U6057 ( .A1(n9552), .A2(n5611), .ZN(n7567) );
  NAND2_X1 U6058 ( .A1(n5353), .A2(n5352), .ZN(n9640) );
  INV_X1 U6059 ( .A(n9640), .ZN(n4532) );
  NAND2_X1 U6060 ( .A1(n6316), .A2(n5833), .ZN(n5834) );
  AND2_X1 U6061 ( .A1(n9822), .A2(n8558), .ZN(n4391) );
  OR2_X1 U6062 ( .A1(n6852), .A2(n8385), .ZN(n9826) );
  INV_X1 U6063 ( .A(n6192), .ZN(n4727) );
  AND2_X1 U6064 ( .A1(n5726), .A2(n9752), .ZN(n4392) );
  NOR2_X1 U6065 ( .A1(n6325), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8894) );
  INV_X1 U6066 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n4639) );
  INV_X1 U6067 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n4475) );
  XNOR2_X1 U6068 ( .A(n5766), .B(n8118), .ZN(n8049) );
  NAND2_X1 U6069 ( .A1(n5622), .A2(n10083), .ZN(n5618) );
  NAND2_X1 U6070 ( .A1(n5614), .A2(n5615), .ZN(n5622) );
  NAND2_X1 U6071 ( .A1(n8217), .A2(n8200), .ZN(n8197) );
  OAI21_X2 U6072 ( .B1(n9204), .B2(n9203), .A(n6171), .ZN(n9187) );
  NAND3_X1 U6073 ( .A1(n7200), .A2(n6619), .A3(n7258), .ZN(n7264) );
  NAND2_X1 U6074 ( .A1(n9230), .A2(n9233), .ZN(n5592) );
  NAND2_X1 U6075 ( .A1(n4926), .A2(n4925), .ZN(n4932) );
  NAND2_X1 U6076 ( .A1(n8711), .A2(n8340), .ZN(n4652) );
  NAND2_X1 U6077 ( .A1(n7903), .A2(n6624), .ZN(n4637) );
  NAND2_X1 U6078 ( .A1(n6631), .A2(n4649), .ZN(n8742) );
  NAND2_X1 U6079 ( .A1(n6643), .A2(n4650), .ZN(n8628) );
  NAND2_X1 U6080 ( .A1(n7926), .A2(n6143), .ZN(n9312) );
  NAND2_X1 U6081 ( .A1(n4614), .A2(n4618), .ZN(n8663) );
  NAND2_X1 U6082 ( .A1(n9520), .A2(n6265), .ZN(n4699) );
  AOI21_X2 U6083 ( .B1(n7317), .B2(n6263), .A(n5581), .ZN(n7090) );
  NAND2_X1 U6084 ( .A1(n9341), .A2(n4393), .ZN(P1_U3549) );
  NAND2_X1 U6085 ( .A1(n4394), .A2(n9541), .ZN(n9176) );
  NAND2_X1 U6086 ( .A1(n9171), .A2(n4356), .ZN(n4394) );
  INV_X4 U6087 ( .A(n5430), .ZN(n6088) );
  INV_X1 U6088 ( .A(n9312), .ZN(n4400) );
  INV_X1 U6089 ( .A(n6107), .ZN(n4399) );
  NAND2_X1 U6090 ( .A1(n4399), .A2(n6101), .ZN(n5583) );
  NAND2_X1 U6091 ( .A1(n5657), .A2(n5656), .ZN(n6322) );
  NAND2_X1 U6092 ( .A1(n8536), .A2(n8537), .ZN(n8535) );
  NAND2_X1 U6093 ( .A1(n4469), .A2(n4467), .ZN(P2_U3201) );
  INV_X1 U6094 ( .A(n5831), .ZN(n4653) );
  NOR2_X1 U6095 ( .A1(n9739), .A2(n5794), .ZN(n7190) );
  NOR2_X1 U6096 ( .A1(n9760), .A2(n5799), .ZN(n7578) );
  NOR2_X1 U6097 ( .A1(n5807), .A2(n8074), .ZN(n8033) );
  NOR2_X1 U6098 ( .A1(n5804), .A2(n7724), .ZN(n8075) );
  NAND2_X1 U6099 ( .A1(n9780), .A2(n5813), .ZN(n8536) );
  NAND2_X1 U6100 ( .A1(n4364), .A2(n4745), .ZN(n4744) );
  INV_X1 U6101 ( .A(n5058), .ZN(n4924) );
  NAND2_X1 U6102 ( .A1(n5061), .A2(n4922), .ZN(n5058) );
  NAND2_X1 U6103 ( .A1(n7502), .A2(n6121), .ZN(n6107) );
  OAI21_X2 U6104 ( .B1(n7807), .B2(n7806), .A(n6135), .ZN(n7927) );
  NAND3_X1 U6105 ( .A1(n4415), .A2(n4414), .A3(n4412), .ZN(n4859) );
  NAND2_X1 U6106 ( .A1(n9004), .A2(n5967), .ZN(n8940) );
  NAND2_X1 U6107 ( .A1(n9006), .A2(n9005), .ZN(n9004) );
  INV_X1 U6108 ( .A(n8941), .ZN(n4417) );
  OAI21_X1 U6109 ( .B1(n7656), .B2(n4423), .A(n4303), .ZN(n5956) );
  NAND2_X1 U6110 ( .A1(n4419), .A2(n4420), .ZN(n4843) );
  NAND2_X1 U6111 ( .A1(n7656), .A2(n4303), .ZN(n4419) );
  NAND3_X1 U6112 ( .A1(n5906), .A2(n7401), .A3(n7476), .ZN(n7399) );
  NAND3_X1 U6113 ( .A1(n4835), .A2(n4308), .A3(n4834), .ZN(n5905) );
  NAND2_X1 U6114 ( .A1(n5476), .A2(n4430), .ZN(n4429) );
  NAND4_X1 U6115 ( .A1(n5001), .A2(n5000), .A3(n4315), .A4(n5006), .ZN(n4444)
         );
  NAND3_X1 U6116 ( .A1(n5001), .A2(n5000), .A3(n4315), .ZN(n4447) );
  NAND3_X1 U6117 ( .A1(n8588), .A2(n6600), .A3(n4550), .ZN(n4548) );
  NAND2_X1 U6118 ( .A1(n4319), .A2(n4306), .ZN(n4450) );
  NAND2_X1 U6119 ( .A1(n5534), .A2(n4455), .ZN(n4454) );
  NAND3_X1 U6120 ( .A1(n4739), .A2(P2_REG1_REG_5__SCAN_IN), .A3(n9728), .ZN(
        n9730) );
  OAI21_X1 U6121 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n4466), .A(n9730), .ZN(
        n9711) );
  NAND2_X1 U6122 ( .A1(n9732), .A2(n5721), .ZN(n5725) );
  INV_X1 U6123 ( .A(n4476), .ZN(n7730) );
  XNOR2_X2 U6124 ( .A(n4482), .B(n5114), .ZN(n5119) );
  NAND3_X1 U6125 ( .A1(n4493), .A2(n4490), .A3(n4489), .ZN(n4488) );
  OAI21_X1 U6126 ( .B1(n4498), .B2(n4497), .A(n4500), .ZN(n4499) );
  INV_X1 U6127 ( .A(n4499), .ZN(n6256) );
  INV_X1 U6128 ( .A(n4715), .ZN(n4502) );
  NAND2_X1 U6129 ( .A1(n6157), .A2(n4512), .ZN(n4509) );
  NAND2_X1 U6130 ( .A1(n4509), .A2(n4510), .ZN(n6163) );
  NAND2_X1 U6131 ( .A1(n6235), .A2(n6096), .ZN(n4519) );
  NAND2_X1 U6132 ( .A1(n7567), .A2(n9573), .ZN(n9529) );
  INV_X1 U6133 ( .A(n4523), .ZN(n7448) );
  NAND2_X1 U6134 ( .A1(n7535), .A2(n4317), .ZN(n7834) );
  AND2_X1 U6135 ( .A1(n9209), .A2(n4537), .ZN(n9161) );
  NAND2_X1 U6136 ( .A1(n7650), .A2(n4539), .ZN(n9317) );
  OAI21_X1 U6137 ( .B1(n8654), .B2(n4553), .A(n4550), .ZN(n4549) );
  NAND2_X1 U6138 ( .A1(n6412), .A2(n4305), .ZN(n4556) );
  INV_X1 U6139 ( .A(n9833), .ZN(n4560) );
  OAI21_X1 U6140 ( .B1(n8344), .B2(n4560), .A(n8193), .ZN(n7212) );
  NAND2_X1 U6141 ( .A1(n8189), .A2(n8193), .ZN(n8344) );
  NAND2_X1 U6142 ( .A1(n7294), .A2(n4562), .ZN(n4561) );
  OAI211_X1 U6143 ( .C1(n4311), .C2(n4565), .A(n4561), .B(n8232), .ZN(n7687)
         );
  NAND2_X1 U6144 ( .A1(n4567), .A2(n4386), .ZN(n6481) );
  NAND2_X1 U6145 ( .A1(n4574), .A2(n4575), .ZN(n8701) );
  INV_X2 U6146 ( .A(n4608), .ZN(n8317) );
  OAI21_X2 U6147 ( .B1(n5595), .B2(n6213), .A(n4586), .ZN(n9148) );
  NAND2_X1 U6148 ( .A1(n5595), .A2(n6288), .ZN(n9172) );
  NAND2_X1 U6149 ( .A1(n9172), .A2(n9173), .ZN(n9171) );
  NAND3_X1 U6150 ( .A1(n4816), .A2(n4817), .A3(n4591), .ZN(n4590) );
  NAND2_X1 U6151 ( .A1(n4590), .A2(n4963), .ZN(n5223) );
  NAND2_X1 U6152 ( .A1(n4590), .A2(n4587), .ZN(n4589) );
  NAND3_X1 U6153 ( .A1(n4816), .A2(n4817), .A3(n4958), .ZN(n5214) );
  OAI21_X2 U6154 ( .B1(n9280), .B2(n4595), .A(n4593), .ZN(n9245) );
  NAND4_X1 U6155 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n5670), .ZN(n5666)
         );
  NAND2_X1 U6156 ( .A1(n4608), .A2(n4607), .ZN(n6355) );
  NAND2_X1 U6157 ( .A1(n4609), .A2(n5759), .ZN(n9766) );
  NAND2_X1 U6158 ( .A1(n7191), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4609) );
  AOI21_X1 U6159 ( .B1(n5759), .B2(n4612), .A(n4611), .ZN(n4610) );
  INV_X1 U6160 ( .A(n9767), .ZN(n4611) );
  INV_X1 U6161 ( .A(n5759), .ZN(n4613) );
  NAND2_X1 U6162 ( .A1(n6640), .A2(n4615), .ZN(n4614) );
  INV_X1 U6163 ( .A(n4621), .ZN(n7771) );
  INV_X1 U6164 ( .A(n5749), .ZN(n4632) );
  NOR2_X1 U6165 ( .A1(n4632), .A2(n9672), .ZN(n4633) );
  NAND3_X1 U6166 ( .A1(n5700), .A2(n4362), .A3(n5699), .ZN(n4634) );
  NAND2_X1 U6167 ( .A1(n4636), .A2(n7017), .ZN(n6890) );
  NAND2_X1 U6168 ( .A1(n4637), .A2(n4361), .ZN(n7967) );
  INV_X1 U6169 ( .A(n4642), .ZN(n7727) );
  NAND2_X1 U6170 ( .A1(n4652), .A2(n4651), .ZN(n8687) );
  OAI22_X2 U6171 ( .A1(n7292), .A2(n6620), .B1(n7433), .B2(n7341), .ZN(n7431)
         );
  MUX2_X1 U6172 ( .A(n8908), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6173 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8908), .S(n6661), .Z(n6939) );
  NAND2_X1 U6174 ( .A1(n5159), .A2(n5160), .ZN(n4952) );
  NAND2_X2 U6175 ( .A1(n5251), .A2(n5250), .ZN(n7495) );
  NAND2_X1 U6176 ( .A1(n8243), .A2(n4658), .ZN(n4655) );
  NAND2_X1 U6177 ( .A1(n4655), .A2(n4656), .ZN(n8258) );
  NAND2_X1 U6178 ( .A1(n8192), .A2(n8310), .ZN(n8195) );
  NAND3_X1 U6179 ( .A1(n4664), .A2(n4663), .A3(n9838), .ZN(n8192) );
  OR2_X1 U6180 ( .A1(n8187), .A2(n8186), .ZN(n4663) );
  NAND2_X1 U6181 ( .A1(n8188), .A2(n8310), .ZN(n4664) );
  OAI21_X1 U6182 ( .B1(n4677), .B2(n8205), .A(n4349), .ZN(n8242) );
  NAND3_X1 U6183 ( .A1(n5631), .A2(n5664), .A3(n4895), .ZN(n5637) );
  NAND4_X1 U6184 ( .A1(n5631), .A2(n5663), .A3(n4895), .A4(n4357), .ZN(n5639)
         );
  NAND3_X1 U6185 ( .A1(n4682), .A2(n8638), .A3(n4681), .ZN(n4680) );
  NAND3_X1 U6186 ( .A1(n8291), .A2(n8335), .A3(n8326), .ZN(n4681) );
  NAND2_X1 U6187 ( .A1(n5657), .A2(n4684), .ZN(n6325) );
  MUX2_X1 U6188 ( .A(n4698), .B(P1_REG2_REG_1__SCAN_IN), .S(n9477), .Z(n9474)
         );
  OR2_X2 U6189 ( .A1(n7562), .A2(n4700), .ZN(n9520) );
  NAND2_X1 U6190 ( .A1(n4701), .A2(n4702), .ZN(n6129) );
  NAND2_X1 U6191 ( .A1(n6123), .A2(n4703), .ZN(n4701) );
  NAND2_X1 U6192 ( .A1(n7090), .A2(n4711), .ZN(n4708) );
  AOI21_X1 U6193 ( .B1(n7090), .B2(n5582), .A(n4713), .ZN(n4710) );
  NAND2_X1 U6194 ( .A1(n6194), .A2(n9535), .ZN(n9534) );
  NAND2_X1 U6195 ( .A1(n5708), .A2(n7008), .ZN(n7010) );
  NAND2_X1 U6196 ( .A1(n7010), .A2(n4738), .ZN(n4739) );
  NAND2_X1 U6197 ( .A1(n4743), .A2(n9752), .ZN(n4741) );
  OR2_X1 U6198 ( .A1(n5619), .A2(n5620), .ZN(P1_U3551) );
  NAND2_X1 U6199 ( .A1(n4750), .A2(n4753), .ZN(n7375) );
  NAND2_X1 U6200 ( .A1(n7491), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U6201 ( .A1(n4757), .A2(n4358), .ZN(n5534) );
  NAND2_X1 U6202 ( .A1(n5493), .A2(n4761), .ZN(n4757) );
  INV_X1 U6203 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4782) );
  INV_X1 U6204 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4783) );
  INV_X1 U6205 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4781) );
  INV_X1 U6206 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4780) );
  NAND3_X1 U6207 ( .A1(n4783), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4778) );
  NAND3_X1 U6208 ( .A1(n4782), .A2(n4781), .A3(n4780), .ZN(n4779) );
  NAND2_X1 U6209 ( .A1(n7310), .A2(n4786), .ZN(n5188) );
  NAND3_X1 U6210 ( .A1(n8277), .A2(n8173), .A3(n8684), .ZN(n4795) );
  NAND3_X1 U6211 ( .A1(n8684), .A2(n8310), .A3(n8278), .ZN(n4788) );
  NAND2_X1 U6212 ( .A1(n4790), .A2(n4789), .ZN(n8281) );
  NAND3_X1 U6213 ( .A1(n4792), .A2(n4794), .A3(n4791), .ZN(n4790) );
  AOI21_X1 U6214 ( .B1(n5411), .B2(n4810), .A(n4808), .ZN(n4799) );
  OAI21_X1 U6215 ( .B1(n5411), .B2(n5011), .A(n5010), .ZN(n5419) );
  NAND2_X1 U6216 ( .A1(n5223), .A2(n5222), .ZN(n5225) );
  NAND3_X1 U6217 ( .A1(n4300), .A2(n4952), .A3(n4312), .ZN(n4817) );
  NAND2_X1 U6218 ( .A1(n4300), .A2(n4955), .ZN(n4818) );
  NAND2_X1 U6219 ( .A1(n5182), .A2(n5183), .ZN(n4819) );
  NAND2_X1 U6220 ( .A1(n5277), .A2(n4827), .ZN(n4824) );
  NAND2_X1 U6221 ( .A1(n5277), .A2(n4979), .ZN(n5292) );
  NAND2_X1 U6222 ( .A1(n5001), .A2(n5000), .ZN(n5383) );
  NAND2_X1 U6223 ( .A1(n7124), .A2(n4830), .ZN(n4835) );
  NAND2_X1 U6224 ( .A1(n7125), .A2(n4836), .ZN(n4834) );
  INV_X1 U6225 ( .A(n5894), .ZN(n4837) );
  NOR2_X1 U6226 ( .A1(n7125), .A2(n7166), .ZN(n4841) );
  NOR2_X2 U6227 ( .A1(n5243), .A2(n4842), .ZN(n5061) );
  NAND4_X1 U6228 ( .A1(n4917), .A2(n4918), .A3(n4916), .A4(n4915), .ZN(n4842)
         );
  NAND2_X1 U6229 ( .A1(n4843), .A2(n4845), .ZN(n7941) );
  NAND2_X1 U6230 ( .A1(n8909), .A2(n4385), .ZN(n4851) );
  NAND2_X1 U6231 ( .A1(n8949), .A2(n5980), .ZN(n8980) );
  OR2_X1 U6232 ( .A1(n8981), .A2(n4862), .ZN(n4861) );
  AND2_X2 U6233 ( .A1(n5119), .A2(n8109), .ZN(n5168) );
  OAI22_X1 U6234 ( .A1(n5119), .A2(P1_U3086), .B1(n9450), .B2(n6183), .ZN(
        n4865) );
  NAND2_X1 U6235 ( .A1(n6706), .A2(n4867), .ZN(n4866) );
  OAI211_X1 U6236 ( .C1(n6706), .C2(n4868), .A(n4866), .B(n6713), .ZN(P1_U3214) );
  NAND2_X1 U6237 ( .A1(n6706), .A2(n4380), .ZN(n6705) );
  NAND2_X1 U6238 ( .A1(n4926), .A2(n4870), .ZN(n5115) );
  INV_X1 U6239 ( .A(n5115), .ZN(n5113) );
  NAND3_X1 U6240 ( .A1(n5838), .A2(n5837), .A3(n6050), .ZN(n5843) );
  NAND4_X1 U6241 ( .A1(n5628), .A2(n5627), .A3(n5710), .A4(n4872), .ZN(n4874)
         );
  OR2_X1 U6242 ( .A1(n6661), .A2(n9682), .ZN(n4875) );
  NAND2_X1 U6243 ( .A1(n8124), .A2(n4877), .ZN(n8441) );
  OAI21_X2 U6244 ( .B1(n7336), .B2(n4880), .A(n4879), .ZN(n7759) );
  NAND2_X1 U6245 ( .A1(n7764), .A2(n7787), .ZN(n4887) );
  NAND2_X1 U6246 ( .A1(n4887), .A2(n4888), .ZN(n7799) );
  NAND2_X1 U6247 ( .A1(n8483), .A2(n8148), .ZN(n4890) );
  NAND2_X1 U6248 ( .A1(n4890), .A2(n8149), .ZN(n4891) );
  NAND3_X1 U6249 ( .A1(n4891), .A2(n4892), .A3(n8487), .ZN(n8400) );
  NAND2_X1 U6250 ( .A1(n8346), .A2(n7137), .ZN(n7136) );
  OAI21_X1 U6251 ( .B1(n8181), .B2(n8346), .A(n8183), .ZN(n9833) );
  NAND2_X1 U6252 ( .A1(n9150), .A2(n9149), .ZN(n9151) );
  INV_X1 U6253 ( .A(n6198), .ZN(n7089) );
  NAND2_X1 U6254 ( .A1(n6325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U6255 ( .A1(n4910), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6256 ( .A1(n5083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6257 ( .A1(n5055), .A2(SI_29_), .ZN(n6080) );
  OR2_X1 U6258 ( .A1(n5055), .A2(SI_29_), .ZN(n5056) );
  OAI211_X4 U6259 ( .C1(n5184), .C2(n4935), .A(n5130), .B(n5129), .ZN(n9549)
         );
  AND2_X1 U6260 ( .A1(n9145), .A2(n9142), .ZN(n5614) );
  OAI211_X1 U6261 ( .C1(n8578), .C2(n9832), .A(n6664), .B(n6663), .ZN(n8577)
         );
  XNOR2_X1 U6262 ( .A(n6078), .B(n6076), .ZN(n5055) );
  INV_X1 U6263 ( .A(n8318), .ZN(n6655) );
  NAND2_X1 U6264 ( .A1(n8318), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6345) );
  OR2_X1 U6265 ( .A1(n8198), .A2(n8197), .ZN(n8220) );
  NAND2_X1 U6266 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5658) );
  AND2_X1 U6267 ( .A1(n7051), .A2(n9834), .ZN(n8586) );
  AND2_X1 U6268 ( .A1(n6346), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4897) );
  AND2_X1 U6269 ( .A1(n6135), .A2(n6095), .ZN(n4898) );
  NOR2_X1 U6270 ( .A1(n9650), .A2(n5623), .ZN(n4899) );
  OR2_X1 U6271 ( .A1(n8582), .A2(n8822), .ZN(n4900) );
  AND2_X1 U6272 ( .A1(n5996), .A2(n5995), .ZN(n4901) );
  AND2_X1 U6273 ( .A1(n6071), .A2(n9007), .ZN(n4902) );
  OR2_X1 U6274 ( .A1(n8582), .A2(n7307), .ZN(n4903) );
  AND2_X2 U6275 ( .A1(n7314), .A2(n9294), .ZN(n9543) );
  INV_X1 U6276 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4935) );
  AND2_X1 U6277 ( .A1(n9650), .A2(n9641), .ZN(n9428) );
  INV_X1 U6278 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5632) );
  INV_X1 U6279 ( .A(n9840), .ZN(n8747) );
  AND2_X1 U6280 ( .A1(n6927), .A2(n8326), .ZN(n9840) );
  NAND2_X1 U6281 ( .A1(n6148), .A2(n6143), .ZN(n4904) );
  OR2_X1 U6282 ( .A1(n9437), .A2(n8918), .ZN(n4905) );
  INV_X1 U6283 ( .A(n5106), .ZN(n5109) );
  AND2_X1 U6284 ( .A1(n9889), .A2(n8527), .ZN(n4906) );
  NOR2_X1 U6285 ( .A1(n8837), .A2(n8656), .ZN(n4907) );
  AND3_X1 U6286 ( .A1(n8206), .A2(n8310), .A3(n8225), .ZN(n4908) );
  INV_X1 U6287 ( .A(n8358), .ZN(n6626) );
  OAI22_X1 U6288 ( .A1(n6194), .A2(n9536), .B1(n9549), .B2(n5844), .ZN(n7565)
         );
  XNOR2_X1 U6289 ( .A(n5850), .B(n5851), .ZN(n6953) );
  INV_X1 U6290 ( .A(n7059), .ZN(n5876) );
  OR2_X1 U6291 ( .A1(n8530), .A2(n7271), .ZN(n4909) );
  XNOR2_X1 U6292 ( .A(n5883), .B(n6034), .ZN(n5888) );
  OAI21_X1 U6293 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8196) );
  OAI211_X1 U6294 ( .C1(n8220), .C2(n8201), .A(n8200), .B(n8221), .ZN(n8202)
         );
  INV_X1 U6295 ( .A(n6307), .ZN(n6096) );
  NAND2_X1 U6296 ( .A1(n6097), .A2(n6096), .ZN(n6105) );
  AOI21_X1 U6297 ( .B1(n6120), .B2(n6112), .A(n6260), .ZN(n6116) );
  NOR2_X1 U6298 ( .A1(n7643), .A2(n6130), .ZN(n6133) );
  INV_X1 U6299 ( .A(n6280), .ZN(n6118) );
  NAND2_X1 U6300 ( .A1(n8269), .A2(n8310), .ZN(n8270) );
  NAND2_X1 U6301 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  INV_X1 U6302 ( .A(n7566), .ZN(n6195) );
  INV_X1 U6303 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5629) );
  INV_X1 U6304 ( .A(n8619), .ZN(n6648) );
  INV_X1 U6305 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U6306 ( .A1(n8770), .A2(n6648), .ZN(n6649) );
  NAND2_X1 U6307 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  INV_X1 U6308 ( .A(n8526), .ZN(n7789) );
  INV_X1 U6309 ( .A(n9377), .ZN(n5612) );
  AND2_X1 U6310 ( .A1(n5346), .A2(n4987), .ZN(n4995) );
  XNOR2_X1 U6311 ( .A(n7224), .B(n7112), .ZN(n7106) );
  NAND2_X1 U6312 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  XNOR2_X1 U6313 ( .A(n5731), .B(n6400), .ZN(n7582) );
  INV_X1 U6314 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5665) );
  INV_X1 U6315 ( .A(n5484), .ZN(n5482) );
  INV_X1 U6316 ( .A(n9261), .ZN(n5461) );
  OR2_X1 U6317 ( .A1(n6736), .A2(n5143), .ZN(n5186) );
  INV_X1 U6318 ( .A(n9161), .ZN(n9177) );
  INV_X1 U6319 ( .A(n5855), .ZN(n5150) );
  NOR2_X1 U6320 ( .A1(n6385), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6405) );
  AND2_X1 U6321 ( .A1(n7869), .A2(n7791), .ZN(n7792) );
  INV_X1 U6322 ( .A(n8476), .ZN(n8140) );
  INV_X1 U6323 ( .A(n8512), .ZN(n8496) );
  NOR2_X1 U6324 ( .A1(n5734), .A2(n8068), .ZN(n8024) );
  NOR2_X1 U6325 ( .A1(n6571), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6582) );
  AND2_X1 U6326 ( .A1(n6493), .A2(n6492), .ZN(n6504) );
  INV_X1 U6327 ( .A(n8355), .ZN(n6411) );
  OR2_X1 U6328 ( .A1(n6729), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6669) );
  INV_X1 U6329 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5670) );
  INV_X1 U6330 ( .A(n5977), .ZN(n5978) );
  OR2_X1 U6331 ( .A1(n5528), .A2(n8997), .ZN(n5540) );
  NAND2_X1 U6332 ( .A1(n5482), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5503) );
  OR2_X1 U6333 ( .A1(n5516), .A2(n8935), .ZN(n5528) );
  NAND2_X1 U6334 ( .A1(n5390), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5404) );
  INV_X1 U6335 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5623) );
  INV_X1 U6336 ( .A(n6092), .ZN(n6132) );
  INV_X1 U6337 ( .A(n7684), .ZN(n5598) );
  AOI21_X1 U6338 ( .B1(n5548), .B2(n5054), .A(n5053), .ZN(n6078) );
  OAI21_X1 U6339 ( .B1(n5464), .B2(n5463), .A(n5026), .ZN(n5478) );
  INV_X1 U6340 ( .A(SI_16_), .ZN(n5380) );
  INV_X1 U6341 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6342 ( .A1(n6435), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6443) );
  OR2_X1 U6343 ( .A1(n6994), .A2(n6993), .ZN(n8499) );
  INV_X1 U6344 ( .A(n8573), .ZN(n8579) );
  OR2_X1 U6345 ( .A1(n6561), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6571) );
  OR2_X1 U6346 ( .A1(n6515), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6525) );
  OR2_X1 U6347 ( .A1(n6465), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6475) );
  OR2_X1 U6348 ( .A1(n6427), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6435) );
  OR2_X1 U6349 ( .A1(n8310), .A2(n6988), .ZN(n7042) );
  INV_X1 U6350 ( .A(n6987), .ZN(n7046) );
  NAND2_X1 U6351 ( .A1(n7908), .A2(n8359), .ZN(n7955) );
  NAND2_X1 U6352 ( .A1(n6993), .A2(n8326), .ZN(n8745) );
  AND2_X1 U6353 ( .A1(n6947), .A2(n6686), .ZN(n6931) );
  INV_X1 U6354 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5634) );
  OR2_X1 U6355 ( .A1(n5683), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U6356 ( .A1(n5964), .A2(n5966), .ZN(n5967) );
  OR2_X1 U6357 ( .A1(n5437), .A2(n10064), .ZN(n5453) );
  OR2_X1 U6358 ( .A1(n5299), .A2(n7858), .ZN(n5321) );
  AND2_X1 U6359 ( .A1(n5540), .A2(n5529), .ZN(n9193) );
  OR2_X1 U6360 ( .A1(n5404), .A2(n5403), .ZN(n5426) );
  INV_X1 U6361 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6977) );
  INV_X1 U6362 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U6363 ( .A1(n9160), .A2(n9159), .ZN(n9336) );
  INV_X1 U6364 ( .A(n6213), .ZN(n9173) );
  OR2_X1 U6365 ( .A1(n9442), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5110) );
  AND2_X1 U6366 ( .A1(n6095), .A2(n6132), .ZN(n7833) );
  OR2_X1 U6367 ( .A1(n6842), .A2(n5598), .ZN(n9620) );
  OR2_X1 U6368 ( .A1(n6307), .A2(n5598), .ZN(n9644) );
  AND2_X1 U6369 ( .A1(n5044), .A2(n5043), .ZN(n5525) );
  INV_X1 U6370 ( .A(n8499), .ZN(n8510) );
  INV_X1 U6371 ( .A(n8503), .ZN(n8508) );
  AND2_X1 U6372 ( .A1(n6599), .A2(n6598), .ZN(n8619) );
  AND4_X1 U6373 ( .A1(n6510), .A2(n6509), .A3(n6508), .A4(n6507), .ZN(n8479)
         );
  INV_X1 U6374 ( .A(n9817), .ZN(n9768) );
  INV_X1 U6375 ( .A(n9737), .ZN(n9808) );
  AOI21_X1 U6376 ( .B1(n5830), .B2(n9822), .A(n5829), .ZN(n5831) );
  OR2_X1 U6377 ( .A1(n6946), .A2(n6937), .ZN(n9834) );
  INV_X2 U6378 ( .A(n8586), .ZN(n8752) );
  AND2_X1 U6379 ( .A1(n9904), .A2(n9865), .ZN(n8809) );
  INV_X1 U6380 ( .A(n7307), .ZN(n8808) );
  AND2_X1 U6381 ( .A1(n8336), .A2(n8335), .ZN(n8655) );
  INV_X1 U6382 ( .A(n8884), .ZN(n8890) );
  AND2_X1 U6383 ( .A1(n7879), .A2(n8328), .ZN(n9890) );
  NAND2_X1 U6384 ( .A1(n9832), .A2(n9885), .ZN(n9865) );
  AND2_X1 U6385 ( .A1(n5677), .A2(n5676), .ZN(n6471) );
  OAI21_X1 U6386 ( .B1(n9409), .B2(n9017), .A(n6711), .ZN(n6712) );
  INV_X1 U6387 ( .A(n9017), .ZN(n8968) );
  OR2_X1 U6388 ( .A1(n9179), .A2(n5563), .ZN(n5546) );
  INV_X1 U6389 ( .A(n5469), .ZN(n5563) );
  INV_X1 U6390 ( .A(n5605), .ZN(n6869) );
  NAND2_X1 U6391 ( .A1(n6772), .A2(n6771), .ZN(n9486) );
  INV_X1 U6392 ( .A(n9486), .ZN(n9116) );
  INV_X1 U6393 ( .A(n9325), .ZN(n9531) );
  INV_X1 U6394 ( .A(n9543), .ZN(n9322) );
  AND2_X1 U6395 ( .A1(n10083), .A2(n9641), .ZN(n9373) );
  AND2_X1 U6396 ( .A1(n5110), .A2(n9444), .ZN(n6044) );
  INV_X1 U6397 ( .A(n6044), .ZN(n7313) );
  XNOR2_X1 U6398 ( .A(n5102), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6741) );
  INV_X1 U6399 ( .A(n9452), .ZN(n7895) );
  OR2_X1 U6400 ( .A1(n6994), .A2(n6927), .ZN(n8512) );
  AND2_X1 U6401 ( .A1(n6933), .A2(n6932), .ZN(n8503) );
  AND2_X1 U6402 ( .A1(n8323), .A2(n6608), .ZN(n8600) );
  INV_X1 U6403 ( .A(n8468), .ZN(n8656) );
  INV_X1 U6404 ( .A(n8746), .ZN(n8722) );
  INV_X1 U6405 ( .A(n9822), .ZN(n9763) );
  INV_X1 U6406 ( .A(n9809), .ZN(n9807) );
  NAND2_X1 U6407 ( .A1(n7053), .A2(n7052), .ZN(n8581) );
  INV_X1 U6408 ( .A(n8809), .ZN(n8806) );
  INV_X1 U6409 ( .A(n9904), .ZN(n9902) );
  OR2_X1 U6410 ( .A1(n9893), .A2(n9879), .ZN(n8884) );
  AND2_X1 U6411 ( .A1(n6689), .A2(n6688), .ZN(n9893) );
  AND2_X1 U6412 ( .A1(n6729), .A2(n6950), .ZN(n6753) );
  INV_X1 U6413 ( .A(n6753), .ZN(n6751) );
  INV_X1 U6414 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8085) );
  INV_X1 U6415 ( .A(n7899), .ZN(n8906) );
  NAND2_X1 U6416 ( .A1(n6072), .A2(n4902), .ZN(n6073) );
  INV_X1 U6417 ( .A(n9007), .ZN(n8988) );
  NAND2_X1 U6418 ( .A1(n5510), .A2(n5509), .ZN(n9026) );
  INV_X1 U6419 ( .A(n9478), .ZN(n9498) );
  OR2_X1 U6420 ( .A1(n9543), .A2(n9119), .ZN(n9272) );
  INV_X1 U6421 ( .A(n9322), .ZN(n9268) );
  INV_X1 U6422 ( .A(n9373), .ZN(n9395) );
  INV_X1 U6423 ( .A(n10083), .ZN(n9670) );
  INV_X1 U6424 ( .A(n9178), .ZN(n9409) );
  INV_X1 U6425 ( .A(n6008), .ZN(n9424) );
  INV_X1 U6426 ( .A(n9650), .ZN(n9648) );
  INV_X1 U6427 ( .A(n9558), .ZN(n9559) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7898) );
  INV_X1 U6429 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7561) );
  INV_X1 U6430 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6819) );
  INV_X1 U6431 ( .A(n9447), .ZN(n9450) );
  AND2_X1 U6432 ( .A1(n6716), .A2(n6715), .ZN(P1_U3973) );
  NOR2_X1 U6433 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4918) );
  NOR2_X1 U6434 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4917) );
  NOR2_X1 U6435 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4916) );
  NAND4_X1 U6436 ( .A1(n5064), .A2(n4919), .A3(n5084), .A4(n5086), .ZN(n4921)
         );
  NAND4_X1 U6437 ( .A1(n5081), .A2(n5088), .A3(n5063), .A4(n5066), .ZN(n4920)
         );
  NOR2_X1 U6438 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  NAND2_X1 U6439 ( .A1(n4924), .A2(n4923), .ZN(n5060) );
  OAI21_X1 U6440 ( .B1(n4927), .B2(n5176), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n4930) );
  NAND2_X1 U6441 ( .A1(n4930), .A2(n4929), .ZN(n4931) );
  NAND2_X1 U6442 ( .A1(n4932), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U6443 ( .A1(n4937), .A2(n4936), .ZN(n4941) );
  INV_X1 U6444 ( .A(n5127), .ZN(n4940) );
  AND2_X1 U6445 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U6446 ( .A1(n6717), .A2(n4938), .ZN(n5137) );
  NAND3_X1 U6447 ( .A1(n6722), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4939) );
  NAND2_X1 U6448 ( .A1(n4940), .A2(n5126), .ZN(n4943) );
  NAND2_X1 U6449 ( .A1(n4941), .A2(SI_1_), .ZN(n4942) );
  NAND2_X1 U6450 ( .A1(n4943), .A2(n4942), .ZN(n5141) );
  INV_X1 U6451 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6725) );
  INV_X1 U6452 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6721) );
  MUX2_X1 U6453 ( .A(n6725), .B(n6721), .S(n6717), .Z(n4944) );
  NAND2_X1 U6454 ( .A1(n5141), .A2(n5142), .ZN(n4947) );
  INV_X1 U6455 ( .A(n4944), .ZN(n4945) );
  NAND2_X1 U6456 ( .A1(n4945), .A2(SI_2_), .ZN(n4946) );
  NAND2_X1 U6457 ( .A1(n4947), .A2(n4946), .ZN(n5159) );
  INV_X1 U6458 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6730) );
  INV_X1 U6459 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6718) );
  XNOR2_X1 U6460 ( .A(n4949), .B(SI_3_), .ZN(n5160) );
  INV_X1 U6461 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6462 ( .A1(n4950), .A2(SI_3_), .ZN(n4951) );
  INV_X1 U6463 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6735) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6719) );
  MUX2_X1 U6465 ( .A(n6735), .B(n6719), .S(n6717), .Z(n4953) );
  XNOR2_X1 U6466 ( .A(n4953), .B(SI_4_), .ZN(n5183) );
  INV_X1 U6467 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6468 ( .A1(n4954), .A2(SI_4_), .ZN(n4955) );
  INV_X1 U6469 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6732) );
  INV_X1 U6470 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4956) );
  MUX2_X1 U6471 ( .A(n6732), .B(n4956), .S(n6717), .Z(n5197) );
  INV_X1 U6472 ( .A(SI_5_), .ZN(n4957) );
  NAND2_X1 U6473 ( .A1(n5197), .A2(n4957), .ZN(n4958) );
  MUX2_X1 U6474 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6717), .Z(n4959) );
  NAND2_X1 U6475 ( .A1(n4959), .A2(SI_6_), .ZN(n4963) );
  INV_X1 U6476 ( .A(n4959), .ZN(n4961) );
  INV_X1 U6477 ( .A(SI_6_), .ZN(n4960) );
  NAND2_X1 U6478 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  NAND2_X1 U6479 ( .A1(n4963), .A2(n4962), .ZN(n5212) );
  MUX2_X1 U6480 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6717), .Z(n4964) );
  INV_X1 U6481 ( .A(n4964), .ZN(n4966) );
  INV_X1 U6482 ( .A(SI_7_), .ZN(n4965) );
  NAND2_X1 U6483 ( .A1(n4966), .A2(n4965), .ZN(n4967) );
  MUX2_X1 U6484 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6717), .Z(n4969) );
  XNOR2_X1 U6485 ( .A(n4969), .B(SI_8_), .ZN(n5241) );
  INV_X1 U6486 ( .A(n4969), .ZN(n4971) );
  INV_X1 U6487 ( .A(SI_8_), .ZN(n4970) );
  MUX2_X1 U6488 ( .A(n6817), .B(n6819), .S(n6717), .Z(n4972) );
  XNOR2_X1 U6489 ( .A(n4972), .B(SI_9_), .ZN(n5262) );
  INV_X1 U6490 ( .A(n4972), .ZN(n4973) );
  MUX2_X1 U6491 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6717), .Z(n4974) );
  NAND2_X1 U6492 ( .A1(n4974), .A2(SI_10_), .ZN(n4979) );
  INV_X1 U6493 ( .A(n4974), .ZN(n4976) );
  INV_X1 U6494 ( .A(SI_10_), .ZN(n4975) );
  NAND2_X1 U6495 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  NAND2_X1 U6496 ( .A1(n4979), .A2(n4977), .ZN(n5275) );
  INV_X1 U6497 ( .A(n5275), .ZN(n4978) );
  MUX2_X1 U6498 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6717), .Z(n4980) );
  XNOR2_X1 U6499 ( .A(n4980), .B(SI_11_), .ZN(n5291) );
  MUX2_X1 U6500 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6717), .Z(n4981) );
  NAND2_X1 U6501 ( .A1(n4981), .A2(SI_12_), .ZN(n4982) );
  OAI21_X1 U6502 ( .B1(n4981), .B2(SI_12_), .A(n4982), .ZN(n5308) );
  MUX2_X1 U6503 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6717), .Z(n4983) );
  NAND2_X1 U6504 ( .A1(n4983), .A2(SI_13_), .ZN(n5346) );
  OAI21_X1 U6505 ( .B1(n4983), .B2(SI_13_), .A(n5346), .ZN(n5331) );
  INV_X1 U6506 ( .A(n5331), .ZN(n4993) );
  MUX2_X1 U6507 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6717), .Z(n5347) );
  INV_X1 U6508 ( .A(n5347), .ZN(n4985) );
  AND2_X1 U6509 ( .A1(n4993), .A2(n4997), .ZN(n4986) );
  INV_X1 U6510 ( .A(n4997), .ZN(n4988) );
  NAND2_X1 U6511 ( .A1(n5347), .A2(SI_14_), .ZN(n4987) );
  NAND2_X1 U6512 ( .A1(n4990), .A2(n4989), .ZN(n5362) );
  NAND2_X1 U6513 ( .A1(n5362), .A2(SI_15_), .ZN(n4992) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6717), .Z(n5363) );
  INV_X1 U6515 ( .A(n5363), .ZN(n4991) );
  NAND2_X1 U6516 ( .A1(n4992), .A2(n4991), .ZN(n5001) );
  INV_X1 U6517 ( .A(SI_15_), .ZN(n4994) );
  NAND2_X1 U6518 ( .A1(n5333), .A2(n4996), .ZN(n4999) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6717), .Z(n5381) );
  MUX2_X1 U6520 ( .A(n7289), .B(n7288), .S(n6717), .Z(n5003) );
  NAND2_X1 U6521 ( .A1(n5003), .A2(n5002), .ZN(n5006) );
  INV_X1 U6522 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6523 ( .A1(n5004), .A2(SI_17_), .ZN(n5005) );
  NAND2_X1 U6524 ( .A1(n5006), .A2(n5005), .ZN(n5398) );
  MUX2_X1 U6525 ( .A(n7349), .B(n5007), .S(n6717), .Z(n5008) );
  XNOR2_X1 U6526 ( .A(n5008), .B(SI_18_), .ZN(n5410) );
  INV_X1 U6527 ( .A(n5410), .ZN(n5011) );
  INV_X1 U6528 ( .A(n5008), .ZN(n5009) );
  NAND2_X1 U6529 ( .A1(n5009), .A2(SI_18_), .ZN(n5010) );
  MUX2_X1 U6530 ( .A(n7558), .B(n7561), .S(n6717), .Z(n5013) );
  INV_X1 U6531 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6532 ( .A1(n5014), .A2(SI_19_), .ZN(n5015) );
  NAND2_X1 U6533 ( .A1(n5018), .A2(n5015), .ZN(n5418) );
  MUX2_X1 U6534 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6717), .Z(n5432) );
  INV_X1 U6535 ( .A(n5432), .ZN(n5016) );
  MUX2_X1 U6536 ( .A(n10021), .B(n7721), .S(n6717), .Z(n5446) );
  NOR2_X1 U6537 ( .A1(n5019), .A2(SI_21_), .ZN(n5021) );
  NAND2_X1 U6538 ( .A1(n5019), .A2(SI_21_), .ZN(n5020) );
  OAI21_X1 U6539 ( .B1(n5448), .B2(n5021), .A(n5020), .ZN(n5464) );
  MUX2_X1 U6540 ( .A(n7878), .B(n7882), .S(n6717), .Z(n5023) );
  INV_X1 U6541 ( .A(SI_22_), .ZN(n5022) );
  NAND2_X1 U6542 ( .A1(n5023), .A2(n5022), .ZN(n5026) );
  INV_X1 U6543 ( .A(n5023), .ZN(n5024) );
  NAND2_X1 U6544 ( .A1(n5024), .A2(SI_22_), .ZN(n5025) );
  NAND2_X1 U6545 ( .A1(n5026), .A2(n5025), .ZN(n5463) );
  MUX2_X1 U6546 ( .A(n7902), .B(n7898), .S(n6717), .Z(n5028) );
  INV_X1 U6547 ( .A(SI_23_), .ZN(n5027) );
  NAND2_X1 U6548 ( .A1(n5028), .A2(n5027), .ZN(n5494) );
  INV_X1 U6549 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6550 ( .A1(n5029), .A2(SI_23_), .ZN(n5030) );
  NAND2_X1 U6551 ( .A1(n5478), .A2(n5477), .ZN(n5476) );
  MUX2_X1 U6552 ( .A(n9961), .B(n7980), .S(n6717), .Z(n5032) );
  INV_X1 U6553 ( .A(SI_24_), .ZN(n5031) );
  NAND2_X1 U6554 ( .A1(n5032), .A2(n5031), .ZN(n5496) );
  AND2_X1 U6555 ( .A1(n5494), .A2(n5496), .ZN(n5035) );
  INV_X1 U6556 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6557 ( .A1(n5033), .A2(SI_24_), .ZN(n5495) );
  INV_X1 U6558 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8115) );
  INV_X1 U6559 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7991) );
  MUX2_X1 U6560 ( .A(n8115), .B(n7991), .S(n6717), .Z(n5036) );
  INV_X1 U6561 ( .A(SI_25_), .ZN(n10049) );
  NAND2_X1 U6562 ( .A1(n5036), .A2(n10049), .ZN(n5039) );
  INV_X1 U6563 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6564 ( .A1(n5037), .A2(SI_25_), .ZN(n5038) );
  MUX2_X1 U6565 ( .A(n8085), .B(n9959), .S(n6717), .Z(n5041) );
  INV_X1 U6566 ( .A(SI_26_), .ZN(n5040) );
  NAND2_X1 U6567 ( .A1(n5041), .A2(n5040), .ZN(n5044) );
  INV_X1 U6568 ( .A(n5041), .ZN(n5042) );
  NAND2_X1 U6569 ( .A1(n5042), .A2(SI_26_), .ZN(n5043) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6578) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8107) );
  MUX2_X1 U6572 ( .A(n6578), .B(n8107), .S(n6717), .Z(n5047) );
  INV_X1 U6573 ( .A(SI_27_), .ZN(n5046) );
  NAND2_X1 U6574 ( .A1(n5047), .A2(n5046), .ZN(n5547) );
  INV_X1 U6575 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6576 ( .A1(n5048), .A2(SI_27_), .ZN(n5049) );
  INV_X1 U6577 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6590) );
  INV_X1 U6578 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8114) );
  MUX2_X1 U6579 ( .A(n6590), .B(n8114), .S(n6717), .Z(n5051) );
  INV_X1 U6580 ( .A(SI_28_), .ZN(n5050) );
  NAND2_X1 U6581 ( .A1(n5051), .A2(n5050), .ZN(n5550) );
  AND2_X1 U6582 ( .A1(n5547), .A2(n5550), .ZN(n5054) );
  INV_X1 U6583 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6584 ( .A1(n5052), .A2(SI_28_), .ZN(n5549) );
  MUX2_X1 U6585 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6717), .Z(n6076) );
  INV_X1 U6586 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8110) );
  OR2_X1 U6587 ( .A1(n5184), .A2(n8110), .ZN(n5057) );
  AND2_X1 U6588 ( .A1(n5058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6589 ( .A1(n7992), .A2(P1_B_REG_SCAN_IN), .ZN(n5068) );
  NAND3_X1 U6590 ( .A1(n5084), .A2(n5086), .A3(n5088), .ZN(n5062) );
  INV_X1 U6591 ( .A(n5064), .ZN(n5065) );
  MUX2_X1 U6592 ( .A(n5068), .B(P1_B_REG_SCAN_IN), .S(n5109), .Z(n5071) );
  NAND2_X1 U6593 ( .A1(n5069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5070) );
  OR2_X1 U6594 ( .A1(n9442), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6595 ( .A1(n7992), .A2(n8088), .ZN(n9443) );
  INV_X1 U6596 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6597 ( .A1(n5400), .A2(n5084), .ZN(n5085) );
  NAND2_X1 U6598 ( .A1(n5412), .A2(n5086), .ZN(n5087) );
  NOR2_X1 U6599 ( .A1(n7311), .A2(n6061), .ZN(n5108) );
  NOR2_X1 U6600 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .ZN(
        n5093) );
  NOR4_X1 U6601 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5092) );
  NOR4_X1 U6602 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5091) );
  NOR4_X1 U6603 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5090) );
  NAND4_X1 U6604 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), .ZN(n5099)
         );
  NOR4_X1 U6605 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5097) );
  NOR4_X1 U6606 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5096) );
  NOR4_X1 U6607 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5095) );
  NOR4_X1 U6608 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5094) );
  NAND4_X1 U6609 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n5098)
         );
  NOR2_X1 U6610 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  OR2_X1 U6611 ( .A1(n9442), .A2(n5100), .ZN(n6043) );
  NAND2_X1 U6612 ( .A1(n6316), .A2(n5572), .ZN(n6742) );
  NAND2_X1 U6613 ( .A1(n5833), .A2(n7684), .ZN(n6305) );
  INV_X1 U6614 ( .A(n6305), .ZN(n5111) );
  NAND2_X1 U6615 ( .A1(n5101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5102) );
  INV_X1 U6616 ( .A(n6741), .ZN(n6715) );
  OAI211_X1 U6617 ( .C1(n6742), .C2(n5111), .A(n6715), .B(n6714), .ZN(n6062)
         );
  NOR2_X1 U6618 ( .A1(n6062), .A2(P1_U3086), .ZN(n5107) );
  NAND2_X1 U6619 ( .A1(n5106), .A2(n8088), .ZN(n9444) );
  INV_X1 U6620 ( .A(n9632), .ZN(n9641) );
  INV_X1 U6621 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6622 ( .A1(n5113), .A2(n5112), .ZN(n5117) );
  NAND2_X1 U6623 ( .A1(n5115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6624 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5116), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5118) );
  NAND2_X1 U6625 ( .A1(n5192), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6626 ( .A1(n4287), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5124) );
  INV_X1 U6627 ( .A(n5119), .ZN(n5121) );
  AND2_X4 U6628 ( .A1(n5121), .A2(n5120), .ZN(n5469) );
  NAND2_X1 U6629 ( .A1(n5469), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6630 ( .A1(n4910), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6631 ( .A1(n4292), .A2(n4327), .ZN(n5130) );
  XNOR2_X2 U6632 ( .A(n5844), .B(n9549), .ZN(n6194) );
  NAND2_X1 U6633 ( .A1(n5469), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6634 ( .A1(n5192), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6635 ( .A1(n4287), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5131) );
  INV_X1 U6636 ( .A(SI_0_), .ZN(n5136) );
  INV_X1 U6637 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5135) );
  OAI21_X1 U6638 ( .B1(n6722), .B2(n5136), .A(n5135), .ZN(n5138) );
  AND2_X1 U6639 ( .A1(n5138), .A2(n5137), .ZN(n9453) );
  AND2_X1 U6640 ( .A1(n6192), .A2(n9548), .ZN(n9536) );
  OR2_X1 U6641 ( .A1(n5174), .A2(n5176), .ZN(n5140) );
  XNOR2_X1 U6642 ( .A(n5140), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6777) );
  INV_X1 U6643 ( .A(n6777), .ZN(n9497) );
  XNOR2_X1 U6644 ( .A(n5141), .B(n5142), .ZN(n6726) );
  NAND2_X1 U6645 ( .A1(n5192), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6646 ( .A1(n4288), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6647 ( .A1(n5469), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6648 ( .A1(n4910), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6649 ( .A1(n5611), .A2(n5150), .ZN(n5578) );
  NAND2_X1 U6650 ( .A1(n5855), .A2(n5151), .ZN(n9519) );
  NAND2_X1 U6651 ( .A1(n5578), .A2(n9519), .ZN(n7566) );
  NAND2_X1 U6652 ( .A1(n7565), .A2(n7566), .ZN(n5153) );
  NAND2_X1 U6653 ( .A1(n5150), .A2(n5151), .ZN(n5152) );
  NAND2_X1 U6654 ( .A1(n5153), .A2(n5152), .ZN(n9527) );
  INV_X1 U6655 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U6656 ( .A1(n5469), .A2(n9524), .ZN(n5157) );
  NAND2_X1 U6657 ( .A1(n5192), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6658 ( .A1(n4910), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5155) );
  INV_X1 U6659 ( .A(n4288), .ZN(n5267) );
  NAND2_X1 U6660 ( .A1(n4288), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5154) );
  INV_X1 U6661 ( .A(n9045), .ZN(n5163) );
  NAND2_X1 U6662 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4330), .ZN(n5158) );
  XNOR2_X1 U6663 ( .A(n5158), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6776) );
  INV_X1 U6664 ( .A(n6776), .ZN(n6800) );
  XNOR2_X1 U6665 ( .A(n5159), .B(n5160), .ZN(n6731) );
  OR2_X1 U6666 ( .A1(n5143), .A2(n6731), .ZN(n5162) );
  OR2_X1 U6667 ( .A1(n5184), .A2(n6718), .ZN(n5161) );
  OAI211_X1 U6668 ( .C1(n6743), .C2(n6800), .A(n5162), .B(n5161), .ZN(n6963)
         );
  NAND2_X1 U6669 ( .A1(n5163), .A2(n6963), .ZN(n5580) );
  NAND2_X1 U6670 ( .A1(n9045), .A2(n9573), .ZN(n5579) );
  NAND2_X1 U6671 ( .A1(n5580), .A2(n5579), .ZN(n9528) );
  NAND2_X1 U6672 ( .A1(n9527), .A2(n9528), .ZN(n5165) );
  NAND2_X1 U6673 ( .A1(n5163), .A2(n9573), .ZN(n5164) );
  NAND2_X1 U6674 ( .A1(n5165), .A2(n5164), .ZN(n7310) );
  NAND2_X1 U6675 ( .A1(n4910), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6676 ( .A1(n5192), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5171) );
  INV_X1 U6677 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6678 ( .A1(n9524), .A2(n5166), .ZN(n5167) );
  NAND2_X1 U6679 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5190) );
  AND2_X1 U6680 ( .A1(n5167), .A2(n5190), .ZN(n7068) );
  NAND2_X1 U6681 ( .A1(n5469), .A2(n7068), .ZN(n5170) );
  NAND2_X1 U6682 ( .A1(n4288), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5169) );
  NOR2_X1 U6683 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5173) );
  AND2_X1 U6684 ( .A1(n5174), .A2(n5173), .ZN(n5179) );
  NOR2_X1 U6685 ( .A1(n5179), .A2(n5176), .ZN(n5175) );
  MUX2_X1 U6686 ( .A(n5176), .B(n5175), .S(P1_IR_REG_4__SCAN_IN), .Z(n5177) );
  INV_X1 U6687 ( .A(n5177), .ZN(n5181) );
  INV_X1 U6688 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5178) );
  INV_X1 U6689 ( .A(n5216), .ZN(n5180) );
  NAND2_X1 U6690 ( .A1(n5181), .A2(n5180), .ZN(n6872) );
  OR2_X1 U6691 ( .A1(n5184), .A2(n6719), .ZN(n5185) );
  NAND2_X1 U6692 ( .A1(n4462), .A2(n7323), .ZN(n5187) );
  NAND2_X1 U6693 ( .A1(n5188), .A2(n5187), .ZN(n7088) );
  NAND2_X1 U6694 ( .A1(n4288), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6695 ( .A1(n6088), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5195) );
  INV_X1 U6696 ( .A(n5190), .ZN(n5189) );
  NAND2_X1 U6697 ( .A1(n5189), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5208) );
  INV_X1 U6698 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U6699 ( .A1(n5190), .A2(n7130), .ZN(n5191) );
  AND2_X1 U6700 ( .A1(n5208), .A2(n5191), .ZN(n7455) );
  NAND2_X1 U6701 ( .A1(n5469), .A2(n7455), .ZN(n5194) );
  NAND2_X1 U6702 ( .A1(n6087), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5193) );
  INV_X1 U6703 ( .A(n9043), .ZN(n5203) );
  XNOR2_X1 U6704 ( .A(n5197), .B(SI_5_), .ZN(n5198) );
  XNOR2_X1 U6705 ( .A(n5199), .B(n5198), .ZN(n6733) );
  OR2_X1 U6706 ( .A1(n6733), .A2(n5143), .ZN(n5202) );
  OR2_X1 U6707 ( .A1(n5216), .A2(n5176), .ZN(n5200) );
  AOI22_X1 U6708 ( .A1(n5420), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4291), .B2(
        n6813), .ZN(n5201) );
  NAND2_X1 U6709 ( .A1(n5203), .A2(n7456), .ZN(n5582) );
  NAND2_X1 U6710 ( .A1(n7131), .A2(n9043), .ZN(n6261) );
  AND2_X1 U6711 ( .A1(n5582), .A2(n6261), .ZN(n6198) );
  NAND2_X1 U6712 ( .A1(n7088), .A2(n7089), .ZN(n5205) );
  NAND2_X1 U6713 ( .A1(n5203), .A2(n7131), .ZN(n5204) );
  NAND2_X1 U6714 ( .A1(n5205), .A2(n5204), .ZN(n7445) );
  NAND2_X1 U6715 ( .A1(n5601), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5211) );
  INV_X1 U6716 ( .A(n5208), .ZN(n5206) );
  NAND2_X1 U6717 ( .A1(n5206), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5232) );
  INV_X1 U6718 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6719 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  AND2_X1 U6720 ( .A1(n5232), .A2(n5209), .ZN(n7449) );
  NAND2_X1 U6721 ( .A1(n5469), .A2(n7449), .ZN(n5210) );
  INV_X1 U6722 ( .A(n5212), .ZN(n5213) );
  XNOR2_X1 U6723 ( .A(n5214), .B(n5213), .ZN(n6728) );
  NAND2_X1 U6724 ( .A1(n6728), .A2(n6182), .ZN(n5218) );
  INV_X1 U6725 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6726 ( .A1(n5216), .A2(n5215), .ZN(n5247) );
  NAND2_X1 U6727 ( .A1(n5247), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6728 ( .A(n5226), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U6729 ( .A1(n5420), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4291), .B2(
        n6824), .ZN(n5217) );
  NAND2_X1 U6730 ( .A1(n5218), .A2(n5217), .ZN(n7450) );
  OR2_X1 U6731 ( .A1(n5219), .A2(n7450), .ZN(n6098) );
  NAND2_X1 U6732 ( .A1(n6098), .A2(n6197), .ZN(n7446) );
  NAND2_X1 U6733 ( .A1(n7445), .A2(n7446), .ZN(n5221) );
  OR2_X1 U6734 ( .A1(n7450), .A2(n9042), .ZN(n5220) );
  NAND2_X1 U6735 ( .A1(n5221), .A2(n5220), .ZN(n9502) );
  OR2_X1 U6736 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  AND2_X1 U6737 ( .A1(n5225), .A2(n5224), .ZN(n6747) );
  NAND2_X1 U6738 ( .A1(n6747), .A2(n6182), .ZN(n5230) );
  INV_X1 U6739 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6740 ( .A1(n5226), .A2(n5245), .ZN(n5227) );
  NAND2_X1 U6741 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6742 ( .A(n5228), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6906) );
  AOI22_X1 U6743 ( .A1(n5420), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4291), .B2(
        n6906), .ZN(n5229) );
  NAND2_X1 U6744 ( .A1(n5230), .A2(n5229), .ZN(n5899) );
  NAND2_X1 U6745 ( .A1(n5601), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6746 ( .A1(n6088), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5236) );
  INV_X1 U6747 ( .A(n5232), .ZN(n5231) );
  NAND2_X1 U6748 ( .A1(n5231), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5254) );
  INV_X1 U6749 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U6750 ( .A1(n5232), .A2(n6828), .ZN(n5233) );
  AND2_X1 U6751 ( .A1(n5254), .A2(n5233), .ZN(n9510) );
  NAND2_X1 U6752 ( .A1(n5469), .A2(n9510), .ZN(n5235) );
  NAND2_X1 U6753 ( .A1(n6087), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5234) );
  NAND4_X1 U6754 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n9041)
         );
  INV_X1 U6755 ( .A(n9041), .ZN(n5238) );
  OR2_X1 U6756 ( .A1(n5899), .A2(n5238), .ZN(n6100) );
  NAND2_X1 U6757 ( .A1(n5899), .A2(n5238), .ZN(n7485) );
  NAND2_X1 U6758 ( .A1(n6100), .A2(n7485), .ZN(n9504) );
  NAND2_X1 U6759 ( .A1(n9502), .A2(n9504), .ZN(n5240) );
  OR2_X1 U6760 ( .A1(n5899), .A2(n9041), .ZN(n5239) );
  NAND2_X1 U6761 ( .A1(n5240), .A2(n5239), .ZN(n7491) );
  NAND2_X1 U6762 ( .A1(n6759), .A2(n6182), .ZN(n5251) );
  NAND2_X1 U6763 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  OAI21_X1 U6764 ( .B1(n5247), .B2(n5246), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5248) );
  MUX2_X1 U6765 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5248), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5249) );
  AND2_X1 U6766 ( .A1(n5243), .A2(n5249), .ZN(n6973) );
  AOI22_X1 U6767 ( .A1(n5420), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4291), .B2(
        n6973), .ZN(n5250) );
  NAND2_X1 U6768 ( .A1(n5601), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6769 ( .A1(n6087), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5258) );
  INV_X1 U6770 ( .A(n5254), .ZN(n5252) );
  NAND2_X1 U6771 ( .A1(n5252), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5268) );
  INV_X1 U6772 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6773 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  AND2_X1 U6774 ( .A1(n5268), .A2(n5255), .ZN(n7494) );
  NAND2_X1 U6775 ( .A1(n5469), .A2(n7494), .ZN(n5257) );
  NAND2_X1 U6776 ( .A1(n6088), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6777 ( .A1(n7495), .A2(n5260), .ZN(n7502) );
  NAND2_X1 U6778 ( .A1(n7495), .A2(n5260), .ZN(n7501) );
  NAND2_X1 U6779 ( .A1(n7502), .A2(n7501), .ZN(n7492) );
  OR2_X1 U6780 ( .A1(n7495), .A2(n9040), .ZN(n5261) );
  XNOR2_X1 U6781 ( .A(n5263), .B(n5262), .ZN(n6816) );
  NAND2_X1 U6782 ( .A1(n6816), .A2(n6182), .ZN(n5266) );
  NAND2_X1 U6783 ( .A1(n5243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5264) );
  XNOR2_X1 U6784 ( .A(n5264), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7076) );
  AOI22_X1 U6785 ( .A1(n5420), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4291), .B2(
        n7076), .ZN(n5265) );
  NAND2_X1 U6786 ( .A1(n6087), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6787 ( .A1(n5601), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6788 ( .A1(n5268), .A2(n6977), .ZN(n5269) );
  AND2_X1 U6789 ( .A1(n5282), .A2(n5269), .ZN(n7517) );
  NAND2_X1 U6790 ( .A1(n5469), .A2(n7517), .ZN(n5271) );
  NAND2_X1 U6791 ( .A1(n6088), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5270) );
  OR2_X1 U6792 ( .A1(n9608), .A2(n5274), .ZN(n6121) );
  NAND2_X1 U6793 ( .A1(n9608), .A2(n5274), .ZN(n6112) );
  NAND2_X1 U6794 ( .A1(n6121), .A2(n6112), .ZN(n7510) );
  NAND2_X1 U6795 ( .A1(n4348), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6796 ( .A1(n5277), .A2(n5276), .ZN(n6821) );
  OR2_X1 U6797 ( .A1(n6821), .A2(n5143), .ZN(n5279) );
  NOR2_X1 U6798 ( .A1(n5243), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6799 ( .A1(n5313), .A2(n5176), .ZN(n5294) );
  XNOR2_X1 U6800 ( .A(n5294), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7241) );
  AOI22_X1 U6801 ( .A1(n5420), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4291), .B2(
        n7241), .ZN(n5278) );
  NAND2_X1 U6802 ( .A1(n5279), .A2(n5278), .ZN(n7751) );
  NAND2_X1 U6803 ( .A1(n6087), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6804 ( .A1(n5601), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5286) );
  INV_X1 U6805 ( .A(n5282), .ZN(n5280) );
  NAND2_X1 U6806 ( .A1(n5280), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5299) );
  INV_X1 U6807 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6808 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AND2_X1 U6809 ( .A1(n5299), .A2(n5283), .ZN(n7377) );
  NAND2_X1 U6810 ( .A1(n5469), .A2(n7377), .ZN(n5285) );
  NAND2_X1 U6811 ( .A1(n6088), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5284) );
  NAND4_X1 U6812 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n9038)
         );
  INV_X1 U6813 ( .A(n9038), .ZN(n5288) );
  NOR2_X1 U6814 ( .A1(n7751), .A2(n5288), .ZN(n6111) );
  INV_X1 U6815 ( .A(n6111), .ZN(n6124) );
  NAND2_X1 U6816 ( .A1(n7751), .A2(n5288), .ZN(n7528) );
  NAND2_X1 U6817 ( .A1(n6124), .A2(n7528), .ZN(n7376) );
  NAND2_X1 U6818 ( .A1(n7375), .A2(n7376), .ZN(n5290) );
  OR2_X1 U6819 ( .A1(n7751), .A2(n9038), .ZN(n5289) );
  NAND2_X1 U6820 ( .A1(n5290), .A2(n5289), .ZN(n7524) );
  XNOR2_X1 U6821 ( .A(n5292), .B(n5291), .ZN(n6859) );
  NAND2_X1 U6822 ( .A1(n6859), .A2(n6182), .ZN(n5298) );
  INV_X1 U6823 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6824 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  NAND2_X1 U6825 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5296) );
  XNOR2_X1 U6826 ( .A(n5296), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U6827 ( .A1(n5420), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4291), .B2(
        n7242), .ZN(n5297) );
  NAND2_X1 U6828 ( .A1(n4288), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6829 ( .A1(n6088), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6830 ( .A1(n5299), .A2(n7858), .ZN(n5300) );
  AND2_X1 U6831 ( .A1(n5321), .A2(n5300), .ZN(n7862) );
  NAND2_X1 U6832 ( .A1(n5469), .A2(n7862), .ZN(n5302) );
  NAND2_X1 U6833 ( .A1(n6087), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5301) );
  NAND4_X1 U6834 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9037)
         );
  INV_X1 U6835 ( .A(n9037), .ZN(n5305) );
  NAND2_X1 U6836 ( .A1(n7536), .A2(n5305), .ZN(n6126) );
  NAND2_X1 U6837 ( .A1(n7524), .A2(n7525), .ZN(n5307) );
  OR2_X1 U6838 ( .A1(n7536), .A2(n9037), .ZN(n5306) );
  NAND2_X1 U6839 ( .A1(n5307), .A2(n5306), .ZN(n7464) );
  NAND2_X1 U6840 ( .A1(n5309), .A2(n5308), .ZN(n5311) );
  NAND2_X1 U6841 ( .A1(n5311), .A2(n5310), .ZN(n6919) );
  NOR2_X1 U6842 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5312) );
  NAND2_X1 U6843 ( .A1(n5313), .A2(n5312), .ZN(n5315) );
  NAND2_X1 U6844 ( .A1(n5315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5314) );
  MUX2_X1 U6845 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5314), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5316) );
  AOI22_X1 U6846 ( .A1(n5420), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4291), .B2(
        n7386), .ZN(n5317) );
  NAND2_X1 U6847 ( .A1(n6087), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6848 ( .A1(n4288), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5325) );
  INV_X1 U6849 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6850 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  AND2_X1 U6851 ( .A1(n5338), .A2(n5322), .ZN(n7658) );
  NAND2_X1 U6852 ( .A1(n5469), .A2(n7658), .ZN(n5324) );
  NAND2_X1 U6853 ( .A1(n6088), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5323) );
  NAND4_X1 U6854 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n7545)
         );
  INV_X1 U6855 ( .A(n7545), .ZN(n5327) );
  NAND2_X1 U6856 ( .A1(n7663), .A2(n5327), .ZN(n6127) );
  INV_X1 U6857 ( .A(n7466), .ZN(n7465) );
  NAND2_X1 U6858 ( .A1(n7464), .A2(n7465), .ZN(n5329) );
  NAND2_X1 U6859 ( .A1(n9626), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6860 ( .A1(n5332), .A2(n5331), .ZN(n5334) );
  NAND2_X1 U6861 ( .A1(n5334), .A2(n5333), .ZN(n8120) );
  NAND2_X1 U6862 ( .A1(n5350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5335) );
  XNOR2_X1 U6863 ( .A(n5335), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7667) );
  AOI22_X1 U6864 ( .A1(n5420), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4291), .B2(
        n7667), .ZN(n5336) );
  NAND2_X1 U6865 ( .A1(n6087), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6866 ( .A1(n4288), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6867 ( .A1(n5338), .A2(n7707), .ZN(n5339) );
  AND2_X1 U6868 ( .A1(n5354), .A2(n5339), .ZN(n7711) );
  NAND2_X1 U6869 ( .A1(n5469), .A2(n7711), .ZN(n5341) );
  NAND2_X1 U6870 ( .A1(n6088), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5340) );
  NAND4_X1 U6871 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n9036)
         );
  NOR2_X1 U6872 ( .A1(n5951), .A2(n9036), .ZN(n5344) );
  NAND2_X1 U6873 ( .A1(n5951), .A2(n9036), .ZN(n5345) );
  NAND2_X1 U6874 ( .A1(n5333), .A2(n5346), .ZN(n5349) );
  XNOR2_X1 U6875 ( .A(n5347), .B(SI_14_), .ZN(n5348) );
  XNOR2_X1 U6876 ( .A(n5349), .B(n5348), .ZN(n7096) );
  NAND2_X1 U6877 ( .A1(n7096), .A2(n6182), .ZN(n5353) );
  NAND2_X1 U6878 ( .A1(n5351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5366) );
  XNOR2_X1 U6879 ( .A(n5366), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7884) );
  AOI22_X1 U6880 ( .A1(n5420), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4291), .B2(
        n7884), .ZN(n5352) );
  NAND2_X1 U6881 ( .A1(n6087), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6882 ( .A1(n5601), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6883 ( .A1(n5354), .A2(n7949), .ZN(n5355) );
  AND2_X1 U6884 ( .A1(n5372), .A2(n5355), .ZN(n7952) );
  NAND2_X1 U6885 ( .A1(n5469), .A2(n7952), .ZN(n5357) );
  NAND2_X1 U6886 ( .A1(n6088), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5356) );
  NAND4_X1 U6887 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n9035)
         );
  AND2_X1 U6888 ( .A1(n9640), .A2(n9035), .ZN(n5361) );
  OR2_X1 U6889 ( .A1(n9640), .A2(n9035), .ZN(n5360) );
  XNOR2_X1 U6890 ( .A(n5363), .B(SI_15_), .ZN(n5364) );
  XNOR2_X1 U6891 ( .A(n5362), .B(n5364), .ZN(n7100) );
  NAND2_X1 U6892 ( .A1(n7100), .A2(n6182), .ZN(n5370) );
  INV_X1 U6893 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6894 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6895 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6896 ( .A(n5368), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9049) );
  AOI22_X1 U6897 ( .A1(n5420), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4291), .B2(
        n9049), .ZN(n5369) );
  INV_X1 U6898 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U6899 ( .A1(n5372), .A2(n9009), .ZN(n5373) );
  AND2_X1 U6900 ( .A1(n5392), .A2(n5373), .ZN(n9014) );
  NAND2_X1 U6901 ( .A1(n9014), .A2(n5469), .ZN(n5377) );
  NAND2_X1 U6902 ( .A1(n5601), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6903 ( .A1(n6088), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6904 ( .A1(n6087), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5374) );
  NAND4_X1 U6905 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n9034)
         );
  NAND2_X1 U6906 ( .A1(n7835), .A2(n9034), .ZN(n5378) );
  OR2_X1 U6907 ( .A1(n7835), .A2(n9034), .ZN(n5379) );
  XNOR2_X1 U6908 ( .A(n5381), .B(n5380), .ZN(n5382) );
  NAND2_X1 U6909 ( .A1(n7151), .A2(n6182), .ZN(n5387) );
  INV_X1 U6910 ( .A(n5061), .ZN(n5384) );
  NAND2_X1 U6911 ( .A1(n5384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U6912 ( .A(n5385), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9070) );
  AOI22_X1 U6913 ( .A1(n5420), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4291), .B2(
        n9070), .ZN(n5386) );
  INV_X1 U6914 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U6915 ( .A1(n5601), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6916 ( .A1(n6087), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5388) );
  AND2_X1 U6917 ( .A1(n5389), .A2(n5388), .ZN(n5395) );
  INV_X1 U6918 ( .A(n5392), .ZN(n5390) );
  INV_X1 U6919 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6920 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U6921 ( .A1(n5404), .A2(n5393), .ZN(n8944) );
  OR2_X1 U6922 ( .A1(n8944), .A2(n5563), .ZN(n5394) );
  OAI211_X1 U6923 ( .C1(n5430), .C2(n7812), .A(n5395), .B(n5394), .ZN(n9033)
         );
  INV_X1 U6924 ( .A(n9033), .ZN(n5396) );
  NAND2_X1 U6925 ( .A1(n8946), .A2(n9033), .ZN(n5397) );
  XNOR2_X1 U6926 ( .A(n5399), .B(n5398), .ZN(n7287) );
  NAND2_X1 U6927 ( .A1(n7287), .A2(n6182), .ZN(n5402) );
  XNOR2_X1 U6928 ( .A(n5400), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9083) );
  AOI22_X1 U6929 ( .A1(n5420), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4291), .B2(
        n9083), .ZN(n5401) );
  INV_X1 U6930 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6931 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U6932 ( .A1(n5426), .A2(n5405), .ZN(n8951) );
  AOI22_X1 U6933 ( .A1(n6087), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n4288), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6934 ( .A1(n6088), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5406) );
  OAI211_X1 U6935 ( .C1(n8951), .C2(n5563), .A(n5407), .B(n5406), .ZN(n9032)
         );
  OR2_X1 U6936 ( .A1(n7933), .A2(n9032), .ZN(n5408) );
  NAND2_X1 U6937 ( .A1(n7933), .A2(n9032), .ZN(n5409) );
  XNOR2_X1 U6938 ( .A(n5411), .B(n5410), .ZN(n7299) );
  NAND2_X1 U6939 ( .A1(n7299), .A2(n6182), .ZN(n5414) );
  XNOR2_X1 U6940 ( .A(n5412), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9111) );
  AOI22_X1 U6941 ( .A1(n5420), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4291), .B2(
        n9111), .ZN(n5413) );
  XNOR2_X1 U6942 ( .A(n5426), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9318) );
  INV_X1 U6943 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U6944 ( .A1(n6088), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6945 ( .A1(n4288), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6946 ( .C1(n5557), .C2(n9389), .A(n5416), .B(n5415), .ZN(n5417)
         );
  AOI21_X1 U6947 ( .B1(n9318), .B2(n5469), .A(n5417), .ZN(n8918) );
  XNOR2_X1 U6948 ( .A(n5419), .B(n5418), .ZN(n7557) );
  NAND2_X1 U6949 ( .A1(n7557), .A2(n6182), .ZN(n5422) );
  AOI22_X1 U6950 ( .A1(n5420), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4291), .B2(
        n9119), .ZN(n5421) );
  INV_X1 U6951 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9109) );
  AND2_X1 U6952 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5423) );
  INV_X1 U6953 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8984) );
  INV_X1 U6954 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5425) );
  OAI21_X1 U6955 ( .B1(n5426), .B2(n8984), .A(n5425), .ZN(n5427) );
  NAND2_X1 U6956 ( .A1(n5437), .A2(n5427), .ZN(n9293) );
  OR2_X1 U6957 ( .A1(n9293), .A2(n5563), .ZN(n5429) );
  AOI22_X1 U6958 ( .A1(n6087), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n4288), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5428) );
  OAI211_X1 U6959 ( .C1(n5430), .C2(n9109), .A(n5429), .B(n5428), .ZN(n9030)
         );
  NAND2_X1 U6960 ( .A1(n9380), .A2(n9030), .ZN(n5431) );
  XNOR2_X1 U6961 ( .A(n5432), .B(n10036), .ZN(n5433) );
  XNOR2_X1 U6962 ( .A(n5434), .B(n5433), .ZN(n7681) );
  NAND2_X1 U6963 ( .A1(n7681), .A2(n6182), .ZN(n5436) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7685) );
  OR2_X1 U6965 ( .A1(n5184), .A2(n7685), .ZN(n5435) );
  NAND2_X1 U6966 ( .A1(n5437), .A2(n10064), .ZN(n5438) );
  AND2_X1 U6967 ( .A1(n5453), .A2(n5438), .ZN(n9286) );
  NAND2_X1 U6968 ( .A1(n9286), .A2(n5469), .ZN(n5444) );
  INV_X1 U6969 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6970 ( .A1(n5601), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6971 ( .A1(n6088), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5439) );
  OAI211_X1 U6972 ( .C1(n5441), .C2(n5557), .A(n5440), .B(n5439), .ZN(n5442)
         );
  INV_X1 U6973 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6974 ( .A1(n5444), .A2(n5443), .ZN(n8926) );
  AND2_X1 U6975 ( .A1(n9377), .A2(n8926), .ZN(n5445) );
  XNOR2_X1 U6976 ( .A(n5446), .B(SI_21_), .ZN(n5447) );
  XNOR2_X1 U6977 ( .A(n5448), .B(n5447), .ZN(n7720) );
  NAND2_X1 U6978 ( .A1(n7720), .A2(n6182), .ZN(n5450) );
  OR2_X1 U6979 ( .A1(n5184), .A2(n7721), .ZN(n5449) );
  INV_X1 U6980 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6981 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  NAND2_X1 U6982 ( .A1(n5467), .A2(n5454), .ZN(n9267) );
  OR2_X1 U6983 ( .A1(n9267), .A2(n5563), .ZN(n5459) );
  INV_X1 U6984 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U6985 ( .A1(n6087), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6986 ( .A1(n6088), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5455) );
  OAI211_X1 U6987 ( .C1(n5267), .C2(n10037), .A(n5456), .B(n5455), .ZN(n5457)
         );
  INV_X1 U6988 ( .A(n5457), .ZN(n5458) );
  NAND2_X1 U6989 ( .A1(n5459), .A2(n5458), .ZN(n9029) );
  INV_X1 U6990 ( .A(n9029), .ZN(n5460) );
  NAND2_X1 U6991 ( .A1(n9427), .A2(n5460), .ZN(n6159) );
  NAND2_X1 U6992 ( .A1(n9427), .A2(n9029), .ZN(n5462) );
  XNOR2_X1 U6993 ( .A(n5464), .B(n5463), .ZN(n7877) );
  NAND2_X1 U6994 ( .A1(n7877), .A2(n6182), .ZN(n5466) );
  OR2_X1 U6995 ( .A1(n5184), .A2(n7882), .ZN(n5465) );
  INV_X1 U6996 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U6997 ( .A1(n5467), .A2(n8976), .ZN(n5468) );
  AND2_X1 U6998 ( .A1(n5484), .A2(n5468), .ZN(n9252) );
  NAND2_X1 U6999 ( .A1(n9252), .A2(n5469), .ZN(n5474) );
  INV_X1 U7000 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U7001 ( .A1(n5601), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7002 ( .A1(n6088), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U7003 ( .C1(n9367), .C2(n5557), .A(n5471), .B(n5470), .ZN(n5472)
         );
  INV_X1 U7004 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U7005 ( .A1(n5474), .A2(n5473), .ZN(n9028) );
  AND2_X1 U7006 ( .A1(n6008), .A2(n9028), .ZN(n5475) );
  OR2_X1 U7007 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  NAND2_X1 U7008 ( .A1(n5476), .A2(n5479), .ZN(n7900) );
  NAND2_X1 U7009 ( .A1(n7900), .A2(n6182), .ZN(n5481) );
  OR2_X1 U7010 ( .A1(n5184), .A2(n7898), .ZN(n5480) );
  INV_X1 U7011 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7012 ( .A1(n5484), .A2(n5483), .ZN(n5485) );
  NAND2_X1 U7013 ( .A1(n5503), .A2(n5485), .ZN(n8911) );
  OR2_X1 U7014 ( .A1(n8911), .A2(n5563), .ZN(n5490) );
  INV_X1 U7015 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U7016 ( .A1(n5601), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7017 ( .A1(n6088), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5486) );
  OAI211_X1 U7018 ( .C1(n5557), .C2(n9362), .A(n5487), .B(n5486), .ZN(n5488)
         );
  INV_X1 U7019 ( .A(n5488), .ZN(n5489) );
  NOR2_X1 U7020 ( .A1(n9235), .A2(n9027), .ZN(n5491) );
  NAND2_X1 U7021 ( .A1(n9235), .A2(n9027), .ZN(n5492) );
  NAND2_X1 U7022 ( .A1(n5476), .A2(n5494), .ZN(n5498) );
  AND2_X1 U7023 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U7024 ( .A1(n7979), .A2(n6182), .ZN(n5500) );
  OR2_X1 U7025 ( .A1(n5184), .A2(n7980), .ZN(n5499) );
  INV_X1 U7026 ( .A(n5503), .ZN(n5501) );
  NAND2_X1 U7027 ( .A1(n5501), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5516) );
  INV_X1 U7028 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7029 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  NAND2_X1 U7030 ( .A1(n5516), .A2(n5504), .ZN(n8959) );
  INV_X1 U7031 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7032 ( .A1(n5601), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7033 ( .A1(n6088), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5505) );
  OAI211_X1 U7034 ( .C1(n5557), .C2(n5507), .A(n5506), .B(n5505), .ZN(n5508)
         );
  INV_X1 U7035 ( .A(n5508), .ZN(n5509) );
  AND2_X1 U7036 ( .A1(n9354), .A2(n9026), .ZN(n5511) );
  XNOR2_X1 U7037 ( .A(n5513), .B(n5512), .ZN(n7990) );
  NAND2_X1 U7038 ( .A1(n7990), .A2(n6182), .ZN(n5515) );
  OR2_X1 U7039 ( .A1(n5184), .A2(n7991), .ZN(n5514) );
  INV_X1 U7040 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U7041 ( .A1(n5516), .A2(n8935), .ZN(n5517) );
  NAND2_X1 U7042 ( .A1(n5528), .A2(n5517), .ZN(n9201) );
  OR2_X1 U7043 ( .A1(n9201), .A2(n5563), .ZN(n5522) );
  INV_X1 U7044 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U7045 ( .A1(n6087), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7046 ( .A1(n6088), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5518) );
  OAI211_X1 U7047 ( .C1(n5267), .C2(n10053), .A(n5519), .B(n5518), .ZN(n5520)
         );
  INV_X1 U7048 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7049 ( .A1(n5522), .A2(n5521), .ZN(n9025) );
  NAND2_X1 U7050 ( .A1(n9348), .A2(n9025), .ZN(n5523) );
  NAND2_X1 U7051 ( .A1(n8084), .A2(n6182), .ZN(n5527) );
  OR2_X1 U7052 ( .A1(n5184), .A2(n9959), .ZN(n5526) );
  INV_X1 U7053 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U7054 ( .A1(n5528), .A2(n8997), .ZN(n5529) );
  INV_X1 U7055 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7056 ( .A1(n6088), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7057 ( .A1(n5601), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5530) );
  OAI211_X1 U7058 ( .C1(n5557), .C2(n9346), .A(n5531), .B(n5530), .ZN(n5532)
         );
  AOI21_X1 U7059 ( .B1(n9193), .B2(n5469), .A(n5532), .ZN(n6032) );
  INV_X1 U7060 ( .A(n6032), .ZN(n9024) );
  NAND2_X1 U7061 ( .A1(n9413), .A2(n9024), .ZN(n6228) );
  NAND2_X1 U7062 ( .A1(n6288), .A2(n6228), .ZN(n9190) );
  OR2_X1 U7063 ( .A1(n9413), .A2(n6032), .ZN(n5533) );
  NAND2_X1 U7064 ( .A1(n8103), .A2(n6182), .ZN(n5538) );
  OR2_X1 U7065 ( .A1(n5184), .A2(n8107), .ZN(n5537) );
  INV_X1 U7066 ( .A(n5540), .ZN(n5539) );
  NAND2_X1 U7067 ( .A1(n5539), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9138) );
  INV_X1 U7068 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7069 ( .A1(n5540), .A2(n6709), .ZN(n5541) );
  NAND2_X1 U7070 ( .A1(n9138), .A2(n5541), .ZN(n9179) );
  INV_X1 U7071 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U7072 ( .A1(n6087), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7073 ( .A1(n6088), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U7074 ( .C1(n5267), .C2(n9407), .A(n5543), .B(n5542), .ZN(n5544)
         );
  INV_X1 U7075 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U7076 ( .A1(n5546), .A2(n5545), .ZN(n9023) );
  INV_X1 U7077 ( .A(n9023), .ZN(n8996) );
  OR2_X1 U7078 ( .A1(n9178), .A2(n8996), .ZN(n6291) );
  NAND2_X1 U7079 ( .A1(n9178), .A2(n8996), .ZN(n9146) );
  NAND2_X1 U7080 ( .A1(n6291), .A2(n9146), .ZN(n6213) );
  NAND2_X1 U7081 ( .A1(n5548), .A2(n5547), .ZN(n5552) );
  AND2_X1 U7082 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7083 ( .A1(n8113), .A2(n6182), .ZN(n5554) );
  OR2_X1 U7084 ( .A1(n5184), .A2(n8114), .ZN(n5553) );
  XNOR2_X1 U7085 ( .A(n9138), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U7086 ( .A1(n9164), .A2(n5469), .ZN(n5560) );
  INV_X1 U7087 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U7088 ( .A1(n6088), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7089 ( .A1(n4288), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5555) );
  OAI211_X1 U7090 ( .C1(n5557), .C2(n9984), .A(n5556), .B(n5555), .ZN(n5558)
         );
  INV_X1 U7091 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7092 ( .A1(n5560), .A2(n5559), .ZN(n9022) );
  INV_X1 U7093 ( .A(n9022), .ZN(n5561) );
  NAND2_X1 U7094 ( .A1(n9404), .A2(n5561), .ZN(n5596) );
  NAND2_X1 U7095 ( .A1(n9149), .A2(n5596), .ZN(n9156) );
  NAND2_X1 U7096 ( .A1(n9155), .A2(n9156), .ZN(n9160) );
  NAND2_X1 U7097 ( .A1(n9404), .A2(n9022), .ZN(n5562) );
  NAND2_X1 U7098 ( .A1(n9160), .A2(n5562), .ZN(n5571) );
  INV_X1 U7099 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5564) );
  OR3_X1 U7100 ( .A1(n9138), .A2(n5564), .A3(n5563), .ZN(n5569) );
  NAND2_X1 U7101 ( .A1(n6088), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7102 ( .A1(n6087), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7103 ( .A1(n4288), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5565) );
  AND3_X1 U7104 ( .A1(n5567), .A2(n5566), .A3(n5565), .ZN(n5568) );
  NAND2_X1 U7105 ( .A1(n5569), .A2(n5568), .ZN(n9021) );
  INV_X1 U7106 ( .A(n9021), .ZN(n5570) );
  NAND2_X1 U7107 ( .A1(n9140), .A2(n5570), .ZN(n6189) );
  NAND2_X1 U7108 ( .A1(n6244), .A2(n6189), .ZN(n6179) );
  XNOR2_X1 U7109 ( .A(n5571), .B(n4489), .ZN(n9135) );
  AND2_X1 U7110 ( .A1(n5834), .A2(n6305), .ZN(n5573) );
  OAI21_X1 U7111 ( .B1(n5834), .B2(n6313), .A(n6842), .ZN(n7350) );
  OR2_X1 U7112 ( .A1(n5573), .A2(n7350), .ZN(n9537) );
  NAND2_X1 U7113 ( .A1(n7880), .A2(n9119), .ZN(n6307) );
  NAND2_X1 U7114 ( .A1(n9135), .A2(n9635), .ZN(n5615) );
  INV_X1 U7115 ( .A(n9190), .ZN(n9186) );
  INV_X1 U7116 ( .A(n8918), .ZN(n9031) );
  NAND2_X1 U7117 ( .A1(n9437), .A2(n9031), .ZN(n6148) );
  INV_X1 U7118 ( .A(n9309), .ZN(n9313) );
  INV_X1 U7119 ( .A(n9032), .ZN(n7809) );
  OR2_X1 U7120 ( .A1(n7933), .A2(n7809), .ZN(n6143) );
  NAND2_X1 U7121 ( .A1(n7933), .A2(n7809), .ZN(n6145) );
  NAND2_X1 U7122 ( .A1(n6143), .A2(n6145), .ZN(n6208) );
  INV_X1 U7123 ( .A(n9035), .ZN(n5574) );
  NAND2_X1 U7124 ( .A1(n9640), .A2(n5574), .ZN(n6131) );
  NAND2_X1 U7125 ( .A1(n7828), .A2(n6131), .ZN(n7643) );
  INV_X1 U7126 ( .A(n9036), .ZN(n5575) );
  INV_X1 U7127 ( .A(n9047), .ZN(n5576) );
  NAND2_X1 U7128 ( .A1(n5576), .A2(n9549), .ZN(n5577) );
  AND2_X1 U7129 ( .A1(n9519), .A2(n5579), .ZN(n6265) );
  INV_X1 U7130 ( .A(n6099), .ZN(n5584) );
  NAND2_X1 U7131 ( .A1(n7501), .A2(n7485), .ZN(n6101) );
  AND2_X1 U7132 ( .A1(n5583), .A2(n6112), .ZN(n6203) );
  NAND2_X1 U7133 ( .A1(n5584), .A2(n6203), .ZN(n6266) );
  NAND2_X1 U7134 ( .A1(n6100), .A2(n6098), .ZN(n5585) );
  OR2_X1 U7135 ( .A1(n6107), .A2(n5585), .ZN(n6201) );
  NAND2_X1 U7136 ( .A1(n6203), .A2(n6201), .ZN(n6270) );
  AND2_X2 U7137 ( .A1(n6266), .A2(n6270), .ZN(n7370) );
  INV_X1 U7138 ( .A(n7376), .ZN(n7371) );
  INV_X1 U7139 ( .A(n7528), .ZN(n5586) );
  NOR2_X1 U7140 ( .A1(n7525), .A2(n5586), .ZN(n5587) );
  NAND2_X1 U7141 ( .A1(n7526), .A2(n6125), .ZN(n7467) );
  NAND2_X1 U7142 ( .A1(n9633), .A2(n9036), .ZN(n6276) );
  INV_X1 U7143 ( .A(n7644), .ZN(n6273) );
  NAND2_X1 U7144 ( .A1(n6276), .A2(n6273), .ZN(n7551) );
  INV_X1 U7145 ( .A(n9034), .ZN(n7808) );
  OR2_X1 U7146 ( .A1(n7835), .A2(n7808), .ZN(n6095) );
  AND2_X1 U7147 ( .A1(n7835), .A2(n7808), .ZN(n6092) );
  NAND3_X1 U7148 ( .A1(n7829), .A2(n7833), .A3(n7828), .ZN(n5588) );
  NAND2_X1 U7149 ( .A1(n5588), .A2(n6132), .ZN(n7807) );
  INV_X1 U7150 ( .A(n7815), .ZN(n7806) );
  NAND2_X1 U7151 ( .A1(n7936), .A2(n7927), .ZN(n7926) );
  INV_X1 U7152 ( .A(n9030), .ZN(n5589) );
  OR2_X1 U7153 ( .A1(n9380), .A2(n5589), .ZN(n6153) );
  NAND2_X1 U7154 ( .A1(n9380), .A2(n5589), .ZN(n6149) );
  INV_X1 U7155 ( .A(n6149), .ZN(n6285) );
  INV_X1 U7156 ( .A(n8926), .ZN(n8919) );
  NAND2_X1 U7157 ( .A1(n9377), .A2(n8919), .ZN(n6158) );
  NAND2_X1 U7158 ( .A1(n6154), .A2(n6158), .ZN(n9276) );
  INV_X1 U7159 ( .A(n9276), .ZN(n9279) );
  INV_X1 U7160 ( .A(n9028), .ZN(n5590) );
  OR2_X1 U7161 ( .A1(n6008), .A2(n5590), .ZN(n6160) );
  NAND2_X1 U7162 ( .A1(n6008), .A2(n5590), .ZN(n6162) );
  NAND2_X1 U7163 ( .A1(n6160), .A2(n6162), .ZN(n9244) );
  INV_X1 U7164 ( .A(n9244), .ZN(n9248) );
  NAND2_X1 U7165 ( .A1(n9245), .A2(n9248), .ZN(n5591) );
  NAND2_X1 U7166 ( .A1(n5591), .A2(n6162), .ZN(n9230) );
  XNOR2_X1 U7167 ( .A(n9235), .B(n9027), .ZN(n9233) );
  INV_X1 U7168 ( .A(n9027), .ZN(n6164) );
  NAND2_X1 U7169 ( .A1(n9235), .A2(n6164), .ZN(n6218) );
  INV_X1 U7170 ( .A(n9026), .ZN(n5593) );
  NAND2_X1 U7171 ( .A1(n9354), .A2(n5593), .ZN(n6233) );
  NAND2_X1 U7172 ( .A1(n6221), .A2(n6233), .ZN(n9220) );
  INV_X1 U7173 ( .A(n9220), .ZN(n5594) );
  INV_X1 U7174 ( .A(n9025), .ZN(n8994) );
  OR2_X1 U7175 ( .A1(n9348), .A2(n8994), .ZN(n6224) );
  AND2_X1 U7176 ( .A1(n9348), .A2(n8994), .ZN(n6236) );
  NAND2_X1 U7177 ( .A1(n6224), .A2(n6171), .ZN(n9203) );
  NAND2_X1 U7178 ( .A1(n9186), .A2(n9187), .ZN(n5595) );
  NAND2_X1 U7179 ( .A1(n5596), .A2(n9146), .ZN(n6242) );
  INV_X1 U7180 ( .A(n6242), .ZN(n6175) );
  NAND2_X1 U7181 ( .A1(n9148), .A2(n9149), .ZN(n5597) );
  XNOR2_X1 U7182 ( .A(n6179), .B(n5597), .ZN(n5610) );
  NAND2_X1 U7183 ( .A1(n6316), .A2(n9119), .ZN(n5600) );
  NAND2_X1 U7184 ( .A1(n5572), .A2(n5598), .ZN(n5599) );
  NAND2_X1 U7185 ( .A1(n6087), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7186 ( .A1(n6088), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7187 ( .A1(n5601), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5602) );
  AND3_X1 U7188 ( .A1(n5604), .A2(n5603), .A3(n5602), .ZN(n6191) );
  INV_X1 U7189 ( .A(n6742), .ZN(n5607) );
  NAND2_X1 U7190 ( .A1(n5607), .A2(n5605), .ZN(n8995) );
  INV_X1 U7191 ( .A(n4294), .ZN(n6866) );
  NAND2_X1 U7192 ( .A1(n6866), .A2(P1_B_REG_SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7193 ( .A1(n8983), .A2(n5606), .ZN(n9124) );
  NAND2_X1 U7194 ( .A1(n9022), .A2(n8982), .ZN(n5608) );
  OAI21_X1 U7195 ( .B1(n6191), .B2(n9124), .A(n5608), .ZN(n5609) );
  AOI21_X2 U7196 ( .B1(n5610), .B2(n9541), .A(n5609), .ZN(n9145) );
  INV_X1 U7197 ( .A(n7450), .ZN(n9589) );
  INV_X1 U7198 ( .A(n5899), .ZN(n9593) );
  NAND2_X1 U7199 ( .A1(n9515), .A2(n9593), .ZN(n9514) );
  OR2_X1 U7200 ( .A1(n9514), .A2(n7495), .ZN(n7511) );
  INV_X1 U7201 ( .A(n7751), .ZN(n9616) );
  AND2_X1 U7202 ( .A1(n7513), .A2(n9616), .ZN(n7535) );
  AOI21_X1 U7203 ( .B1(n9140), .B2(n9162), .A(n9620), .ZN(n5613) );
  NAND2_X1 U7204 ( .A1(n5613), .A2(n9128), .ZN(n9142) );
  INV_X1 U7205 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5616) );
  OR2_X1 U7206 ( .A1(n10083), .A2(n5616), .ZN(n5617) );
  NAND2_X1 U7207 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  INV_X1 U7208 ( .A(n9428), .ZN(n5626) );
  INV_X1 U7209 ( .A(n9140), .ZN(n5625) );
  AOI21_X1 U7210 ( .B1(n5622), .B2(n9650), .A(n4899), .ZN(n5624) );
  OAI21_X1 U7211 ( .B1(n5626), .B2(n5625), .A(n5624), .ZN(P1_U3519) );
  NOR2_X4 U7212 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5693) );
  NOR2_X1 U7213 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5628) );
  NAND3_X1 U7214 ( .A1(n5665), .A2(n5629), .A3(n5668), .ZN(n5630) );
  NAND2_X1 U7215 ( .A1(n5650), .A2(n5649), .ZN(n5633) );
  INV_X1 U7216 ( .A(n8117), .ZN(n5648) );
  NAND2_X1 U7217 ( .A1(n5639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5638) );
  MUX2_X1 U7218 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5638), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5642) );
  INV_X1 U7219 ( .A(n5639), .ZN(n5641) );
  INV_X1 U7220 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7221 ( .A1(n5644), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5646) );
  NOR2_X1 U7222 ( .A1(n8086), .A2(n8172), .ZN(n5647) );
  INV_X1 U7223 ( .A(n6950), .ZN(n5651) );
  NAND2_X1 U7224 ( .A1(n4363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7225 ( .A1(n5653), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7226 ( .A1(n6698), .A2(n8310), .ZN(n5655) );
  NAND2_X1 U7227 ( .A1(n5655), .A2(n5826), .ZN(n5824) );
  INV_X1 U7228 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7229 ( .A1(n5659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5660) );
  NAND2_X4 U7230 ( .A1(n5661), .A2(n6322), .ZN(n6847) );
  NAND2_X1 U7231 ( .A1(n5824), .A2(n6661), .ZN(n5662) );
  NAND2_X1 U7232 ( .A1(n5662), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U7233 ( .A1(n5664), .A2(n5665), .ZN(n5687) );
  INV_X1 U7234 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7235 ( .A1(n5687), .A2(n5667), .ZN(n5743) );
  OAI21_X1 U7236 ( .B1(n5743), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U7237 ( .A(n7559), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7238 ( .A1(n5687), .A2(n5670), .ZN(n5689) );
  NOR2_X1 U7239 ( .A1(n5680), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5678) );
  INV_X1 U7240 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7241 ( .A1(n5678), .A2(n5671), .ZN(n5672) );
  NAND2_X1 U7242 ( .A1(n5672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5675) );
  INV_X1 U7243 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7244 ( .A1(n5675), .A2(n5674), .ZN(n5677) );
  NAND2_X1 U7245 ( .A1(n5677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U7246 ( .A(n5673), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9810) );
  OR2_X1 U7247 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  INV_X1 U7248 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5694) );
  OR2_X1 U7249 ( .A1(n5678), .A2(n5694), .ZN(n5679) );
  XNOR2_X1 U7250 ( .A(n5679), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U7251 ( .A1(n5680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5682) );
  INV_X1 U7252 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5681) );
  XNOR2_X1 U7253 ( .A(n5682), .B(n5681), .ZN(n9790) );
  NAND2_X1 U7254 ( .A1(n5683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  XNOR2_X1 U7255 ( .A(n5684), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U7256 ( .A1(n5689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5686) );
  INV_X1 U7257 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U7258 ( .A(n5686), .B(n5685), .ZN(n6918) );
  NOR2_X1 U7259 ( .A1(n5687), .A2(n5694), .ZN(n5688) );
  MUX2_X1 U7260 ( .A(n5694), .B(n5688), .S(P2_IR_REG_11__SCAN_IN), .Z(n5691)
         );
  INV_X1 U7261 ( .A(n5689), .ZN(n5690) );
  OR2_X1 U7262 ( .A1(n5664), .A2(n5694), .ZN(n5692) );
  XNOR2_X1 U7263 ( .A(n5692), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6413) );
  INV_X1 U7264 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5697) );
  XNOR2_X1 U7265 ( .A(n6727), .B(n5697), .ZN(n9697) );
  INV_X1 U7266 ( .A(n5693), .ZN(n5699) );
  AND2_X1 U7267 ( .A1(n6850), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7268 ( .A1(n5693), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U7269 ( .B1(n6724), .B2(n5701), .A(n5702), .ZN(n9677) );
  INV_X1 U7270 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9676) );
  OR2_X1 U7271 ( .A1(n9677), .A2(n9676), .ZN(n9679) );
  NAND2_X1 U7272 ( .A1(n9679), .A2(n5702), .ZN(n9696) );
  NAND2_X1 U7273 ( .A1(n9697), .A2(n9696), .ZN(n9695) );
  NAND2_X1 U7274 ( .A1(n6727), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7275 ( .A1(n9695), .A2(n5703), .ZN(n5705) );
  NAND2_X1 U7276 ( .A1(n5695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  XNOR2_X1 U7277 ( .A(n5704), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6352) );
  INV_X1 U7278 ( .A(n6352), .ZN(n6896) );
  NAND2_X1 U7279 ( .A1(n5705), .A2(n6896), .ZN(n7007) );
  OAI21_X1 U7280 ( .B1(n5705), .B2(n6896), .A(n7007), .ZN(n6887) );
  INV_X1 U7281 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U7282 ( .A1(n7012), .A2(n7007), .ZN(n5708) );
  INV_X1 U7283 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5707) );
  INV_X1 U7284 ( .A(n5706), .ZN(n5711) );
  NAND2_X1 U7285 ( .A1(n5711), .A2(n5710), .ZN(n5713) );
  NAND2_X1 U7286 ( .A1(n5713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5712) );
  XNOR2_X1 U7287 ( .A(n5712), .B(n5714), .ZN(n6734) );
  NAND2_X1 U7288 ( .A1(n9730), .A2(n9728), .ZN(n5720) );
  INV_X1 U7289 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5719) );
  INV_X1 U7290 ( .A(n5713), .ZN(n5715) );
  NAND2_X1 U7291 ( .A1(n5715), .A2(n5714), .ZN(n5717) );
  NAND2_X1 U7292 ( .A1(n5717), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5716) );
  MUX2_X1 U7293 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5716), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5718) );
  MUX2_X1 U7294 ( .A(n5719), .B(P2_REG1_REG_6__SCAN_IN), .S(n9726), .Z(n9727)
         );
  INV_X1 U7295 ( .A(n9726), .ZN(n6739) );
  NAND2_X1 U7296 ( .A1(n6739), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7297 ( .A1(n5723), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5722) );
  MUX2_X1 U7298 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5722), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5724) );
  NAND2_X1 U7299 ( .A1(n5725), .A2(n7195), .ZN(n9752) );
  INV_X1 U7300 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U7301 ( .A1(n5729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U7302 ( .A(n5727), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9757) );
  MUX2_X1 U7303 ( .A(n9987), .B(P2_REG1_REG_8__SCAN_IN), .S(n9757), .Z(n9751)
         );
  INV_X1 U7304 ( .A(n9757), .ZN(n6763) );
  NAND2_X1 U7305 ( .A1(n6763), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7306 ( .A1(n9756), .A2(n5728), .ZN(n5731) );
  OAI21_X1 U7307 ( .B1(n5729), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U7308 ( .A(n5730), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6400) );
  INV_X1 U7309 ( .A(n6400), .ZN(n7587) );
  NAND2_X1 U7310 ( .A1(n5731), .A2(n7587), .ZN(n5732) );
  INV_X1 U7311 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5781) );
  AOI22_X1 U7312 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6413), .B1(n7734), .B2(
        n5781), .ZN(n7731) );
  NOR2_X1 U7313 ( .A1(n6424), .A2(n5733), .ZN(n5734) );
  INV_X1 U7314 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8070) );
  NOR2_X1 U7315 ( .A1(n8070), .A2(n8069), .ZN(n8068) );
  NAND2_X1 U7316 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6918), .ZN(n5735) );
  OAI21_X1 U7317 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6918), .A(n5735), .ZN(
        n8023) );
  NOR2_X1 U7318 ( .A1(n8024), .A2(n8023), .ZN(n8022) );
  NOR2_X1 U7319 ( .A1(n8118), .A2(n5736), .ZN(n5737) );
  INV_X1 U7320 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8055) );
  XNOR2_X1 U7321 ( .A(n5736), .B(n8118), .ZN(n8054) );
  NOR2_X1 U7322 ( .A1(n8055), .A2(n8054), .ZN(n8053) );
  NAND2_X1 U7323 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9790), .ZN(n5738) );
  OAI21_X1 U7324 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9790), .A(n5738), .ZN(
        n9775) );
  NOR2_X1 U7325 ( .A1(n8538), .A2(n5739), .ZN(n5740) );
  INV_X1 U7326 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8544) );
  INV_X1 U7327 ( .A(n8538), .ZN(n7102) );
  INV_X1 U7328 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8807) );
  AOI22_X1 U7329 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n6471), .B1(n9806), .B2(
        n8807), .ZN(n9792) );
  NOR2_X1 U7330 ( .A1(n9810), .A2(n5741), .ZN(n5742) );
  INV_X1 U7331 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U7332 ( .A1(n5743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U7333 ( .A(n5744), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8567) );
  INV_X1 U7334 ( .A(n8567), .ZN(n8558) );
  NAND2_X1 U7335 ( .A1(n8558), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U7336 ( .B1(n8558), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5745), .ZN(
        n8564) );
  INV_X1 U7337 ( .A(n5745), .ZN(n5746) );
  NOR2_X1 U7338 ( .A1(n8563), .A2(n5746), .ZN(n5747) );
  NOR2_X1 U7339 ( .A1(n8384), .A2(P2_U3151), .ZN(n8903) );
  NAND2_X1 U7340 ( .A1(n5824), .A2(n8903), .ZN(n6852) );
  INV_X1 U7341 ( .A(n6847), .ZN(n8385) );
  INV_X1 U7342 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U7343 ( .A(n6727), .B(n5748), .ZN(n9694) );
  NAND2_X1 U7344 ( .A1(n5693), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5749) );
  INV_X1 U7345 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U7346 ( .A1(n9694), .A2(n9693), .ZN(n9692) );
  NAND2_X1 U7347 ( .A1(n6727), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7348 ( .A1(n9692), .A2(n5750), .ZN(n5751) );
  NAND2_X1 U7349 ( .A1(n5751), .A2(n6896), .ZN(n7017) );
  INV_X1 U7350 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6889) );
  INV_X1 U7351 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U7352 ( .A(n7026), .B(n5752), .ZN(n7016) );
  NAND2_X1 U7353 ( .A1(n7026), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7354 ( .A1(n7021), .A2(n5753), .ZN(n5754) );
  INV_X1 U7355 ( .A(n6734), .ZN(n9710) );
  NAND2_X1 U7356 ( .A1(n9720), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U7357 ( .A1(n5754), .A2(n6734), .ZN(n5755) );
  NAND2_X1 U7358 ( .A1(n9719), .A2(n5755), .ZN(n9744) );
  INV_X1 U7359 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5756) );
  MUX2_X1 U7360 ( .A(n5756), .B(P2_REG2_REG_6__SCAN_IN), .S(n9726), .Z(n9745)
         );
  NAND2_X1 U7361 ( .A1(n9744), .A2(n9745), .ZN(n9743) );
  NAND2_X1 U7362 ( .A1(n6739), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7363 ( .A1(n9743), .A2(n5757), .ZN(n5758) );
  XNOR2_X1 U7364 ( .A(n5758), .B(n6391), .ZN(n7191) );
  NAND2_X1 U7365 ( .A1(n5758), .A2(n7195), .ZN(n5759) );
  INV_X1 U7366 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U7367 ( .A(n9983), .B(P2_REG2_REG_8__SCAN_IN), .S(n9757), .Z(n9767)
         );
  NAND2_X1 U7368 ( .A1(n6763), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7369 ( .A(n5761), .B(n6400), .ZN(n7580) );
  NAND2_X1 U7370 ( .A1(n5761), .A2(n7587), .ZN(n5762) );
  INV_X1 U7371 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U7372 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6413), .B1(n7734), .B2(
        n10008), .ZN(n7728) );
  NOR2_X1 U7373 ( .A1(n6424), .A2(n5763), .ZN(n5764) );
  INV_X1 U7374 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8067) );
  XOR2_X1 U7375 ( .A(n8073), .B(n5763), .Z(n8066) );
  NOR2_X1 U7376 ( .A1(n8067), .A2(n8066), .ZN(n8065) );
  NOR2_X1 U7377 ( .A1(n5764), .A2(n8065), .ZN(n8018) );
  NAND2_X1 U7378 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6918), .ZN(n5765) );
  OAI21_X1 U7379 ( .B1(n6918), .B2(P2_REG2_REG_12__SCAN_IN), .A(n5765), .ZN(
        n8017) );
  NOR2_X1 U7380 ( .A1(n8018), .A2(n8017), .ZN(n8016) );
  NOR2_X1 U7381 ( .A1(n8118), .A2(n5766), .ZN(n5767) );
  INV_X1 U7382 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U7383 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9790), .ZN(n5768) );
  OAI21_X1 U7384 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9790), .A(n5768), .ZN(
        n9778) );
  NOR2_X1 U7385 ( .A1(n8538), .A2(n5769), .ZN(n5770) );
  INV_X1 U7386 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10033) );
  INV_X1 U7387 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8753) );
  AOI22_X1 U7388 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6471), .B1(n9806), .B2(
        n8753), .ZN(n9794) );
  NOR2_X1 U7389 ( .A1(n9810), .A2(n5771), .ZN(n5772) );
  INV_X1 U7390 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9816) );
  INV_X1 U7391 ( .A(n9810), .ZN(n7291) );
  XOR2_X1 U7392 ( .A(n7291), .B(n5771), .Z(n9815) );
  NOR2_X1 U7393 ( .A1(n9816), .A2(n9815), .ZN(n9814) );
  NOR2_X1 U7394 ( .A1(n5772), .A2(n9814), .ZN(n8553) );
  NAND2_X1 U7395 ( .A1(n8558), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5773) );
  OAI21_X1 U7396 ( .B1(n8558), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5773), .ZN(
        n8552) );
  NOR2_X1 U7397 ( .A1(n8553), .A2(n8552), .ZN(n8551) );
  INV_X1 U7398 ( .A(n5773), .ZN(n5774) );
  NOR2_X1 U7399 ( .A1(n8551), .A2(n5774), .ZN(n5776) );
  XNOR2_X1 U7400 ( .A(n7559), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5821) );
  INV_X1 U7401 ( .A(n5821), .ZN(n5775) );
  MUX2_X1 U7402 ( .A(n9816), .B(n9813), .S(n6847), .Z(n5817) );
  XNOR2_X1 U7403 ( .A(n5817), .B(n7291), .ZN(n9821) );
  MUX2_X1 U7404 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6847), .Z(n5777) );
  OR2_X1 U7405 ( .A1(n5777), .A2(n9806), .ZN(n5815) );
  XNOR2_X1 U7406 ( .A(n5777), .B(n6471), .ZN(n9798) );
  MUX2_X1 U7407 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6847), .Z(n5778) );
  OR2_X1 U7408 ( .A1(n5778), .A2(n7102), .ZN(n5814) );
  XNOR2_X1 U7409 ( .A(n5778), .B(n8538), .ZN(n8537) );
  MUX2_X1 U7410 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6847), .Z(n5779) );
  OR2_X1 U7411 ( .A1(n5779), .A2(n9790), .ZN(n5813) );
  INV_X1 U7412 ( .A(n9790), .ZN(n6452) );
  XNOR2_X1 U7413 ( .A(n5779), .B(n6452), .ZN(n9782) );
  MUX2_X1 U7414 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6847), .Z(n5811) );
  INV_X1 U7415 ( .A(n5811), .ZN(n5780) );
  NAND2_X1 U7416 ( .A1(n8118), .A2(n5780), .ZN(n5812) );
  MUX2_X1 U7417 ( .A(n8067), .B(n8070), .S(n6847), .Z(n5806) );
  AND2_X1 U7418 ( .A1(n5806), .A2(n6424), .ZN(n5807) );
  MUX2_X1 U7419 ( .A(n10008), .B(n5781), .S(n6847), .Z(n5803) );
  AND2_X1 U7420 ( .A1(n5803), .A2(n6413), .ZN(n5804) );
  MUX2_X1 U7421 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6847), .Z(n5800) );
  INV_X1 U7422 ( .A(n5800), .ZN(n5801) );
  MUX2_X1 U7423 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6847), .Z(n5795) );
  INV_X1 U7424 ( .A(n5795), .ZN(n5796) );
  MUX2_X1 U7425 ( .A(n5752), .B(n5707), .S(n6847), .Z(n5788) );
  INV_X1 U7426 ( .A(n5788), .ZN(n5789) );
  MUX2_X1 U7427 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6847), .Z(n5787) );
  INV_X1 U7428 ( .A(n6724), .ZN(n9682) );
  XNOR2_X1 U7429 ( .A(n5785), .B(n9682), .ZN(n9688) );
  INV_X1 U7430 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5783) );
  INV_X1 U7431 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5782) );
  MUX2_X1 U7432 ( .A(n5783), .B(n5782), .S(n6847), .Z(n5784) );
  INV_X1 U7433 ( .A(n9687), .ZN(n6848) );
  OAI22_X1 U7434 ( .A1(n9688), .A2(n6848), .B1(n9682), .B2(n5785), .ZN(n9705)
         );
  MUX2_X1 U7435 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6847), .Z(n5786) );
  INV_X1 U7436 ( .A(n6727), .ZN(n9700) );
  XNOR2_X1 U7437 ( .A(n5786), .B(n9700), .ZN(n9706) );
  AOI22_X1 U7438 ( .A1(n9705), .A2(n9706), .B1(n5786), .B2(n6727), .ZN(n6884)
         );
  XNOR2_X1 U7439 ( .A(n5787), .B(n6352), .ZN(n6883) );
  NAND2_X1 U7440 ( .A1(n6884), .A2(n6883), .ZN(n6882) );
  OAI21_X1 U7441 ( .B1(n5787), .B2(n6896), .A(n6882), .ZN(n7004) );
  XOR2_X1 U7442 ( .A(n7026), .B(n5788), .Z(n7005) );
  NOR2_X1 U7443 ( .A1(n7004), .A2(n7005), .ZN(n7003) );
  MUX2_X1 U7444 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6847), .Z(n5790) );
  XNOR2_X1 U7445 ( .A(n5790), .B(n6734), .ZN(n9717) );
  INV_X1 U7446 ( .A(n5790), .ZN(n5791) );
  OAI22_X1 U7447 ( .A1(n9716), .A2(n9717), .B1(n9710), .B2(n5791), .ZN(n9741)
         );
  MUX2_X1 U7448 ( .A(n5756), .B(n5719), .S(n6847), .Z(n5792) );
  NAND2_X1 U7449 ( .A1(n5792), .A2(n9726), .ZN(n5793) );
  OAI21_X1 U7450 ( .B1(n5792), .B2(n9726), .A(n5793), .ZN(n9740) );
  NOR2_X1 U7451 ( .A1(n9741), .A2(n9740), .ZN(n9739) );
  INV_X1 U7452 ( .A(n5793), .ZN(n5794) );
  XOR2_X1 U7453 ( .A(n6391), .B(n5795), .Z(n7189) );
  NOR2_X1 U7454 ( .A1(n7190), .A2(n7189), .ZN(n7188) );
  AOI21_X1 U7455 ( .B1(n6391), .B2(n5796), .A(n7188), .ZN(n9762) );
  MUX2_X1 U7456 ( .A(n9983), .B(n9987), .S(n6847), .Z(n5797) );
  NAND2_X1 U7457 ( .A1(n5797), .A2(n9757), .ZN(n5798) );
  OAI21_X1 U7458 ( .B1(n5797), .B2(n9757), .A(n5798), .ZN(n9761) );
  NOR2_X1 U7459 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  INV_X1 U7460 ( .A(n5798), .ZN(n5799) );
  XOR2_X1 U7461 ( .A(n6400), .B(n5800), .Z(n7577) );
  NOR2_X1 U7462 ( .A1(n7578), .A2(n7577), .ZN(n7576) );
  AOI21_X1 U7463 ( .B1(n6400), .B2(n5801), .A(n7576), .ZN(n7726) );
  INV_X1 U7464 ( .A(n5804), .ZN(n5802) );
  OAI21_X1 U7465 ( .B1(n6413), .B2(n5803), .A(n5802), .ZN(n7725) );
  NOR2_X1 U7466 ( .A1(n7726), .A2(n7725), .ZN(n7724) );
  INV_X1 U7467 ( .A(n5807), .ZN(n5805) );
  OAI21_X1 U7468 ( .B1(n6424), .B2(n5806), .A(n5805), .ZN(n8076) );
  NOR2_X1 U7469 ( .A1(n8075), .A2(n8076), .ZN(n8074) );
  INV_X1 U7470 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5808) );
  INV_X1 U7471 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7961) );
  MUX2_X1 U7472 ( .A(n5808), .B(n7961), .S(n6847), .Z(n5809) );
  INV_X1 U7473 ( .A(n6918), .ZN(n8028) );
  NAND2_X1 U7474 ( .A1(n5809), .A2(n8028), .ZN(n8030) );
  MUX2_X1 U7475 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6847), .Z(n5810) );
  AND2_X1 U7476 ( .A1(n5810), .A2(n6918), .ZN(n8029) );
  AOI21_X1 U7477 ( .B1(n8033), .B2(n8030), .A(n8029), .ZN(n8061) );
  XNOR2_X1 U7478 ( .A(n5811), .B(n8118), .ZN(n8060) );
  NAND2_X1 U7479 ( .A1(n8061), .A2(n8060), .ZN(n8059) );
  NAND2_X1 U7480 ( .A1(n5812), .A2(n8059), .ZN(n9781) );
  NAND2_X1 U7481 ( .A1(n9782), .A2(n9781), .ZN(n9780) );
  NAND2_X1 U7482 ( .A1(n5814), .A2(n8535), .ZN(n9797) );
  NAND2_X1 U7483 ( .A1(n9798), .A2(n9797), .ZN(n9796) );
  NAND2_X1 U7484 ( .A1(n5815), .A2(n9796), .ZN(n9820) );
  NAND2_X1 U7485 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  INV_X1 U7486 ( .A(n9819), .ZN(n5816) );
  MUX2_X1 U7487 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6847), .Z(n5818) );
  NAND2_X1 U7488 ( .A1(n5819), .A2(n5818), .ZN(n8555) );
  OAI21_X1 U7489 ( .B1(n8554), .B2(n8567), .A(n8555), .ZN(n5823) );
  MUX2_X1 U7490 ( .A(n5821), .B(n5820), .S(n6847), .Z(n5822) );
  XNOR2_X1 U7491 ( .A(n5823), .B(n5822), .ZN(n5830) );
  INV_X1 U7492 ( .A(n8384), .ZN(n6659) );
  NOR2_X2 U7493 ( .A1(n8557), .A2(n6659), .ZN(n9822) );
  NOR2_X1 U7494 ( .A1(n6847), .A2(P2_U3151), .ZN(n8104) );
  AND2_X1 U7495 ( .A1(n5824), .A2(n8104), .ZN(n5825) );
  MUX2_X1 U7496 ( .A(P2_U3893), .B(n5825), .S(n8384), .Z(n9809) );
  NAND2_X1 U7497 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8411) );
  INV_X1 U7498 ( .A(n5826), .ZN(n7116) );
  NOR2_X1 U7499 ( .A1(n6698), .A2(n7116), .ZN(n5827) );
  NAND2_X1 U7500 ( .A1(n9808), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5828) );
  OAI211_X1 U7501 ( .C1(n9807), .C2(n7559), .A(n8411), .B(n5828), .ZN(n5829)
         );
  OAI211_X2 U7502 ( .C1(n6316), .C2(n6305), .A(n6714), .B(n9513), .ZN(n6031)
         );
  OAI22_X1 U7503 ( .A1(n9437), .A2(n5865), .B1(n8918), .B2(n6031), .ZN(n5981)
         );
  INV_X1 U7504 ( .A(n5981), .ZN(n5984) );
  NAND2_X4 U7505 ( .A1(n5835), .A2(n6714), .ZN(n6034) );
  OAI22_X1 U7506 ( .A1(n9437), .A2(n6033), .B1(n8918), .B2(n5865), .ZN(n5836)
         );
  XNOR2_X1 U7507 ( .A(n5836), .B(n6034), .ZN(n5982) );
  INV_X1 U7508 ( .A(n5982), .ZN(n5983) );
  NAND2_X1 U7509 ( .A1(n6192), .A2(n6052), .ZN(n5838) );
  NAND2_X1 U7510 ( .A1(n4290), .A2(n9548), .ZN(n5837) );
  INV_X1 U7511 ( .A(n6714), .ZN(n6046) );
  NAND2_X1 U7512 ( .A1(n6046), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7513 ( .A1(n6192), .A2(n5848), .ZN(n5842) );
  NOR2_X1 U7514 ( .A1(n6714), .A2(n4726), .ZN(n5840) );
  AOI21_X1 U7515 ( .B1(n9548), .B2(n6052), .A(n5840), .ZN(n5841) );
  NAND2_X1 U7516 ( .A1(n5842), .A2(n5841), .ZN(n6864) );
  NAND2_X1 U7517 ( .A1(n6865), .A2(n6864), .ZN(n6863) );
  AND2_X1 U7518 ( .A1(n6863), .A2(n5843), .ZN(n6955) );
  NAND2_X1 U7519 ( .A1(n9549), .A2(n4289), .ZN(n5846) );
  NAND2_X1 U7520 ( .A1(n5844), .A2(n5854), .ZN(n5845) );
  XNOR2_X1 U7521 ( .A(n5847), .B(n6034), .ZN(n5850) );
  AND2_X1 U7522 ( .A1(n9549), .A2(n6052), .ZN(n5849) );
  NAND2_X1 U7523 ( .A1(n6955), .A2(n6953), .ZN(n6954) );
  INV_X1 U7524 ( .A(n5850), .ZN(n5852) );
  NAND2_X1 U7525 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U7526 ( .A1(n6954), .A2(n5853), .ZN(n6897) );
  NAND2_X1 U7527 ( .A1(n5855), .A2(n5968), .ZN(n5858) );
  NAND2_X1 U7528 ( .A1(n5611), .A2(n5856), .ZN(n5857) );
  NAND2_X1 U7529 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  XNOR2_X1 U7530 ( .A(n5859), .B(n6034), .ZN(n5860) );
  AOI22_X1 U7531 ( .A1(n5855), .A2(n5848), .B1(n6052), .B2(n5611), .ZN(n5861)
         );
  XNOR2_X1 U7532 ( .A(n5860), .B(n5861), .ZN(n6898) );
  NAND2_X1 U7533 ( .A1(n6897), .A2(n6898), .ZN(n5864) );
  INV_X1 U7534 ( .A(n5860), .ZN(n5862) );
  NAND2_X1 U7535 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U7536 ( .A1(n5864), .A2(n5863), .ZN(n6961) );
  INV_X2 U7537 ( .A(n5865), .ZN(n5997) );
  NAND2_X1 U7538 ( .A1(n9045), .A2(n5997), .ZN(n5867) );
  NAND2_X1 U7539 ( .A1(n6963), .A2(n5856), .ZN(n5866) );
  NAND2_X1 U7540 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  XNOR2_X1 U7541 ( .A(n5868), .B(n6034), .ZN(n5870) );
  AND2_X1 U7542 ( .A1(n6963), .A2(n6052), .ZN(n5869) );
  AOI21_X1 U7543 ( .B1(n9045), .B2(n5848), .A(n5869), .ZN(n5871) );
  XNOR2_X1 U7544 ( .A(n5870), .B(n5871), .ZN(n6962) );
  NAND2_X1 U7545 ( .A1(n6961), .A2(n6962), .ZN(n7061) );
  INV_X1 U7546 ( .A(n5870), .ZN(n5872) );
  NAND2_X1 U7547 ( .A1(n5872), .A2(n5871), .ZN(n7062) );
  NAND2_X1 U7548 ( .A1(n9044), .A2(n5997), .ZN(n5874) );
  XNOR2_X1 U7549 ( .A(n7060), .B(n5876), .ZN(n5877) );
  AND2_X1 U7550 ( .A1(n7062), .A2(n5877), .ZN(n5878) );
  INV_X1 U7551 ( .A(n7060), .ZN(n5879) );
  NAND2_X1 U7552 ( .A1(n5879), .A2(n5876), .ZN(n5880) );
  NAND2_X1 U7553 ( .A1(n9043), .A2(n5997), .ZN(n5882) );
  NAND2_X1 U7554 ( .A1(n7456), .A2(n4290), .ZN(n5881) );
  NAND2_X1 U7555 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  AND2_X1 U7556 ( .A1(n5887), .A2(n5888), .ZN(n7125) );
  NAND2_X1 U7557 ( .A1(n7450), .A2(n4290), .ZN(n5885) );
  NAND2_X1 U7558 ( .A1(n9042), .A2(n5997), .ZN(n5884) );
  NAND2_X1 U7559 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  XNOR2_X1 U7560 ( .A(n5886), .B(n6050), .ZN(n5893) );
  AOI22_X1 U7561 ( .A1(n7450), .A2(n5997), .B1(n5848), .B2(n9042), .ZN(n5892)
         );
  XNOR2_X1 U7562 ( .A(n5893), .B(n5892), .ZN(n7166) );
  NAND2_X1 U7563 ( .A1(n9043), .A2(n5848), .ZN(n5891) );
  NAND2_X1 U7564 ( .A1(n7456), .A2(n5997), .ZN(n5890) );
  NAND2_X1 U7565 ( .A1(n5891), .A2(n5890), .ZN(n7127) );
  NAND2_X1 U7566 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7567 ( .A1(n5899), .A2(n5856), .ZN(n5896) );
  NAND2_X1 U7568 ( .A1(n9041), .A2(n5997), .ZN(n5895) );
  NAND2_X1 U7569 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  XNOR2_X1 U7570 ( .A(n5897), .B(n6050), .ZN(n7177) );
  AND2_X1 U7571 ( .A1(n9041), .A2(n5848), .ZN(n5898) );
  AOI21_X1 U7572 ( .B1(n5899), .B2(n5997), .A(n5898), .ZN(n7178) );
  AND2_X1 U7573 ( .A1(n7177), .A2(n7178), .ZN(n5900) );
  NAND2_X1 U7574 ( .A1(n7495), .A2(n5856), .ZN(n5902) );
  NAND2_X1 U7575 ( .A1(n9040), .A2(n5997), .ZN(n5901) );
  NAND2_X1 U7576 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  XNOR2_X1 U7577 ( .A(n5903), .B(n6034), .ZN(n5904) );
  NAND2_X1 U7578 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  AND2_X1 U7579 ( .A1(n9040), .A2(n5848), .ZN(n5907) );
  AOI21_X1 U7580 ( .B1(n7495), .B2(n5997), .A(n5907), .ZN(n7401) );
  NAND2_X1 U7581 ( .A1(n9608), .A2(n5856), .ZN(n5909) );
  NAND2_X1 U7582 ( .A1(n9039), .A2(n5997), .ZN(n5908) );
  NAND2_X1 U7583 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  XNOR2_X1 U7584 ( .A(n5910), .B(n6034), .ZN(n5927) );
  INV_X1 U7585 ( .A(n5927), .ZN(n5914) );
  NAND2_X1 U7586 ( .A1(n9608), .A2(n5968), .ZN(n5912) );
  NAND2_X1 U7587 ( .A1(n9039), .A2(n5848), .ZN(n5911) );
  NAND2_X1 U7588 ( .A1(n5912), .A2(n5911), .ZN(n5926) );
  INV_X1 U7589 ( .A(n5926), .ZN(n5913) );
  NAND2_X1 U7590 ( .A1(n5914), .A2(n5913), .ZN(n7477) );
  AND2_X1 U7591 ( .A1(n7476), .A2(n7477), .ZN(n5915) );
  NAND2_X1 U7592 ( .A1(n7536), .A2(n5856), .ZN(n5917) );
  NAND2_X1 U7593 ( .A1(n9037), .A2(n5968), .ZN(n5916) );
  NAND2_X1 U7594 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  XNOR2_X1 U7595 ( .A(n5918), .B(n6034), .ZN(n7855) );
  NAND2_X1 U7596 ( .A1(n7536), .A2(n5968), .ZN(n5920) );
  NAND2_X1 U7597 ( .A1(n9037), .A2(n5848), .ZN(n5919) );
  NAND2_X1 U7598 ( .A1(n5920), .A2(n5919), .ZN(n5933) );
  NAND2_X1 U7599 ( .A1(n7751), .A2(n4290), .ZN(n5922) );
  NAND2_X1 U7600 ( .A1(n9038), .A2(n5968), .ZN(n5921) );
  NAND2_X1 U7601 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  XNOR2_X1 U7602 ( .A(n5923), .B(n6034), .ZN(n5930) );
  NAND2_X1 U7603 ( .A1(n7751), .A2(n5968), .ZN(n5925) );
  NAND2_X1 U7604 ( .A1(n9038), .A2(n5848), .ZN(n5924) );
  NAND2_X1 U7605 ( .A1(n5925), .A2(n5924), .ZN(n7745) );
  AOI22_X1 U7606 ( .A1(n7855), .A2(n5933), .B1(n5930), .B2(n7745), .ZN(n5928)
         );
  NAND2_X1 U7607 ( .A1(n5927), .A2(n5926), .ZN(n7743) );
  AND2_X1 U7608 ( .A1(n5928), .A2(n7743), .ZN(n5929) );
  NAND2_X1 U7609 ( .A1(n7744), .A2(n5929), .ZN(n5938) );
  INV_X1 U7610 ( .A(n7855), .ZN(n5936) );
  INV_X1 U7611 ( .A(n5930), .ZN(n7853) );
  INV_X1 U7612 ( .A(n7745), .ZN(n5931) );
  NAND2_X1 U7613 ( .A1(n7853), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U7614 ( .A1(n5932), .A2(n5933), .ZN(n5935) );
  INV_X1 U7615 ( .A(n5932), .ZN(n5934) );
  INV_X1 U7616 ( .A(n5933), .ZN(n7854) );
  AOI22_X1 U7617 ( .A1(n5936), .A2(n5935), .B1(n5934), .B2(n7854), .ZN(n5937)
         );
  NAND2_X1 U7618 ( .A1(n5938), .A2(n5937), .ZN(n7656) );
  NAND2_X1 U7619 ( .A1(n7663), .A2(n4290), .ZN(n5940) );
  NAND2_X1 U7620 ( .A1(n7545), .A2(n5968), .ZN(n5939) );
  NAND2_X1 U7621 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  XNOR2_X1 U7622 ( .A(n5941), .B(n6034), .ZN(n5943) );
  AND2_X1 U7623 ( .A1(n7545), .A2(n5848), .ZN(n5942) );
  AOI21_X1 U7624 ( .B1(n7663), .B2(n6052), .A(n5942), .ZN(n5944) );
  XNOR2_X1 U7625 ( .A(n5943), .B(n5944), .ZN(n7657) );
  INV_X1 U7626 ( .A(n5943), .ZN(n5945) );
  NAND2_X1 U7627 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7628 ( .A1(n5951), .A2(n5856), .ZN(n5948) );
  NAND2_X1 U7629 ( .A1(n9036), .A2(n5968), .ZN(n5947) );
  NAND2_X1 U7630 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  XNOR2_X1 U7631 ( .A(n5949), .B(n6034), .ZN(n5952) );
  AND2_X1 U7632 ( .A1(n9036), .A2(n5848), .ZN(n5950) );
  AOI21_X1 U7633 ( .B1(n5951), .B2(n6052), .A(n5950), .ZN(n5953) );
  XNOR2_X1 U7634 ( .A(n5952), .B(n5953), .ZN(n7706) );
  INV_X1 U7635 ( .A(n5952), .ZN(n5954) );
  NAND2_X1 U7636 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7637 ( .A1(n9640), .A2(n4290), .ZN(n5958) );
  NAND2_X1 U7638 ( .A1(n9035), .A2(n5968), .ZN(n5957) );
  NAND2_X1 U7639 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7640 ( .A(n5959), .B(n6050), .ZN(n5960) );
  AOI22_X1 U7641 ( .A1(n9640), .A2(n5997), .B1(n5848), .B2(n9035), .ZN(n7944)
         );
  NAND2_X1 U7642 ( .A1(n7835), .A2(n5856), .ZN(n5962) );
  NAND2_X1 U7643 ( .A1(n9034), .A2(n5997), .ZN(n5961) );
  NAND2_X1 U7644 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  XNOR2_X1 U7645 ( .A(n5963), .B(n6034), .ZN(n5965) );
  XNOR2_X1 U7646 ( .A(n5964), .B(n5965), .ZN(n9006) );
  AOI22_X1 U7647 ( .A1(n7835), .A2(n5997), .B1(n5848), .B2(n9034), .ZN(n9005)
         );
  INV_X1 U7648 ( .A(n5964), .ZN(n7947) );
  INV_X1 U7649 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7650 ( .A1(n8946), .A2(n5856), .ZN(n5970) );
  NAND2_X1 U7651 ( .A1(n9033), .A2(n5968), .ZN(n5969) );
  NAND2_X1 U7652 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  XNOR2_X1 U7653 ( .A(n5971), .B(n6034), .ZN(n5972) );
  AOI22_X1 U7654 ( .A1(n8946), .A2(n5997), .B1(n5848), .B2(n9033), .ZN(n5973)
         );
  XNOR2_X1 U7655 ( .A(n5972), .B(n5973), .ZN(n8941) );
  INV_X1 U7656 ( .A(n5972), .ZN(n5974) );
  AOI22_X1 U7657 ( .A1(n7933), .A2(n5997), .B1(n5848), .B2(n9032), .ZN(n5977)
         );
  AOI22_X1 U7658 ( .A1(n7933), .A2(n5856), .B1(n6052), .B2(n9032), .ZN(n5975)
         );
  XNOR2_X1 U7659 ( .A(n5975), .B(n6034), .ZN(n5976) );
  XOR2_X1 U7660 ( .A(n5977), .B(n5976), .Z(n8950) );
  INV_X1 U7661 ( .A(n5976), .ZN(n5979) );
  NAND2_X1 U7662 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7663 ( .A(n5982), .B(n5981), .ZN(n8981) );
  AOI22_X1 U7664 ( .A1(n9380), .A2(n5997), .B1(n5848), .B2(n9030), .ZN(n5988)
         );
  NAND2_X1 U7665 ( .A1(n9380), .A2(n4290), .ZN(n5986) );
  NAND2_X1 U7666 ( .A1(n9030), .A2(n5997), .ZN(n5985) );
  NAND2_X1 U7667 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  XNOR2_X1 U7668 ( .A(n5987), .B(n6034), .ZN(n5990) );
  XOR2_X1 U7669 ( .A(n5988), .B(n5990), .Z(n8917) );
  INV_X1 U7670 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7671 ( .A1(n9377), .A2(n4290), .ZN(n5992) );
  NAND2_X1 U7672 ( .A1(n8926), .A2(n5997), .ZN(n5991) );
  NAND2_X1 U7673 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  XNOR2_X1 U7674 ( .A(n5993), .B(n6034), .ZN(n5994) );
  AOI22_X1 U7675 ( .A1(n9377), .A2(n6052), .B1(n5848), .B2(n8926), .ZN(n5995)
         );
  XNOR2_X1 U7676 ( .A(n5994), .B(n5995), .ZN(n8965) );
  INV_X1 U7677 ( .A(n5994), .ZN(n5996) );
  AOI22_X1 U7678 ( .A1(n9427), .A2(n6052), .B1(n5848), .B2(n9029), .ZN(n6001)
         );
  NAND2_X1 U7679 ( .A1(n9427), .A2(n5856), .ZN(n5999) );
  NAND2_X1 U7680 ( .A1(n9029), .A2(n5997), .ZN(n5998) );
  NAND2_X1 U7681 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  XNOR2_X1 U7682 ( .A(n6000), .B(n6034), .ZN(n6003) );
  XOR2_X1 U7683 ( .A(n6001), .B(n6003), .Z(n8924) );
  INV_X1 U7684 ( .A(n6001), .ZN(n6002) );
  OR2_X1 U7685 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7686 ( .A1(n6008), .A2(n4290), .ZN(n6006) );
  NAND2_X1 U7687 ( .A1(n9028), .A2(n5968), .ZN(n6005) );
  NAND2_X1 U7688 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  XNOR2_X1 U7689 ( .A(n6007), .B(n6034), .ZN(n6010) );
  AOI22_X1 U7690 ( .A1(n6008), .A2(n5997), .B1(n5848), .B2(n9028), .ZN(n8974)
         );
  NAND2_X1 U7691 ( .A1(n8973), .A2(n8974), .ZN(n8972) );
  INV_X1 U7692 ( .A(n6009), .ZN(n6011) );
  NAND2_X1 U7693 ( .A1(n9235), .A2(n4290), .ZN(n6014) );
  NAND2_X1 U7694 ( .A1(n9027), .A2(n5997), .ZN(n6013) );
  NAND2_X1 U7695 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  XNOR2_X1 U7696 ( .A(n6015), .B(n6034), .ZN(n6016) );
  AOI22_X1 U7697 ( .A1(n9235), .A2(n6052), .B1(n5848), .B2(n9027), .ZN(n6017)
         );
  XNOR2_X1 U7698 ( .A(n6016), .B(n6017), .ZN(n8910) );
  INV_X1 U7699 ( .A(n6016), .ZN(n6018) );
  AOI22_X1 U7700 ( .A1(n9354), .A2(n6052), .B1(n5848), .B2(n9026), .ZN(n6022)
         );
  NAND2_X1 U7701 ( .A1(n9354), .A2(n4290), .ZN(n6020) );
  NAND2_X1 U7702 ( .A1(n9026), .A2(n5997), .ZN(n6019) );
  NAND2_X1 U7703 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7704 ( .A(n6021), .B(n6034), .ZN(n6024) );
  XOR2_X1 U7705 ( .A(n6022), .B(n6024), .Z(n8957) );
  INV_X1 U7706 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7707 ( .A1(n9348), .A2(n5856), .ZN(n6026) );
  NAND2_X1 U7708 ( .A1(n9025), .A2(n5997), .ZN(n6025) );
  NAND2_X1 U7709 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7710 ( .A(n6027), .B(n6034), .ZN(n6028) );
  AOI22_X1 U7711 ( .A1(n9348), .A2(n5968), .B1(n5848), .B2(n9025), .ZN(n6029)
         );
  XNOR2_X1 U7712 ( .A(n6028), .B(n6029), .ZN(n8934) );
  INV_X1 U7713 ( .A(n6028), .ZN(n6030) );
  OAI22_X1 U7714 ( .A1(n9413), .A2(n5865), .B1(n6032), .B2(n6031), .ZN(n6037)
         );
  OAI22_X1 U7715 ( .A1(n9413), .A2(n6033), .B1(n6032), .B2(n5865), .ZN(n6035)
         );
  XNOR2_X1 U7716 ( .A(n6035), .B(n6034), .ZN(n6036) );
  XOR2_X1 U7717 ( .A(n6037), .B(n6036), .Z(n8991) );
  NAND2_X1 U7718 ( .A1(n6036), .A2(n6037), .ZN(n6038) );
  AND2_X1 U7719 ( .A1(n9023), .A2(n5848), .ZN(n6039) );
  AOI21_X1 U7720 ( .B1(n9178), .B2(n5968), .A(n6039), .ZN(n6055) );
  NAND2_X1 U7721 ( .A1(n9178), .A2(n5856), .ZN(n6041) );
  NAND2_X1 U7722 ( .A1(n9023), .A2(n5997), .ZN(n6040) );
  NAND2_X1 U7723 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  XNOR2_X1 U7724 ( .A(n6042), .B(n6034), .ZN(n6057) );
  NAND3_X1 U7725 ( .A1(n6044), .A2(n7311), .A3(n6043), .ZN(n6064) );
  OR2_X1 U7726 ( .A1(n6064), .A2(n6740), .ZN(n6060) );
  NAND2_X1 U7727 ( .A1(n9632), .A2(n6742), .ZN(n6047) );
  NAND2_X1 U7728 ( .A1(n9404), .A2(n5856), .ZN(n6049) );
  NAND2_X1 U7729 ( .A1(n9022), .A2(n5968), .ZN(n6048) );
  NAND2_X1 U7730 ( .A1(n6049), .A2(n6048), .ZN(n6051) );
  XNOR2_X1 U7731 ( .A(n6051), .B(n6050), .ZN(n6054) );
  AOI22_X1 U7732 ( .A1(n9404), .A2(n6052), .B1(n5848), .B2(n9022), .ZN(n6053)
         );
  XNOR2_X1 U7733 ( .A(n6054), .B(n6053), .ZN(n6070) );
  INV_X1 U7734 ( .A(n6055), .ZN(n6056) );
  OR2_X1 U7735 ( .A1(n6057), .A2(n6056), .ZN(n6067) );
  NAND4_X1 U7736 ( .A1(n6705), .A2(n9007), .A3(n6070), .A4(n6067), .ZN(n6075)
         );
  INV_X1 U7737 ( .A(n6060), .ZN(n6059) );
  OR2_X1 U7738 ( .A1(n6842), .A2(n7684), .ZN(n7321) );
  INV_X1 U7739 ( .A(n7321), .ZN(n6058) );
  AOI21_X2 U7740 ( .B1(n6059), .B2(n6058), .A(n9542), .ZN(n9017) );
  AOI22_X1 U7741 ( .A1(n9023), .A2(n8982), .B1(n8983), .B2(n9021), .ZN(n9153)
         );
  NOR2_X2 U7742 ( .A1(n6060), .A2(n6305), .ZN(n9001) );
  INV_X1 U7743 ( .A(n6061), .ZN(n6063) );
  AOI21_X1 U7744 ( .B1(n6064), .B2(n6063), .A(n6062), .ZN(n6065) );
  AOI22_X1 U7745 ( .A1(n9164), .A2(n9013), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6066) );
  OAI21_X1 U7746 ( .B1(n9153), .B2(n9011), .A(n6066), .ZN(n6069) );
  NOR3_X1 U7747 ( .A1(n6070), .A2(n8988), .A3(n6067), .ZN(n6068) );
  AOI211_X1 U7748 ( .C1(n9404), .C2(n8968), .A(n6069), .B(n6068), .ZN(n6074)
         );
  INV_X1 U7749 ( .A(n6705), .ZN(n6072) );
  INV_X1 U7750 ( .A(n6070), .ZN(n6071) );
  NAND3_X1 U7751 ( .A1(n6075), .A2(n6074), .A3(n6073), .ZN(P1_U3220) );
  INV_X1 U7752 ( .A(n6076), .ZN(n6077) );
  MUX2_X1 U7753 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6722), .Z(n6081) );
  XNOR2_X1 U7754 ( .A(n6081), .B(SI_30_), .ZN(n6180) );
  OAI22_X1 U7755 ( .A1(n6181), .A2(n6180), .B1(SI_30_), .B2(n6081), .ZN(n6085)
         );
  INV_X1 U7756 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6082) );
  INV_X1 U7757 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U7758 ( .A(n6082), .B(n8315), .S(n6722), .Z(n6083) );
  XNOR2_X1 U7759 ( .A(n6083), .B(SI_31_), .ZN(n6084) );
  XNOR2_X1 U7760 ( .A(n6085), .B(n6084), .ZN(n8314) );
  MUX2_X1 U7761 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8314), .S(n6717), .Z(n6086) );
  INV_X1 U7762 ( .A(n6191), .ZN(n9020) );
  NAND2_X1 U7763 ( .A1(n6087), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7764 ( .A1(n4288), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7765 ( .A1(n6088), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6089) );
  AND3_X1 U7766 ( .A1(n6091), .A2(n6090), .A3(n6089), .ZN(n9125) );
  INV_X1 U7767 ( .A(n9125), .ZN(n9019) );
  OAI21_X1 U7768 ( .B1(n9398), .B2(n9020), .A(n9019), .ZN(n6188) );
  INV_X1 U7769 ( .A(n6155), .ZN(n6235) );
  NAND2_X1 U7770 ( .A1(n6135), .A2(n6092), .ZN(n6094) );
  OR2_X1 U7771 ( .A1(n7835), .A2(n6307), .ZN(n6093) );
  NAND2_X1 U7772 ( .A1(n6094), .A2(n6093), .ZN(n6140) );
  AOI211_X1 U7773 ( .C1(n4710), .C2(n6098), .A(n4712), .B(n9504), .ZN(n6097)
         );
  NOR2_X1 U7774 ( .A1(n9505), .A2(n9504), .ZN(n9503) );
  NAND2_X1 U7775 ( .A1(n7502), .A2(n6100), .ZN(n6102) );
  MUX2_X1 U7776 ( .A(n6102), .B(n6101), .S(n6307), .Z(n6103) );
  AOI21_X1 U7777 ( .B1(n9503), .B2(n6307), .A(n6103), .ZN(n6104) );
  NAND2_X1 U7778 ( .A1(n6105), .A2(n6104), .ZN(n6110) );
  NAND2_X1 U7779 ( .A1(n6112), .A2(n7501), .ZN(n6106) );
  MUX2_X1 U7780 ( .A(n6107), .B(n6106), .S(n6096), .Z(n6108) );
  INV_X1 U7781 ( .A(n6108), .ZN(n6109) );
  NAND2_X1 U7782 ( .A1(n6128), .A2(n6125), .ZN(n6114) );
  OR2_X1 U7783 ( .A1(n6114), .A2(n6111), .ZN(n6260) );
  AND2_X1 U7784 ( .A1(n6126), .A2(n7528), .ZN(n6113) );
  OR2_X1 U7785 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  NAND2_X1 U7786 ( .A1(n6115), .A2(n6127), .ZN(n6272) );
  INV_X1 U7787 ( .A(n6120), .ZN(n6123) );
  INV_X1 U7788 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7789 ( .A1(n6129), .A2(n6273), .ZN(n6134) );
  INV_X1 U7790 ( .A(n6276), .ZN(n6130) );
  NAND2_X1 U7791 ( .A1(n6132), .A2(n6131), .ZN(n6259) );
  AOI21_X1 U7792 ( .B1(n6134), .B2(n6133), .A(n6259), .ZN(n6137) );
  INV_X1 U7793 ( .A(n6135), .ZN(n6136) );
  AOI21_X1 U7794 ( .B1(n6137), .B2(n6118), .A(n6136), .ZN(n6138) );
  MUX2_X1 U7795 ( .A(n6139), .B(n6138), .S(n6096), .Z(n6142) );
  NAND3_X1 U7796 ( .A1(n6140), .A2(n6118), .A3(n9034), .ZN(n6141) );
  AOI21_X1 U7797 ( .B1(n6142), .B2(n6141), .A(n6208), .ZN(n6147) );
  INV_X1 U7798 ( .A(n6144), .ZN(n6152) );
  NAND2_X1 U7799 ( .A1(n6146), .A2(n6145), .ZN(n6282) );
  NOR2_X1 U7800 ( .A1(n6147), .A2(n6282), .ZN(n6150) );
  NAND2_X1 U7801 ( .A1(n6153), .A2(n6148), .ZN(n6258) );
  OAI211_X1 U7802 ( .C1(n6150), .C2(n6258), .A(n6158), .B(n6149), .ZN(n6151)
         );
  MUX2_X1 U7803 ( .A(n6152), .B(n6151), .S(n6307), .Z(n6157) );
  AOI21_X1 U7804 ( .B1(n6154), .B2(n6153), .A(n6307), .ZN(n6156) );
  AND2_X1 U7805 ( .A1(n6155), .A2(n6154), .ZN(n6225) );
  NAND2_X1 U7806 ( .A1(n6159), .A2(n6158), .ZN(n6230) );
  OR2_X1 U7807 ( .A1(n9235), .A2(n6164), .ZN(n6161) );
  NAND2_X1 U7808 ( .A1(n6218), .A2(n6162), .ZN(n6231) );
  AOI22_X1 U7809 ( .A1(n6163), .A2(n6218), .B1(n6231), .B2(n6307), .ZN(n6166)
         );
  NOR3_X1 U7810 ( .A1(n9235), .A2(n6164), .A3(n6096), .ZN(n6165) );
  INV_X1 U7811 ( .A(n6233), .ZN(n6168) );
  INV_X1 U7812 ( .A(n6221), .ZN(n6167) );
  MUX2_X1 U7813 ( .A(n6168), .B(n6167), .S(n6096), .Z(n6169) );
  INV_X1 U7814 ( .A(n6224), .ZN(n6170) );
  AOI21_X1 U7815 ( .B1(n6177), .B2(n6171), .A(n6170), .ZN(n6173) );
  INV_X1 U7816 ( .A(n6288), .ZN(n6176) );
  NAND2_X1 U7817 ( .A1(n6291), .A2(n6228), .ZN(n6240) );
  INV_X1 U7818 ( .A(n6240), .ZN(n6172) );
  INV_X1 U7819 ( .A(n9149), .ZN(n6174) );
  MUX2_X1 U7820 ( .A(n6244), .B(n6189), .S(n6096), .Z(n6178) );
  NAND2_X1 U7821 ( .A1(n8898), .A2(n6182), .ZN(n6185) );
  INV_X1 U7822 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6183) );
  OR2_X1 U7823 ( .A1(n5184), .A2(n6183), .ZN(n6184) );
  OR2_X1 U7824 ( .A1(n9401), .A2(n6191), .ZN(n6248) );
  NAND2_X1 U7825 ( .A1(n6308), .A2(n6248), .ZN(n6300) );
  INV_X1 U7826 ( .A(n6244), .ZN(n6216) );
  NAND2_X1 U7827 ( .A1(n9398), .A2(n9019), .ZN(n6301) );
  INV_X1 U7828 ( .A(n6189), .ZN(n6190) );
  AOI21_X1 U7829 ( .B1(n9401), .B2(n6191), .A(n6190), .ZN(n6257) );
  NAND2_X1 U7830 ( .A1(n6301), .A2(n6257), .ZN(n6245) );
  INV_X1 U7831 ( .A(n7643), .ZN(n6206) );
  INV_X1 U7832 ( .A(n9535), .ZN(n6193) );
  NAND2_X1 U7833 ( .A1(n6192), .A2(n6841), .ZN(n6262) );
  AND2_X1 U7834 ( .A1(n6193), .A2(n6262), .ZN(n7351) );
  NAND4_X1 U7835 ( .A1(n6195), .A2(n7351), .A3(n6194), .A4(n7723), .ZN(n6196)
         );
  NOR2_X1 U7836 ( .A1(n6196), .A2(n9528), .ZN(n6199) );
  NAND4_X1 U7837 ( .A1(n6199), .A2(n6198), .A3(n7316), .A4(n6197), .ZN(n6200)
         );
  NOR3_X1 U7838 ( .A1(n7376), .A2(n6201), .A3(n6200), .ZN(n6202) );
  NAND4_X1 U7839 ( .A1(n7466), .A2(n7527), .A3(n6203), .A4(n6202), .ZN(n6204)
         );
  NOR2_X1 U7840 ( .A1(n7551), .A2(n6204), .ZN(n6205) );
  NAND4_X1 U7841 ( .A1(n7815), .A2(n7833), .A3(n6206), .A4(n6205), .ZN(n6207)
         );
  NOR2_X1 U7842 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND3_X1 U7843 ( .A1(n9298), .A2(n9309), .A3(n6209), .ZN(n6210) );
  NOR2_X1 U7844 ( .A1(n9276), .A2(n6210), .ZN(n6211) );
  NAND4_X1 U7845 ( .A1(n9233), .A2(n9248), .A3(n9261), .A4(n6211), .ZN(n6212)
         );
  OR3_X1 U7846 ( .A1(n9203), .A2(n9220), .A3(n6212), .ZN(n6214) );
  OR4_X1 U7847 ( .A1(n6214), .A2(n9156), .A3(n6213), .A4(n9190), .ZN(n6215) );
  INV_X1 U7848 ( .A(n6217), .ZN(n6219) );
  NAND2_X1 U7849 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7850 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  NAND2_X1 U7851 ( .A1(n6222), .A2(n6233), .ZN(n6223) );
  AND2_X1 U7852 ( .A1(n6224), .A2(n6223), .ZN(n6238) );
  INV_X1 U7853 ( .A(n6238), .ZN(n6227) );
  INV_X1 U7854 ( .A(n6225), .ZN(n6226) );
  NOR2_X1 U7855 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  NAND2_X1 U7856 ( .A1(n6229), .A2(n6228), .ZN(n6290) );
  OAI21_X1 U7857 ( .B1(n6290), .B2(n9280), .A(n6288), .ZN(n6243) );
  INV_X1 U7858 ( .A(n6230), .ZN(n6234) );
  INV_X1 U7859 ( .A(n6231), .ZN(n6232) );
  OAI211_X1 U7860 ( .C1(n6235), .C2(n6234), .A(n6233), .B(n6232), .ZN(n6237)
         );
  AOI21_X1 U7861 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(n6239) );
  NOR2_X1 U7862 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  OR2_X1 U7863 ( .A1(n6242), .A2(n6241), .ZN(n6294) );
  AOI21_X1 U7864 ( .B1(n6291), .B2(n6243), .A(n6294), .ZN(n6247) );
  NAND2_X1 U7865 ( .A1(n6244), .A2(n9149), .ZN(n6296) );
  INV_X1 U7866 ( .A(n6245), .ZN(n6246) );
  OAI21_X1 U7867 ( .B1(n6247), .B2(n6296), .A(n6246), .ZN(n6252) );
  INV_X1 U7868 ( .A(n6248), .ZN(n6250) );
  INV_X1 U7869 ( .A(n9398), .ZN(n6249) );
  OAI21_X1 U7870 ( .B1(n9125), .B2(n6250), .A(n6249), .ZN(n6251) );
  AOI22_X1 U7871 ( .A1(n6252), .A2(n6251), .B1(n9398), .B2(n9401), .ZN(n6254)
         );
  OAI21_X1 U7872 ( .B1(n6254), .B2(n6742), .A(n6253), .ZN(n6255) );
  NOR2_X1 U7873 ( .A1(n6256), .A2(n7684), .ZN(n6321) );
  INV_X1 U7874 ( .A(n6257), .ZN(n6298) );
  INV_X1 U7875 ( .A(n6258), .ZN(n6287) );
  INV_X1 U7876 ( .A(n6259), .ZN(n6279) );
  INV_X1 U7877 ( .A(n6260), .ZN(n6271) );
  INV_X1 U7878 ( .A(n9549), .ZN(n9561) );
  AOI21_X1 U7879 ( .B1(n9047), .B2(n9561), .A(n7723), .ZN(n6264) );
  NAND4_X1 U7880 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n6268)
         );
  INV_X1 U7881 ( .A(n6266), .ZN(n6267) );
  OAI21_X1 U7882 ( .B1(n4713), .B2(n6268), .A(n6267), .ZN(n6269) );
  NAND3_X1 U7883 ( .A1(n6271), .A2(n6270), .A3(n6269), .ZN(n6275) );
  INV_X1 U7884 ( .A(n6272), .ZN(n6274) );
  NAND3_X1 U7885 ( .A1(n6275), .A2(n6274), .A3(n6273), .ZN(n6277) );
  NAND3_X1 U7886 ( .A1(n6277), .A2(n7828), .A3(n6276), .ZN(n6278) );
  NAND2_X1 U7887 ( .A1(n6279), .A2(n6278), .ZN(n6281) );
  AOI21_X1 U7888 ( .B1(n4898), .B2(n6281), .A(n6280), .ZN(n6284) );
  INV_X1 U7889 ( .A(n6282), .ZN(n6283) );
  OAI21_X1 U7890 ( .B1(n4904), .B2(n6284), .A(n6283), .ZN(n6286) );
  AOI21_X1 U7891 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(n6289) );
  OAI21_X1 U7892 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6292) );
  AND2_X1 U7893 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NOR2_X1 U7894 ( .A1(n6294), .A2(n6293), .ZN(n6295) );
  NOR2_X1 U7895 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  NOR2_X1 U7896 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  OR2_X1 U7897 ( .A1(n6300), .A2(n6299), .ZN(n6302) );
  NAND2_X1 U7898 ( .A1(n6302), .A2(n6301), .ZN(n6306) );
  NAND3_X1 U7899 ( .A1(n6306), .A2(n9119), .A3(n7684), .ZN(n6304) );
  NAND2_X1 U7900 ( .A1(n6741), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7896) );
  INV_X1 U7901 ( .A(n7896), .ZN(n6303) );
  OAI211_X1 U7902 ( .C1(n6306), .C2(n6305), .A(n6304), .B(n6303), .ZN(n6320)
         );
  NOR2_X1 U7903 ( .A1(n6308), .A2(n6307), .ZN(n6311) );
  NOR4_X1 U7904 ( .A1(n7896), .A2(n6316), .A3(n7723), .A4(n7684), .ZN(n6310)
         );
  NAND3_X1 U7905 ( .A1(n9398), .A2(n9119), .A3(n9019), .ZN(n6309) );
  OAI211_X1 U7906 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n6309), .ZN(n6318)
         );
  NOR4_X1 U7907 ( .A1(n5834), .A2(n6313), .A3(n5605), .A4(n4294), .ZN(n6314)
         );
  NAND2_X1 U7908 ( .A1(n6314), .A2(n9441), .ZN(n6315) );
  OAI211_X1 U7909 ( .C1(n6316), .C2(n7896), .A(n6315), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6317) );
  OAI21_X1 U7910 ( .B1(n6321), .B2(n6320), .A(n6319), .ZN(P1_U3242) );
  INV_X1 U7911 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U7912 ( .A1(n6376), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6334) );
  AND2_X4 U7913 ( .A1(n8902), .A2(n6329), .ZN(n8318) );
  NAND2_X1 U7914 ( .A1(n8318), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7915 ( .A1(n4297), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7916 ( .A1(n6346), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7917 ( .A1(n6351), .A2(n6725), .ZN(n6335) );
  OAI211_X1 U7918 ( .C1(n6661), .C2(n6727), .A(n6336), .B(n6335), .ZN(n7034)
         );
  NAND2_X1 U7919 ( .A1(n7033), .A2(n7034), .ZN(n8193) );
  INV_X1 U7920 ( .A(n7033), .ZN(n7138) );
  NAND2_X1 U7921 ( .A1(n7138), .A2(n9854), .ZN(n8189) );
  NAND2_X1 U7922 ( .A1(n6346), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7923 ( .A1(n8318), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7924 ( .A1(n4297), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7925 ( .A1(n6376), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7926 ( .A1(n6722), .A2(SI_0_), .ZN(n6341) );
  XNOR2_X1 U7927 ( .A(n6341), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U7928 ( .A1(n4295), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6344) );
  NOR2_X1 U7929 ( .A1(n6342), .A2(n4897), .ZN(n6343) );
  OR2_X2 U7930 ( .A1(n6615), .A2(n6992), .ZN(n8183) );
  NAND2_X1 U7931 ( .A1(n4293), .A2(n6992), .ZN(n8184) );
  NAND2_X2 U7932 ( .A1(n8183), .A2(n8184), .ZN(n8346) );
  NAND2_X1 U7933 ( .A1(n8318), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7934 ( .A1(n6376), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7935 ( .A1(n4298), .A2(n7233), .ZN(n6348) );
  NAND2_X1 U7936 ( .A1(n6346), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6347) );
  OR2_X1 U7937 ( .A1(n6351), .A2(n6730), .ZN(n6354) );
  NAND2_X1 U7938 ( .A1(n6499), .A2(n6352), .ZN(n6353) );
  OR2_X1 U7939 ( .A1(n9842), .A2(n7224), .ZN(n8216) );
  NAND2_X1 U7940 ( .A1(n9842), .A2(n7224), .ZN(n8199) );
  INV_X1 U7941 ( .A(n8343), .ZN(n7215) );
  NAND2_X1 U7942 ( .A1(n7212), .A2(n7215), .ZN(n7211) );
  NAND2_X1 U7943 ( .A1(n7211), .A2(n8216), .ZN(n7208) );
  NAND2_X1 U7944 ( .A1(n6376), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7945 ( .A1(n8318), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6363) );
  NOR2_X1 U7946 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6366) );
  INV_X1 U7947 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U7948 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6357) );
  NAND2_X1 U7949 ( .A1(n6367), .A2(n6357), .ZN(n7115) );
  NAND2_X1 U7950 ( .A1(n4297), .A2(n7115), .ZN(n6361) );
  NAND2_X1 U7951 ( .A1(n6346), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6360) );
  NAND4_X1 U7952 ( .A1(n6362), .A2(n6363), .A3(n6361), .A4(n6360), .ZN(n8531)
         );
  OR2_X1 U7953 ( .A1(n6351), .A2(n6735), .ZN(n6358) );
  OAI211_X1 U7954 ( .C1(n6661), .C2(n7026), .A(n6359), .B(n6358), .ZN(n7118)
         );
  NAND2_X1 U7955 ( .A1(n8531), .A2(n9863), .ZN(n8217) );
  NAND2_X1 U7956 ( .A1(n7147), .A2(n7118), .ZN(n8200) );
  NAND2_X1 U7957 ( .A1(n7208), .A2(n6618), .ZN(n6364) );
  NAND2_X1 U7958 ( .A1(n6364), .A2(n8200), .ZN(n7254) );
  NAND2_X1 U7959 ( .A1(n6346), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7960 ( .A1(n6376), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6371) );
  INV_X1 U7961 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7962 ( .A1(n6366), .A2(n6365), .ZN(n6377) );
  NAND2_X1 U7963 ( .A1(n6367), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7964 ( .A1(n6377), .A2(n6368), .ZN(n7267) );
  NAND2_X1 U7965 ( .A1(n4297), .A2(n7267), .ZN(n6370) );
  NAND2_X1 U7966 ( .A1(n8318), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6369) );
  NAND4_X1 U7967 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n8530)
         );
  OR2_X1 U7968 ( .A1(n8317), .A2(n6733), .ZN(n6374) );
  OR2_X1 U7969 ( .A1(n8316), .A2(n6732), .ZN(n6373) );
  OAI211_X1 U7970 ( .C1(n6661), .C2(n6734), .A(n6374), .B(n6373), .ZN(n7271)
         );
  INV_X1 U7971 ( .A(n7271), .ZN(n9868) );
  NAND2_X1 U7972 ( .A1(n8530), .A2(n9868), .ZN(n8218) );
  NAND2_X1 U7973 ( .A1(n7254), .A2(n8218), .ZN(n6375) );
  INV_X1 U7974 ( .A(n8530), .ZN(n7331) );
  NAND2_X1 U7975 ( .A1(n7331), .A2(n7271), .ZN(n8221) );
  NAND2_X1 U7976 ( .A1(n6375), .A2(n8221), .ZN(n7294) );
  INV_X1 U7977 ( .A(n6474), .ZN(n6514) );
  NAND2_X1 U7978 ( .A1(n6514), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7979 ( .A1(n6376), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7980 ( .A1(n6377), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7981 ( .A1(n6385), .A2(n6378), .ZN(n7340) );
  NAND2_X1 U7982 ( .A1(n4298), .A2(n7340), .ZN(n6380) );
  NAND2_X1 U7983 ( .A1(n8318), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6379) );
  NAND4_X1 U7984 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n7433)
         );
  INV_X1 U7985 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U7986 ( .A1(n8307), .A2(n6728), .ZN(n6384) );
  NAND2_X1 U7987 ( .A1(n6499), .A2(n9726), .ZN(n6383) );
  OAI211_X1 U7988 ( .C1(n8316), .C2(n6737), .A(n6384), .B(n6383), .ZN(n7341)
         );
  INV_X1 U7989 ( .A(n7341), .ZN(n7304) );
  NOR2_X1 U7990 ( .A1(n7433), .A2(n7304), .ZN(n8203) );
  NAND2_X1 U7991 ( .A1(n7433), .A2(n7304), .ZN(n8226) );
  NAND2_X1 U7992 ( .A1(n6553), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7993 ( .A1(n6376), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6389) );
  INV_X1 U7994 ( .A(n6405), .ZN(n6403) );
  NAND2_X1 U7995 ( .A1(n6385), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7996 ( .A1(n6403), .A2(n6386), .ZN(n7436) );
  NAND2_X1 U7997 ( .A1(n4297), .A2(n7436), .ZN(n6388) );
  NAND2_X1 U7998 ( .A1(n8318), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6387) );
  NAND4_X1 U7999 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n8529)
         );
  INV_X1 U8000 ( .A(n8529), .ZN(n7422) );
  NAND2_X1 U8001 ( .A1(n6747), .A2(n8307), .ZN(n6393) );
  AOI22_X1 U8002 ( .A1(n6500), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6499), .B2(
        n6391), .ZN(n6392) );
  NAND2_X1 U8003 ( .A1(n6393), .A2(n6392), .ZN(n7437) );
  NAND2_X1 U8004 ( .A1(n7422), .A2(n7437), .ZN(n8231) );
  INV_X1 U8005 ( .A(n7437), .ZN(n9874) );
  NAND2_X1 U8006 ( .A1(n8529), .A2(n9874), .ZN(n7418) );
  NAND2_X1 U8007 ( .A1(n6759), .A2(n8307), .ZN(n6395) );
  AOI22_X1 U8008 ( .A1(n6500), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6499), .B2(
        n9757), .ZN(n6394) );
  NAND2_X1 U8009 ( .A1(n6395), .A2(n6394), .ZN(n9883) );
  NAND2_X1 U8010 ( .A1(n6553), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8011 ( .A1(n6376), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6398) );
  XNOR2_X1 U8012 ( .A(n6403), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U8013 ( .A1(n4298), .A2(n7423), .ZN(n6397) );
  NAND2_X1 U8014 ( .A1(n8318), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6396) );
  NAND4_X1 U8015 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n8528)
         );
  OR2_X1 U8016 ( .A1(n9883), .A2(n7760), .ZN(n8224) );
  NAND2_X1 U8017 ( .A1(n9883), .A2(n7760), .ZN(n8232) );
  INV_X1 U8018 ( .A(n7687), .ZN(n6412) );
  NAND2_X1 U8019 ( .A1(n6816), .A2(n8307), .ZN(n6402) );
  AOI22_X1 U8020 ( .A1(n6500), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6499), .B2(
        n6400), .ZN(n6401) );
  NAND2_X1 U8021 ( .A1(n6402), .A2(n6401), .ZN(n9889) );
  NAND2_X1 U8022 ( .A1(n6376), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8023 ( .A1(n8318), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6409) );
  OAI21_X1 U8024 ( .B1(n6403), .B2(P2_REG3_REG_8__SCAN_IN), .A(
        P2_REG3_REG_9__SCAN_IN), .ZN(n6406) );
  NOR2_X1 U8025 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n6404) );
  INV_X1 U8026 ( .A(n6417), .ZN(n6418) );
  NAND2_X1 U8027 ( .A1(n6406), .A2(n6418), .ZN(n7755) );
  NAND2_X1 U8028 ( .A1(n4298), .A2(n7755), .ZN(n6408) );
  NAND2_X1 U8029 ( .A1(n6553), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6407) );
  NAND4_X1 U8030 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n8527)
         );
  NAND2_X1 U8031 ( .A1(n9889), .A2(n7820), .ZN(n8228) );
  NAND2_X1 U8032 ( .A1(n8225), .A2(n8228), .ZN(n8355) );
  OR2_X1 U8033 ( .A1(n6821), .A2(n8317), .ZN(n6415) );
  AOI22_X1 U8034 ( .A1(n6500), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6499), .B2(
        n6413), .ZN(n6414) );
  NAND2_X1 U8035 ( .A1(n6514), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8036 ( .A1(n6376), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6422) );
  INV_X1 U8037 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8038 ( .A1(n6417), .A2(n6416), .ZN(n6427) );
  NAND2_X1 U8039 ( .A1(n6418), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8040 ( .A1(n6427), .A2(n6419), .ZN(n7825) );
  NAND2_X1 U8041 ( .A1(n4298), .A2(n7825), .ZN(n6421) );
  NAND2_X1 U8042 ( .A1(n8318), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6420) );
  NAND4_X1 U8043 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n8526)
         );
  OR2_X1 U8044 ( .A1(n8207), .A2(n7789), .ZN(n8206) );
  NAND2_X1 U8045 ( .A1(n8207), .A2(n7789), .ZN(n8229) );
  NAND2_X1 U8046 ( .A1(n6859), .A2(n8307), .ZN(n6426) );
  AOI22_X1 U8047 ( .A1(n6500), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6499), .B2(
        n6424), .ZN(n6425) );
  NAND2_X1 U8048 ( .A1(n6426), .A2(n6425), .ZN(n8211) );
  NAND2_X1 U8049 ( .A1(n6553), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8050 ( .A1(n6376), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8051 ( .A1(n6427), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8052 ( .A1(n6435), .A2(n6428), .ZN(n7871) );
  NAND2_X1 U8053 ( .A1(n4297), .A2(n7871), .ZN(n6430) );
  NAND2_X1 U8054 ( .A1(n8318), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8055 ( .A1(n8211), .A2(n8209), .ZN(n8236) );
  OR2_X1 U8056 ( .A1(n6919), .A2(n8317), .ZN(n6434) );
  AOI22_X1 U8057 ( .A1(n6500), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6499), .B2(
        n8028), .ZN(n6433) );
  INV_X1 U8058 ( .A(n7958), .ZN(n8245) );
  NAND2_X1 U8059 ( .A1(n6376), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8060 ( .A1(n8318), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8061 ( .A1(n6435), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8062 ( .A1(n6443), .A2(n6436), .ZN(n7909) );
  NAND2_X1 U8063 ( .A1(n4297), .A2(n7909), .ZN(n6438) );
  NAND2_X1 U8064 ( .A1(n6514), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6437) );
  XNOR2_X1 U8065 ( .A(n8245), .B(n8524), .ZN(n8359) );
  NAND2_X1 U8066 ( .A1(n7958), .A2(n8524), .ZN(n8246) );
  NAND2_X1 U8067 ( .A1(n7955), .A2(n8246), .ZN(n7966) );
  OR2_X1 U8068 ( .A1(n8120), .A2(n8317), .ZN(n6442) );
  AOI22_X1 U8069 ( .A1(n6500), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6499), .B2(
        n8118), .ZN(n6441) );
  NAND2_X1 U8070 ( .A1(n6376), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8071 ( .A1(n6514), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6447) );
  INV_X1 U8072 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U8073 ( .A1(n6443), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8074 ( .A1(n6457), .A2(n6444), .ZN(n7975) );
  NAND2_X1 U8075 ( .A1(n4298), .A2(n7975), .ZN(n6446) );
  NAND2_X1 U8076 ( .A1(n8318), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U8077 ( .A1(n8249), .A2(n7995), .ZN(n6449) );
  NAND2_X1 U8078 ( .A1(n7966), .A2(n6449), .ZN(n6451) );
  NAND2_X1 U8079 ( .A1(n7921), .A2(n8523), .ZN(n6450) );
  NAND2_X1 U8080 ( .A1(n6451), .A2(n6450), .ZN(n7999) );
  NAND2_X1 U8081 ( .A1(n7096), .A2(n8307), .ZN(n6454) );
  AOI22_X1 U8082 ( .A1(n6500), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6499), .B2(
        n6452), .ZN(n6453) );
  NAND2_X1 U8083 ( .A1(n6376), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8084 ( .A1(n8318), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6461) );
  INV_X1 U8085 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U8086 ( .A1(n6456), .A2(n6455), .ZN(n6465) );
  NAND2_X1 U8087 ( .A1(n6457), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8088 ( .A1(n6465), .A2(n6458), .ZN(n8043) );
  NAND2_X1 U8089 ( .A1(n4298), .A2(n8043), .ZN(n6460) );
  NAND2_X1 U8090 ( .A1(n6553), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6459) );
  NAND4_X1 U8091 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .ZN(n8522)
         );
  INV_X1 U8092 ( .A(n8522), .ZN(n8005) );
  NOR2_X1 U8093 ( .A1(n8038), .A2(n8005), .ZN(n8255) );
  NAND2_X1 U8094 ( .A1(n8038), .A2(n8005), .ZN(n7994) );
  NAND2_X1 U8095 ( .A1(n7100), .A2(n8307), .ZN(n6464) );
  AOI22_X1 U8096 ( .A1(n6500), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6499), .B2(
        n8538), .ZN(n6463) );
  NAND2_X1 U8097 ( .A1(n6553), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8098 ( .A1(n6376), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U8099 ( .A1(n6465), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8100 ( .A1(n6475), .A2(n6466), .ZN(n8098) );
  NAND2_X1 U8101 ( .A1(n4298), .A2(n8098), .ZN(n6468) );
  NAND2_X1 U8102 ( .A1(n8318), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8103 ( .A1(n8099), .A2(n8748), .ZN(n8264) );
  NAND2_X1 U8104 ( .A1(n7151), .A2(n8307), .ZN(n6473) );
  AOI22_X1 U8105 ( .A1(n6500), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6499), .B2(
        n6471), .ZN(n6472) );
  NAND2_X1 U8106 ( .A1(n6514), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8107 ( .A1(n6376), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6479) );
  INV_X1 U8108 ( .A(n6493), .ZN(n6491) );
  NAND2_X1 U8109 ( .A1(n6475), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8110 ( .A1(n6491), .A2(n6476), .ZN(n8754) );
  NAND2_X1 U8111 ( .A1(n4298), .A2(n8754), .ZN(n6478) );
  NAND2_X1 U8112 ( .A1(n8318), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8113 ( .A1(n8888), .A2(n8457), .ZN(n8265) );
  NAND2_X1 U8114 ( .A1(n6481), .A2(n8267), .ZN(n8730) );
  NAND2_X1 U8115 ( .A1(n7287), .A2(n8307), .ZN(n6483) );
  AOI22_X1 U8116 ( .A1(n6500), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6499), .B2(
        n9810), .ZN(n6482) );
  NAND2_X1 U8117 ( .A1(n6553), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8118 ( .A1(n6376), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6486) );
  XNOR2_X1 U8119 ( .A(n6491), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U8120 ( .A1(n4297), .A2(n8738), .ZN(n6485) );
  NAND2_X1 U8121 ( .A1(n8318), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6484) );
  INV_X1 U8122 ( .A(n8178), .ZN(n6488) );
  NAND2_X1 U8123 ( .A1(n8881), .A2(n8746), .ZN(n8176) );
  NAND2_X1 U8124 ( .A1(n7299), .A2(n8307), .ZN(n6490) );
  AOI22_X1 U8125 ( .A1(n6500), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6499), .B2(
        n8567), .ZN(n6489) );
  NAND2_X1 U8126 ( .A1(n6514), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8127 ( .A1(n6376), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6497) );
  OAI21_X1 U8128 ( .B1(n6491), .B2(P2_REG3_REG_17__SCAN_IN), .A(
        P2_REG3_REG_18__SCAN_IN), .ZN(n6494) );
  NOR2_X1 U8129 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6492) );
  INV_X1 U8130 ( .A(n6504), .ZN(n6505) );
  NAND2_X1 U8131 ( .A1(n6494), .A2(n6505), .ZN(n8726) );
  NAND2_X1 U8132 ( .A1(n4297), .A2(n8726), .ZN(n6496) );
  NAND2_X1 U8133 ( .A1(n8318), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6495) );
  NAND4_X1 U8134 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n8734)
         );
  INV_X1 U8135 ( .A(n8734), .ZN(n8413) );
  NAND2_X1 U8136 ( .A1(n8875), .A2(n8413), .ZN(n8177) );
  NAND2_X1 U8137 ( .A1(n8709), .A2(n8177), .ZN(n8339) );
  NAND2_X1 U8138 ( .A1(n7557), .A2(n8307), .ZN(n6502) );
  AOI22_X1 U8139 ( .A1(n6500), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8382), .B2(
        n6499), .ZN(n6501) );
  NAND2_X1 U8140 ( .A1(n6376), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8141 ( .A1(n6514), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6509) );
  INV_X1 U8142 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8143 ( .A1(n6505), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8144 ( .A1(n6515), .A2(n6506), .ZN(n8716) );
  NAND2_X1 U8145 ( .A1(n4298), .A2(n8716), .ZN(n6508) );
  NAND2_X1 U8146 ( .A1(n8318), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6507) );
  OR2_X1 U8147 ( .A1(n8869), .A2(n8479), .ZN(n8173) );
  AND2_X1 U8148 ( .A1(n8173), .A2(n8709), .ZN(n8175) );
  NAND2_X1 U8149 ( .A1(n8869), .A2(n8479), .ZN(n8273) );
  NAND2_X1 U8150 ( .A1(n7681), .A2(n8307), .ZN(n6513) );
  INV_X1 U8151 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6511) );
  OR2_X1 U8152 ( .A1(n8316), .A2(n6511), .ZN(n6512) );
  NAND2_X1 U8153 ( .A1(n6514), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8154 ( .A1(n6376), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U8155 ( .A1(n6515), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8156 ( .A1(n6525), .A2(n6516), .ZN(n8706) );
  NAND2_X1 U8157 ( .A1(n4298), .A2(n8706), .ZN(n6518) );
  NAND2_X1 U8158 ( .A1(n8318), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8159 ( .A1(n8701), .A2(n8277), .ZN(n8685) );
  NAND2_X1 U8160 ( .A1(n7720), .A2(n8307), .ZN(n6522) );
  OR2_X1 U8161 ( .A1(n8316), .A2(n10021), .ZN(n6521) );
  NAND2_X1 U8162 ( .A1(n6376), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8163 ( .A1(n6553), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6523) );
  AND2_X1 U8164 ( .A1(n6524), .A2(n6523), .ZN(n6529) );
  INV_X1 U8165 ( .A(n6534), .ZN(n6535) );
  NAND2_X1 U8166 ( .A1(n6525), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8167 ( .A1(n6535), .A2(n6526), .ZN(n8695) );
  NAND2_X1 U8168 ( .A1(n8695), .A2(n4297), .ZN(n6528) );
  NAND2_X1 U8169 ( .A1(n8318), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8170 ( .A1(n8864), .A2(n8693), .ZN(n8684) );
  NAND2_X1 U8171 ( .A1(n8685), .A2(n4387), .ZN(n6530) );
  NAND2_X1 U8172 ( .A1(n7877), .A2(n8307), .ZN(n6532) );
  OR2_X1 U8173 ( .A1(n8316), .A2(n7878), .ZN(n6531) );
  INV_X1 U8174 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8788) );
  INV_X1 U8175 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6533) );
  INV_X1 U8176 ( .A(n6543), .ZN(n6544) );
  NAND2_X1 U8177 ( .A1(n6535), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8178 ( .A1(n6544), .A2(n6536), .ZN(n8681) );
  NAND2_X1 U8179 ( .A1(n8681), .A2(n4298), .ZN(n6538) );
  AOI22_X1 U8180 ( .A1(n6514), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6376), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6537) );
  OAI211_X1 U8181 ( .C1(n6655), .C2(n8788), .A(n6538), .B(n6537), .ZN(n8665)
         );
  INV_X1 U8182 ( .A(n8665), .ZN(n8694) );
  NAND2_X1 U8183 ( .A1(n8854), .A2(n8694), .ZN(n6539) );
  NAND2_X1 U8184 ( .A1(n7900), .A2(n8307), .ZN(n6541) );
  OR2_X1 U8185 ( .A1(n8316), .A2(n7902), .ZN(n6540) );
  INV_X1 U8186 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8785) );
  INV_X1 U8187 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8188 ( .A1(n6544), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8189 ( .A1(n6551), .A2(n6545), .ZN(n8669) );
  NAND2_X1 U8190 ( .A1(n8669), .A2(n4297), .ZN(n6547) );
  AOI22_X1 U8191 ( .A1(n6553), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n6376), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6546) );
  OAI211_X1 U8192 ( .C1(n6655), .C2(n8785), .A(n6547), .B(n6546), .ZN(n8678)
         );
  INV_X1 U8193 ( .A(n8678), .ZN(n8487) );
  NAND2_X1 U8194 ( .A1(n8662), .A2(n8338), .ZN(n6548) );
  NAND2_X1 U8195 ( .A1(n8848), .A2(n8487), .ZN(n8337) );
  NAND2_X1 U8196 ( .A1(n6548), .A2(n8337), .ZN(n8654) );
  NAND2_X1 U8197 ( .A1(n7979), .A2(n8307), .ZN(n6550) );
  OR2_X1 U8198 ( .A1(n8316), .A2(n9961), .ZN(n6549) );
  NAND2_X1 U8199 ( .A1(n6551), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8200 ( .A1(n6561), .A2(n6552), .ZN(n8659) );
  NAND2_X1 U8201 ( .A1(n8659), .A2(n4298), .ZN(n6558) );
  INV_X1 U8202 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U8203 ( .A1(n6553), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U8204 ( .A1(n4295), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6554) );
  OAI211_X1 U8205 ( .C1(n8782), .C2(n6655), .A(n6555), .B(n6554), .ZN(n6556)
         );
  INV_X1 U8206 ( .A(n6556), .ZN(n6557) );
  AND2_X1 U8207 ( .A1(n8843), .A2(n8436), .ZN(n8289) );
  NAND2_X1 U8208 ( .A1(n7990), .A2(n8307), .ZN(n6560) );
  OR2_X1 U8209 ( .A1(n8316), .A2(n8115), .ZN(n6559) );
  NAND2_X1 U8210 ( .A1(n6561), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8211 ( .A1(n6571), .A2(n6562), .ZN(n8651) );
  NAND2_X1 U8212 ( .A1(n8651), .A2(n4298), .ZN(n6567) );
  INV_X1 U8213 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U8214 ( .A1(n6553), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U8215 ( .A1(n8318), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6563) );
  OAI211_X1 U8216 ( .C1(n4296), .C2(n10005), .A(n6564), .B(n6563), .ZN(n6565)
         );
  INV_X1 U8217 ( .A(n6565), .ZN(n6566) );
  NAND2_X1 U8218 ( .A1(n8837), .A2(n8468), .ZN(n8297) );
  INV_X1 U8219 ( .A(n8296), .ZN(n6568) );
  NAND2_X1 U8220 ( .A1(n8084), .A2(n8307), .ZN(n6570) );
  OR2_X1 U8221 ( .A1(n8316), .A2(n8085), .ZN(n6569) );
  INV_X1 U8222 ( .A(n6582), .ZN(n6583) );
  NAND2_X1 U8223 ( .A1(n6571), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U8224 ( .A1(n6583), .A2(n6572), .ZN(n8635) );
  NAND2_X1 U8225 ( .A1(n8635), .A2(n4297), .ZN(n6577) );
  INV_X1 U8226 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U8227 ( .A1(n6553), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8228 ( .A1(n6376), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U8229 ( .C1(n8776), .C2(n6655), .A(n6574), .B(n6573), .ZN(n6575)
         );
  INV_X1 U8230 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U8231 ( .A1(n8103), .A2(n8307), .ZN(n6580) );
  OR2_X1 U8232 ( .A1(n8316), .A2(n6578), .ZN(n6579) );
  INV_X1 U8233 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U8234 ( .A1(n6582), .A2(n6581), .ZN(n6593) );
  NAND2_X1 U8235 ( .A1(n6583), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8236 ( .A1(n6593), .A2(n6584), .ZN(n8624) );
  NAND2_X1 U8237 ( .A1(n8624), .A2(n4297), .ZN(n6589) );
  INV_X1 U8238 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U8239 ( .A1(n4295), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U8240 ( .A1(n6514), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6585) );
  OAI211_X1 U8241 ( .C1(n6655), .C2(n8773), .A(n6586), .B(n6585), .ZN(n6587)
         );
  INV_X1 U8242 ( .A(n6587), .ZN(n6588) );
  AND2_X1 U8243 ( .A1(n8608), .A2(n8302), .ZN(n8588) );
  NAND2_X1 U8244 ( .A1(n8113), .A2(n8307), .ZN(n6592) );
  OR2_X1 U8245 ( .A1(n8316), .A2(n6590), .ZN(n6591) );
  NAND2_X1 U8246 ( .A1(n6593), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8247 ( .A1(n8573), .A2(n6594), .ZN(n8604) );
  NAND2_X1 U8248 ( .A1(n8604), .A2(n4298), .ZN(n6599) );
  INV_X1 U8249 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U8250 ( .A1(n6553), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8251 ( .A1(n6376), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6595) );
  OAI211_X1 U8252 ( .C1(n9962), .C2(n6655), .A(n6596), .B(n6595), .ZN(n6597)
         );
  INV_X1 U8253 ( .A(n6597), .ZN(n6598) );
  OR2_X1 U8254 ( .A1(n8770), .A2(n8619), .ZN(n6600) );
  INV_X1 U8255 ( .A(n6600), .ZN(n6602) );
  INV_X1 U8256 ( .A(n8302), .ZN(n6601) );
  NAND2_X1 U8257 ( .A1(n8832), .A2(n8618), .ZN(n8609) );
  NAND2_X1 U8258 ( .A1(n8826), .A2(n8599), .ZN(n8303) );
  AND2_X1 U8259 ( .A1(n8609), .A2(n8616), .ZN(n8610) );
  XNOR2_X1 U8260 ( .A(n8770), .B(n8619), .ZN(n8597) );
  INV_X1 U8261 ( .A(n8597), .ZN(n8590) );
  AND2_X1 U8262 ( .A1(n8589), .A2(n8590), .ZN(n8592) );
  INV_X1 U8263 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8111) );
  OR2_X1 U8264 ( .A1(n8316), .A2(n8111), .ZN(n6603) );
  NAND2_X1 U8265 ( .A1(n8579), .A2(n4297), .ZN(n8323) );
  INV_X1 U8266 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8267 ( .A1(n6376), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8268 ( .A1(n6514), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6605) );
  OAI211_X1 U8269 ( .C1(n6655), .C2(n6703), .A(n6606), .B(n6605), .ZN(n6607)
         );
  INV_X1 U8270 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8271 ( .A1(n6691), .A2(n8600), .ZN(n8330) );
  INV_X1 U8272 ( .A(n6609), .ZN(n6610) );
  NAND2_X1 U8273 ( .A1(n6610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U8274 ( .A1(n7559), .A2(n7682), .ZN(n6988) );
  NAND2_X1 U8275 ( .A1(n8342), .A2(n7682), .ZN(n7156) );
  NAND2_X1 U8276 ( .A1(n7879), .A2(n7156), .ZN(n6613) );
  NAND2_X1 U8277 ( .A1(n6613), .A2(n7559), .ZN(n6693) );
  INV_X1 U8278 ( .A(n6693), .ZN(n6614) );
  NAND2_X1 U8279 ( .A1(n8532), .A2(n6939), .ZN(n7137) );
  INV_X1 U8280 ( .A(n4293), .ZN(n7030) );
  NAND2_X1 U8281 ( .A1(n7030), .A2(n6992), .ZN(n9837) );
  NAND2_X1 U8282 ( .A1(n7136), .A2(n9837), .ZN(n6616) );
  NAND2_X1 U8283 ( .A1(n6616), .A2(n8344), .ZN(n7213) );
  NAND2_X1 U8284 ( .A1(n7033), .A2(n9854), .ZN(n7214) );
  NAND2_X1 U8285 ( .A1(n7213), .A2(n7214), .ZN(n7201) );
  AND2_X1 U8286 ( .A1(n8197), .A2(n8343), .ZN(n6617) );
  NAND2_X1 U8287 ( .A1(n7201), .A2(n6617), .ZN(n7200) );
  NAND2_X1 U8288 ( .A1(n7147), .A2(n9863), .ZN(n7257) );
  AND2_X1 U8289 ( .A1(n4909), .A2(n7257), .ZN(n6619) );
  INV_X1 U8290 ( .A(n8197), .ZN(n6618) );
  INV_X1 U8291 ( .A(n9842), .ZN(n7036) );
  NAND2_X1 U8292 ( .A1(n7036), .A2(n7224), .ZN(n7202) );
  OR2_X1 U8293 ( .A1(n6618), .A2(n7202), .ZN(n7258) );
  NAND2_X1 U8294 ( .A1(n8530), .A2(n7271), .ZN(n7256) );
  AND2_X1 U8295 ( .A1(n7433), .A2(n7341), .ZN(n6620) );
  NAND2_X1 U8296 ( .A1(n8529), .A2(n7437), .ZN(n6621) );
  NAND2_X1 U8297 ( .A1(n8207), .A2(n8526), .ZN(n6622) );
  NAND2_X1 U8298 ( .A1(n7771), .A2(n8357), .ZN(n7770) );
  INV_X1 U8299 ( .A(n8209), .ZN(n8525) );
  NAND2_X1 U8300 ( .A1(n8211), .A2(n8525), .ZN(n6623) );
  NAND2_X1 U8301 ( .A1(n7770), .A2(n6623), .ZN(n7903) );
  NAND2_X1 U8302 ( .A1(n7958), .A2(n8244), .ZN(n6624) );
  NAND2_X1 U8303 ( .A1(n8245), .A2(n8524), .ZN(n6625) );
  NAND2_X1 U8304 ( .A1(n7921), .A2(n7995), .ZN(n8252) );
  NAND2_X1 U8305 ( .A1(n8249), .A2(n8523), .ZN(n8250) );
  NAND2_X1 U8306 ( .A1(n8252), .A2(n8250), .ZN(n8358) );
  NAND2_X1 U8307 ( .A1(n7967), .A2(n8252), .ZN(n7993) );
  NAND2_X1 U8308 ( .A1(n8038), .A2(n8522), .ZN(n6627) );
  NAND2_X1 U8309 ( .A1(n7993), .A2(n6627), .ZN(n6629) );
  OR2_X1 U8310 ( .A1(n8038), .A2(n8522), .ZN(n6628) );
  NAND2_X1 U8311 ( .A1(n6629), .A2(n6628), .ZN(n8090) );
  NAND2_X1 U8312 ( .A1(n8261), .A2(n8264), .ZN(n8362) );
  NAND2_X1 U8313 ( .A1(n8090), .A2(n8362), .ZN(n6631) );
  OR2_X1 U8314 ( .A1(n8099), .A2(n8521), .ZN(n6630) );
  INV_X1 U8315 ( .A(n8457), .ZN(n8735) );
  NAND2_X1 U8316 ( .A1(n8888), .A2(n8735), .ZN(n6633) );
  NAND2_X1 U8317 ( .A1(n8178), .A2(n8176), .ZN(n8732) );
  NAND2_X1 U8318 ( .A1(n8733), .A2(n8732), .ZN(n8731) );
  NAND2_X1 U8319 ( .A1(n8881), .A2(n8722), .ZN(n6634) );
  NAND2_X1 U8320 ( .A1(n8731), .A2(n6634), .ZN(n8720) );
  OR2_X1 U8321 ( .A1(n8875), .A2(n8734), .ZN(n6635) );
  NAND2_X1 U8322 ( .A1(n8720), .A2(n6635), .ZN(n6637) );
  NAND2_X1 U8323 ( .A1(n8875), .A2(n8734), .ZN(n6636) );
  NAND2_X1 U8324 ( .A1(n6637), .A2(n6636), .ZN(n8711) );
  NAND2_X1 U8325 ( .A1(n8173), .A2(n8273), .ZN(n8340) );
  NAND2_X1 U8326 ( .A1(n8869), .A2(n8723), .ZN(n6638) );
  INV_X1 U8327 ( .A(n8702), .ZN(n6639) );
  INV_X1 U8328 ( .A(n8693), .ZN(n8713) );
  OR2_X1 U8329 ( .A1(n8864), .A2(n8713), .ZN(n8689) );
  NAND2_X1 U8330 ( .A1(n8687), .A2(n8689), .ZN(n6640) );
  NAND2_X1 U8331 ( .A1(n8279), .A2(n8278), .ZN(n8688) );
  OR2_X1 U8332 ( .A1(n8792), .A2(n8703), .ZN(n8675) );
  OR2_X1 U8333 ( .A1(n8854), .A2(n8665), .ZN(n8282) );
  NAND2_X1 U8334 ( .A1(n8854), .A2(n8665), .ZN(n8287) );
  NAND2_X1 U8335 ( .A1(n8848), .A2(n8678), .ZN(n6641) );
  NAND2_X1 U8336 ( .A1(n8663), .A2(n6641), .ZN(n6643) );
  OR2_X1 U8337 ( .A1(n8848), .A2(n8678), .ZN(n6642) );
  NOR2_X1 U8338 ( .A1(n8843), .A2(n8666), .ZN(n8641) );
  NAND2_X1 U8339 ( .A1(n8843), .A2(n8666), .ZN(n8642) );
  INV_X1 U8340 ( .A(n8638), .ZN(n8646) );
  AND2_X1 U8341 ( .A1(n8642), .A2(n8646), .ZN(n8643) );
  NAND2_X1 U8342 ( .A1(n8832), .A2(n8648), .ZN(n6644) );
  AND2_X1 U8343 ( .A1(n8629), .A2(n6644), .ZN(n6645) );
  INV_X1 U8344 ( .A(n8616), .ZN(n8367) );
  OR2_X1 U8345 ( .A1(n8832), .A2(n8648), .ZN(n8614) );
  AND2_X1 U8346 ( .A1(n8367), .A2(n8614), .ZN(n6646) );
  NAND2_X1 U8347 ( .A1(n8615), .A2(n6646), .ZN(n8621) );
  NAND2_X1 U8348 ( .A1(n8826), .A2(n8632), .ZN(n6647) );
  NAND2_X1 U8349 ( .A1(n8621), .A2(n6647), .ZN(n8598) );
  NAND2_X1 U8350 ( .A1(n8598), .A2(n8597), .ZN(n8596) );
  INV_X1 U8351 ( .A(n8770), .ZN(n8823) );
  NAND2_X1 U8352 ( .A1(n8596), .A2(n6649), .ZN(n6650) );
  XNOR2_X1 U8353 ( .A(n6650), .B(n4676), .ZN(n6652) );
  OR2_X1 U8354 ( .A1(n7879), .A2(n7559), .ZN(n6682) );
  INV_X1 U8355 ( .A(n7682), .ZN(n8375) );
  NAND2_X1 U8356 ( .A1(n8342), .A2(n8375), .ZN(n6651) );
  NAND2_X1 U8357 ( .A1(n6652), .A2(n9844), .ZN(n6664) );
  INV_X1 U8358 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8359 ( .A1(n6514), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8360 ( .A1(n6376), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6653) );
  OAI211_X1 U8361 ( .C1(n6656), .C2(n6655), .A(n6654), .B(n6653), .ZN(n6657)
         );
  INV_X1 U8362 ( .A(n6657), .ZN(n6658) );
  NAND2_X1 U8363 ( .A1(n8323), .A2(n6658), .ZN(n8520) );
  NAND2_X1 U8364 ( .A1(n6659), .A2(n8385), .ZN(n6660) );
  NAND2_X1 U8365 ( .A1(n6661), .A2(n6660), .ZN(n6993) );
  AND2_X1 U8366 ( .A1(n6661), .A2(P2_B_REG_SCAN_IN), .ZN(n6662) );
  NOR2_X1 U8367 ( .A1(n8745), .A2(n6662), .ZN(n8570) );
  INV_X1 U8368 ( .A(n6993), .ZN(n6927) );
  AOI22_X1 U8369 ( .A1(n8520), .A2(n8570), .B1(n6648), .B2(n9840), .ZN(n6663)
         );
  NAND2_X1 U8370 ( .A1(n8382), .A2(n7682), .ZN(n6687) );
  NOR2_X1 U8371 ( .A1(n8577), .A2(n6665), .ZN(n6702) );
  XNOR2_X1 U8372 ( .A(n8172), .B(P2_B_REG_SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8373 ( .A1(n8117), .A2(n6666), .ZN(n6668) );
  NAND2_X1 U8374 ( .A1(n8117), .A2(n8086), .ZN(n6754) );
  NAND2_X1 U8375 ( .A1(n8086), .A2(n8172), .ZN(n6757) );
  NAND2_X1 U8376 ( .A1(n7045), .A2(n7046), .ZN(n6700) );
  NOR2_X1 U8377 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .ZN(
        n6673) );
  NOR4_X1 U8378 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6672) );
  NOR4_X1 U8379 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6671) );
  NOR4_X1 U8380 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6670) );
  NAND4_X1 U8381 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n6679)
         );
  NOR4_X1 U8382 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6677) );
  NOR4_X1 U8383 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6676) );
  NOR4_X1 U8384 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6675) );
  NOR4_X1 U8385 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6674) );
  NAND4_X1 U8386 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6678)
         );
  NOR2_X1 U8387 ( .A1(n6679), .A2(n6678), .ZN(n6680) );
  INV_X1 U8388 ( .A(n6699), .ZN(n6681) );
  INV_X1 U8389 ( .A(n6682), .ZN(n6683) );
  NOR2_X1 U8390 ( .A1(n8342), .A2(n7682), .ZN(n6985) );
  NAND2_X1 U8391 ( .A1(n6683), .A2(n6985), .ZN(n6944) );
  NAND2_X1 U8392 ( .A1(n6944), .A2(n7042), .ZN(n6684) );
  NAND2_X1 U8393 ( .A1(n6935), .A2(n6684), .ZN(n6689) );
  NAND2_X1 U8394 ( .A1(n6987), .A2(n6699), .ZN(n6685) );
  INV_X1 U8395 ( .A(n6946), .ZN(n6686) );
  INV_X1 U8396 ( .A(n8342), .ZN(n8328) );
  NAND3_X1 U8397 ( .A1(n6944), .A2(n8310), .A3(n9873), .ZN(n6928) );
  NAND2_X1 U8398 ( .A1(n9890), .A2(n6687), .ZN(n9836) );
  NAND2_X1 U8399 ( .A1(n6928), .A2(n9836), .ZN(n6940) );
  NAND2_X1 U8400 ( .A1(n6931), .A2(n6940), .ZN(n6688) );
  MUX2_X1 U8401 ( .A(n6690), .B(n6702), .S(n9891), .Z(n6692) );
  INV_X1 U8402 ( .A(n6691), .ZN(n8582) );
  NAND2_X1 U8403 ( .A1(n6692), .A2(n4900), .ZN(P2_U3456) );
  OR2_X1 U8404 ( .A1(n6693), .A2(n7682), .ZN(n6694) );
  NAND2_X1 U8405 ( .A1(n6694), .A2(n8310), .ZN(n6696) );
  NAND2_X1 U8406 ( .A1(n7045), .A2(n6696), .ZN(n6695) );
  OAI21_X1 U8407 ( .B1(n6696), .B2(n6987), .A(n6695), .ZN(n7048) );
  NAND2_X1 U8408 ( .A1(n8326), .A2(n6988), .ZN(n6697) );
  AND2_X1 U8409 ( .A1(n6698), .A2(n6697), .ZN(n6943) );
  NAND3_X1 U8410 ( .A1(n6699), .A2(n6950), .A3(n6943), .ZN(n7043) );
  NOR2_X1 U8411 ( .A1(n9885), .A2(n8342), .ZN(n6936) );
  NOR2_X1 U8412 ( .A1(n7043), .A2(n6936), .ZN(n6701) );
  MUX2_X1 U8413 ( .A(n6703), .B(n6702), .S(n9904), .Z(n6704) );
  NAND2_X1 U8414 ( .A1(n9904), .A2(n9890), .ZN(n7307) );
  NAND2_X1 U8415 ( .A1(n6704), .A2(n4903), .ZN(P2_U3488) );
  NAND2_X1 U8416 ( .A1(n9022), .A2(n8983), .ZN(n6708) );
  NAND2_X1 U8417 ( .A1(n9024), .A2(n8982), .ZN(n6707) );
  NAND2_X1 U8418 ( .A1(n6708), .A2(n6707), .ZN(n9174) );
  OAI22_X1 U8419 ( .A1(n9179), .A2(n8998), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6709), .ZN(n6710) );
  AOI21_X1 U8420 ( .B1(n9174), .B2(n9001), .A(n6710), .ZN(n6711) );
  INV_X1 U8421 ( .A(n6712), .ZN(n6713) );
  NOR2_X1 U8422 ( .A1(n6714), .A2(P1_U3086), .ZN(n6716) );
  NAND2_X1 U8423 ( .A1(n6722), .A2(P1_U3086), .ZN(n8108) );
  NAND2_X2 U8424 ( .A1(n6717), .A2(P1_U3086), .ZN(n9452) );
  OAI222_X1 U8425 ( .A1(n8108), .A2(n4935), .B1(n9452), .B2(n4327), .C1(
        P1_U3086), .C2(n6778), .ZN(P1_U3354) );
  OAI222_X1 U8426 ( .A1(n8108), .A2(n6718), .B1(n9452), .B2(n6731), .C1(
        P1_U3086), .C2(n6800), .ZN(P1_U3352) );
  OAI222_X1 U8427 ( .A1(n8108), .A2(n6719), .B1(n9452), .B2(n6736), .C1(
        P1_U3086), .C2(n6872), .ZN(P1_U3351) );
  INV_X1 U8428 ( .A(n8108), .ZN(n9447) );
  AOI22_X1 U8429 ( .A1(n6813), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9447), .ZN(n6720) );
  OAI21_X1 U8430 ( .B1(n6733), .B2(n9452), .A(n6720), .ZN(P1_U3350) );
  OAI222_X1 U8431 ( .A1(n9450), .A2(n6721), .B1(n9452), .B2(n6726), .C1(
        P1_U3086), .C2(n9497), .ZN(P1_U3353) );
  NAND2_X1 U8432 ( .A1(n6722), .A2(P2_U3151), .ZN(n8901) );
  INV_X1 U8433 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6723) );
  NOR2_X1 U8434 ( .A1(n6722), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8904) );
  INV_X2 U8435 ( .A(n8904), .ZN(n8899) );
  OAI222_X1 U8436 ( .A1(P2_U3151), .A2(n6724), .B1(n8901), .B2(n4327), .C1(
        n6723), .C2(n8899), .ZN(P2_U3294) );
  OAI222_X1 U8437 ( .A1(n6727), .A2(P2_U3151), .B1(n8901), .B2(n6726), .C1(
        n6725), .C2(n8899), .ZN(P2_U3293) );
  INV_X1 U8438 ( .A(n6824), .ZN(n6830) );
  INV_X1 U8439 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6858) );
  INV_X1 U8440 ( .A(n6728), .ZN(n6738) );
  OAI222_X1 U8441 ( .A1(P1_U3086), .A2(n6830), .B1(n9450), .B2(n6858), .C1(
        n6738), .C2(n9452), .ZN(P1_U3349) );
  INV_X1 U8442 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U8443 ( .A1(n6753), .A2(n10027), .ZN(P2_U3253) );
  INV_X1 U8444 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10023) );
  NOR2_X1 U8445 ( .A1(n6753), .A2(n10023), .ZN(P2_U3237) );
  INV_X1 U8446 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U8447 ( .A1(n6753), .A2(n10018), .ZN(P2_U3256) );
  INV_X1 U8448 ( .A(n8901), .ZN(n7899) );
  OAI222_X1 U8449 ( .A1(n6896), .A2(P2_U3151), .B1(n8906), .B2(n6731), .C1(
        n6730), .C2(n8899), .ZN(P2_U3292) );
  OAI222_X1 U8450 ( .A1(n6734), .A2(P2_U3151), .B1(n8906), .B2(n6733), .C1(
        n6732), .C2(n8899), .ZN(P2_U3290) );
  OAI222_X1 U8451 ( .A1(n7026), .A2(P2_U3151), .B1(n8906), .B2(n6736), .C1(
        n6735), .C2(n8899), .ZN(P2_U3291) );
  OAI222_X1 U8452 ( .A1(P2_U3151), .A2(n6739), .B1(n8906), .B2(n6738), .C1(
        n6737), .C2(n8899), .ZN(P2_U3289) );
  NAND2_X1 U8453 ( .A1(n6740), .A2(n7896), .ZN(n6770) );
  INV_X1 U8454 ( .A(n6770), .ZN(n6745) );
  OR2_X1 U8455 ( .A1(n6742), .A2(n6741), .ZN(n6744) );
  NOR2_X2 U8456 ( .A1(n6745), .A2(n6769), .ZN(n9490) );
  NOR2_X1 U8457 ( .A1(n9490), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8458 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U8459 ( .A1(n6192), .A2(P1_U3973), .ZN(n6746) );
  OAI21_X1 U8460 ( .B1(P1_U3973), .B2(n9956), .A(n6746), .ZN(P1_U3554) );
  INV_X1 U8461 ( .A(n6747), .ZN(n6749) );
  INV_X1 U8462 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6748) );
  OAI222_X1 U8463 ( .A1(P2_U3151), .A2(n7195), .B1(n8906), .B2(n6749), .C1(
        n6748), .C2(n8899), .ZN(P2_U3288) );
  INV_X1 U8464 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6750) );
  INV_X1 U8465 ( .A(n6906), .ZN(n6836) );
  OAI222_X1 U8466 ( .A1(n8108), .A2(n6750), .B1(n9452), .B2(n6749), .C1(n6836), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  AND2_X1 U8467 ( .A1(n6751), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8468 ( .A1(n6751), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8469 ( .A1(n6751), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8470 ( .A1(n6751), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8471 ( .A1(n6751), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8472 ( .A1(n6751), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8473 ( .A1(n6751), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8474 ( .A1(n6751), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8475 ( .A1(n6751), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8476 ( .A1(n6751), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8477 ( .A1(n6751), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8478 ( .A1(n6751), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8479 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8480 ( .A1(n7545), .A2(P1_U3973), .ZN(n6752) );
  OAI21_X1 U8481 ( .B1(n6917), .B2(P1_U3973), .A(n6752), .ZN(P1_U3566) );
  INV_X1 U8482 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6756) );
  INV_X1 U8483 ( .A(n6754), .ZN(n6755) );
  AOI22_X1 U8484 ( .A1(n6751), .A2(n6756), .B1(n6950), .B2(n6755), .ZN(
        P2_U3377) );
  INV_X1 U8485 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9986) );
  INV_X1 U8486 ( .A(n6757), .ZN(n6758) );
  AOI22_X1 U8487 ( .A1(n6751), .A2(n9986), .B1(n6950), .B2(n6758), .ZN(
        P2_U3376) );
  INV_X1 U8488 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6760) );
  INV_X1 U8489 ( .A(n6759), .ZN(n6762) );
  INV_X1 U8490 ( .A(n6973), .ZN(n6914) );
  OAI222_X1 U8491 ( .A1(n8108), .A2(n6760), .B1(n9452), .B2(n6762), .C1(
        P1_U3086), .C2(n6914), .ZN(P1_U3347) );
  INV_X1 U8492 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6761) );
  OAI222_X1 U8493 ( .A1(n6763), .A2(P2_U3151), .B1(n8906), .B2(n6762), .C1(
        n6761), .C2(n8899), .ZN(P2_U3287) );
  INV_X1 U8494 ( .A(n6872), .ZN(n6766) );
  NAND2_X1 U8495 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9475) );
  NOR2_X1 U8496 ( .A1(n9474), .A2(n9475), .ZN(n9473) );
  AOI21_X1 U8497 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9477), .A(n9473), .ZN(
        n9489) );
  INV_X1 U8498 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9999) );
  AOI22_X1 U8499 ( .A1(n6777), .A2(n9999), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n9497), .ZN(n9488) );
  NOR2_X1 U8500 ( .A1(n9489), .A2(n9488), .ZN(n9487) );
  INV_X1 U8501 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U8502 ( .A1(n6776), .A2(n6764), .B1(P1_REG2_REG_3__SCAN_IN), .B2(
        n6800), .ZN(n6792) );
  INV_X1 U8503 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6765) );
  MUX2_X1 U8504 ( .A(n6765), .B(P1_REG2_REG_4__SCAN_IN), .S(n6872), .Z(n6877)
         );
  NAND2_X1 U8505 ( .A1(n6876), .A2(n6877), .ZN(n6875) );
  NAND2_X1 U8506 ( .A1(n6813), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U8507 ( .B1(n6813), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6767), .ZN(
        n6809) );
  INV_X1 U8508 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6768) );
  AOI22_X1 U8509 ( .A1(n6824), .A2(n6768), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n6830), .ZN(n6773) );
  NOR2_X1 U8510 ( .A1(n6774), .A2(n6773), .ZN(n6823) );
  NAND2_X1 U8511 ( .A1(n6770), .A2(n6769), .ZN(n9472) );
  INV_X1 U8512 ( .A(n9472), .ZN(n6772) );
  NOR2_X1 U8513 ( .A1(n5605), .A2(n4294), .ZN(n6771) );
  AOI211_X1 U8514 ( .C1(n6774), .C2(n6773), .A(n6823), .B(n9486), .ZN(n6790)
         );
  AND2_X1 U8515 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6775) );
  AOI21_X1 U8516 ( .B1(n9490), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6775), .ZN(
        n6788) );
  NAND2_X1 U8517 ( .A1(n6813), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6783) );
  INV_X1 U8518 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U8519 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9657), .S(n6872), .Z(n6874)
         );
  INV_X1 U8520 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U8521 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9655), .S(n6776), .Z(n6796)
         );
  INV_X1 U8522 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9653) );
  MUX2_X1 U8523 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9653), .S(n6777), .Z(n9493)
         );
  INV_X1 U8524 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9651) );
  MUX2_X1 U8525 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9651), .S(n9477), .Z(n9481)
         );
  NAND3_X1 U8526 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n9481), .ZN(n9480) );
  OAI21_X1 U8527 ( .B1(n6778), .B2(n9651), .A(n9480), .ZN(n9494) );
  NAND2_X1 U8528 ( .A1(n9493), .A2(n9494), .ZN(n9491) );
  OAI21_X1 U8529 ( .B1(n9497), .B2(n9653), .A(n9491), .ZN(n6797) );
  NAND2_X1 U8530 ( .A1(n6796), .A2(n6797), .ZN(n6795) );
  OAI21_X1 U8531 ( .B1(n9655), .B2(n6800), .A(n6795), .ZN(n6873) );
  INV_X1 U8532 ( .A(n6873), .ZN(n6779) );
  OAI22_X1 U8533 ( .A1(n6874), .A2(n6779), .B1(n9657), .B2(n6872), .ZN(n6803)
         );
  INV_X1 U8534 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6780) );
  MUX2_X1 U8535 ( .A(n6780), .B(P1_REG1_REG_5__SCAN_IN), .S(n6813), .Z(n6804)
         );
  INV_X1 U8536 ( .A(n6804), .ZN(n6781) );
  NAND2_X1 U8537 ( .A1(n6803), .A2(n6781), .ZN(n6782) );
  NAND2_X1 U8538 ( .A1(n6783), .A2(n6782), .ZN(n6786) );
  INV_X1 U8539 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6784) );
  MUX2_X1 U8540 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6784), .S(n6824), .Z(n6785)
         );
  NOR2_X2 U8541 ( .A1(n9472), .A2(n6866), .ZN(n9492) );
  NAND2_X1 U8542 ( .A1(n6785), .A2(n6786), .ZN(n6829) );
  OAI211_X1 U8543 ( .C1(n6786), .C2(n6785), .A(n9492), .B(n6829), .ZN(n6787)
         );
  OAI211_X1 U8544 ( .C1(n9498), .C2(n6830), .A(n6788), .B(n6787), .ZN(n6789)
         );
  OR2_X1 U8545 ( .A1(n6790), .A2(n6789), .ZN(P1_U3249) );
  AOI211_X1 U8546 ( .C1(n6793), .C2(n6792), .A(n6791), .B(n9486), .ZN(n6802)
         );
  AND2_X1 U8547 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6794) );
  AOI21_X1 U8548 ( .B1(n9490), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6794), .ZN(
        n6799) );
  OAI211_X1 U8549 ( .C1(n6797), .C2(n6796), .A(n9492), .B(n6795), .ZN(n6798)
         );
  OAI211_X1 U8550 ( .C1(n9498), .C2(n6800), .A(n6799), .B(n6798), .ZN(n6801)
         );
  OR2_X1 U8551 ( .A1(n6802), .A2(n6801), .ZN(P1_U3246) );
  AND2_X1 U8552 ( .A1(n6751), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8553 ( .A1(n6751), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8554 ( .A1(n6751), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8555 ( .A1(n6751), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8556 ( .A1(n6751), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8557 ( .A1(n6751), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8558 ( .A1(n6751), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8559 ( .A1(n6751), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8560 ( .A1(n6751), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8561 ( .A1(n6751), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8562 ( .A1(n6751), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8563 ( .A1(n6751), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8564 ( .A1(n6751), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8565 ( .A1(n6751), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8566 ( .A1(n6751), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8567 ( .A(n9492), .ZN(n9067) );
  XOR2_X1 U8568 ( .A(n6804), .B(n6803), .Z(n6807) );
  NOR2_X1 U8569 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7130), .ZN(n6805) );
  AOI21_X1 U8570 ( .B1(n9490), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6805), .ZN(
        n6806) );
  OAI21_X1 U8571 ( .B1(n9067), .B2(n6807), .A(n6806), .ZN(n6812) );
  AOI211_X1 U8572 ( .C1(n6810), .C2(n6809), .A(n6808), .B(n9486), .ZN(n6811)
         );
  AOI211_X1 U8573 ( .C1(n9478), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  INV_X1 U8574 ( .A(n6814), .ZN(P1_U3248) );
  NAND2_X1 U8575 ( .A1(n8926), .A2(P1_U3973), .ZN(n6815) );
  OAI21_X1 U8576 ( .B1(n6511), .B2(P1_U3973), .A(n6815), .ZN(P1_U3574) );
  INV_X1 U8577 ( .A(n6816), .ZN(n6818) );
  OAI222_X1 U8578 ( .A1(P2_U3151), .A2(n7587), .B1(n8901), .B2(n6818), .C1(
        n6817), .C2(n8899), .ZN(P2_U3286) );
  INV_X1 U8579 ( .A(n7076), .ZN(n6978) );
  OAI222_X1 U8580 ( .A1(n9450), .A2(n6819), .B1(n9452), .B2(n6818), .C1(n6978), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8581 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6820) );
  OAI222_X1 U8582 ( .A1(P2_U3151), .A2(n7734), .B1(n8901), .B2(n6821), .C1(
        n6820), .C2(n8899), .ZN(P2_U3285) );
  INV_X1 U8583 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6822) );
  INV_X1 U8584 ( .A(n7241), .ZN(n7085) );
  OAI222_X1 U8585 ( .A1(n9450), .A2(n6822), .B1(n9452), .B2(n6821), .C1(n7085), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  AOI21_X1 U8586 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6824), .A(n6823), .ZN(
        n6827) );
  NAND2_X1 U8587 ( .A1(n6906), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6825) );
  OAI21_X1 U8588 ( .B1(n6906), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6825), .ZN(
        n6826) );
  NOR2_X1 U8589 ( .A1(n6827), .A2(n6826), .ZN(n6902) );
  AOI211_X1 U8590 ( .C1(n6827), .C2(n6826), .A(n6902), .B(n9486), .ZN(n6838)
         );
  NOR2_X1 U8591 ( .A1(n6828), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7182) );
  AOI21_X1 U8592 ( .B1(n9490), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7182), .ZN(
        n6835) );
  OAI21_X1 U8593 ( .B1(n6830), .B2(n6784), .A(n6829), .ZN(n6833) );
  INV_X1 U8594 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6831) );
  MUX2_X1 U8595 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6831), .S(n6906), .Z(n6832)
         );
  NAND2_X1 U8596 ( .A1(n6832), .A2(n6833), .ZN(n6907) );
  OAI211_X1 U8597 ( .C1(n6833), .C2(n6832), .A(n9492), .B(n6907), .ZN(n6834)
         );
  OAI211_X1 U8598 ( .C1(n9498), .C2(n6836), .A(n6835), .B(n6834), .ZN(n6837)
         );
  OR2_X1 U8599 ( .A1(n6838), .A2(n6837), .ZN(P1_U3250) );
  INV_X1 U8600 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9479) );
  INV_X1 U8601 ( .A(n7351), .ZN(n6839) );
  OAI21_X1 U8602 ( .B1(n9541), .B2(n9635), .A(n6839), .ZN(n6840) );
  NAND2_X1 U8603 ( .A1(n9047), .A2(n8983), .ZN(n7352) );
  OAI211_X1 U8604 ( .C1(n6842), .C2(n6841), .A(n6840), .B(n7352), .ZN(n6844)
         );
  NAND2_X1 U8605 ( .A1(n6844), .A2(n10083), .ZN(n6843) );
  OAI21_X1 U8606 ( .B1(n10083), .B2(n9479), .A(n6843), .ZN(P1_U3522) );
  INV_X1 U8607 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8608 ( .A1(n6844), .A2(n9650), .ZN(n6845) );
  OAI21_X1 U8609 ( .B1(n9650), .B2(n6846), .A(n6845), .ZN(P1_U3453) );
  INV_X1 U8610 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6856) );
  MUX2_X1 U8611 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n6847), .Z(n6849) );
  AOI21_X1 U8612 ( .B1(n6850), .B2(n6849), .A(n6848), .ZN(n6851) );
  AOI21_X1 U8613 ( .B1(n6852), .B2(n9763), .A(n6851), .ZN(n6853) );
  AOI21_X1 U8614 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6853), .ZN(
        n6855) );
  OAI211_X1 U8615 ( .C1(n9737), .C2(n6856), .A(n6855), .B(n6854), .ZN(P2_U3182) );
  NAND2_X1 U8616 ( .A1(n7433), .A2(P2_U3893), .ZN(n6857) );
  OAI21_X1 U8617 ( .B1(P2_U3893), .B2(n6858), .A(n6857), .ZN(P2_U3497) );
  INV_X1 U8618 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6860) );
  INV_X1 U8619 ( .A(n6859), .ZN(n6862) );
  INV_X1 U8620 ( .A(n7242), .ZN(n7286) );
  OAI222_X1 U8621 ( .A1(n9450), .A2(n6860), .B1(n9452), .B2(n6862), .C1(
        P1_U3086), .C2(n7286), .ZN(P1_U3344) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6861) );
  OAI222_X1 U8623 ( .A1(n8073), .A2(P2_U3151), .B1(n8901), .B2(n6862), .C1(
        n6861), .C2(n8899), .ZN(P2_U3284) );
  OAI21_X1 U8624 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6922) );
  INV_X1 U8625 ( .A(n9475), .ZN(n6867) );
  MUX2_X1 U8626 ( .A(n6922), .B(n6867), .S(n6866), .Z(n6870) );
  NOR2_X1 U8627 ( .A1(n4294), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6868) );
  NOR2_X1 U8628 ( .A1(n5605), .A2(n6868), .ZN(n9465) );
  NOR2_X1 U8629 ( .A1(n9465), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9463) );
  AOI211_X1 U8630 ( .C1(n6870), .C2(n6869), .A(n9463), .B(n9046), .ZN(n9501)
         );
  NAND2_X1 U8631 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8632 ( .A1(n9490), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6871) );
  OAI211_X1 U8633 ( .C1(n9498), .C2(n6872), .A(n7067), .B(n6871), .ZN(n6881)
         );
  XOR2_X1 U8634 ( .A(n6874), .B(n6873), .Z(n6879) );
  OAI211_X1 U8635 ( .C1(n6877), .C2(n6876), .A(n9116), .B(n6875), .ZN(n6878)
         );
  OAI21_X1 U8636 ( .B1(n6879), .B2(n9067), .A(n6878), .ZN(n6880) );
  OR3_X1 U8637 ( .A1(n9501), .A2(n6881), .A3(n6880), .ZN(P1_U3247) );
  OAI21_X1 U8638 ( .B1(n6884), .B2(n6883), .A(n6882), .ZN(n6885) );
  NAND2_X1 U8639 ( .A1(n6885), .A2(n9822), .ZN(n6895) );
  INV_X1 U8640 ( .A(n7012), .ZN(n6886) );
  AOI21_X1 U8641 ( .B1(n9895), .B2(n6887), .A(n6886), .ZN(n6888) );
  NAND2_X1 U8642 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n7222) );
  OAI21_X1 U8643 ( .B1(n9826), .B2(n6888), .A(n7222), .ZN(n6893) );
  NAND2_X1 U8644 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  AOI21_X1 U8645 ( .B1(n7019), .B2(n6891), .A(n9817), .ZN(n6892) );
  AOI211_X1 U8646 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9808), .A(n6893), .B(
        n6892), .ZN(n6894) );
  OAI211_X1 U8647 ( .C1(n9807), .C2(n6896), .A(n6895), .B(n6894), .ZN(P2_U3185) );
  XOR2_X1 U8648 ( .A(n6898), .B(n6897), .Z(n6901) );
  NAND2_X1 U8649 ( .A1(n8998), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6921) );
  AOI22_X1 U8650 ( .A1(n8982), .A2(n9047), .B1(n9045), .B2(n8983), .ZN(n7563)
         );
  OAI22_X1 U8651 ( .A1(n5151), .A2(n9017), .B1(n9011), .B2(n7563), .ZN(n6899)
         );
  AOI21_X1 U8652 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6921), .A(n6899), .ZN(
        n6900) );
  OAI21_X1 U8653 ( .B1(n6901), .B2(n8988), .A(n6900), .ZN(P1_U3237) );
  NAND2_X1 U8654 ( .A1(n6973), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6903) );
  OAI21_X1 U8655 ( .B1(n6973), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6903), .ZN(
        n6904) );
  AOI211_X1 U8656 ( .C1(n6905), .C2(n6904), .A(n6972), .B(n9486), .ZN(n6916)
         );
  NAND2_X1 U8657 ( .A1(n6906), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U8658 ( .A1(n6908), .A2(n6907), .ZN(n6911) );
  INV_X1 U8659 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6909) );
  MUX2_X1 U8660 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6909), .S(n6973), .Z(n6910)
         );
  NAND2_X1 U8661 ( .A1(n6910), .A2(n6911), .ZN(n6967) );
  OAI211_X1 U8662 ( .C1(n6911), .C2(n6910), .A(n9492), .B(n6967), .ZN(n6913)
         );
  AND2_X1 U8663 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7404) );
  AOI21_X1 U8664 ( .B1(n9490), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7404), .ZN(
        n6912) );
  OAI211_X1 U8665 ( .C1(n9498), .C2(n6914), .A(n6913), .B(n6912), .ZN(n6915)
         );
  OR2_X1 U8666 ( .A1(n6916), .A2(n6915), .ZN(P1_U3251) );
  OAI222_X1 U8667 ( .A1(n6918), .A2(P2_U3151), .B1(n8899), .B2(n6917), .C1(
        n6919), .C2(n8906), .ZN(P2_U3283) );
  INV_X1 U8668 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6920) );
  INV_X1 U8669 ( .A(n7386), .ZN(n7391) );
  OAI222_X1 U8670 ( .A1(n9450), .A2(n6920), .B1(n9452), .B2(n6919), .C1(n7391), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8671 ( .A(n6921), .ZN(n6960) );
  INV_X1 U8672 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6925) );
  OAI22_X1 U8673 ( .A1(n8988), .A2(n6922), .B1(n9011), .B2(n7352), .ZN(n6923)
         );
  AOI21_X1 U8674 ( .B1(n9548), .B2(n8968), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8675 ( .B1(n6960), .B2(n6925), .A(n6924), .ZN(P1_U3232) );
  INV_X1 U8676 ( .A(n7042), .ZN(n6926) );
  NAND2_X1 U8677 ( .A1(n6931), .A2(n6926), .ZN(n6994) );
  INV_X1 U8678 ( .A(n6928), .ZN(n6929) );
  NAND2_X1 U8679 ( .A1(n6935), .A2(n6929), .ZN(n6933) );
  INV_X1 U8680 ( .A(n6944), .ZN(n6930) );
  NAND2_X1 U8681 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  AND2_X1 U8682 ( .A1(n8532), .A2(n7055), .ZN(n8182) );
  INV_X1 U8683 ( .A(n8182), .ZN(n6934) );
  NAND2_X1 U8684 ( .A1(n8181), .A2(n6934), .ZN(n8345) );
  NAND2_X1 U8685 ( .A1(n6935), .A2(n9890), .ZN(n6938) );
  INV_X1 U8686 ( .A(n6936), .ZN(n6937) );
  AOI22_X1 U8687 ( .A1(n8508), .A2(n8345), .B1(n6939), .B2(n8501), .ZN(n6952)
         );
  NAND2_X1 U8688 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  OAI211_X1 U8689 ( .C1(n6947), .C2(n6944), .A(n6943), .B(n6942), .ZN(n6945)
         );
  NAND2_X1 U8690 ( .A1(n6945), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6949) );
  OR2_X1 U8691 ( .A1(n6946), .A2(n7042), .ZN(n8386) );
  OR2_X1 U8692 ( .A1(n6947), .A2(n8386), .ZN(n6948) );
  AND2_X1 U8693 ( .A1(n6949), .A2(n6948), .ZN(n7117) );
  NAND2_X1 U8694 ( .A1(n7117), .A2(n6950), .ZN(n7038) );
  NAND2_X1 U8695 ( .A1(n7038), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6951) );
  OAI211_X1 U8696 ( .C1(n7030), .C2(n8512), .A(n6952), .B(n6951), .ZN(P2_U3172) );
  INV_X1 U8697 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6959) );
  INV_X1 U8698 ( .A(n8982), .ZN(n8993) );
  OAI22_X1 U8699 ( .A1(n4727), .A2(n8993), .B1(n5150), .B2(n8995), .ZN(n9539)
         );
  AOI22_X1 U8700 ( .A1(n8968), .A2(n9549), .B1(n9001), .B2(n9539), .ZN(n6958)
         );
  OAI21_X1 U8701 ( .B1(n6953), .B2(n6955), .A(n6954), .ZN(n6956) );
  NAND2_X1 U8702 ( .A1(n6956), .A2(n9007), .ZN(n6957) );
  OAI211_X1 U8703 ( .C1(n6960), .C2(n6959), .A(n6958), .B(n6957), .ZN(P1_U3222) );
  XOR2_X1 U8704 ( .A(n6962), .B(n6961), .Z(n6966) );
  OAI22_X1 U8705 ( .A1(n5150), .A2(n8993), .B1(n4462), .B2(n8995), .ZN(n9522)
         );
  AOI22_X1 U8706 ( .A1(n8968), .A2(n6963), .B1(n9001), .B2(n9522), .ZN(n6965)
         );
  MUX2_X1 U8707 ( .A(n8998), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6964) );
  OAI211_X1 U8708 ( .C1(n6966), .C2(n8988), .A(n6965), .B(n6964), .ZN(P1_U3218) );
  INV_X1 U8709 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9662) );
  AOI22_X1 U8710 ( .A1(n7076), .A2(n9662), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6978), .ZN(n6970) );
  NAND2_X1 U8711 ( .A1(n6973), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U8712 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  NOR2_X1 U8713 ( .A1(n6970), .A2(n6969), .ZN(n7078) );
  AOI21_X1 U8714 ( .B1(n6970), .B2(n6969), .A(n7078), .ZN(n6982) );
  INV_X1 U8715 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U8716 ( .A1(n7076), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6971), .B2(
        n6978), .ZN(n6975) );
  OAI21_X1 U8717 ( .B1(n6975), .B2(n6974), .A(n7073), .ZN(n6976) );
  NAND2_X1 U8718 ( .A1(n6976), .A2(n9116), .ZN(n6981) );
  NOR2_X1 U8719 ( .A1(n6977), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7481) );
  NOR2_X1 U8720 ( .A1(n9498), .A2(n6978), .ZN(n6979) );
  AOI211_X1 U8721 ( .C1(n9490), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7481), .B(
        n6979), .ZN(n6980) );
  OAI211_X1 U8722 ( .C1(n6982), .C2(n9067), .A(n6981), .B(n6980), .ZN(P1_U3252) );
  OAI21_X1 U8723 ( .B1(n9844), .B2(n9865), .A(n8345), .ZN(n6983) );
  NAND2_X1 U8724 ( .A1(n4293), .A2(n9841), .ZN(n7049) );
  OAI211_X1 U8725 ( .C1(n9873), .C2(n7055), .A(n6983), .B(n7049), .ZN(n7001)
         );
  NAND2_X1 U8726 ( .A1(n7001), .A2(n9904), .ZN(n6984) );
  OAI21_X1 U8727 ( .B1(n9904), .B2(n5782), .A(n6984), .ZN(P2_U3459) );
  INV_X1 U8728 ( .A(n6985), .ZN(n6986) );
  AND2_X1 U8729 ( .A1(n6988), .A2(n7156), .ZN(n6989) );
  NAND2_X1 U8730 ( .A1(n7795), .A2(n7055), .ZN(n6991) );
  NAND2_X1 U8731 ( .A1(n8181), .A2(n6991), .ZN(n7028) );
  INV_X1 U8732 ( .A(n6992), .ZN(n6995) );
  XNOR2_X1 U8733 ( .A(n7029), .B(n4293), .ZN(n7027) );
  XOR2_X1 U8734 ( .A(n7028), .B(n7027), .Z(n6999) );
  AOI22_X1 U8735 ( .A1(n8510), .A2(n8532), .B1(n8501), .B2(n6995), .ZN(n6996)
         );
  OAI21_X1 U8736 ( .B1(n7033), .B2(n8512), .A(n6996), .ZN(n6997) );
  AOI21_X1 U8737 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7038), .A(n6997), .ZN(
        n6998) );
  OAI21_X1 U8738 ( .B1(n8503), .B2(n6999), .A(n6998), .ZN(P2_U3162) );
  INV_X1 U8739 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7000) );
  INV_X1 U8740 ( .A(n7667), .ZN(n7673) );
  OAI222_X1 U8741 ( .A1(n9450), .A2(n7000), .B1(n9452), .B2(n8120), .C1(n7673), 
        .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U8742 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U8743 ( .A1(n7001), .A2(n9891), .ZN(n7002) );
  OAI21_X1 U8744 ( .B1(n9891), .B2(n10034), .A(n7002), .ZN(P2_U3390) );
  AOI211_X1 U8745 ( .C1(n7005), .C2(n7004), .A(n9763), .B(n7003), .ZN(n7006)
         );
  INV_X1 U8746 ( .A(n7006), .ZN(n7025) );
  INV_X1 U8747 ( .A(n7007), .ZN(n7009) );
  NOR2_X1 U8748 ( .A1(n7009), .A2(n7008), .ZN(n7013) );
  INV_X1 U8749 ( .A(n7010), .ZN(n7011) );
  AOI21_X1 U8750 ( .B1(n7013), .B2(n7012), .A(n7011), .ZN(n7015) );
  NAND2_X1 U8751 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3151), .ZN(n7014) );
  OAI21_X1 U8752 ( .B1(n9826), .B2(n7015), .A(n7014), .ZN(n7023) );
  INV_X1 U8753 ( .A(n7016), .ZN(n7018) );
  NAND3_X1 U8754 ( .A1(n7019), .A2(n7018), .A3(n7017), .ZN(n7020) );
  AOI21_X1 U8755 ( .B1(n7021), .B2(n7020), .A(n9817), .ZN(n7022) );
  AOI211_X1 U8756 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9808), .A(n7023), .B(
        n7022), .ZN(n7024) );
  OAI211_X1 U8757 ( .C1(n9807), .C2(n7026), .A(n7025), .B(n7024), .ZN(P2_U3186) );
  NAND2_X1 U8758 ( .A1(n7028), .A2(n7027), .ZN(n7032) );
  NAND2_X1 U8759 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  NAND2_X1 U8760 ( .A1(n7032), .A2(n7031), .ZN(n7227) );
  XNOR2_X1 U8761 ( .A(n7105), .B(n7033), .ZN(n7226) );
  XOR2_X1 U8762 ( .A(n7227), .B(n7226), .Z(n7040) );
  AOI22_X1 U8763 ( .A1(n8510), .A2(n4293), .B1(n8501), .B2(n7034), .ZN(n7035)
         );
  OAI21_X1 U8764 ( .B1(n7036), .B2(n8512), .A(n7035), .ZN(n7037) );
  AOI21_X1 U8765 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7038), .A(n7037), .ZN(
        n7039) );
  OAI21_X1 U8766 ( .B1(n7040), .B2(n8503), .A(n7039), .ZN(P2_U3177) );
  NAND2_X1 U8767 ( .A1(n8557), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7041) );
  OAI21_X1 U8768 ( .B1(n8600), .B2(n8557), .A(n7041), .ZN(P2_U3520) );
  NAND3_X1 U8769 ( .A1(n8345), .A2(n7042), .A3(n9873), .ZN(n7050) );
  INV_X1 U8770 ( .A(n7043), .ZN(n7044) );
  OAI21_X1 U8771 ( .B1(n7046), .B2(n7045), .A(n7044), .ZN(n7047) );
  AOI21_X1 U8772 ( .B1(n7050), .B2(n7049), .A(n8586), .ZN(n7058) );
  NOR2_X1 U8773 ( .A1(n8752), .A2(n5783), .ZN(n7057) );
  INV_X1 U8774 ( .A(n7051), .ZN(n7053) );
  INV_X1 U8775 ( .A(n9836), .ZN(n7052) );
  INV_X1 U8776 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7054) );
  OAI22_X1 U8777 ( .A1(n8581), .A2(n7055), .B1(n7054), .B2(n9834), .ZN(n7056)
         );
  OR3_X1 U8778 ( .A1(n7058), .A2(n7057), .A3(n7056), .ZN(P2_U3233) );
  XNOR2_X1 U8779 ( .A(n7060), .B(n7059), .ZN(n7066) );
  NAND2_X1 U8780 ( .A1(n7061), .A2(n7062), .ZN(n7065) );
  INV_X1 U8781 ( .A(n7063), .ZN(n7064) );
  AOI211_X1 U8782 ( .C1(n7066), .C2(n7065), .A(n8988), .B(n7064), .ZN(n7071)
         );
  AOI22_X1 U8783 ( .A1(n8982), .A2(n9045), .B1(n9043), .B2(n8983), .ZN(n7318)
         );
  OAI21_X1 U8784 ( .B1(n9011), .B2(n7318), .A(n7067), .ZN(n7070) );
  INV_X1 U8785 ( .A(n7068), .ZN(n7322) );
  OAI22_X1 U8786 ( .A1(n9017), .A2(n7323), .B1(n8998), .B2(n7322), .ZN(n7069)
         );
  OR3_X1 U8787 ( .A1(n7071), .A2(n7070), .A3(n7069), .ZN(P1_U3230) );
  NAND2_X1 U8788 ( .A1(n7241), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7072) );
  OAI21_X1 U8789 ( .B1(n7241), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7072), .ZN(
        n7075) );
  OAI21_X1 U8790 ( .B1(n7076), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7073), .ZN(
        n7074) );
  NOR2_X1 U8791 ( .A1(n7075), .A2(n7074), .ZN(n7240) );
  AOI211_X1 U8792 ( .C1(n7075), .C2(n7074), .A(n7240), .B(n9486), .ZN(n7087)
         );
  NOR2_X1 U8793 ( .A1(n7076), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U8794 ( .A1(n7078), .A2(n7077), .ZN(n7081) );
  INV_X1 U8795 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7079) );
  MUX2_X1 U8796 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7079), .S(n7241), .Z(n7080)
         );
  NAND2_X1 U8797 ( .A1(n7080), .A2(n7081), .ZN(n7235) );
  OAI211_X1 U8798 ( .C1(n7081), .C2(n7080), .A(n7235), .B(n9492), .ZN(n7084)
         );
  AND2_X1 U8799 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7082) );
  AOI21_X1 U8800 ( .B1(n9490), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7082), .ZN(
        n7083) );
  OAI211_X1 U8801 ( .C1(n9498), .C2(n7085), .A(n7084), .B(n7083), .ZN(n7086)
         );
  OR2_X1 U8802 ( .A1(n7087), .A2(n7086), .ZN(P1_U3253) );
  XNOR2_X1 U8803 ( .A(n7088), .B(n7089), .ZN(n7461) );
  XNOR2_X1 U8804 ( .A(n7090), .B(n7089), .ZN(n7093) );
  NAND2_X1 U8805 ( .A1(n9044), .A2(n8982), .ZN(n7092) );
  NAND2_X1 U8806 ( .A1(n9042), .A2(n8983), .ZN(n7091) );
  NAND2_X1 U8807 ( .A1(n7092), .A2(n7091), .ZN(n7128) );
  AOI21_X1 U8808 ( .B1(n7093), .B2(n9541), .A(n7128), .ZN(n7463) );
  OAI211_X1 U8809 ( .C1(n7131), .C2(n4318), .A(n4523), .B(n9551), .ZN(n7459)
         );
  OAI211_X1 U8810 ( .C1(n7131), .C2(n9632), .A(n7463), .B(n7459), .ZN(n7094)
         );
  AOI21_X1 U8811 ( .B1(n9635), .B2(n7461), .A(n7094), .ZN(n10081) );
  NAND2_X1 U8812 ( .A1(n9648), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7095) );
  OAI21_X1 U8813 ( .B1(n10081), .B2(n9648), .A(n7095), .ZN(P1_U3468) );
  INV_X1 U8814 ( .A(n7096), .ZN(n7098) );
  INV_X1 U8815 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7097) );
  OAI222_X1 U8816 ( .A1(n9790), .A2(P2_U3151), .B1(n8901), .B2(n7098), .C1(
        n7097), .C2(n8899), .ZN(P2_U3281) );
  INV_X1 U8817 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7099) );
  INV_X1 U8818 ( .A(n7884), .ZN(n7889) );
  OAI222_X1 U8819 ( .A1(n8108), .A2(n7099), .B1(n9452), .B2(n7098), .C1(
        P1_U3086), .C2(n7889), .ZN(P1_U3341) );
  INV_X1 U8820 ( .A(n7100), .ZN(n7103) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7101) );
  OAI222_X1 U8822 ( .A1(n7102), .A2(P2_U3151), .B1(n8901), .B2(n7103), .C1(
        n7101), .C2(n8899), .ZN(P2_U3280) );
  INV_X1 U8823 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7104) );
  OAI222_X1 U8824 ( .A1(n8108), .A2(n7104), .B1(n9452), .B2(n7103), .C1(
        P1_U3086), .C2(n9055), .ZN(P1_U3340) );
  INV_X1 U8825 ( .A(n7228), .ZN(n7107) );
  XNOR2_X1 U8826 ( .A(n7106), .B(n9842), .ZN(n7225) );
  NAND2_X1 U8827 ( .A1(n7106), .A2(n9842), .ZN(n7108) );
  OAI21_X1 U8828 ( .B1(n7107), .B2(n7225), .A(n7108), .ZN(n7111) );
  AND2_X1 U8829 ( .A1(n7226), .A2(n7108), .ZN(n7109) );
  NAND2_X1 U8830 ( .A1(n7109), .A2(n7227), .ZN(n7110) );
  NAND2_X1 U8831 ( .A1(n7111), .A2(n7110), .ZN(n7113) );
  INV_X2 U8832 ( .A(n7112), .ZN(n7795) );
  XNOR2_X1 U8833 ( .A(n9863), .B(n7112), .ZN(n7142) );
  XNOR2_X1 U8834 ( .A(n7147), .B(n7142), .ZN(n7114) );
  NAND2_X1 U8835 ( .A1(n7113), .A2(n7114), .ZN(n7145) );
  OAI21_X1 U8836 ( .B1(n7113), .B2(n7114), .A(n7145), .ZN(n7122) );
  INV_X1 U8837 ( .A(n7115), .ZN(n7206) );
  NAND2_X1 U8838 ( .A1(n7116), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8390) );
  INV_X1 U8839 ( .A(n8514), .ZN(n8466) );
  AOI22_X1 U8840 ( .A1(n8496), .A2(n8530), .B1(n8510), .B2(n9842), .ZN(n7120)
         );
  AOI22_X1 U8841 ( .A1(n8501), .A2(n7118), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3151), .ZN(n7119) );
  OAI211_X1 U8842 ( .C1(n7206), .C2(n8466), .A(n7120), .B(n7119), .ZN(n7121)
         );
  AOI21_X1 U8843 ( .B1(n7122), .B2(n8508), .A(n7121), .ZN(n7123) );
  INV_X1 U8844 ( .A(n7123), .ZN(P2_U3170) );
  INV_X1 U8845 ( .A(n7125), .ZN(n7165) );
  NAND2_X1 U8846 ( .A1(n7124), .A2(n7165), .ZN(n7126) );
  XOR2_X1 U8847 ( .A(n7127), .B(n7126), .Z(n7135) );
  NAND2_X1 U8848 ( .A1(n9001), .A2(n7128), .ZN(n7129) );
  OAI21_X1 U8849 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7130), .A(n7129), .ZN(n7133) );
  NOR2_X1 U8850 ( .A1(n9017), .A2(n7131), .ZN(n7132) );
  AOI211_X1 U8851 ( .C1(n9013), .C2(n7455), .A(n7133), .B(n7132), .ZN(n7134)
         );
  OAI21_X1 U8852 ( .B1(n7135), .B2(n8988), .A(n7134), .ZN(P1_U3227) );
  XNOR2_X1 U8853 ( .A(n8346), .B(n8181), .ZN(n7155) );
  OAI21_X1 U8854 ( .B1(n7137), .B2(n8346), .A(n7136), .ZN(n7139) );
  AOI222_X1 U8855 ( .A1(n9844), .A2(n7139), .B1(n7138), .B2(n9841), .C1(n8532), 
        .C2(n9840), .ZN(n7159) );
  OAI21_X1 U8856 ( .B1(n6992), .B2(n9873), .A(n7159), .ZN(n7140) );
  AOI21_X1 U8857 ( .B1(n9865), .B2(n7155), .A(n7140), .ZN(n9851) );
  NAND2_X1 U8858 ( .A1(n9902), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U8859 ( .B1(n9851), .B2(n9902), .A(n7141), .ZN(P2_U3460) );
  INV_X1 U8860 ( .A(n7142), .ZN(n7143) );
  NAND2_X1 U8861 ( .A1(n7147), .A2(n7143), .ZN(n7144) );
  NAND2_X1 U8862 ( .A1(n7145), .A2(n7144), .ZN(n7329) );
  XNOR2_X1 U8863 ( .A(n8161), .B(n7271), .ZN(n7330) );
  XNOR2_X1 U8864 ( .A(n7330), .B(n8530), .ZN(n7328) );
  XOR2_X1 U8865 ( .A(n7329), .B(n7328), .Z(n7150) );
  AOI22_X1 U8866 ( .A1(n8496), .A2(n7433), .B1(n8501), .B2(n7271), .ZN(n7146)
         );
  NAND2_X1 U8867 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n9724) );
  OAI211_X1 U8868 ( .C1(n7147), .C2(n8499), .A(n7146), .B(n9724), .ZN(n7148)
         );
  AOI21_X1 U8869 ( .B1(n7267), .B2(n8514), .A(n7148), .ZN(n7149) );
  OAI21_X1 U8870 ( .B1(n7150), .B2(n8503), .A(n7149), .ZN(P2_U3167) );
  INV_X1 U8871 ( .A(n7151), .ZN(n7153) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7152) );
  OAI222_X1 U8873 ( .A1(P2_U3151), .A2(n9806), .B1(n8901), .B2(n7153), .C1(
        n7152), .C2(n8899), .ZN(P2_U3279) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7154) );
  INV_X1 U8875 ( .A(n9070), .ZN(n9078) );
  OAI222_X1 U8876 ( .A1(n8108), .A2(n7154), .B1(n9452), .B2(n7153), .C1(n9078), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8877 ( .A(n7155), .ZN(n7163) );
  OR2_X1 U8878 ( .A1(n7156), .A2(n7559), .ZN(n7255) );
  NAND2_X1 U8879 ( .A1(n9832), .A2(n7255), .ZN(n7157) );
  INV_X1 U8880 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7158) );
  OAI22_X1 U8881 ( .A1(n8581), .A2(n6992), .B1(n7158), .B2(n9834), .ZN(n7161)
         );
  NOR2_X1 U8882 ( .A1(n7159), .A2(n8586), .ZN(n7160) );
  AOI211_X1 U8883 ( .C1(n8586), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7161), .B(
        n7160), .ZN(n7162) );
  OAI21_X1 U8884 ( .B1(n7163), .B2(n8741), .A(n7162), .ZN(P2_U3232) );
  NAND2_X1 U8885 ( .A1(n7164), .A2(n7165), .ZN(n7167) );
  NAND2_X1 U8886 ( .A1(n7167), .A2(n7166), .ZN(n7168) );
  AOI21_X1 U8887 ( .B1(n7169), .B2(n7168), .A(n8988), .ZN(n7175) );
  NAND2_X1 U8888 ( .A1(n9043), .A2(n8982), .ZN(n7171) );
  NAND2_X1 U8889 ( .A1(n9041), .A2(n8983), .ZN(n7170) );
  NAND2_X1 U8890 ( .A1(n7171), .A2(n7170), .ZN(n7443) );
  AOI22_X1 U8891 ( .A1(n9001), .A2(n7443), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7173) );
  NAND2_X1 U8892 ( .A1(n9013), .A2(n7449), .ZN(n7172) );
  OAI211_X1 U8893 ( .C1(n9017), .C2(n9589), .A(n7173), .B(n7172), .ZN(n7174)
         );
  OR2_X1 U8894 ( .A1(n7175), .A2(n7174), .ZN(P1_U3239) );
  XOR2_X1 U8895 ( .A(n7178), .B(n7177), .Z(n7179) );
  XNOR2_X1 U8896 ( .A(n7176), .B(n7179), .ZN(n7186) );
  NAND2_X1 U8897 ( .A1(n9042), .A2(n8982), .ZN(n7181) );
  NAND2_X1 U8898 ( .A1(n9040), .A2(n8983), .ZN(n7180) );
  NAND2_X1 U8899 ( .A1(n7181), .A2(n7180), .ZN(n9509) );
  AOI21_X1 U8900 ( .B1(n9001), .B2(n9509), .A(n7182), .ZN(n7184) );
  NAND2_X1 U8901 ( .A1(n9013), .A2(n9510), .ZN(n7183) );
  OAI211_X1 U8902 ( .C1(n9017), .C2(n9593), .A(n7184), .B(n7183), .ZN(n7185)
         );
  AOI21_X1 U8903 ( .B1(n7186), .B2(n9007), .A(n7185), .ZN(n7187) );
  INV_X1 U8904 ( .A(n7187), .ZN(P1_U3213) );
  AOI21_X1 U8905 ( .B1(n7190), .B2(n7189), .A(n7188), .ZN(n7199) );
  XNOR2_X1 U8906 ( .A(n7191), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7197) );
  OAI21_X1 U8907 ( .B1(n4392), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9754), .ZN(
        n7192) );
  INV_X1 U8908 ( .A(n9826), .ZN(n9758) );
  NAND2_X1 U8909 ( .A1(n7192), .A2(n9758), .ZN(n7194) );
  AND2_X1 U8910 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7364) );
  AOI21_X1 U8911 ( .B1(n9808), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7364), .ZN(
        n7193) );
  OAI211_X1 U8912 ( .C1(n9807), .C2(n7195), .A(n7194), .B(n7193), .ZN(n7196)
         );
  AOI21_X1 U8913 ( .B1(n9768), .B2(n7197), .A(n7196), .ZN(n7198) );
  OAI21_X1 U8914 ( .B1(n7199), .B2(n9763), .A(n7198), .ZN(P2_U3189) );
  AND2_X1 U8915 ( .A1(n7200), .A2(n7258), .ZN(n7204) );
  NAND2_X1 U8916 ( .A1(n7201), .A2(n8343), .ZN(n7217) );
  NAND3_X1 U8917 ( .A1(n7217), .A2(n6618), .A3(n7202), .ZN(n7203) );
  NAND2_X1 U8918 ( .A1(n7204), .A2(n7203), .ZN(n7205) );
  AOI222_X1 U8919 ( .A1(n9844), .A2(n7205), .B1(n9842), .B2(n9840), .C1(n8530), 
        .C2(n9841), .ZN(n9862) );
  OAI22_X1 U8920 ( .A1(n8581), .A2(n9863), .B1(n7206), .B2(n9834), .ZN(n7207)
         );
  AOI21_X1 U8921 ( .B1(n8586), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7207), .ZN(
        n7210) );
  XNOR2_X1 U8922 ( .A(n7208), .B(n6618), .ZN(n9866) );
  INV_X1 U8923 ( .A(n8741), .ZN(n8759) );
  NAND2_X1 U8924 ( .A1(n9866), .A2(n8759), .ZN(n7209) );
  OAI211_X1 U8925 ( .C1(n9862), .C2(n8586), .A(n7210), .B(n7209), .ZN(P2_U3229) );
  OAI21_X1 U8926 ( .B1(n7212), .B2(n7215), .A(n7211), .ZN(n9858) );
  INV_X1 U8927 ( .A(n9858), .ZN(n7221) );
  NAND3_X1 U8928 ( .A1(n7213), .A2(n7215), .A3(n7214), .ZN(n7216) );
  NAND2_X1 U8929 ( .A1(n7217), .A2(n7216), .ZN(n7218) );
  AOI222_X1 U8930 ( .A1(n9844), .A2(n7218), .B1(n8531), .B2(n9841), .C1(n7138), 
        .C2(n9840), .ZN(n9860) );
  MUX2_X1 U8931 ( .A(n6889), .B(n9860), .S(n8752), .Z(n7220) );
  INV_X1 U8932 ( .A(n7224), .ZN(n9857) );
  INV_X1 U8933 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7233) );
  AOI22_X1 U8934 ( .A1(n8756), .A2(n9857), .B1(n7233), .B2(n8755), .ZN(n7219)
         );
  OAI211_X1 U8935 ( .C1(n7221), .C2(n8741), .A(n7220), .B(n7219), .ZN(P2_U3230) );
  INV_X1 U8936 ( .A(n8501), .ZN(n8517) );
  AOI22_X1 U8937 ( .A1(n8510), .A2(n7138), .B1(n8496), .B2(n8531), .ZN(n7223)
         );
  OAI211_X1 U8938 ( .C1(n7224), .C2(n8517), .A(n7223), .B(n7222), .ZN(n7232)
         );
  NAND2_X1 U8939 ( .A1(n7227), .A2(n7226), .ZN(n7229) );
  NAND2_X1 U8940 ( .A1(n7229), .A2(n7228), .ZN(n7230) );
  AOI211_X1 U8941 ( .C1(n7225), .C2(n7230), .A(n8503), .B(n4389), .ZN(n7231)
         );
  AOI211_X1 U8942 ( .C1(n7233), .C2(n8514), .A(n7232), .B(n7231), .ZN(n7234)
         );
  INV_X1 U8943 ( .A(n7234), .ZN(P2_U3158) );
  INV_X1 U8944 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U8945 ( .A1(n7241), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8946 ( .A1(n7236), .A2(n7235), .ZN(n7280) );
  NAND2_X1 U8947 ( .A1(n7242), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7237) );
  OAI211_X1 U8948 ( .C1(n7242), .C2(P1_REG1_REG_11__SCAN_IN), .A(n7280), .B(
        n7237), .ZN(n7283) );
  OAI21_X1 U8949 ( .B1(n10050), .B2(n7286), .A(n7283), .ZN(n7239) );
  INV_X1 U8950 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U8951 ( .A1(n7386), .A2(n9666), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n7391), .ZN(n7238) );
  NOR2_X1 U8952 ( .A1(n7239), .A2(n7238), .ZN(n7390) );
  AOI21_X1 U8953 ( .B1(n7239), .B2(n7238), .A(n7390), .ZN(n7253) );
  AOI21_X1 U8954 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7241), .A(n7240), .ZN(
        n7277) );
  NAND2_X1 U8955 ( .A1(n7242), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7244) );
  OR2_X1 U8956 ( .A1(n7242), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7243) );
  NAND2_X1 U8957 ( .A1(n7244), .A2(n7243), .ZN(n7276) );
  NOR2_X1 U8958 ( .A1(n7386), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7245) );
  AOI21_X1 U8959 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7386), .A(n7245), .ZN(
        n7246) );
  NAND2_X1 U8960 ( .A1(n7246), .A2(n7247), .ZN(n7385) );
  OAI21_X1 U8961 ( .B1(n7247), .B2(n7246), .A(n7385), .ZN(n7248) );
  NAND2_X1 U8962 ( .A1(n7248), .A2(n9116), .ZN(n7252) );
  INV_X1 U8963 ( .A(n9490), .ZN(n9122) );
  INV_X1 U8964 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U8965 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7660) );
  OAI21_X1 U8966 ( .B1(n9122), .B2(n7249), .A(n7660), .ZN(n7250) );
  AOI21_X1 U8967 ( .B1(n7386), .B2(n9478), .A(n7250), .ZN(n7251) );
  OAI211_X1 U8968 ( .C1(n7253), .C2(n9067), .A(n7252), .B(n7251), .ZN(P1_U3255) );
  XNOR2_X1 U8969 ( .A(n8530), .B(n9868), .ZN(n8352) );
  XNOR2_X1 U8970 ( .A(n7254), .B(n8352), .ZN(n9869) );
  NOR2_X1 U8971 ( .A1(n8586), .A2(n7255), .ZN(n9848) );
  INV_X1 U8972 ( .A(n9848), .ZN(n7697) );
  AOI22_X1 U8973 ( .A1(n8531), .A2(n9840), .B1(n9841), .B2(n7433), .ZN(n7266)
         );
  INV_X1 U8974 ( .A(n7256), .ZN(n7263) );
  AND2_X1 U8975 ( .A1(n7258), .A2(n7257), .ZN(n7259) );
  NAND2_X1 U8976 ( .A1(n7200), .A2(n7259), .ZN(n7261) );
  INV_X1 U8977 ( .A(n8352), .ZN(n7260) );
  INV_X1 U8978 ( .A(n9844), .ZN(n8692) );
  AOI21_X1 U8979 ( .B1(n7261), .B2(n7260), .A(n8692), .ZN(n7262) );
  OAI21_X1 U8980 ( .B1(n7264), .B2(n7263), .A(n7262), .ZN(n7265) );
  OAI211_X1 U8981 ( .C1(n9869), .C2(n9832), .A(n7266), .B(n7265), .ZN(n9871)
         );
  NAND2_X1 U8982 ( .A1(n9871), .A2(n8752), .ZN(n7273) );
  INV_X1 U8983 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7269) );
  INV_X1 U8984 ( .A(n7267), .ZN(n7268) );
  OAI22_X1 U8985 ( .A1(n8752), .A2(n7269), .B1(n7268), .B2(n9834), .ZN(n7270)
         );
  AOI21_X1 U8986 ( .B1(n8756), .B2(n7271), .A(n7270), .ZN(n7272) );
  OAI211_X1 U8987 ( .C1(n9869), .C2(n7697), .A(n7273), .B(n7272), .ZN(P2_U3228) );
  NOR2_X1 U8988 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7858), .ZN(n7279) );
  INV_X1 U8989 ( .A(n7274), .ZN(n7275) );
  AOI211_X1 U8990 ( .C1(n7277), .C2(n7276), .A(n7275), .B(n9486), .ZN(n7278)
         );
  AOI211_X1 U8991 ( .C1(n9490), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7279), .B(
        n7278), .ZN(n7285) );
  AOI21_X1 U8992 ( .B1(n7286), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7280), .ZN(
        n7281) );
  OAI21_X1 U8993 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7286), .A(n7281), .ZN(
        n7282) );
  NAND3_X1 U8994 ( .A1(n9492), .A2(n7283), .A3(n7282), .ZN(n7284) );
  OAI211_X1 U8995 ( .C1(n9498), .C2(n7286), .A(n7285), .B(n7284), .ZN(P1_U3254) );
  INV_X1 U8996 ( .A(n7287), .ZN(n7290) );
  INV_X1 U8997 ( .A(n9083), .ZN(n9098) );
  OAI222_X1 U8998 ( .A1(n8108), .A2(n7288), .B1(n9452), .B2(n7290), .C1(
        P1_U3086), .C2(n9098), .ZN(P1_U3338) );
  OAI222_X1 U8999 ( .A1(n7291), .A2(P2_U3151), .B1(n8901), .B2(n7290), .C1(
        n7289), .C2(n8899), .ZN(P2_U3278) );
  XNOR2_X1 U9000 ( .A(n7433), .B(n7304), .ZN(n8351) );
  XNOR2_X1 U9001 ( .A(n7292), .B(n8351), .ZN(n7293) );
  OAI222_X1 U9002 ( .A1(n8747), .A2(n7331), .B1(n8745), .B2(n7422), .C1(n8692), 
        .C2(n7293), .ZN(n7301) );
  INV_X1 U9003 ( .A(n7301), .ZN(n7298) );
  XOR2_X1 U9004 ( .A(n8351), .B(n7294), .Z(n7302) );
  AOI22_X1 U9005 ( .A1(n8586), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n8755), .B2(
        n7340), .ZN(n7295) );
  OAI21_X1 U9006 ( .B1(n7304), .B2(n8581), .A(n7295), .ZN(n7296) );
  AOI21_X1 U9007 ( .B1(n7302), .B2(n8759), .A(n7296), .ZN(n7297) );
  OAI21_X1 U9008 ( .B1(n7298), .B2(n8586), .A(n7297), .ZN(P2_U3227) );
  INV_X1 U9009 ( .A(n7299), .ZN(n7348) );
  AOI22_X1 U9010 ( .A1(n9111), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9447), .ZN(n7300) );
  OAI21_X1 U9011 ( .B1(n7348), .B2(n9452), .A(n7300), .ZN(P1_U3337) );
  AOI21_X1 U9012 ( .B1(n9865), .B2(n7302), .A(n7301), .ZN(n7309) );
  INV_X1 U9013 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7303) );
  OAI22_X1 U9014 ( .A1(n7304), .A2(n8822), .B1(n9891), .B2(n7303), .ZN(n7305)
         );
  INV_X1 U9015 ( .A(n7305), .ZN(n7306) );
  OAI21_X1 U9016 ( .B1(n7309), .B2(n9893), .A(n7306), .ZN(P2_U3408) );
  AOI22_X1 U9017 ( .A1(n8808), .A2(n7341), .B1(n9902), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7308) );
  OAI21_X1 U9018 ( .B1(n7309), .B2(n9902), .A(n7308), .ZN(P2_U3465) );
  XNOR2_X1 U9019 ( .A(n7310), .B(n7316), .ZN(n9584) );
  NAND3_X1 U9020 ( .A1(n7313), .A2(n7312), .A3(n7311), .ZN(n7314) );
  AND2_X1 U9021 ( .A1(n9537), .A2(n9513), .ZN(n7315) );
  XNOR2_X1 U9022 ( .A(n7317), .B(n7316), .ZN(n7320) );
  INV_X1 U9023 ( .A(n7318), .ZN(n7319) );
  AOI21_X1 U9024 ( .B1(n7320), .B2(n9541), .A(n7319), .ZN(n9581) );
  MUX2_X1 U9025 ( .A(n9581), .B(n6765), .S(n9543), .Z(n7326) );
  AOI211_X1 U9026 ( .C1(n9580), .C2(n9529), .A(n9620), .B(n4318), .ZN(n9579)
         );
  OAI22_X1 U9027 ( .A1(n9545), .A2(n7323), .B1(n9294), .B2(n7322), .ZN(n7324)
         );
  AOI21_X1 U9028 ( .B1(n9579), .B2(n9554), .A(n7324), .ZN(n7325) );
  OAI211_X1 U9029 ( .C1(n9584), .C2(n9325), .A(n7326), .B(n7325), .ZN(P1_U3289) );
  INV_X1 U9030 ( .A(n7433), .ZN(n7327) );
  XNOR2_X1 U9031 ( .A(n8161), .B(n7341), .ZN(n7358) );
  XNOR2_X1 U9032 ( .A(n7327), .B(n7358), .ZN(n7338) );
  NAND2_X1 U9033 ( .A1(n7329), .A2(n7328), .ZN(n7333) );
  NAND2_X1 U9034 ( .A1(n7331), .A2(n7330), .ZN(n7332) );
  NAND2_X1 U9035 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  INV_X1 U9036 ( .A(n7334), .ZN(n7336) );
  INV_X1 U9037 ( .A(n7361), .ZN(n7337) );
  AOI211_X1 U9038 ( .C1(n7338), .C2(n7334), .A(n8503), .B(n7337), .ZN(n7347)
         );
  NAND2_X1 U9039 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9749) );
  INV_X1 U9040 ( .A(n9749), .ZN(n7339) );
  AOI21_X1 U9041 ( .B1(n8510), .B2(n8530), .A(n7339), .ZN(n7345) );
  NAND2_X1 U9042 ( .A1(n8514), .A2(n7340), .ZN(n7344) );
  NAND2_X1 U9043 ( .A1(n8501), .A2(n7341), .ZN(n7343) );
  OR2_X1 U9044 ( .A1(n8512), .A2(n7422), .ZN(n7342) );
  NAND4_X1 U9045 ( .A1(n7345), .A2(n7344), .A3(n7343), .A4(n7342), .ZN(n7346)
         );
  OR2_X1 U9046 ( .A1(n7347), .A2(n7346), .ZN(P2_U3179) );
  OAI222_X1 U9047 ( .A1(n8899), .A2(n7349), .B1(n8901), .B2(n7348), .C1(
        P2_U3151), .C2(n8558), .ZN(P2_U3277) );
  INV_X1 U9048 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7357) );
  NOR2_X1 U9049 ( .A1(n9272), .A2(n9620), .ZN(n9228) );
  OAI21_X1 U9050 ( .B1(n9228), .B2(n9296), .A(n9548), .ZN(n7356) );
  NOR2_X1 U9051 ( .A1(n7351), .A2(n7350), .ZN(n7354) );
  OAI21_X1 U9052 ( .B1(n9294), .B2(n6925), .A(n7352), .ZN(n7353) );
  OAI21_X1 U9053 ( .B1(n7354), .B2(n7353), .A(n9322), .ZN(n7355) );
  OAI211_X1 U9054 ( .C1(n9322), .C2(n7357), .A(n7356), .B(n7355), .ZN(P1_U3293) );
  INV_X1 U9055 ( .A(n7436), .ZN(n7369) );
  INV_X1 U9056 ( .A(n7358), .ZN(n7359) );
  NAND2_X1 U9057 ( .A1(n7359), .A2(n7433), .ZN(n7360) );
  XNOR2_X1 U9058 ( .A(n7437), .B(n8161), .ZN(n7410) );
  XNOR2_X1 U9059 ( .A(n7410), .B(n8529), .ZN(n7362) );
  OAI21_X1 U9060 ( .B1(n4390), .B2(n7362), .A(n7411), .ZN(n7363) );
  NAND2_X1 U9061 ( .A1(n7363), .A2(n8508), .ZN(n7368) );
  AOI21_X1 U9062 ( .B1(n8510), .B2(n7433), .A(n7364), .ZN(n7365) );
  OAI21_X1 U9063 ( .B1(n7760), .B2(n8512), .A(n7365), .ZN(n7366) );
  AOI21_X1 U9064 ( .B1(n7437), .B2(n8501), .A(n7366), .ZN(n7367) );
  OAI211_X1 U9065 ( .C1(n7369), .C2(n8466), .A(n7368), .B(n7367), .ZN(P2_U3153) );
  OAI21_X1 U9066 ( .B1(n7371), .B2(n7370), .A(n7529), .ZN(n7374) );
  NAND2_X1 U9067 ( .A1(n9039), .A2(n8982), .ZN(n7373) );
  NAND2_X1 U9068 ( .A1(n9037), .A2(n8983), .ZN(n7372) );
  NAND2_X1 U9069 ( .A1(n7373), .A2(n7372), .ZN(n7747) );
  AOI21_X1 U9070 ( .B1(n7374), .B2(n9541), .A(n7747), .ZN(n9615) );
  XNOR2_X1 U9071 ( .A(n7375), .B(n7376), .ZN(n9618) );
  NAND2_X1 U9072 ( .A1(n9618), .A2(n9531), .ZN(n7383) );
  INV_X1 U9073 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7378) );
  INV_X1 U9074 ( .A(n7377), .ZN(n7749) );
  OAI22_X1 U9075 ( .A1(n9322), .A2(n7378), .B1(n7749), .B2(n9294), .ZN(n7381)
         );
  INV_X1 U9076 ( .A(n7535), .ZN(n7379) );
  OAI211_X1 U9077 ( .C1(n9616), .C2(n7513), .A(n7379), .B(n9551), .ZN(n9614)
         );
  NOR2_X1 U9078 ( .A1(n9614), .A2(n9272), .ZN(n7380) );
  AOI211_X1 U9079 ( .C1(n9296), .C2(n7751), .A(n7381), .B(n7380), .ZN(n7382)
         );
  OAI211_X1 U9080 ( .C1(n9543), .C2(n9615), .A(n7383), .B(n7382), .ZN(P1_U3283) );
  NAND2_X1 U9081 ( .A1(n7667), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7384) );
  OAI21_X1 U9082 ( .B1(n7667), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7384), .ZN(
        n7388) );
  OAI21_X1 U9083 ( .B1(n7386), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7385), .ZN(
        n7387) );
  NOR2_X1 U9084 ( .A1(n7388), .A2(n7387), .ZN(n7666) );
  AOI211_X1 U9085 ( .C1(n7388), .C2(n7387), .A(n7666), .B(n9486), .ZN(n7398)
         );
  AND2_X1 U9086 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7389) );
  AOI21_X1 U9087 ( .B1(n9490), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7389), .ZN(
        n7396) );
  AOI21_X1 U9088 ( .B1(n7391), .B2(n9666), .A(n7390), .ZN(n7394) );
  NOR2_X1 U9089 ( .A1(n7667), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7392) );
  AOI21_X1 U9090 ( .B1(n7667), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7392), .ZN(
        n7393) );
  NAND2_X1 U9091 ( .A1(n7393), .A2(n7394), .ZN(n7672) );
  OAI211_X1 U9092 ( .C1(n7394), .C2(n7393), .A(n9492), .B(n7672), .ZN(n7395)
         );
  OAI211_X1 U9093 ( .C1(n9498), .C2(n7673), .A(n7396), .B(n7395), .ZN(n7397)
         );
  OR2_X1 U9094 ( .A1(n7398), .A2(n7397), .ZN(P1_U3256) );
  OAI21_X1 U9095 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n7408) );
  INV_X1 U9096 ( .A(n7495), .ZN(n9602) );
  NAND2_X1 U9097 ( .A1(n9041), .A2(n8982), .ZN(n7403) );
  NAND2_X1 U9098 ( .A1(n9039), .A2(n8983), .ZN(n7402) );
  NAND2_X1 U9099 ( .A1(n7403), .A2(n7402), .ZN(n7488) );
  AOI21_X1 U9100 ( .B1(n9001), .B2(n7488), .A(n7404), .ZN(n7406) );
  NAND2_X1 U9101 ( .A1(n9013), .A2(n7494), .ZN(n7405) );
  OAI211_X1 U9102 ( .C1(n9602), .C2(n9017), .A(n7406), .B(n7405), .ZN(n7407)
         );
  AOI21_X1 U9103 ( .B1(n7408), .B2(n9007), .A(n7407), .ZN(n7409) );
  INV_X1 U9104 ( .A(n7409), .ZN(P1_U3221) );
  XNOR2_X1 U9105 ( .A(n9883), .B(n8161), .ZN(n7761) );
  XNOR2_X1 U9106 ( .A(n7761), .B(n8528), .ZN(n7758) );
  XOR2_X1 U9107 ( .A(n7759), .B(n7758), .Z(n7417) );
  NAND2_X1 U9108 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9772) );
  INV_X1 U9109 ( .A(n9772), .ZN(n7412) );
  AOI21_X1 U9110 ( .B1(n8510), .B2(n8529), .A(n7412), .ZN(n7414) );
  NAND2_X1 U9111 ( .A1(n8514), .A2(n7423), .ZN(n7413) );
  OAI211_X1 U9112 ( .C1(n7820), .C2(n8512), .A(n7414), .B(n7413), .ZN(n7415)
         );
  AOI21_X1 U9113 ( .B1(n9883), .B2(n8501), .A(n7415), .ZN(n7416) );
  OAI21_X1 U9114 ( .B1(n7417), .B2(n8503), .A(n7416), .ZN(P2_U3161) );
  NAND2_X1 U9115 ( .A1(n8224), .A2(n8232), .ZN(n8350) );
  NAND2_X1 U9116 ( .A1(n7430), .A2(n7418), .ZN(n7419) );
  XOR2_X1 U9117 ( .A(n8350), .B(n7419), .Z(n9880) );
  XNOR2_X1 U9118 ( .A(n7420), .B(n8350), .ZN(n7421) );
  OAI222_X1 U9119 ( .A1(n8747), .A2(n7422), .B1(n8745), .B2(n7820), .C1(n7421), 
        .C2(n8692), .ZN(n9881) );
  NAND2_X1 U9120 ( .A1(n9881), .A2(n8752), .ZN(n7427) );
  INV_X1 U9121 ( .A(n7423), .ZN(n7424) );
  OAI22_X1 U9122 ( .A1(n8752), .A2(n9983), .B1(n7424), .B2(n9834), .ZN(n7425)
         );
  AOI21_X1 U9123 ( .B1(n8756), .B2(n9883), .A(n7425), .ZN(n7426) );
  OAI211_X1 U9124 ( .C1(n9880), .C2(n8741), .A(n7427), .B(n7426), .ZN(P2_U3225) );
  OR2_X1 U9125 ( .A1(n7428), .A2(n8348), .ZN(n7429) );
  NAND2_X1 U9126 ( .A1(n7430), .A2(n7429), .ZN(n9875) );
  XOR2_X1 U9127 ( .A(n7431), .B(n8348), .Z(n7432) );
  NAND2_X1 U9128 ( .A1(n7432), .A2(n9844), .ZN(n7435) );
  AOI22_X1 U9129 ( .A1(n9840), .A2(n7433), .B1(n8528), .B2(n9841), .ZN(n7434)
         );
  OAI211_X1 U9130 ( .C1(n9832), .C2(n9875), .A(n7435), .B(n7434), .ZN(n9877)
         );
  AOI22_X1 U9131 ( .A1(n8586), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8755), .B2(
        n7436), .ZN(n7439) );
  NAND2_X1 U9132 ( .A1(n8756), .A2(n7437), .ZN(n7438) );
  OAI211_X1 U9133 ( .C1(n9875), .C2(n7697), .A(n7439), .B(n7438), .ZN(n7440)
         );
  AOI21_X1 U9134 ( .B1(n9877), .B2(n8752), .A(n7440), .ZN(n7441) );
  INV_X1 U9135 ( .A(n7441), .ZN(P2_U3226) );
  XNOR2_X1 U9136 ( .A(n7442), .B(n7446), .ZN(n7444) );
  AOI21_X1 U9137 ( .B1(n7444), .B2(n9541), .A(n7443), .ZN(n9588) );
  XNOR2_X1 U9138 ( .A(n7445), .B(n7446), .ZN(n9591) );
  INV_X1 U9139 ( .A(n9515), .ZN(n7447) );
  OAI211_X1 U9140 ( .C1(n9589), .C2(n7448), .A(n7447), .B(n9551), .ZN(n9587)
         );
  AOI22_X1 U9141 ( .A1(n9268), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7449), .B2(
        n9542), .ZN(n7452) );
  NAND2_X1 U9142 ( .A1(n9296), .A2(n7450), .ZN(n7451) );
  OAI211_X1 U9143 ( .C1(n9587), .C2(n9272), .A(n7452), .B(n7451), .ZN(n7453)
         );
  AOI21_X1 U9144 ( .B1(n9591), .B2(n9531), .A(n7453), .ZN(n7454) );
  OAI21_X1 U9145 ( .B1(n9588), .B2(n9268), .A(n7454), .ZN(P1_U3287) );
  AOI22_X1 U9146 ( .A1(n9268), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7455), .B2(
        n9542), .ZN(n7458) );
  NAND2_X1 U9147 ( .A1(n9296), .A2(n7456), .ZN(n7457) );
  OAI211_X1 U9148 ( .C1(n7459), .C2(n9272), .A(n7458), .B(n7457), .ZN(n7460)
         );
  AOI21_X1 U9149 ( .B1(n7461), .B2(n9531), .A(n7460), .ZN(n7462) );
  OAI21_X1 U9150 ( .B1(n7463), .B2(n9268), .A(n7462), .ZN(P1_U3288) );
  XNOR2_X1 U9151 ( .A(n7464), .B(n7465), .ZN(n9629) );
  INV_X1 U9152 ( .A(n9629), .ZN(n7475) );
  XNOR2_X1 U9153 ( .A(n7467), .B(n7466), .ZN(n7468) );
  AOI22_X1 U9154 ( .A1(n8982), .A2(n9037), .B1(n9036), .B2(n8983), .ZN(n7661)
         );
  OAI21_X1 U9155 ( .B1(n7468), .B2(n9506), .A(n7661), .ZN(n9627) );
  NAND2_X1 U9156 ( .A1(n7534), .A2(n7663), .ZN(n7469) );
  NAND2_X1 U9157 ( .A1(n7469), .A2(n9551), .ZN(n7470) );
  OR2_X1 U9158 ( .A1(n7470), .A2(n4388), .ZN(n9625) );
  AOI22_X1 U9159 ( .A1(n9268), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7658), .B2(
        n9542), .ZN(n7472) );
  NAND2_X1 U9160 ( .A1(n7663), .A2(n9296), .ZN(n7471) );
  OAI211_X1 U9161 ( .C1(n9625), .C2(n9272), .A(n7472), .B(n7471), .ZN(n7473)
         );
  AOI21_X1 U9162 ( .B1(n9627), .B2(n9322), .A(n7473), .ZN(n7474) );
  OAI21_X1 U9163 ( .B1(n7475), .B2(n9325), .A(n7474), .ZN(P1_U3281) );
  NAND2_X1 U9164 ( .A1(n7399), .A2(n7476), .ZN(n7479) );
  NAND2_X1 U9165 ( .A1(n7743), .A2(n7477), .ZN(n7478) );
  XNOR2_X1 U9166 ( .A(n7479), .B(n7478), .ZN(n7484) );
  NAND2_X1 U9167 ( .A1(n9038), .A2(n8983), .ZN(n7515) );
  NAND2_X1 U9168 ( .A1(n9040), .A2(n8982), .ZN(n7507) );
  AOI21_X1 U9169 ( .B1(n7515), .B2(n7507), .A(n9011), .ZN(n7480) );
  AOI211_X1 U9170 ( .C1(n9013), .C2(n7517), .A(n7481), .B(n7480), .ZN(n7483)
         );
  NAND2_X1 U9171 ( .A1(n9608), .A2(n8968), .ZN(n7482) );
  OAI211_X1 U9172 ( .C1(n7484), .C2(n8988), .A(n7483), .B(n7482), .ZN(P1_U3231) );
  INV_X1 U9173 ( .A(n7485), .ZN(n7486) );
  OR2_X1 U9174 ( .A1(n9503), .A2(n7486), .ZN(n7504) );
  XNOR2_X1 U9175 ( .A(n7504), .B(n4752), .ZN(n7487) );
  NAND2_X1 U9176 ( .A1(n7487), .A2(n9541), .ZN(n7490) );
  INV_X1 U9177 ( .A(n7488), .ZN(n7489) );
  NAND2_X1 U9178 ( .A1(n7490), .A2(n7489), .ZN(n9605) );
  INV_X1 U9179 ( .A(n9605), .ZN(n7500) );
  XNOR2_X1 U9180 ( .A(n7491), .B(n7492), .ZN(n9600) );
  AOI21_X1 U9181 ( .B1(n9514), .B2(n7495), .A(n9620), .ZN(n7493) );
  NAND2_X1 U9182 ( .A1(n7493), .A2(n7511), .ZN(n9601) );
  AOI22_X1 U9183 ( .A1(n9543), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7494), .B2(
        n9542), .ZN(n7497) );
  NAND2_X1 U9184 ( .A1(n9296), .A2(n7495), .ZN(n7496) );
  OAI211_X1 U9185 ( .C1(n9601), .C2(n9272), .A(n7497), .B(n7496), .ZN(n7498)
         );
  AOI21_X1 U9186 ( .B1(n9600), .B2(n9531), .A(n7498), .ZN(n7499) );
  OAI21_X1 U9187 ( .B1(n7500), .B2(n9268), .A(n7499), .ZN(P1_U3285) );
  INV_X1 U9188 ( .A(n7501), .ZN(n7503) );
  OAI21_X1 U9189 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7505) );
  XNOR2_X1 U9190 ( .A(n7505), .B(n7510), .ZN(n7506) );
  NAND2_X1 U9191 ( .A1(n7506), .A2(n9541), .ZN(n7508) );
  NAND2_X1 U9192 ( .A1(n7508), .A2(n7507), .ZN(n9612) );
  INV_X1 U9193 ( .A(n9612), .ZN(n7523) );
  XNOR2_X1 U9194 ( .A(n7509), .B(n7510), .ZN(n9607) );
  INV_X1 U9195 ( .A(n9608), .ZN(n7520) );
  NAND2_X1 U9196 ( .A1(n7511), .A2(n9608), .ZN(n7512) );
  NAND2_X1 U9197 ( .A1(n7512), .A2(n9551), .ZN(n7514) );
  OR2_X1 U9198 ( .A1(n7514), .A2(n7513), .ZN(n7516) );
  NAND2_X1 U9199 ( .A1(n7516), .A2(n7515), .ZN(n9609) );
  NAND2_X1 U9200 ( .A1(n9609), .A2(n9554), .ZN(n7519) );
  AOI22_X1 U9201 ( .A1(n9543), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7517), .B2(
        n9542), .ZN(n7518) );
  OAI211_X1 U9202 ( .C1(n7520), .C2(n9545), .A(n7519), .B(n7518), .ZN(n7521)
         );
  AOI21_X1 U9203 ( .B1(n9607), .B2(n9531), .A(n7521), .ZN(n7522) );
  OAI21_X1 U9204 ( .B1(n7523), .B2(n9543), .A(n7522), .ZN(P1_U3284) );
  XNOR2_X1 U9205 ( .A(n7524), .B(n7525), .ZN(n9624) );
  INV_X1 U9206 ( .A(n9624), .ZN(n7542) );
  NAND2_X1 U9207 ( .A1(n7526), .A2(n9541), .ZN(n7533) );
  AOI21_X1 U9208 ( .B1(n7529), .B2(n7528), .A(n7527), .ZN(n7532) );
  NAND2_X1 U9209 ( .A1(n9038), .A2(n8982), .ZN(n7531) );
  NAND2_X1 U9210 ( .A1(n7545), .A2(n8983), .ZN(n7530) );
  AND2_X1 U9211 ( .A1(n7531), .A2(n7530), .ZN(n7859) );
  OAI21_X1 U9212 ( .B1(n7533), .B2(n7532), .A(n7859), .ZN(n9622) );
  OAI21_X1 U9213 ( .B1(n7535), .B2(n4596), .A(n7534), .ZN(n9621) );
  INV_X1 U9214 ( .A(n9228), .ZN(n7539) );
  AOI22_X1 U9215 ( .A1(n9543), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7862), .B2(
        n9542), .ZN(n7538) );
  NAND2_X1 U9216 ( .A1(n7536), .A2(n9296), .ZN(n7537) );
  OAI211_X1 U9217 ( .C1(n9621), .C2(n7539), .A(n7538), .B(n7537), .ZN(n7540)
         );
  AOI21_X1 U9218 ( .B1(n9622), .B2(n9322), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9219 ( .B1(n7542), .B2(n9325), .A(n7541), .ZN(P1_U3282) );
  NAND2_X1 U9220 ( .A1(n7543), .A2(n7551), .ZN(n7544) );
  NAND2_X1 U9221 ( .A1(n7642), .A2(n7544), .ZN(n7549) );
  NAND2_X1 U9222 ( .A1(n7545), .A2(n8982), .ZN(n7547) );
  NAND2_X1 U9223 ( .A1(n9035), .A2(n8983), .ZN(n7546) );
  AND2_X1 U9224 ( .A1(n7547), .A2(n7546), .ZN(n7708) );
  INV_X1 U9225 ( .A(n7708), .ZN(n7548) );
  AOI21_X1 U9226 ( .B1(n7549), .B2(n9541), .A(n7548), .ZN(n9631) );
  XNOR2_X1 U9227 ( .A(n7550), .B(n7551), .ZN(n9636) );
  NAND2_X1 U9228 ( .A1(n9636), .A2(n9531), .ZN(n7556) );
  OAI211_X1 U9229 ( .C1(n9633), .C2(n4388), .A(n9551), .B(n7651), .ZN(n9630)
         );
  INV_X1 U9230 ( .A(n9630), .ZN(n7554) );
  AOI22_X1 U9231 ( .A1(n9543), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7711), .B2(
        n9542), .ZN(n7552) );
  OAI21_X1 U9232 ( .B1(n9633), .B2(n9545), .A(n7552), .ZN(n7553) );
  AOI21_X1 U9233 ( .B1(n7554), .B2(n9554), .A(n7553), .ZN(n7555) );
  OAI211_X1 U9234 ( .C1(n9543), .C2(n9631), .A(n7556), .B(n7555), .ZN(P1_U3280) );
  INV_X1 U9235 ( .A(n7557), .ZN(n7560) );
  OAI222_X1 U9236 ( .A1(P2_U3151), .A2(n7559), .B1(n8901), .B2(n7560), .C1(
        n7558), .C2(n8899), .ZN(P2_U3276) );
  OAI222_X1 U9237 ( .A1(n8108), .A2(n7561), .B1(n9452), .B2(n7560), .C1(
        P1_U3086), .C2(n5833), .ZN(P1_U3336) );
  XNOR2_X1 U9238 ( .A(n7562), .B(n7566), .ZN(n7564) );
  OAI21_X1 U9239 ( .B1(n7564), .B2(n9506), .A(n7563), .ZN(n9568) );
  INV_X1 U9240 ( .A(n9568), .ZN(n7575) );
  XNOR2_X1 U9241 ( .A(n7566), .B(n7565), .ZN(n9570) );
  INV_X1 U9242 ( .A(n9552), .ZN(n7569) );
  INV_X1 U9243 ( .A(n7567), .ZN(n7568) );
  OAI211_X1 U9244 ( .C1(n5151), .C2(n7569), .A(n7568), .B(n9551), .ZN(n9567)
         );
  INV_X1 U9245 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7570) );
  OAI22_X1 U9246 ( .A1(n9322), .A2(n9999), .B1(n7570), .B2(n9294), .ZN(n7571)
         );
  AOI21_X1 U9247 ( .B1(n9296), .B2(n5611), .A(n7571), .ZN(n7572) );
  OAI21_X1 U9248 ( .B1(n9272), .B2(n9567), .A(n7572), .ZN(n7573) );
  AOI21_X1 U9249 ( .B1(n9531), .B2(n9570), .A(n7573), .ZN(n7574) );
  OAI21_X1 U9250 ( .B1(n9543), .B2(n7575), .A(n7574), .ZN(P1_U3291) );
  AOI21_X1 U9251 ( .B1(n7578), .B2(n7577), .A(n7576), .ZN(n7591) );
  OAI21_X1 U9252 ( .B1(n7580), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7579), .ZN(
        n7589) );
  OAI21_X1 U9253 ( .B1(n7582), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7581), .ZN(
        n7583) );
  NAND2_X1 U9254 ( .A1(n7583), .A2(n9758), .ZN(n7586) );
  INV_X1 U9255 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7584) );
  NOR2_X1 U9256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7584), .ZN(n7754) );
  AOI21_X1 U9257 ( .B1(n9808), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7754), .ZN(
        n7585) );
  OAI211_X1 U9258 ( .C1(n9807), .C2(n7587), .A(n7586), .B(n7585), .ZN(n7588)
         );
  AOI21_X1 U9259 ( .B1(n9768), .B2(n7589), .A(n7588), .ZN(n7590) );
  OAI21_X1 U9260 ( .B1(n7591), .B2(n9763), .A(n7590), .ZN(P2_U3191) );
  NOR2_X1 U9261 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7636) );
  NOR2_X1 U9262 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7633) );
  NOR2_X1 U9263 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7631) );
  NOR2_X1 U9264 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7628) );
  NOR2_X1 U9265 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7626) );
  NOR2_X1 U9266 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7623) );
  NOR2_X1 U9267 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7621) );
  NOR2_X1 U9268 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7618) );
  NOR2_X1 U9269 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7615) );
  NOR2_X1 U9270 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7611) );
  NOR2_X1 U9271 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7608) );
  NOR2_X1 U9272 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7604) );
  NOR2_X1 U9273 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7602) );
  NOR2_X1 U9274 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7600) );
  NAND2_X1 U9275 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7598) );
  XOR2_X1 U9276 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10099) );
  NAND2_X1 U9277 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7596) );
  AOI21_X1 U9278 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9906) );
  INV_X1 U9279 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9280 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7592) );
  NOR2_X1 U9281 ( .A1(n7593), .A2(n7592), .ZN(n9905) );
  NOR2_X1 U9282 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9905), .ZN(n7594) );
  NOR2_X1 U9283 ( .A1(n9906), .A2(n7594), .ZN(n10097) );
  XOR2_X1 U9284 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10096) );
  NAND2_X1 U9285 ( .A1(n10097), .A2(n10096), .ZN(n7595) );
  NAND2_X1 U9286 ( .A1(n7596), .A2(n7595), .ZN(n10098) );
  NAND2_X1 U9287 ( .A1(n10099), .A2(n10098), .ZN(n7597) );
  NAND2_X1 U9288 ( .A1(n7598), .A2(n7597), .ZN(n10101) );
  XNOR2_X1 U9289 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10100) );
  NOR2_X1 U9290 ( .A1(n10101), .A2(n10100), .ZN(n7599) );
  NOR2_X1 U9291 ( .A1(n7600), .A2(n7599), .ZN(n10089) );
  XNOR2_X1 U9292 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10088) );
  NOR2_X1 U9293 ( .A1(n10089), .A2(n10088), .ZN(n7601) );
  NOR2_X1 U9294 ( .A1(n7602), .A2(n7601), .ZN(n10087) );
  XNOR2_X1 U9295 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10086) );
  NOR2_X1 U9296 ( .A1(n10087), .A2(n10086), .ZN(n7603) );
  NOR2_X1 U9297 ( .A1(n7604), .A2(n7603), .ZN(n10093) );
  INV_X1 U9298 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7606) );
  INV_X1 U9299 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7605) );
  AOI22_X1 U9300 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n7606), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n7605), .ZN(n10092) );
  NOR2_X1 U9301 ( .A1(n10093), .A2(n10092), .ZN(n7607) );
  NOR2_X1 U9302 ( .A1(n7608), .A2(n7607), .ZN(n10095) );
  INV_X1 U9303 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7609) );
  INV_X1 U9304 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U9305 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7609), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10024), .ZN(n10094) );
  NOR2_X1 U9306 ( .A1(n10095), .A2(n10094), .ZN(n7610) );
  NOR2_X1 U9307 ( .A1(n7611), .A2(n7610), .ZN(n10091) );
  INV_X1 U9308 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7613) );
  INV_X1 U9309 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7612) );
  AOI22_X1 U9310 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7613), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7612), .ZN(n10090) );
  NOR2_X1 U9311 ( .A1(n10091), .A2(n10090), .ZN(n7614) );
  NOR2_X1 U9312 ( .A1(n7615), .A2(n7614), .ZN(n9926) );
  INV_X1 U9313 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7616) );
  INV_X1 U9314 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U9315 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7616), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10007), .ZN(n9925) );
  NOR2_X1 U9316 ( .A1(n9926), .A2(n9925), .ZN(n7617) );
  NOR2_X1 U9317 ( .A1(n7618), .A2(n7617), .ZN(n9924) );
  INV_X1 U9318 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7619) );
  INV_X1 U9319 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8072) );
  AOI22_X1 U9320 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7619), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n8072), .ZN(n9923) );
  NOR2_X1 U9321 ( .A1(n9924), .A2(n9923), .ZN(n7620) );
  NOR2_X1 U9322 ( .A1(n7621), .A2(n7620), .ZN(n9922) );
  INV_X1 U9323 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8021) );
  AOI22_X1 U9324 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7249), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n8021), .ZN(n9921) );
  NOR2_X1 U9325 ( .A1(n9922), .A2(n9921), .ZN(n7622) );
  NOR2_X1 U9326 ( .A1(n7623), .A2(n7622), .ZN(n9920) );
  INV_X1 U9327 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7624) );
  INV_X1 U9328 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U9329 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7624), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9971), .ZN(n9919) );
  NOR2_X1 U9330 ( .A1(n9920), .A2(n9919), .ZN(n7625) );
  NOR2_X1 U9331 ( .A1(n7626), .A2(n7625), .ZN(n9918) );
  XNOR2_X1 U9332 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9917) );
  NOR2_X1 U9333 ( .A1(n9918), .A2(n9917), .ZN(n7627) );
  NOR2_X1 U9334 ( .A1(n7628), .A2(n7627), .ZN(n9916) );
  INV_X1 U9335 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7629) );
  INV_X1 U9336 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8541) );
  AOI22_X1 U9337 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7629), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8541), .ZN(n9915) );
  NOR2_X1 U9338 ( .A1(n9916), .A2(n9915), .ZN(n7630) );
  NOR2_X1 U9339 ( .A1(n7631), .A2(n7630), .ZN(n9914) );
  XNOR2_X1 U9340 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9913) );
  NOR2_X1 U9341 ( .A1(n9914), .A2(n9913), .ZN(n7632) );
  NOR2_X1 U9342 ( .A1(n7633), .A2(n7632), .ZN(n9912) );
  INV_X1 U9343 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7634) );
  INV_X1 U9344 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U9345 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7634), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9992), .ZN(n9911) );
  NOR2_X1 U9346 ( .A1(n9912), .A2(n9911), .ZN(n7635) );
  NOR2_X1 U9347 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  NOR2_X1 U9348 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7637), .ZN(n9908) );
  AND2_X1 U9349 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7637), .ZN(n9909) );
  NOR2_X1 U9350 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9909), .ZN(n7638) );
  NOR2_X1 U9351 ( .A1(n9908), .A2(n7638), .ZN(n7640) );
  XNOR2_X1 U9352 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7639) );
  XNOR2_X1 U9353 ( .A(n7640), .B(n7639), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9354 ( .A(n7641), .B(n7643), .ZN(n9643) );
  INV_X1 U9355 ( .A(n7642), .ZN(n7645) );
  OAI21_X1 U9356 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7646) );
  NAND3_X1 U9357 ( .A1(n7646), .A2(n7829), .A3(n9541), .ZN(n7649) );
  NAND2_X1 U9358 ( .A1(n9036), .A2(n8982), .ZN(n7648) );
  NAND2_X1 U9359 ( .A1(n9034), .A2(n8983), .ZN(n7647) );
  AND2_X1 U9360 ( .A1(n7648), .A2(n7647), .ZN(n7950) );
  NAND2_X1 U9361 ( .A1(n7649), .A2(n7950), .ZN(n9638) );
  AOI211_X1 U9362 ( .C1(n9640), .C2(n7651), .A(n9620), .B(n7650), .ZN(n9639)
         );
  NAND2_X1 U9363 ( .A1(n9639), .A2(n9554), .ZN(n7653) );
  AOI22_X1 U9364 ( .A1(n9543), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7952), .B2(
        n9542), .ZN(n7652) );
  OAI211_X1 U9365 ( .C1(n4532), .C2(n9545), .A(n7653), .B(n7652), .ZN(n7654)
         );
  AOI21_X1 U9366 ( .B1(n9322), .B2(n9638), .A(n7654), .ZN(n7655) );
  OAI21_X1 U9367 ( .B1(n9325), .B2(n9643), .A(n7655), .ZN(P1_U3279) );
  XOR2_X1 U9368 ( .A(n7656), .B(n7657), .Z(n7665) );
  NAND2_X1 U9369 ( .A1(n9013), .A2(n7658), .ZN(n7659) );
  OAI211_X1 U9370 ( .C1(n9011), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7662)
         );
  AOI21_X1 U9371 ( .B1(n7663), .B2(n8968), .A(n7662), .ZN(n7664) );
  OAI21_X1 U9372 ( .B1(n7665), .B2(n8988), .A(n7664), .ZN(P1_U3224) );
  INV_X1 U9373 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7668) );
  AOI22_X1 U9374 ( .A1(n7884), .A2(n7668), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7889), .ZN(n7669) );
  AOI211_X1 U9375 ( .C1(n7670), .C2(n7669), .A(n7883), .B(n9486), .ZN(n7680)
         );
  AND2_X1 U9376 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7671) );
  AOI21_X1 U9377 ( .B1(n9490), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7671), .ZN(
        n7678) );
  INV_X1 U9378 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9668) );
  OAI21_X1 U9379 ( .B1(n7673), .B2(n9668), .A(n7672), .ZN(n7676) );
  INV_X1 U9380 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7674) );
  MUX2_X1 U9381 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7674), .S(n7884), .Z(n7675)
         );
  NAND2_X1 U9382 ( .A1(n7675), .A2(n7676), .ZN(n7888) );
  OAI211_X1 U9383 ( .C1(n7676), .C2(n7675), .A(n9492), .B(n7888), .ZN(n7677)
         );
  OAI211_X1 U9384 ( .C1(n9498), .C2(n7889), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OR2_X1 U9385 ( .A1(n7680), .A2(n7679), .ZN(P1_U3257) );
  INV_X1 U9386 ( .A(n7681), .ZN(n7683) );
  OAI222_X1 U9387 ( .A1(P2_U3151), .A2(n7682), .B1(n8899), .B2(n6511), .C1(
        n7683), .C2(n8906), .ZN(P2_U3275) );
  OAI222_X1 U9388 ( .A1(n8108), .A2(n7685), .B1(P1_U3086), .B2(n7684), .C1(
        n9452), .C2(n7683), .ZN(P1_U3335) );
  NAND2_X1 U9389 ( .A1(n7687), .A2(n8355), .ZN(n7688) );
  NAND2_X1 U9390 ( .A1(n7686), .A2(n7688), .ZN(n9886) );
  XNOR2_X1 U9391 ( .A(n7689), .B(n8355), .ZN(n7690) );
  NAND2_X1 U9392 ( .A1(n7690), .A2(n9844), .ZN(n7692) );
  AOI22_X1 U9393 ( .A1(n9840), .A2(n8528), .B1(n8526), .B2(n9841), .ZN(n7691)
         );
  OAI211_X1 U9394 ( .C1(n9832), .C2(n9886), .A(n7692), .B(n7691), .ZN(n9887)
         );
  NAND2_X1 U9395 ( .A1(n9887), .A2(n8752), .ZN(n7696) );
  INV_X1 U9396 ( .A(n7755), .ZN(n7693) );
  OAI22_X1 U9397 ( .A1(n8752), .A2(n4639), .B1(n7693), .B2(n9834), .ZN(n7694)
         );
  AOI21_X1 U9398 ( .B1(n8756), .B2(n9889), .A(n7694), .ZN(n7695) );
  OAI211_X1 U9399 ( .C1(n9886), .C2(n7697), .A(n7696), .B(n7695), .ZN(P2_U3224) );
  NAND2_X1 U9400 ( .A1(n8206), .A2(n8229), .ZN(n8356) );
  XNOR2_X1 U9401 ( .A(n7698), .B(n8356), .ZN(n7699) );
  AOI222_X1 U9402 ( .A1(n9844), .A2(n7699), .B1(n8525), .B2(n9841), .C1(n8527), 
        .C2(n9840), .ZN(n7719) );
  NAND2_X1 U9403 ( .A1(n7686), .A2(n8225), .ZN(n7700) );
  XNOR2_X1 U9404 ( .A(n7700), .B(n8356), .ZN(n7716) );
  NAND2_X1 U9405 ( .A1(n8207), .A2(n8756), .ZN(n7702) );
  AOI22_X1 U9406 ( .A1(n8586), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8755), .B2(
        n7825), .ZN(n7701) );
  NAND2_X1 U9407 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  AOI21_X1 U9408 ( .B1(n7716), .B2(n8759), .A(n7703), .ZN(n7704) );
  OAI21_X1 U9409 ( .B1(n7719), .B2(n8586), .A(n7704), .ZN(P2_U3223) );
  XOR2_X1 U9410 ( .A(n7705), .B(n7706), .Z(n7713) );
  OAI22_X1 U9411 ( .A1(n9011), .A2(n7708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7707), .ZN(n7710) );
  NOR2_X1 U9412 ( .A1(n9633), .A2(n9017), .ZN(n7709) );
  AOI211_X1 U9413 ( .C1(n9013), .C2(n7711), .A(n7710), .B(n7709), .ZN(n7712)
         );
  OAI21_X1 U9414 ( .B1(n7713), .B2(n8988), .A(n7712), .ZN(P1_U3234) );
  AOI22_X1 U9415 ( .A1(n8207), .A2(n8808), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n9902), .ZN(n7715) );
  NAND2_X1 U9416 ( .A1(n7716), .A2(n8809), .ZN(n7714) );
  OAI211_X1 U9417 ( .C1(n7719), .C2(n9902), .A(n7715), .B(n7714), .ZN(P2_U3469) );
  AOI22_X1 U9418 ( .A1(n8889), .A2(n8207), .B1(n9893), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n7718) );
  INV_X1 U9419 ( .A(n9865), .ZN(n9879) );
  NAND2_X1 U9420 ( .A1(n7716), .A2(n8890), .ZN(n7717) );
  OAI211_X1 U9421 ( .C1(n7719), .C2(n9893), .A(n7718), .B(n7717), .ZN(P2_U3420) );
  INV_X1 U9422 ( .A(n7720), .ZN(n7722) );
  OAI222_X1 U9423 ( .A1(n8328), .A2(P2_U3151), .B1(n8901), .B2(n7722), .C1(
        n10021), .C2(n8899), .ZN(P2_U3274) );
  OAI222_X1 U9424 ( .A1(P1_U3086), .A2(n7723), .B1(n9452), .B2(n7722), .C1(
        n7721), .C2(n9450), .ZN(P1_U3334) );
  AOI21_X1 U9425 ( .B1(n7726), .B2(n7725), .A(n7724), .ZN(n7742) );
  AOI21_X1 U9426 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7739) );
  AOI21_X1 U9427 ( .B1(n7732), .B2(n7731), .A(n7730), .ZN(n7733) );
  OR2_X1 U9428 ( .A1(n7733), .A2(n9826), .ZN(n7738) );
  OAI22_X1 U9429 ( .A1(n9807), .A2(n7734), .B1(n9737), .B2(n10007), .ZN(n7736)
         );
  NAND2_X1 U9430 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7821) );
  INV_X1 U9431 ( .A(n7821), .ZN(n7735) );
  NOR2_X1 U9432 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  OAI211_X1 U9433 ( .C1(n7739), .C2(n9817), .A(n7738), .B(n7737), .ZN(n7740)
         );
  INV_X1 U9434 ( .A(n7740), .ZN(n7741) );
  OAI21_X1 U9435 ( .B1(n7742), .B2(n9763), .A(n7741), .ZN(P2_U3192) );
  AND2_X1 U9436 ( .A1(n7744), .A2(n7743), .ZN(n7852) );
  XNOR2_X1 U9437 ( .A(n7852), .B(n7853), .ZN(n7746) );
  NOR2_X1 U9438 ( .A1(n7746), .A2(n7745), .ZN(n7851) );
  AOI21_X1 U9439 ( .B1(n7746), .B2(n7745), .A(n7851), .ZN(n7753) );
  AOI22_X1 U9440 ( .A1(n9001), .A2(n7747), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7748) );
  OAI21_X1 U9441 ( .B1(n7749), .B2(n8998), .A(n7748), .ZN(n7750) );
  AOI21_X1 U9442 ( .B1(n7751), .B2(n8968), .A(n7750), .ZN(n7752) );
  OAI21_X1 U9443 ( .B1(n7753), .B2(n8988), .A(n7752), .ZN(P1_U3217) );
  AOI21_X1 U9444 ( .B1(n8510), .B2(n8528), .A(n7754), .ZN(n7757) );
  NAND2_X1 U9445 ( .A1(n8514), .A2(n7755), .ZN(n7756) );
  OAI211_X1 U9446 ( .C1(n7789), .C2(n8512), .A(n7757), .B(n7756), .ZN(n7768)
         );
  XNOR2_X1 U9447 ( .A(n9889), .B(n8161), .ZN(n7785) );
  XNOR2_X1 U9448 ( .A(n7785), .B(n7820), .ZN(n7766) );
  NAND2_X1 U9449 ( .A1(n7759), .A2(n7758), .ZN(n7763) );
  NAND2_X1 U9450 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  NAND2_X1 U9451 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  INV_X1 U9452 ( .A(n7788), .ZN(n7765) );
  AOI211_X1 U9453 ( .C1(n7766), .C2(n7764), .A(n8503), .B(n7765), .ZN(n7767)
         );
  AOI211_X1 U9454 ( .C1(n9889), .C2(n8501), .A(n7768), .B(n7767), .ZN(n7769)
         );
  INV_X1 U9455 ( .A(n7769), .ZN(P2_U3171) );
  INV_X1 U9456 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7774) );
  OAI211_X1 U9457 ( .C1(n7771), .C2(n8357), .A(n7770), .B(n9844), .ZN(n7773)
         );
  AOI22_X1 U9458 ( .A1(n8524), .A2(n9841), .B1(n9840), .B2(n8526), .ZN(n7772)
         );
  AND2_X1 U9459 ( .A1(n7773), .A2(n7772), .ZN(n7781) );
  MUX2_X1 U9460 ( .A(n7774), .B(n7781), .S(n9891), .Z(n7777) );
  XOR2_X1 U9461 ( .A(n8357), .B(n7775), .Z(n7780) );
  AOI22_X1 U9462 ( .A1(n7780), .A2(n8890), .B1(n8889), .B2(n8211), .ZN(n7776)
         );
  NAND2_X1 U9463 ( .A1(n7777), .A2(n7776), .ZN(P2_U3423) );
  MUX2_X1 U9464 ( .A(n8070), .B(n7781), .S(n9904), .Z(n7779) );
  AOI22_X1 U9465 ( .A1(n7780), .A2(n8809), .B1(n8808), .B2(n8211), .ZN(n7778)
         );
  NAND2_X1 U9466 ( .A1(n7779), .A2(n7778), .ZN(P2_U3470) );
  INV_X1 U9467 ( .A(n7780), .ZN(n7784) );
  MUX2_X1 U9468 ( .A(n8067), .B(n7781), .S(n8752), .Z(n7783) );
  AOI22_X1 U9469 ( .A1(n8211), .A2(n8756), .B1(n8755), .B2(n7871), .ZN(n7782)
         );
  OAI211_X1 U9470 ( .C1(n7784), .C2(n8741), .A(n7783), .B(n7782), .ZN(P2_U3222) );
  INV_X1 U9471 ( .A(n7785), .ZN(n7786) );
  NAND2_X1 U9472 ( .A1(n7786), .A2(n8527), .ZN(n7787) );
  XNOR2_X1 U9473 ( .A(n8357), .B(n7795), .ZN(n7869) );
  XNOR2_X1 U9474 ( .A(n8207), .B(n7795), .ZN(n7866) );
  INV_X1 U9475 ( .A(n7866), .ZN(n7790) );
  OR2_X1 U9476 ( .A1(n8209), .A2(n8161), .ZN(n7793) );
  OAI21_X1 U9477 ( .B1(n8206), .B2(n7795), .A(n7793), .ZN(n7797) );
  NAND3_X1 U9478 ( .A1(n8207), .A2(n7795), .A3(n8526), .ZN(n7794) );
  OAI211_X1 U9479 ( .C1(n8209), .C2(n7795), .A(n8357), .B(n7794), .ZN(n7796)
         );
  OAI21_X1 U9480 ( .B1(n8357), .B2(n7797), .A(n7796), .ZN(n7798) );
  NAND2_X1 U9481 ( .A1(n7799), .A2(n7798), .ZN(n7801) );
  XNOR2_X1 U9482 ( .A(n7958), .B(n8161), .ZN(n7914) );
  XNOR2_X1 U9483 ( .A(n7914), .B(n8244), .ZN(n7800) );
  NAND2_X1 U9484 ( .A1(n7801), .A2(n7800), .ZN(n7916) );
  OAI211_X1 U9485 ( .C1(n7801), .C2(n7800), .A(n7916), .B(n8508), .ZN(n7805)
         );
  AND2_X1 U9486 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8019) );
  AOI21_X1 U9487 ( .B1(n8496), .B2(n8523), .A(n8019), .ZN(n7802) );
  OAI21_X1 U9488 ( .B1(n8209), .B2(n8499), .A(n7802), .ZN(n7803) );
  AOI21_X1 U9489 ( .B1(n7909), .B2(n8514), .A(n7803), .ZN(n7804) );
  OAI211_X1 U9490 ( .C1(n7958), .C2(n8517), .A(n7805), .B(n7804), .ZN(P2_U3164) );
  XNOR2_X1 U9491 ( .A(n7807), .B(n7806), .ZN(n7811) );
  OAI22_X1 U9492 ( .A1(n7809), .A2(n8995), .B1(n7808), .B2(n8993), .ZN(n8942)
         );
  INV_X1 U9493 ( .A(n8942), .ZN(n7810) );
  OAI21_X1 U9494 ( .B1(n7811), .B2(n9506), .A(n7810), .ZN(n9458) );
  INV_X1 U9495 ( .A(n9458), .ZN(n7819) );
  OAI22_X1 U9496 ( .A1(n9322), .A2(n7812), .B1(n8944), .B2(n9294), .ZN(n7814)
         );
  INV_X1 U9497 ( .A(n8946), .ZN(n9457) );
  OAI211_X1 U9498 ( .C1(n9457), .C2(n4365), .A(n9551), .B(n7932), .ZN(n9455)
         );
  NOR2_X1 U9499 ( .A1(n9455), .A2(n9272), .ZN(n7813) );
  AOI211_X1 U9500 ( .C1(n9296), .C2(n8946), .A(n7814), .B(n7813), .ZN(n7818)
         );
  NAND2_X1 U9501 ( .A1(n7816), .A2(n7815), .ZN(n9454) );
  NAND3_X1 U9502 ( .A1(n4319), .A2(n9454), .A3(n9531), .ZN(n7817) );
  OAI211_X1 U9503 ( .C1(n7819), .C2(n9543), .A(n7818), .B(n7817), .ZN(P1_U3277) );
  XNOR2_X1 U9504 ( .A(n7865), .B(n8526), .ZN(n7867) );
  XOR2_X1 U9505 ( .A(n7866), .B(n7867), .Z(n7827) );
  OR2_X1 U9506 ( .A1(n8499), .A2(n7820), .ZN(n7822) );
  OAI211_X1 U9507 ( .C1(n8209), .C2(n8512), .A(n7822), .B(n7821), .ZN(n7824)
         );
  INV_X1 U9508 ( .A(n8207), .ZN(n8215) );
  NOR2_X1 U9509 ( .A1(n8215), .A2(n8517), .ZN(n7823) );
  AOI211_X1 U9510 ( .C1(n7825), .C2(n8514), .A(n7824), .B(n7823), .ZN(n7826)
         );
  OAI21_X1 U9511 ( .B1(n7827), .B2(n8503), .A(n7826), .ZN(P2_U3157) );
  NAND2_X1 U9512 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  XNOR2_X1 U9513 ( .A(n7830), .B(n7833), .ZN(n7831) );
  AOI22_X1 U9514 ( .A1(n9033), .A2(n8983), .B1(n9035), .B2(n8982), .ZN(n9010)
         );
  OAI21_X1 U9515 ( .B1(n7831), .B2(n9506), .A(n9010), .ZN(n7841) );
  INV_X1 U9516 ( .A(n7841), .ZN(n7840) );
  XOR2_X1 U9517 ( .A(n7832), .B(n7833), .Z(n7843) );
  AOI211_X1 U9518 ( .C1(n7835), .C2(n7834), .A(n9620), .B(n4365), .ZN(n7842)
         );
  NAND2_X1 U9519 ( .A1(n7842), .A2(n9554), .ZN(n7837) );
  AOI22_X1 U9520 ( .A1(n9543), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9014), .B2(
        n9542), .ZN(n7836) );
  OAI211_X1 U9521 ( .C1(n9018), .C2(n9545), .A(n7837), .B(n7836), .ZN(n7838)
         );
  AOI21_X1 U9522 ( .B1(n7843), .B2(n9531), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9523 ( .B1(n9543), .B2(n7840), .A(n7839), .ZN(P1_U3278) );
  AOI211_X1 U9524 ( .C1(n7843), .C2(n9635), .A(n7842), .B(n7841), .ZN(n7850)
         );
  INV_X1 U9525 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7844) );
  OAI22_X1 U9526 ( .A1(n9018), .A2(n9395), .B1(n10083), .B2(n7844), .ZN(n7845)
         );
  INV_X1 U9527 ( .A(n7845), .ZN(n7846) );
  OAI21_X1 U9528 ( .B1(n7850), .B2(n9670), .A(n7846), .ZN(P1_U3537) );
  INV_X1 U9529 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7847) );
  OAI22_X1 U9530 ( .A1(n9018), .A2(n5626), .B1(n9650), .B2(n7847), .ZN(n7848)
         );
  INV_X1 U9531 ( .A(n7848), .ZN(n7849) );
  OAI21_X1 U9532 ( .B1(n7850), .B2(n9648), .A(n7849), .ZN(P1_U3498) );
  AOI21_X1 U9533 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(n7857) );
  XNOR2_X1 U9534 ( .A(n7855), .B(n7854), .ZN(n7856) );
  XNOR2_X1 U9535 ( .A(n7857), .B(n7856), .ZN(n7864) );
  OAI22_X1 U9536 ( .A1(n9011), .A2(n7859), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7858), .ZN(n7861) );
  NOR2_X1 U9537 ( .A1(n4596), .A2(n9017), .ZN(n7860) );
  AOI211_X1 U9538 ( .C1(n9013), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  OAI21_X1 U9539 ( .B1(n7864), .B2(n8988), .A(n7863), .ZN(P1_U3236) );
  OAI22_X1 U9540 ( .A1(n7867), .A2(n7866), .B1(n8526), .B2(n7865), .ZN(n7868)
         );
  XOR2_X1 U9541 ( .A(n7869), .B(n7868), .Z(n7876) );
  INV_X1 U9542 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7870) );
  NOR2_X1 U9543 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7870), .ZN(n8080) );
  AOI21_X1 U9544 ( .B1(n8510), .B2(n8526), .A(n8080), .ZN(n7873) );
  NAND2_X1 U9545 ( .A1(n8514), .A2(n7871), .ZN(n7872) );
  OAI211_X1 U9546 ( .C1(n8244), .C2(n8512), .A(n7873), .B(n7872), .ZN(n7874)
         );
  AOI21_X1 U9547 ( .B1(n8211), .B2(n8501), .A(n7874), .ZN(n7875) );
  OAI21_X1 U9548 ( .B1(n7876), .B2(n8503), .A(n7875), .ZN(P2_U3176) );
  INV_X1 U9549 ( .A(n7877), .ZN(n7881) );
  OAI222_X1 U9550 ( .A1(P2_U3151), .A2(n7879), .B1(n8901), .B2(n7881), .C1(
        n7878), .C2(n8899), .ZN(P2_U3273) );
  OAI222_X1 U9551 ( .A1(n8108), .A2(n7882), .B1(n9452), .B2(n7881), .C1(
        P1_U3086), .C2(n7880), .ZN(P1_U3333) );
  INV_X1 U9552 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7886) );
  NOR2_X1 U9553 ( .A1(n7886), .A2(n7885), .ZN(n9057) );
  AOI211_X1 U9554 ( .C1(n7886), .C2(n7885), .A(n9057), .B(n9486), .ZN(n7894)
         );
  AND2_X1 U9555 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7887) );
  AOI21_X1 U9556 ( .B1(n9490), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7887), .ZN(
        n7892) );
  OAI21_X1 U9557 ( .B1(n7674), .B2(n7889), .A(n7888), .ZN(n9048) );
  XNOR2_X1 U9558 ( .A(n9055), .B(n9048), .ZN(n7890) );
  NAND2_X1 U9559 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7890), .ZN(n9050) );
  OAI211_X1 U9560 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7890), .A(n9492), .B(
        n9050), .ZN(n7891) );
  OAI211_X1 U9561 ( .C1(n9498), .C2(n9055), .A(n7892), .B(n7891), .ZN(n7893)
         );
  OR2_X1 U9562 ( .A1(n7894), .A2(n7893), .ZN(P1_U3258) );
  NAND2_X1 U9563 ( .A1(n7900), .A2(n7895), .ZN(n7897) );
  OAI211_X1 U9564 ( .C1(n7898), .C2(n8108), .A(n7897), .B(n7896), .ZN(P1_U3332) );
  NAND2_X1 U9565 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  OAI211_X1 U9566 ( .C1(n7902), .C2(n8899), .A(n7901), .B(n8390), .ZN(P2_U3272) );
  XNOR2_X1 U9567 ( .A(n7903), .B(n8359), .ZN(n7904) );
  NAND2_X1 U9568 ( .A1(n7904), .A2(n9844), .ZN(n7907) );
  OAI22_X1 U9569 ( .A1(n7995), .A2(n8745), .B1(n8209), .B2(n8747), .ZN(n7905)
         );
  INV_X1 U9570 ( .A(n7905), .ZN(n7906) );
  NAND2_X1 U9571 ( .A1(n7907), .A2(n7906), .ZN(n7960) );
  OR2_X1 U9572 ( .A1(n7908), .A2(n8359), .ZN(n7956) );
  NAND3_X1 U9573 ( .A1(n7956), .A2(n8759), .A3(n7955), .ZN(n7911) );
  AOI22_X1 U9574 ( .A1(n8586), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8755), .B2(
        n7909), .ZN(n7910) );
  OAI211_X1 U9575 ( .C1(n7958), .C2(n8581), .A(n7911), .B(n7910), .ZN(n7912)
         );
  AOI21_X1 U9576 ( .B1(n7960), .B2(n8752), .A(n7912), .ZN(n7913) );
  INV_X1 U9577 ( .A(n7913), .ZN(P2_U3221) );
  XNOR2_X1 U9578 ( .A(n7921), .B(n8161), .ZN(n7981) );
  XNOR2_X1 U9579 ( .A(n7981), .B(n8523), .ZN(n7919) );
  NAND2_X1 U9580 ( .A1(n7914), .A2(n8524), .ZN(n7915) );
  INV_X1 U9581 ( .A(n7984), .ZN(n7917) );
  AOI21_X1 U9582 ( .B1(n7919), .B2(n7918), .A(n7917), .ZN(n7925) );
  NAND2_X1 U9583 ( .A1(n8510), .A2(n8524), .ZN(n7920) );
  NAND2_X1 U9584 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8052) );
  OAI211_X1 U9585 ( .C1(n8005), .C2(n8512), .A(n7920), .B(n8052), .ZN(n7923)
         );
  NOR2_X1 U9586 ( .A1(n7921), .A2(n8517), .ZN(n7922) );
  AOI211_X1 U9587 ( .C1(n7975), .C2(n8514), .A(n7923), .B(n7922), .ZN(n7924)
         );
  OAI21_X1 U9588 ( .B1(n7925), .B2(n8503), .A(n7924), .ZN(P2_U3174) );
  OAI211_X1 U9589 ( .C1(n7936), .C2(n7927), .A(n9541), .B(n7926), .ZN(n7931)
         );
  OR2_X1 U9590 ( .A1(n8918), .A2(n8995), .ZN(n7929) );
  NAND2_X1 U9591 ( .A1(n9033), .A2(n8982), .ZN(n7928) );
  NAND2_X1 U9592 ( .A1(n7929), .A2(n7928), .ZN(n8953) );
  INV_X1 U9593 ( .A(n8953), .ZN(n7930) );
  NAND2_X1 U9594 ( .A1(n7931), .A2(n7930), .ZN(n9392) );
  INV_X1 U9595 ( .A(n9392), .ZN(n7940) );
  AOI211_X1 U9596 ( .C1(n7933), .C2(n7932), .A(n9620), .B(n4369), .ZN(n9391)
         );
  NOR2_X1 U9597 ( .A1(n4542), .A2(n9545), .ZN(n7935) );
  INV_X1 U9598 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9088) );
  OAI22_X1 U9599 ( .A1(n9322), .A2(n9088), .B1(n8951), .B2(n9294), .ZN(n7934)
         );
  AOI211_X1 U9600 ( .C1(n9391), .C2(n9554), .A(n7935), .B(n7934), .ZN(n7939)
         );
  XNOR2_X1 U9601 ( .A(n7937), .B(n7936), .ZN(n9393) );
  NAND2_X1 U9602 ( .A1(n9393), .A2(n9531), .ZN(n7938) );
  OAI211_X1 U9603 ( .C1(n9543), .C2(n7940), .A(n7939), .B(n7938), .ZN(P1_U3276) );
  INV_X1 U9604 ( .A(n7941), .ZN(n7943) );
  NOR2_X1 U9605 ( .A1(n7943), .A2(n7942), .ZN(n7945) );
  OAI22_X1 U9606 ( .A1(n7947), .A2(n7946), .B1(n7945), .B2(n7944), .ZN(n7948)
         );
  NAND2_X1 U9607 ( .A1(n7948), .A2(n9007), .ZN(n7954) );
  OAI22_X1 U9608 ( .A1(n9011), .A2(n7950), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7949), .ZN(n7951) );
  AOI21_X1 U9609 ( .B1(n7952), .B2(n9013), .A(n7951), .ZN(n7953) );
  OAI211_X1 U9610 ( .C1(n4532), .C2(n9017), .A(n7954), .B(n7953), .ZN(P1_U3215) );
  NAND3_X1 U9611 ( .A1(n7956), .A2(n7955), .A3(n9865), .ZN(n7957) );
  OAI21_X1 U9612 ( .B1(n7958), .B2(n9873), .A(n7957), .ZN(n7959) );
  NOR2_X1 U9613 ( .A1(n7960), .A2(n7959), .ZN(n7963) );
  MUX2_X1 U9614 ( .A(n7961), .B(n7963), .S(n9904), .Z(n7962) );
  INV_X1 U9615 ( .A(n7962), .ZN(P2_U3471) );
  INV_X1 U9616 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7964) );
  MUX2_X1 U9617 ( .A(n7964), .B(n7963), .S(n9891), .Z(n7965) );
  INV_X1 U9618 ( .A(n7965), .ZN(P2_U3426) );
  XNOR2_X1 U9619 ( .A(n7966), .B(n8358), .ZN(n7978) );
  OAI21_X1 U9620 ( .B1(n4376), .B2(n6626), .A(n7967), .ZN(n7968) );
  AOI222_X1 U9621 ( .A1(n9844), .A2(n7968), .B1(n8522), .B2(n9841), .C1(n8524), 
        .C2(n9840), .ZN(n7974) );
  MUX2_X1 U9622 ( .A(n8055), .B(n7974), .S(n9904), .Z(n7970) );
  NAND2_X1 U9623 ( .A1(n8249), .A2(n8808), .ZN(n7969) );
  OAI211_X1 U9624 ( .C1(n8806), .C2(n7978), .A(n7970), .B(n7969), .ZN(P2_U3472) );
  INV_X1 U9625 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7971) );
  MUX2_X1 U9626 ( .A(n7971), .B(n7974), .S(n9891), .Z(n7973) );
  NAND2_X1 U9627 ( .A1(n8249), .A2(n8889), .ZN(n7972) );
  OAI211_X1 U9628 ( .C1(n7978), .C2(n8884), .A(n7973), .B(n7972), .ZN(P2_U3429) );
  MUX2_X1 U9629 ( .A(n8048), .B(n7974), .S(n8752), .Z(n7977) );
  AOI22_X1 U9630 ( .A1(n8249), .A2(n8756), .B1(n8755), .B2(n7975), .ZN(n7976)
         );
  OAI211_X1 U9631 ( .C1(n7978), .C2(n8741), .A(n7977), .B(n7976), .ZN(P2_U3220) );
  INV_X1 U9632 ( .A(n7979), .ZN(n8171) );
  OAI222_X1 U9633 ( .A1(n5106), .A2(P1_U3086), .B1(n9452), .B2(n8171), .C1(
        n7980), .C2(n9450), .ZN(P1_U3331) );
  INV_X1 U9634 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U9635 ( .A1(n7982), .A2(n7995), .ZN(n7983) );
  XNOR2_X1 U9636 ( .A(n8038), .B(n8161), .ZN(n8006) );
  XNOR2_X1 U9637 ( .A(n8006), .B(n8522), .ZN(n8007) );
  XOR2_X1 U9638 ( .A(n8008), .B(n8007), .Z(n7989) );
  AOI22_X1 U9639 ( .A1(n8496), .A2(n8521), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7986) );
  NAND2_X1 U9640 ( .A1(n8514), .A2(n8043), .ZN(n7985) );
  OAI211_X1 U9641 ( .C1(n7995), .C2(n8499), .A(n7986), .B(n7985), .ZN(n7987)
         );
  AOI21_X1 U9642 ( .B1(n8038), .B2(n8501), .A(n7987), .ZN(n7988) );
  OAI21_X1 U9643 ( .B1(n7989), .B2(n8503), .A(n7988), .ZN(P2_U3155) );
  INV_X1 U9644 ( .A(n7990), .ZN(n8116) );
  OAI222_X1 U9645 ( .A1(n7992), .A2(P1_U3086), .B1(n9452), .B2(n8116), .C1(
        n7991), .C2(n9450), .ZN(P1_U3330) );
  INV_X1 U9646 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7998) );
  INV_X1 U9647 ( .A(n7994), .ZN(n8256) );
  XNOR2_X1 U9648 ( .A(n7993), .B(n8341), .ZN(n7997) );
  OAI22_X1 U9649 ( .A1(n7995), .A2(n8747), .B1(n8748), .B2(n8745), .ZN(n7996)
         );
  AOI21_X1 U9650 ( .B1(n7997), .B2(n9844), .A(n7996), .ZN(n8040) );
  MUX2_X1 U9651 ( .A(n7998), .B(n8040), .S(n9891), .Z(n8001) );
  XNOR2_X1 U9652 ( .A(n7999), .B(n8341), .ZN(n8044) );
  AOI22_X1 U9653 ( .A1(n8044), .A2(n8890), .B1(n8889), .B2(n8038), .ZN(n8000)
         );
  NAND2_X1 U9654 ( .A1(n8001), .A2(n8000), .ZN(P2_U3432) );
  INV_X1 U9655 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8002) );
  MUX2_X1 U9656 ( .A(n8002), .B(n8040), .S(n9904), .Z(n8004) );
  AOI22_X1 U9657 ( .A1(n8044), .A2(n8809), .B1(n8808), .B2(n8038), .ZN(n8003)
         );
  NAND2_X1 U9658 ( .A1(n8004), .A2(n8003), .ZN(P2_U3473) );
  INV_X1 U9659 ( .A(n8099), .ZN(n8015) );
  XNOR2_X1 U9660 ( .A(n8099), .B(n8161), .ZN(n8121) );
  XNOR2_X1 U9661 ( .A(n8121), .B(n8521), .ZN(n8009) );
  NAND2_X1 U9662 ( .A1(n8010), .A2(n8009), .ZN(n8124) );
  OAI211_X1 U9663 ( .C1(n8010), .C2(n8009), .A(n8124), .B(n8508), .ZN(n8014)
         );
  NAND2_X1 U9664 ( .A1(n8510), .A2(n8522), .ZN(n8011) );
  NAND2_X1 U9665 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8539) );
  OAI211_X1 U9666 ( .C1(n8457), .C2(n8512), .A(n8011), .B(n8539), .ZN(n8012)
         );
  AOI21_X1 U9667 ( .B1(n8098), .B2(n8514), .A(n8012), .ZN(n8013) );
  OAI211_X1 U9668 ( .C1(n8015), .C2(n8517), .A(n8014), .B(n8013), .ZN(P2_U3181) );
  AOI21_X1 U9669 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8037) );
  INV_X1 U9670 ( .A(n8019), .ZN(n8020) );
  OAI21_X1 U9671 ( .B1(n9737), .B2(n8021), .A(n8020), .ZN(n8027) );
  AOI21_X1 U9672 ( .B1(n8024), .B2(n8023), .A(n8022), .ZN(n8025) );
  NOR2_X1 U9673 ( .A1(n8025), .A2(n9826), .ZN(n8026) );
  AOI211_X1 U9674 ( .C1(n9809), .C2(n8028), .A(n8027), .B(n8026), .ZN(n8036)
         );
  INV_X1 U9675 ( .A(n8029), .ZN(n8031) );
  NAND2_X1 U9676 ( .A1(n8031), .A2(n8030), .ZN(n8032) );
  XNOR2_X1 U9677 ( .A(n8033), .B(n8032), .ZN(n8034) );
  NAND2_X1 U9678 ( .A1(n8034), .A2(n9822), .ZN(n8035) );
  OAI211_X1 U9679 ( .C1(n8037), .C2(n9817), .A(n8036), .B(n8035), .ZN(P2_U3194) );
  INV_X1 U9680 ( .A(n8038), .ZN(n8039) );
  NOR2_X1 U9681 ( .A1(n8039), .A2(n9836), .ZN(n8042) );
  INV_X1 U9682 ( .A(n8040), .ZN(n8041) );
  AOI211_X1 U9683 ( .C1(n8755), .C2(n8043), .A(n8042), .B(n8041), .ZN(n8046)
         );
  AOI22_X1 U9684 ( .A1(n8044), .A2(n8759), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8586), .ZN(n8045) );
  OAI21_X1 U9685 ( .B1(n8046), .B2(n8586), .A(n8045), .ZN(P2_U3219) );
  AOI21_X1 U9686 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8050) );
  OR2_X1 U9687 ( .A1(n9817), .A2(n8050), .ZN(n8051) );
  OAI211_X1 U9688 ( .C1(n9737), .C2(n9971), .A(n8052), .B(n8051), .ZN(n8058)
         );
  AOI21_X1 U9689 ( .B1(n8055), .B2(n8054), .A(n8053), .ZN(n8056) );
  NOR2_X1 U9690 ( .A1(n8056), .A2(n9826), .ZN(n8057) );
  AOI211_X1 U9691 ( .C1(n9809), .C2(n8118), .A(n8058), .B(n8057), .ZN(n8064)
         );
  OAI21_X1 U9692 ( .B1(n8061), .B2(n8060), .A(n8059), .ZN(n8062) );
  NAND2_X1 U9693 ( .A1(n8062), .A2(n9822), .ZN(n8063) );
  NAND2_X1 U9694 ( .A1(n8064), .A2(n8063), .ZN(P2_U3195) );
  AOI21_X1 U9695 ( .B1(n8067), .B2(n8066), .A(n8065), .ZN(n8083) );
  AOI21_X1 U9696 ( .B1(n8070), .B2(n8069), .A(n8068), .ZN(n8071) );
  NOR2_X1 U9697 ( .A1(n8071), .A2(n9826), .ZN(n8081) );
  OAI22_X1 U9698 ( .A1(n9807), .A2(n8073), .B1(n9737), .B2(n8072), .ZN(n8079)
         );
  AOI21_X1 U9699 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(n8077) );
  NOR2_X1 U9700 ( .A1(n8077), .A2(n9763), .ZN(n8078) );
  NOR4_X1 U9701 ( .A1(n8081), .A2(n8080), .A3(n8079), .A4(n8078), .ZN(n8082)
         );
  OAI21_X1 U9702 ( .B1(n8083), .B2(n9817), .A(n8082), .ZN(P2_U3193) );
  INV_X1 U9703 ( .A(n8084), .ZN(n8087) );
  OAI222_X1 U9704 ( .A1(n8086), .A2(P2_U3151), .B1(n8906), .B2(n8087), .C1(
        n8085), .C2(n8899), .ZN(P2_U3269) );
  OAI222_X1 U9705 ( .A1(n8088), .A2(P1_U3086), .B1(n9452), .B2(n8087), .C1(
        n9959), .C2(n9450), .ZN(P1_U3329) );
  XNOR2_X1 U9706 ( .A(n8089), .B(n8362), .ZN(n8102) );
  XNOR2_X1 U9707 ( .A(n8090), .B(n8362), .ZN(n8091) );
  AOI222_X1 U9708 ( .A1(n9844), .A2(n8091), .B1(n8735), .B2(n9841), .C1(n8522), 
        .C2(n9840), .ZN(n8097) );
  MUX2_X1 U9709 ( .A(n8544), .B(n8097), .S(n9904), .Z(n8093) );
  NAND2_X1 U9710 ( .A1(n8099), .A2(n8808), .ZN(n8092) );
  OAI211_X1 U9711 ( .C1(n8806), .C2(n8102), .A(n8093), .B(n8092), .ZN(P2_U3474) );
  INV_X1 U9712 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8094) );
  MUX2_X1 U9713 ( .A(n8094), .B(n8097), .S(n9891), .Z(n8096) );
  NAND2_X1 U9714 ( .A1(n8099), .A2(n8889), .ZN(n8095) );
  OAI211_X1 U9715 ( .C1(n8102), .C2(n8884), .A(n8096), .B(n8095), .ZN(P2_U3435) );
  MUX2_X1 U9716 ( .A(n10033), .B(n8097), .S(n8752), .Z(n8101) );
  AOI22_X1 U9717 ( .A1(n8099), .A2(n8756), .B1(n8755), .B2(n8098), .ZN(n8100)
         );
  OAI211_X1 U9718 ( .C1(n8102), .C2(n8741), .A(n8101), .B(n8100), .ZN(P2_U3218) );
  INV_X1 U9719 ( .A(n8103), .ZN(n8106) );
  AOI21_X1 U9720 ( .B1(n8904), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8104), .ZN(
        n8105) );
  OAI21_X1 U9721 ( .B1(n8106), .B2(n8906), .A(n8105), .ZN(P2_U3268) );
  OAI222_X1 U9722 ( .A1(n8108), .A2(n8107), .B1(P1_U3086), .B2(n4294), .C1(
        n9452), .C2(n8106), .ZN(P1_U3328) );
  OAI222_X1 U9723 ( .A1(n9450), .A2(n8110), .B1(P1_U3086), .B2(n8109), .C1(
        n9452), .C2(n8112), .ZN(P1_U3326) );
  OAI222_X1 U9724 ( .A1(P2_U3151), .A2(n6328), .B1(n8906), .B2(n8112), .C1(
        n8111), .C2(n8899), .ZN(P2_U3266) );
  INV_X1 U9725 ( .A(n8113), .ZN(n8907) );
  OAI222_X1 U9726 ( .A1(n8117), .A2(P2_U3151), .B1(n8906), .B2(n8116), .C1(
        n8115), .C2(n8899), .ZN(P2_U3270) );
  AOI22_X1 U9727 ( .A1(n8118), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8904), .ZN(n8119) );
  OAI21_X1 U9728 ( .B1(n8120), .B2(n8906), .A(n8119), .ZN(P2_U3282) );
  INV_X1 U9729 ( .A(n8121), .ZN(n8122) );
  NAND2_X1 U9730 ( .A1(n8122), .A2(n8521), .ZN(n8123) );
  XNOR2_X1 U9731 ( .A(n8888), .B(n8161), .ZN(n8125) );
  XNOR2_X1 U9732 ( .A(n8125), .B(n8457), .ZN(n8443) );
  NAND2_X1 U9733 ( .A1(n8125), .A2(n8457), .ZN(n8451) );
  XNOR2_X1 U9734 ( .A(n8881), .B(n8161), .ZN(n8128) );
  NAND2_X1 U9735 ( .A1(n8128), .A2(n8746), .ZN(n8127) );
  AND2_X1 U9736 ( .A1(n8451), .A2(n8127), .ZN(n8126) );
  XNOR2_X1 U9737 ( .A(n8875), .B(n8161), .ZN(n8131) );
  XNOR2_X1 U9738 ( .A(n8131), .B(n8734), .ZN(n8495) );
  INV_X1 U9739 ( .A(n8127), .ZN(n8129) );
  XNOR2_X1 U9740 ( .A(n8128), .B(n8722), .ZN(n8452) );
  OR2_X1 U9741 ( .A1(n8129), .A2(n8452), .ZN(n8492) );
  AND2_X1 U9742 ( .A1(n8495), .A2(n8492), .ZN(n8130) );
  NAND2_X1 U9743 ( .A1(n8493), .A2(n8130), .ZN(n8133) );
  NAND2_X1 U9744 ( .A1(n8131), .A2(n8413), .ZN(n8132) );
  XNOR2_X1 U9745 ( .A(n8869), .B(n8161), .ZN(n8408) );
  AND2_X1 U9746 ( .A1(n8408), .A2(n8479), .ZN(n8134) );
  INV_X1 U9747 ( .A(n8408), .ZN(n8135) );
  NAND2_X1 U9748 ( .A1(n8135), .A2(n8723), .ZN(n8136) );
  XNOR2_X1 U9749 ( .A(n8864), .B(n8161), .ZN(n8137) );
  NAND2_X1 U9750 ( .A1(n8137), .A2(n8693), .ZN(n8419) );
  INV_X1 U9751 ( .A(n8137), .ZN(n8138) );
  NAND2_X1 U9752 ( .A1(n8138), .A2(n8713), .ZN(n8139) );
  NAND2_X1 U9753 ( .A1(n8419), .A2(n8139), .ZN(n8476) );
  NAND2_X1 U9754 ( .A1(n8141), .A2(n8140), .ZN(n8418) );
  NAND2_X1 U9755 ( .A1(n8418), .A2(n8419), .ZN(n8142) );
  XNOR2_X1 U9756 ( .A(n8792), .B(n7112), .ZN(n8144) );
  XNOR2_X1 U9757 ( .A(n8144), .B(n8703), .ZN(n8420) );
  NAND2_X1 U9758 ( .A1(n8142), .A2(n8420), .ZN(n8422) );
  NAND2_X1 U9759 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  XNOR2_X1 U9760 ( .A(n8854), .B(n8161), .ZN(n8146) );
  XNOR2_X1 U9761 ( .A(n8146), .B(n8665), .ZN(n8484) );
  INV_X1 U9762 ( .A(n8146), .ZN(n8147) );
  NAND2_X1 U9763 ( .A1(n8147), .A2(n8665), .ZN(n8148) );
  XNOR2_X1 U9764 ( .A(n8848), .B(n7795), .ZN(n8149) );
  XNOR2_X1 U9765 ( .A(n8843), .B(n8161), .ZN(n8150) );
  NAND2_X1 U9766 ( .A1(n8150), .A2(n8436), .ZN(n8153) );
  INV_X1 U9767 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U9768 ( .A1(n8151), .A2(n8666), .ZN(n8152) );
  NAND2_X1 U9769 ( .A1(n8153), .A2(n8152), .ZN(n8462) );
  AOI21_X2 U9770 ( .B1(n8400), .B2(n4892), .A(n8462), .ZN(n8464) );
  INV_X1 U9771 ( .A(n8153), .ZN(n8432) );
  XNOR2_X1 U9772 ( .A(n8837), .B(n8161), .ZN(n8154) );
  NAND2_X1 U9773 ( .A1(n8154), .A2(n8468), .ZN(n8506) );
  INV_X1 U9774 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U9775 ( .A1(n8155), .A2(n8656), .ZN(n8156) );
  AND2_X1 U9776 ( .A1(n8506), .A2(n8156), .ZN(n8431) );
  XNOR2_X1 U9777 ( .A(n8832), .B(n8161), .ZN(n8157) );
  XNOR2_X1 U9778 ( .A(n8157), .B(n8618), .ZN(n8507) );
  NOR2_X1 U9779 ( .A1(n8505), .A2(n8158), .ZN(n8394) );
  XNOR2_X1 U9780 ( .A(n8826), .B(n8161), .ZN(n8159) );
  XNOR2_X1 U9781 ( .A(n8159), .B(n8632), .ZN(n8393) );
  NAND2_X1 U9782 ( .A1(n8394), .A2(n8393), .ZN(n8392) );
  NAND2_X1 U9783 ( .A1(n8392), .A2(n8160), .ZN(n8163) );
  XNOR2_X1 U9784 ( .A(n8590), .B(n8161), .ZN(n8162) );
  XNOR2_X1 U9785 ( .A(n8163), .B(n8162), .ZN(n8170) );
  INV_X1 U9786 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8164) );
  OAI22_X1 U9787 ( .A1(n8599), .A2(n8499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8164), .ZN(n8165) );
  INV_X1 U9788 ( .A(n8165), .ZN(n8167) );
  NAND2_X1 U9789 ( .A1(n8604), .A2(n8514), .ZN(n8166) );
  OAI211_X1 U9790 ( .C1(n8600), .C2(n8512), .A(n8167), .B(n8166), .ZN(n8168)
         );
  AOI21_X1 U9791 ( .B1(n8770), .B2(n8501), .A(n8168), .ZN(n8169) );
  OAI21_X1 U9792 ( .B1(n8170), .B2(n8503), .A(n8169), .ZN(P2_U3160) );
  OAI222_X1 U9793 ( .A1(n8172), .A2(P2_U3151), .B1(n8906), .B2(n8171), .C1(
        n9961), .C2(n8899), .ZN(P2_U3271) );
  MUX2_X1 U9794 ( .A(n8619), .B(n8823), .S(n8310), .Z(n8311) );
  NAND2_X1 U9795 ( .A1(n8684), .A2(n8273), .ZN(n8174) );
  MUX2_X1 U9796 ( .A(n8177), .B(n8175), .S(n8326), .Z(n8276) );
  AND2_X1 U9797 ( .A1(n8177), .A2(n8176), .ZN(n8180) );
  AND2_X1 U9798 ( .A1(n8709), .A2(n8178), .ZN(n8179) );
  MUX2_X1 U9799 ( .A(n8180), .B(n8179), .S(n8310), .Z(n8275) );
  INV_X1 U9800 ( .A(n8181), .ZN(n8187) );
  NAND2_X1 U9801 ( .A1(n8183), .A2(n8328), .ZN(n8186) );
  NAND2_X1 U9802 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  NOR2_X1 U9803 ( .A1(n8188), .A2(n8310), .ZN(n8191) );
  AND2_X1 U9804 ( .A1(n8199), .A2(n8189), .ZN(n8190) );
  AOI21_X1 U9805 ( .B1(n8193), .B2(n8216), .A(n8326), .ZN(n8194) );
  AOI21_X1 U9806 ( .B1(n8196), .B2(n8195), .A(n8194), .ZN(n8198) );
  INV_X1 U9807 ( .A(n8199), .ZN(n8201) );
  NAND3_X1 U9808 ( .A1(n8202), .A2(n8226), .A3(n8218), .ZN(n8204) );
  INV_X1 U9809 ( .A(n8203), .ZN(n8222) );
  NAND2_X1 U9810 ( .A1(n8228), .A2(n8232), .ZN(n8205) );
  NAND4_X1 U9811 ( .A1(n8208), .A2(n7789), .A3(n8310), .A4(n8207), .ZN(n8214)
         );
  NOR2_X1 U9812 ( .A1(n8209), .A2(n8310), .ZN(n8212) );
  OAI21_X1 U9813 ( .B1(n8326), .B2(n8525), .A(n8211), .ZN(n8210) );
  OAI21_X1 U9814 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8213) );
  AND2_X1 U9815 ( .A1(n8214), .A2(n8213), .ZN(n8241) );
  NAND4_X1 U9816 ( .A1(n8236), .A2(n8326), .A3(n8215), .A4(n8526), .ZN(n8240)
         );
  INV_X1 U9817 ( .A(n8216), .ZN(n8219) );
  OAI211_X1 U9818 ( .C1(n8220), .C2(n8219), .A(n8218), .B(n8217), .ZN(n8223)
         );
  NAND3_X1 U9819 ( .A1(n8223), .A2(n8222), .A3(n8221), .ZN(n8227) );
  AND2_X1 U9820 ( .A1(n8225), .A2(n8224), .ZN(n8230) );
  NAND4_X1 U9821 ( .A1(n8227), .A2(n8348), .A3(n8230), .A4(n8226), .ZN(n8238)
         );
  AND3_X1 U9822 ( .A1(n8229), .A2(n8326), .A3(n8228), .ZN(n8237) );
  INV_X1 U9823 ( .A(n8230), .ZN(n8234) );
  AND2_X1 U9824 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  OR2_X1 U9825 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  NAND4_X1 U9826 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n8239)
         );
  NAND4_X1 U9827 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n8243)
         );
  NAND2_X1 U9828 ( .A1(n8245), .A2(n8244), .ZN(n8247) );
  MUX2_X1 U9829 ( .A(n8247), .B(n8246), .S(n8326), .Z(n8248) );
  MUX2_X1 U9830 ( .A(n8249), .B(n8523), .S(n8310), .Z(n8251) );
  INV_X1 U9831 ( .A(n8251), .ZN(n8253) );
  NAND2_X1 U9832 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  MUX2_X1 U9833 ( .A(n8256), .B(n8255), .S(n8326), .Z(n8257) );
  OR2_X1 U9834 ( .A1(n8258), .A2(n8257), .ZN(n8260) );
  INV_X1 U9835 ( .A(n8362), .ZN(n8259) );
  NAND2_X1 U9836 ( .A1(n8260), .A2(n8259), .ZN(n8266) );
  NAND3_X1 U9837 ( .A1(n8266), .A2(n8267), .A3(n8261), .ZN(n8262) );
  NAND3_X1 U9838 ( .A1(n8266), .A2(n8265), .A3(n8264), .ZN(n8268) );
  NAND2_X1 U9839 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  INV_X1 U9840 ( .A(n8732), .ZN(n8729) );
  INV_X1 U9841 ( .A(n8273), .ZN(n8274) );
  MUX2_X1 U9842 ( .A(n8279), .B(n8278), .S(n8326), .Z(n8280) );
  NAND2_X1 U9843 ( .A1(n8281), .A2(n8280), .ZN(n8288) );
  INV_X1 U9844 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U9845 ( .A1(n8288), .A2(n8283), .ZN(n8285) );
  INV_X1 U9846 ( .A(n8854), .ZN(n8491) );
  MUX2_X1 U9847 ( .A(n8694), .B(n8491), .S(n8326), .Z(n8284) );
  NAND2_X1 U9848 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  OAI21_X1 U9849 ( .B1(n8288), .B2(n8287), .A(n8286), .ZN(n8293) );
  INV_X1 U9850 ( .A(n8338), .ZN(n8290) );
  INV_X1 U9851 ( .A(n8289), .ZN(n8336) );
  OAI211_X1 U9852 ( .C1(n8293), .C2(n8290), .A(n8336), .B(n8337), .ZN(n8291)
         );
  INV_X1 U9853 ( .A(n8337), .ZN(n8292) );
  AOI21_X1 U9854 ( .B1(n8293), .B2(n8338), .A(n8292), .ZN(n8295) );
  INV_X1 U9855 ( .A(n8335), .ZN(n8294) );
  MUX2_X1 U9856 ( .A(n8297), .B(n8296), .S(n8326), .Z(n8298) );
  MUX2_X1 U9857 ( .A(n8609), .B(n8608), .S(n8326), .Z(n8299) );
  NAND2_X1 U9858 ( .A1(n8616), .A2(n8299), .ZN(n8300) );
  AOI21_X1 U9859 ( .B1(n8301), .B2(n8631), .A(n8300), .ZN(n8305) );
  MUX2_X1 U9860 ( .A(n8303), .B(n8302), .S(n8310), .Z(n8304) );
  INV_X1 U9861 ( .A(n8306), .ZN(n8332) );
  NAND2_X1 U9862 ( .A1(n8898), .A2(n8307), .ZN(n8309) );
  INV_X1 U9863 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8900) );
  OR2_X1 U9864 ( .A1(n8316), .A2(n8900), .ZN(n8308) );
  AND2_X1 U9865 ( .A1(n8817), .A2(n8520), .ZN(n8369) );
  NOR2_X1 U9866 ( .A1(n8817), .A2(n8520), .ZN(n8329) );
  INV_X1 U9867 ( .A(n8329), .ZN(n8370) );
  OAI21_X1 U9868 ( .B1(n8369), .B2(n8326), .A(n8370), .ZN(n8324) );
  INV_X1 U9869 ( .A(n8314), .ZN(n9449) );
  OAI22_X1 U9870 ( .A1(n9449), .A2(n8317), .B1(n8316), .B2(n8315), .ZN(n8763)
         );
  NAND2_X1 U9871 ( .A1(n8318), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U9872 ( .A1(n6514), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U9873 ( .A1(n6376), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8319) );
  AND3_X1 U9874 ( .A1(n8321), .A2(n8320), .A3(n8319), .ZN(n8322) );
  NOR2_X1 U9875 ( .A1(n8763), .A2(n8572), .ZN(n8334) );
  AOI211_X1 U9876 ( .C1(n8325), .C2(n8324), .A(n8334), .B(n8375), .ZN(n8381)
         );
  INV_X1 U9877 ( .A(n8325), .ZN(n8327) );
  NAND2_X1 U9878 ( .A1(n8327), .A2(n8326), .ZN(n8380) );
  INV_X1 U9879 ( .A(n8763), .ZN(n8814) );
  INV_X1 U9880 ( .A(n8572), .ZN(n8519) );
  NOR2_X1 U9881 ( .A1(n8814), .A2(n8519), .ZN(n8373) );
  AOI211_X1 U9882 ( .C1(n8369), .C2(n8763), .A(n8328), .B(n8373), .ZN(n8378)
         );
  INV_X1 U9883 ( .A(n8817), .ZN(n8767) );
  OAI22_X1 U9884 ( .A1(n8814), .A2(n8329), .B1(n8519), .B2(n8767), .ZN(n8331)
         );
  OAI211_X1 U9885 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8330), .ZN(n8377)
         );
  INV_X1 U9886 ( .A(n8334), .ZN(n8372) );
  NAND2_X1 U9887 ( .A1(n8338), .A2(n8337), .ZN(n8664) );
  INV_X1 U9888 ( .A(n8339), .ZN(n8721) );
  INV_X1 U9889 ( .A(n8340), .ZN(n8712) );
  NOR3_X1 U9890 ( .A1(n8344), .A2(n8343), .A3(n8342), .ZN(n8349) );
  NOR2_X1 U9891 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NAND4_X1 U9892 ( .A1(n8349), .A2(n6618), .A3(n8348), .A4(n8347), .ZN(n8353)
         );
  OR4_X1 U9893 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n8354) );
  NOR4_X1 U9894 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n8360)
         );
  NAND4_X1 U9895 ( .A1(n4661), .A2(n8360), .A3(n8359), .A4(n8358), .ZN(n8361)
         );
  NOR4_X1 U9896 ( .A1(n8732), .A2(n6632), .A3(n8362), .A4(n8361), .ZN(n8363)
         );
  NAND4_X1 U9897 ( .A1(n8702), .A2(n8721), .A3(n8712), .A4(n8363), .ZN(n8364)
         );
  NOR4_X1 U9898 ( .A1(n8664), .A2(n8674), .A3(n8688), .A4(n8364), .ZN(n8365)
         );
  NAND4_X1 U9899 ( .A1(n8631), .A2(n8638), .A3(n8655), .A4(n8365), .ZN(n8366)
         );
  NOR4_X1 U9900 ( .A1(n8368), .A2(n8597), .A3(n8367), .A4(n8366), .ZN(n8371)
         );
  NAND4_X1 U9901 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n4670), .ZN(n8374)
         );
  AOI21_X1 U9902 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8376) );
  AOI21_X1 U9903 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8379) );
  AOI21_X1 U9904 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8383) );
  XNOR2_X1 U9905 ( .A(n8383), .B(n8382), .ZN(n8391) );
  NOR3_X1 U9906 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(n8389) );
  OAI21_X1 U9907 ( .B1(n8390), .B2(n8387), .A(P2_B_REG_SCAN_IN), .ZN(n8388) );
  OAI22_X1 U9908 ( .A1(n8391), .A2(n8390), .B1(n8389), .B2(n8388), .ZN(
        P2_U3296) );
  INV_X1 U9909 ( .A(n8826), .ZN(n8399) );
  OAI211_X1 U9910 ( .C1(n8394), .C2(n8393), .A(n8392), .B(n8508), .ZN(n8398)
         );
  AOI22_X1 U9911 ( .A1(n8648), .A2(n8510), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8395) );
  OAI21_X1 U9912 ( .B1(n8619), .B2(n8512), .A(n8395), .ZN(n8396) );
  AOI21_X1 U9913 ( .B1(n8624), .B2(n8514), .A(n8396), .ZN(n8397) );
  OAI211_X1 U9914 ( .C1(n8399), .C2(n8517), .A(n8398), .B(n8397), .ZN(P2_U3154) );
  INV_X1 U9915 ( .A(n8848), .ZN(n8407) );
  OAI21_X1 U9916 ( .B1(n8487), .B2(n8401), .A(n8400), .ZN(n8402) );
  NAND2_X1 U9917 ( .A1(n8402), .A2(n8508), .ZN(n8406) );
  AOI22_X1 U9918 ( .A1(n8666), .A2(n8496), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8403) );
  OAI21_X1 U9919 ( .B1(n8694), .B2(n8499), .A(n8403), .ZN(n8404) );
  AOI21_X1 U9920 ( .B1(n8669), .B2(n8514), .A(n8404), .ZN(n8405) );
  OAI211_X1 U9921 ( .C1(n8407), .C2(n8517), .A(n8406), .B(n8405), .ZN(P2_U3156) );
  XNOR2_X1 U9922 ( .A(n8408), .B(n8479), .ZN(n8409) );
  XNOR2_X1 U9923 ( .A(n8410), .B(n8409), .ZN(n8417) );
  NAND2_X1 U9924 ( .A1(n8496), .A2(n8713), .ZN(n8412) );
  OAI211_X1 U9925 ( .C1(n8413), .C2(n8499), .A(n8412), .B(n8411), .ZN(n8414)
         );
  AOI21_X1 U9926 ( .B1(n8716), .B2(n8514), .A(n8414), .ZN(n8416) );
  NAND2_X1 U9927 ( .A1(n8869), .A2(n8501), .ZN(n8415) );
  OAI211_X1 U9928 ( .C1(n8417), .C2(n8503), .A(n8416), .B(n8415), .ZN(P2_U3159) );
  INV_X1 U9929 ( .A(n8792), .ZN(n8429) );
  INV_X1 U9930 ( .A(n8418), .ZN(n8474) );
  INV_X1 U9931 ( .A(n8419), .ZN(n8421) );
  NOR3_X1 U9932 ( .A1(n8474), .A2(n8421), .A3(n8420), .ZN(n8424) );
  INV_X1 U9933 ( .A(n8422), .ZN(n8423) );
  OAI21_X1 U9934 ( .B1(n8424), .B2(n8423), .A(n8508), .ZN(n8428) );
  AOI22_X1 U9935 ( .A1(n8496), .A2(n8665), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8425) );
  OAI21_X1 U9936 ( .B1(n8693), .B2(n8499), .A(n8425), .ZN(n8426) );
  AOI21_X1 U9937 ( .B1(n8695), .B2(n8514), .A(n8426), .ZN(n8427) );
  OAI211_X1 U9938 ( .C1(n8429), .C2(n8517), .A(n8428), .B(n8427), .ZN(P2_U3163) );
  INV_X1 U9939 ( .A(n8837), .ZN(n8440) );
  INV_X1 U9940 ( .A(n8430), .ZN(n8434) );
  NOR3_X1 U9941 ( .A1(n8464), .A2(n8432), .A3(n8431), .ZN(n8433) );
  OAI21_X1 U9942 ( .B1(n8434), .B2(n8433), .A(n8508), .ZN(n8439) );
  AOI22_X1 U9943 ( .A1(n8648), .A2(n8496), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8435) );
  OAI21_X1 U9944 ( .B1(n8436), .B2(n8499), .A(n8435), .ZN(n8437) );
  AOI21_X1 U9945 ( .B1(n8651), .B2(n8514), .A(n8437), .ZN(n8438) );
  OAI211_X1 U9946 ( .C1(n8440), .C2(n8517), .A(n8439), .B(n8438), .ZN(P2_U3165) );
  INV_X1 U9947 ( .A(n8441), .ZN(n8450) );
  AOI21_X1 U9948 ( .B1(n8443), .B2(n8442), .A(n8450), .ZN(n8448) );
  AOI22_X1 U9949 ( .A1(n8496), .A2(n8722), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8445) );
  NAND2_X1 U9950 ( .A1(n8514), .A2(n8754), .ZN(n8444) );
  OAI211_X1 U9951 ( .C1(n8748), .C2(n8499), .A(n8445), .B(n8444), .ZN(n8446)
         );
  AOI21_X1 U9952 ( .B1(n8888), .B2(n8501), .A(n8446), .ZN(n8447) );
  OAI21_X1 U9953 ( .B1(n8448), .B2(n8503), .A(n8447), .ZN(P2_U3166) );
  INV_X1 U9954 ( .A(n8881), .ZN(n8461) );
  INV_X1 U9955 ( .A(n8451), .ZN(n8449) );
  NOR3_X1 U9956 ( .A1(n8450), .A2(n8449), .A3(n8452), .ZN(n8455) );
  NAND2_X1 U9957 ( .A1(n8441), .A2(n8451), .ZN(n8453) );
  AND2_X1 U9958 ( .A1(n8453), .A2(n8452), .ZN(n8454) );
  OAI21_X1 U9959 ( .B1(n8455), .B2(n8454), .A(n8508), .ZN(n8460) );
  AOI22_X1 U9960 ( .A1(n8496), .A2(n8734), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8456) );
  OAI21_X1 U9961 ( .B1(n8457), .B2(n8499), .A(n8456), .ZN(n8458) );
  AOI21_X1 U9962 ( .B1(n8738), .B2(n8514), .A(n8458), .ZN(n8459) );
  OAI211_X1 U9963 ( .C1(n8461), .C2(n8517), .A(n8460), .B(n8459), .ZN(P2_U3168) );
  INV_X1 U9964 ( .A(n8843), .ZN(n8473) );
  AND3_X1 U9965 ( .A1(n8400), .A2(n4892), .A3(n8462), .ZN(n8463) );
  OAI21_X1 U9966 ( .B1(n8464), .B2(n8463), .A(n8508), .ZN(n8472) );
  INV_X1 U9967 ( .A(n8659), .ZN(n8465) );
  NOR2_X1 U9968 ( .A1(n8466), .A2(n8465), .ZN(n8470) );
  INV_X1 U9969 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8467) );
  OAI22_X1 U9970 ( .A1(n8468), .A2(n8512), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8467), .ZN(n8469) );
  AOI211_X1 U9971 ( .C1(n8510), .C2(n8678), .A(n8470), .B(n8469), .ZN(n8471)
         );
  OAI211_X1 U9972 ( .C1(n8473), .C2(n8517), .A(n8472), .B(n8471), .ZN(P2_U3169) );
  AOI21_X1 U9973 ( .B1(n8476), .B2(n8475), .A(n8474), .ZN(n8482) );
  AOI22_X1 U9974 ( .A1(n8496), .A2(n8703), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8478) );
  NAND2_X1 U9975 ( .A1(n8514), .A2(n8706), .ZN(n8477) );
  OAI211_X1 U9976 ( .C1(n8479), .C2(n8499), .A(n8478), .B(n8477), .ZN(n8480)
         );
  AOI21_X1 U9977 ( .B1(n8864), .B2(n8501), .A(n8480), .ZN(n8481) );
  OAI21_X1 U9978 ( .B1(n8482), .B2(n8503), .A(n8481), .ZN(P2_U3173) );
  OAI211_X1 U9979 ( .C1(n8485), .C2(n8484), .A(n8483), .B(n8508), .ZN(n8490)
         );
  AOI22_X1 U9980 ( .A1(n8510), .A2(n8703), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8486) );
  OAI21_X1 U9981 ( .B1(n8487), .B2(n8512), .A(n8486), .ZN(n8488) );
  AOI21_X1 U9982 ( .B1(n8681), .B2(n8514), .A(n8488), .ZN(n8489) );
  OAI211_X1 U9983 ( .C1(n8491), .C2(n8517), .A(n8490), .B(n8489), .ZN(P2_U3175) );
  AND2_X1 U9984 ( .A1(n8493), .A2(n8492), .ZN(n8494) );
  XOR2_X1 U9985 ( .A(n8495), .B(n8494), .Z(n8504) );
  AOI22_X1 U9986 ( .A1(n8496), .A2(n8723), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8498) );
  NAND2_X1 U9987 ( .A1(n8514), .A2(n8726), .ZN(n8497) );
  OAI211_X1 U9988 ( .C1(n8746), .C2(n8499), .A(n8498), .B(n8497), .ZN(n8500)
         );
  AOI21_X1 U9989 ( .B1(n8875), .B2(n8501), .A(n8500), .ZN(n8502) );
  OAI21_X1 U9990 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(P2_U3178) );
  INV_X1 U9991 ( .A(n8832), .ZN(n8518) );
  AND3_X1 U9992 ( .A1(n8430), .A2(n8507), .A3(n8506), .ZN(n8509) );
  OAI21_X1 U9993 ( .B1(n8505), .B2(n8509), .A(n8508), .ZN(n8516) );
  AOI22_X1 U9994 ( .A1(n8656), .A2(n8510), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8511) );
  OAI21_X1 U9995 ( .B1(n8599), .B2(n8512), .A(n8511), .ZN(n8513) );
  AOI21_X1 U9996 ( .B1(n8635), .B2(n8514), .A(n8513), .ZN(n8515) );
  OAI211_X1 U9997 ( .C1(n8518), .C2(n8517), .A(n8516), .B(n8515), .ZN(P2_U3180) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8519), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8520), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n6648), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8632), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8648), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10003 ( .A(n8656), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8557), .Z(
        P2_U3516) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8666), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8678), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8665), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8703), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8713), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10009 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8723), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10010 ( .A(n8734), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8557), .Z(
        P2_U3509) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8722), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8735), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8521), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10014 ( .A(n8522), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8557), .Z(
        P2_U3505) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8523), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8524), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8525), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10018 ( .A(n8526), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8557), .Z(
        P2_U3501) );
  MUX2_X1 U10019 ( .A(n8527), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8557), .Z(
        P2_U3500) );
  MUX2_X1 U10020 ( .A(n8528), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8557), .Z(
        P2_U3499) );
  MUX2_X1 U10021 ( .A(n8529), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8557), .Z(
        P2_U3498) );
  MUX2_X1 U10022 ( .A(n8530), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8557), .Z(
        P2_U3496) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8531), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10024 ( .A(n9842), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8557), .Z(
        P2_U3494) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7138), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10026 ( .A(n4293), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8557), .Z(
        P2_U3492) );
  MUX2_X1 U10027 ( .A(n8532), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8557), .Z(
        P2_U3491) );
  AOI21_X1 U10028 ( .B1(n8534), .B2(n10033), .A(n8533), .ZN(n8550) );
  OAI21_X1 U10029 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8548) );
  NAND2_X1 U10030 ( .A1(n9809), .A2(n8538), .ZN(n8540) );
  OAI211_X1 U10031 ( .C1(n8541), .C2(n9737), .A(n8540), .B(n8539), .ZN(n8547)
         );
  AOI21_X1 U10032 ( .B1(n8544), .B2(n8543), .A(n8542), .ZN(n8545) );
  NOR2_X1 U10033 ( .A1(n8545), .A2(n9826), .ZN(n8546) );
  AOI211_X1 U10034 ( .C1(n9822), .C2(n8548), .A(n8547), .B(n8546), .ZN(n8549)
         );
  OAI21_X1 U10035 ( .B1(n8550), .B2(n9817), .A(n8549), .ZN(P2_U3197) );
  AOI21_X1 U10036 ( .B1(n8553), .B2(n8552), .A(n8551), .ZN(n8569) );
  INV_X1 U10037 ( .A(n8554), .ZN(n8556) );
  NAND2_X1 U10038 ( .A1(n8556), .A2(n8555), .ZN(n8559) );
  OAI21_X1 U10039 ( .B1(n8559), .B2(n8557), .A(n9807), .ZN(n8566) );
  INV_X1 U10040 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8562) );
  INV_X1 U10041 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8560) );
  OR2_X1 U10042 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8560), .ZN(n8561) );
  OAI21_X1 U10043 ( .B1(n8569), .B2(n9817), .A(n8568), .ZN(P2_U3200) );
  INV_X1 U10044 ( .A(n8570), .ZN(n8571) );
  OAI22_X1 U10045 ( .A1(n8586), .A2(n8812), .B1(n8573), .B2(n9834), .ZN(n8575)
         );
  AOI21_X1 U10046 ( .B1(n8586), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8575), .ZN(
        n8574) );
  OAI21_X1 U10047 ( .B1(n8814), .B2(n8581), .A(n8574), .ZN(P2_U3202) );
  AOI21_X1 U10048 ( .B1(n8586), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8575), .ZN(
        n8576) );
  OAI21_X1 U10049 ( .B1(n8817), .B2(n8581), .A(n8576), .ZN(P2_U3203) );
  INV_X1 U10050 ( .A(n8577), .ZN(n8587) );
  INV_X1 U10051 ( .A(n8578), .ZN(n8584) );
  AOI22_X1 U10052 ( .A1(n8579), .A2(n8755), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8586), .ZN(n8580) );
  OAI21_X1 U10053 ( .B1(n8582), .B2(n8581), .A(n8580), .ZN(n8583) );
  AOI21_X1 U10054 ( .B1(n8584), .B2(n9848), .A(n8583), .ZN(n8585) );
  OAI21_X1 U10055 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(P2_U3204) );
  NAND2_X1 U10056 ( .A1(n8627), .A2(n8588), .ZN(n8593) );
  AND2_X1 U10057 ( .A1(n8593), .A2(n8589), .ZN(n8591) );
  NAND2_X1 U10058 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  INV_X1 U10059 ( .A(n8819), .ZN(n8607) );
  INV_X1 U10060 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9991) );
  OAI211_X1 U10061 ( .C1(n8598), .C2(n8597), .A(n8596), .B(n9844), .ZN(n8603)
         );
  OAI22_X1 U10062 ( .A1(n8600), .A2(n8745), .B1(n8599), .B2(n8747), .ZN(n8601)
         );
  INV_X1 U10063 ( .A(n8601), .ZN(n8602) );
  MUX2_X1 U10064 ( .A(n9991), .B(n8818), .S(n8752), .Z(n8606) );
  AOI22_X1 U10065 ( .A1(n8770), .A2(n8756), .B1(n8755), .B2(n8604), .ZN(n8605)
         );
  OAI211_X1 U10066 ( .C1(n8607), .C2(n8741), .A(n8606), .B(n8605), .ZN(
        P2_U3205) );
  NAND2_X1 U10067 ( .A1(n8627), .A2(n8608), .ZN(n8611) );
  AND2_X1 U10068 ( .A1(n8611), .A2(n8609), .ZN(n8613) );
  NAND2_X1 U10069 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  OAI21_X1 U10070 ( .B1(n8613), .B2(n8616), .A(n8612), .ZN(n8829) );
  INV_X1 U10071 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U10072 ( .A1(n8615), .A2(n8614), .ZN(n8617) );
  AOI21_X1 U10073 ( .B1(n8617), .B2(n8616), .A(n8692), .ZN(n8622) );
  OAI22_X1 U10074 ( .A1(n8619), .A2(n8745), .B1(n8618), .B2(n8747), .ZN(n8620)
         );
  AOI21_X1 U10075 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8824) );
  MUX2_X1 U10076 ( .A(n8623), .B(n8824), .S(n8752), .Z(n8626) );
  AOI22_X1 U10077 ( .A1(n8826), .A2(n8756), .B1(n8755), .B2(n8624), .ZN(n8625)
         );
  OAI211_X1 U10078 ( .C1(n8829), .C2(n8741), .A(n8626), .B(n8625), .ZN(
        P2_U3206) );
  XOR2_X1 U10079 ( .A(n8627), .B(n8631), .Z(n8835) );
  INV_X1 U10080 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8634) );
  XOR2_X1 U10081 ( .A(n8631), .B(n8630), .Z(n8633) );
  AOI222_X1 U10082 ( .A1(n9844), .A2(n8633), .B1(n8632), .B2(n9841), .C1(n8656), .C2(n9840), .ZN(n8830) );
  MUX2_X1 U10083 ( .A(n8634), .B(n8830), .S(n8752), .Z(n8637) );
  AOI22_X1 U10084 ( .A1(n8832), .A2(n8756), .B1(n8755), .B2(n8635), .ZN(n8636)
         );
  OAI211_X1 U10085 ( .C1(n8835), .C2(n8741), .A(n8637), .B(n8636), .ZN(
        P2_U3207) );
  XNOR2_X1 U10086 ( .A(n8639), .B(n8638), .ZN(n8840) );
  INV_X1 U10087 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8650) );
  OR2_X1 U10088 ( .A1(n8640), .A2(n8641), .ZN(n8644) );
  AND2_X1 U10089 ( .A1(n8644), .A2(n8642), .ZN(n8647) );
  NAND2_X1 U10090 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  OAI21_X1 U10091 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8649) );
  AOI222_X1 U10092 ( .A1(n9844), .A2(n8649), .B1(n8648), .B2(n9841), .C1(n8666), .C2(n9840), .ZN(n8836) );
  MUX2_X1 U10093 ( .A(n8650), .B(n8836), .S(n8752), .Z(n8653) );
  AOI22_X1 U10094 ( .A1(n8837), .A2(n8756), .B1(n8755), .B2(n8651), .ZN(n8652)
         );
  OAI211_X1 U10095 ( .C1(n8840), .C2(n8741), .A(n8653), .B(n8652), .ZN(
        P2_U3208) );
  XOR2_X1 U10096 ( .A(n8654), .B(n8655), .Z(n8846) );
  INV_X1 U10097 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8658) );
  XOR2_X1 U10098 ( .A(n8655), .B(n8640), .Z(n8657) );
  AOI222_X1 U10099 ( .A1(n9844), .A2(n8657), .B1(n8656), .B2(n9841), .C1(n8678), .C2(n9840), .ZN(n8841) );
  MUX2_X1 U10100 ( .A(n8658), .B(n8841), .S(n8752), .Z(n8661) );
  AOI22_X1 U10101 ( .A1(n8843), .A2(n8756), .B1(n8755), .B2(n8659), .ZN(n8660)
         );
  OAI211_X1 U10102 ( .C1(n8846), .C2(n8741), .A(n8661), .B(n8660), .ZN(
        P2_U3209) );
  XNOR2_X1 U10103 ( .A(n8662), .B(n8664), .ZN(n8851) );
  INV_X1 U10104 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U10105 ( .A(n8663), .B(n8664), .ZN(n8667) );
  AOI222_X1 U10106 ( .A1(n9844), .A2(n8667), .B1(n8666), .B2(n9841), .C1(n8665), .C2(n9840), .ZN(n8847) );
  MUX2_X1 U10107 ( .A(n8668), .B(n8847), .S(n8752), .Z(n8671) );
  AOI22_X1 U10108 ( .A1(n8848), .A2(n8756), .B1(n8755), .B2(n8669), .ZN(n8670)
         );
  OAI211_X1 U10109 ( .C1(n8851), .C2(n8741), .A(n8671), .B(n8670), .ZN(
        P2_U3210) );
  XOR2_X1 U10110 ( .A(n8674), .B(n8672), .Z(n8857) );
  INV_X1 U10111 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8680) );
  NAND3_X1 U10112 ( .A1(n8673), .A2(n4620), .A3(n8675), .ZN(n8676) );
  NAND2_X1 U10113 ( .A1(n8677), .A2(n8676), .ZN(n8679) );
  AOI222_X1 U10114 ( .A1(n9844), .A2(n8679), .B1(n8678), .B2(n9841), .C1(n8703), .C2(n9840), .ZN(n8852) );
  MUX2_X1 U10115 ( .A(n8680), .B(n8852), .S(n8752), .Z(n8683) );
  AOI22_X1 U10116 ( .A1(n8854), .A2(n8756), .B1(n8755), .B2(n8681), .ZN(n8682)
         );
  OAI211_X1 U10117 ( .C1(n8857), .C2(n8741), .A(n8683), .B(n8682), .ZN(
        P2_U3211) );
  NAND2_X1 U10118 ( .A1(n8685), .A2(n8684), .ZN(n8686) );
  XNOR2_X1 U10119 ( .A(n8686), .B(n8688), .ZN(n8861) );
  NAND3_X1 U10120 ( .A1(n8687), .A2(n4616), .A3(n8689), .ZN(n8690) );
  AND2_X1 U10121 ( .A1(n8673), .A2(n8690), .ZN(n8691) );
  OAI222_X1 U10122 ( .A1(n8745), .A2(n8694), .B1(n8747), .B2(n8693), .C1(n8692), .C2(n8691), .ZN(n8791) );
  NAND2_X1 U10123 ( .A1(n8791), .A2(n8752), .ZN(n8700) );
  INV_X1 U10124 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8697) );
  INV_X1 U10125 ( .A(n8695), .ZN(n8696) );
  OAI22_X1 U10126 ( .A1(n8752), .A2(n8697), .B1(n8696), .B2(n9834), .ZN(n8698)
         );
  AOI21_X1 U10127 ( .B1(n8792), .B2(n8756), .A(n8698), .ZN(n8699) );
  OAI211_X1 U10128 ( .C1(n8861), .C2(n8741), .A(n8700), .B(n8699), .ZN(
        P2_U3212) );
  XOR2_X1 U10129 ( .A(n8701), .B(n8702), .Z(n8867) );
  INV_X1 U10130 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8705) );
  OAI21_X1 U10131 ( .B1(n4309), .B2(n6639), .A(n8687), .ZN(n8704) );
  AOI222_X1 U10132 ( .A1(n9844), .A2(n8704), .B1(n8703), .B2(n9841), .C1(n8723), .C2(n9840), .ZN(n8862) );
  MUX2_X1 U10133 ( .A(n8705), .B(n8862), .S(n8752), .Z(n8708) );
  AOI22_X1 U10134 ( .A1(n8864), .A2(n8756), .B1(n8755), .B2(n8706), .ZN(n8707)
         );
  OAI211_X1 U10135 ( .C1(n8867), .C2(n8741), .A(n8708), .B(n8707), .ZN(
        P2_U3213) );
  NAND2_X1 U10136 ( .A1(n8719), .A2(n8709), .ZN(n8710) );
  XNOR2_X1 U10137 ( .A(n8710), .B(n8712), .ZN(n8872) );
  INV_X1 U10138 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8715) );
  XNOR2_X1 U10139 ( .A(n8711), .B(n8712), .ZN(n8714) );
  AOI222_X1 U10140 ( .A1(n9844), .A2(n8714), .B1(n8734), .B2(n9840), .C1(n8713), .C2(n9841), .ZN(n8868) );
  MUX2_X1 U10141 ( .A(n8715), .B(n8868), .S(n8752), .Z(n8718) );
  AOI22_X1 U10142 ( .A1(n8869), .A2(n8756), .B1(n8755), .B2(n8716), .ZN(n8717)
         );
  OAI211_X1 U10143 ( .C1(n8872), .C2(n8741), .A(n8718), .B(n8717), .ZN(
        P2_U3214) );
  OAI21_X1 U10144 ( .B1(n4375), .B2(n8721), .A(n8719), .ZN(n8878) );
  INV_X1 U10145 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U10146 ( .A(n8720), .B(n8721), .ZN(n8724) );
  AOI222_X1 U10147 ( .A1(n9844), .A2(n8724), .B1(n8723), .B2(n9841), .C1(n8722), .C2(n9840), .ZN(n8873) );
  MUX2_X1 U10148 ( .A(n8725), .B(n8873), .S(n8752), .Z(n8728) );
  AOI22_X1 U10149 ( .A1(n8875), .A2(n8756), .B1(n8755), .B2(n8726), .ZN(n8727)
         );
  OAI211_X1 U10150 ( .C1(n8878), .C2(n8741), .A(n8728), .B(n8727), .ZN(
        P2_U3215) );
  XNOR2_X1 U10151 ( .A(n8730), .B(n8729), .ZN(n8885) );
  OAI211_X1 U10152 ( .C1(n8733), .C2(n8732), .A(n8731), .B(n9844), .ZN(n8737)
         );
  AOI22_X1 U10153 ( .A1(n8735), .A2(n9840), .B1(n9841), .B2(n8734), .ZN(n8736)
         );
  MUX2_X1 U10154 ( .A(n9816), .B(n8879), .S(n8752), .Z(n8740) );
  AOI22_X1 U10155 ( .A1(n8881), .A2(n8756), .B1(n8755), .B2(n8738), .ZN(n8739)
         );
  OAI211_X1 U10156 ( .C1(n8885), .C2(n8741), .A(n8740), .B(n8739), .ZN(
        P2_U3216) );
  NAND2_X1 U10157 ( .A1(n8743), .A2(n8757), .ZN(n8744) );
  NAND3_X1 U10158 ( .A1(n8742), .A2(n9844), .A3(n8744), .ZN(n8751) );
  OAI22_X1 U10159 ( .A1(n8748), .A2(n8747), .B1(n8746), .B2(n8745), .ZN(n8749)
         );
  INV_X1 U10160 ( .A(n8749), .ZN(n8750) );
  MUX2_X1 U10161 ( .A(n8753), .B(n8886), .S(n8752), .Z(n8762) );
  AOI22_X1 U10162 ( .A1(n8888), .A2(n8756), .B1(n8755), .B2(n8754), .ZN(n8761)
         );
  XNOR2_X1 U10163 ( .A(n8758), .B(n8757), .ZN(n8891) );
  NAND2_X1 U10164 ( .A1(n8891), .A2(n8759), .ZN(n8760) );
  NAND3_X1 U10165 ( .A1(n8762), .A2(n8761), .A3(n8760), .ZN(P2_U3217) );
  INV_X1 U10166 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U10167 ( .A1(n8763), .A2(n8808), .ZN(n8765) );
  INV_X1 U10168 ( .A(n8812), .ZN(n8764) );
  NAND2_X1 U10169 ( .A1(n8764), .A2(n9904), .ZN(n8768) );
  OAI211_X1 U10170 ( .C1(n9904), .C2(n8766), .A(n8765), .B(n8768), .ZN(
        P2_U3490) );
  NAND2_X1 U10171 ( .A1(n8767), .A2(n8808), .ZN(n8769) );
  OAI211_X1 U10172 ( .C1(n9904), .C2(n6656), .A(n8769), .B(n8768), .ZN(
        P2_U3489) );
  MUX2_X1 U10173 ( .A(n9962), .B(n8818), .S(n9904), .Z(n8772) );
  AOI22_X1 U10174 ( .A1(n8819), .A2(n8809), .B1(n8808), .B2(n8770), .ZN(n8771)
         );
  NAND2_X1 U10175 ( .A1(n8772), .A2(n8771), .ZN(P2_U3487) );
  MUX2_X1 U10176 ( .A(n8773), .B(n8824), .S(n9904), .Z(n8775) );
  NAND2_X1 U10177 ( .A1(n8826), .A2(n8808), .ZN(n8774) );
  OAI211_X1 U10178 ( .C1(n8806), .C2(n8829), .A(n8775), .B(n8774), .ZN(
        P2_U3486) );
  MUX2_X1 U10179 ( .A(n8776), .B(n8830), .S(n9904), .Z(n8778) );
  NAND2_X1 U10180 ( .A1(n8832), .A2(n8808), .ZN(n8777) );
  OAI211_X1 U10181 ( .C1(n8835), .C2(n8806), .A(n8778), .B(n8777), .ZN(
        P2_U3485) );
  INV_X1 U10182 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8779) );
  MUX2_X1 U10183 ( .A(n8779), .B(n8836), .S(n9904), .Z(n8781) );
  NAND2_X1 U10184 ( .A1(n8837), .A2(n8808), .ZN(n8780) );
  OAI211_X1 U10185 ( .C1(n8840), .C2(n8806), .A(n8781), .B(n8780), .ZN(
        P2_U3484) );
  MUX2_X1 U10186 ( .A(n8782), .B(n8841), .S(n9904), .Z(n8784) );
  NAND2_X1 U10187 ( .A1(n8843), .A2(n8808), .ZN(n8783) );
  OAI211_X1 U10188 ( .C1(n8806), .C2(n8846), .A(n8784), .B(n8783), .ZN(
        P2_U3483) );
  MUX2_X1 U10189 ( .A(n8785), .B(n8847), .S(n9904), .Z(n8787) );
  NAND2_X1 U10190 ( .A1(n8848), .A2(n8808), .ZN(n8786) );
  OAI211_X1 U10191 ( .C1(n8806), .C2(n8851), .A(n8787), .B(n8786), .ZN(
        P2_U3482) );
  MUX2_X1 U10192 ( .A(n8788), .B(n8852), .S(n9904), .Z(n8790) );
  NAND2_X1 U10193 ( .A1(n8854), .A2(n8808), .ZN(n8789) );
  OAI211_X1 U10194 ( .C1(n8806), .C2(n8857), .A(n8790), .B(n8789), .ZN(
        P2_U3481) );
  INV_X1 U10195 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8793) );
  AOI21_X1 U10196 ( .B1(n9890), .B2(n8792), .A(n8791), .ZN(n8858) );
  MUX2_X1 U10197 ( .A(n8793), .B(n8858), .S(n9904), .Z(n8794) );
  OAI21_X1 U10198 ( .B1(n8806), .B2(n8861), .A(n8794), .ZN(P2_U3480) );
  INV_X1 U10199 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8795) );
  MUX2_X1 U10200 ( .A(n8795), .B(n8862), .S(n9904), .Z(n8797) );
  NAND2_X1 U10201 ( .A1(n8864), .A2(n8808), .ZN(n8796) );
  OAI211_X1 U10202 ( .C1(n8806), .C2(n8867), .A(n8797), .B(n8796), .ZN(
        P2_U3479) );
  INV_X1 U10203 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8798) );
  MUX2_X1 U10204 ( .A(n8798), .B(n8868), .S(n9904), .Z(n8800) );
  NAND2_X1 U10205 ( .A1(n8869), .A2(n8808), .ZN(n8799) );
  OAI211_X1 U10206 ( .C1(n8872), .C2(n8806), .A(n8800), .B(n8799), .ZN(
        P2_U3478) );
  INV_X1 U10207 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U10208 ( .A(n8801), .B(n8873), .S(n9904), .Z(n8803) );
  NAND2_X1 U10209 ( .A1(n8875), .A2(n8808), .ZN(n8802) );
  OAI211_X1 U10210 ( .C1(n8806), .C2(n8878), .A(n8803), .B(n8802), .ZN(
        P2_U3477) );
  MUX2_X1 U10211 ( .A(n9813), .B(n8879), .S(n9904), .Z(n8805) );
  NAND2_X1 U10212 ( .A1(n8881), .A2(n8808), .ZN(n8804) );
  OAI211_X1 U10213 ( .C1(n8885), .C2(n8806), .A(n8805), .B(n8804), .ZN(
        P2_U3476) );
  MUX2_X1 U10214 ( .A(n8807), .B(n8886), .S(n9904), .Z(n8811) );
  AOI22_X1 U10215 ( .A1(n8891), .A2(n8809), .B1(n8808), .B2(n8888), .ZN(n8810)
         );
  NAND2_X1 U10216 ( .A1(n8811), .A2(n8810), .ZN(P2_U3475) );
  NOR2_X1 U10217 ( .A1(n8812), .A2(n9893), .ZN(n8815) );
  AOI21_X1 U10218 ( .B1(n9893), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8815), .ZN(
        n8813) );
  OAI21_X1 U10219 ( .B1(n8814), .B2(n8822), .A(n8813), .ZN(P2_U3458) );
  AOI21_X1 U10220 ( .B1(n9893), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8815), .ZN(
        n8816) );
  OAI21_X1 U10221 ( .B1(n8817), .B2(n8822), .A(n8816), .ZN(P2_U3457) );
  INV_X1 U10222 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10047) );
  MUX2_X1 U10223 ( .A(n10047), .B(n8818), .S(n9891), .Z(n8821) );
  NAND2_X1 U10224 ( .A1(n8819), .A2(n8890), .ZN(n8820) );
  OAI211_X1 U10225 ( .C1(n8823), .C2(n8822), .A(n8821), .B(n8820), .ZN(
        P2_U3455) );
  INV_X1 U10226 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8825) );
  MUX2_X1 U10227 ( .A(n8825), .B(n8824), .S(n9891), .Z(n8828) );
  NAND2_X1 U10228 ( .A1(n8826), .A2(n8889), .ZN(n8827) );
  OAI211_X1 U10229 ( .C1(n8829), .C2(n8884), .A(n8828), .B(n8827), .ZN(
        P2_U3454) );
  INV_X1 U10230 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U10231 ( .A(n8831), .B(n8830), .S(n9891), .Z(n8834) );
  NAND2_X1 U10232 ( .A1(n8832), .A2(n8889), .ZN(n8833) );
  OAI211_X1 U10233 ( .C1(n8835), .C2(n8884), .A(n8834), .B(n8833), .ZN(
        P2_U3453) );
  MUX2_X1 U10234 ( .A(n10005), .B(n8836), .S(n9891), .Z(n8839) );
  NAND2_X1 U10235 ( .A1(n8837), .A2(n8889), .ZN(n8838) );
  OAI211_X1 U10236 ( .C1(n8840), .C2(n8884), .A(n8839), .B(n8838), .ZN(
        P2_U3452) );
  INV_X1 U10237 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U10238 ( .A(n8842), .B(n8841), .S(n9891), .Z(n8845) );
  NAND2_X1 U10239 ( .A1(n8843), .A2(n8889), .ZN(n8844) );
  OAI211_X1 U10240 ( .C1(n8846), .C2(n8884), .A(n8845), .B(n8844), .ZN(
        P2_U3451) );
  INV_X1 U10241 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U10242 ( .A(n9970), .B(n8847), .S(n9891), .Z(n8850) );
  NAND2_X1 U10243 ( .A1(n8848), .A2(n8889), .ZN(n8849) );
  OAI211_X1 U10244 ( .C1(n8851), .C2(n8884), .A(n8850), .B(n8849), .ZN(
        P2_U3450) );
  INV_X1 U10245 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8853) );
  MUX2_X1 U10246 ( .A(n8853), .B(n8852), .S(n9891), .Z(n8856) );
  NAND2_X1 U10247 ( .A1(n8854), .A2(n8889), .ZN(n8855) );
  OAI211_X1 U10248 ( .C1(n8857), .C2(n8884), .A(n8856), .B(n8855), .ZN(
        P2_U3449) );
  INV_X1 U10249 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8859) );
  MUX2_X1 U10250 ( .A(n8859), .B(n8858), .S(n9891), .Z(n8860) );
  OAI21_X1 U10251 ( .B1(n8861), .B2(n8884), .A(n8860), .ZN(P2_U3448) );
  INV_X1 U10252 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8863) );
  MUX2_X1 U10253 ( .A(n8863), .B(n8862), .S(n9891), .Z(n8866) );
  NAND2_X1 U10254 ( .A1(n8864), .A2(n8889), .ZN(n8865) );
  OAI211_X1 U10255 ( .C1(n8867), .C2(n8884), .A(n8866), .B(n8865), .ZN(
        P2_U3447) );
  INV_X1 U10256 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U10257 ( .A(n9998), .B(n8868), .S(n9891), .Z(n8871) );
  NAND2_X1 U10258 ( .A1(n8869), .A2(n8889), .ZN(n8870) );
  OAI211_X1 U10259 ( .C1(n8872), .C2(n8884), .A(n8871), .B(n8870), .ZN(
        P2_U3446) );
  INV_X1 U10260 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8874) );
  MUX2_X1 U10261 ( .A(n8874), .B(n8873), .S(n9891), .Z(n8877) );
  NAND2_X1 U10262 ( .A1(n8875), .A2(n8889), .ZN(n8876) );
  OAI211_X1 U10263 ( .C1(n8878), .C2(n8884), .A(n8877), .B(n8876), .ZN(
        P2_U3444) );
  INV_X1 U10264 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U10265 ( .A(n8880), .B(n8879), .S(n9891), .Z(n8883) );
  NAND2_X1 U10266 ( .A1(n8881), .A2(n8889), .ZN(n8882) );
  OAI211_X1 U10267 ( .C1(n8885), .C2(n8884), .A(n8883), .B(n8882), .ZN(
        P2_U3441) );
  INV_X1 U10268 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8887) );
  MUX2_X1 U10269 ( .A(n8887), .B(n8886), .S(n9891), .Z(n8893) );
  AOI22_X1 U10270 ( .A1(n8891), .A2(n8890), .B1(n8889), .B2(n8888), .ZN(n8892)
         );
  NAND2_X1 U10271 ( .A1(n8893), .A2(n8892), .ZN(P2_U3438) );
  INV_X1 U10272 ( .A(n8894), .ZN(n8895) );
  NOR4_X1 U10273 ( .A1(n8895), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5694), .ZN(n8896) );
  AOI21_X1 U10274 ( .B1(n8904), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8896), .ZN(
        n8897) );
  OAI21_X1 U10275 ( .B1(n9449), .B2(n8906), .A(n8897), .ZN(P2_U3264) );
  INV_X1 U10276 ( .A(n8898), .ZN(n9451) );
  OAI222_X1 U10277 ( .A1(n8902), .A2(P2_U3151), .B1(n8901), .B2(n9451), .C1(
        n8900), .C2(n8899), .ZN(P2_U3265) );
  AOI21_X1 U10278 ( .B1(n8904), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8903), .ZN(
        n8905) );
  OAI21_X1 U10279 ( .B1(n8907), .B2(n8906), .A(n8905), .ZN(P2_U3267) );
  XOR2_X1 U10280 ( .A(n8910), .B(n8909), .Z(n8915) );
  AOI22_X1 U10281 ( .A1(n9026), .A2(n8983), .B1(n8982), .B2(n9028), .ZN(n9231)
         );
  INV_X1 U10282 ( .A(n8911), .ZN(n9238) );
  AOI22_X1 U10283 ( .A1(n9238), .A2(n9013), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8912) );
  OAI21_X1 U10284 ( .B1(n9231), .B2(n9011), .A(n8912), .ZN(n8913) );
  AOI21_X1 U10285 ( .B1(n9235), .B2(n8968), .A(n8913), .ZN(n8914) );
  OAI21_X1 U10286 ( .B1(n8915), .B2(n8988), .A(n8914), .ZN(P1_U3216) );
  XOR2_X1 U10287 ( .A(n8917), .B(n8916), .Z(n8923) );
  OAI22_X1 U10288 ( .A1(n8919), .A2(n8995), .B1(n8918), .B2(n8993), .ZN(n9299)
         );
  AOI22_X1 U10289 ( .A1(n9299), .A2(n9001), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8920) );
  OAI21_X1 U10290 ( .B1(n9293), .B2(n8998), .A(n8920), .ZN(n8921) );
  AOI21_X1 U10291 ( .B1(n9380), .B2(n8968), .A(n8921), .ZN(n8922) );
  OAI21_X1 U10292 ( .B1(n8923), .B2(n8988), .A(n8922), .ZN(P1_U3219) );
  XOR2_X1 U10293 ( .A(n8925), .B(n8924), .Z(n8932) );
  NAND2_X1 U10294 ( .A1(n9028), .A2(n8983), .ZN(n8928) );
  NAND2_X1 U10295 ( .A1(n8926), .A2(n8982), .ZN(n8927) );
  NAND2_X1 U10296 ( .A1(n8928), .A2(n8927), .ZN(n9259) );
  AOI22_X1 U10297 ( .A1(n9259), .A2(n9001), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8929) );
  OAI21_X1 U10298 ( .B1(n9267), .B2(n8998), .A(n8929), .ZN(n8930) );
  AOI21_X1 U10299 ( .B1(n9427), .B2(n8968), .A(n8930), .ZN(n8931) );
  OAI21_X1 U10300 ( .B1(n8932), .B2(n8988), .A(n8931), .ZN(P1_U3223) );
  XOR2_X1 U10301 ( .A(n8934), .B(n8933), .Z(n8939) );
  AOI22_X1 U10302 ( .A1(n9024), .A2(n8983), .B1(n8982), .B2(n9026), .ZN(n9205)
         );
  NOR2_X1 U10303 ( .A1(n9205), .A2(n9011), .ZN(n8937) );
  OAI22_X1 U10304 ( .A1(n9201), .A2(n8998), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8935), .ZN(n8936) );
  AOI211_X1 U10305 ( .C1(n9348), .C2(n8968), .A(n8937), .B(n8936), .ZN(n8938)
         );
  OAI21_X1 U10306 ( .B1(n8939), .B2(n8988), .A(n8938), .ZN(P1_U3225) );
  XOR2_X1 U10307 ( .A(n8941), .B(n8940), .Z(n8948) );
  AOI22_X1 U10308 ( .A1(n8942), .A2(n9001), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n8943) );
  OAI21_X1 U10309 ( .B1(n8944), .B2(n8998), .A(n8943), .ZN(n8945) );
  AOI21_X1 U10310 ( .B1(n8946), .B2(n8968), .A(n8945), .ZN(n8947) );
  OAI21_X1 U10311 ( .B1(n8948), .B2(n8988), .A(n8947), .ZN(P1_U3226) );
  OAI211_X1 U10312 ( .C1(n4371), .C2(n8950), .A(n8949), .B(n9007), .ZN(n8955)
         );
  AND2_X1 U10313 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9074) );
  NOR2_X1 U10314 ( .A1(n8998), .A2(n8951), .ZN(n8952) );
  AOI211_X1 U10315 ( .C1(n9001), .C2(n8953), .A(n9074), .B(n8952), .ZN(n8954)
         );
  OAI211_X1 U10316 ( .C1(n4542), .C2(n9017), .A(n8955), .B(n8954), .ZN(
        P1_U3228) );
  XOR2_X1 U10317 ( .A(n8957), .B(n8956), .Z(n8963) );
  AND2_X1 U10318 ( .A1(n9027), .A2(n8982), .ZN(n8958) );
  AOI21_X1 U10319 ( .B1(n9025), .B2(n8983), .A(n8958), .ZN(n9222) );
  INV_X1 U10320 ( .A(n8959), .ZN(n9218) );
  AOI22_X1 U10321 ( .A1(n9218), .A2(n9013), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8960) );
  OAI21_X1 U10322 ( .B1(n9222), .B2(n9011), .A(n8960), .ZN(n8961) );
  AOI21_X1 U10323 ( .B1(n9354), .B2(n8968), .A(n8961), .ZN(n8962) );
  OAI21_X1 U10324 ( .B1(n8963), .B2(n8988), .A(n8962), .ZN(P1_U3229) );
  XOR2_X1 U10325 ( .A(n8965), .B(n8964), .Z(n8971) );
  AND2_X1 U10326 ( .A1(n9030), .A2(n8982), .ZN(n8966) );
  AOI21_X1 U10327 ( .B1(n9029), .B2(n8983), .A(n8966), .ZN(n9281) );
  OAI22_X1 U10328 ( .A1(n9281), .A2(n9011), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10064), .ZN(n8967) );
  AOI21_X1 U10329 ( .B1(n9286), .B2(n9013), .A(n8967), .ZN(n8970) );
  NAND2_X1 U10330 ( .A1(n9377), .A2(n8968), .ZN(n8969) );
  OAI211_X1 U10331 ( .C1(n8971), .C2(n8988), .A(n8970), .B(n8969), .ZN(
        P1_U3233) );
  OAI21_X1 U10332 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8975) );
  NAND2_X1 U10333 ( .A1(n8975), .A2(n9007), .ZN(n8979) );
  AOI22_X1 U10334 ( .A1(n9027), .A2(n8983), .B1(n8982), .B2(n9029), .ZN(n9246)
         );
  OAI22_X1 U10335 ( .A1(n9246), .A2(n9011), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8976), .ZN(n8977) );
  AOI21_X1 U10336 ( .B1(n9252), .B2(n9013), .A(n8977), .ZN(n8978) );
  OAI211_X1 U10337 ( .C1(n9424), .C2(n9017), .A(n8979), .B(n8978), .ZN(
        P1_U3235) );
  AOI21_X1 U10338 ( .B1(n8981), .B2(n8980), .A(n4378), .ZN(n8989) );
  AOI22_X1 U10339 ( .A1(n9030), .A2(n8983), .B1(n8982), .B2(n9032), .ZN(n9314)
         );
  OAI22_X1 U10340 ( .A1(n9011), .A2(n9314), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8984), .ZN(n8986) );
  NOR2_X1 U10341 ( .A1(n9437), .A2(n9017), .ZN(n8985) );
  AOI211_X1 U10342 ( .C1(n9013), .C2(n9318), .A(n8986), .B(n8985), .ZN(n8987)
         );
  OAI21_X1 U10343 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(P1_U3238) );
  OAI211_X1 U10344 ( .C1(n8992), .C2(n8991), .A(n8990), .B(n9007), .ZN(n9003)
         );
  OAI22_X1 U10345 ( .A1(n8996), .A2(n8995), .B1(n8994), .B2(n8993), .ZN(n9188)
         );
  INV_X1 U10346 ( .A(n9193), .ZN(n8999) );
  OAI22_X1 U10347 ( .A1(n8999), .A2(n8998), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8997), .ZN(n9000) );
  AOI21_X1 U10348 ( .B1(n9188), .B2(n9001), .A(n9000), .ZN(n9002) );
  OAI211_X1 U10349 ( .C1(n9413), .C2(n9017), .A(n9003), .B(n9002), .ZN(
        P1_U3240) );
  OAI21_X1 U10350 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9008) );
  NAND2_X1 U10351 ( .A1(n9008), .A2(n9007), .ZN(n9016) );
  OAI22_X1 U10352 ( .A1(n9011), .A2(n9010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9009), .ZN(n9012) );
  AOI21_X1 U10353 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9015) );
  OAI211_X1 U10354 ( .C1(n9018), .C2(n9017), .A(n9016), .B(n9015), .ZN(
        P1_U3241) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9019), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9020), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9021), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9022), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9023), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9024), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9025), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9026), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9027), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9028), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10365 ( .A(n9029), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9046), .Z(
        P1_U3575) );
  MUX2_X1 U10366 ( .A(n9030), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9046), .Z(
        P1_U3573) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9031), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9032), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10369 ( .A(n9033), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9046), .Z(
        P1_U3570) );
  MUX2_X1 U10370 ( .A(n9034), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9046), .Z(
        P1_U3569) );
  MUX2_X1 U10371 ( .A(n9035), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9046), .Z(
        P1_U3568) );
  MUX2_X1 U10372 ( .A(n9036), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9046), .Z(
        P1_U3567) );
  MUX2_X1 U10373 ( .A(n9037), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9046), .Z(
        P1_U3565) );
  MUX2_X1 U10374 ( .A(n9038), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9046), .Z(
        P1_U3564) );
  MUX2_X1 U10375 ( .A(n9039), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9046), .Z(
        P1_U3563) );
  MUX2_X1 U10376 ( .A(n9040), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9046), .Z(
        P1_U3562) );
  MUX2_X1 U10377 ( .A(n9041), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9046), .Z(
        P1_U3561) );
  MUX2_X1 U10378 ( .A(n9042), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9046), .Z(
        P1_U3560) );
  MUX2_X1 U10379 ( .A(n9043), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9046), .Z(
        P1_U3559) );
  MUX2_X1 U10380 ( .A(n9044), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9046), .Z(
        P1_U3558) );
  MUX2_X1 U10381 ( .A(n9045), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9046), .Z(
        P1_U3557) );
  MUX2_X1 U10382 ( .A(n5855), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9046), .Z(
        P1_U3556) );
  MUX2_X1 U10383 ( .A(n9047), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9046), .Z(
        P1_U3555) );
  NAND2_X1 U10384 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  NAND2_X1 U10385 ( .A1(n9051), .A2(n9050), .ZN(n9054) );
  INV_X1 U10386 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9460) );
  NOR2_X1 U10387 ( .A1(n9070), .A2(n9460), .ZN(n9052) );
  AOI21_X1 U10388 ( .B1(n9070), .B2(n9460), .A(n9052), .ZN(n9053) );
  NOR2_X1 U10389 ( .A1(n9053), .A2(n9054), .ZN(n9077) );
  AOI21_X1 U10390 ( .B1(n9054), .B2(n9053), .A(n9077), .ZN(n9068) );
  NOR2_X1 U10391 ( .A1(n9056), .A2(n9055), .ZN(n9058) );
  NOR2_X1 U10392 ( .A1(n9058), .A2(n9057), .ZN(n9061) );
  NAND2_X1 U10393 ( .A1(n9070), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9059) );
  OAI21_X1 U10394 ( .B1(n9070), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9059), .ZN(
        n9060) );
  NOR2_X1 U10395 ( .A1(n9061), .A2(n9060), .ZN(n9069) );
  AOI211_X1 U10396 ( .C1(n9061), .C2(n9060), .A(n9069), .B(n9486), .ZN(n9062)
         );
  INV_X1 U10397 ( .A(n9062), .ZN(n9066) );
  AND2_X1 U10398 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9064) );
  NOR2_X1 U10399 ( .A1(n9498), .A2(n9078), .ZN(n9063) );
  AOI211_X1 U10400 ( .C1(n9490), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9064), .B(
        n9063), .ZN(n9065) );
  OAI211_X1 U10401 ( .C1(n9068), .C2(n9067), .A(n9066), .B(n9065), .ZN(
        P1_U3259) );
  AOI21_X1 U10402 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9070), .A(n9069), .ZN(
        n9072) );
  MUX2_X1 U10403 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n9088), .S(n9083), .Z(n9071) );
  NAND2_X1 U10404 ( .A1(n9072), .A2(n9071), .ZN(n9090) );
  OAI21_X1 U10405 ( .B1(n9072), .B2(n9071), .A(n9090), .ZN(n9073) );
  NAND2_X1 U10406 ( .A1(n9073), .A2(n9116), .ZN(n9087) );
  AOI21_X1 U10407 ( .B1(n9490), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9074), .ZN(
        n9086) );
  INV_X1 U10408 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U10409 ( .A1(n9083), .A2(n9076), .ZN(n9075) );
  OAI21_X1 U10410 ( .B1(n9083), .B2(n9076), .A(n9075), .ZN(n9081) );
  AOI21_X1 U10411 ( .B1(n9078), .B2(n9460), .A(n9077), .ZN(n9079) );
  INV_X1 U10412 ( .A(n9079), .ZN(n9080) );
  NAND2_X1 U10413 ( .A1(n9081), .A2(n9080), .ZN(n9100) );
  OAI21_X1 U10414 ( .B1(n9081), .B2(n9080), .A(n9100), .ZN(n9082) );
  NAND2_X1 U10415 ( .A1(n9492), .A2(n9082), .ZN(n9085) );
  NAND2_X1 U10416 ( .A1(n9478), .A2(n9083), .ZN(n9084) );
  NAND4_X1 U10417 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(
        P1_U3260) );
  INV_X1 U10418 ( .A(n9111), .ZN(n9106) );
  AND2_X1 U10419 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U10420 ( .A1(n9098), .A2(n9088), .ZN(n9089) );
  NAND2_X1 U10421 ( .A1(n9090), .A2(n9089), .ZN(n9095) );
  INV_X1 U10422 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9091) );
  OR2_X1 U10423 ( .A1(n9111), .A2(n9091), .ZN(n9093) );
  NAND2_X1 U10424 ( .A1(n9111), .A2(n9091), .ZN(n9092) );
  AND2_X1 U10425 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  NOR2_X1 U10426 ( .A1(n9095), .A2(n9094), .ZN(n9108) );
  AOI211_X1 U10427 ( .C1(n9095), .C2(n9094), .A(n9108), .B(n9486), .ZN(n9096)
         );
  AOI211_X1 U10428 ( .C1(n9490), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9097), .B(
        n9096), .ZN(n9105) );
  NAND2_X1 U10429 ( .A1(n9098), .A2(n9076), .ZN(n9099) );
  NAND2_X1 U10430 ( .A1(n9100), .A2(n9099), .ZN(n9102) );
  XNOR2_X1 U10431 ( .A(n9111), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10432 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  NAND3_X1 U10433 ( .A1(n9492), .A2(n9113), .A3(n9103), .ZN(n9104) );
  OAI211_X1 U10434 ( .C1(n9498), .C2(n9106), .A(n9105), .B(n9104), .ZN(
        P1_U3261) );
  AND2_X1 U10435 ( .A1(n9111), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9107) );
  OR2_X1 U10436 ( .A1(n9108), .A2(n9107), .ZN(n9110) );
  XNOR2_X1 U10437 ( .A(n9110), .B(n9109), .ZN(n9117) );
  NAND2_X1 U10438 ( .A1(n9111), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10439 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  XNOR2_X1 U10440 ( .A(n9114), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9118) );
  INV_X1 U10441 ( .A(n9118), .ZN(n9115) );
  AOI22_X1 U10442 ( .A1(n9117), .A2(n9116), .B1(n9492), .B2(n9115), .ZN(n9120)
         );
  NAND2_X1 U10443 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9121) );
  XNOR2_X1 U10444 ( .A(n9131), .B(n9398), .ZN(n9123) );
  NAND2_X1 U10445 ( .A1(n9327), .A2(n9554), .ZN(n9127) );
  NOR2_X1 U10446 ( .A1(n9125), .A2(n9124), .ZN(n9326) );
  INV_X1 U10447 ( .A(n9326), .ZN(n9330) );
  NOR2_X1 U10448 ( .A1(n9543), .A2(n9330), .ZN(n9132) );
  AOI21_X1 U10449 ( .B1(n9543), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9132), .ZN(
        n9126) );
  OAI211_X1 U10450 ( .C1(n9398), .C2(n9545), .A(n9127), .B(n9126), .ZN(
        P1_U3263) );
  NAND2_X1 U10451 ( .A1(n9401), .A2(n9128), .ZN(n9129) );
  NAND2_X1 U10452 ( .A1(n9129), .A2(n9551), .ZN(n9130) );
  AOI21_X1 U10453 ( .B1(n9543), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9132), .ZN(
        n9134) );
  NAND2_X1 U10454 ( .A1(n9401), .A2(n9296), .ZN(n9133) );
  OAI211_X1 U10455 ( .C1(n9331), .C2(n9272), .A(n9134), .B(n9133), .ZN(
        P1_U3264) );
  NAND2_X1 U10456 ( .A1(n9542), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9137) );
  INV_X1 U10457 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9136) );
  OAI22_X1 U10458 ( .A1(n9138), .A2(n9137), .B1(n9136), .B2(n9322), .ZN(n9139)
         );
  AOI21_X1 U10459 ( .B1(n9140), .B2(n9296), .A(n9139), .ZN(n9141) );
  OAI21_X1 U10460 ( .B1(n9142), .B2(n9272), .A(n9141), .ZN(n9143) );
  AOI21_X1 U10461 ( .B1(n9135), .B2(n9531), .A(n9143), .ZN(n9144) );
  OAI21_X1 U10462 ( .B1(n9543), .B2(n9145), .A(n9144), .ZN(P1_U3356) );
  NAND2_X1 U10463 ( .A1(n9171), .A2(n9146), .ZN(n9147) );
  NAND2_X1 U10464 ( .A1(n9147), .A2(n9156), .ZN(n9152) );
  NAND3_X1 U10465 ( .A1(n9152), .A2(n9151), .A3(n9541), .ZN(n9154) );
  INV_X1 U10466 ( .A(n9156), .ZN(n9157) );
  NAND2_X1 U10467 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  INV_X1 U10468 ( .A(n9336), .ZN(n9168) );
  AOI21_X1 U10469 ( .B1(n9404), .B2(n9177), .A(n9620), .ZN(n9163) );
  NAND2_X1 U10470 ( .A1(n9163), .A2(n9162), .ZN(n9334) );
  AOI22_X1 U10471 ( .A1(n9164), .A2(n9542), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9268), .ZN(n9166) );
  NAND2_X1 U10472 ( .A1(n9404), .A2(n9296), .ZN(n9165) );
  OAI211_X1 U10473 ( .C1(n9334), .C2(n9272), .A(n9166), .B(n9165), .ZN(n9167)
         );
  AOI21_X1 U10474 ( .B1(n9168), .B2(n9531), .A(n9167), .ZN(n9169) );
  OAI21_X1 U10475 ( .B1(n9543), .B2(n9335), .A(n9169), .ZN(P1_U3265) );
  XNOR2_X1 U10476 ( .A(n9170), .B(n9173), .ZN(n9339) );
  INV_X1 U10477 ( .A(n9339), .ZN(n9185) );
  INV_X1 U10478 ( .A(n9174), .ZN(n9175) );
  NAND2_X1 U10479 ( .A1(n9176), .A2(n9175), .ZN(n9337) );
  AOI211_X1 U10480 ( .C1(n9178), .C2(n9192), .A(n9620), .B(n9161), .ZN(n9338)
         );
  NAND2_X1 U10481 ( .A1(n9338), .A2(n9554), .ZN(n9182) );
  INV_X1 U10482 ( .A(n9179), .ZN(n9180) );
  AOI22_X1 U10483 ( .A1(n9180), .A2(n9542), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9268), .ZN(n9181) );
  OAI211_X1 U10484 ( .C1(n9409), .C2(n9545), .A(n9182), .B(n9181), .ZN(n9183)
         );
  AOI21_X1 U10485 ( .B1(n9322), .B2(n9337), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10486 ( .B1(n9325), .B2(n9185), .A(n9184), .ZN(P1_U3266) );
  XNOR2_X1 U10487 ( .A(n9187), .B(n9186), .ZN(n9189) );
  AOI21_X1 U10488 ( .B1(n9189), .B2(n9541), .A(n9188), .ZN(n9343) );
  XNOR2_X1 U10489 ( .A(n9191), .B(n9190), .ZN(n9344) );
  INV_X1 U10490 ( .A(n9344), .ZN(n9197) );
  OAI211_X1 U10491 ( .C1(n9413), .C2(n9209), .A(n9551), .B(n9192), .ZN(n9342)
         );
  NOR2_X1 U10492 ( .A1(n9342), .A2(n9272), .ZN(n9196) );
  AOI22_X1 U10493 ( .A1(n9193), .A2(n9542), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9268), .ZN(n9194) );
  OAI21_X1 U10494 ( .B1(n9413), .B2(n9545), .A(n9194), .ZN(n9195) );
  AOI211_X1 U10495 ( .C1(n9197), .C2(n9531), .A(n9196), .B(n9195), .ZN(n9198)
         );
  OAI21_X1 U10496 ( .B1(n9543), .B2(n9343), .A(n9198), .ZN(P1_U3267) );
  XNOR2_X1 U10497 ( .A(n9199), .B(n9203), .ZN(n9351) );
  NAND2_X1 U10498 ( .A1(n9351), .A2(n9531), .ZN(n9213) );
  INV_X1 U10499 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9200) );
  OAI22_X1 U10500 ( .A1(n9201), .A2(n9294), .B1(n9200), .B2(n9322), .ZN(n9202)
         );
  AOI21_X1 U10501 ( .B1(n9348), .B2(n9296), .A(n9202), .ZN(n9212) );
  XOR2_X1 U10502 ( .A(n9204), .B(n9203), .Z(n9206) );
  OAI21_X1 U10503 ( .B1(n9206), .B2(n9506), .A(n9205), .ZN(n9349) );
  NAND2_X1 U10504 ( .A1(n9349), .A2(n9322), .ZN(n9211) );
  NAND2_X1 U10505 ( .A1(n9348), .A2(n9216), .ZN(n9207) );
  NAND2_X1 U10506 ( .A1(n9207), .A2(n9551), .ZN(n9208) );
  NOR2_X1 U10507 ( .A1(n9209), .A2(n9208), .ZN(n9350) );
  NAND2_X1 U10508 ( .A1(n9350), .A2(n9554), .ZN(n9210) );
  NAND4_X1 U10509 ( .A1(n9213), .A2(n9212), .A3(n9211), .A4(n9210), .ZN(
        P1_U3268) );
  XNOR2_X1 U10510 ( .A(n9214), .B(n9220), .ZN(n9358) );
  INV_X1 U10511 ( .A(n9215), .ZN(n9236) );
  INV_X1 U10512 ( .A(n9216), .ZN(n9217) );
  AOI21_X1 U10513 ( .B1(n9354), .B2(n9236), .A(n9217), .ZN(n9355) );
  AOI22_X1 U10514 ( .A1(n9218), .A2(n9542), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9268), .ZN(n9219) );
  OAI21_X1 U10515 ( .B1(n4767), .B2(n9545), .A(n9219), .ZN(n9227) );
  AOI21_X1 U10516 ( .B1(n9221), .B2(n9220), .A(n9506), .ZN(n9225) );
  INV_X1 U10517 ( .A(n9222), .ZN(n9223) );
  AOI21_X1 U10518 ( .B1(n9225), .B2(n9224), .A(n9223), .ZN(n9357) );
  NOR2_X1 U10519 ( .A1(n9357), .A2(n9543), .ZN(n9226) );
  AOI211_X1 U10520 ( .C1(n9355), .C2(n9228), .A(n9227), .B(n9226), .ZN(n9229)
         );
  OAI21_X1 U10521 ( .B1(n9325), .B2(n9358), .A(n9229), .ZN(P1_U3269) );
  XOR2_X1 U10522 ( .A(n9230), .B(n9233), .Z(n9232) );
  OAI21_X1 U10523 ( .B1(n9232), .B2(n9506), .A(n9231), .ZN(n9359) );
  INV_X1 U10524 ( .A(n9359), .ZN(n9243) );
  XOR2_X1 U10525 ( .A(n9234), .B(n9233), .Z(n9361) );
  AOI21_X1 U10526 ( .B1(n9251), .B2(n9235), .A(n9620), .ZN(n9237) );
  AND2_X1 U10527 ( .A1(n9237), .A2(n9236), .ZN(n9360) );
  NAND2_X1 U10528 ( .A1(n9360), .A2(n9554), .ZN(n9240) );
  AOI22_X1 U10529 ( .A1(n9238), .A2(n9542), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9268), .ZN(n9239) );
  OAI211_X1 U10530 ( .C1(n4525), .C2(n9545), .A(n9240), .B(n9239), .ZN(n9241)
         );
  AOI21_X1 U10531 ( .B1(n9361), .B2(n9531), .A(n9241), .ZN(n9242) );
  OAI21_X1 U10532 ( .B1(n9543), .B2(n9243), .A(n9242), .ZN(P1_U3270) );
  XNOR2_X1 U10533 ( .A(n9245), .B(n9244), .ZN(n9247) );
  OAI21_X1 U10534 ( .B1(n9247), .B2(n9506), .A(n9246), .ZN(n9364) );
  INV_X1 U10535 ( .A(n9364), .ZN(n9257) );
  XNOR2_X1 U10536 ( .A(n9249), .B(n9248), .ZN(n9366) );
  OR2_X1 U10537 ( .A1(n9424), .A2(n4372), .ZN(n9250) );
  AND3_X1 U10538 ( .A1(n9251), .A2(n9250), .A3(n9551), .ZN(n9365) );
  NAND2_X1 U10539 ( .A1(n9365), .A2(n9554), .ZN(n9254) );
  AOI22_X1 U10540 ( .A1(n9252), .A2(n9542), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9268), .ZN(n9253) );
  OAI211_X1 U10541 ( .C1(n9424), .C2(n9545), .A(n9254), .B(n9253), .ZN(n9255)
         );
  AOI21_X1 U10542 ( .B1(n9366), .B2(n9531), .A(n9255), .ZN(n9256) );
  OAI21_X1 U10543 ( .B1(n9543), .B2(n9257), .A(n9256), .ZN(P1_U3271) );
  XNOR2_X1 U10544 ( .A(n9258), .B(n9261), .ZN(n9260) );
  AOI21_X1 U10545 ( .B1(n9260), .B2(n9541), .A(n9259), .ZN(n9370) );
  NAND2_X1 U10546 ( .A1(n9262), .A2(n9261), .ZN(n9263) );
  NAND2_X1 U10547 ( .A1(n9264), .A2(n9263), .ZN(n9371) );
  INV_X1 U10548 ( .A(n9371), .ZN(n9274) );
  NAND2_X1 U10549 ( .A1(n9427), .A2(n9284), .ZN(n9265) );
  NAND2_X1 U10550 ( .A1(n9265), .A2(n9551), .ZN(n9266) );
  OR2_X1 U10551 ( .A1(n4372), .A2(n9266), .ZN(n9369) );
  INV_X1 U10552 ( .A(n9267), .ZN(n9269) );
  AOI22_X1 U10553 ( .A1(n9269), .A2(n9542), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9268), .ZN(n9271) );
  NAND2_X1 U10554 ( .A1(n9427), .A2(n9296), .ZN(n9270) );
  OAI211_X1 U10555 ( .C1(n9369), .C2(n9272), .A(n9271), .B(n9270), .ZN(n9273)
         );
  AOI21_X1 U10556 ( .B1(n9274), .B2(n9531), .A(n9273), .ZN(n9275) );
  OAI21_X1 U10557 ( .B1(n9543), .B2(n9370), .A(n9275), .ZN(P1_U3272) );
  XNOR2_X1 U10558 ( .A(n9277), .B(n9276), .ZN(n9379) );
  OAI211_X1 U10559 ( .C1(n9280), .C2(n9279), .A(n9278), .B(n9541), .ZN(n9282)
         );
  NAND2_X1 U10560 ( .A1(n9282), .A2(n9281), .ZN(n9376) );
  INV_X1 U10561 ( .A(n9283), .ZN(n9302) );
  INV_X1 U10562 ( .A(n9284), .ZN(n9285) );
  AOI211_X1 U10563 ( .C1(n9377), .C2(n9302), .A(n9620), .B(n9285), .ZN(n9375)
         );
  NAND2_X1 U10564 ( .A1(n9375), .A2(n9554), .ZN(n9288) );
  AOI22_X1 U10565 ( .A1(n9543), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9286), .B2(
        n9542), .ZN(n9287) );
  OAI211_X1 U10566 ( .C1(n5612), .C2(n9545), .A(n9288), .B(n9287), .ZN(n9289)
         );
  AOI21_X1 U10567 ( .B1(n9322), .B2(n9376), .A(n9289), .ZN(n9290) );
  OAI21_X1 U10568 ( .B1(n9325), .B2(n9379), .A(n9290), .ZN(P1_U3273) );
  XOR2_X1 U10569 ( .A(n9291), .B(n9298), .Z(n9383) );
  NAND2_X1 U10570 ( .A1(n9383), .A2(n9531), .ZN(n9307) );
  NAND2_X1 U10571 ( .A1(n9543), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9292) );
  OAI21_X1 U10572 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9295) );
  AOI21_X1 U10573 ( .B1(n9380), .B2(n9296), .A(n9295), .ZN(n9306) );
  XOR2_X1 U10574 ( .A(n9298), .B(n9297), .Z(n9301) );
  INV_X1 U10575 ( .A(n9299), .ZN(n9300) );
  OAI21_X1 U10576 ( .B1(n9301), .B2(n9506), .A(n9300), .ZN(n9381) );
  NAND2_X1 U10577 ( .A1(n9381), .A2(n9322), .ZN(n9305) );
  AOI21_X1 U10578 ( .B1(n9380), .B2(n9317), .A(n9620), .ZN(n9303) );
  AND2_X1 U10579 ( .A1(n9303), .A2(n9302), .ZN(n9382) );
  NAND2_X1 U10580 ( .A1(n9382), .A2(n9554), .ZN(n9304) );
  NAND4_X1 U10581 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(
        P1_U3274) );
  XNOR2_X1 U10582 ( .A(n9308), .B(n9309), .ZN(n9388) );
  INV_X1 U10583 ( .A(n9388), .ZN(n9324) );
  INV_X1 U10584 ( .A(n9310), .ZN(n9311) );
  AOI21_X1 U10585 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9315) );
  OAI21_X1 U10586 ( .B1(n9315), .B2(n9506), .A(n9314), .ZN(n9386) );
  OR2_X1 U10587 ( .A1(n9437), .A2(n4369), .ZN(n9316) );
  AND3_X1 U10588 ( .A1(n9317), .A2(n9551), .A3(n9316), .ZN(n9387) );
  NAND2_X1 U10589 ( .A1(n9387), .A2(n9554), .ZN(n9320) );
  AOI22_X1 U10590 ( .A1(n9543), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9318), .B2(
        n9542), .ZN(n9319) );
  OAI211_X1 U10591 ( .C1(n9437), .C2(n9545), .A(n9320), .B(n9319), .ZN(n9321)
         );
  AOI21_X1 U10592 ( .B1(n9386), .B2(n9322), .A(n9321), .ZN(n9323) );
  OAI21_X1 U10593 ( .B1(n9325), .B2(n9324), .A(n9323), .ZN(P1_U3275) );
  INV_X1 U10594 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9328) );
  NOR2_X1 U10595 ( .A1(n9327), .A2(n9326), .ZN(n9396) );
  MUX2_X1 U10596 ( .A(n9328), .B(n9396), .S(n10083), .Z(n9329) );
  OAI21_X1 U10597 ( .B1(n9398), .B2(n9395), .A(n9329), .ZN(P1_U3553) );
  NAND2_X1 U10598 ( .A1(n9331), .A2(n9330), .ZN(n9399) );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9399), .S(n10083), .Z(
        n9332) );
  AOI21_X1 U10600 ( .B1(n9373), .B2(n9401), .A(n9332), .ZN(n9333) );
  INV_X1 U10601 ( .A(n9333), .ZN(P1_U3552) );
  INV_X1 U10602 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9340) );
  MUX2_X1 U10603 ( .A(n9340), .B(n9406), .S(n10083), .Z(n9341) );
  OAI211_X1 U10604 ( .C1(n9344), .C2(n9583), .A(n9343), .B(n9342), .ZN(n9345)
         );
  INV_X1 U10605 ( .A(n9345), .ZN(n9410) );
  MUX2_X1 U10606 ( .A(n9346), .B(n9410), .S(n10083), .Z(n9347) );
  OAI21_X1 U10607 ( .B1(n9413), .B2(n9395), .A(n9347), .ZN(P1_U3548) );
  INV_X1 U10608 ( .A(n9348), .ZN(n9416) );
  INV_X1 U10609 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9352) );
  AOI211_X1 U10610 ( .C1(n9635), .C2(n9351), .A(n9350), .B(n9349), .ZN(n9414)
         );
  MUX2_X1 U10611 ( .A(n9352), .B(n9414), .S(n10083), .Z(n9353) );
  OAI21_X1 U10612 ( .B1(n9416), .B2(n9395), .A(n9353), .ZN(P1_U3547) );
  AOI22_X1 U10613 ( .A1(n9355), .A2(n9551), .B1(n9641), .B2(n9354), .ZN(n9356)
         );
  OAI211_X1 U10614 ( .C1(n9358), .C2(n9583), .A(n9357), .B(n9356), .ZN(n9417)
         );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9417), .S(n10083), .Z(
        P1_U3546) );
  AOI211_X1 U10616 ( .C1(n9361), .C2(n9635), .A(n9360), .B(n9359), .ZN(n9418)
         );
  MUX2_X1 U10617 ( .A(n9362), .B(n9418), .S(n10083), .Z(n9363) );
  OAI21_X1 U10618 ( .B1(n4525), .B2(n9395), .A(n9363), .ZN(P1_U3545) );
  AOI211_X1 U10619 ( .C1(n9366), .C2(n9635), .A(n9365), .B(n9364), .ZN(n9421)
         );
  MUX2_X1 U10620 ( .A(n9367), .B(n9421), .S(n10083), .Z(n9368) );
  OAI21_X1 U10621 ( .B1(n9424), .B2(n9395), .A(n9368), .ZN(P1_U3544) );
  OAI211_X1 U10622 ( .C1(n9371), .C2(n9583), .A(n9370), .B(n9369), .ZN(n9425)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9425), .S(n10083), .Z(
        n9372) );
  AOI21_X1 U10624 ( .B1(n9373), .B2(n9427), .A(n9372), .ZN(n9374) );
  INV_X1 U10625 ( .A(n9374), .ZN(P1_U3543) );
  AOI211_X1 U10626 ( .C1(n9641), .C2(n9377), .A(n9376), .B(n9375), .ZN(n9378)
         );
  OAI21_X1 U10627 ( .B1(n9583), .B2(n9379), .A(n9378), .ZN(n9430) );
  MUX2_X1 U10628 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9430), .S(n10083), .Z(
        P1_U3542) );
  INV_X1 U10629 ( .A(n9380), .ZN(n9433) );
  INV_X1 U10630 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9384) );
  AOI211_X1 U10631 ( .C1(n9383), .C2(n9635), .A(n9382), .B(n9381), .ZN(n9431)
         );
  MUX2_X1 U10632 ( .A(n9384), .B(n9431), .S(n10083), .Z(n9385) );
  OAI21_X1 U10633 ( .B1(n9433), .B2(n9395), .A(n9385), .ZN(P1_U3541) );
  AOI211_X1 U10634 ( .C1(n9388), .C2(n9635), .A(n9387), .B(n9386), .ZN(n9434)
         );
  MUX2_X1 U10635 ( .A(n9389), .B(n9434), .S(n10083), .Z(n9390) );
  OAI21_X1 U10636 ( .B1(n9437), .B2(n9395), .A(n9390), .ZN(P1_U3540) );
  AOI211_X1 U10637 ( .C1(n9393), .C2(n9635), .A(n9392), .B(n9391), .ZN(n9438)
         );
  MUX2_X1 U10638 ( .A(n9076), .B(n9438), .S(n10083), .Z(n9394) );
  OAI21_X1 U10639 ( .B1(n4542), .B2(n9395), .A(n9394), .ZN(P1_U3539) );
  INV_X1 U10640 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U10641 ( .A(n10061), .B(n9396), .S(n9650), .Z(n9397) );
  OAI21_X1 U10642 ( .B1(n9398), .B2(n5626), .A(n9397), .ZN(P1_U3521) );
  MUX2_X1 U10643 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9399), .S(n9650), .Z(n9400) );
  AOI21_X1 U10644 ( .B1(n9428), .B2(n9401), .A(n9400), .ZN(n9402) );
  INV_X1 U10645 ( .A(n9402), .ZN(P1_U3520) );
  INV_X1 U10646 ( .A(n9405), .ZN(P1_U3518) );
  MUX2_X1 U10647 ( .A(n9407), .B(n9406), .S(n9650), .Z(n9408) );
  OAI21_X1 U10648 ( .B1(n9409), .B2(n5626), .A(n9408), .ZN(P1_U3517) );
  INV_X1 U10649 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U10650 ( .A(n9411), .B(n9410), .S(n9650), .Z(n9412) );
  OAI21_X1 U10651 ( .B1(n9413), .B2(n5626), .A(n9412), .ZN(P1_U3516) );
  MUX2_X1 U10652 ( .A(n10053), .B(n9414), .S(n9650), .Z(n9415) );
  OAI21_X1 U10653 ( .B1(n9416), .B2(n5626), .A(n9415), .ZN(P1_U3515) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9417), .S(n9650), .Z(
        P1_U3514) );
  INV_X1 U10655 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9419) );
  MUX2_X1 U10656 ( .A(n9419), .B(n9418), .S(n9650), .Z(n9420) );
  OAI21_X1 U10657 ( .B1(n4525), .B2(n5626), .A(n9420), .ZN(P1_U3513) );
  INV_X1 U10658 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9422) );
  MUX2_X1 U10659 ( .A(n9422), .B(n9421), .S(n9650), .Z(n9423) );
  OAI21_X1 U10660 ( .B1(n9424), .B2(n5626), .A(n9423), .ZN(P1_U3512) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9425), .S(n9650), .Z(n9426) );
  AOI21_X1 U10662 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9429) );
  INV_X1 U10663 ( .A(n9429), .ZN(P1_U3511) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9430), .S(n9650), .Z(
        P1_U3510) );
  INV_X1 U10665 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U10666 ( .A(n10002), .B(n9431), .S(n9650), .Z(n9432) );
  OAI21_X1 U10667 ( .B1(n9433), .B2(n5626), .A(n9432), .ZN(P1_U3509) );
  INV_X1 U10668 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9435) );
  MUX2_X1 U10669 ( .A(n9435), .B(n9434), .S(n9650), .Z(n9436) );
  OAI21_X1 U10670 ( .B1(n9437), .B2(n5626), .A(n9436), .ZN(P1_U3507) );
  INV_X1 U10671 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9439) );
  MUX2_X1 U10672 ( .A(n9439), .B(n9438), .S(n9650), .Z(n9440) );
  OAI21_X1 U10673 ( .B1(n4542), .B2(n5626), .A(n9440), .ZN(P1_U3504) );
  MUX2_X1 U10674 ( .A(P1_D_REG_1__SCAN_IN), .B(n9443), .S(n9558), .Z(P1_U3440)
         );
  MUX2_X1 U10675 ( .A(P1_D_REG_0__SCAN_IN), .B(n9444), .S(n9558), .Z(P1_U3439)
         );
  NOR4_X1 U10676 ( .A1(n9445), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5176), .A4(
        P1_U3086), .ZN(n9446) );
  AOI21_X1 U10677 ( .B1(n9447), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9446), .ZN(
        n9448) );
  OAI21_X1 U10678 ( .B1(n9449), .B2(n9452), .A(n9448), .ZN(P1_U3324) );
  MUX2_X1 U10679 ( .A(n9453), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NAND3_X1 U10680 ( .A1(n4319), .A2(n9454), .A3(n9635), .ZN(n9456) );
  OAI211_X1 U10681 ( .C1(n9457), .C2(n9632), .A(n9456), .B(n9455), .ZN(n9459)
         );
  NOR2_X1 U10682 ( .A1(n9459), .A2(n9458), .ZN(n9462) );
  AOI22_X1 U10683 ( .A1(n10083), .A2(n9462), .B1(n9460), .B2(n9670), .ZN(
        P1_U3538) );
  INV_X1 U10684 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9461) );
  AOI22_X1 U10685 ( .A1(n9650), .A2(n9462), .B1(n9461), .B2(n9648), .ZN(
        P1_U3501) );
  XNOR2_X1 U10686 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10687 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10688 ( .A(n9463), .ZN(n9469) );
  NAND2_X1 U10689 ( .A1(n4294), .A2(n9479), .ZN(n9467) );
  NAND2_X1 U10690 ( .A1(n9465), .A2(n9467), .ZN(n9466) );
  MUX2_X1 U10691 ( .A(n9467), .B(n9466), .S(P1_IR_REG_0__SCAN_IN), .Z(n9468)
         );
  NAND2_X1 U10692 ( .A1(n9469), .A2(n9468), .ZN(n9471) );
  AOI22_X1 U10693 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9490), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9470) );
  OAI21_X1 U10694 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(P1_U3243) );
  AOI22_X1 U10695 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9490), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9485) );
  AOI211_X1 U10696 ( .C1(n9475), .C2(n9474), .A(n9473), .B(n9486), .ZN(n9476)
         );
  AOI21_X1 U10697 ( .B1(n9478), .B2(n9477), .A(n9476), .ZN(n9484) );
  NOR2_X1 U10698 ( .A1(n4726), .A2(n9479), .ZN(n9482) );
  OAI211_X1 U10699 ( .C1(n9482), .C2(n9481), .A(n9492), .B(n9480), .ZN(n9483)
         );
  NAND3_X1 U10700 ( .A1(n9485), .A2(n9484), .A3(n9483), .ZN(P1_U3244) );
  AOI211_X1 U10701 ( .C1(n9489), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9500)
         );
  AOI22_X1 U10702 ( .A1(n9490), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9496) );
  OAI211_X1 U10703 ( .C1(n9494), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9495)
         );
  OAI211_X1 U10704 ( .C1(n9498), .C2(n9497), .A(n9496), .B(n9495), .ZN(n9499)
         );
  OR3_X1 U10705 ( .A1(n9501), .A2(n9500), .A3(n9499), .ZN(P1_U3245) );
  INV_X1 U10706 ( .A(n9537), .ZN(n9647) );
  XNOR2_X1 U10707 ( .A(n9502), .B(n9504), .ZN(n9597) );
  AOI21_X1 U10708 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9507) );
  NOR2_X1 U10709 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  AOI211_X1 U10710 ( .C1(n9647), .C2(n9597), .A(n9509), .B(n9508), .ZN(n9594)
         );
  AOI22_X1 U10711 ( .A1(n9543), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9510), .B2(
        n9542), .ZN(n9511) );
  OAI21_X1 U10712 ( .B1(n9545), .B2(n9593), .A(n9511), .ZN(n9512) );
  INV_X1 U10713 ( .A(n9512), .ZN(n9518) );
  NOR2_X1 U10714 ( .A1(n9543), .A2(n9513), .ZN(n9555) );
  OAI211_X1 U10715 ( .C1(n9515), .C2(n9593), .A(n9551), .B(n9514), .ZN(n9592)
         );
  INV_X1 U10716 ( .A(n9592), .ZN(n9516) );
  AOI22_X1 U10717 ( .A1(n9597), .A2(n9555), .B1(n9554), .B2(n9516), .ZN(n9517)
         );
  OAI211_X1 U10718 ( .C1(n9543), .C2(n9594), .A(n9518), .B(n9517), .ZN(
        P1_U3286) );
  NAND2_X1 U10719 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  XNOR2_X1 U10720 ( .A(n9521), .B(n9528), .ZN(n9523) );
  AOI21_X1 U10721 ( .B1(n9523), .B2(n9541), .A(n9522), .ZN(n9574) );
  AOI22_X1 U10722 ( .A1(n9543), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9542), .B2(
        n9524), .ZN(n9525) );
  OAI21_X1 U10723 ( .B1(n9545), .B2(n9573), .A(n9525), .ZN(n9526) );
  INV_X1 U10724 ( .A(n9526), .ZN(n9533) );
  XNOR2_X1 U10725 ( .A(n9528), .B(n9527), .ZN(n9577) );
  OAI211_X1 U10726 ( .C1(n7567), .C2(n9573), .A(n9529), .B(n9551), .ZN(n9572)
         );
  INV_X1 U10727 ( .A(n9572), .ZN(n9530) );
  AOI22_X1 U10728 ( .A1(n9577), .A2(n9531), .B1(n9554), .B2(n9530), .ZN(n9532)
         );
  OAI211_X1 U10729 ( .C1(n9543), .C2(n9574), .A(n9533), .B(n9532), .ZN(
        P1_U3290) );
  OAI21_X1 U10730 ( .B1(n9535), .B2(n6194), .A(n9534), .ZN(n9540) );
  XOR2_X1 U10731 ( .A(n9536), .B(n6194), .Z(n9547) );
  NOR2_X1 U10732 ( .A1(n9547), .A2(n9537), .ZN(n9538) );
  AOI211_X1 U10733 ( .C1(n9541), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9562)
         );
  AOI22_X1 U10734 ( .A1(n9543), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9542), .ZN(n9544) );
  OAI21_X1 U10735 ( .B1(n9545), .B2(n9561), .A(n9544), .ZN(n9546) );
  INV_X1 U10736 ( .A(n9546), .ZN(n9557) );
  INV_X1 U10737 ( .A(n9547), .ZN(n9565) );
  NAND2_X1 U10738 ( .A1(n9549), .A2(n9548), .ZN(n9550) );
  NAND3_X1 U10739 ( .A1(n9552), .A2(n9551), .A3(n9550), .ZN(n9560) );
  INV_X1 U10740 ( .A(n9560), .ZN(n9553) );
  AOI22_X1 U10741 ( .A1(n9565), .A2(n9555), .B1(n9554), .B2(n9553), .ZN(n9556)
         );
  OAI211_X1 U10742 ( .C1(n9543), .C2(n9562), .A(n9557), .B(n9556), .ZN(
        P1_U3292) );
  INV_X1 U10743 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U10744 ( .A1(n9558), .A2(n10026), .ZN(P1_U3294) );
  AND2_X1 U10745 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9559), .ZN(P1_U3295) );
  AND2_X1 U10746 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9559), .ZN(P1_U3296) );
  AND2_X1 U10747 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9559), .ZN(P1_U3297) );
  AND2_X1 U10748 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9559), .ZN(P1_U3298) );
  AND2_X1 U10749 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9559), .ZN(P1_U3299) );
  AND2_X1 U10750 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9559), .ZN(P1_U3300) );
  AND2_X1 U10751 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9559), .ZN(P1_U3301) );
  AND2_X1 U10752 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9559), .ZN(P1_U3302) );
  AND2_X1 U10753 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9559), .ZN(P1_U3303) );
  AND2_X1 U10754 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9559), .ZN(P1_U3304) );
  AND2_X1 U10755 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9559), .ZN(P1_U3305) );
  INV_X1 U10756 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U10757 ( .A1(n9558), .A2(n10062), .ZN(P1_U3306) );
  INV_X1 U10758 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U10759 ( .A1(n9558), .A2(n10046), .ZN(P1_U3307) );
  AND2_X1 U10760 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9559), .ZN(P1_U3308) );
  AND2_X1 U10761 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9559), .ZN(P1_U3309) );
  AND2_X1 U10762 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9559), .ZN(P1_U3310) );
  AND2_X1 U10763 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9559), .ZN(P1_U3311) );
  AND2_X1 U10764 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9559), .ZN(P1_U3312) );
  AND2_X1 U10765 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9559), .ZN(P1_U3313) );
  AND2_X1 U10766 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9559), .ZN(P1_U3314) );
  AND2_X1 U10767 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9559), .ZN(P1_U3315) );
  AND2_X1 U10768 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9559), .ZN(P1_U3316) );
  AND2_X1 U10769 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9559), .ZN(P1_U3317) );
  AND2_X1 U10770 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9559), .ZN(P1_U3318) );
  AND2_X1 U10771 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9559), .ZN(P1_U3319) );
  AND2_X1 U10772 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9559), .ZN(P1_U3320) );
  AND2_X1 U10773 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9559), .ZN(P1_U3321) );
  AND2_X1 U10774 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9559), .ZN(P1_U3322) );
  AND2_X1 U10775 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9559), .ZN(P1_U3323) );
  INV_X1 U10776 ( .A(n9644), .ZN(n9598) );
  OAI21_X1 U10777 ( .B1(n9561), .B2(n9632), .A(n9560), .ZN(n9564) );
  INV_X1 U10778 ( .A(n9562), .ZN(n9563) );
  AOI211_X1 U10779 ( .C1(n9598), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9652)
         );
  INV_X1 U10780 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U10781 ( .A1(n9650), .A2(n9652), .B1(n9566), .B2(n9648), .ZN(
        P1_U3456) );
  OAI21_X1 U10782 ( .B1(n5151), .B2(n9632), .A(n9567), .ZN(n9569) );
  AOI211_X1 U10783 ( .C1(n9635), .C2(n9570), .A(n9569), .B(n9568), .ZN(n9654)
         );
  INV_X1 U10784 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9571) );
  AOI22_X1 U10785 ( .A1(n9650), .A2(n9654), .B1(n9571), .B2(n9648), .ZN(
        P1_U3459) );
  OAI21_X1 U10786 ( .B1(n9573), .B2(n9632), .A(n9572), .ZN(n9576) );
  INV_X1 U10787 ( .A(n9574), .ZN(n9575) );
  AOI211_X1 U10788 ( .C1(n9635), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9656)
         );
  INV_X1 U10789 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9578) );
  AOI22_X1 U10790 ( .A1(n9650), .A2(n9656), .B1(n9578), .B2(n9648), .ZN(
        P1_U3462) );
  AOI21_X1 U10791 ( .B1(n9641), .B2(n9580), .A(n9579), .ZN(n9582) );
  OAI211_X1 U10792 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9585)
         );
  INV_X1 U10793 ( .A(n9585), .ZN(n9658) );
  INV_X1 U10794 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U10795 ( .A1(n9650), .A2(n9658), .B1(n9586), .B2(n9648), .ZN(
        P1_U3465) );
  OAI211_X1 U10796 ( .C1(n9589), .C2(n9632), .A(n9588), .B(n9587), .ZN(n9590)
         );
  AOI21_X1 U10797 ( .B1(n9635), .B2(n9591), .A(n9590), .ZN(n9659) );
  INV_X1 U10798 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U10799 ( .A1(n9650), .A2(n9659), .B1(n10004), .B2(n9648), .ZN(
        P1_U3471) );
  OAI21_X1 U10800 ( .B1(n9593), .B2(n9632), .A(n9592), .ZN(n9596) );
  INV_X1 U10801 ( .A(n9594), .ZN(n9595) );
  AOI211_X1 U10802 ( .C1(n9598), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9660)
         );
  INV_X1 U10803 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U10804 ( .A1(n9650), .A2(n9660), .B1(n9599), .B2(n9648), .ZN(
        P1_U3474) );
  AND2_X1 U10805 ( .A1(n9600), .A2(n9635), .ZN(n9604) );
  OAI21_X1 U10806 ( .B1(n9602), .B2(n9632), .A(n9601), .ZN(n9603) );
  NOR3_X1 U10807 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n9661) );
  INV_X1 U10808 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9606) );
  AOI22_X1 U10809 ( .A1(n9650), .A2(n9661), .B1(n9606), .B2(n9648), .ZN(
        P1_U3477) );
  AND2_X1 U10810 ( .A1(n9607), .A2(n9635), .ZN(n9611) );
  AND2_X1 U10811 ( .A1(n9608), .A2(n9641), .ZN(n9610) );
  NOR4_X1 U10812 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9663)
         );
  INV_X1 U10813 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9613) );
  AOI22_X1 U10814 ( .A1(n9650), .A2(n9663), .B1(n9613), .B2(n9648), .ZN(
        P1_U3480) );
  OAI211_X1 U10815 ( .C1(n9616), .C2(n9632), .A(n9615), .B(n9614), .ZN(n9617)
         );
  AOI21_X1 U10816 ( .B1(n9635), .B2(n9618), .A(n9617), .ZN(n9664) );
  INV_X1 U10817 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9619) );
  AOI22_X1 U10818 ( .A1(n9650), .A2(n9664), .B1(n9619), .B2(n9648), .ZN(
        P1_U3483) );
  OAI22_X1 U10819 ( .A1(n9621), .A2(n9620), .B1(n4596), .B2(n9632), .ZN(n9623)
         );
  AOI211_X1 U10820 ( .C1(n9624), .C2(n9635), .A(n9623), .B(n9622), .ZN(n9665)
         );
  INV_X1 U10821 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U10822 ( .A1(n9650), .A2(n9665), .B1(n9972), .B2(n9648), .ZN(
        P1_U3486) );
  OAI21_X1 U10823 ( .B1(n9626), .B2(n9632), .A(n9625), .ZN(n9628) );
  AOI211_X1 U10824 ( .C1(n9629), .C2(n9635), .A(n9628), .B(n9627), .ZN(n9667)
         );
  INV_X1 U10825 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U10826 ( .A1(n9650), .A2(n9667), .B1(n9955), .B2(n9648), .ZN(
        P1_U3489) );
  OAI211_X1 U10827 ( .C1(n9633), .C2(n9632), .A(n9631), .B(n9630), .ZN(n9634)
         );
  AOI21_X1 U10828 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9669) );
  INV_X1 U10829 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9637) );
  AOI22_X1 U10830 ( .A1(n9650), .A2(n9669), .B1(n9637), .B2(n9648), .ZN(
        P1_U3492) );
  INV_X1 U10831 ( .A(n9643), .ZN(n9646) );
  AOI211_X1 U10832 ( .C1(n9641), .C2(n9640), .A(n9639), .B(n9638), .ZN(n9642)
         );
  OAI21_X1 U10833 ( .B1(n9644), .B2(n9643), .A(n9642), .ZN(n9645) );
  AOI21_X1 U10834 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9671) );
  INV_X1 U10835 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9649) );
  AOI22_X1 U10836 ( .A1(n9650), .A2(n9671), .B1(n9649), .B2(n9648), .ZN(
        P1_U3495) );
  AOI22_X1 U10837 ( .A1(n10083), .A2(n9652), .B1(n9651), .B2(n9670), .ZN(
        P1_U3523) );
  AOI22_X1 U10838 ( .A1(n10083), .A2(n9654), .B1(n9653), .B2(n9670), .ZN(
        P1_U3524) );
  AOI22_X1 U10839 ( .A1(n10083), .A2(n9656), .B1(n9655), .B2(n9670), .ZN(
        P1_U3525) );
  AOI22_X1 U10840 ( .A1(n10083), .A2(n9658), .B1(n9657), .B2(n9670), .ZN(
        P1_U3526) );
  AOI22_X1 U10841 ( .A1(n10083), .A2(n9659), .B1(n6784), .B2(n9670), .ZN(
        P1_U3528) );
  AOI22_X1 U10842 ( .A1(n10083), .A2(n9660), .B1(n6831), .B2(n9670), .ZN(
        P1_U3529) );
  AOI22_X1 U10843 ( .A1(n10083), .A2(n9661), .B1(n6909), .B2(n9670), .ZN(
        P1_U3530) );
  AOI22_X1 U10844 ( .A1(n10083), .A2(n9663), .B1(n9662), .B2(n9670), .ZN(
        P1_U3531) );
  AOI22_X1 U10845 ( .A1(n10083), .A2(n9664), .B1(n7079), .B2(n9670), .ZN(
        P1_U3532) );
  AOI22_X1 U10846 ( .A1(n10083), .A2(n9665), .B1(n10050), .B2(n9670), .ZN(
        P1_U3533) );
  AOI22_X1 U10847 ( .A1(n10083), .A2(n9667), .B1(n9666), .B2(n9670), .ZN(
        P1_U3534) );
  AOI22_X1 U10848 ( .A1(n10083), .A2(n9669), .B1(n9668), .B2(n9670), .ZN(
        P1_U3535) );
  AOI22_X1 U10849 ( .A1(n10083), .A2(n9671), .B1(n7674), .B2(n9670), .ZN(
        P1_U3536) );
  INV_X1 U10850 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U10851 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  NAND2_X1 U10852 ( .A1(n9675), .A2(n9674), .ZN(n9681) );
  NAND2_X1 U10853 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  NAND2_X1 U10854 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  AOI22_X1 U10855 ( .A1(n9768), .A2(n9681), .B1(n9758), .B2(n9680), .ZN(n9684)
         );
  NAND2_X1 U10856 ( .A1(n9809), .A2(n9682), .ZN(n9683) );
  OAI211_X1 U10857 ( .C1(n9737), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9686)
         );
  INV_X1 U10858 ( .A(n9686), .ZN(n9691) );
  XNOR2_X1 U10859 ( .A(n9688), .B(n9687), .ZN(n9689) );
  NAND2_X1 U10860 ( .A1(n9689), .A2(n9822), .ZN(n9690) );
  OAI211_X1 U10861 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7158), .A(n9691), .B(
        n9690), .ZN(P2_U3183) );
  INV_X1 U10862 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9835) );
  INV_X1 U10863 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9703) );
  OAI21_X1 U10864 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9699) );
  OAI21_X1 U10865 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9698) );
  AOI22_X1 U10866 ( .A1(n9768), .A2(n9699), .B1(n9758), .B2(n9698), .ZN(n9702)
         );
  NAND2_X1 U10867 ( .A1(n9809), .A2(n9700), .ZN(n9701) );
  OAI211_X1 U10868 ( .C1(n9737), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9704)
         );
  INV_X1 U10869 ( .A(n9704), .ZN(n9709) );
  XOR2_X1 U10870 ( .A(n9705), .B(n9706), .Z(n9707) );
  NAND2_X1 U10871 ( .A1(n9707), .A2(n9822), .ZN(n9708) );
  OAI211_X1 U10872 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9835), .A(n9709), .B(
        n9708), .ZN(P2_U3184) );
  AND2_X1 U10873 ( .A1(n9809), .A2(n9710), .ZN(n9715) );
  INV_X1 U10874 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9713) );
  INV_X1 U10875 ( .A(n9711), .ZN(n9712) );
  OAI22_X1 U10876 ( .A1(n9737), .A2(n9713), .B1(n9826), .B2(n9712), .ZN(n9714)
         );
  NOR2_X1 U10877 ( .A1(n9715), .A2(n9714), .ZN(n9725) );
  XOR2_X1 U10878 ( .A(n9717), .B(n9716), .Z(n9718) );
  NAND2_X1 U10879 ( .A1(n9718), .A2(n9822), .ZN(n9723) );
  OAI21_X1 U10880 ( .B1(n9720), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9719), .ZN(
        n9721) );
  NAND2_X1 U10881 ( .A1(n9768), .A2(n9721), .ZN(n9722) );
  NAND4_X1 U10882 ( .A1(n9725), .A2(n9724), .A3(n9723), .A4(n9722), .ZN(
        P2_U3187) );
  INV_X1 U10883 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U10884 ( .A1(n9809), .A2(n9726), .ZN(n9735) );
  INV_X1 U10885 ( .A(n9727), .ZN(n9729) );
  NAND3_X1 U10886 ( .A1(n9730), .A2(n9729), .A3(n9728), .ZN(n9731) );
  NAND2_X1 U10887 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U10888 ( .A1(n9758), .A2(n9733), .ZN(n9734) );
  OAI211_X1 U10889 ( .C1(n9737), .C2(n9736), .A(n9735), .B(n9734), .ZN(n9738)
         );
  INV_X1 U10890 ( .A(n9738), .ZN(n9750) );
  AOI21_X1 U10891 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  OR2_X1 U10892 ( .A1(n9742), .A2(n9763), .ZN(n9748) );
  OAI21_X1 U10893 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  NAND2_X1 U10894 ( .A1(n9768), .A2(n9746), .ZN(n9747) );
  NAND4_X1 U10895 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(
        P2_U3188) );
  INV_X1 U10896 ( .A(n9751), .ZN(n9753) );
  NAND3_X1 U10897 ( .A1(n9754), .A2(n9753), .A3(n9752), .ZN(n9755) );
  NAND2_X1 U10898 ( .A1(n9756), .A2(n9755), .ZN(n9759) );
  AOI222_X1 U10899 ( .A1(n9759), .A2(n9758), .B1(n9808), .B2(
        P2_ADDR_REG_8__SCAN_IN), .C1(n9757), .C2(n9809), .ZN(n9773) );
  AOI21_X1 U10900 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9764) );
  OR2_X1 U10901 ( .A1(n9764), .A2(n9763), .ZN(n9771) );
  OAI21_X1 U10902 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9769) );
  NAND2_X1 U10903 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  NAND4_X1 U10904 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(
        P2_U3190) );
  AOI22_X1 U10905 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9808), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n9789) );
  AOI21_X1 U10906 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9786) );
  AOI21_X1 U10907 ( .B1(n4374), .B2(n9778), .A(n9777), .ZN(n9779) );
  OR2_X1 U10908 ( .A1(n9779), .A2(n9817), .ZN(n9785) );
  OAI21_X1 U10909 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9783) );
  NAND2_X1 U10910 ( .A1(n9783), .A2(n9822), .ZN(n9784) );
  OAI211_X1 U10911 ( .C1(n9786), .C2(n9826), .A(n9785), .B(n9784), .ZN(n9787)
         );
  INV_X1 U10912 ( .A(n9787), .ZN(n9788) );
  OAI211_X1 U10913 ( .C1(n9807), .C2(n9790), .A(n9789), .B(n9788), .ZN(
        P2_U3196) );
  AOI22_X1 U10914 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9808), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3151), .ZN(n9805) );
  AOI21_X1 U10915 ( .B1(n4337), .B2(n9792), .A(n9791), .ZN(n9802) );
  AOI21_X1 U10916 ( .B1(n4338), .B2(n9794), .A(n9793), .ZN(n9795) );
  OR2_X1 U10917 ( .A1(n9795), .A2(n9817), .ZN(n9801) );
  OAI21_X1 U10918 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9799) );
  NAND2_X1 U10919 ( .A1(n9799), .A2(n9822), .ZN(n9800) );
  OAI211_X1 U10920 ( .C1(n9802), .C2(n9826), .A(n9801), .B(n9800), .ZN(n9803)
         );
  INV_X1 U10921 ( .A(n9803), .ZN(n9804) );
  OAI211_X1 U10922 ( .C1(n9807), .C2(n9806), .A(n9805), .B(n9804), .ZN(
        P2_U3198) );
  INV_X1 U10923 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U10924 ( .A1(n9810), .A2(n9809), .B1(n9808), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9830) );
  AOI21_X1 U10925 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9827) );
  AOI21_X1 U10926 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9818) );
  OR2_X1 U10927 ( .A1(n9818), .A2(n9817), .ZN(n9825) );
  OAI21_X1 U10928 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9823) );
  NAND2_X1 U10929 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  OAI211_X1 U10930 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n9824), .ZN(n9828)
         );
  INV_X1 U10931 ( .A(n9828), .ZN(n9829) );
  OAI211_X1 U10932 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9831), .A(n9830), .B(
        n9829), .ZN(P2_U3199) );
  INV_X1 U10933 ( .A(n9832), .ZN(n9847) );
  XNOR2_X1 U10934 ( .A(n9833), .B(n9838), .ZN(n9856) );
  OAI22_X1 U10935 ( .A1(n9854), .A2(n9836), .B1(n9835), .B2(n9834), .ZN(n9846)
         );
  NAND3_X1 U10936 ( .A1(n9838), .A2(n9837), .A3(n7136), .ZN(n9839) );
  NAND2_X1 U10937 ( .A1(n7213), .A2(n9839), .ZN(n9843) );
  AOI222_X1 U10938 ( .A1(n9844), .A2(n9843), .B1(n9842), .B2(n9841), .C1(n4293), .C2(n9840), .ZN(n9853) );
  INV_X1 U10939 ( .A(n9853), .ZN(n9845) );
  AOI211_X1 U10940 ( .C1(n9847), .C2(n9856), .A(n9846), .B(n9845), .ZN(n9850)
         );
  AOI22_X1 U10941 ( .A1(n9856), .A2(n9848), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n8586), .ZN(n9849) );
  OAI21_X1 U10942 ( .B1(n8586), .B2(n9850), .A(n9849), .ZN(P2_U3231) );
  INV_X1 U10943 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9852) );
  AOI22_X1 U10944 ( .A1(n9893), .A2(n9852), .B1(n9851), .B2(n9891), .ZN(
        P2_U3393) );
  INV_X1 U10945 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10065) );
  OAI21_X1 U10946 ( .B1(n9854), .B2(n9873), .A(n9853), .ZN(n9855) );
  AOI21_X1 U10947 ( .B1(n9856), .B2(n9865), .A(n9855), .ZN(n9894) );
  AOI22_X1 U10948 ( .A1(n9893), .A2(n10065), .B1(n9894), .B2(n9891), .ZN(
        P2_U3396) );
  INV_X1 U10949 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U10950 ( .A1(n9858), .A2(n9865), .B1(n9890), .B2(n9857), .ZN(n9859)
         );
  AND2_X1 U10951 ( .A1(n9860), .A2(n9859), .ZN(n9896) );
  AOI22_X1 U10952 ( .A1(n9893), .A2(n9861), .B1(n9896), .B2(n9891), .ZN(
        P2_U3399) );
  INV_X1 U10953 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9867) );
  OAI21_X1 U10954 ( .B1(n9863), .B2(n9873), .A(n9862), .ZN(n9864) );
  AOI21_X1 U10955 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9897) );
  AOI22_X1 U10956 ( .A1(n9893), .A2(n9867), .B1(n9897), .B2(n9891), .ZN(
        P2_U3402) );
  INV_X1 U10957 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9872) );
  OAI22_X1 U10958 ( .A1(n9869), .A2(n9885), .B1(n9868), .B2(n9873), .ZN(n9870)
         );
  NOR2_X1 U10959 ( .A1(n9871), .A2(n9870), .ZN(n9899) );
  AOI22_X1 U10960 ( .A1(n9893), .A2(n9872), .B1(n9899), .B2(n9891), .ZN(
        P2_U3405) );
  INV_X1 U10961 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9878) );
  OAI22_X1 U10962 ( .A1(n9875), .A2(n9885), .B1(n9874), .B2(n9873), .ZN(n9876)
         );
  NOR2_X1 U10963 ( .A1(n9877), .A2(n9876), .ZN(n9900) );
  AOI22_X1 U10964 ( .A1(n9893), .A2(n9878), .B1(n9900), .B2(n9891), .ZN(
        P2_U3411) );
  INV_X1 U10965 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9884) );
  NOR2_X1 U10966 ( .A1(n9880), .A2(n9879), .ZN(n9882) );
  AOI211_X1 U10967 ( .C1(n9890), .C2(n9883), .A(n9882), .B(n9881), .ZN(n9901)
         );
  AOI22_X1 U10968 ( .A1(n9893), .A2(n9884), .B1(n9901), .B2(n9891), .ZN(
        P2_U3414) );
  INV_X1 U10969 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9892) );
  NOR2_X1 U10970 ( .A1(n9886), .A2(n9885), .ZN(n9888) );
  AOI211_X1 U10971 ( .C1(n9890), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9903)
         );
  AOI22_X1 U10972 ( .A1(n9893), .A2(n9892), .B1(n9903), .B2(n9891), .ZN(
        P2_U3417) );
  AOI22_X1 U10973 ( .A1(n9904), .A2(n9894), .B1(n5697), .B2(n9902), .ZN(
        P2_U3461) );
  AOI22_X1 U10974 ( .A1(n9904), .A2(n9896), .B1(n9895), .B2(n9902), .ZN(
        P2_U3462) );
  AOI22_X1 U10975 ( .A1(n9904), .A2(n9897), .B1(n5707), .B2(n9902), .ZN(
        P2_U3463) );
  INV_X1 U10976 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U10977 ( .A1(n9904), .A2(n9899), .B1(n9898), .B2(n9902), .ZN(
        P2_U3464) );
  INV_X1 U10978 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U10979 ( .A1(n9904), .A2(n9900), .B1(n9973), .B2(n9902), .ZN(
        P2_U3466) );
  AOI22_X1 U10980 ( .A1(n9904), .A2(n9901), .B1(n9987), .B2(n9902), .ZN(
        P2_U3467) );
  AOI22_X1 U10981 ( .A1(n9904), .A2(n9903), .B1(n4475), .B2(n9902), .ZN(
        P2_U3468) );
  NOR2_X1 U10982 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  XOR2_X1 U10983 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9907), .Z(ADD_1068_U5) );
  XOR2_X1 U10984 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10985 ( .A1(n9909), .A2(n9908), .ZN(n9910) );
  XOR2_X1 U10986 ( .A(n9910), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55) );
  XNOR2_X1 U10987 ( .A(n9912), .B(n9911), .ZN(ADD_1068_U56) );
  XNOR2_X1 U10988 ( .A(n9914), .B(n9913), .ZN(ADD_1068_U57) );
  XNOR2_X1 U10989 ( .A(n9916), .B(n9915), .ZN(ADD_1068_U58) );
  XNOR2_X1 U10990 ( .A(n9918), .B(n9917), .ZN(ADD_1068_U59) );
  XNOR2_X1 U10991 ( .A(n9920), .B(n9919), .ZN(ADD_1068_U60) );
  XNOR2_X1 U10992 ( .A(n9922), .B(n9921), .ZN(ADD_1068_U61) );
  XNOR2_X1 U10993 ( .A(n9924), .B(n9923), .ZN(ADD_1068_U62) );
  XNOR2_X1 U10994 ( .A(n9926), .B(n9925), .ZN(ADD_1068_U63) );
  NAND2_X1 U10995 ( .A1(keyinput47), .A2(keyinput63), .ZN(n9932) );
  NOR2_X1 U10996 ( .A1(keyinput8), .A2(keyinput59), .ZN(n9930) );
  NAND3_X1 U10997 ( .A1(keyinput34), .A2(keyinput22), .A3(keyinput52), .ZN(
        n9928) );
  NAND3_X1 U10998 ( .A1(keyinput25), .A2(keyinput16), .A3(keyinput54), .ZN(
        n9927) );
  NOR4_X1 U10999 ( .A1(keyinput39), .A2(keyinput44), .A3(n9928), .A4(n9927), 
        .ZN(n9929) );
  NAND4_X1 U11000 ( .A1(keyinput42), .A2(keyinput40), .A3(n9930), .A4(n9929), 
        .ZN(n9931) );
  NOR4_X1 U11001 ( .A1(keyinput32), .A2(keyinput4), .A3(n9932), .A4(n9931), 
        .ZN(n10080) );
  NOR3_X1 U11002 ( .A1(keyinput14), .A2(keyinput57), .A3(keyinput46), .ZN(
        n9938) );
  INV_X1 U11003 ( .A(keyinput38), .ZN(n9933) );
  NOR4_X1 U11004 ( .A1(keyinput13), .A2(keyinput45), .A3(keyinput23), .A4(
        n9933), .ZN(n9937) );
  NAND4_X1 U11005 ( .A1(keyinput11), .A2(keyinput50), .A3(keyinput24), .A4(
        keyinput10), .ZN(n9935) );
  NAND2_X1 U11006 ( .A1(keyinput60), .A2(keyinput37), .ZN(n9934) );
  NOR4_X1 U11007 ( .A1(keyinput7), .A2(keyinput36), .A3(n9935), .A4(n9934), 
        .ZN(n9936) );
  NAND4_X1 U11008 ( .A1(keyinput1), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(
        n9953) );
  NOR2_X1 U11009 ( .A1(keyinput27), .A2(keyinput19), .ZN(n9944) );
  NAND2_X1 U11010 ( .A1(keyinput58), .A2(keyinput31), .ZN(n9942) );
  NOR3_X1 U11011 ( .A1(keyinput5), .A2(keyinput20), .A3(keyinput9), .ZN(n9940)
         );
  NOR3_X1 U11012 ( .A1(keyinput2), .A2(keyinput48), .A3(keyinput53), .ZN(n9939) );
  NAND4_X1 U11013 ( .A1(keyinput15), .A2(n9940), .A3(keyinput43), .A4(n9939), 
        .ZN(n9941) );
  NOR4_X1 U11014 ( .A1(keyinput12), .A2(keyinput29), .A3(n9942), .A4(n9941), 
        .ZN(n9943) );
  NAND4_X1 U11015 ( .A1(keyinput17), .A2(keyinput49), .A3(n9944), .A4(n9943), 
        .ZN(n9952) );
  NOR2_X1 U11016 ( .A1(keyinput28), .A2(keyinput56), .ZN(n9947) );
  INV_X1 U11017 ( .A(keyinput33), .ZN(n9945) );
  NOR4_X1 U11018 ( .A1(keyinput55), .A2(keyinput30), .A3(keyinput62), .A4(
        n9945), .ZN(n9946) );
  NAND4_X1 U11019 ( .A1(keyinput3), .A2(keyinput0), .A3(n9947), .A4(n9946), 
        .ZN(n9951) );
  NOR2_X1 U11020 ( .A1(keyinput51), .A2(keyinput35), .ZN(n9949) );
  NOR4_X1 U11021 ( .A1(keyinput41), .A2(keyinput6), .A3(keyinput21), .A4(
        keyinput18), .ZN(n9948) );
  NAND4_X1 U11022 ( .A1(keyinput26), .A2(keyinput61), .A3(n9949), .A4(n9948), 
        .ZN(n9950) );
  NOR4_X1 U11023 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n10079)
         );
  AOI22_X1 U11024 ( .A1(n9956), .A2(keyinput1), .B1(keyinput46), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11025 ( .B1(n9956), .B2(keyinput1), .C1(n9955), .C2(keyinput46), 
        .A(n9954), .ZN(n9968) );
  INV_X1 U11026 ( .A(keyinput14), .ZN(n9958) );
  AOI22_X1 U11027 ( .A1(n9959), .A2(keyinput57), .B1(P1_ADDR_REG_2__SCAN_IN), 
        .B2(n9958), .ZN(n9957) );
  OAI221_X1 U11028 ( .B1(n9959), .B2(keyinput57), .C1(n9958), .C2(
        P1_ADDR_REG_2__SCAN_IN), .A(n9957), .ZN(n9967) );
  AOI22_X1 U11029 ( .A1(n9962), .A2(keyinput11), .B1(keyinput50), .B2(n9961), 
        .ZN(n9960) );
  OAI221_X1 U11030 ( .B1(n9962), .B2(keyinput11), .C1(n9961), .C2(keyinput50), 
        .A(n9960), .ZN(n9966) );
  XNOR2_X1 U11031 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput24), .ZN(n9964) );
  XNOR2_X1 U11032 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput10), .ZN(n9963) );
  NAND2_X1 U11033 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  NOR4_X1 U11034 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n10016)
         );
  AOI22_X1 U11035 ( .A1(n9971), .A2(keyinput7), .B1(n9970), .B2(keyinput37), 
        .ZN(n9969) );
  OAI221_X1 U11036 ( .B1(n9971), .B2(keyinput7), .C1(n9970), .C2(keyinput37), 
        .A(n9969), .ZN(n9981) );
  XNOR2_X1 U11037 ( .A(keyinput60), .B(n9972), .ZN(n9980) );
  XNOR2_X1 U11038 ( .A(keyinput13), .B(n9973), .ZN(n9979) );
  XNOR2_X1 U11039 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput38), .ZN(n9977) );
  XNOR2_X1 U11040 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput36), .ZN(n9976) );
  XNOR2_X1 U11041 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput45), .ZN(n9975) );
  XNOR2_X1 U11042 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput23), .ZN(n9974) );
  NAND4_X1 U11043 ( .A1(n9977), .A2(n9976), .A3(n9975), .A4(n9974), .ZN(n9978)
         );
  NOR4_X1 U11044 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n10015)
         );
  AOI22_X1 U11045 ( .A1(n9984), .A2(keyinput5), .B1(n9983), .B2(keyinput15), 
        .ZN(n9982) );
  OAI221_X1 U11046 ( .B1(n9984), .B2(keyinput5), .C1(n9983), .C2(keyinput15), 
        .A(n9982), .ZN(n9996) );
  AOI22_X1 U11047 ( .A1(n9987), .A2(keyinput20), .B1(n9986), .B2(keyinput9), 
        .ZN(n9985) );
  OAI221_X1 U11048 ( .B1(n9987), .B2(keyinput20), .C1(n9986), .C2(keyinput9), 
        .A(n9985), .ZN(n9995) );
  INV_X1 U11049 ( .A(SI_13_), .ZN(n9989) );
  AOI22_X1 U11050 ( .A1(n9989), .A2(keyinput2), .B1(keyinput43), .B2(n8650), 
        .ZN(n9988) );
  OAI221_X1 U11051 ( .B1(n9989), .B2(keyinput2), .C1(n8650), .C2(keyinput43), 
        .A(n9988), .ZN(n9994) );
  AOI22_X1 U11052 ( .A1(n9992), .A2(keyinput48), .B1(n9991), .B2(keyinput53), 
        .ZN(n9990) );
  OAI221_X1 U11053 ( .B1(n9992), .B2(keyinput48), .C1(n9991), .C2(keyinput53), 
        .A(n9990), .ZN(n9993) );
  NOR4_X1 U11054 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n10014)
         );
  AOI22_X1 U11055 ( .A1(n9999), .A2(keyinput27), .B1(n9998), .B2(keyinput17), 
        .ZN(n9997) );
  OAI221_X1 U11056 ( .B1(n9999), .B2(keyinput27), .C1(n9998), .C2(keyinput17), 
        .A(n9997), .ZN(n10012) );
  INV_X1 U11057 ( .A(SI_21_), .ZN(n10001) );
  AOI22_X1 U11058 ( .A1(n10002), .A2(keyinput49), .B1(n10001), .B2(keyinput19), 
        .ZN(n10000) );
  OAI221_X1 U11059 ( .B1(n10002), .B2(keyinput49), .C1(n10001), .C2(keyinput19), .A(n10000), .ZN(n10011) );
  AOI22_X1 U11060 ( .A1(n10005), .A2(keyinput58), .B1(keyinput12), .B2(n10004), 
        .ZN(n10003) );
  OAI221_X1 U11061 ( .B1(n10005), .B2(keyinput58), .C1(n10004), .C2(keyinput12), .A(n10003), .ZN(n10010) );
  AOI22_X1 U11062 ( .A1(n10008), .A2(keyinput31), .B1(keyinput29), .B2(n10007), 
        .ZN(n10006) );
  OAI221_X1 U11063 ( .B1(n10008), .B2(keyinput31), .C1(n10007), .C2(keyinput29), .A(n10006), .ZN(n10009) );
  NOR4_X1 U11064 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10013) );
  NAND4_X1 U11065 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10078) );
  INV_X1 U11066 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10019) );
  AOI22_X1 U11067 ( .A1(n10019), .A2(keyinput8), .B1(n10018), .B2(keyinput59), 
        .ZN(n10017) );
  OAI221_X1 U11068 ( .B1(n10019), .B2(keyinput8), .C1(n10018), .C2(keyinput59), 
        .A(n10017), .ZN(n10031) );
  AOI22_X1 U11069 ( .A1(n10021), .A2(keyinput42), .B1(keyinput40), .B2(n7674), 
        .ZN(n10020) );
  OAI221_X1 U11070 ( .B1(n10021), .B2(keyinput42), .C1(n7674), .C2(keyinput40), 
        .A(n10020), .ZN(n10030) );
  AOI22_X1 U11071 ( .A1(n10024), .A2(keyinput54), .B1(n10023), .B2(keyinput44), 
        .ZN(n10022) );
  OAI221_X1 U11072 ( .B1(n10024), .B2(keyinput54), .C1(n10023), .C2(keyinput44), .A(n10022), .ZN(n10029) );
  AOI22_X1 U11073 ( .A1(n10027), .A2(keyinput25), .B1(keyinput16), .B2(n10026), 
        .ZN(n10025) );
  OAI221_X1 U11074 ( .B1(n10027), .B2(keyinput25), .C1(n10026), .C2(keyinput16), .A(n10025), .ZN(n10028) );
  NOR4_X1 U11075 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10076) );
  AOI22_X1 U11076 ( .A1(n10034), .A2(keyinput47), .B1(n10033), .B2(keyinput32), 
        .ZN(n10032) );
  OAI221_X1 U11077 ( .B1(n10034), .B2(keyinput47), .C1(n10033), .C2(keyinput32), .A(n10032), .ZN(n10044) );
  AOI22_X1 U11078 ( .A1(n10037), .A2(keyinput4), .B1(n10036), .B2(keyinput63), 
        .ZN(n10035) );
  OAI221_X1 U11079 ( .B1(n10037), .B2(keyinput4), .C1(n10036), .C2(keyinput63), 
        .A(n10035), .ZN(n10043) );
  XNOR2_X1 U11080 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput52), .ZN(n10041)
         );
  XNOR2_X1 U11081 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput22), .ZN(n10040) );
  XNOR2_X1 U11082 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput34), .ZN(n10039)
         );
  XNOR2_X1 U11083 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput39), .ZN(n10038) );
  NAND4_X1 U11084 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10042) );
  NOR3_X1 U11085 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10075) );
  AOI22_X1 U11086 ( .A1(n10047), .A2(keyinput0), .B1(keyinput56), .B2(n10046), 
        .ZN(n10045) );
  OAI221_X1 U11087 ( .B1(n10047), .B2(keyinput0), .C1(n10046), .C2(keyinput56), 
        .A(n10045), .ZN(n10059) );
  AOI22_X1 U11088 ( .A1(n10050), .A2(keyinput3), .B1(n10049), .B2(keyinput28), 
        .ZN(n10048) );
  OAI221_X1 U11089 ( .B1(n10050), .B2(keyinput3), .C1(n10049), .C2(keyinput28), 
        .A(n10048), .ZN(n10058) );
  INV_X1 U11090 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U11091 ( .A1(n10053), .A2(keyinput33), .B1(n10052), .B2(keyinput30), 
        .ZN(n10051) );
  OAI221_X1 U11092 ( .B1(n10053), .B2(keyinput33), .C1(n10052), .C2(keyinput30), .A(n10051), .ZN(n10057) );
  XNOR2_X1 U11093 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput62), .ZN(n10055)
         );
  XNOR2_X1 U11094 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput55), .ZN(n10054)
         );
  NAND2_X1 U11095 ( .A1(n10055), .A2(n10054), .ZN(n10056) );
  NOR4_X1 U11096 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10074) );
  AOI22_X1 U11097 ( .A1(n10062), .A2(keyinput35), .B1(keyinput61), .B2(n10061), 
        .ZN(n10060) );
  OAI221_X1 U11098 ( .B1(n10062), .B2(keyinput35), .C1(n10061), .C2(keyinput61), .A(n10060), .ZN(n10072) );
  AOI22_X1 U11099 ( .A1(n10065), .A2(keyinput26), .B1(keyinput51), .B2(n10064), 
        .ZN(n10063) );
  OAI221_X1 U11100 ( .B1(n10065), .B2(keyinput26), .C1(n10064), .C2(keyinput51), .A(n10063), .ZN(n10071) );
  XNOR2_X1 U11101 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput18), .ZN(n10069) );
  XNOR2_X1 U11102 ( .A(P2_REG1_REG_29__SCAN_IN), .B(keyinput21), .ZN(n10068)
         );
  XNOR2_X1 U11103 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput41), .ZN(n10067) );
  XNOR2_X1 U11104 ( .A(P1_REG0_REG_27__SCAN_IN), .B(keyinput6), .ZN(n10066) );
  NAND4_X1 U11105 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10070) );
  NOR3_X1 U11106 ( .A1(n10072), .A2(n10071), .A3(n10070), .ZN(n10073) );
  NAND4_X1 U11107 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10077) );
  AOI211_X1 U11108 ( .C1(n10080), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10085) );
  NAND2_X1 U11109 ( .A1(n10081), .A2(n10083), .ZN(n10082) );
  OAI21_X1 U11110 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10083), .A(n10082), .ZN(
        n10084) );
  XNOR2_X1 U11111 ( .A(n10085), .B(n10084), .ZN(P1_U3527) );
  XNOR2_X1 U11112 ( .A(n10087), .B(n10086), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11113 ( .A(n10089), .B(n10088), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11114 ( .A(n10091), .B(n10090), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11115 ( .A(n10093), .B(n10092), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11116 ( .A(n10095), .B(n10094), .ZN(ADD_1068_U48) );
  XOR2_X1 U11117 ( .A(n10097), .B(n10096), .Z(ADD_1068_U54) );
  XOR2_X1 U11118 ( .A(n10099), .B(n10098), .Z(ADD_1068_U53) );
  XNOR2_X1 U11119 ( .A(n10101), .B(n10100), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4844 ( .A(n5128), .Z(n4291) );
endmodule

